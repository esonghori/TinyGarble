
module hamming_N16000_CC8_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  XOR U19 ( .A(A[13]), .B(n19), .Z(SUM[13]) );
  ANDN U20 ( .B(A[12]), .A(n20), .Z(n19) );
  XNOR U21 ( .A(A[12]), .B(n20), .Z(SUM[12]) );
  NANDN U22 ( .A(n21), .B(A[11]), .Z(n20) );
  XNOR U23 ( .A(A[11]), .B(n21), .Z(SUM[11]) );
  AND U24 ( .A(n22), .B(n23), .Z(n21) );
  NAND U25 ( .A(n24), .B(B[10]), .Z(n23) );
  NANDN U26 ( .A(A[10]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(n25), .B(A[10]), .Z(n22) );
  XOR U28 ( .A(n25), .B(n26), .Z(SUM[10]) );
  XNOR U29 ( .A(B[10]), .B(A[10]), .Z(n26) );
  AND U30 ( .A(n27), .B(n28), .Z(n25) );
  NAND U31 ( .A(n29), .B(B[9]), .Z(n28) );
  NANDN U32 ( .A(A[9]), .B(n1), .Z(n29) );
  NANDN U33 ( .A(n1), .B(A[9]), .Z(n27) );
  AND U34 ( .A(n30), .B(n31), .Z(n1) );
  NAND U35 ( .A(n32), .B(B[8]), .Z(n31) );
  NANDN U36 ( .A(A[8]), .B(n3), .Z(n32) );
  NANDN U37 ( .A(n3), .B(A[8]), .Z(n30) );
  AND U38 ( .A(n33), .B(n34), .Z(n3) );
  NAND U39 ( .A(n35), .B(B[7]), .Z(n34) );
  NANDN U40 ( .A(A[7]), .B(n5), .Z(n35) );
  NANDN U41 ( .A(n5), .B(A[7]), .Z(n33) );
  AND U42 ( .A(n36), .B(n37), .Z(n5) );
  NAND U43 ( .A(n38), .B(B[6]), .Z(n37) );
  NANDN U44 ( .A(A[6]), .B(n7), .Z(n38) );
  NANDN U45 ( .A(n7), .B(A[6]), .Z(n36) );
  AND U46 ( .A(n39), .B(n40), .Z(n7) );
  NAND U47 ( .A(n41), .B(B[5]), .Z(n40) );
  NANDN U48 ( .A(A[5]), .B(n9), .Z(n41) );
  NANDN U49 ( .A(n9), .B(A[5]), .Z(n39) );
  AND U50 ( .A(n42), .B(n43), .Z(n9) );
  NAND U51 ( .A(n44), .B(B[4]), .Z(n43) );
  NANDN U52 ( .A(A[4]), .B(n11), .Z(n44) );
  NANDN U53 ( .A(n11), .B(A[4]), .Z(n42) );
  AND U54 ( .A(n45), .B(n46), .Z(n11) );
  NAND U55 ( .A(n47), .B(B[3]), .Z(n46) );
  NANDN U56 ( .A(A[3]), .B(n13), .Z(n47) );
  NANDN U57 ( .A(n13), .B(A[3]), .Z(n45) );
  AND U58 ( .A(n48), .B(n49), .Z(n13) );
  NAND U59 ( .A(n50), .B(B[2]), .Z(n49) );
  NANDN U60 ( .A(A[2]), .B(n15), .Z(n50) );
  NANDN U61 ( .A(n15), .B(A[2]), .Z(n48) );
  AND U62 ( .A(n51), .B(n52), .Z(n15) );
  NAND U63 ( .A(n53), .B(B[1]), .Z(n52) );
  OR U64 ( .A(n17), .B(A[1]), .Z(n53) );
  NAND U65 ( .A(n17), .B(A[1]), .Z(n51) );
  AND U66 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U67 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_1 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  IV U1 ( .A(B[10]), .Z(n1) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  XOR U20 ( .A(n20), .B(n1), .Z(SUM[10]) );
  AND U21 ( .A(n21), .B(n22), .Z(n20) );
  NAND U22 ( .A(n23), .B(B[9]), .Z(n22) );
  NANDN U23 ( .A(A[9]), .B(n2), .Z(n23) );
  NANDN U24 ( .A(n2), .B(A[9]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n2) );
  NAND U26 ( .A(n26), .B(B[8]), .Z(n25) );
  NANDN U27 ( .A(A[8]), .B(n4), .Z(n26) );
  NANDN U28 ( .A(n4), .B(A[8]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n4) );
  NAND U30 ( .A(n29), .B(B[7]), .Z(n28) );
  NANDN U31 ( .A(A[7]), .B(n6), .Z(n29) );
  NANDN U32 ( .A(n6), .B(A[7]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n6) );
  NAND U34 ( .A(n32), .B(B[6]), .Z(n31) );
  NANDN U35 ( .A(A[6]), .B(n8), .Z(n32) );
  NANDN U36 ( .A(n8), .B(A[6]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n8) );
  NAND U38 ( .A(n35), .B(B[5]), .Z(n34) );
  NANDN U39 ( .A(A[5]), .B(n10), .Z(n35) );
  NANDN U40 ( .A(n10), .B(A[5]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n10) );
  NAND U42 ( .A(n38), .B(B[4]), .Z(n37) );
  NANDN U43 ( .A(A[4]), .B(n12), .Z(n38) );
  NANDN U44 ( .A(n12), .B(A[4]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n12) );
  NAND U46 ( .A(n41), .B(B[3]), .Z(n40) );
  NANDN U47 ( .A(A[3]), .B(n14), .Z(n41) );
  NANDN U48 ( .A(n14), .B(A[3]), .Z(n39) );
  AND U49 ( .A(n42), .B(n43), .Z(n14) );
  NAND U50 ( .A(n44), .B(B[2]), .Z(n43) );
  NANDN U51 ( .A(A[2]), .B(n16), .Z(n44) );
  NANDN U52 ( .A(n16), .B(A[2]), .Z(n42) );
  AND U53 ( .A(n45), .B(n46), .Z(n16) );
  NAND U54 ( .A(n47), .B(B[1]), .Z(n46) );
  OR U55 ( .A(n18), .B(A[1]), .Z(n47) );
  NAND U56 ( .A(n18), .B(A[1]), .Z(n45) );
  AND U57 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U58 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_2 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(n22), .B(B[9]), .Z(n21) );
  NANDN U21 ( .A(A[9]), .B(n2), .Z(n22) );
  NANDN U22 ( .A(n2), .B(A[9]), .Z(n20) );
  AND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(n25), .B(B[8]), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(n28), .B(B[7]), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(n31), .B(B[6]), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(n34), .B(B[5]), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(n37), .B(B[4]), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(n40), .B(B[3]), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(n43), .B(B[2]), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(n46), .B(B[1]), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(n18), .B(A[1]), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_3 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_4 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n18), .B(n19), .Z(SUM[9]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[8]) );
  XNOR U3 ( .A(B[8]), .B(A[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[7]) );
  XNOR U5 ( .A(B[7]), .B(A[7]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U7 ( .A(B[6]), .B(A[6]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U9 ( .A(B[5]), .B(A[5]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U11 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[3]) );
  XNOR U13 ( .A(B[3]), .B(A[3]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[2]) );
  XNOR U15 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[1]) );
  XOR U17 ( .A(B[1]), .B(A[1]), .Z(n17) );
  NAND U18 ( .A(n20), .B(B[8]), .Z(n19) );
  NANDN U19 ( .A(A[8]), .B(n2), .Z(n20) );
  NANDN U20 ( .A(n2), .B(A[8]), .Z(n18) );
  AND U21 ( .A(n21), .B(n22), .Z(n2) );
  NAND U22 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U23 ( .A(A[7]), .B(n4), .Z(n23) );
  NANDN U24 ( .A(n4), .B(A[7]), .Z(n21) );
  AND U25 ( .A(n24), .B(n25), .Z(n4) );
  NAND U26 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U27 ( .A(A[6]), .B(n6), .Z(n26) );
  NANDN U28 ( .A(n6), .B(A[6]), .Z(n24) );
  AND U29 ( .A(n27), .B(n28), .Z(n6) );
  NAND U30 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U31 ( .A(A[5]), .B(n8), .Z(n29) );
  NANDN U32 ( .A(n8), .B(A[5]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n8) );
  NAND U34 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U35 ( .A(A[4]), .B(n10), .Z(n32) );
  NANDN U36 ( .A(n10), .B(A[4]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(n10) );
  NAND U38 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U39 ( .A(A[3]), .B(n12), .Z(n35) );
  NANDN U40 ( .A(n12), .B(A[3]), .Z(n33) );
  AND U41 ( .A(n36), .B(n37), .Z(n12) );
  NAND U42 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U43 ( .A(A[2]), .B(n14), .Z(n38) );
  NANDN U44 ( .A(n14), .B(A[2]), .Z(n36) );
  AND U45 ( .A(n39), .B(n40), .Z(n14) );
  NAND U46 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U47 ( .A(n16), .B(A[1]), .Z(n41) );
  NAND U48 ( .A(n16), .B(A[1]), .Z(n39) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n16) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_5 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39;

  AND U1 ( .A(n2), .B(B[8]), .Z(SUM[9]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[8]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[8]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  AND U19 ( .A(n19), .B(n20), .Z(n4) );
  NAND U20 ( .A(n21), .B(B[7]), .Z(n20) );
  NANDN U21 ( .A(A[7]), .B(n5), .Z(n21) );
  NANDN U22 ( .A(n5), .B(A[7]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n5) );
  NAND U24 ( .A(n24), .B(B[6]), .Z(n23) );
  NANDN U25 ( .A(A[6]), .B(n7), .Z(n24) );
  NANDN U26 ( .A(n7), .B(A[6]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n7) );
  NAND U28 ( .A(n27), .B(B[5]), .Z(n26) );
  NANDN U29 ( .A(A[5]), .B(n9), .Z(n27) );
  NANDN U30 ( .A(n9), .B(A[5]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n9) );
  NAND U32 ( .A(n30), .B(B[4]), .Z(n29) );
  NANDN U33 ( .A(A[4]), .B(n11), .Z(n30) );
  NANDN U34 ( .A(n11), .B(A[4]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n11) );
  NAND U36 ( .A(n33), .B(B[3]), .Z(n32) );
  NANDN U37 ( .A(A[3]), .B(n13), .Z(n33) );
  NANDN U38 ( .A(n13), .B(A[3]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n13) );
  NAND U40 ( .A(n36), .B(B[2]), .Z(n35) );
  NANDN U41 ( .A(A[2]), .B(n15), .Z(n36) );
  NANDN U42 ( .A(n15), .B(A[2]), .Z(n34) );
  AND U43 ( .A(n37), .B(n38), .Z(n15) );
  NAND U44 ( .A(n39), .B(B[1]), .Z(n38) );
  OR U45 ( .A(n17), .B(A[1]), .Z(n39) );
  NAND U46 ( .A(n17), .B(A[1]), .Z(n37) );
  AND U47 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U48 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_6 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_7 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_8 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_9 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(n18), .B(B[7]), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(n21), .B(B[6]), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(n24), .B(B[5]), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(n27), .B(B[4]), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(n33), .B(B[2]), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(n36), .B(B[1]), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(n14), .B(A[1]), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_10 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34;

  AND U1 ( .A(n2), .B(B[7]), .Z(SUM[8]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[7]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  AND U17 ( .A(n17), .B(n18), .Z(n4) );
  NAND U18 ( .A(n19), .B(B[6]), .Z(n18) );
  NANDN U19 ( .A(A[6]), .B(n5), .Z(n19) );
  NANDN U20 ( .A(n5), .B(A[6]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n5) );
  NAND U22 ( .A(n22), .B(B[5]), .Z(n21) );
  NANDN U23 ( .A(A[5]), .B(n7), .Z(n22) );
  NANDN U24 ( .A(n7), .B(A[5]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n7) );
  NAND U26 ( .A(n25), .B(B[4]), .Z(n24) );
  NANDN U27 ( .A(A[4]), .B(n9), .Z(n25) );
  NANDN U28 ( .A(n9), .B(A[4]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n9) );
  NAND U30 ( .A(n28), .B(B[3]), .Z(n27) );
  NANDN U31 ( .A(A[3]), .B(n11), .Z(n28) );
  NANDN U32 ( .A(n11), .B(A[3]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n11) );
  NAND U34 ( .A(n31), .B(B[2]), .Z(n30) );
  NANDN U35 ( .A(A[2]), .B(n13), .Z(n31) );
  NANDN U36 ( .A(n13), .B(A[2]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n13) );
  NAND U38 ( .A(n34), .B(B[1]), .Z(n33) );
  OR U39 ( .A(n15), .B(A[1]), .Z(n34) );
  NAND U40 ( .A(n15), .B(A[1]), .Z(n32) );
  AND U41 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U42 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_11 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_12 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_13 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_14 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_15 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_16 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_17 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_18 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_19 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_20 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(n16), .B(B[6]), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(n22), .B(B[4]), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(n25), .B(B[3]), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(n28), .B(B[2]), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(n31), .B(B[1]), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(n12), .B(A[1]), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_21 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_22 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_23 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_24 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_25 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_26 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_27 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_28 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_29 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_30 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_31 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_32 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_33 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_34 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_35 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_36 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_37 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_38 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_39 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_40 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_41 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(n23), .B(B[2]), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(n26), .B(B[1]), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(n10), .B(A[1]), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_42 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_43 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_44 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_45 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_46 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_47 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_48 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_49 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_50 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_51 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_52 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_53 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_54 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_55 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_56 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_57 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_58 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_59 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_60 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_61 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_62 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_63 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_64 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_65 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_66 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_67 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_68 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_69 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_70 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_71 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_72 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_73 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_74 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_75 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_76 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_77 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_78 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_79 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_80 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_81 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_82 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(n15), .B(B[3]), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(n18), .B(B[2]), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(n21), .B(B[1]), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(n8), .B(A[1]), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8_DW01_add_83 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;

  AND U1 ( .A(n2), .B(B[4]), .Z(SUM[5]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[4]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[3]) );
  XNOR U6 ( .A(B[3]), .B(A[3]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[2]) );
  XNOR U8 ( .A(B[2]), .B(A[2]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[1]) );
  XOR U10 ( .A(B[1]), .B(A[1]), .Z(n10) );
  AND U11 ( .A(n11), .B(n12), .Z(n4) );
  NAND U12 ( .A(n13), .B(B[3]), .Z(n12) );
  NANDN U13 ( .A(A[3]), .B(n5), .Z(n13) );
  NANDN U14 ( .A(n5), .B(A[3]), .Z(n11) );
  AND U15 ( .A(n14), .B(n15), .Z(n5) );
  NAND U16 ( .A(n16), .B(B[2]), .Z(n15) );
  NANDN U17 ( .A(A[2]), .B(n7), .Z(n16) );
  NANDN U18 ( .A(n7), .B(A[2]), .Z(n14) );
  AND U19 ( .A(n17), .B(n18), .Z(n7) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n9), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n9), .B(A[1]), .Z(n17) );
  AND U23 ( .A(B[0]), .B(A[0]), .Z(n9) );
  XOR U24 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC8 ( clk, rst, x, y, o );
  input [1999:0] x;
  input [1999:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N12770, N12771, N12772, N12773, N12781, N12782, N12783, N12784,
         N12785, N12792, N12793, N12794, N12795, N12796, N12803, N12804,
         N12805, N12806, N12807, N12814, N12815, N12816, N12817, N12818,
         N12825, N12826, N12827, N12828, N12829, N12836, N12837, N12838,
         N12839, N12840, N12847, N12848, N12849, N12850, N12851, N12858,
         N12859, N12860, N12861, N12862, N12869, N12870, N12871, N12872,
         N12873, N12880, N12881, N12882, N12883, N12884, N12891, N12892,
         N12893, N12894, N12895, N12902, N12903, N12904, N12905, N12906,
         N12913, N12914, N12915, N12916, N12917, N12924, N12925, N12926,
         N12927, N12928, N12935, N12936, N12937, N12938, N12939, N12946,
         N12947, N12948, N12949, N12950, N12957, N12958, N12959, N12960,
         N12961, N12968, N12969, N12970, N12971, N12972, N12979, N12980,
         N12981, N12982, N12983, N12990, N12991, N12992, N12993, N12994,
         N13001, N13002, N13003, N13004, N13005, N13012, N13013, N13014,
         N13015, N13016, N13023, N13024, N13025, N13026, N13027, N13034,
         N13035, N13036, N13037, N13038, N13045, N13046, N13047, N13048,
         N13049, N13056, N13057, N13058, N13059, N13060, N13067, N13068,
         N13069, N13070, N13071, N13078, N13079, N13080, N13081, N13082,
         N13089, N13090, N13091, N13092, N13093, N13100, N13101, N13102,
         N13103, N13104, N13111, N13112, N13113, N13114, N13115, N13122,
         N13123, N13124, N13125, N13126, N13133, N13134, N13135, N13136,
         N13137, N13144, N13145, N13146, N13147, N13148, N13155, N13156,
         N13157, N13158, N13159, N13166, N13167, N13168, N13169, N13170,
         N13177, N13178, N13179, N13180, N13181, N13188, N13189, N13190,
         N13191, N13192, N13199, N13200, N13201, N13202, N13203, N13210,
         N13211, N13212, N13213, N13214, N13221, N13222, N13223, N13224,
         N13225, N13232, N13233, N13234, N13235, N13236, N13243, N13244,
         N13245, N13246, N13247, N13254, N13255, N13256, N13257, N13258,
         N13265, N13266, N13267, N13268, N13269, N13276, N13277, N13278,
         N13279, N13280, N13287, N13288, N13289, N13290, N13291, N13298,
         N13299, N13300, N13301, N13302, N13309, N13310, N13311, N13312,
         N13313, N13320, N13321, N13322, N13323, N13324, N13331, N13332,
         N13333, N13334, N13335, N13342, N13343, N13344, N13345, N13346,
         N13353, N13354, N13355, N13356, N13357, N13364, N13365, N13366,
         N13367, N13368, N13375, N13376, N13377, N13378, N13379, N13386,
         N13387, N13388, N13389, N13390, N13397, N13398, N13399, N13400,
         N13401, N13408, N13409, N13410, N13411, N13412, N13419, N13420,
         N13421, N13422, N13423, N13430, N13431, N13432, N13433, N13434,
         N13441, N13442, N13443, N13444, N13445, N13452, N13453, N13454,
         N13455, N13456, N13463, N13464, N13465, N13466, N13467, N13474,
         N13475, N13476, N13477, N13478, N13485, N13486, N13487, N13488,
         N13489, N13496, N13497, N13498, N13499, N13500, N13507, N13508,
         N13509, N13510, N13511, N13518, N13519, N13520, N13521, N13522,
         N13529, N13530, N13531, N13532, N13533, N13540, N13541, N13542,
         N13543, N13544, N13551, N13552, N13553, N13554, N13555, N13562,
         N13563, N13564, N13565, N13566, N13573, N13574, N13575, N13576,
         N13577, N13584, N13585, N13586, N13587, N13588, N13595, N13596,
         N13597, N13598, N13599, N13606, N13607, N13608, N13609, N13610,
         N13617, N13618, N13619, N13620, N13621, N13628, N13629, N13630,
         N13631, N13632, N13639, N13640, N13641, N13642, N13643, N13650,
         N13651, N13652, N13653, N13654, N13661, N13662, N13663, N13664,
         N13665, N13672, N13673, N13674, N13675, N13676, N13683, N13684,
         N13685, N13686, N13687, N13694, N13695, N13696, N13697, N13698,
         N13699, N13705, N13706, N13707, N13708, N13709, N13710, N13716,
         N13717, N13718, N13719, N13720, N13721, N13727, N13728, N13729,
         N13730, N13731, N13732, N13738, N13739, N13740, N13741, N13742,
         N13743, N13749, N13750, N13751, N13752, N13753, N13754, N13760,
         N13761, N13762, N13763, N13764, N13765, N13771, N13772, N13773,
         N13774, N13775, N13776, N13782, N13783, N13784, N13785, N13786,
         N13787, N13793, N13794, N13795, N13796, N13797, N13798, N13804,
         N13805, N13806, N13807, N13808, N13809, N13815, N13816, N13817,
         N13818, N13819, N13820, N13826, N13827, N13828, N13829, N13830,
         N13831, N13837, N13838, N13839, N13840, N13841, N13842, N13848,
         N13849, N13850, N13851, N13852, N13853, N13859, N13860, N13861,
         N13862, N13863, N13864, N13870, N13871, N13872, N13873, N13874,
         N13875, N13881, N13882, N13883, N13884, N13885, N13886, N13892,
         N13893, N13894, N13895, N13896, N13897, N13903, N13904, N13905,
         N13906, N13907, N13908, N13914, N13915, N13916, N13917, N13918,
         N13919, N13925, N13926, N13927, N13928, N13929, N13930, N13936,
         N13937, N13938, N13939, N13940, N13941, N13947, N13948, N13949,
         N13950, N13951, N13952, N13958, N13959, N13960, N13961, N13962,
         N13963, N13969, N13970, N13971, N13972, N13973, N13974, N13980,
         N13981, N13982, N13983, N13984, N13985, N13991, N13992, N13993,
         N13994, N13995, N13996, N14002, N14003, N14004, N14005, N14006,
         N14007, N14013, N14014, N14015, N14016, N14017, N14018, N14024,
         N14025, N14026, N14027, N14028, N14029, N14035, N14036, N14037,
         N14038, N14039, N14040, N14046, N14047, N14048, N14049, N14050,
         N14051, N14057, N14058, N14059, N14060, N14061, N14062, N14068,
         N14069, N14070, N14071, N14072, N14073, N14079, N14080, N14081,
         N14082, N14083, N14084, N14090, N14091, N14092, N14093, N14094,
         N14095, N14101, N14102, N14103, N14104, N14105, N14106, N14112,
         N14113, N14114, N14115, N14116, N14117, N14123, N14124, N14125,
         N14126, N14127, N14128, N14134, N14135, N14136, N14137, N14138,
         N14139, N14145, N14146, N14147, N14148, N14149, N14150, N14156,
         N14157, N14158, N14159, N14160, N14161, N14162, N14167, N14168,
         N14169, N14170, N14171, N14172, N14173, N14178, N14179, N14180,
         N14181, N14182, N14183, N14184, N14189, N14190, N14191, N14192,
         N14193, N14194, N14195, N14200, N14201, N14202, N14203, N14204,
         N14205, N14206, N14211, N14212, N14213, N14214, N14215, N14216,
         N14217, N14222, N14223, N14224, N14225, N14226, N14227, N14228,
         N14233, N14234, N14235, N14236, N14237, N14238, N14239, N14244,
         N14245, N14246, N14247, N14248, N14249, N14250, N14255, N14256,
         N14257, N14258, N14259, N14260, N14261, N14266, N14267, N14268,
         N14269, N14270, N14271, N14272, N14277, N14278, N14279, N14280,
         N14281, N14282, N14283, N14288, N14289, N14290, N14291, N14292,
         N14293, N14294, N14299, N14300, N14301, N14302, N14303, N14304,
         N14305, N14310, N14311, N14312, N14313, N14314, N14315, N14316,
         N14321, N14322, N14323, N14324, N14325, N14326, N14327, N14332,
         N14333, N14334, N14335, N14336, N14337, N14338, N14343, N14344,
         N14345, N14346, N14347, N14348, N14349, N14354, N14355, N14356,
         N14357, N14358, N14359, N14360, N14365, N14366, N14367, N14368,
         N14369, N14370, N14371, N14376, N14377, N14378, N14379, N14380,
         N14381, N14382, N14387, N14388, N14389, N14390, N14391, N14392,
         N14393, N14394, N14398, N14399, N14400, N14401, N14402, N14403,
         N14404, N14405, N14409, N14410, N14411, N14412, N14413, N14414,
         N14415, N14416, N14420, N14421, N14422, N14423, N14424, N14425,
         N14426, N14427, N14431, N14432, N14433, N14434, N14435, N14436,
         N14437, N14438, N14442, N14443, N14444, N14445, N14446, N14447,
         N14448, N14449, N14453, N14454, N14455, N14456, N14457, N14458,
         N14459, N14460, N14464, N14465, N14466, N14467, N14468, N14469,
         N14470, N14471, N14475, N14476, N14477, N14478, N14479, N14480,
         N14481, N14482, N14486, N14487, N14488, N14489, N14490, N14491,
         N14492, N14493, N14497, N14498, N14499, N14500, N14501, N14502,
         N14503, N14504, N14505, N14508, N14509, N14510, N14511, N14512,
         N14513, N14514, N14515, N14516, N14519, N14520, N14521, N14522,
         N14523, N14524, N14525, N14526, N14527, N14530, N14531, N14532,
         N14533, N14534, N14535, N14536, N14537, N14538, N14541, N14542,
         N14543, N14544, N14545, N14546, N14547, N14548, N14549, N14552,
         N14553, N14554, N14555, N14556, N14557, N14558, N14559, N14560,
         N14561, N14563, N14564, N14565, N14566, N14567, N14568, N14569,
         N14570, N14571, N14572, N14574, N14575, N14576, N14577, N14578,
         N14579, N14580, N14581, N14582, N14583, N14585, N14586, N14587,
         N14588, N14589, N14590, N14591, N14592, N14593, N14594, N14595, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588;
  wire   [10:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC8_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, 1'b0, 1'b0, 
        olocal}), .CI(1'b0), .SUM(o) );
  hamming_N16000_CC8_DW01_add_1 add_667_root_add_71_I976 ( .A({1'b0, N14583, 
        N14582, N14581, N14580, N14579, N14578, N14577, N14576, N14575, N14574}), .B({N14595, N14594, N14593, N14592, N14591, N14590, N14589, N14588, N14587, 
        N14586, N14585}), .CI(1'b0), .SUM(olocal) );
  hamming_N16000_CC8_DW01_add_2 add_668_root_add_71_I976 ( .A({1'b0, N14561, 
        N14560, N14559, N14558, N14557, N14556, N14555, N14554, N14553, N14552}), .B({1'b0, N14572, N14571, N14570, N14569, N14568, N14567, N14566, N14565, 
        N14564, N14563}), .CI(1'b0), .SUM({N14595, N14594, N14593, N14592, 
        N14591, N14590, N14589, N14588, N14587, N14586, N14585}) );
  hamming_N16000_CC8_DW01_add_3 add_669_root_add_71_I976 ( .A({1'b0, 1'b0, 
        N14538, N14537, N14536, N14535, N14534, N14533, N14532, N14531, N14530}), .B({1'b0, 1'b0, N14549, N14548, N14547, N14546, N14545, N14544, N14543, 
        N14542, N14541}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, N14583, 
        N14582, N14581, N14580, N14579, N14578, N14577, N14576, N14575, N14574}) );
  hamming_N16000_CC8_DW01_add_4 add_670_root_add_71_I976 ( .A({1'b0, 1'b0, 
        N14516, N14515, N14514, N14513, N14512, N14511, N14510, N14509, N14508}), .B({1'b0, 1'b0, N14527, N14526, N14525, N14524, N14523, N14522, N14521, 
        N14520, N14519}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__1, N14572, 
        N14571, N14570, N14569, N14568, N14567, N14566, N14565, N14564, N14563}) );
  hamming_N16000_CC8_DW01_add_5 add_671_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, N14493, N14492, N14491, N14490, N14489, N14488, N14487, N14486}), 
        .B({1'b0, 1'b0, N14505, N14504, N14503, N14502, N14501, N14500, N14499, 
        N14498, N14497}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__2, N14561, 
        N14560, N14559, N14558, N14557, N14556, N14555, N14554, N14553, N14552}) );
  hamming_N16000_CC8_DW01_add_6 add_672_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, N14471, N14470, N14469, N14468, N14467, N14466, N14465, N14464}), 
        .B({1'b0, 1'b0, 1'b0, N14482, N14481, N14480, N14479, N14478, N14477, 
        N14476, N14475}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, N14549, N14548, N14547, N14546, N14545, 
        N14544, N14543, N14542, N14541}) );
  hamming_N16000_CC8_DW01_add_7 add_673_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, N14449, N14448, N14447, N14446, N14445, N14444, N14443, N14442}), 
        .B({1'b0, 1'b0, 1'b0, N14460, N14459, N14458, N14457, N14456, N14455, 
        N14454, N14453}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, N14538, N14537, N14536, N14535, N14534, 
        N14533, N14532, N14531, N14530}) );
  hamming_N16000_CC8_DW01_add_8 add_674_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, N14427, N14426, N14425, N14424, N14423, N14422, N14421, N14420}), 
        .B({1'b0, 1'b0, 1'b0, N14438, N14437, N14436, N14435, N14434, N14433, 
        N14432, N14431}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, N14527, N14526, N14525, N14524, N14523, 
        N14522, N14521, N14520, N14519}) );
  hamming_N16000_CC8_DW01_add_9 add_675_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, N14405, N14404, N14403, N14402, N14401, N14400, N14399, N14398}), 
        .B({1'b0, 1'b0, 1'b0, N14416, N14415, N14414, N14413, N14412, N14411, 
        N14410, N14409}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, N14516, N14515, N14514, N14513, N14512, 
        N14511, N14510, N14509, N14508}) );
  hamming_N16000_CC8_DW01_add_10 add_676_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14382, N14381, N14380, N14379, N14378, N14377, N14376}), 
        .B({1'b0, 1'b0, 1'b0, N14394, N14393, N14392, N14391, N14390, N14389, 
        N14388, N14387}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, N14505, N14504, N14503, N14502, N14501, 
        N14500, N14499, N14498, N14497}) );
  hamming_N16000_CC8_DW01_add_11 add_677_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14360, N14359, N14358, N14357, N14356, N14355, N14354}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14371, N14370, N14369, N14368, N14367, 
        N14366, N14365}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, N14493, N14492, 
        N14491, N14490, N14489, N14488, N14487, N14486}) );
  hamming_N16000_CC8_DW01_add_12 add_678_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14338, N14337, N14336, N14335, N14334, N14333, N14332}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14349, N14348, N14347, N14346, N14345, 
        N14344, N14343}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, N14482, N14481, 
        N14480, N14479, N14478, N14477, N14476, N14475}) );
  hamming_N16000_CC8_DW01_add_13 add_679_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14316, N14315, N14314, N14313, N14312, N14311, N14310}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14327, N14326, N14325, N14324, N14323, 
        N14322, N14321}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, N14471, N14470, 
        N14469, N14468, N14467, N14466, N14465, N14464}) );
  hamming_N16000_CC8_DW01_add_14 add_680_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14294, N14293, N14292, N14291, N14290, N14289, N14288}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14305, N14304, N14303, N14302, N14301, 
        N14300, N14299}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, N14460, N14459, 
        N14458, N14457, N14456, N14455, N14454, N14453}) );
  hamming_N16000_CC8_DW01_add_15 add_681_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14272, N14271, N14270, N14269, N14268, N14267, N14266}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14283, N14282, N14281, N14280, N14279, 
        N14278, N14277}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, N14449, N14448, 
        N14447, N14446, N14445, N14444, N14443, N14442}) );
  hamming_N16000_CC8_DW01_add_16 add_682_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14250, N14249, N14248, N14247, N14246, N14245, N14244}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14261, N14260, N14259, N14258, N14257, 
        N14256, N14255}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, N14438, N14437, 
        N14436, N14435, N14434, N14433, N14432, N14431}) );
  hamming_N16000_CC8_DW01_add_17 add_683_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14228, N14227, N14226, N14225, N14224, N14223, N14222}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14239, N14238, N14237, N14236, N14235, 
        N14234, N14233}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, N14427, N14426, 
        N14425, N14424, N14423, N14422, N14421, N14420}) );
  hamming_N16000_CC8_DW01_add_18 add_684_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14206, N14205, N14204, N14203, N14202, N14201, N14200}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14217, N14216, N14215, N14214, N14213, 
        N14212, N14211}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, N14416, N14415, 
        N14414, N14413, N14412, N14411, N14410, N14409}) );
  hamming_N16000_CC8_DW01_add_19 add_685_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14184, N14183, N14182, N14181, N14180, N14179, N14178}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14195, N14194, N14193, N14192, N14191, 
        N14190, N14189}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, N14405, N14404, 
        N14403, N14402, N14401, N14400, N14399, N14398}) );
  hamming_N16000_CC8_DW01_add_20 add_686_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N14162, N14161, N14160, N14159, N14158, N14157, N14156}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, N14173, N14172, N14171, N14170, N14169, 
        N14168, N14167}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, N14394, N14393, 
        N14392, N14391, N14390, N14389, N14388, N14387}) );
  hamming_N16000_CC8_DW01_add_21 add_687_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N14139, N14138, N14137, N14136, N14135, N14134}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N14150, N14149, N14148, N14147, 
        N14146, N14145}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, N14382, N14381, N14380, N14379, N14378, 
        N14377, N14376}) );
  hamming_N16000_CC8_DW01_add_22 add_688_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N14117, N14116, N14115, N14114, N14113, N14112}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N14128, N14127, N14126, N14125, 
        N14124, N14123}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, N14371, N14370, N14369, N14368, N14367, 
        N14366, N14365}) );
  hamming_N16000_CC8_DW01_add_23 add_689_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N14095, N14094, N14093, N14092, N14091, N14090}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N14106, N14105, N14104, N14103, 
        N14102, N14101}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, N14360, N14359, N14358, N14357, N14356, 
        N14355, N14354}) );
  hamming_N16000_CC8_DW01_add_24 add_690_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N14073, N14072, N14071, N14070, N14069, N14068}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N14084, N14083, N14082, N14081, 
        N14080, N14079}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, N14349, N14348, N14347, N14346, N14345, 
        N14344, N14343}) );
  hamming_N16000_CC8_DW01_add_25 add_691_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N14051, N14050, N14049, N14048, N14047, N14046}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N14062, N14061, N14060, N14059, 
        N14058, N14057}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, N14338, N14337, N14336, N14335, N14334, 
        N14333, N14332}) );
  hamming_N16000_CC8_DW01_add_26 add_692_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N14029, N14028, N14027, N14026, N14025, N14024}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N14040, N14039, N14038, N14037, 
        N14036, N14035}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, N14327, N14326, N14325, N14324, N14323, 
        N14322, N14321}) );
  hamming_N16000_CC8_DW01_add_27 add_693_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N14007, N14006, N14005, N14004, N14003, N14002}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N14018, N14017, N14016, N14015, 
        N14014, N14013}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, N14316, N14315, N14314, N14313, N14312, 
        N14311, N14310}) );
  hamming_N16000_CC8_DW01_add_28 add_694_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13985, N13984, N13983, N13982, N13981, N13980}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13996, N13995, N13994, N13993, 
        N13992, N13991}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, N14305, N14304, N14303, N14302, N14301, 
        N14300, N14299}) );
  hamming_N16000_CC8_DW01_add_29 add_695_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13963, N13962, N13961, N13960, N13959, N13958}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13974, N13973, N13972, N13971, 
        N13970, N13969}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, N14294, N14293, N14292, N14291, N14290, 
        N14289, N14288}) );
  hamming_N16000_CC8_DW01_add_30 add_696_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13941, N13940, N13939, N13938, N13937, N13936}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13952, N13951, N13950, N13949, 
        N13948, N13947}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, N14283, N14282, N14281, N14280, N14279, 
        N14278, N14277}) );
  hamming_N16000_CC8_DW01_add_31 add_697_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13919, N13918, N13917, N13916, N13915, N13914}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13930, N13929, N13928, N13927, 
        N13926, N13925}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, N14272, N14271, N14270, N14269, N14268, 
        N14267, N14266}) );
  hamming_N16000_CC8_DW01_add_32 add_698_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13897, N13896, N13895, N13894, N13893, N13892}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13908, N13907, N13906, N13905, 
        N13904, N13903}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, N14261, N14260, N14259, N14258, N14257, 
        N14256, N14255}) );
  hamming_N16000_CC8_DW01_add_33 add_699_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13875, N13874, N13873, N13872, N13871, N13870}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13886, N13885, N13884, N13883, 
        N13882, N13881}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, N14250, N14249, N14248, N14247, N14246, 
        N14245, N14244}) );
  hamming_N16000_CC8_DW01_add_34 add_700_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13853, N13852, N13851, N13850, N13849, N13848}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13864, N13863, N13862, N13861, 
        N13860, N13859}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, N14239, N14238, N14237, N14236, N14235, 
        N14234, N14233}) );
  hamming_N16000_CC8_DW01_add_35 add_701_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13831, N13830, N13829, N13828, N13827, N13826}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13842, N13841, N13840, N13839, 
        N13838, N13837}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, N14228, N14227, N14226, N14225, N14224, 
        N14223, N14222}) );
  hamming_N16000_CC8_DW01_add_36 add_702_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13809, N13808, N13807, N13806, N13805, N13804}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13820, N13819, N13818, N13817, 
        N13816, N13815}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, N14217, N14216, N14215, N14214, N14213, 
        N14212, N14211}) );
  hamming_N16000_CC8_DW01_add_37 add_703_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13787, N13786, N13785, N13784, N13783, N13782}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13798, N13797, N13796, N13795, 
        N13794, N13793}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, N14206, N14205, N14204, N14203, N14202, 
        N14201, N14200}) );
  hamming_N16000_CC8_DW01_add_38 add_704_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13765, N13764, N13763, N13762, N13761, N13760}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13776, N13775, N13774, N13773, 
        N13772, N13771}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, N14195, N14194, N14193, N14192, N14191, 
        N14190, N14189}) );
  hamming_N16000_CC8_DW01_add_39 add_705_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13743, N13742, N13741, N13740, N13739, N13738}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13754, N13753, N13752, N13751, 
        N13750, N13749}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, N14184, N14183, N14182, N14181, N14180, 
        N14179, N14178}) );
  hamming_N16000_CC8_DW01_add_40 add_706_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13721, N13720, N13719, N13718, N13717, N13716}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13732, N13731, N13730, N13729, 
        N13728, N13727}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, N14173, N14172, N14171, N14170, N14169, 
        N14168, N14167}) );
  hamming_N16000_CC8_DW01_add_41 add_707_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N13699, N13698, N13697, N13696, N13695, N13694}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13710, N13709, N13708, N13707, 
        N13706, N13705}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, N14162, N14161, N14160, N14159, N14158, 
        N14157, N14156}) );
  hamming_N16000_CC8_DW01_add_42 add_708_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13676, N13675, N13674, N13673, N13672}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13687, N13686, N13685, N13684, 
        N13683}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, N14150, N14149, 
        N14148, N14147, N14146, N14145}) );
  hamming_N16000_CC8_DW01_add_43 add_709_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13654, N13653, N13652, N13651, N13650}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13665, N13664, N13663, N13662, 
        N13661}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, N14139, N14138, 
        N14137, N14136, N14135, N14134}) );
  hamming_N16000_CC8_DW01_add_44 add_710_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13632, N13631, N13630, N13629, N13628}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13643, N13642, N13641, N13640, 
        N13639}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, N14128, N14127, 
        N14126, N14125, N14124, N14123}) );
  hamming_N16000_CC8_DW01_add_45 add_711_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13610, N13609, N13608, N13607, N13606}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13621, N13620, N13619, N13618, 
        N13617}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, N14117, N14116, 
        N14115, N14114, N14113, N14112}) );
  hamming_N16000_CC8_DW01_add_46 add_712_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13588, N13587, N13586, N13585, N13584}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13599, N13598, N13597, N13596, 
        N13595}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, N14106, N14105, 
        N14104, N14103, N14102, N14101}) );
  hamming_N16000_CC8_DW01_add_47 add_713_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13566, N13565, N13564, N13563, N13562}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13577, N13576, N13575, N13574, 
        N13573}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, N14095, N14094, 
        N14093, N14092, N14091, N14090}) );
  hamming_N16000_CC8_DW01_add_48 add_714_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13544, N13543, N13542, N13541, N13540}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13555, N13554, N13553, N13552, 
        N13551}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, N14084, N14083, 
        N14082, N14081, N14080, N14079}) );
  hamming_N16000_CC8_DW01_add_49 add_715_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13522, N13521, N13520, N13519, N13518}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13533, N13532, N13531, N13530, 
        N13529}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, N14073, N14072, 
        N14071, N14070, N14069, N14068}) );
  hamming_N16000_CC8_DW01_add_50 add_716_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13500, N13499, N13498, N13497, N13496}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13511, N13510, N13509, N13508, 
        N13507}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, N14062, N14061, 
        N14060, N14059, N14058, N14057}) );
  hamming_N16000_CC8_DW01_add_51 add_717_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13478, N13477, N13476, N13475, N13474}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13489, N13488, N13487, N13486, 
        N13485}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, N14051, N14050, 
        N14049, N14048, N14047, N14046}) );
  hamming_N16000_CC8_DW01_add_52 add_718_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13456, N13455, N13454, N13453, N13452}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13467, N13466, N13465, N13464, 
        N13463}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, N14040, N14039, 
        N14038, N14037, N14036, N14035}) );
  hamming_N16000_CC8_DW01_add_53 add_719_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13434, N13433, N13432, N13431, N13430}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13445, N13444, N13443, N13442, 
        N13441}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, SYNOPSYS_UNCONNECTED__186, N14029, N14028, 
        N14027, N14026, N14025, N14024}) );
  hamming_N16000_CC8_DW01_add_54 add_720_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13412, N13411, N13410, N13409, N13408}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13423, N13422, N13421, N13420, 
        N13419}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, N14018, N14017, 
        N14016, N14015, N14014, N14013}) );
  hamming_N16000_CC8_DW01_add_55 add_721_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13390, N13389, N13388, N13387, N13386}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13401, N13400, N13399, N13398, 
        N13397}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__192, 
        SYNOPSYS_UNCONNECTED__193, SYNOPSYS_UNCONNECTED__194, 
        SYNOPSYS_UNCONNECTED__195, SYNOPSYS_UNCONNECTED__196, N14007, N14006, 
        N14005, N14004, N14003, N14002}) );
  hamming_N16000_CC8_DW01_add_56 add_722_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13368, N13367, N13366, N13365, N13364}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13379, N13378, N13377, N13376, 
        N13375}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, N13996, N13995, 
        N13994, N13993, N13992, N13991}) );
  hamming_N16000_CC8_DW01_add_57 add_723_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13346, N13345, N13344, N13343, N13342}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13357, N13356, N13355, N13354, 
        N13353}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__202, 
        SYNOPSYS_UNCONNECTED__203, SYNOPSYS_UNCONNECTED__204, 
        SYNOPSYS_UNCONNECTED__205, SYNOPSYS_UNCONNECTED__206, N13985, N13984, 
        N13983, N13982, N13981, N13980}) );
  hamming_N16000_CC8_DW01_add_58 add_724_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13324, N13323, N13322, N13321, N13320}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13335, N13334, N13333, N13332, 
        N13331}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, N13974, N13973, 
        N13972, N13971, N13970, N13969}) );
  hamming_N16000_CC8_DW01_add_59 add_725_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13302, N13301, N13300, N13299, N13298}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13313, N13312, N13311, N13310, 
        N13309}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__212, 
        SYNOPSYS_UNCONNECTED__213, SYNOPSYS_UNCONNECTED__214, 
        SYNOPSYS_UNCONNECTED__215, SYNOPSYS_UNCONNECTED__216, N13963, N13962, 
        N13961, N13960, N13959, N13958}) );
  hamming_N16000_CC8_DW01_add_60 add_726_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13280, N13279, N13278, N13277, N13276}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13291, N13290, N13289, N13288, 
        N13287}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, N13952, N13951, 
        N13950, N13949, N13948, N13947}) );
  hamming_N16000_CC8_DW01_add_61 add_727_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13258, N13257, N13256, N13255, N13254}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13269, N13268, N13267, N13266, 
        N13265}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__222, 
        SYNOPSYS_UNCONNECTED__223, SYNOPSYS_UNCONNECTED__224, 
        SYNOPSYS_UNCONNECTED__225, SYNOPSYS_UNCONNECTED__226, N13941, N13940, 
        N13939, N13938, N13937, N13936}) );
  hamming_N16000_CC8_DW01_add_62 add_728_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13236, N13235, N13234, N13233, N13232}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13247, N13246, N13245, N13244, 
        N13243}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, N13930, N13929, 
        N13928, N13927, N13926, N13925}) );
  hamming_N16000_CC8_DW01_add_63 add_729_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13214, N13213, N13212, N13211, N13210}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13225, N13224, N13223, N13222, 
        N13221}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__232, 
        SYNOPSYS_UNCONNECTED__233, SYNOPSYS_UNCONNECTED__234, 
        SYNOPSYS_UNCONNECTED__235, SYNOPSYS_UNCONNECTED__236, N13919, N13918, 
        N13917, N13916, N13915, N13914}) );
  hamming_N16000_CC8_DW01_add_64 add_730_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13192, N13191, N13190, N13189, N13188}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13203, N13202, N13201, N13200, 
        N13199}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, N13908, N13907, 
        N13906, N13905, N13904, N13903}) );
  hamming_N16000_CC8_DW01_add_65 add_731_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13170, N13169, N13168, N13167, N13166}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13181, N13180, N13179, N13178, 
        N13177}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__242, 
        SYNOPSYS_UNCONNECTED__243, SYNOPSYS_UNCONNECTED__244, 
        SYNOPSYS_UNCONNECTED__245, SYNOPSYS_UNCONNECTED__246, N13897, N13896, 
        N13895, N13894, N13893, N13892}) );
  hamming_N16000_CC8_DW01_add_66 add_732_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13148, N13147, N13146, N13145, N13144}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13159, N13158, N13157, N13156, 
        N13155}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, N13886, N13885, 
        N13884, N13883, N13882, N13881}) );
  hamming_N16000_CC8_DW01_add_67 add_733_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13126, N13125, N13124, N13123, N13122}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13137, N13136, N13135, N13134, 
        N13133}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__252, 
        SYNOPSYS_UNCONNECTED__253, SYNOPSYS_UNCONNECTED__254, 
        SYNOPSYS_UNCONNECTED__255, SYNOPSYS_UNCONNECTED__256, N13875, N13874, 
        N13873, N13872, N13871, N13870}) );
  hamming_N16000_CC8_DW01_add_68 add_734_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13104, N13103, N13102, N13101, N13100}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13115, N13114, N13113, N13112, 
        N13111}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, N13864, N13863, 
        N13862, N13861, N13860, N13859}) );
  hamming_N16000_CC8_DW01_add_69 add_735_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13082, N13081, N13080, N13079, N13078}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13093, N13092, N13091, N13090, 
        N13089}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__262, 
        SYNOPSYS_UNCONNECTED__263, SYNOPSYS_UNCONNECTED__264, 
        SYNOPSYS_UNCONNECTED__265, SYNOPSYS_UNCONNECTED__266, N13853, N13852, 
        N13851, N13850, N13849, N13848}) );
  hamming_N16000_CC8_DW01_add_70 add_736_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13060, N13059, N13058, N13057, N13056}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13071, N13070, N13069, N13068, 
        N13067}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, N13842, N13841, 
        N13840, N13839, N13838, N13837}) );
  hamming_N16000_CC8_DW01_add_71 add_737_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13038, N13037, N13036, N13035, N13034}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13049, N13048, N13047, N13046, 
        N13045}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__272, 
        SYNOPSYS_UNCONNECTED__273, SYNOPSYS_UNCONNECTED__274, 
        SYNOPSYS_UNCONNECTED__275, SYNOPSYS_UNCONNECTED__276, N13831, N13830, 
        N13829, N13828, N13827, N13826}) );
  hamming_N16000_CC8_DW01_add_72 add_738_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N13016, N13015, N13014, N13013, N13012}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13027, N13026, N13025, N13024, 
        N13023}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, N13820, N13819, 
        N13818, N13817, N13816, N13815}) );
  hamming_N16000_CC8_DW01_add_73 add_739_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12994, N12993, N12992, N12991, N12990}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N13005, N13004, N13003, N13002, 
        N13001}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__282, 
        SYNOPSYS_UNCONNECTED__283, SYNOPSYS_UNCONNECTED__284, 
        SYNOPSYS_UNCONNECTED__285, SYNOPSYS_UNCONNECTED__286, N13809, N13808, 
        N13807, N13806, N13805, N13804}) );
  hamming_N16000_CC8_DW01_add_74 add_740_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12972, N12971, N12970, N12969, N12968}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12983, N12982, N12981, N12980, 
        N12979}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, N13798, N13797, 
        N13796, N13795, N13794, N13793}) );
  hamming_N16000_CC8_DW01_add_75 add_741_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12950, N12949, N12948, N12947, N12946}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12961, N12960, N12959, N12958, 
        N12957}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__292, 
        SYNOPSYS_UNCONNECTED__293, SYNOPSYS_UNCONNECTED__294, 
        SYNOPSYS_UNCONNECTED__295, SYNOPSYS_UNCONNECTED__296, N13787, N13786, 
        N13785, N13784, N13783, N13782}) );
  hamming_N16000_CC8_DW01_add_76 add_742_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12928, N12927, N12926, N12925, N12924}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12939, N12938, N12937, N12936, 
        N12935}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, N13776, N13775, 
        N13774, N13773, N13772, N13771}) );
  hamming_N16000_CC8_DW01_add_77 add_743_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12906, N12905, N12904, N12903, N12902}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12917, N12916, N12915, N12914, 
        N12913}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__302, 
        SYNOPSYS_UNCONNECTED__303, SYNOPSYS_UNCONNECTED__304, 
        SYNOPSYS_UNCONNECTED__305, SYNOPSYS_UNCONNECTED__306, N13765, N13764, 
        N13763, N13762, N13761, N13760}) );
  hamming_N16000_CC8_DW01_add_78 add_744_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12884, N12883, N12882, N12881, N12880}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12895, N12894, N12893, N12892, 
        N12891}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, N13754, N13753, 
        N13752, N13751, N13750, N13749}) );
  hamming_N16000_CC8_DW01_add_79 add_745_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12862, N12861, N12860, N12859, N12858}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12873, N12872, N12871, N12870, 
        N12869}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__312, 
        SYNOPSYS_UNCONNECTED__313, SYNOPSYS_UNCONNECTED__314, 
        SYNOPSYS_UNCONNECTED__315, SYNOPSYS_UNCONNECTED__316, N13743, N13742, 
        N13741, N13740, N13739, N13738}) );
  hamming_N16000_CC8_DW01_add_80 add_746_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12840, N12839, N12838, N12837, N12836}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12851, N12850, N12849, N12848, 
        N12847}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, N13732, N13731, 
        N13730, N13729, N13728, N13727}) );
  hamming_N16000_CC8_DW01_add_81 add_747_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12818, N12817, N12816, N12815, N12814}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12829, N12828, N12827, N12826, 
        N12825}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__322, 
        SYNOPSYS_UNCONNECTED__323, SYNOPSYS_UNCONNECTED__324, 
        SYNOPSYS_UNCONNECTED__325, SYNOPSYS_UNCONNECTED__326, N13721, N13720, 
        N13719, N13718, N13717, N13716}) );
  hamming_N16000_CC8_DW01_add_82 add_748_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N12796, N12795, N12794, N12793, N12792}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12807, N12806, N12805, N12804, 
        N12803}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, N13710, N13709, 
        N13708, N13707, N13706, N13705}) );
  hamming_N16000_CC8_DW01_add_83 add_749_root_add_71_I976 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12773, N12772, N12771, N12770}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N12785, N12784, N12783, N12782, 
        N12781}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__332, 
        SYNOPSYS_UNCONNECTED__333, SYNOPSYS_UNCONNECTED__334, 
        SYNOPSYS_UNCONNECTED__335, SYNOPSYS_UNCONNECTED__336, N13699, N13698, 
        N13697, N13696, N13695, N13694}) );
  NAND U3353 ( .A(n1354), .B(n1355), .Z(N13687) );
  NANDN U3354 ( .A(n1356), .B(n1357), .Z(n1355) );
  OR U3355 ( .A(n1358), .B(n1359), .Z(n1357) );
  NAND U3356 ( .A(n1358), .B(n1359), .Z(n1354) );
  XOR U3357 ( .A(n1358), .B(n1360), .Z(N13686) );
  XNOR U3358 ( .A(n1356), .B(n1359), .Z(n1360) );
  AND U3359 ( .A(n1361), .B(n1362), .Z(n1359) );
  NANDN U3360 ( .A(n1363), .B(n1364), .Z(n1362) );
  NANDN U3361 ( .A(n1365), .B(n1366), .Z(n1364) );
  NANDN U3362 ( .A(n1366), .B(n1365), .Z(n1361) );
  NAND U3363 ( .A(n1367), .B(n1368), .Z(n1356) );
  NANDN U3364 ( .A(n1369), .B(n1370), .Z(n1368) );
  OR U3365 ( .A(n1371), .B(n1372), .Z(n1370) );
  NAND U3366 ( .A(n1372), .B(n1371), .Z(n1367) );
  AND U3367 ( .A(n1373), .B(n1374), .Z(n1358) );
  NANDN U3368 ( .A(n1375), .B(n1376), .Z(n1374) );
  NANDN U3369 ( .A(n1377), .B(n1378), .Z(n1376) );
  NANDN U3370 ( .A(n1378), .B(n1377), .Z(n1373) );
  XOR U3371 ( .A(n1372), .B(n1379), .Z(N13685) );
  XOR U3372 ( .A(n1369), .B(n1371), .Z(n1379) );
  XNOR U3373 ( .A(n1365), .B(n1380), .Z(n1371) );
  XNOR U3374 ( .A(n1363), .B(n1366), .Z(n1380) );
  NAND U3375 ( .A(n1381), .B(n1382), .Z(n1366) );
  NAND U3376 ( .A(n1383), .B(n1384), .Z(n1382) );
  OR U3377 ( .A(n1385), .B(n1386), .Z(n1383) );
  NANDN U3378 ( .A(n1387), .B(n1385), .Z(n1381) );
  IV U3379 ( .A(n1386), .Z(n1387) );
  NAND U3380 ( .A(n1388), .B(n1389), .Z(n1363) );
  NAND U3381 ( .A(n1390), .B(n1391), .Z(n1389) );
  NANDN U3382 ( .A(n1392), .B(n1393), .Z(n1390) );
  NANDN U3383 ( .A(n1393), .B(n1392), .Z(n1388) );
  AND U3384 ( .A(n1394), .B(n1395), .Z(n1365) );
  NAND U3385 ( .A(n1396), .B(n1397), .Z(n1395) );
  OR U3386 ( .A(n1398), .B(n1399), .Z(n1396) );
  NANDN U3387 ( .A(n1400), .B(n1398), .Z(n1394) );
  NAND U3388 ( .A(n1401), .B(n1402), .Z(n1369) );
  NANDN U3389 ( .A(n1403), .B(n1404), .Z(n1402) );
  OR U3390 ( .A(n1405), .B(n1406), .Z(n1404) );
  NANDN U3391 ( .A(n1407), .B(n1405), .Z(n1401) );
  IV U3392 ( .A(n1406), .Z(n1407) );
  XNOR U3393 ( .A(n1377), .B(n1408), .Z(n1372) );
  XNOR U3394 ( .A(n1375), .B(n1378), .Z(n1408) );
  NAND U3395 ( .A(n1409), .B(n1410), .Z(n1378) );
  NAND U3396 ( .A(n1411), .B(n1412), .Z(n1410) );
  OR U3397 ( .A(n1413), .B(n1414), .Z(n1411) );
  NANDN U3398 ( .A(n1415), .B(n1413), .Z(n1409) );
  IV U3399 ( .A(n1414), .Z(n1415) );
  NAND U3400 ( .A(n1416), .B(n1417), .Z(n1375) );
  NAND U3401 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U3402 ( .A(n1420), .B(n1421), .Z(n1418) );
  NANDN U3403 ( .A(n1421), .B(n1420), .Z(n1416) );
  AND U3404 ( .A(n1422), .B(n1423), .Z(n1377) );
  NAND U3405 ( .A(n1424), .B(n1425), .Z(n1423) );
  OR U3406 ( .A(n1426), .B(n1427), .Z(n1424) );
  NANDN U3407 ( .A(n1428), .B(n1426), .Z(n1422) );
  XNOR U3408 ( .A(n1403), .B(n1429), .Z(N13684) );
  XOR U3409 ( .A(n1405), .B(n1406), .Z(n1429) );
  XNOR U3410 ( .A(n1419), .B(n1430), .Z(n1406) );
  XOR U3411 ( .A(n1420), .B(n1421), .Z(n1430) );
  XOR U3412 ( .A(n1426), .B(n1431), .Z(n1421) );
  XOR U3413 ( .A(n1425), .B(n1428), .Z(n1431) );
  IV U3414 ( .A(n1427), .Z(n1428) );
  NAND U3415 ( .A(n1432), .B(n1433), .Z(n1427) );
  OR U3416 ( .A(n1434), .B(n1435), .Z(n1433) );
  OR U3417 ( .A(n1436), .B(n1437), .Z(n1432) );
  NAND U3418 ( .A(n1438), .B(n1439), .Z(n1425) );
  OR U3419 ( .A(n1440), .B(n1441), .Z(n1439) );
  OR U3420 ( .A(n1442), .B(n1443), .Z(n1438) );
  NOR U3421 ( .A(n1444), .B(n1445), .Z(n1426) );
  ANDN U3422 ( .B(n1446), .A(n1447), .Z(n1420) );
  XNOR U3423 ( .A(n1413), .B(n1448), .Z(n1419) );
  XNOR U3424 ( .A(n1412), .B(n1414), .Z(n1448) );
  NAND U3425 ( .A(n1449), .B(n1450), .Z(n1414) );
  OR U3426 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U3427 ( .A(n1453), .B(n1454), .Z(n1449) );
  NAND U3428 ( .A(n1455), .B(n1456), .Z(n1412) );
  OR U3429 ( .A(n1457), .B(n1458), .Z(n1456) );
  OR U3430 ( .A(n1459), .B(n1460), .Z(n1455) );
  ANDN U3431 ( .B(n1461), .A(n1462), .Z(n1413) );
  IV U3432 ( .A(n1463), .Z(n1461) );
  ANDN U3433 ( .B(n1464), .A(n1465), .Z(n1405) );
  XOR U3434 ( .A(n1391), .B(n1466), .Z(n1403) );
  XOR U3435 ( .A(n1392), .B(n1393), .Z(n1466) );
  XOR U3436 ( .A(n1398), .B(n1467), .Z(n1393) );
  XOR U3437 ( .A(n1397), .B(n1400), .Z(n1467) );
  IV U3438 ( .A(n1399), .Z(n1400) );
  NAND U3439 ( .A(n1468), .B(n1469), .Z(n1399) );
  OR U3440 ( .A(n1470), .B(n1471), .Z(n1469) );
  OR U3441 ( .A(n1472), .B(n1473), .Z(n1468) );
  NAND U3442 ( .A(n1474), .B(n1475), .Z(n1397) );
  OR U3443 ( .A(n1476), .B(n1477), .Z(n1475) );
  OR U3444 ( .A(n1478), .B(n1479), .Z(n1474) );
  NOR U3445 ( .A(n1480), .B(n1481), .Z(n1398) );
  ANDN U3446 ( .B(n1482), .A(n1483), .Z(n1392) );
  IV U3447 ( .A(n1484), .Z(n1482) );
  XNOR U3448 ( .A(n1385), .B(n1485), .Z(n1391) );
  XNOR U3449 ( .A(n1384), .B(n1386), .Z(n1485) );
  NAND U3450 ( .A(n1486), .B(n1487), .Z(n1386) );
  OR U3451 ( .A(n1488), .B(n1489), .Z(n1487) );
  OR U3452 ( .A(n1490), .B(n1491), .Z(n1486) );
  NAND U3453 ( .A(n1492), .B(n1493), .Z(n1384) );
  OR U3454 ( .A(n1494), .B(n1495), .Z(n1493) );
  OR U3455 ( .A(n1496), .B(n1497), .Z(n1492) );
  ANDN U3456 ( .B(n1498), .A(n1499), .Z(n1385) );
  IV U3457 ( .A(n1500), .Z(n1498) );
  XNOR U3458 ( .A(n1465), .B(n1464), .Z(N13683) );
  XOR U3459 ( .A(n1484), .B(n1483), .Z(n1464) );
  XNOR U3460 ( .A(n1499), .B(n1500), .Z(n1483) );
  XNOR U3461 ( .A(n1494), .B(n1495), .Z(n1500) );
  XNOR U3462 ( .A(n1496), .B(n1497), .Z(n1495) );
  XNOR U3463 ( .A(y[1981]), .B(x[1981]), .Z(n1497) );
  XNOR U3464 ( .A(y[1982]), .B(x[1982]), .Z(n1496) );
  XNOR U3465 ( .A(y[1980]), .B(x[1980]), .Z(n1494) );
  XNOR U3466 ( .A(n1488), .B(n1489), .Z(n1499) );
  XNOR U3467 ( .A(y[1977]), .B(x[1977]), .Z(n1489) );
  XNOR U3468 ( .A(n1490), .B(n1491), .Z(n1488) );
  XNOR U3469 ( .A(y[1978]), .B(x[1978]), .Z(n1491) );
  XNOR U3470 ( .A(y[1979]), .B(x[1979]), .Z(n1490) );
  XNOR U3471 ( .A(n1481), .B(n1480), .Z(n1484) );
  XNOR U3472 ( .A(n1476), .B(n1477), .Z(n1480) );
  XNOR U3473 ( .A(y[1974]), .B(x[1974]), .Z(n1477) );
  XNOR U3474 ( .A(n1478), .B(n1479), .Z(n1476) );
  XNOR U3475 ( .A(y[1975]), .B(x[1975]), .Z(n1479) );
  XNOR U3476 ( .A(y[1976]), .B(x[1976]), .Z(n1478) );
  XNOR U3477 ( .A(n1470), .B(n1471), .Z(n1481) );
  XNOR U3478 ( .A(y[1971]), .B(x[1971]), .Z(n1471) );
  XNOR U3479 ( .A(n1472), .B(n1473), .Z(n1470) );
  XNOR U3480 ( .A(y[1972]), .B(x[1972]), .Z(n1473) );
  XNOR U3481 ( .A(y[1973]), .B(x[1973]), .Z(n1472) );
  XOR U3482 ( .A(n1446), .B(n1447), .Z(n1465) );
  XNOR U3483 ( .A(n1462), .B(n1463), .Z(n1447) );
  XNOR U3484 ( .A(n1457), .B(n1458), .Z(n1463) );
  XNOR U3485 ( .A(n1459), .B(n1460), .Z(n1458) );
  XNOR U3486 ( .A(y[1969]), .B(x[1969]), .Z(n1460) );
  XNOR U3487 ( .A(y[1970]), .B(x[1970]), .Z(n1459) );
  XNOR U3488 ( .A(y[1968]), .B(x[1968]), .Z(n1457) );
  XNOR U3489 ( .A(n1451), .B(n1452), .Z(n1462) );
  XNOR U3490 ( .A(y[1965]), .B(x[1965]), .Z(n1452) );
  XNOR U3491 ( .A(n1453), .B(n1454), .Z(n1451) );
  XNOR U3492 ( .A(y[1966]), .B(x[1966]), .Z(n1454) );
  XNOR U3493 ( .A(y[1967]), .B(x[1967]), .Z(n1453) );
  XOR U3494 ( .A(n1445), .B(n1444), .Z(n1446) );
  XNOR U3495 ( .A(n1440), .B(n1441), .Z(n1444) );
  XNOR U3496 ( .A(y[1962]), .B(x[1962]), .Z(n1441) );
  XNOR U3497 ( .A(n1442), .B(n1443), .Z(n1440) );
  XNOR U3498 ( .A(y[1963]), .B(x[1963]), .Z(n1443) );
  XNOR U3499 ( .A(y[1964]), .B(x[1964]), .Z(n1442) );
  XNOR U3500 ( .A(n1434), .B(n1435), .Z(n1445) );
  XNOR U3501 ( .A(y[1959]), .B(x[1959]), .Z(n1435) );
  XNOR U3502 ( .A(n1436), .B(n1437), .Z(n1434) );
  XNOR U3503 ( .A(y[1960]), .B(x[1960]), .Z(n1437) );
  XNOR U3504 ( .A(y[1961]), .B(x[1961]), .Z(n1436) );
  NAND U3505 ( .A(n1501), .B(n1502), .Z(N13676) );
  NANDN U3506 ( .A(n1503), .B(n1504), .Z(n1502) );
  OR U3507 ( .A(n1505), .B(n1506), .Z(n1504) );
  NAND U3508 ( .A(n1505), .B(n1506), .Z(n1501) );
  XOR U3509 ( .A(n1505), .B(n1507), .Z(N13675) );
  XNOR U3510 ( .A(n1503), .B(n1506), .Z(n1507) );
  AND U3511 ( .A(n1508), .B(n1509), .Z(n1506) );
  NANDN U3512 ( .A(n1510), .B(n1511), .Z(n1509) );
  NANDN U3513 ( .A(n1512), .B(n1513), .Z(n1511) );
  NANDN U3514 ( .A(n1513), .B(n1512), .Z(n1508) );
  NAND U3515 ( .A(n1514), .B(n1515), .Z(n1503) );
  NANDN U3516 ( .A(n1516), .B(n1517), .Z(n1515) );
  OR U3517 ( .A(n1518), .B(n1519), .Z(n1517) );
  NAND U3518 ( .A(n1519), .B(n1518), .Z(n1514) );
  AND U3519 ( .A(n1520), .B(n1521), .Z(n1505) );
  NANDN U3520 ( .A(n1522), .B(n1523), .Z(n1521) );
  NANDN U3521 ( .A(n1524), .B(n1525), .Z(n1523) );
  NANDN U3522 ( .A(n1525), .B(n1524), .Z(n1520) );
  XOR U3523 ( .A(n1519), .B(n1526), .Z(N13674) );
  XOR U3524 ( .A(n1516), .B(n1518), .Z(n1526) );
  XNOR U3525 ( .A(n1512), .B(n1527), .Z(n1518) );
  XNOR U3526 ( .A(n1510), .B(n1513), .Z(n1527) );
  NAND U3527 ( .A(n1528), .B(n1529), .Z(n1513) );
  NAND U3528 ( .A(n1530), .B(n1531), .Z(n1529) );
  OR U3529 ( .A(n1532), .B(n1533), .Z(n1530) );
  NANDN U3530 ( .A(n1534), .B(n1532), .Z(n1528) );
  IV U3531 ( .A(n1533), .Z(n1534) );
  NAND U3532 ( .A(n1535), .B(n1536), .Z(n1510) );
  NAND U3533 ( .A(n1537), .B(n1538), .Z(n1536) );
  NANDN U3534 ( .A(n1539), .B(n1540), .Z(n1537) );
  NANDN U3535 ( .A(n1540), .B(n1539), .Z(n1535) );
  AND U3536 ( .A(n1541), .B(n1542), .Z(n1512) );
  NAND U3537 ( .A(n1543), .B(n1544), .Z(n1542) );
  OR U3538 ( .A(n1545), .B(n1546), .Z(n1543) );
  NANDN U3539 ( .A(n1547), .B(n1545), .Z(n1541) );
  NAND U3540 ( .A(n1548), .B(n1549), .Z(n1516) );
  NANDN U3541 ( .A(n1550), .B(n1551), .Z(n1549) );
  OR U3542 ( .A(n1552), .B(n1553), .Z(n1551) );
  NANDN U3543 ( .A(n1554), .B(n1552), .Z(n1548) );
  IV U3544 ( .A(n1553), .Z(n1554) );
  XNOR U3545 ( .A(n1524), .B(n1555), .Z(n1519) );
  XNOR U3546 ( .A(n1522), .B(n1525), .Z(n1555) );
  NAND U3547 ( .A(n1556), .B(n1557), .Z(n1525) );
  NAND U3548 ( .A(n1558), .B(n1559), .Z(n1557) );
  OR U3549 ( .A(n1560), .B(n1561), .Z(n1558) );
  NANDN U3550 ( .A(n1562), .B(n1560), .Z(n1556) );
  IV U3551 ( .A(n1561), .Z(n1562) );
  NAND U3552 ( .A(n1563), .B(n1564), .Z(n1522) );
  NAND U3553 ( .A(n1565), .B(n1566), .Z(n1564) );
  NANDN U3554 ( .A(n1567), .B(n1568), .Z(n1565) );
  NANDN U3555 ( .A(n1568), .B(n1567), .Z(n1563) );
  AND U3556 ( .A(n1569), .B(n1570), .Z(n1524) );
  NAND U3557 ( .A(n1571), .B(n1572), .Z(n1570) );
  OR U3558 ( .A(n1573), .B(n1574), .Z(n1571) );
  NANDN U3559 ( .A(n1575), .B(n1573), .Z(n1569) );
  XNOR U3560 ( .A(n1550), .B(n1576), .Z(N13673) );
  XOR U3561 ( .A(n1552), .B(n1553), .Z(n1576) );
  XNOR U3562 ( .A(n1566), .B(n1577), .Z(n1553) );
  XOR U3563 ( .A(n1567), .B(n1568), .Z(n1577) );
  XOR U3564 ( .A(n1573), .B(n1578), .Z(n1568) );
  XOR U3565 ( .A(n1572), .B(n1575), .Z(n1578) );
  IV U3566 ( .A(n1574), .Z(n1575) );
  NAND U3567 ( .A(n1579), .B(n1580), .Z(n1574) );
  OR U3568 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U3569 ( .A(n1583), .B(n1584), .Z(n1579) );
  NAND U3570 ( .A(n1585), .B(n1586), .Z(n1572) );
  OR U3571 ( .A(n1587), .B(n1588), .Z(n1586) );
  OR U3572 ( .A(n1589), .B(n1590), .Z(n1585) );
  NOR U3573 ( .A(n1591), .B(n1592), .Z(n1573) );
  ANDN U3574 ( .B(n1593), .A(n1594), .Z(n1567) );
  XNOR U3575 ( .A(n1560), .B(n1595), .Z(n1566) );
  XNOR U3576 ( .A(n1559), .B(n1561), .Z(n1595) );
  NAND U3577 ( .A(n1596), .B(n1597), .Z(n1561) );
  OR U3578 ( .A(n1598), .B(n1599), .Z(n1597) );
  OR U3579 ( .A(n1600), .B(n1601), .Z(n1596) );
  NAND U3580 ( .A(n1602), .B(n1603), .Z(n1559) );
  OR U3581 ( .A(n1604), .B(n1605), .Z(n1603) );
  OR U3582 ( .A(n1606), .B(n1607), .Z(n1602) );
  ANDN U3583 ( .B(n1608), .A(n1609), .Z(n1560) );
  IV U3584 ( .A(n1610), .Z(n1608) );
  ANDN U3585 ( .B(n1611), .A(n1612), .Z(n1552) );
  XOR U3586 ( .A(n1538), .B(n1613), .Z(n1550) );
  XOR U3587 ( .A(n1539), .B(n1540), .Z(n1613) );
  XOR U3588 ( .A(n1545), .B(n1614), .Z(n1540) );
  XOR U3589 ( .A(n1544), .B(n1547), .Z(n1614) );
  IV U3590 ( .A(n1546), .Z(n1547) );
  NAND U3591 ( .A(n1615), .B(n1616), .Z(n1546) );
  OR U3592 ( .A(n1617), .B(n1618), .Z(n1616) );
  OR U3593 ( .A(n1619), .B(n1620), .Z(n1615) );
  NAND U3594 ( .A(n1621), .B(n1622), .Z(n1544) );
  OR U3595 ( .A(n1623), .B(n1624), .Z(n1622) );
  OR U3596 ( .A(n1625), .B(n1626), .Z(n1621) );
  NOR U3597 ( .A(n1627), .B(n1628), .Z(n1545) );
  ANDN U3598 ( .B(n1629), .A(n1630), .Z(n1539) );
  IV U3599 ( .A(n1631), .Z(n1629) );
  XNOR U3600 ( .A(n1532), .B(n1632), .Z(n1538) );
  XNOR U3601 ( .A(n1531), .B(n1533), .Z(n1632) );
  NAND U3602 ( .A(n1633), .B(n1634), .Z(n1533) );
  OR U3603 ( .A(n1635), .B(n1636), .Z(n1634) );
  OR U3604 ( .A(n1637), .B(n1638), .Z(n1633) );
  NAND U3605 ( .A(n1639), .B(n1640), .Z(n1531) );
  OR U3606 ( .A(n1641), .B(n1642), .Z(n1640) );
  OR U3607 ( .A(n1643), .B(n1644), .Z(n1639) );
  ANDN U3608 ( .B(n1645), .A(n1646), .Z(n1532) );
  IV U3609 ( .A(n1647), .Z(n1645) );
  XNOR U3610 ( .A(n1612), .B(n1611), .Z(N13672) );
  XOR U3611 ( .A(n1631), .B(n1630), .Z(n1611) );
  XNOR U3612 ( .A(n1646), .B(n1647), .Z(n1630) );
  XNOR U3613 ( .A(n1641), .B(n1642), .Z(n1647) );
  XNOR U3614 ( .A(n1643), .B(n1644), .Z(n1642) );
  XNOR U3615 ( .A(y[1957]), .B(x[1957]), .Z(n1644) );
  XNOR U3616 ( .A(y[1958]), .B(x[1958]), .Z(n1643) );
  XNOR U3617 ( .A(y[1956]), .B(x[1956]), .Z(n1641) );
  XNOR U3618 ( .A(n1635), .B(n1636), .Z(n1646) );
  XNOR U3619 ( .A(y[1953]), .B(x[1953]), .Z(n1636) );
  XNOR U3620 ( .A(n1637), .B(n1638), .Z(n1635) );
  XNOR U3621 ( .A(y[1954]), .B(x[1954]), .Z(n1638) );
  XNOR U3622 ( .A(y[1955]), .B(x[1955]), .Z(n1637) );
  XNOR U3623 ( .A(n1628), .B(n1627), .Z(n1631) );
  XNOR U3624 ( .A(n1623), .B(n1624), .Z(n1627) );
  XNOR U3625 ( .A(y[1950]), .B(x[1950]), .Z(n1624) );
  XNOR U3626 ( .A(n1625), .B(n1626), .Z(n1623) );
  XNOR U3627 ( .A(y[1951]), .B(x[1951]), .Z(n1626) );
  XNOR U3628 ( .A(y[1952]), .B(x[1952]), .Z(n1625) );
  XNOR U3629 ( .A(n1617), .B(n1618), .Z(n1628) );
  XNOR U3630 ( .A(y[1947]), .B(x[1947]), .Z(n1618) );
  XNOR U3631 ( .A(n1619), .B(n1620), .Z(n1617) );
  XNOR U3632 ( .A(y[1948]), .B(x[1948]), .Z(n1620) );
  XNOR U3633 ( .A(y[1949]), .B(x[1949]), .Z(n1619) );
  XOR U3634 ( .A(n1593), .B(n1594), .Z(n1612) );
  XNOR U3635 ( .A(n1609), .B(n1610), .Z(n1594) );
  XNOR U3636 ( .A(n1604), .B(n1605), .Z(n1610) );
  XNOR U3637 ( .A(n1606), .B(n1607), .Z(n1605) );
  XNOR U3638 ( .A(y[1945]), .B(x[1945]), .Z(n1607) );
  XNOR U3639 ( .A(y[1946]), .B(x[1946]), .Z(n1606) );
  XNOR U3640 ( .A(y[1944]), .B(x[1944]), .Z(n1604) );
  XNOR U3641 ( .A(n1598), .B(n1599), .Z(n1609) );
  XNOR U3642 ( .A(y[1941]), .B(x[1941]), .Z(n1599) );
  XNOR U3643 ( .A(n1600), .B(n1601), .Z(n1598) );
  XNOR U3644 ( .A(y[1942]), .B(x[1942]), .Z(n1601) );
  XNOR U3645 ( .A(y[1943]), .B(x[1943]), .Z(n1600) );
  XOR U3646 ( .A(n1592), .B(n1591), .Z(n1593) );
  XNOR U3647 ( .A(n1587), .B(n1588), .Z(n1591) );
  XNOR U3648 ( .A(y[1938]), .B(x[1938]), .Z(n1588) );
  XNOR U3649 ( .A(n1589), .B(n1590), .Z(n1587) );
  XNOR U3650 ( .A(y[1939]), .B(x[1939]), .Z(n1590) );
  XNOR U3651 ( .A(y[1940]), .B(x[1940]), .Z(n1589) );
  XNOR U3652 ( .A(n1581), .B(n1582), .Z(n1592) );
  XNOR U3653 ( .A(y[1935]), .B(x[1935]), .Z(n1582) );
  XNOR U3654 ( .A(n1583), .B(n1584), .Z(n1581) );
  XNOR U3655 ( .A(y[1936]), .B(x[1936]), .Z(n1584) );
  XNOR U3656 ( .A(y[1937]), .B(x[1937]), .Z(n1583) );
  NAND U3657 ( .A(n1648), .B(n1649), .Z(N13665) );
  NANDN U3658 ( .A(n1650), .B(n1651), .Z(n1649) );
  OR U3659 ( .A(n1652), .B(n1653), .Z(n1651) );
  NAND U3660 ( .A(n1652), .B(n1653), .Z(n1648) );
  XOR U3661 ( .A(n1652), .B(n1654), .Z(N13664) );
  XNOR U3662 ( .A(n1650), .B(n1653), .Z(n1654) );
  AND U3663 ( .A(n1655), .B(n1656), .Z(n1653) );
  NANDN U3664 ( .A(n1657), .B(n1658), .Z(n1656) );
  NANDN U3665 ( .A(n1659), .B(n1660), .Z(n1658) );
  NANDN U3666 ( .A(n1660), .B(n1659), .Z(n1655) );
  NAND U3667 ( .A(n1661), .B(n1662), .Z(n1650) );
  NANDN U3668 ( .A(n1663), .B(n1664), .Z(n1662) );
  OR U3669 ( .A(n1665), .B(n1666), .Z(n1664) );
  NAND U3670 ( .A(n1666), .B(n1665), .Z(n1661) );
  AND U3671 ( .A(n1667), .B(n1668), .Z(n1652) );
  NANDN U3672 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U3673 ( .A(n1671), .B(n1672), .Z(n1670) );
  NANDN U3674 ( .A(n1672), .B(n1671), .Z(n1667) );
  XOR U3675 ( .A(n1666), .B(n1673), .Z(N13663) );
  XOR U3676 ( .A(n1663), .B(n1665), .Z(n1673) );
  XNOR U3677 ( .A(n1659), .B(n1674), .Z(n1665) );
  XNOR U3678 ( .A(n1657), .B(n1660), .Z(n1674) );
  NAND U3679 ( .A(n1675), .B(n1676), .Z(n1660) );
  NAND U3680 ( .A(n1677), .B(n1678), .Z(n1676) );
  OR U3681 ( .A(n1679), .B(n1680), .Z(n1677) );
  NANDN U3682 ( .A(n1681), .B(n1679), .Z(n1675) );
  IV U3683 ( .A(n1680), .Z(n1681) );
  NAND U3684 ( .A(n1682), .B(n1683), .Z(n1657) );
  NAND U3685 ( .A(n1684), .B(n1685), .Z(n1683) );
  NANDN U3686 ( .A(n1686), .B(n1687), .Z(n1684) );
  NANDN U3687 ( .A(n1687), .B(n1686), .Z(n1682) );
  AND U3688 ( .A(n1688), .B(n1689), .Z(n1659) );
  NAND U3689 ( .A(n1690), .B(n1691), .Z(n1689) );
  OR U3690 ( .A(n1692), .B(n1693), .Z(n1690) );
  NANDN U3691 ( .A(n1694), .B(n1692), .Z(n1688) );
  NAND U3692 ( .A(n1695), .B(n1696), .Z(n1663) );
  NANDN U3693 ( .A(n1697), .B(n1698), .Z(n1696) );
  OR U3694 ( .A(n1699), .B(n1700), .Z(n1698) );
  NANDN U3695 ( .A(n1701), .B(n1699), .Z(n1695) );
  IV U3696 ( .A(n1700), .Z(n1701) );
  XNOR U3697 ( .A(n1671), .B(n1702), .Z(n1666) );
  XNOR U3698 ( .A(n1669), .B(n1672), .Z(n1702) );
  NAND U3699 ( .A(n1703), .B(n1704), .Z(n1672) );
  NAND U3700 ( .A(n1705), .B(n1706), .Z(n1704) );
  OR U3701 ( .A(n1707), .B(n1708), .Z(n1705) );
  NANDN U3702 ( .A(n1709), .B(n1707), .Z(n1703) );
  IV U3703 ( .A(n1708), .Z(n1709) );
  NAND U3704 ( .A(n1710), .B(n1711), .Z(n1669) );
  NAND U3705 ( .A(n1712), .B(n1713), .Z(n1711) );
  NANDN U3706 ( .A(n1714), .B(n1715), .Z(n1712) );
  NANDN U3707 ( .A(n1715), .B(n1714), .Z(n1710) );
  AND U3708 ( .A(n1716), .B(n1717), .Z(n1671) );
  NAND U3709 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U3710 ( .A(n1720), .B(n1721), .Z(n1718) );
  NANDN U3711 ( .A(n1722), .B(n1720), .Z(n1716) );
  XNOR U3712 ( .A(n1697), .B(n1723), .Z(N13662) );
  XOR U3713 ( .A(n1699), .B(n1700), .Z(n1723) );
  XNOR U3714 ( .A(n1713), .B(n1724), .Z(n1700) );
  XOR U3715 ( .A(n1714), .B(n1715), .Z(n1724) );
  XOR U3716 ( .A(n1720), .B(n1725), .Z(n1715) );
  XOR U3717 ( .A(n1719), .B(n1722), .Z(n1725) );
  IV U3718 ( .A(n1721), .Z(n1722) );
  NAND U3719 ( .A(n1726), .B(n1727), .Z(n1721) );
  OR U3720 ( .A(n1728), .B(n1729), .Z(n1727) );
  OR U3721 ( .A(n1730), .B(n1731), .Z(n1726) );
  NAND U3722 ( .A(n1732), .B(n1733), .Z(n1719) );
  OR U3723 ( .A(n1734), .B(n1735), .Z(n1733) );
  OR U3724 ( .A(n1736), .B(n1737), .Z(n1732) );
  NOR U3725 ( .A(n1738), .B(n1739), .Z(n1720) );
  ANDN U3726 ( .B(n1740), .A(n1741), .Z(n1714) );
  XNOR U3727 ( .A(n1707), .B(n1742), .Z(n1713) );
  XNOR U3728 ( .A(n1706), .B(n1708), .Z(n1742) );
  NAND U3729 ( .A(n1743), .B(n1744), .Z(n1708) );
  OR U3730 ( .A(n1745), .B(n1746), .Z(n1744) );
  OR U3731 ( .A(n1747), .B(n1748), .Z(n1743) );
  NAND U3732 ( .A(n1749), .B(n1750), .Z(n1706) );
  OR U3733 ( .A(n1751), .B(n1752), .Z(n1750) );
  OR U3734 ( .A(n1753), .B(n1754), .Z(n1749) );
  ANDN U3735 ( .B(n1755), .A(n1756), .Z(n1707) );
  IV U3736 ( .A(n1757), .Z(n1755) );
  ANDN U3737 ( .B(n1758), .A(n1759), .Z(n1699) );
  XOR U3738 ( .A(n1685), .B(n1760), .Z(n1697) );
  XOR U3739 ( .A(n1686), .B(n1687), .Z(n1760) );
  XOR U3740 ( .A(n1692), .B(n1761), .Z(n1687) );
  XOR U3741 ( .A(n1691), .B(n1694), .Z(n1761) );
  IV U3742 ( .A(n1693), .Z(n1694) );
  NAND U3743 ( .A(n1762), .B(n1763), .Z(n1693) );
  OR U3744 ( .A(n1764), .B(n1765), .Z(n1763) );
  OR U3745 ( .A(n1766), .B(n1767), .Z(n1762) );
  NAND U3746 ( .A(n1768), .B(n1769), .Z(n1691) );
  OR U3747 ( .A(n1770), .B(n1771), .Z(n1769) );
  OR U3748 ( .A(n1772), .B(n1773), .Z(n1768) );
  NOR U3749 ( .A(n1774), .B(n1775), .Z(n1692) );
  ANDN U3750 ( .B(n1776), .A(n1777), .Z(n1686) );
  IV U3751 ( .A(n1778), .Z(n1776) );
  XNOR U3752 ( .A(n1679), .B(n1779), .Z(n1685) );
  XNOR U3753 ( .A(n1678), .B(n1680), .Z(n1779) );
  NAND U3754 ( .A(n1780), .B(n1781), .Z(n1680) );
  OR U3755 ( .A(n1782), .B(n1783), .Z(n1781) );
  OR U3756 ( .A(n1784), .B(n1785), .Z(n1780) );
  NAND U3757 ( .A(n1786), .B(n1787), .Z(n1678) );
  OR U3758 ( .A(n1788), .B(n1789), .Z(n1787) );
  OR U3759 ( .A(n1790), .B(n1791), .Z(n1786) );
  ANDN U3760 ( .B(n1792), .A(n1793), .Z(n1679) );
  IV U3761 ( .A(n1794), .Z(n1792) );
  XNOR U3762 ( .A(n1759), .B(n1758), .Z(N13661) );
  XOR U3763 ( .A(n1778), .B(n1777), .Z(n1758) );
  XNOR U3764 ( .A(n1793), .B(n1794), .Z(n1777) );
  XNOR U3765 ( .A(n1788), .B(n1789), .Z(n1794) );
  XNOR U3766 ( .A(n1790), .B(n1791), .Z(n1789) );
  XNOR U3767 ( .A(y[1933]), .B(x[1933]), .Z(n1791) );
  XNOR U3768 ( .A(y[1934]), .B(x[1934]), .Z(n1790) );
  XNOR U3769 ( .A(y[1932]), .B(x[1932]), .Z(n1788) );
  XNOR U3770 ( .A(n1782), .B(n1783), .Z(n1793) );
  XNOR U3771 ( .A(y[1929]), .B(x[1929]), .Z(n1783) );
  XNOR U3772 ( .A(n1784), .B(n1785), .Z(n1782) );
  XNOR U3773 ( .A(y[1930]), .B(x[1930]), .Z(n1785) );
  XNOR U3774 ( .A(y[1931]), .B(x[1931]), .Z(n1784) );
  XNOR U3775 ( .A(n1775), .B(n1774), .Z(n1778) );
  XNOR U3776 ( .A(n1770), .B(n1771), .Z(n1774) );
  XNOR U3777 ( .A(y[1926]), .B(x[1926]), .Z(n1771) );
  XNOR U3778 ( .A(n1772), .B(n1773), .Z(n1770) );
  XNOR U3779 ( .A(y[1927]), .B(x[1927]), .Z(n1773) );
  XNOR U3780 ( .A(y[1928]), .B(x[1928]), .Z(n1772) );
  XNOR U3781 ( .A(n1764), .B(n1765), .Z(n1775) );
  XNOR U3782 ( .A(y[1923]), .B(x[1923]), .Z(n1765) );
  XNOR U3783 ( .A(n1766), .B(n1767), .Z(n1764) );
  XNOR U3784 ( .A(y[1924]), .B(x[1924]), .Z(n1767) );
  XNOR U3785 ( .A(y[1925]), .B(x[1925]), .Z(n1766) );
  XOR U3786 ( .A(n1740), .B(n1741), .Z(n1759) );
  XNOR U3787 ( .A(n1756), .B(n1757), .Z(n1741) );
  XNOR U3788 ( .A(n1751), .B(n1752), .Z(n1757) );
  XNOR U3789 ( .A(n1753), .B(n1754), .Z(n1752) );
  XNOR U3790 ( .A(y[1921]), .B(x[1921]), .Z(n1754) );
  XNOR U3791 ( .A(y[1922]), .B(x[1922]), .Z(n1753) );
  XNOR U3792 ( .A(y[1920]), .B(x[1920]), .Z(n1751) );
  XNOR U3793 ( .A(n1745), .B(n1746), .Z(n1756) );
  XNOR U3794 ( .A(y[1917]), .B(x[1917]), .Z(n1746) );
  XNOR U3795 ( .A(n1747), .B(n1748), .Z(n1745) );
  XNOR U3796 ( .A(y[1918]), .B(x[1918]), .Z(n1748) );
  XNOR U3797 ( .A(y[1919]), .B(x[1919]), .Z(n1747) );
  XOR U3798 ( .A(n1739), .B(n1738), .Z(n1740) );
  XNOR U3799 ( .A(n1734), .B(n1735), .Z(n1738) );
  XNOR U3800 ( .A(y[1914]), .B(x[1914]), .Z(n1735) );
  XNOR U3801 ( .A(n1736), .B(n1737), .Z(n1734) );
  XNOR U3802 ( .A(y[1915]), .B(x[1915]), .Z(n1737) );
  XNOR U3803 ( .A(y[1916]), .B(x[1916]), .Z(n1736) );
  XNOR U3804 ( .A(n1728), .B(n1729), .Z(n1739) );
  XNOR U3805 ( .A(y[1911]), .B(x[1911]), .Z(n1729) );
  XNOR U3806 ( .A(n1730), .B(n1731), .Z(n1728) );
  XNOR U3807 ( .A(y[1912]), .B(x[1912]), .Z(n1731) );
  XNOR U3808 ( .A(y[1913]), .B(x[1913]), .Z(n1730) );
  NAND U3809 ( .A(n1795), .B(n1796), .Z(N13654) );
  NANDN U3810 ( .A(n1797), .B(n1798), .Z(n1796) );
  OR U3811 ( .A(n1799), .B(n1800), .Z(n1798) );
  NAND U3812 ( .A(n1799), .B(n1800), .Z(n1795) );
  XOR U3813 ( .A(n1799), .B(n1801), .Z(N13653) );
  XNOR U3814 ( .A(n1797), .B(n1800), .Z(n1801) );
  AND U3815 ( .A(n1802), .B(n1803), .Z(n1800) );
  NANDN U3816 ( .A(n1804), .B(n1805), .Z(n1803) );
  NANDN U3817 ( .A(n1806), .B(n1807), .Z(n1805) );
  NANDN U3818 ( .A(n1807), .B(n1806), .Z(n1802) );
  NAND U3819 ( .A(n1808), .B(n1809), .Z(n1797) );
  NANDN U3820 ( .A(n1810), .B(n1811), .Z(n1809) );
  OR U3821 ( .A(n1812), .B(n1813), .Z(n1811) );
  NAND U3822 ( .A(n1813), .B(n1812), .Z(n1808) );
  AND U3823 ( .A(n1814), .B(n1815), .Z(n1799) );
  NANDN U3824 ( .A(n1816), .B(n1817), .Z(n1815) );
  NANDN U3825 ( .A(n1818), .B(n1819), .Z(n1817) );
  NANDN U3826 ( .A(n1819), .B(n1818), .Z(n1814) );
  XOR U3827 ( .A(n1813), .B(n1820), .Z(N13652) );
  XOR U3828 ( .A(n1810), .B(n1812), .Z(n1820) );
  XNOR U3829 ( .A(n1806), .B(n1821), .Z(n1812) );
  XNOR U3830 ( .A(n1804), .B(n1807), .Z(n1821) );
  NAND U3831 ( .A(n1822), .B(n1823), .Z(n1807) );
  NAND U3832 ( .A(n1824), .B(n1825), .Z(n1823) );
  OR U3833 ( .A(n1826), .B(n1827), .Z(n1824) );
  NANDN U3834 ( .A(n1828), .B(n1826), .Z(n1822) );
  IV U3835 ( .A(n1827), .Z(n1828) );
  NAND U3836 ( .A(n1829), .B(n1830), .Z(n1804) );
  NAND U3837 ( .A(n1831), .B(n1832), .Z(n1830) );
  NANDN U3838 ( .A(n1833), .B(n1834), .Z(n1831) );
  NANDN U3839 ( .A(n1834), .B(n1833), .Z(n1829) );
  AND U3840 ( .A(n1835), .B(n1836), .Z(n1806) );
  NAND U3841 ( .A(n1837), .B(n1838), .Z(n1836) );
  OR U3842 ( .A(n1839), .B(n1840), .Z(n1837) );
  NANDN U3843 ( .A(n1841), .B(n1839), .Z(n1835) );
  NAND U3844 ( .A(n1842), .B(n1843), .Z(n1810) );
  NANDN U3845 ( .A(n1844), .B(n1845), .Z(n1843) );
  OR U3846 ( .A(n1846), .B(n1847), .Z(n1845) );
  NANDN U3847 ( .A(n1848), .B(n1846), .Z(n1842) );
  IV U3848 ( .A(n1847), .Z(n1848) );
  XNOR U3849 ( .A(n1818), .B(n1849), .Z(n1813) );
  XNOR U3850 ( .A(n1816), .B(n1819), .Z(n1849) );
  NAND U3851 ( .A(n1850), .B(n1851), .Z(n1819) );
  NAND U3852 ( .A(n1852), .B(n1853), .Z(n1851) );
  OR U3853 ( .A(n1854), .B(n1855), .Z(n1852) );
  NANDN U3854 ( .A(n1856), .B(n1854), .Z(n1850) );
  IV U3855 ( .A(n1855), .Z(n1856) );
  NAND U3856 ( .A(n1857), .B(n1858), .Z(n1816) );
  NAND U3857 ( .A(n1859), .B(n1860), .Z(n1858) );
  NANDN U3858 ( .A(n1861), .B(n1862), .Z(n1859) );
  NANDN U3859 ( .A(n1862), .B(n1861), .Z(n1857) );
  AND U3860 ( .A(n1863), .B(n1864), .Z(n1818) );
  NAND U3861 ( .A(n1865), .B(n1866), .Z(n1864) );
  OR U3862 ( .A(n1867), .B(n1868), .Z(n1865) );
  NANDN U3863 ( .A(n1869), .B(n1867), .Z(n1863) );
  XNOR U3864 ( .A(n1844), .B(n1870), .Z(N13651) );
  XOR U3865 ( .A(n1846), .B(n1847), .Z(n1870) );
  XNOR U3866 ( .A(n1860), .B(n1871), .Z(n1847) );
  XOR U3867 ( .A(n1861), .B(n1862), .Z(n1871) );
  XOR U3868 ( .A(n1867), .B(n1872), .Z(n1862) );
  XOR U3869 ( .A(n1866), .B(n1869), .Z(n1872) );
  IV U3870 ( .A(n1868), .Z(n1869) );
  NAND U3871 ( .A(n1873), .B(n1874), .Z(n1868) );
  OR U3872 ( .A(n1875), .B(n1876), .Z(n1874) );
  OR U3873 ( .A(n1877), .B(n1878), .Z(n1873) );
  NAND U3874 ( .A(n1879), .B(n1880), .Z(n1866) );
  OR U3875 ( .A(n1881), .B(n1882), .Z(n1880) );
  OR U3876 ( .A(n1883), .B(n1884), .Z(n1879) );
  NOR U3877 ( .A(n1885), .B(n1886), .Z(n1867) );
  ANDN U3878 ( .B(n1887), .A(n1888), .Z(n1861) );
  XNOR U3879 ( .A(n1854), .B(n1889), .Z(n1860) );
  XNOR U3880 ( .A(n1853), .B(n1855), .Z(n1889) );
  NAND U3881 ( .A(n1890), .B(n1891), .Z(n1855) );
  OR U3882 ( .A(n1892), .B(n1893), .Z(n1891) );
  OR U3883 ( .A(n1894), .B(n1895), .Z(n1890) );
  NAND U3884 ( .A(n1896), .B(n1897), .Z(n1853) );
  OR U3885 ( .A(n1898), .B(n1899), .Z(n1897) );
  OR U3886 ( .A(n1900), .B(n1901), .Z(n1896) );
  ANDN U3887 ( .B(n1902), .A(n1903), .Z(n1854) );
  IV U3888 ( .A(n1904), .Z(n1902) );
  ANDN U3889 ( .B(n1905), .A(n1906), .Z(n1846) );
  XOR U3890 ( .A(n1832), .B(n1907), .Z(n1844) );
  XOR U3891 ( .A(n1833), .B(n1834), .Z(n1907) );
  XOR U3892 ( .A(n1839), .B(n1908), .Z(n1834) );
  XOR U3893 ( .A(n1838), .B(n1841), .Z(n1908) );
  IV U3894 ( .A(n1840), .Z(n1841) );
  NAND U3895 ( .A(n1909), .B(n1910), .Z(n1840) );
  OR U3896 ( .A(n1911), .B(n1912), .Z(n1910) );
  OR U3897 ( .A(n1913), .B(n1914), .Z(n1909) );
  NAND U3898 ( .A(n1915), .B(n1916), .Z(n1838) );
  OR U3899 ( .A(n1917), .B(n1918), .Z(n1916) );
  OR U3900 ( .A(n1919), .B(n1920), .Z(n1915) );
  NOR U3901 ( .A(n1921), .B(n1922), .Z(n1839) );
  ANDN U3902 ( .B(n1923), .A(n1924), .Z(n1833) );
  IV U3903 ( .A(n1925), .Z(n1923) );
  XNOR U3904 ( .A(n1826), .B(n1926), .Z(n1832) );
  XNOR U3905 ( .A(n1825), .B(n1827), .Z(n1926) );
  NAND U3906 ( .A(n1927), .B(n1928), .Z(n1827) );
  OR U3907 ( .A(n1929), .B(n1930), .Z(n1928) );
  OR U3908 ( .A(n1931), .B(n1932), .Z(n1927) );
  NAND U3909 ( .A(n1933), .B(n1934), .Z(n1825) );
  OR U3910 ( .A(n1935), .B(n1936), .Z(n1934) );
  OR U3911 ( .A(n1937), .B(n1938), .Z(n1933) );
  ANDN U3912 ( .B(n1939), .A(n1940), .Z(n1826) );
  IV U3913 ( .A(n1941), .Z(n1939) );
  XNOR U3914 ( .A(n1906), .B(n1905), .Z(N13650) );
  XOR U3915 ( .A(n1925), .B(n1924), .Z(n1905) );
  XNOR U3916 ( .A(n1940), .B(n1941), .Z(n1924) );
  XNOR U3917 ( .A(n1935), .B(n1936), .Z(n1941) );
  XNOR U3918 ( .A(n1937), .B(n1938), .Z(n1936) );
  XNOR U3919 ( .A(y[1909]), .B(x[1909]), .Z(n1938) );
  XNOR U3920 ( .A(y[1910]), .B(x[1910]), .Z(n1937) );
  XNOR U3921 ( .A(y[1908]), .B(x[1908]), .Z(n1935) );
  XNOR U3922 ( .A(n1929), .B(n1930), .Z(n1940) );
  XNOR U3923 ( .A(y[1905]), .B(x[1905]), .Z(n1930) );
  XNOR U3924 ( .A(n1931), .B(n1932), .Z(n1929) );
  XNOR U3925 ( .A(y[1906]), .B(x[1906]), .Z(n1932) );
  XNOR U3926 ( .A(y[1907]), .B(x[1907]), .Z(n1931) );
  XNOR U3927 ( .A(n1922), .B(n1921), .Z(n1925) );
  XNOR U3928 ( .A(n1917), .B(n1918), .Z(n1921) );
  XNOR U3929 ( .A(y[1902]), .B(x[1902]), .Z(n1918) );
  XNOR U3930 ( .A(n1919), .B(n1920), .Z(n1917) );
  XNOR U3931 ( .A(y[1903]), .B(x[1903]), .Z(n1920) );
  XNOR U3932 ( .A(y[1904]), .B(x[1904]), .Z(n1919) );
  XNOR U3933 ( .A(n1911), .B(n1912), .Z(n1922) );
  XNOR U3934 ( .A(y[1899]), .B(x[1899]), .Z(n1912) );
  XNOR U3935 ( .A(n1913), .B(n1914), .Z(n1911) );
  XNOR U3936 ( .A(y[1900]), .B(x[1900]), .Z(n1914) );
  XNOR U3937 ( .A(y[1901]), .B(x[1901]), .Z(n1913) );
  XOR U3938 ( .A(n1887), .B(n1888), .Z(n1906) );
  XNOR U3939 ( .A(n1903), .B(n1904), .Z(n1888) );
  XNOR U3940 ( .A(n1898), .B(n1899), .Z(n1904) );
  XNOR U3941 ( .A(n1900), .B(n1901), .Z(n1899) );
  XNOR U3942 ( .A(y[1897]), .B(x[1897]), .Z(n1901) );
  XNOR U3943 ( .A(y[1898]), .B(x[1898]), .Z(n1900) );
  XNOR U3944 ( .A(y[1896]), .B(x[1896]), .Z(n1898) );
  XNOR U3945 ( .A(n1892), .B(n1893), .Z(n1903) );
  XNOR U3946 ( .A(y[1893]), .B(x[1893]), .Z(n1893) );
  XNOR U3947 ( .A(n1894), .B(n1895), .Z(n1892) );
  XNOR U3948 ( .A(y[1894]), .B(x[1894]), .Z(n1895) );
  XNOR U3949 ( .A(y[1895]), .B(x[1895]), .Z(n1894) );
  XOR U3950 ( .A(n1886), .B(n1885), .Z(n1887) );
  XNOR U3951 ( .A(n1881), .B(n1882), .Z(n1885) );
  XNOR U3952 ( .A(y[1890]), .B(x[1890]), .Z(n1882) );
  XNOR U3953 ( .A(n1883), .B(n1884), .Z(n1881) );
  XNOR U3954 ( .A(y[1891]), .B(x[1891]), .Z(n1884) );
  XNOR U3955 ( .A(y[1892]), .B(x[1892]), .Z(n1883) );
  XNOR U3956 ( .A(n1875), .B(n1876), .Z(n1886) );
  XNOR U3957 ( .A(y[1887]), .B(x[1887]), .Z(n1876) );
  XNOR U3958 ( .A(n1877), .B(n1878), .Z(n1875) );
  XNOR U3959 ( .A(y[1888]), .B(x[1888]), .Z(n1878) );
  XNOR U3960 ( .A(y[1889]), .B(x[1889]), .Z(n1877) );
  NAND U3961 ( .A(n1942), .B(n1943), .Z(N13643) );
  NANDN U3962 ( .A(n1944), .B(n1945), .Z(n1943) );
  OR U3963 ( .A(n1946), .B(n1947), .Z(n1945) );
  NAND U3964 ( .A(n1946), .B(n1947), .Z(n1942) );
  XOR U3965 ( .A(n1946), .B(n1948), .Z(N13642) );
  XNOR U3966 ( .A(n1944), .B(n1947), .Z(n1948) );
  AND U3967 ( .A(n1949), .B(n1950), .Z(n1947) );
  NANDN U3968 ( .A(n1951), .B(n1952), .Z(n1950) );
  NANDN U3969 ( .A(n1953), .B(n1954), .Z(n1952) );
  NANDN U3970 ( .A(n1954), .B(n1953), .Z(n1949) );
  NAND U3971 ( .A(n1955), .B(n1956), .Z(n1944) );
  NANDN U3972 ( .A(n1957), .B(n1958), .Z(n1956) );
  OR U3973 ( .A(n1959), .B(n1960), .Z(n1958) );
  NAND U3974 ( .A(n1960), .B(n1959), .Z(n1955) );
  AND U3975 ( .A(n1961), .B(n1962), .Z(n1946) );
  NANDN U3976 ( .A(n1963), .B(n1964), .Z(n1962) );
  NANDN U3977 ( .A(n1965), .B(n1966), .Z(n1964) );
  NANDN U3978 ( .A(n1966), .B(n1965), .Z(n1961) );
  XOR U3979 ( .A(n1960), .B(n1967), .Z(N13641) );
  XOR U3980 ( .A(n1957), .B(n1959), .Z(n1967) );
  XNOR U3981 ( .A(n1953), .B(n1968), .Z(n1959) );
  XNOR U3982 ( .A(n1951), .B(n1954), .Z(n1968) );
  NAND U3983 ( .A(n1969), .B(n1970), .Z(n1954) );
  NAND U3984 ( .A(n1971), .B(n1972), .Z(n1970) );
  OR U3985 ( .A(n1973), .B(n1974), .Z(n1971) );
  NANDN U3986 ( .A(n1975), .B(n1973), .Z(n1969) );
  IV U3987 ( .A(n1974), .Z(n1975) );
  NAND U3988 ( .A(n1976), .B(n1977), .Z(n1951) );
  NAND U3989 ( .A(n1978), .B(n1979), .Z(n1977) );
  NANDN U3990 ( .A(n1980), .B(n1981), .Z(n1978) );
  NANDN U3991 ( .A(n1981), .B(n1980), .Z(n1976) );
  AND U3992 ( .A(n1982), .B(n1983), .Z(n1953) );
  NAND U3993 ( .A(n1984), .B(n1985), .Z(n1983) );
  OR U3994 ( .A(n1986), .B(n1987), .Z(n1984) );
  NANDN U3995 ( .A(n1988), .B(n1986), .Z(n1982) );
  NAND U3996 ( .A(n1989), .B(n1990), .Z(n1957) );
  NANDN U3997 ( .A(n1991), .B(n1992), .Z(n1990) );
  OR U3998 ( .A(n1993), .B(n1994), .Z(n1992) );
  NANDN U3999 ( .A(n1995), .B(n1993), .Z(n1989) );
  IV U4000 ( .A(n1994), .Z(n1995) );
  XNOR U4001 ( .A(n1965), .B(n1996), .Z(n1960) );
  XNOR U4002 ( .A(n1963), .B(n1966), .Z(n1996) );
  NAND U4003 ( .A(n1997), .B(n1998), .Z(n1966) );
  NAND U4004 ( .A(n1999), .B(n2000), .Z(n1998) );
  OR U4005 ( .A(n2001), .B(n2002), .Z(n1999) );
  NANDN U4006 ( .A(n2003), .B(n2001), .Z(n1997) );
  IV U4007 ( .A(n2002), .Z(n2003) );
  NAND U4008 ( .A(n2004), .B(n2005), .Z(n1963) );
  NAND U4009 ( .A(n2006), .B(n2007), .Z(n2005) );
  NANDN U4010 ( .A(n2008), .B(n2009), .Z(n2006) );
  NANDN U4011 ( .A(n2009), .B(n2008), .Z(n2004) );
  AND U4012 ( .A(n2010), .B(n2011), .Z(n1965) );
  NAND U4013 ( .A(n2012), .B(n2013), .Z(n2011) );
  OR U4014 ( .A(n2014), .B(n2015), .Z(n2012) );
  NANDN U4015 ( .A(n2016), .B(n2014), .Z(n2010) );
  XNOR U4016 ( .A(n1991), .B(n2017), .Z(N13640) );
  XOR U4017 ( .A(n1993), .B(n1994), .Z(n2017) );
  XNOR U4018 ( .A(n2007), .B(n2018), .Z(n1994) );
  XOR U4019 ( .A(n2008), .B(n2009), .Z(n2018) );
  XOR U4020 ( .A(n2014), .B(n2019), .Z(n2009) );
  XOR U4021 ( .A(n2013), .B(n2016), .Z(n2019) );
  IV U4022 ( .A(n2015), .Z(n2016) );
  NAND U4023 ( .A(n2020), .B(n2021), .Z(n2015) );
  OR U4024 ( .A(n2022), .B(n2023), .Z(n2021) );
  OR U4025 ( .A(n2024), .B(n2025), .Z(n2020) );
  NAND U4026 ( .A(n2026), .B(n2027), .Z(n2013) );
  OR U4027 ( .A(n2028), .B(n2029), .Z(n2027) );
  OR U4028 ( .A(n2030), .B(n2031), .Z(n2026) );
  NOR U4029 ( .A(n2032), .B(n2033), .Z(n2014) );
  ANDN U4030 ( .B(n2034), .A(n2035), .Z(n2008) );
  XNOR U4031 ( .A(n2001), .B(n2036), .Z(n2007) );
  XNOR U4032 ( .A(n2000), .B(n2002), .Z(n2036) );
  NAND U4033 ( .A(n2037), .B(n2038), .Z(n2002) );
  OR U4034 ( .A(n2039), .B(n2040), .Z(n2038) );
  OR U4035 ( .A(n2041), .B(n2042), .Z(n2037) );
  NAND U4036 ( .A(n2043), .B(n2044), .Z(n2000) );
  OR U4037 ( .A(n2045), .B(n2046), .Z(n2044) );
  OR U4038 ( .A(n2047), .B(n2048), .Z(n2043) );
  ANDN U4039 ( .B(n2049), .A(n2050), .Z(n2001) );
  IV U4040 ( .A(n2051), .Z(n2049) );
  ANDN U4041 ( .B(n2052), .A(n2053), .Z(n1993) );
  XOR U4042 ( .A(n1979), .B(n2054), .Z(n1991) );
  XOR U4043 ( .A(n1980), .B(n1981), .Z(n2054) );
  XOR U4044 ( .A(n1986), .B(n2055), .Z(n1981) );
  XOR U4045 ( .A(n1985), .B(n1988), .Z(n2055) );
  IV U4046 ( .A(n1987), .Z(n1988) );
  NAND U4047 ( .A(n2056), .B(n2057), .Z(n1987) );
  OR U4048 ( .A(n2058), .B(n2059), .Z(n2057) );
  OR U4049 ( .A(n2060), .B(n2061), .Z(n2056) );
  NAND U4050 ( .A(n2062), .B(n2063), .Z(n1985) );
  OR U4051 ( .A(n2064), .B(n2065), .Z(n2063) );
  OR U4052 ( .A(n2066), .B(n2067), .Z(n2062) );
  NOR U4053 ( .A(n2068), .B(n2069), .Z(n1986) );
  ANDN U4054 ( .B(n2070), .A(n2071), .Z(n1980) );
  IV U4055 ( .A(n2072), .Z(n2070) );
  XNOR U4056 ( .A(n1973), .B(n2073), .Z(n1979) );
  XNOR U4057 ( .A(n1972), .B(n1974), .Z(n2073) );
  NAND U4058 ( .A(n2074), .B(n2075), .Z(n1974) );
  OR U4059 ( .A(n2076), .B(n2077), .Z(n2075) );
  OR U4060 ( .A(n2078), .B(n2079), .Z(n2074) );
  NAND U4061 ( .A(n2080), .B(n2081), .Z(n1972) );
  OR U4062 ( .A(n2082), .B(n2083), .Z(n2081) );
  OR U4063 ( .A(n2084), .B(n2085), .Z(n2080) );
  ANDN U4064 ( .B(n2086), .A(n2087), .Z(n1973) );
  IV U4065 ( .A(n2088), .Z(n2086) );
  XNOR U4066 ( .A(n2053), .B(n2052), .Z(N13639) );
  XOR U4067 ( .A(n2072), .B(n2071), .Z(n2052) );
  XNOR U4068 ( .A(n2087), .B(n2088), .Z(n2071) );
  XNOR U4069 ( .A(n2082), .B(n2083), .Z(n2088) );
  XNOR U4070 ( .A(n2084), .B(n2085), .Z(n2083) );
  XNOR U4071 ( .A(y[1885]), .B(x[1885]), .Z(n2085) );
  XNOR U4072 ( .A(y[1886]), .B(x[1886]), .Z(n2084) );
  XNOR U4073 ( .A(y[1884]), .B(x[1884]), .Z(n2082) );
  XNOR U4074 ( .A(n2076), .B(n2077), .Z(n2087) );
  XNOR U4075 ( .A(y[1881]), .B(x[1881]), .Z(n2077) );
  XNOR U4076 ( .A(n2078), .B(n2079), .Z(n2076) );
  XNOR U4077 ( .A(y[1882]), .B(x[1882]), .Z(n2079) );
  XNOR U4078 ( .A(y[1883]), .B(x[1883]), .Z(n2078) );
  XNOR U4079 ( .A(n2069), .B(n2068), .Z(n2072) );
  XNOR U4080 ( .A(n2064), .B(n2065), .Z(n2068) );
  XNOR U4081 ( .A(y[1878]), .B(x[1878]), .Z(n2065) );
  XNOR U4082 ( .A(n2066), .B(n2067), .Z(n2064) );
  XNOR U4083 ( .A(y[1879]), .B(x[1879]), .Z(n2067) );
  XNOR U4084 ( .A(y[1880]), .B(x[1880]), .Z(n2066) );
  XNOR U4085 ( .A(n2058), .B(n2059), .Z(n2069) );
  XNOR U4086 ( .A(y[1875]), .B(x[1875]), .Z(n2059) );
  XNOR U4087 ( .A(n2060), .B(n2061), .Z(n2058) );
  XNOR U4088 ( .A(y[1876]), .B(x[1876]), .Z(n2061) );
  XNOR U4089 ( .A(y[1877]), .B(x[1877]), .Z(n2060) );
  XOR U4090 ( .A(n2034), .B(n2035), .Z(n2053) );
  XNOR U4091 ( .A(n2050), .B(n2051), .Z(n2035) );
  XNOR U4092 ( .A(n2045), .B(n2046), .Z(n2051) );
  XNOR U4093 ( .A(n2047), .B(n2048), .Z(n2046) );
  XNOR U4094 ( .A(y[1873]), .B(x[1873]), .Z(n2048) );
  XNOR U4095 ( .A(y[1874]), .B(x[1874]), .Z(n2047) );
  XNOR U4096 ( .A(y[1872]), .B(x[1872]), .Z(n2045) );
  XNOR U4097 ( .A(n2039), .B(n2040), .Z(n2050) );
  XNOR U4098 ( .A(y[1869]), .B(x[1869]), .Z(n2040) );
  XNOR U4099 ( .A(n2041), .B(n2042), .Z(n2039) );
  XNOR U4100 ( .A(y[1870]), .B(x[1870]), .Z(n2042) );
  XNOR U4101 ( .A(y[1871]), .B(x[1871]), .Z(n2041) );
  XOR U4102 ( .A(n2033), .B(n2032), .Z(n2034) );
  XNOR U4103 ( .A(n2028), .B(n2029), .Z(n2032) );
  XNOR U4104 ( .A(y[1866]), .B(x[1866]), .Z(n2029) );
  XNOR U4105 ( .A(n2030), .B(n2031), .Z(n2028) );
  XNOR U4106 ( .A(y[1867]), .B(x[1867]), .Z(n2031) );
  XNOR U4107 ( .A(y[1868]), .B(x[1868]), .Z(n2030) );
  XNOR U4108 ( .A(n2022), .B(n2023), .Z(n2033) );
  XNOR U4109 ( .A(y[1863]), .B(x[1863]), .Z(n2023) );
  XNOR U4110 ( .A(n2024), .B(n2025), .Z(n2022) );
  XNOR U4111 ( .A(y[1864]), .B(x[1864]), .Z(n2025) );
  XNOR U4112 ( .A(y[1865]), .B(x[1865]), .Z(n2024) );
  NAND U4113 ( .A(n2089), .B(n2090), .Z(N13632) );
  NANDN U4114 ( .A(n2091), .B(n2092), .Z(n2090) );
  OR U4115 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U4116 ( .A(n2093), .B(n2094), .Z(n2089) );
  XOR U4117 ( .A(n2093), .B(n2095), .Z(N13631) );
  XNOR U4118 ( .A(n2091), .B(n2094), .Z(n2095) );
  AND U4119 ( .A(n2096), .B(n2097), .Z(n2094) );
  NANDN U4120 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U4121 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U4122 ( .A(n2101), .B(n2100), .Z(n2096) );
  NAND U4123 ( .A(n2102), .B(n2103), .Z(n2091) );
  NANDN U4124 ( .A(n2104), .B(n2105), .Z(n2103) );
  OR U4125 ( .A(n2106), .B(n2107), .Z(n2105) );
  NAND U4126 ( .A(n2107), .B(n2106), .Z(n2102) );
  AND U4127 ( .A(n2108), .B(n2109), .Z(n2093) );
  NANDN U4128 ( .A(n2110), .B(n2111), .Z(n2109) );
  NANDN U4129 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U4130 ( .A(n2113), .B(n2112), .Z(n2108) );
  XOR U4131 ( .A(n2107), .B(n2114), .Z(N13630) );
  XOR U4132 ( .A(n2104), .B(n2106), .Z(n2114) );
  XNOR U4133 ( .A(n2100), .B(n2115), .Z(n2106) );
  XNOR U4134 ( .A(n2098), .B(n2101), .Z(n2115) );
  NAND U4135 ( .A(n2116), .B(n2117), .Z(n2101) );
  NAND U4136 ( .A(n2118), .B(n2119), .Z(n2117) );
  OR U4137 ( .A(n2120), .B(n2121), .Z(n2118) );
  NANDN U4138 ( .A(n2122), .B(n2120), .Z(n2116) );
  IV U4139 ( .A(n2121), .Z(n2122) );
  NAND U4140 ( .A(n2123), .B(n2124), .Z(n2098) );
  NAND U4141 ( .A(n2125), .B(n2126), .Z(n2124) );
  NANDN U4142 ( .A(n2127), .B(n2128), .Z(n2125) );
  NANDN U4143 ( .A(n2128), .B(n2127), .Z(n2123) );
  AND U4144 ( .A(n2129), .B(n2130), .Z(n2100) );
  NAND U4145 ( .A(n2131), .B(n2132), .Z(n2130) );
  OR U4146 ( .A(n2133), .B(n2134), .Z(n2131) );
  NANDN U4147 ( .A(n2135), .B(n2133), .Z(n2129) );
  NAND U4148 ( .A(n2136), .B(n2137), .Z(n2104) );
  NANDN U4149 ( .A(n2138), .B(n2139), .Z(n2137) );
  OR U4150 ( .A(n2140), .B(n2141), .Z(n2139) );
  NANDN U4151 ( .A(n2142), .B(n2140), .Z(n2136) );
  IV U4152 ( .A(n2141), .Z(n2142) );
  XNOR U4153 ( .A(n2112), .B(n2143), .Z(n2107) );
  XNOR U4154 ( .A(n2110), .B(n2113), .Z(n2143) );
  NAND U4155 ( .A(n2144), .B(n2145), .Z(n2113) );
  NAND U4156 ( .A(n2146), .B(n2147), .Z(n2145) );
  OR U4157 ( .A(n2148), .B(n2149), .Z(n2146) );
  NANDN U4158 ( .A(n2150), .B(n2148), .Z(n2144) );
  IV U4159 ( .A(n2149), .Z(n2150) );
  NAND U4160 ( .A(n2151), .B(n2152), .Z(n2110) );
  NAND U4161 ( .A(n2153), .B(n2154), .Z(n2152) );
  NANDN U4162 ( .A(n2155), .B(n2156), .Z(n2153) );
  NANDN U4163 ( .A(n2156), .B(n2155), .Z(n2151) );
  AND U4164 ( .A(n2157), .B(n2158), .Z(n2112) );
  NAND U4165 ( .A(n2159), .B(n2160), .Z(n2158) );
  OR U4166 ( .A(n2161), .B(n2162), .Z(n2159) );
  NANDN U4167 ( .A(n2163), .B(n2161), .Z(n2157) );
  XNOR U4168 ( .A(n2138), .B(n2164), .Z(N13629) );
  XOR U4169 ( .A(n2140), .B(n2141), .Z(n2164) );
  XNOR U4170 ( .A(n2154), .B(n2165), .Z(n2141) );
  XOR U4171 ( .A(n2155), .B(n2156), .Z(n2165) );
  XOR U4172 ( .A(n2161), .B(n2166), .Z(n2156) );
  XOR U4173 ( .A(n2160), .B(n2163), .Z(n2166) );
  IV U4174 ( .A(n2162), .Z(n2163) );
  NAND U4175 ( .A(n2167), .B(n2168), .Z(n2162) );
  OR U4176 ( .A(n2169), .B(n2170), .Z(n2168) );
  OR U4177 ( .A(n2171), .B(n2172), .Z(n2167) );
  NAND U4178 ( .A(n2173), .B(n2174), .Z(n2160) );
  OR U4179 ( .A(n2175), .B(n2176), .Z(n2174) );
  OR U4180 ( .A(n2177), .B(n2178), .Z(n2173) );
  NOR U4181 ( .A(n2179), .B(n2180), .Z(n2161) );
  ANDN U4182 ( .B(n2181), .A(n2182), .Z(n2155) );
  XNOR U4183 ( .A(n2148), .B(n2183), .Z(n2154) );
  XNOR U4184 ( .A(n2147), .B(n2149), .Z(n2183) );
  NAND U4185 ( .A(n2184), .B(n2185), .Z(n2149) );
  OR U4186 ( .A(n2186), .B(n2187), .Z(n2185) );
  OR U4187 ( .A(n2188), .B(n2189), .Z(n2184) );
  NAND U4188 ( .A(n2190), .B(n2191), .Z(n2147) );
  OR U4189 ( .A(n2192), .B(n2193), .Z(n2191) );
  OR U4190 ( .A(n2194), .B(n2195), .Z(n2190) );
  ANDN U4191 ( .B(n2196), .A(n2197), .Z(n2148) );
  IV U4192 ( .A(n2198), .Z(n2196) );
  ANDN U4193 ( .B(n2199), .A(n2200), .Z(n2140) );
  XOR U4194 ( .A(n2126), .B(n2201), .Z(n2138) );
  XOR U4195 ( .A(n2127), .B(n2128), .Z(n2201) );
  XOR U4196 ( .A(n2133), .B(n2202), .Z(n2128) );
  XOR U4197 ( .A(n2132), .B(n2135), .Z(n2202) );
  IV U4198 ( .A(n2134), .Z(n2135) );
  NAND U4199 ( .A(n2203), .B(n2204), .Z(n2134) );
  OR U4200 ( .A(n2205), .B(n2206), .Z(n2204) );
  OR U4201 ( .A(n2207), .B(n2208), .Z(n2203) );
  NAND U4202 ( .A(n2209), .B(n2210), .Z(n2132) );
  OR U4203 ( .A(n2211), .B(n2212), .Z(n2210) );
  OR U4204 ( .A(n2213), .B(n2214), .Z(n2209) );
  NOR U4205 ( .A(n2215), .B(n2216), .Z(n2133) );
  ANDN U4206 ( .B(n2217), .A(n2218), .Z(n2127) );
  IV U4207 ( .A(n2219), .Z(n2217) );
  XNOR U4208 ( .A(n2120), .B(n2220), .Z(n2126) );
  XNOR U4209 ( .A(n2119), .B(n2121), .Z(n2220) );
  NAND U4210 ( .A(n2221), .B(n2222), .Z(n2121) );
  OR U4211 ( .A(n2223), .B(n2224), .Z(n2222) );
  OR U4212 ( .A(n2225), .B(n2226), .Z(n2221) );
  NAND U4213 ( .A(n2227), .B(n2228), .Z(n2119) );
  OR U4214 ( .A(n2229), .B(n2230), .Z(n2228) );
  OR U4215 ( .A(n2231), .B(n2232), .Z(n2227) );
  ANDN U4216 ( .B(n2233), .A(n2234), .Z(n2120) );
  IV U4217 ( .A(n2235), .Z(n2233) );
  XNOR U4218 ( .A(n2200), .B(n2199), .Z(N13628) );
  XOR U4219 ( .A(n2219), .B(n2218), .Z(n2199) );
  XNOR U4220 ( .A(n2234), .B(n2235), .Z(n2218) );
  XNOR U4221 ( .A(n2229), .B(n2230), .Z(n2235) );
  XNOR U4222 ( .A(n2231), .B(n2232), .Z(n2230) );
  XNOR U4223 ( .A(y[1861]), .B(x[1861]), .Z(n2232) );
  XNOR U4224 ( .A(y[1862]), .B(x[1862]), .Z(n2231) );
  XNOR U4225 ( .A(y[1860]), .B(x[1860]), .Z(n2229) );
  XNOR U4226 ( .A(n2223), .B(n2224), .Z(n2234) );
  XNOR U4227 ( .A(y[1857]), .B(x[1857]), .Z(n2224) );
  XNOR U4228 ( .A(n2225), .B(n2226), .Z(n2223) );
  XNOR U4229 ( .A(y[1858]), .B(x[1858]), .Z(n2226) );
  XNOR U4230 ( .A(y[1859]), .B(x[1859]), .Z(n2225) );
  XNOR U4231 ( .A(n2216), .B(n2215), .Z(n2219) );
  XNOR U4232 ( .A(n2211), .B(n2212), .Z(n2215) );
  XNOR U4233 ( .A(y[1854]), .B(x[1854]), .Z(n2212) );
  XNOR U4234 ( .A(n2213), .B(n2214), .Z(n2211) );
  XNOR U4235 ( .A(y[1855]), .B(x[1855]), .Z(n2214) );
  XNOR U4236 ( .A(y[1856]), .B(x[1856]), .Z(n2213) );
  XNOR U4237 ( .A(n2205), .B(n2206), .Z(n2216) );
  XNOR U4238 ( .A(y[1851]), .B(x[1851]), .Z(n2206) );
  XNOR U4239 ( .A(n2207), .B(n2208), .Z(n2205) );
  XNOR U4240 ( .A(y[1852]), .B(x[1852]), .Z(n2208) );
  XNOR U4241 ( .A(y[1853]), .B(x[1853]), .Z(n2207) );
  XOR U4242 ( .A(n2181), .B(n2182), .Z(n2200) );
  XNOR U4243 ( .A(n2197), .B(n2198), .Z(n2182) );
  XNOR U4244 ( .A(n2192), .B(n2193), .Z(n2198) );
  XNOR U4245 ( .A(n2194), .B(n2195), .Z(n2193) );
  XNOR U4246 ( .A(y[1849]), .B(x[1849]), .Z(n2195) );
  XNOR U4247 ( .A(y[1850]), .B(x[1850]), .Z(n2194) );
  XNOR U4248 ( .A(y[1848]), .B(x[1848]), .Z(n2192) );
  XNOR U4249 ( .A(n2186), .B(n2187), .Z(n2197) );
  XNOR U4250 ( .A(y[1845]), .B(x[1845]), .Z(n2187) );
  XNOR U4251 ( .A(n2188), .B(n2189), .Z(n2186) );
  XNOR U4252 ( .A(y[1846]), .B(x[1846]), .Z(n2189) );
  XNOR U4253 ( .A(y[1847]), .B(x[1847]), .Z(n2188) );
  XOR U4254 ( .A(n2180), .B(n2179), .Z(n2181) );
  XNOR U4255 ( .A(n2175), .B(n2176), .Z(n2179) );
  XNOR U4256 ( .A(y[1842]), .B(x[1842]), .Z(n2176) );
  XNOR U4257 ( .A(n2177), .B(n2178), .Z(n2175) );
  XNOR U4258 ( .A(y[1843]), .B(x[1843]), .Z(n2178) );
  XNOR U4259 ( .A(y[1844]), .B(x[1844]), .Z(n2177) );
  XNOR U4260 ( .A(n2169), .B(n2170), .Z(n2180) );
  XNOR U4261 ( .A(y[1839]), .B(x[1839]), .Z(n2170) );
  XNOR U4262 ( .A(n2171), .B(n2172), .Z(n2169) );
  XNOR U4263 ( .A(y[1840]), .B(x[1840]), .Z(n2172) );
  XNOR U4264 ( .A(y[1841]), .B(x[1841]), .Z(n2171) );
  NAND U4265 ( .A(n2236), .B(n2237), .Z(N13621) );
  NANDN U4266 ( .A(n2238), .B(n2239), .Z(n2237) );
  OR U4267 ( .A(n2240), .B(n2241), .Z(n2239) );
  NAND U4268 ( .A(n2240), .B(n2241), .Z(n2236) );
  XOR U4269 ( .A(n2240), .B(n2242), .Z(N13620) );
  XNOR U4270 ( .A(n2238), .B(n2241), .Z(n2242) );
  AND U4271 ( .A(n2243), .B(n2244), .Z(n2241) );
  NANDN U4272 ( .A(n2245), .B(n2246), .Z(n2244) );
  NANDN U4273 ( .A(n2247), .B(n2248), .Z(n2246) );
  NANDN U4274 ( .A(n2248), .B(n2247), .Z(n2243) );
  NAND U4275 ( .A(n2249), .B(n2250), .Z(n2238) );
  NANDN U4276 ( .A(n2251), .B(n2252), .Z(n2250) );
  OR U4277 ( .A(n2253), .B(n2254), .Z(n2252) );
  NAND U4278 ( .A(n2254), .B(n2253), .Z(n2249) );
  AND U4279 ( .A(n2255), .B(n2256), .Z(n2240) );
  NANDN U4280 ( .A(n2257), .B(n2258), .Z(n2256) );
  NANDN U4281 ( .A(n2259), .B(n2260), .Z(n2258) );
  NANDN U4282 ( .A(n2260), .B(n2259), .Z(n2255) );
  XOR U4283 ( .A(n2254), .B(n2261), .Z(N13619) );
  XOR U4284 ( .A(n2251), .B(n2253), .Z(n2261) );
  XNOR U4285 ( .A(n2247), .B(n2262), .Z(n2253) );
  XNOR U4286 ( .A(n2245), .B(n2248), .Z(n2262) );
  NAND U4287 ( .A(n2263), .B(n2264), .Z(n2248) );
  NAND U4288 ( .A(n2265), .B(n2266), .Z(n2264) );
  OR U4289 ( .A(n2267), .B(n2268), .Z(n2265) );
  NANDN U4290 ( .A(n2269), .B(n2267), .Z(n2263) );
  IV U4291 ( .A(n2268), .Z(n2269) );
  NAND U4292 ( .A(n2270), .B(n2271), .Z(n2245) );
  NAND U4293 ( .A(n2272), .B(n2273), .Z(n2271) );
  NANDN U4294 ( .A(n2274), .B(n2275), .Z(n2272) );
  NANDN U4295 ( .A(n2275), .B(n2274), .Z(n2270) );
  AND U4296 ( .A(n2276), .B(n2277), .Z(n2247) );
  NAND U4297 ( .A(n2278), .B(n2279), .Z(n2277) );
  OR U4298 ( .A(n2280), .B(n2281), .Z(n2278) );
  NANDN U4299 ( .A(n2282), .B(n2280), .Z(n2276) );
  NAND U4300 ( .A(n2283), .B(n2284), .Z(n2251) );
  NANDN U4301 ( .A(n2285), .B(n2286), .Z(n2284) );
  OR U4302 ( .A(n2287), .B(n2288), .Z(n2286) );
  NANDN U4303 ( .A(n2289), .B(n2287), .Z(n2283) );
  IV U4304 ( .A(n2288), .Z(n2289) );
  XNOR U4305 ( .A(n2259), .B(n2290), .Z(n2254) );
  XNOR U4306 ( .A(n2257), .B(n2260), .Z(n2290) );
  NAND U4307 ( .A(n2291), .B(n2292), .Z(n2260) );
  NAND U4308 ( .A(n2293), .B(n2294), .Z(n2292) );
  OR U4309 ( .A(n2295), .B(n2296), .Z(n2293) );
  NANDN U4310 ( .A(n2297), .B(n2295), .Z(n2291) );
  IV U4311 ( .A(n2296), .Z(n2297) );
  NAND U4312 ( .A(n2298), .B(n2299), .Z(n2257) );
  NAND U4313 ( .A(n2300), .B(n2301), .Z(n2299) );
  NANDN U4314 ( .A(n2302), .B(n2303), .Z(n2300) );
  NANDN U4315 ( .A(n2303), .B(n2302), .Z(n2298) );
  AND U4316 ( .A(n2304), .B(n2305), .Z(n2259) );
  NAND U4317 ( .A(n2306), .B(n2307), .Z(n2305) );
  OR U4318 ( .A(n2308), .B(n2309), .Z(n2306) );
  NANDN U4319 ( .A(n2310), .B(n2308), .Z(n2304) );
  XNOR U4320 ( .A(n2285), .B(n2311), .Z(N13618) );
  XOR U4321 ( .A(n2287), .B(n2288), .Z(n2311) );
  XNOR U4322 ( .A(n2301), .B(n2312), .Z(n2288) );
  XOR U4323 ( .A(n2302), .B(n2303), .Z(n2312) );
  XOR U4324 ( .A(n2308), .B(n2313), .Z(n2303) );
  XOR U4325 ( .A(n2307), .B(n2310), .Z(n2313) );
  IV U4326 ( .A(n2309), .Z(n2310) );
  NAND U4327 ( .A(n2314), .B(n2315), .Z(n2309) );
  OR U4328 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U4329 ( .A(n2318), .B(n2319), .Z(n2314) );
  NAND U4330 ( .A(n2320), .B(n2321), .Z(n2307) );
  OR U4331 ( .A(n2322), .B(n2323), .Z(n2321) );
  OR U4332 ( .A(n2324), .B(n2325), .Z(n2320) );
  NOR U4333 ( .A(n2326), .B(n2327), .Z(n2308) );
  ANDN U4334 ( .B(n2328), .A(n2329), .Z(n2302) );
  XNOR U4335 ( .A(n2295), .B(n2330), .Z(n2301) );
  XNOR U4336 ( .A(n2294), .B(n2296), .Z(n2330) );
  NAND U4337 ( .A(n2331), .B(n2332), .Z(n2296) );
  OR U4338 ( .A(n2333), .B(n2334), .Z(n2332) );
  OR U4339 ( .A(n2335), .B(n2336), .Z(n2331) );
  NAND U4340 ( .A(n2337), .B(n2338), .Z(n2294) );
  OR U4341 ( .A(n2339), .B(n2340), .Z(n2338) );
  OR U4342 ( .A(n2341), .B(n2342), .Z(n2337) );
  ANDN U4343 ( .B(n2343), .A(n2344), .Z(n2295) );
  IV U4344 ( .A(n2345), .Z(n2343) );
  ANDN U4345 ( .B(n2346), .A(n2347), .Z(n2287) );
  XOR U4346 ( .A(n2273), .B(n2348), .Z(n2285) );
  XOR U4347 ( .A(n2274), .B(n2275), .Z(n2348) );
  XOR U4348 ( .A(n2280), .B(n2349), .Z(n2275) );
  XOR U4349 ( .A(n2279), .B(n2282), .Z(n2349) );
  IV U4350 ( .A(n2281), .Z(n2282) );
  NAND U4351 ( .A(n2350), .B(n2351), .Z(n2281) );
  OR U4352 ( .A(n2352), .B(n2353), .Z(n2351) );
  OR U4353 ( .A(n2354), .B(n2355), .Z(n2350) );
  NAND U4354 ( .A(n2356), .B(n2357), .Z(n2279) );
  OR U4355 ( .A(n2358), .B(n2359), .Z(n2357) );
  OR U4356 ( .A(n2360), .B(n2361), .Z(n2356) );
  NOR U4357 ( .A(n2362), .B(n2363), .Z(n2280) );
  ANDN U4358 ( .B(n2364), .A(n2365), .Z(n2274) );
  IV U4359 ( .A(n2366), .Z(n2364) );
  XNOR U4360 ( .A(n2267), .B(n2367), .Z(n2273) );
  XNOR U4361 ( .A(n2266), .B(n2268), .Z(n2367) );
  NAND U4362 ( .A(n2368), .B(n2369), .Z(n2268) );
  OR U4363 ( .A(n2370), .B(n2371), .Z(n2369) );
  OR U4364 ( .A(n2372), .B(n2373), .Z(n2368) );
  NAND U4365 ( .A(n2374), .B(n2375), .Z(n2266) );
  OR U4366 ( .A(n2376), .B(n2377), .Z(n2375) );
  OR U4367 ( .A(n2378), .B(n2379), .Z(n2374) );
  ANDN U4368 ( .B(n2380), .A(n2381), .Z(n2267) );
  IV U4369 ( .A(n2382), .Z(n2380) );
  XNOR U4370 ( .A(n2347), .B(n2346), .Z(N13617) );
  XOR U4371 ( .A(n2366), .B(n2365), .Z(n2346) );
  XNOR U4372 ( .A(n2381), .B(n2382), .Z(n2365) );
  XNOR U4373 ( .A(n2376), .B(n2377), .Z(n2382) );
  XNOR U4374 ( .A(n2378), .B(n2379), .Z(n2377) );
  XNOR U4375 ( .A(y[1837]), .B(x[1837]), .Z(n2379) );
  XNOR U4376 ( .A(y[1838]), .B(x[1838]), .Z(n2378) );
  XNOR U4377 ( .A(y[1836]), .B(x[1836]), .Z(n2376) );
  XNOR U4378 ( .A(n2370), .B(n2371), .Z(n2381) );
  XNOR U4379 ( .A(y[1833]), .B(x[1833]), .Z(n2371) );
  XNOR U4380 ( .A(n2372), .B(n2373), .Z(n2370) );
  XNOR U4381 ( .A(y[1834]), .B(x[1834]), .Z(n2373) );
  XNOR U4382 ( .A(y[1835]), .B(x[1835]), .Z(n2372) );
  XNOR U4383 ( .A(n2363), .B(n2362), .Z(n2366) );
  XNOR U4384 ( .A(n2358), .B(n2359), .Z(n2362) );
  XNOR U4385 ( .A(y[1830]), .B(x[1830]), .Z(n2359) );
  XNOR U4386 ( .A(n2360), .B(n2361), .Z(n2358) );
  XNOR U4387 ( .A(y[1831]), .B(x[1831]), .Z(n2361) );
  XNOR U4388 ( .A(y[1832]), .B(x[1832]), .Z(n2360) );
  XNOR U4389 ( .A(n2352), .B(n2353), .Z(n2363) );
  XNOR U4390 ( .A(y[1827]), .B(x[1827]), .Z(n2353) );
  XNOR U4391 ( .A(n2354), .B(n2355), .Z(n2352) );
  XNOR U4392 ( .A(y[1828]), .B(x[1828]), .Z(n2355) );
  XNOR U4393 ( .A(y[1829]), .B(x[1829]), .Z(n2354) );
  XOR U4394 ( .A(n2328), .B(n2329), .Z(n2347) );
  XNOR U4395 ( .A(n2344), .B(n2345), .Z(n2329) );
  XNOR U4396 ( .A(n2339), .B(n2340), .Z(n2345) );
  XNOR U4397 ( .A(n2341), .B(n2342), .Z(n2340) );
  XNOR U4398 ( .A(y[1825]), .B(x[1825]), .Z(n2342) );
  XNOR U4399 ( .A(y[1826]), .B(x[1826]), .Z(n2341) );
  XNOR U4400 ( .A(y[1824]), .B(x[1824]), .Z(n2339) );
  XNOR U4401 ( .A(n2333), .B(n2334), .Z(n2344) );
  XNOR U4402 ( .A(y[1821]), .B(x[1821]), .Z(n2334) );
  XNOR U4403 ( .A(n2335), .B(n2336), .Z(n2333) );
  XNOR U4404 ( .A(y[1822]), .B(x[1822]), .Z(n2336) );
  XNOR U4405 ( .A(y[1823]), .B(x[1823]), .Z(n2335) );
  XOR U4406 ( .A(n2327), .B(n2326), .Z(n2328) );
  XNOR U4407 ( .A(n2322), .B(n2323), .Z(n2326) );
  XNOR U4408 ( .A(y[1818]), .B(x[1818]), .Z(n2323) );
  XNOR U4409 ( .A(n2324), .B(n2325), .Z(n2322) );
  XNOR U4410 ( .A(y[1819]), .B(x[1819]), .Z(n2325) );
  XNOR U4411 ( .A(y[1820]), .B(x[1820]), .Z(n2324) );
  XNOR U4412 ( .A(n2316), .B(n2317), .Z(n2327) );
  XNOR U4413 ( .A(y[1815]), .B(x[1815]), .Z(n2317) );
  XNOR U4414 ( .A(n2318), .B(n2319), .Z(n2316) );
  XNOR U4415 ( .A(y[1816]), .B(x[1816]), .Z(n2319) );
  XNOR U4416 ( .A(y[1817]), .B(x[1817]), .Z(n2318) );
  NAND U4417 ( .A(n2383), .B(n2384), .Z(N13610) );
  NANDN U4418 ( .A(n2385), .B(n2386), .Z(n2384) );
  OR U4419 ( .A(n2387), .B(n2388), .Z(n2386) );
  NAND U4420 ( .A(n2387), .B(n2388), .Z(n2383) );
  XOR U4421 ( .A(n2387), .B(n2389), .Z(N13609) );
  XNOR U4422 ( .A(n2385), .B(n2388), .Z(n2389) );
  AND U4423 ( .A(n2390), .B(n2391), .Z(n2388) );
  NANDN U4424 ( .A(n2392), .B(n2393), .Z(n2391) );
  NANDN U4425 ( .A(n2394), .B(n2395), .Z(n2393) );
  NANDN U4426 ( .A(n2395), .B(n2394), .Z(n2390) );
  NAND U4427 ( .A(n2396), .B(n2397), .Z(n2385) );
  NANDN U4428 ( .A(n2398), .B(n2399), .Z(n2397) );
  OR U4429 ( .A(n2400), .B(n2401), .Z(n2399) );
  NAND U4430 ( .A(n2401), .B(n2400), .Z(n2396) );
  AND U4431 ( .A(n2402), .B(n2403), .Z(n2387) );
  NANDN U4432 ( .A(n2404), .B(n2405), .Z(n2403) );
  NANDN U4433 ( .A(n2406), .B(n2407), .Z(n2405) );
  NANDN U4434 ( .A(n2407), .B(n2406), .Z(n2402) );
  XOR U4435 ( .A(n2401), .B(n2408), .Z(N13608) );
  XOR U4436 ( .A(n2398), .B(n2400), .Z(n2408) );
  XNOR U4437 ( .A(n2394), .B(n2409), .Z(n2400) );
  XNOR U4438 ( .A(n2392), .B(n2395), .Z(n2409) );
  NAND U4439 ( .A(n2410), .B(n2411), .Z(n2395) );
  NAND U4440 ( .A(n2412), .B(n2413), .Z(n2411) );
  OR U4441 ( .A(n2414), .B(n2415), .Z(n2412) );
  NANDN U4442 ( .A(n2416), .B(n2414), .Z(n2410) );
  IV U4443 ( .A(n2415), .Z(n2416) );
  NAND U4444 ( .A(n2417), .B(n2418), .Z(n2392) );
  NAND U4445 ( .A(n2419), .B(n2420), .Z(n2418) );
  NANDN U4446 ( .A(n2421), .B(n2422), .Z(n2419) );
  NANDN U4447 ( .A(n2422), .B(n2421), .Z(n2417) );
  AND U4448 ( .A(n2423), .B(n2424), .Z(n2394) );
  NAND U4449 ( .A(n2425), .B(n2426), .Z(n2424) );
  OR U4450 ( .A(n2427), .B(n2428), .Z(n2425) );
  NANDN U4451 ( .A(n2429), .B(n2427), .Z(n2423) );
  NAND U4452 ( .A(n2430), .B(n2431), .Z(n2398) );
  NANDN U4453 ( .A(n2432), .B(n2433), .Z(n2431) );
  OR U4454 ( .A(n2434), .B(n2435), .Z(n2433) );
  NANDN U4455 ( .A(n2436), .B(n2434), .Z(n2430) );
  IV U4456 ( .A(n2435), .Z(n2436) );
  XNOR U4457 ( .A(n2406), .B(n2437), .Z(n2401) );
  XNOR U4458 ( .A(n2404), .B(n2407), .Z(n2437) );
  NAND U4459 ( .A(n2438), .B(n2439), .Z(n2407) );
  NAND U4460 ( .A(n2440), .B(n2441), .Z(n2439) );
  OR U4461 ( .A(n2442), .B(n2443), .Z(n2440) );
  NANDN U4462 ( .A(n2444), .B(n2442), .Z(n2438) );
  IV U4463 ( .A(n2443), .Z(n2444) );
  NAND U4464 ( .A(n2445), .B(n2446), .Z(n2404) );
  NAND U4465 ( .A(n2447), .B(n2448), .Z(n2446) );
  NANDN U4466 ( .A(n2449), .B(n2450), .Z(n2447) );
  NANDN U4467 ( .A(n2450), .B(n2449), .Z(n2445) );
  AND U4468 ( .A(n2451), .B(n2452), .Z(n2406) );
  NAND U4469 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U4470 ( .A(n2455), .B(n2456), .Z(n2453) );
  NANDN U4471 ( .A(n2457), .B(n2455), .Z(n2451) );
  XNOR U4472 ( .A(n2432), .B(n2458), .Z(N13607) );
  XOR U4473 ( .A(n2434), .B(n2435), .Z(n2458) );
  XNOR U4474 ( .A(n2448), .B(n2459), .Z(n2435) );
  XOR U4475 ( .A(n2449), .B(n2450), .Z(n2459) );
  XOR U4476 ( .A(n2455), .B(n2460), .Z(n2450) );
  XOR U4477 ( .A(n2454), .B(n2457), .Z(n2460) );
  IV U4478 ( .A(n2456), .Z(n2457) );
  NAND U4479 ( .A(n2461), .B(n2462), .Z(n2456) );
  OR U4480 ( .A(n2463), .B(n2464), .Z(n2462) );
  OR U4481 ( .A(n2465), .B(n2466), .Z(n2461) );
  NAND U4482 ( .A(n2467), .B(n2468), .Z(n2454) );
  OR U4483 ( .A(n2469), .B(n2470), .Z(n2468) );
  OR U4484 ( .A(n2471), .B(n2472), .Z(n2467) );
  NOR U4485 ( .A(n2473), .B(n2474), .Z(n2455) );
  ANDN U4486 ( .B(n2475), .A(n2476), .Z(n2449) );
  XNOR U4487 ( .A(n2442), .B(n2477), .Z(n2448) );
  XNOR U4488 ( .A(n2441), .B(n2443), .Z(n2477) );
  NAND U4489 ( .A(n2478), .B(n2479), .Z(n2443) );
  OR U4490 ( .A(n2480), .B(n2481), .Z(n2479) );
  OR U4491 ( .A(n2482), .B(n2483), .Z(n2478) );
  NAND U4492 ( .A(n2484), .B(n2485), .Z(n2441) );
  OR U4493 ( .A(n2486), .B(n2487), .Z(n2485) );
  OR U4494 ( .A(n2488), .B(n2489), .Z(n2484) );
  ANDN U4495 ( .B(n2490), .A(n2491), .Z(n2442) );
  IV U4496 ( .A(n2492), .Z(n2490) );
  ANDN U4497 ( .B(n2493), .A(n2494), .Z(n2434) );
  XOR U4498 ( .A(n2420), .B(n2495), .Z(n2432) );
  XOR U4499 ( .A(n2421), .B(n2422), .Z(n2495) );
  XOR U4500 ( .A(n2427), .B(n2496), .Z(n2422) );
  XOR U4501 ( .A(n2426), .B(n2429), .Z(n2496) );
  IV U4502 ( .A(n2428), .Z(n2429) );
  NAND U4503 ( .A(n2497), .B(n2498), .Z(n2428) );
  OR U4504 ( .A(n2499), .B(n2500), .Z(n2498) );
  OR U4505 ( .A(n2501), .B(n2502), .Z(n2497) );
  NAND U4506 ( .A(n2503), .B(n2504), .Z(n2426) );
  OR U4507 ( .A(n2505), .B(n2506), .Z(n2504) );
  OR U4508 ( .A(n2507), .B(n2508), .Z(n2503) );
  NOR U4509 ( .A(n2509), .B(n2510), .Z(n2427) );
  ANDN U4510 ( .B(n2511), .A(n2512), .Z(n2421) );
  IV U4511 ( .A(n2513), .Z(n2511) );
  XNOR U4512 ( .A(n2414), .B(n2514), .Z(n2420) );
  XNOR U4513 ( .A(n2413), .B(n2415), .Z(n2514) );
  NAND U4514 ( .A(n2515), .B(n2516), .Z(n2415) );
  OR U4515 ( .A(n2517), .B(n2518), .Z(n2516) );
  OR U4516 ( .A(n2519), .B(n2520), .Z(n2515) );
  NAND U4517 ( .A(n2521), .B(n2522), .Z(n2413) );
  OR U4518 ( .A(n2523), .B(n2524), .Z(n2522) );
  OR U4519 ( .A(n2525), .B(n2526), .Z(n2521) );
  ANDN U4520 ( .B(n2527), .A(n2528), .Z(n2414) );
  IV U4521 ( .A(n2529), .Z(n2527) );
  XNOR U4522 ( .A(n2494), .B(n2493), .Z(N13606) );
  XOR U4523 ( .A(n2513), .B(n2512), .Z(n2493) );
  XNOR U4524 ( .A(n2528), .B(n2529), .Z(n2512) );
  XNOR U4525 ( .A(n2523), .B(n2524), .Z(n2529) );
  XNOR U4526 ( .A(n2525), .B(n2526), .Z(n2524) );
  XNOR U4527 ( .A(y[1813]), .B(x[1813]), .Z(n2526) );
  XNOR U4528 ( .A(y[1814]), .B(x[1814]), .Z(n2525) );
  XNOR U4529 ( .A(y[1812]), .B(x[1812]), .Z(n2523) );
  XNOR U4530 ( .A(n2517), .B(n2518), .Z(n2528) );
  XNOR U4531 ( .A(y[1809]), .B(x[1809]), .Z(n2518) );
  XNOR U4532 ( .A(n2519), .B(n2520), .Z(n2517) );
  XNOR U4533 ( .A(y[1810]), .B(x[1810]), .Z(n2520) );
  XNOR U4534 ( .A(y[1811]), .B(x[1811]), .Z(n2519) );
  XNOR U4535 ( .A(n2510), .B(n2509), .Z(n2513) );
  XNOR U4536 ( .A(n2505), .B(n2506), .Z(n2509) );
  XNOR U4537 ( .A(y[1806]), .B(x[1806]), .Z(n2506) );
  XNOR U4538 ( .A(n2507), .B(n2508), .Z(n2505) );
  XNOR U4539 ( .A(y[1807]), .B(x[1807]), .Z(n2508) );
  XNOR U4540 ( .A(y[1808]), .B(x[1808]), .Z(n2507) );
  XNOR U4541 ( .A(n2499), .B(n2500), .Z(n2510) );
  XNOR U4542 ( .A(y[1803]), .B(x[1803]), .Z(n2500) );
  XNOR U4543 ( .A(n2501), .B(n2502), .Z(n2499) );
  XNOR U4544 ( .A(y[1804]), .B(x[1804]), .Z(n2502) );
  XNOR U4545 ( .A(y[1805]), .B(x[1805]), .Z(n2501) );
  XOR U4546 ( .A(n2475), .B(n2476), .Z(n2494) );
  XNOR U4547 ( .A(n2491), .B(n2492), .Z(n2476) );
  XNOR U4548 ( .A(n2486), .B(n2487), .Z(n2492) );
  XNOR U4549 ( .A(n2488), .B(n2489), .Z(n2487) );
  XNOR U4550 ( .A(y[1801]), .B(x[1801]), .Z(n2489) );
  XNOR U4551 ( .A(y[1802]), .B(x[1802]), .Z(n2488) );
  XNOR U4552 ( .A(y[1800]), .B(x[1800]), .Z(n2486) );
  XNOR U4553 ( .A(n2480), .B(n2481), .Z(n2491) );
  XNOR U4554 ( .A(y[1797]), .B(x[1797]), .Z(n2481) );
  XNOR U4555 ( .A(n2482), .B(n2483), .Z(n2480) );
  XNOR U4556 ( .A(y[1798]), .B(x[1798]), .Z(n2483) );
  XNOR U4557 ( .A(y[1799]), .B(x[1799]), .Z(n2482) );
  XOR U4558 ( .A(n2474), .B(n2473), .Z(n2475) );
  XNOR U4559 ( .A(n2469), .B(n2470), .Z(n2473) );
  XNOR U4560 ( .A(y[1794]), .B(x[1794]), .Z(n2470) );
  XNOR U4561 ( .A(n2471), .B(n2472), .Z(n2469) );
  XNOR U4562 ( .A(y[1795]), .B(x[1795]), .Z(n2472) );
  XNOR U4563 ( .A(y[1796]), .B(x[1796]), .Z(n2471) );
  XNOR U4564 ( .A(n2463), .B(n2464), .Z(n2474) );
  XNOR U4565 ( .A(y[1791]), .B(x[1791]), .Z(n2464) );
  XNOR U4566 ( .A(n2465), .B(n2466), .Z(n2463) );
  XNOR U4567 ( .A(y[1792]), .B(x[1792]), .Z(n2466) );
  XNOR U4568 ( .A(y[1793]), .B(x[1793]), .Z(n2465) );
  NAND U4569 ( .A(n2530), .B(n2531), .Z(N13599) );
  NANDN U4570 ( .A(n2532), .B(n2533), .Z(n2531) );
  OR U4571 ( .A(n2534), .B(n2535), .Z(n2533) );
  NAND U4572 ( .A(n2534), .B(n2535), .Z(n2530) );
  XOR U4573 ( .A(n2534), .B(n2536), .Z(N13598) );
  XNOR U4574 ( .A(n2532), .B(n2535), .Z(n2536) );
  AND U4575 ( .A(n2537), .B(n2538), .Z(n2535) );
  NANDN U4576 ( .A(n2539), .B(n2540), .Z(n2538) );
  NANDN U4577 ( .A(n2541), .B(n2542), .Z(n2540) );
  NANDN U4578 ( .A(n2542), .B(n2541), .Z(n2537) );
  NAND U4579 ( .A(n2543), .B(n2544), .Z(n2532) );
  NANDN U4580 ( .A(n2545), .B(n2546), .Z(n2544) );
  OR U4581 ( .A(n2547), .B(n2548), .Z(n2546) );
  NAND U4582 ( .A(n2548), .B(n2547), .Z(n2543) );
  AND U4583 ( .A(n2549), .B(n2550), .Z(n2534) );
  NANDN U4584 ( .A(n2551), .B(n2552), .Z(n2550) );
  NANDN U4585 ( .A(n2553), .B(n2554), .Z(n2552) );
  NANDN U4586 ( .A(n2554), .B(n2553), .Z(n2549) );
  XOR U4587 ( .A(n2548), .B(n2555), .Z(N13597) );
  XOR U4588 ( .A(n2545), .B(n2547), .Z(n2555) );
  XNOR U4589 ( .A(n2541), .B(n2556), .Z(n2547) );
  XNOR U4590 ( .A(n2539), .B(n2542), .Z(n2556) );
  NAND U4591 ( .A(n2557), .B(n2558), .Z(n2542) );
  NAND U4592 ( .A(n2559), .B(n2560), .Z(n2558) );
  OR U4593 ( .A(n2561), .B(n2562), .Z(n2559) );
  NANDN U4594 ( .A(n2563), .B(n2561), .Z(n2557) );
  IV U4595 ( .A(n2562), .Z(n2563) );
  NAND U4596 ( .A(n2564), .B(n2565), .Z(n2539) );
  NAND U4597 ( .A(n2566), .B(n2567), .Z(n2565) );
  NANDN U4598 ( .A(n2568), .B(n2569), .Z(n2566) );
  NANDN U4599 ( .A(n2569), .B(n2568), .Z(n2564) );
  AND U4600 ( .A(n2570), .B(n2571), .Z(n2541) );
  NAND U4601 ( .A(n2572), .B(n2573), .Z(n2571) );
  OR U4602 ( .A(n2574), .B(n2575), .Z(n2572) );
  NANDN U4603 ( .A(n2576), .B(n2574), .Z(n2570) );
  NAND U4604 ( .A(n2577), .B(n2578), .Z(n2545) );
  NANDN U4605 ( .A(n2579), .B(n2580), .Z(n2578) );
  OR U4606 ( .A(n2581), .B(n2582), .Z(n2580) );
  NANDN U4607 ( .A(n2583), .B(n2581), .Z(n2577) );
  IV U4608 ( .A(n2582), .Z(n2583) );
  XNOR U4609 ( .A(n2553), .B(n2584), .Z(n2548) );
  XNOR U4610 ( .A(n2551), .B(n2554), .Z(n2584) );
  NAND U4611 ( .A(n2585), .B(n2586), .Z(n2554) );
  NAND U4612 ( .A(n2587), .B(n2588), .Z(n2586) );
  OR U4613 ( .A(n2589), .B(n2590), .Z(n2587) );
  NANDN U4614 ( .A(n2591), .B(n2589), .Z(n2585) );
  IV U4615 ( .A(n2590), .Z(n2591) );
  NAND U4616 ( .A(n2592), .B(n2593), .Z(n2551) );
  NAND U4617 ( .A(n2594), .B(n2595), .Z(n2593) );
  NANDN U4618 ( .A(n2596), .B(n2597), .Z(n2594) );
  NANDN U4619 ( .A(n2597), .B(n2596), .Z(n2592) );
  AND U4620 ( .A(n2598), .B(n2599), .Z(n2553) );
  NAND U4621 ( .A(n2600), .B(n2601), .Z(n2599) );
  OR U4622 ( .A(n2602), .B(n2603), .Z(n2600) );
  NANDN U4623 ( .A(n2604), .B(n2602), .Z(n2598) );
  XNOR U4624 ( .A(n2579), .B(n2605), .Z(N13596) );
  XOR U4625 ( .A(n2581), .B(n2582), .Z(n2605) );
  XNOR U4626 ( .A(n2595), .B(n2606), .Z(n2582) );
  XOR U4627 ( .A(n2596), .B(n2597), .Z(n2606) );
  XOR U4628 ( .A(n2602), .B(n2607), .Z(n2597) );
  XOR U4629 ( .A(n2601), .B(n2604), .Z(n2607) );
  IV U4630 ( .A(n2603), .Z(n2604) );
  NAND U4631 ( .A(n2608), .B(n2609), .Z(n2603) );
  OR U4632 ( .A(n2610), .B(n2611), .Z(n2609) );
  OR U4633 ( .A(n2612), .B(n2613), .Z(n2608) );
  NAND U4634 ( .A(n2614), .B(n2615), .Z(n2601) );
  OR U4635 ( .A(n2616), .B(n2617), .Z(n2615) );
  OR U4636 ( .A(n2618), .B(n2619), .Z(n2614) );
  NOR U4637 ( .A(n2620), .B(n2621), .Z(n2602) );
  ANDN U4638 ( .B(n2622), .A(n2623), .Z(n2596) );
  XNOR U4639 ( .A(n2589), .B(n2624), .Z(n2595) );
  XNOR U4640 ( .A(n2588), .B(n2590), .Z(n2624) );
  NAND U4641 ( .A(n2625), .B(n2626), .Z(n2590) );
  OR U4642 ( .A(n2627), .B(n2628), .Z(n2626) );
  OR U4643 ( .A(n2629), .B(n2630), .Z(n2625) );
  NAND U4644 ( .A(n2631), .B(n2632), .Z(n2588) );
  OR U4645 ( .A(n2633), .B(n2634), .Z(n2632) );
  OR U4646 ( .A(n2635), .B(n2636), .Z(n2631) );
  ANDN U4647 ( .B(n2637), .A(n2638), .Z(n2589) );
  IV U4648 ( .A(n2639), .Z(n2637) );
  ANDN U4649 ( .B(n2640), .A(n2641), .Z(n2581) );
  XOR U4650 ( .A(n2567), .B(n2642), .Z(n2579) );
  XOR U4651 ( .A(n2568), .B(n2569), .Z(n2642) );
  XOR U4652 ( .A(n2574), .B(n2643), .Z(n2569) );
  XOR U4653 ( .A(n2573), .B(n2576), .Z(n2643) );
  IV U4654 ( .A(n2575), .Z(n2576) );
  NAND U4655 ( .A(n2644), .B(n2645), .Z(n2575) );
  OR U4656 ( .A(n2646), .B(n2647), .Z(n2645) );
  OR U4657 ( .A(n2648), .B(n2649), .Z(n2644) );
  NAND U4658 ( .A(n2650), .B(n2651), .Z(n2573) );
  OR U4659 ( .A(n2652), .B(n2653), .Z(n2651) );
  OR U4660 ( .A(n2654), .B(n2655), .Z(n2650) );
  NOR U4661 ( .A(n2656), .B(n2657), .Z(n2574) );
  ANDN U4662 ( .B(n2658), .A(n2659), .Z(n2568) );
  IV U4663 ( .A(n2660), .Z(n2658) );
  XNOR U4664 ( .A(n2561), .B(n2661), .Z(n2567) );
  XNOR U4665 ( .A(n2560), .B(n2562), .Z(n2661) );
  NAND U4666 ( .A(n2662), .B(n2663), .Z(n2562) );
  OR U4667 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U4668 ( .A(n2666), .B(n2667), .Z(n2662) );
  NAND U4669 ( .A(n2668), .B(n2669), .Z(n2560) );
  OR U4670 ( .A(n2670), .B(n2671), .Z(n2669) );
  OR U4671 ( .A(n2672), .B(n2673), .Z(n2668) );
  ANDN U4672 ( .B(n2674), .A(n2675), .Z(n2561) );
  IV U4673 ( .A(n2676), .Z(n2674) );
  XNOR U4674 ( .A(n2641), .B(n2640), .Z(N13595) );
  XOR U4675 ( .A(n2660), .B(n2659), .Z(n2640) );
  XNOR U4676 ( .A(n2675), .B(n2676), .Z(n2659) );
  XNOR U4677 ( .A(n2670), .B(n2671), .Z(n2676) );
  XNOR U4678 ( .A(n2672), .B(n2673), .Z(n2671) );
  XNOR U4679 ( .A(y[1789]), .B(x[1789]), .Z(n2673) );
  XNOR U4680 ( .A(y[1790]), .B(x[1790]), .Z(n2672) );
  XNOR U4681 ( .A(y[1788]), .B(x[1788]), .Z(n2670) );
  XNOR U4682 ( .A(n2664), .B(n2665), .Z(n2675) );
  XNOR U4683 ( .A(y[1785]), .B(x[1785]), .Z(n2665) );
  XNOR U4684 ( .A(n2666), .B(n2667), .Z(n2664) );
  XNOR U4685 ( .A(y[1786]), .B(x[1786]), .Z(n2667) );
  XNOR U4686 ( .A(y[1787]), .B(x[1787]), .Z(n2666) );
  XNOR U4687 ( .A(n2657), .B(n2656), .Z(n2660) );
  XNOR U4688 ( .A(n2652), .B(n2653), .Z(n2656) );
  XNOR U4689 ( .A(y[1782]), .B(x[1782]), .Z(n2653) );
  XNOR U4690 ( .A(n2654), .B(n2655), .Z(n2652) );
  XNOR U4691 ( .A(y[1783]), .B(x[1783]), .Z(n2655) );
  XNOR U4692 ( .A(y[1784]), .B(x[1784]), .Z(n2654) );
  XNOR U4693 ( .A(n2646), .B(n2647), .Z(n2657) );
  XNOR U4694 ( .A(y[1779]), .B(x[1779]), .Z(n2647) );
  XNOR U4695 ( .A(n2648), .B(n2649), .Z(n2646) );
  XNOR U4696 ( .A(y[1780]), .B(x[1780]), .Z(n2649) );
  XNOR U4697 ( .A(y[1781]), .B(x[1781]), .Z(n2648) );
  XOR U4698 ( .A(n2622), .B(n2623), .Z(n2641) );
  XNOR U4699 ( .A(n2638), .B(n2639), .Z(n2623) );
  XNOR U4700 ( .A(n2633), .B(n2634), .Z(n2639) );
  XNOR U4701 ( .A(n2635), .B(n2636), .Z(n2634) );
  XNOR U4702 ( .A(y[1777]), .B(x[1777]), .Z(n2636) );
  XNOR U4703 ( .A(y[1778]), .B(x[1778]), .Z(n2635) );
  XNOR U4704 ( .A(y[1776]), .B(x[1776]), .Z(n2633) );
  XNOR U4705 ( .A(n2627), .B(n2628), .Z(n2638) );
  XNOR U4706 ( .A(y[1773]), .B(x[1773]), .Z(n2628) );
  XNOR U4707 ( .A(n2629), .B(n2630), .Z(n2627) );
  XNOR U4708 ( .A(y[1774]), .B(x[1774]), .Z(n2630) );
  XNOR U4709 ( .A(y[1775]), .B(x[1775]), .Z(n2629) );
  XOR U4710 ( .A(n2621), .B(n2620), .Z(n2622) );
  XNOR U4711 ( .A(n2616), .B(n2617), .Z(n2620) );
  XNOR U4712 ( .A(y[1770]), .B(x[1770]), .Z(n2617) );
  XNOR U4713 ( .A(n2618), .B(n2619), .Z(n2616) );
  XNOR U4714 ( .A(y[1771]), .B(x[1771]), .Z(n2619) );
  XNOR U4715 ( .A(y[1772]), .B(x[1772]), .Z(n2618) );
  XNOR U4716 ( .A(n2610), .B(n2611), .Z(n2621) );
  XNOR U4717 ( .A(y[1767]), .B(x[1767]), .Z(n2611) );
  XNOR U4718 ( .A(n2612), .B(n2613), .Z(n2610) );
  XNOR U4719 ( .A(y[1768]), .B(x[1768]), .Z(n2613) );
  XNOR U4720 ( .A(y[1769]), .B(x[1769]), .Z(n2612) );
  NAND U4721 ( .A(n2677), .B(n2678), .Z(N13588) );
  NANDN U4722 ( .A(n2679), .B(n2680), .Z(n2678) );
  OR U4723 ( .A(n2681), .B(n2682), .Z(n2680) );
  NAND U4724 ( .A(n2681), .B(n2682), .Z(n2677) );
  XOR U4725 ( .A(n2681), .B(n2683), .Z(N13587) );
  XNOR U4726 ( .A(n2679), .B(n2682), .Z(n2683) );
  AND U4727 ( .A(n2684), .B(n2685), .Z(n2682) );
  NANDN U4728 ( .A(n2686), .B(n2687), .Z(n2685) );
  NANDN U4729 ( .A(n2688), .B(n2689), .Z(n2687) );
  NANDN U4730 ( .A(n2689), .B(n2688), .Z(n2684) );
  NAND U4731 ( .A(n2690), .B(n2691), .Z(n2679) );
  NANDN U4732 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U4733 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U4734 ( .A(n2695), .B(n2694), .Z(n2690) );
  AND U4735 ( .A(n2696), .B(n2697), .Z(n2681) );
  NANDN U4736 ( .A(n2698), .B(n2699), .Z(n2697) );
  NANDN U4737 ( .A(n2700), .B(n2701), .Z(n2699) );
  NANDN U4738 ( .A(n2701), .B(n2700), .Z(n2696) );
  XOR U4739 ( .A(n2695), .B(n2702), .Z(N13586) );
  XOR U4740 ( .A(n2692), .B(n2694), .Z(n2702) );
  XNOR U4741 ( .A(n2688), .B(n2703), .Z(n2694) );
  XNOR U4742 ( .A(n2686), .B(n2689), .Z(n2703) );
  NAND U4743 ( .A(n2704), .B(n2705), .Z(n2689) );
  NAND U4744 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U4745 ( .A(n2708), .B(n2709), .Z(n2706) );
  NANDN U4746 ( .A(n2710), .B(n2708), .Z(n2704) );
  IV U4747 ( .A(n2709), .Z(n2710) );
  NAND U4748 ( .A(n2711), .B(n2712), .Z(n2686) );
  NAND U4749 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U4750 ( .A(n2715), .B(n2716), .Z(n2713) );
  NANDN U4751 ( .A(n2716), .B(n2715), .Z(n2711) );
  AND U4752 ( .A(n2717), .B(n2718), .Z(n2688) );
  NAND U4753 ( .A(n2719), .B(n2720), .Z(n2718) );
  OR U4754 ( .A(n2721), .B(n2722), .Z(n2719) );
  NANDN U4755 ( .A(n2723), .B(n2721), .Z(n2717) );
  NAND U4756 ( .A(n2724), .B(n2725), .Z(n2692) );
  NANDN U4757 ( .A(n2726), .B(n2727), .Z(n2725) );
  OR U4758 ( .A(n2728), .B(n2729), .Z(n2727) );
  NANDN U4759 ( .A(n2730), .B(n2728), .Z(n2724) );
  IV U4760 ( .A(n2729), .Z(n2730) );
  XNOR U4761 ( .A(n2700), .B(n2731), .Z(n2695) );
  XNOR U4762 ( .A(n2698), .B(n2701), .Z(n2731) );
  NAND U4763 ( .A(n2732), .B(n2733), .Z(n2701) );
  NAND U4764 ( .A(n2734), .B(n2735), .Z(n2733) );
  OR U4765 ( .A(n2736), .B(n2737), .Z(n2734) );
  NANDN U4766 ( .A(n2738), .B(n2736), .Z(n2732) );
  IV U4767 ( .A(n2737), .Z(n2738) );
  NAND U4768 ( .A(n2739), .B(n2740), .Z(n2698) );
  NAND U4769 ( .A(n2741), .B(n2742), .Z(n2740) );
  NANDN U4770 ( .A(n2743), .B(n2744), .Z(n2741) );
  NANDN U4771 ( .A(n2744), .B(n2743), .Z(n2739) );
  AND U4772 ( .A(n2745), .B(n2746), .Z(n2700) );
  NAND U4773 ( .A(n2747), .B(n2748), .Z(n2746) );
  OR U4774 ( .A(n2749), .B(n2750), .Z(n2747) );
  NANDN U4775 ( .A(n2751), .B(n2749), .Z(n2745) );
  XNOR U4776 ( .A(n2726), .B(n2752), .Z(N13585) );
  XOR U4777 ( .A(n2728), .B(n2729), .Z(n2752) );
  XNOR U4778 ( .A(n2742), .B(n2753), .Z(n2729) );
  XOR U4779 ( .A(n2743), .B(n2744), .Z(n2753) );
  XOR U4780 ( .A(n2749), .B(n2754), .Z(n2744) );
  XOR U4781 ( .A(n2748), .B(n2751), .Z(n2754) );
  IV U4782 ( .A(n2750), .Z(n2751) );
  NAND U4783 ( .A(n2755), .B(n2756), .Z(n2750) );
  OR U4784 ( .A(n2757), .B(n2758), .Z(n2756) );
  OR U4785 ( .A(n2759), .B(n2760), .Z(n2755) );
  NAND U4786 ( .A(n2761), .B(n2762), .Z(n2748) );
  OR U4787 ( .A(n2763), .B(n2764), .Z(n2762) );
  OR U4788 ( .A(n2765), .B(n2766), .Z(n2761) );
  NOR U4789 ( .A(n2767), .B(n2768), .Z(n2749) );
  ANDN U4790 ( .B(n2769), .A(n2770), .Z(n2743) );
  XNOR U4791 ( .A(n2736), .B(n2771), .Z(n2742) );
  XNOR U4792 ( .A(n2735), .B(n2737), .Z(n2771) );
  NAND U4793 ( .A(n2772), .B(n2773), .Z(n2737) );
  OR U4794 ( .A(n2774), .B(n2775), .Z(n2773) );
  OR U4795 ( .A(n2776), .B(n2777), .Z(n2772) );
  NAND U4796 ( .A(n2778), .B(n2779), .Z(n2735) );
  OR U4797 ( .A(n2780), .B(n2781), .Z(n2779) );
  OR U4798 ( .A(n2782), .B(n2783), .Z(n2778) );
  ANDN U4799 ( .B(n2784), .A(n2785), .Z(n2736) );
  IV U4800 ( .A(n2786), .Z(n2784) );
  ANDN U4801 ( .B(n2787), .A(n2788), .Z(n2728) );
  XOR U4802 ( .A(n2714), .B(n2789), .Z(n2726) );
  XOR U4803 ( .A(n2715), .B(n2716), .Z(n2789) );
  XOR U4804 ( .A(n2721), .B(n2790), .Z(n2716) );
  XOR U4805 ( .A(n2720), .B(n2723), .Z(n2790) );
  IV U4806 ( .A(n2722), .Z(n2723) );
  NAND U4807 ( .A(n2791), .B(n2792), .Z(n2722) );
  OR U4808 ( .A(n2793), .B(n2794), .Z(n2792) );
  OR U4809 ( .A(n2795), .B(n2796), .Z(n2791) );
  NAND U4810 ( .A(n2797), .B(n2798), .Z(n2720) );
  OR U4811 ( .A(n2799), .B(n2800), .Z(n2798) );
  OR U4812 ( .A(n2801), .B(n2802), .Z(n2797) );
  NOR U4813 ( .A(n2803), .B(n2804), .Z(n2721) );
  ANDN U4814 ( .B(n2805), .A(n2806), .Z(n2715) );
  IV U4815 ( .A(n2807), .Z(n2805) );
  XNOR U4816 ( .A(n2708), .B(n2808), .Z(n2714) );
  XNOR U4817 ( .A(n2707), .B(n2709), .Z(n2808) );
  NAND U4818 ( .A(n2809), .B(n2810), .Z(n2709) );
  OR U4819 ( .A(n2811), .B(n2812), .Z(n2810) );
  OR U4820 ( .A(n2813), .B(n2814), .Z(n2809) );
  NAND U4821 ( .A(n2815), .B(n2816), .Z(n2707) );
  OR U4822 ( .A(n2817), .B(n2818), .Z(n2816) );
  OR U4823 ( .A(n2819), .B(n2820), .Z(n2815) );
  ANDN U4824 ( .B(n2821), .A(n2822), .Z(n2708) );
  IV U4825 ( .A(n2823), .Z(n2821) );
  XNOR U4826 ( .A(n2788), .B(n2787), .Z(N13584) );
  XOR U4827 ( .A(n2807), .B(n2806), .Z(n2787) );
  XNOR U4828 ( .A(n2822), .B(n2823), .Z(n2806) );
  XNOR U4829 ( .A(n2817), .B(n2818), .Z(n2823) );
  XNOR U4830 ( .A(n2819), .B(n2820), .Z(n2818) );
  XNOR U4831 ( .A(y[1765]), .B(x[1765]), .Z(n2820) );
  XNOR U4832 ( .A(y[1766]), .B(x[1766]), .Z(n2819) );
  XNOR U4833 ( .A(y[1764]), .B(x[1764]), .Z(n2817) );
  XNOR U4834 ( .A(n2811), .B(n2812), .Z(n2822) );
  XNOR U4835 ( .A(y[1761]), .B(x[1761]), .Z(n2812) );
  XNOR U4836 ( .A(n2813), .B(n2814), .Z(n2811) );
  XNOR U4837 ( .A(y[1762]), .B(x[1762]), .Z(n2814) );
  XNOR U4838 ( .A(y[1763]), .B(x[1763]), .Z(n2813) );
  XNOR U4839 ( .A(n2804), .B(n2803), .Z(n2807) );
  XNOR U4840 ( .A(n2799), .B(n2800), .Z(n2803) );
  XNOR U4841 ( .A(y[1758]), .B(x[1758]), .Z(n2800) );
  XNOR U4842 ( .A(n2801), .B(n2802), .Z(n2799) );
  XNOR U4843 ( .A(y[1759]), .B(x[1759]), .Z(n2802) );
  XNOR U4844 ( .A(y[1760]), .B(x[1760]), .Z(n2801) );
  XNOR U4845 ( .A(n2793), .B(n2794), .Z(n2804) );
  XNOR U4846 ( .A(y[1755]), .B(x[1755]), .Z(n2794) );
  XNOR U4847 ( .A(n2795), .B(n2796), .Z(n2793) );
  XNOR U4848 ( .A(y[1756]), .B(x[1756]), .Z(n2796) );
  XNOR U4849 ( .A(y[1757]), .B(x[1757]), .Z(n2795) );
  XOR U4850 ( .A(n2769), .B(n2770), .Z(n2788) );
  XNOR U4851 ( .A(n2785), .B(n2786), .Z(n2770) );
  XNOR U4852 ( .A(n2780), .B(n2781), .Z(n2786) );
  XNOR U4853 ( .A(n2782), .B(n2783), .Z(n2781) );
  XNOR U4854 ( .A(y[1753]), .B(x[1753]), .Z(n2783) );
  XNOR U4855 ( .A(y[1754]), .B(x[1754]), .Z(n2782) );
  XNOR U4856 ( .A(y[1752]), .B(x[1752]), .Z(n2780) );
  XNOR U4857 ( .A(n2774), .B(n2775), .Z(n2785) );
  XNOR U4858 ( .A(y[1749]), .B(x[1749]), .Z(n2775) );
  XNOR U4859 ( .A(n2776), .B(n2777), .Z(n2774) );
  XNOR U4860 ( .A(y[1750]), .B(x[1750]), .Z(n2777) );
  XNOR U4861 ( .A(y[1751]), .B(x[1751]), .Z(n2776) );
  XOR U4862 ( .A(n2768), .B(n2767), .Z(n2769) );
  XNOR U4863 ( .A(n2763), .B(n2764), .Z(n2767) );
  XNOR U4864 ( .A(y[1746]), .B(x[1746]), .Z(n2764) );
  XNOR U4865 ( .A(n2765), .B(n2766), .Z(n2763) );
  XNOR U4866 ( .A(y[1747]), .B(x[1747]), .Z(n2766) );
  XNOR U4867 ( .A(y[1748]), .B(x[1748]), .Z(n2765) );
  XNOR U4868 ( .A(n2757), .B(n2758), .Z(n2768) );
  XNOR U4869 ( .A(y[1743]), .B(x[1743]), .Z(n2758) );
  XNOR U4870 ( .A(n2759), .B(n2760), .Z(n2757) );
  XNOR U4871 ( .A(y[1744]), .B(x[1744]), .Z(n2760) );
  XNOR U4872 ( .A(y[1745]), .B(x[1745]), .Z(n2759) );
  NAND U4873 ( .A(n2824), .B(n2825), .Z(N13577) );
  NANDN U4874 ( .A(n2826), .B(n2827), .Z(n2825) );
  OR U4875 ( .A(n2828), .B(n2829), .Z(n2827) );
  NAND U4876 ( .A(n2828), .B(n2829), .Z(n2824) );
  XOR U4877 ( .A(n2828), .B(n2830), .Z(N13576) );
  XNOR U4878 ( .A(n2826), .B(n2829), .Z(n2830) );
  AND U4879 ( .A(n2831), .B(n2832), .Z(n2829) );
  NANDN U4880 ( .A(n2833), .B(n2834), .Z(n2832) );
  NANDN U4881 ( .A(n2835), .B(n2836), .Z(n2834) );
  NANDN U4882 ( .A(n2836), .B(n2835), .Z(n2831) );
  NAND U4883 ( .A(n2837), .B(n2838), .Z(n2826) );
  NANDN U4884 ( .A(n2839), .B(n2840), .Z(n2838) );
  OR U4885 ( .A(n2841), .B(n2842), .Z(n2840) );
  NAND U4886 ( .A(n2842), .B(n2841), .Z(n2837) );
  AND U4887 ( .A(n2843), .B(n2844), .Z(n2828) );
  NANDN U4888 ( .A(n2845), .B(n2846), .Z(n2844) );
  NANDN U4889 ( .A(n2847), .B(n2848), .Z(n2846) );
  NANDN U4890 ( .A(n2848), .B(n2847), .Z(n2843) );
  XOR U4891 ( .A(n2842), .B(n2849), .Z(N13575) );
  XOR U4892 ( .A(n2839), .B(n2841), .Z(n2849) );
  XNOR U4893 ( .A(n2835), .B(n2850), .Z(n2841) );
  XNOR U4894 ( .A(n2833), .B(n2836), .Z(n2850) );
  NAND U4895 ( .A(n2851), .B(n2852), .Z(n2836) );
  NAND U4896 ( .A(n2853), .B(n2854), .Z(n2852) );
  OR U4897 ( .A(n2855), .B(n2856), .Z(n2853) );
  NANDN U4898 ( .A(n2857), .B(n2855), .Z(n2851) );
  IV U4899 ( .A(n2856), .Z(n2857) );
  NAND U4900 ( .A(n2858), .B(n2859), .Z(n2833) );
  NAND U4901 ( .A(n2860), .B(n2861), .Z(n2859) );
  NANDN U4902 ( .A(n2862), .B(n2863), .Z(n2860) );
  NANDN U4903 ( .A(n2863), .B(n2862), .Z(n2858) );
  AND U4904 ( .A(n2864), .B(n2865), .Z(n2835) );
  NAND U4905 ( .A(n2866), .B(n2867), .Z(n2865) );
  OR U4906 ( .A(n2868), .B(n2869), .Z(n2866) );
  NANDN U4907 ( .A(n2870), .B(n2868), .Z(n2864) );
  NAND U4908 ( .A(n2871), .B(n2872), .Z(n2839) );
  NANDN U4909 ( .A(n2873), .B(n2874), .Z(n2872) );
  OR U4910 ( .A(n2875), .B(n2876), .Z(n2874) );
  NANDN U4911 ( .A(n2877), .B(n2875), .Z(n2871) );
  IV U4912 ( .A(n2876), .Z(n2877) );
  XNOR U4913 ( .A(n2847), .B(n2878), .Z(n2842) );
  XNOR U4914 ( .A(n2845), .B(n2848), .Z(n2878) );
  NAND U4915 ( .A(n2879), .B(n2880), .Z(n2848) );
  NAND U4916 ( .A(n2881), .B(n2882), .Z(n2880) );
  OR U4917 ( .A(n2883), .B(n2884), .Z(n2881) );
  NANDN U4918 ( .A(n2885), .B(n2883), .Z(n2879) );
  IV U4919 ( .A(n2884), .Z(n2885) );
  NAND U4920 ( .A(n2886), .B(n2887), .Z(n2845) );
  NAND U4921 ( .A(n2888), .B(n2889), .Z(n2887) );
  NANDN U4922 ( .A(n2890), .B(n2891), .Z(n2888) );
  NANDN U4923 ( .A(n2891), .B(n2890), .Z(n2886) );
  AND U4924 ( .A(n2892), .B(n2893), .Z(n2847) );
  NAND U4925 ( .A(n2894), .B(n2895), .Z(n2893) );
  OR U4926 ( .A(n2896), .B(n2897), .Z(n2894) );
  NANDN U4927 ( .A(n2898), .B(n2896), .Z(n2892) );
  XNOR U4928 ( .A(n2873), .B(n2899), .Z(N13574) );
  XOR U4929 ( .A(n2875), .B(n2876), .Z(n2899) );
  XNOR U4930 ( .A(n2889), .B(n2900), .Z(n2876) );
  XOR U4931 ( .A(n2890), .B(n2891), .Z(n2900) );
  XOR U4932 ( .A(n2896), .B(n2901), .Z(n2891) );
  XOR U4933 ( .A(n2895), .B(n2898), .Z(n2901) );
  IV U4934 ( .A(n2897), .Z(n2898) );
  NAND U4935 ( .A(n2902), .B(n2903), .Z(n2897) );
  OR U4936 ( .A(n2904), .B(n2905), .Z(n2903) );
  OR U4937 ( .A(n2906), .B(n2907), .Z(n2902) );
  NAND U4938 ( .A(n2908), .B(n2909), .Z(n2895) );
  OR U4939 ( .A(n2910), .B(n2911), .Z(n2909) );
  OR U4940 ( .A(n2912), .B(n2913), .Z(n2908) );
  NOR U4941 ( .A(n2914), .B(n2915), .Z(n2896) );
  ANDN U4942 ( .B(n2916), .A(n2917), .Z(n2890) );
  XNOR U4943 ( .A(n2883), .B(n2918), .Z(n2889) );
  XNOR U4944 ( .A(n2882), .B(n2884), .Z(n2918) );
  NAND U4945 ( .A(n2919), .B(n2920), .Z(n2884) );
  OR U4946 ( .A(n2921), .B(n2922), .Z(n2920) );
  OR U4947 ( .A(n2923), .B(n2924), .Z(n2919) );
  NAND U4948 ( .A(n2925), .B(n2926), .Z(n2882) );
  OR U4949 ( .A(n2927), .B(n2928), .Z(n2926) );
  OR U4950 ( .A(n2929), .B(n2930), .Z(n2925) );
  ANDN U4951 ( .B(n2931), .A(n2932), .Z(n2883) );
  IV U4952 ( .A(n2933), .Z(n2931) );
  ANDN U4953 ( .B(n2934), .A(n2935), .Z(n2875) );
  XOR U4954 ( .A(n2861), .B(n2936), .Z(n2873) );
  XOR U4955 ( .A(n2862), .B(n2863), .Z(n2936) );
  XOR U4956 ( .A(n2868), .B(n2937), .Z(n2863) );
  XOR U4957 ( .A(n2867), .B(n2870), .Z(n2937) );
  IV U4958 ( .A(n2869), .Z(n2870) );
  NAND U4959 ( .A(n2938), .B(n2939), .Z(n2869) );
  OR U4960 ( .A(n2940), .B(n2941), .Z(n2939) );
  OR U4961 ( .A(n2942), .B(n2943), .Z(n2938) );
  NAND U4962 ( .A(n2944), .B(n2945), .Z(n2867) );
  OR U4963 ( .A(n2946), .B(n2947), .Z(n2945) );
  OR U4964 ( .A(n2948), .B(n2949), .Z(n2944) );
  NOR U4965 ( .A(n2950), .B(n2951), .Z(n2868) );
  ANDN U4966 ( .B(n2952), .A(n2953), .Z(n2862) );
  IV U4967 ( .A(n2954), .Z(n2952) );
  XNOR U4968 ( .A(n2855), .B(n2955), .Z(n2861) );
  XNOR U4969 ( .A(n2854), .B(n2856), .Z(n2955) );
  NAND U4970 ( .A(n2956), .B(n2957), .Z(n2856) );
  OR U4971 ( .A(n2958), .B(n2959), .Z(n2957) );
  OR U4972 ( .A(n2960), .B(n2961), .Z(n2956) );
  NAND U4973 ( .A(n2962), .B(n2963), .Z(n2854) );
  OR U4974 ( .A(n2964), .B(n2965), .Z(n2963) );
  OR U4975 ( .A(n2966), .B(n2967), .Z(n2962) );
  ANDN U4976 ( .B(n2968), .A(n2969), .Z(n2855) );
  IV U4977 ( .A(n2970), .Z(n2968) );
  XNOR U4978 ( .A(n2935), .B(n2934), .Z(N13573) );
  XOR U4979 ( .A(n2954), .B(n2953), .Z(n2934) );
  XNOR U4980 ( .A(n2969), .B(n2970), .Z(n2953) );
  XNOR U4981 ( .A(n2964), .B(n2965), .Z(n2970) );
  XNOR U4982 ( .A(n2966), .B(n2967), .Z(n2965) );
  XNOR U4983 ( .A(y[1741]), .B(x[1741]), .Z(n2967) );
  XNOR U4984 ( .A(y[1742]), .B(x[1742]), .Z(n2966) );
  XNOR U4985 ( .A(y[1740]), .B(x[1740]), .Z(n2964) );
  XNOR U4986 ( .A(n2958), .B(n2959), .Z(n2969) );
  XNOR U4987 ( .A(y[1737]), .B(x[1737]), .Z(n2959) );
  XNOR U4988 ( .A(n2960), .B(n2961), .Z(n2958) );
  XNOR U4989 ( .A(y[1738]), .B(x[1738]), .Z(n2961) );
  XNOR U4990 ( .A(y[1739]), .B(x[1739]), .Z(n2960) );
  XNOR U4991 ( .A(n2951), .B(n2950), .Z(n2954) );
  XNOR U4992 ( .A(n2946), .B(n2947), .Z(n2950) );
  XNOR U4993 ( .A(y[1734]), .B(x[1734]), .Z(n2947) );
  XNOR U4994 ( .A(n2948), .B(n2949), .Z(n2946) );
  XNOR U4995 ( .A(y[1735]), .B(x[1735]), .Z(n2949) );
  XNOR U4996 ( .A(y[1736]), .B(x[1736]), .Z(n2948) );
  XNOR U4997 ( .A(n2940), .B(n2941), .Z(n2951) );
  XNOR U4998 ( .A(y[1731]), .B(x[1731]), .Z(n2941) );
  XNOR U4999 ( .A(n2942), .B(n2943), .Z(n2940) );
  XNOR U5000 ( .A(y[1732]), .B(x[1732]), .Z(n2943) );
  XNOR U5001 ( .A(y[1733]), .B(x[1733]), .Z(n2942) );
  XOR U5002 ( .A(n2916), .B(n2917), .Z(n2935) );
  XNOR U5003 ( .A(n2932), .B(n2933), .Z(n2917) );
  XNOR U5004 ( .A(n2927), .B(n2928), .Z(n2933) );
  XNOR U5005 ( .A(n2929), .B(n2930), .Z(n2928) );
  XNOR U5006 ( .A(y[1729]), .B(x[1729]), .Z(n2930) );
  XNOR U5007 ( .A(y[1730]), .B(x[1730]), .Z(n2929) );
  XNOR U5008 ( .A(y[1728]), .B(x[1728]), .Z(n2927) );
  XNOR U5009 ( .A(n2921), .B(n2922), .Z(n2932) );
  XNOR U5010 ( .A(y[1725]), .B(x[1725]), .Z(n2922) );
  XNOR U5011 ( .A(n2923), .B(n2924), .Z(n2921) );
  XNOR U5012 ( .A(y[1726]), .B(x[1726]), .Z(n2924) );
  XNOR U5013 ( .A(y[1727]), .B(x[1727]), .Z(n2923) );
  XOR U5014 ( .A(n2915), .B(n2914), .Z(n2916) );
  XNOR U5015 ( .A(n2910), .B(n2911), .Z(n2914) );
  XNOR U5016 ( .A(y[1722]), .B(x[1722]), .Z(n2911) );
  XNOR U5017 ( .A(n2912), .B(n2913), .Z(n2910) );
  XNOR U5018 ( .A(y[1723]), .B(x[1723]), .Z(n2913) );
  XNOR U5019 ( .A(y[1724]), .B(x[1724]), .Z(n2912) );
  XNOR U5020 ( .A(n2904), .B(n2905), .Z(n2915) );
  XNOR U5021 ( .A(y[1719]), .B(x[1719]), .Z(n2905) );
  XNOR U5022 ( .A(n2906), .B(n2907), .Z(n2904) );
  XNOR U5023 ( .A(y[1720]), .B(x[1720]), .Z(n2907) );
  XNOR U5024 ( .A(y[1721]), .B(x[1721]), .Z(n2906) );
  NAND U5025 ( .A(n2971), .B(n2972), .Z(N13566) );
  NANDN U5026 ( .A(n2973), .B(n2974), .Z(n2972) );
  OR U5027 ( .A(n2975), .B(n2976), .Z(n2974) );
  NAND U5028 ( .A(n2975), .B(n2976), .Z(n2971) );
  XOR U5029 ( .A(n2975), .B(n2977), .Z(N13565) );
  XNOR U5030 ( .A(n2973), .B(n2976), .Z(n2977) );
  AND U5031 ( .A(n2978), .B(n2979), .Z(n2976) );
  NANDN U5032 ( .A(n2980), .B(n2981), .Z(n2979) );
  NANDN U5033 ( .A(n2982), .B(n2983), .Z(n2981) );
  NANDN U5034 ( .A(n2983), .B(n2982), .Z(n2978) );
  NAND U5035 ( .A(n2984), .B(n2985), .Z(n2973) );
  NANDN U5036 ( .A(n2986), .B(n2987), .Z(n2985) );
  OR U5037 ( .A(n2988), .B(n2989), .Z(n2987) );
  NAND U5038 ( .A(n2989), .B(n2988), .Z(n2984) );
  AND U5039 ( .A(n2990), .B(n2991), .Z(n2975) );
  NANDN U5040 ( .A(n2992), .B(n2993), .Z(n2991) );
  NANDN U5041 ( .A(n2994), .B(n2995), .Z(n2993) );
  NANDN U5042 ( .A(n2995), .B(n2994), .Z(n2990) );
  XOR U5043 ( .A(n2989), .B(n2996), .Z(N13564) );
  XOR U5044 ( .A(n2986), .B(n2988), .Z(n2996) );
  XNOR U5045 ( .A(n2982), .B(n2997), .Z(n2988) );
  XNOR U5046 ( .A(n2980), .B(n2983), .Z(n2997) );
  NAND U5047 ( .A(n2998), .B(n2999), .Z(n2983) );
  NAND U5048 ( .A(n3000), .B(n3001), .Z(n2999) );
  OR U5049 ( .A(n3002), .B(n3003), .Z(n3000) );
  NANDN U5050 ( .A(n3004), .B(n3002), .Z(n2998) );
  IV U5051 ( .A(n3003), .Z(n3004) );
  NAND U5052 ( .A(n3005), .B(n3006), .Z(n2980) );
  NAND U5053 ( .A(n3007), .B(n3008), .Z(n3006) );
  NANDN U5054 ( .A(n3009), .B(n3010), .Z(n3007) );
  NANDN U5055 ( .A(n3010), .B(n3009), .Z(n3005) );
  AND U5056 ( .A(n3011), .B(n3012), .Z(n2982) );
  NAND U5057 ( .A(n3013), .B(n3014), .Z(n3012) );
  OR U5058 ( .A(n3015), .B(n3016), .Z(n3013) );
  NANDN U5059 ( .A(n3017), .B(n3015), .Z(n3011) );
  NAND U5060 ( .A(n3018), .B(n3019), .Z(n2986) );
  NANDN U5061 ( .A(n3020), .B(n3021), .Z(n3019) );
  OR U5062 ( .A(n3022), .B(n3023), .Z(n3021) );
  NANDN U5063 ( .A(n3024), .B(n3022), .Z(n3018) );
  IV U5064 ( .A(n3023), .Z(n3024) );
  XNOR U5065 ( .A(n2994), .B(n3025), .Z(n2989) );
  XNOR U5066 ( .A(n2992), .B(n2995), .Z(n3025) );
  NAND U5067 ( .A(n3026), .B(n3027), .Z(n2995) );
  NAND U5068 ( .A(n3028), .B(n3029), .Z(n3027) );
  OR U5069 ( .A(n3030), .B(n3031), .Z(n3028) );
  NANDN U5070 ( .A(n3032), .B(n3030), .Z(n3026) );
  IV U5071 ( .A(n3031), .Z(n3032) );
  NAND U5072 ( .A(n3033), .B(n3034), .Z(n2992) );
  NAND U5073 ( .A(n3035), .B(n3036), .Z(n3034) );
  NANDN U5074 ( .A(n3037), .B(n3038), .Z(n3035) );
  NANDN U5075 ( .A(n3038), .B(n3037), .Z(n3033) );
  AND U5076 ( .A(n3039), .B(n3040), .Z(n2994) );
  NAND U5077 ( .A(n3041), .B(n3042), .Z(n3040) );
  OR U5078 ( .A(n3043), .B(n3044), .Z(n3041) );
  NANDN U5079 ( .A(n3045), .B(n3043), .Z(n3039) );
  XNOR U5080 ( .A(n3020), .B(n3046), .Z(N13563) );
  XOR U5081 ( .A(n3022), .B(n3023), .Z(n3046) );
  XNOR U5082 ( .A(n3036), .B(n3047), .Z(n3023) );
  XOR U5083 ( .A(n3037), .B(n3038), .Z(n3047) );
  XOR U5084 ( .A(n3043), .B(n3048), .Z(n3038) );
  XOR U5085 ( .A(n3042), .B(n3045), .Z(n3048) );
  IV U5086 ( .A(n3044), .Z(n3045) );
  NAND U5087 ( .A(n3049), .B(n3050), .Z(n3044) );
  OR U5088 ( .A(n3051), .B(n3052), .Z(n3050) );
  OR U5089 ( .A(n3053), .B(n3054), .Z(n3049) );
  NAND U5090 ( .A(n3055), .B(n3056), .Z(n3042) );
  OR U5091 ( .A(n3057), .B(n3058), .Z(n3056) );
  OR U5092 ( .A(n3059), .B(n3060), .Z(n3055) );
  NOR U5093 ( .A(n3061), .B(n3062), .Z(n3043) );
  ANDN U5094 ( .B(n3063), .A(n3064), .Z(n3037) );
  XNOR U5095 ( .A(n3030), .B(n3065), .Z(n3036) );
  XNOR U5096 ( .A(n3029), .B(n3031), .Z(n3065) );
  NAND U5097 ( .A(n3066), .B(n3067), .Z(n3031) );
  OR U5098 ( .A(n3068), .B(n3069), .Z(n3067) );
  OR U5099 ( .A(n3070), .B(n3071), .Z(n3066) );
  NAND U5100 ( .A(n3072), .B(n3073), .Z(n3029) );
  OR U5101 ( .A(n3074), .B(n3075), .Z(n3073) );
  OR U5102 ( .A(n3076), .B(n3077), .Z(n3072) );
  ANDN U5103 ( .B(n3078), .A(n3079), .Z(n3030) );
  IV U5104 ( .A(n3080), .Z(n3078) );
  ANDN U5105 ( .B(n3081), .A(n3082), .Z(n3022) );
  XOR U5106 ( .A(n3008), .B(n3083), .Z(n3020) );
  XOR U5107 ( .A(n3009), .B(n3010), .Z(n3083) );
  XOR U5108 ( .A(n3015), .B(n3084), .Z(n3010) );
  XOR U5109 ( .A(n3014), .B(n3017), .Z(n3084) );
  IV U5110 ( .A(n3016), .Z(n3017) );
  NAND U5111 ( .A(n3085), .B(n3086), .Z(n3016) );
  OR U5112 ( .A(n3087), .B(n3088), .Z(n3086) );
  OR U5113 ( .A(n3089), .B(n3090), .Z(n3085) );
  NAND U5114 ( .A(n3091), .B(n3092), .Z(n3014) );
  OR U5115 ( .A(n3093), .B(n3094), .Z(n3092) );
  OR U5116 ( .A(n3095), .B(n3096), .Z(n3091) );
  NOR U5117 ( .A(n3097), .B(n3098), .Z(n3015) );
  ANDN U5118 ( .B(n3099), .A(n3100), .Z(n3009) );
  IV U5119 ( .A(n3101), .Z(n3099) );
  XNOR U5120 ( .A(n3002), .B(n3102), .Z(n3008) );
  XNOR U5121 ( .A(n3001), .B(n3003), .Z(n3102) );
  NAND U5122 ( .A(n3103), .B(n3104), .Z(n3003) );
  OR U5123 ( .A(n3105), .B(n3106), .Z(n3104) );
  OR U5124 ( .A(n3107), .B(n3108), .Z(n3103) );
  NAND U5125 ( .A(n3109), .B(n3110), .Z(n3001) );
  OR U5126 ( .A(n3111), .B(n3112), .Z(n3110) );
  OR U5127 ( .A(n3113), .B(n3114), .Z(n3109) );
  ANDN U5128 ( .B(n3115), .A(n3116), .Z(n3002) );
  IV U5129 ( .A(n3117), .Z(n3115) );
  XNOR U5130 ( .A(n3082), .B(n3081), .Z(N13562) );
  XOR U5131 ( .A(n3101), .B(n3100), .Z(n3081) );
  XNOR U5132 ( .A(n3116), .B(n3117), .Z(n3100) );
  XNOR U5133 ( .A(n3111), .B(n3112), .Z(n3117) );
  XNOR U5134 ( .A(n3113), .B(n3114), .Z(n3112) );
  XNOR U5135 ( .A(y[1717]), .B(x[1717]), .Z(n3114) );
  XNOR U5136 ( .A(y[1718]), .B(x[1718]), .Z(n3113) );
  XNOR U5137 ( .A(y[1716]), .B(x[1716]), .Z(n3111) );
  XNOR U5138 ( .A(n3105), .B(n3106), .Z(n3116) );
  XNOR U5139 ( .A(y[1713]), .B(x[1713]), .Z(n3106) );
  XNOR U5140 ( .A(n3107), .B(n3108), .Z(n3105) );
  XNOR U5141 ( .A(y[1714]), .B(x[1714]), .Z(n3108) );
  XNOR U5142 ( .A(y[1715]), .B(x[1715]), .Z(n3107) );
  XNOR U5143 ( .A(n3098), .B(n3097), .Z(n3101) );
  XNOR U5144 ( .A(n3093), .B(n3094), .Z(n3097) );
  XNOR U5145 ( .A(y[1710]), .B(x[1710]), .Z(n3094) );
  XNOR U5146 ( .A(n3095), .B(n3096), .Z(n3093) );
  XNOR U5147 ( .A(y[1711]), .B(x[1711]), .Z(n3096) );
  XNOR U5148 ( .A(y[1712]), .B(x[1712]), .Z(n3095) );
  XNOR U5149 ( .A(n3087), .B(n3088), .Z(n3098) );
  XNOR U5150 ( .A(y[1707]), .B(x[1707]), .Z(n3088) );
  XNOR U5151 ( .A(n3089), .B(n3090), .Z(n3087) );
  XNOR U5152 ( .A(y[1708]), .B(x[1708]), .Z(n3090) );
  XNOR U5153 ( .A(y[1709]), .B(x[1709]), .Z(n3089) );
  XOR U5154 ( .A(n3063), .B(n3064), .Z(n3082) );
  XNOR U5155 ( .A(n3079), .B(n3080), .Z(n3064) );
  XNOR U5156 ( .A(n3074), .B(n3075), .Z(n3080) );
  XNOR U5157 ( .A(n3076), .B(n3077), .Z(n3075) );
  XNOR U5158 ( .A(y[1705]), .B(x[1705]), .Z(n3077) );
  XNOR U5159 ( .A(y[1706]), .B(x[1706]), .Z(n3076) );
  XNOR U5160 ( .A(y[1704]), .B(x[1704]), .Z(n3074) );
  XNOR U5161 ( .A(n3068), .B(n3069), .Z(n3079) );
  XNOR U5162 ( .A(y[1701]), .B(x[1701]), .Z(n3069) );
  XNOR U5163 ( .A(n3070), .B(n3071), .Z(n3068) );
  XNOR U5164 ( .A(y[1702]), .B(x[1702]), .Z(n3071) );
  XNOR U5165 ( .A(y[1703]), .B(x[1703]), .Z(n3070) );
  XOR U5166 ( .A(n3062), .B(n3061), .Z(n3063) );
  XNOR U5167 ( .A(n3057), .B(n3058), .Z(n3061) );
  XNOR U5168 ( .A(y[1698]), .B(x[1698]), .Z(n3058) );
  XNOR U5169 ( .A(n3059), .B(n3060), .Z(n3057) );
  XNOR U5170 ( .A(y[1699]), .B(x[1699]), .Z(n3060) );
  XNOR U5171 ( .A(y[1700]), .B(x[1700]), .Z(n3059) );
  XNOR U5172 ( .A(n3051), .B(n3052), .Z(n3062) );
  XNOR U5173 ( .A(y[1695]), .B(x[1695]), .Z(n3052) );
  XNOR U5174 ( .A(n3053), .B(n3054), .Z(n3051) );
  XNOR U5175 ( .A(y[1696]), .B(x[1696]), .Z(n3054) );
  XNOR U5176 ( .A(y[1697]), .B(x[1697]), .Z(n3053) );
  NAND U5177 ( .A(n3118), .B(n3119), .Z(N13555) );
  NANDN U5178 ( .A(n3120), .B(n3121), .Z(n3119) );
  OR U5179 ( .A(n3122), .B(n3123), .Z(n3121) );
  NAND U5180 ( .A(n3122), .B(n3123), .Z(n3118) );
  XOR U5181 ( .A(n3122), .B(n3124), .Z(N13554) );
  XNOR U5182 ( .A(n3120), .B(n3123), .Z(n3124) );
  AND U5183 ( .A(n3125), .B(n3126), .Z(n3123) );
  NANDN U5184 ( .A(n3127), .B(n3128), .Z(n3126) );
  NANDN U5185 ( .A(n3129), .B(n3130), .Z(n3128) );
  NANDN U5186 ( .A(n3130), .B(n3129), .Z(n3125) );
  NAND U5187 ( .A(n3131), .B(n3132), .Z(n3120) );
  NANDN U5188 ( .A(n3133), .B(n3134), .Z(n3132) );
  OR U5189 ( .A(n3135), .B(n3136), .Z(n3134) );
  NAND U5190 ( .A(n3136), .B(n3135), .Z(n3131) );
  AND U5191 ( .A(n3137), .B(n3138), .Z(n3122) );
  NANDN U5192 ( .A(n3139), .B(n3140), .Z(n3138) );
  NANDN U5193 ( .A(n3141), .B(n3142), .Z(n3140) );
  NANDN U5194 ( .A(n3142), .B(n3141), .Z(n3137) );
  XOR U5195 ( .A(n3136), .B(n3143), .Z(N13553) );
  XOR U5196 ( .A(n3133), .B(n3135), .Z(n3143) );
  XNOR U5197 ( .A(n3129), .B(n3144), .Z(n3135) );
  XNOR U5198 ( .A(n3127), .B(n3130), .Z(n3144) );
  NAND U5199 ( .A(n3145), .B(n3146), .Z(n3130) );
  NAND U5200 ( .A(n3147), .B(n3148), .Z(n3146) );
  OR U5201 ( .A(n3149), .B(n3150), .Z(n3147) );
  NANDN U5202 ( .A(n3151), .B(n3149), .Z(n3145) );
  IV U5203 ( .A(n3150), .Z(n3151) );
  NAND U5204 ( .A(n3152), .B(n3153), .Z(n3127) );
  NAND U5205 ( .A(n3154), .B(n3155), .Z(n3153) );
  NANDN U5206 ( .A(n3156), .B(n3157), .Z(n3154) );
  NANDN U5207 ( .A(n3157), .B(n3156), .Z(n3152) );
  AND U5208 ( .A(n3158), .B(n3159), .Z(n3129) );
  NAND U5209 ( .A(n3160), .B(n3161), .Z(n3159) );
  OR U5210 ( .A(n3162), .B(n3163), .Z(n3160) );
  NANDN U5211 ( .A(n3164), .B(n3162), .Z(n3158) );
  NAND U5212 ( .A(n3165), .B(n3166), .Z(n3133) );
  NANDN U5213 ( .A(n3167), .B(n3168), .Z(n3166) );
  OR U5214 ( .A(n3169), .B(n3170), .Z(n3168) );
  NANDN U5215 ( .A(n3171), .B(n3169), .Z(n3165) );
  IV U5216 ( .A(n3170), .Z(n3171) );
  XNOR U5217 ( .A(n3141), .B(n3172), .Z(n3136) );
  XNOR U5218 ( .A(n3139), .B(n3142), .Z(n3172) );
  NAND U5219 ( .A(n3173), .B(n3174), .Z(n3142) );
  NAND U5220 ( .A(n3175), .B(n3176), .Z(n3174) );
  OR U5221 ( .A(n3177), .B(n3178), .Z(n3175) );
  NANDN U5222 ( .A(n3179), .B(n3177), .Z(n3173) );
  IV U5223 ( .A(n3178), .Z(n3179) );
  NAND U5224 ( .A(n3180), .B(n3181), .Z(n3139) );
  NAND U5225 ( .A(n3182), .B(n3183), .Z(n3181) );
  NANDN U5226 ( .A(n3184), .B(n3185), .Z(n3182) );
  NANDN U5227 ( .A(n3185), .B(n3184), .Z(n3180) );
  AND U5228 ( .A(n3186), .B(n3187), .Z(n3141) );
  NAND U5229 ( .A(n3188), .B(n3189), .Z(n3187) );
  OR U5230 ( .A(n3190), .B(n3191), .Z(n3188) );
  NANDN U5231 ( .A(n3192), .B(n3190), .Z(n3186) );
  XNOR U5232 ( .A(n3167), .B(n3193), .Z(N13552) );
  XOR U5233 ( .A(n3169), .B(n3170), .Z(n3193) );
  XNOR U5234 ( .A(n3183), .B(n3194), .Z(n3170) );
  XOR U5235 ( .A(n3184), .B(n3185), .Z(n3194) );
  XOR U5236 ( .A(n3190), .B(n3195), .Z(n3185) );
  XOR U5237 ( .A(n3189), .B(n3192), .Z(n3195) );
  IV U5238 ( .A(n3191), .Z(n3192) );
  NAND U5239 ( .A(n3196), .B(n3197), .Z(n3191) );
  OR U5240 ( .A(n3198), .B(n3199), .Z(n3197) );
  OR U5241 ( .A(n3200), .B(n3201), .Z(n3196) );
  NAND U5242 ( .A(n3202), .B(n3203), .Z(n3189) );
  OR U5243 ( .A(n3204), .B(n3205), .Z(n3203) );
  OR U5244 ( .A(n3206), .B(n3207), .Z(n3202) );
  NOR U5245 ( .A(n3208), .B(n3209), .Z(n3190) );
  ANDN U5246 ( .B(n3210), .A(n3211), .Z(n3184) );
  XNOR U5247 ( .A(n3177), .B(n3212), .Z(n3183) );
  XNOR U5248 ( .A(n3176), .B(n3178), .Z(n3212) );
  NAND U5249 ( .A(n3213), .B(n3214), .Z(n3178) );
  OR U5250 ( .A(n3215), .B(n3216), .Z(n3214) );
  OR U5251 ( .A(n3217), .B(n3218), .Z(n3213) );
  NAND U5252 ( .A(n3219), .B(n3220), .Z(n3176) );
  OR U5253 ( .A(n3221), .B(n3222), .Z(n3220) );
  OR U5254 ( .A(n3223), .B(n3224), .Z(n3219) );
  ANDN U5255 ( .B(n3225), .A(n3226), .Z(n3177) );
  IV U5256 ( .A(n3227), .Z(n3225) );
  ANDN U5257 ( .B(n3228), .A(n3229), .Z(n3169) );
  XOR U5258 ( .A(n3155), .B(n3230), .Z(n3167) );
  XOR U5259 ( .A(n3156), .B(n3157), .Z(n3230) );
  XOR U5260 ( .A(n3162), .B(n3231), .Z(n3157) );
  XOR U5261 ( .A(n3161), .B(n3164), .Z(n3231) );
  IV U5262 ( .A(n3163), .Z(n3164) );
  NAND U5263 ( .A(n3232), .B(n3233), .Z(n3163) );
  OR U5264 ( .A(n3234), .B(n3235), .Z(n3233) );
  OR U5265 ( .A(n3236), .B(n3237), .Z(n3232) );
  NAND U5266 ( .A(n3238), .B(n3239), .Z(n3161) );
  OR U5267 ( .A(n3240), .B(n3241), .Z(n3239) );
  OR U5268 ( .A(n3242), .B(n3243), .Z(n3238) );
  NOR U5269 ( .A(n3244), .B(n3245), .Z(n3162) );
  ANDN U5270 ( .B(n3246), .A(n3247), .Z(n3156) );
  IV U5271 ( .A(n3248), .Z(n3246) );
  XNOR U5272 ( .A(n3149), .B(n3249), .Z(n3155) );
  XNOR U5273 ( .A(n3148), .B(n3150), .Z(n3249) );
  NAND U5274 ( .A(n3250), .B(n3251), .Z(n3150) );
  OR U5275 ( .A(n3252), .B(n3253), .Z(n3251) );
  OR U5276 ( .A(n3254), .B(n3255), .Z(n3250) );
  NAND U5277 ( .A(n3256), .B(n3257), .Z(n3148) );
  OR U5278 ( .A(n3258), .B(n3259), .Z(n3257) );
  OR U5279 ( .A(n3260), .B(n3261), .Z(n3256) );
  ANDN U5280 ( .B(n3262), .A(n3263), .Z(n3149) );
  IV U5281 ( .A(n3264), .Z(n3262) );
  XNOR U5282 ( .A(n3229), .B(n3228), .Z(N13551) );
  XOR U5283 ( .A(n3248), .B(n3247), .Z(n3228) );
  XNOR U5284 ( .A(n3263), .B(n3264), .Z(n3247) );
  XNOR U5285 ( .A(n3258), .B(n3259), .Z(n3264) );
  XNOR U5286 ( .A(n3260), .B(n3261), .Z(n3259) );
  XNOR U5287 ( .A(y[1693]), .B(x[1693]), .Z(n3261) );
  XNOR U5288 ( .A(y[1694]), .B(x[1694]), .Z(n3260) );
  XNOR U5289 ( .A(y[1692]), .B(x[1692]), .Z(n3258) );
  XNOR U5290 ( .A(n3252), .B(n3253), .Z(n3263) );
  XNOR U5291 ( .A(y[1689]), .B(x[1689]), .Z(n3253) );
  XNOR U5292 ( .A(n3254), .B(n3255), .Z(n3252) );
  XNOR U5293 ( .A(y[1690]), .B(x[1690]), .Z(n3255) );
  XNOR U5294 ( .A(y[1691]), .B(x[1691]), .Z(n3254) );
  XNOR U5295 ( .A(n3245), .B(n3244), .Z(n3248) );
  XNOR U5296 ( .A(n3240), .B(n3241), .Z(n3244) );
  XNOR U5297 ( .A(y[1686]), .B(x[1686]), .Z(n3241) );
  XNOR U5298 ( .A(n3242), .B(n3243), .Z(n3240) );
  XNOR U5299 ( .A(y[1687]), .B(x[1687]), .Z(n3243) );
  XNOR U5300 ( .A(y[1688]), .B(x[1688]), .Z(n3242) );
  XNOR U5301 ( .A(n3234), .B(n3235), .Z(n3245) );
  XNOR U5302 ( .A(y[1683]), .B(x[1683]), .Z(n3235) );
  XNOR U5303 ( .A(n3236), .B(n3237), .Z(n3234) );
  XNOR U5304 ( .A(y[1684]), .B(x[1684]), .Z(n3237) );
  XNOR U5305 ( .A(y[1685]), .B(x[1685]), .Z(n3236) );
  XOR U5306 ( .A(n3210), .B(n3211), .Z(n3229) );
  XNOR U5307 ( .A(n3226), .B(n3227), .Z(n3211) );
  XNOR U5308 ( .A(n3221), .B(n3222), .Z(n3227) );
  XNOR U5309 ( .A(n3223), .B(n3224), .Z(n3222) );
  XNOR U5310 ( .A(y[1681]), .B(x[1681]), .Z(n3224) );
  XNOR U5311 ( .A(y[1682]), .B(x[1682]), .Z(n3223) );
  XNOR U5312 ( .A(y[1680]), .B(x[1680]), .Z(n3221) );
  XNOR U5313 ( .A(n3215), .B(n3216), .Z(n3226) );
  XNOR U5314 ( .A(y[1677]), .B(x[1677]), .Z(n3216) );
  XNOR U5315 ( .A(n3217), .B(n3218), .Z(n3215) );
  XNOR U5316 ( .A(y[1678]), .B(x[1678]), .Z(n3218) );
  XNOR U5317 ( .A(y[1679]), .B(x[1679]), .Z(n3217) );
  XOR U5318 ( .A(n3209), .B(n3208), .Z(n3210) );
  XNOR U5319 ( .A(n3204), .B(n3205), .Z(n3208) );
  XNOR U5320 ( .A(y[1674]), .B(x[1674]), .Z(n3205) );
  XNOR U5321 ( .A(n3206), .B(n3207), .Z(n3204) );
  XNOR U5322 ( .A(y[1675]), .B(x[1675]), .Z(n3207) );
  XNOR U5323 ( .A(y[1676]), .B(x[1676]), .Z(n3206) );
  XNOR U5324 ( .A(n3198), .B(n3199), .Z(n3209) );
  XNOR U5325 ( .A(y[1671]), .B(x[1671]), .Z(n3199) );
  XNOR U5326 ( .A(n3200), .B(n3201), .Z(n3198) );
  XNOR U5327 ( .A(y[1672]), .B(x[1672]), .Z(n3201) );
  XNOR U5328 ( .A(y[1673]), .B(x[1673]), .Z(n3200) );
  NAND U5329 ( .A(n3265), .B(n3266), .Z(N13544) );
  NANDN U5330 ( .A(n3267), .B(n3268), .Z(n3266) );
  OR U5331 ( .A(n3269), .B(n3270), .Z(n3268) );
  NAND U5332 ( .A(n3269), .B(n3270), .Z(n3265) );
  XOR U5333 ( .A(n3269), .B(n3271), .Z(N13543) );
  XNOR U5334 ( .A(n3267), .B(n3270), .Z(n3271) );
  AND U5335 ( .A(n3272), .B(n3273), .Z(n3270) );
  NANDN U5336 ( .A(n3274), .B(n3275), .Z(n3273) );
  NANDN U5337 ( .A(n3276), .B(n3277), .Z(n3275) );
  NANDN U5338 ( .A(n3277), .B(n3276), .Z(n3272) );
  NAND U5339 ( .A(n3278), .B(n3279), .Z(n3267) );
  NANDN U5340 ( .A(n3280), .B(n3281), .Z(n3279) );
  OR U5341 ( .A(n3282), .B(n3283), .Z(n3281) );
  NAND U5342 ( .A(n3283), .B(n3282), .Z(n3278) );
  AND U5343 ( .A(n3284), .B(n3285), .Z(n3269) );
  NANDN U5344 ( .A(n3286), .B(n3287), .Z(n3285) );
  NANDN U5345 ( .A(n3288), .B(n3289), .Z(n3287) );
  NANDN U5346 ( .A(n3289), .B(n3288), .Z(n3284) );
  XOR U5347 ( .A(n3283), .B(n3290), .Z(N13542) );
  XOR U5348 ( .A(n3280), .B(n3282), .Z(n3290) );
  XNOR U5349 ( .A(n3276), .B(n3291), .Z(n3282) );
  XNOR U5350 ( .A(n3274), .B(n3277), .Z(n3291) );
  NAND U5351 ( .A(n3292), .B(n3293), .Z(n3277) );
  NAND U5352 ( .A(n3294), .B(n3295), .Z(n3293) );
  OR U5353 ( .A(n3296), .B(n3297), .Z(n3294) );
  NANDN U5354 ( .A(n3298), .B(n3296), .Z(n3292) );
  IV U5355 ( .A(n3297), .Z(n3298) );
  NAND U5356 ( .A(n3299), .B(n3300), .Z(n3274) );
  NAND U5357 ( .A(n3301), .B(n3302), .Z(n3300) );
  NANDN U5358 ( .A(n3303), .B(n3304), .Z(n3301) );
  NANDN U5359 ( .A(n3304), .B(n3303), .Z(n3299) );
  AND U5360 ( .A(n3305), .B(n3306), .Z(n3276) );
  NAND U5361 ( .A(n3307), .B(n3308), .Z(n3306) );
  OR U5362 ( .A(n3309), .B(n3310), .Z(n3307) );
  NANDN U5363 ( .A(n3311), .B(n3309), .Z(n3305) );
  NAND U5364 ( .A(n3312), .B(n3313), .Z(n3280) );
  NANDN U5365 ( .A(n3314), .B(n3315), .Z(n3313) );
  OR U5366 ( .A(n3316), .B(n3317), .Z(n3315) );
  NANDN U5367 ( .A(n3318), .B(n3316), .Z(n3312) );
  IV U5368 ( .A(n3317), .Z(n3318) );
  XNOR U5369 ( .A(n3288), .B(n3319), .Z(n3283) );
  XNOR U5370 ( .A(n3286), .B(n3289), .Z(n3319) );
  NAND U5371 ( .A(n3320), .B(n3321), .Z(n3289) );
  NAND U5372 ( .A(n3322), .B(n3323), .Z(n3321) );
  OR U5373 ( .A(n3324), .B(n3325), .Z(n3322) );
  NANDN U5374 ( .A(n3326), .B(n3324), .Z(n3320) );
  IV U5375 ( .A(n3325), .Z(n3326) );
  NAND U5376 ( .A(n3327), .B(n3328), .Z(n3286) );
  NAND U5377 ( .A(n3329), .B(n3330), .Z(n3328) );
  NANDN U5378 ( .A(n3331), .B(n3332), .Z(n3329) );
  NANDN U5379 ( .A(n3332), .B(n3331), .Z(n3327) );
  AND U5380 ( .A(n3333), .B(n3334), .Z(n3288) );
  NAND U5381 ( .A(n3335), .B(n3336), .Z(n3334) );
  OR U5382 ( .A(n3337), .B(n3338), .Z(n3335) );
  NANDN U5383 ( .A(n3339), .B(n3337), .Z(n3333) );
  XNOR U5384 ( .A(n3314), .B(n3340), .Z(N13541) );
  XOR U5385 ( .A(n3316), .B(n3317), .Z(n3340) );
  XNOR U5386 ( .A(n3330), .B(n3341), .Z(n3317) );
  XOR U5387 ( .A(n3331), .B(n3332), .Z(n3341) );
  XOR U5388 ( .A(n3337), .B(n3342), .Z(n3332) );
  XOR U5389 ( .A(n3336), .B(n3339), .Z(n3342) );
  IV U5390 ( .A(n3338), .Z(n3339) );
  NAND U5391 ( .A(n3343), .B(n3344), .Z(n3338) );
  OR U5392 ( .A(n3345), .B(n3346), .Z(n3344) );
  OR U5393 ( .A(n3347), .B(n3348), .Z(n3343) );
  NAND U5394 ( .A(n3349), .B(n3350), .Z(n3336) );
  OR U5395 ( .A(n3351), .B(n3352), .Z(n3350) );
  OR U5396 ( .A(n3353), .B(n3354), .Z(n3349) );
  NOR U5397 ( .A(n3355), .B(n3356), .Z(n3337) );
  ANDN U5398 ( .B(n3357), .A(n3358), .Z(n3331) );
  XNOR U5399 ( .A(n3324), .B(n3359), .Z(n3330) );
  XNOR U5400 ( .A(n3323), .B(n3325), .Z(n3359) );
  NAND U5401 ( .A(n3360), .B(n3361), .Z(n3325) );
  OR U5402 ( .A(n3362), .B(n3363), .Z(n3361) );
  OR U5403 ( .A(n3364), .B(n3365), .Z(n3360) );
  NAND U5404 ( .A(n3366), .B(n3367), .Z(n3323) );
  OR U5405 ( .A(n3368), .B(n3369), .Z(n3367) );
  OR U5406 ( .A(n3370), .B(n3371), .Z(n3366) );
  ANDN U5407 ( .B(n3372), .A(n3373), .Z(n3324) );
  IV U5408 ( .A(n3374), .Z(n3372) );
  ANDN U5409 ( .B(n3375), .A(n3376), .Z(n3316) );
  XOR U5410 ( .A(n3302), .B(n3377), .Z(n3314) );
  XOR U5411 ( .A(n3303), .B(n3304), .Z(n3377) );
  XOR U5412 ( .A(n3309), .B(n3378), .Z(n3304) );
  XOR U5413 ( .A(n3308), .B(n3311), .Z(n3378) );
  IV U5414 ( .A(n3310), .Z(n3311) );
  NAND U5415 ( .A(n3379), .B(n3380), .Z(n3310) );
  OR U5416 ( .A(n3381), .B(n3382), .Z(n3380) );
  OR U5417 ( .A(n3383), .B(n3384), .Z(n3379) );
  NAND U5418 ( .A(n3385), .B(n3386), .Z(n3308) );
  OR U5419 ( .A(n3387), .B(n3388), .Z(n3386) );
  OR U5420 ( .A(n3389), .B(n3390), .Z(n3385) );
  NOR U5421 ( .A(n3391), .B(n3392), .Z(n3309) );
  ANDN U5422 ( .B(n3393), .A(n3394), .Z(n3303) );
  IV U5423 ( .A(n3395), .Z(n3393) );
  XNOR U5424 ( .A(n3296), .B(n3396), .Z(n3302) );
  XNOR U5425 ( .A(n3295), .B(n3297), .Z(n3396) );
  NAND U5426 ( .A(n3397), .B(n3398), .Z(n3297) );
  OR U5427 ( .A(n3399), .B(n3400), .Z(n3398) );
  OR U5428 ( .A(n3401), .B(n3402), .Z(n3397) );
  NAND U5429 ( .A(n3403), .B(n3404), .Z(n3295) );
  OR U5430 ( .A(n3405), .B(n3406), .Z(n3404) );
  OR U5431 ( .A(n3407), .B(n3408), .Z(n3403) );
  ANDN U5432 ( .B(n3409), .A(n3410), .Z(n3296) );
  IV U5433 ( .A(n3411), .Z(n3409) );
  XNOR U5434 ( .A(n3376), .B(n3375), .Z(N13540) );
  XOR U5435 ( .A(n3395), .B(n3394), .Z(n3375) );
  XNOR U5436 ( .A(n3410), .B(n3411), .Z(n3394) );
  XNOR U5437 ( .A(n3405), .B(n3406), .Z(n3411) );
  XNOR U5438 ( .A(n3407), .B(n3408), .Z(n3406) );
  XNOR U5439 ( .A(y[1669]), .B(x[1669]), .Z(n3408) );
  XNOR U5440 ( .A(y[1670]), .B(x[1670]), .Z(n3407) );
  XNOR U5441 ( .A(y[1668]), .B(x[1668]), .Z(n3405) );
  XNOR U5442 ( .A(n3399), .B(n3400), .Z(n3410) );
  XNOR U5443 ( .A(y[1665]), .B(x[1665]), .Z(n3400) );
  XNOR U5444 ( .A(n3401), .B(n3402), .Z(n3399) );
  XNOR U5445 ( .A(y[1666]), .B(x[1666]), .Z(n3402) );
  XNOR U5446 ( .A(y[1667]), .B(x[1667]), .Z(n3401) );
  XNOR U5447 ( .A(n3392), .B(n3391), .Z(n3395) );
  XNOR U5448 ( .A(n3387), .B(n3388), .Z(n3391) );
  XNOR U5449 ( .A(y[1662]), .B(x[1662]), .Z(n3388) );
  XNOR U5450 ( .A(n3389), .B(n3390), .Z(n3387) );
  XNOR U5451 ( .A(y[1663]), .B(x[1663]), .Z(n3390) );
  XNOR U5452 ( .A(y[1664]), .B(x[1664]), .Z(n3389) );
  XNOR U5453 ( .A(n3381), .B(n3382), .Z(n3392) );
  XNOR U5454 ( .A(y[1659]), .B(x[1659]), .Z(n3382) );
  XNOR U5455 ( .A(n3383), .B(n3384), .Z(n3381) );
  XNOR U5456 ( .A(y[1660]), .B(x[1660]), .Z(n3384) );
  XNOR U5457 ( .A(y[1661]), .B(x[1661]), .Z(n3383) );
  XOR U5458 ( .A(n3357), .B(n3358), .Z(n3376) );
  XNOR U5459 ( .A(n3373), .B(n3374), .Z(n3358) );
  XNOR U5460 ( .A(n3368), .B(n3369), .Z(n3374) );
  XNOR U5461 ( .A(n3370), .B(n3371), .Z(n3369) );
  XNOR U5462 ( .A(y[1657]), .B(x[1657]), .Z(n3371) );
  XNOR U5463 ( .A(y[1658]), .B(x[1658]), .Z(n3370) );
  XNOR U5464 ( .A(y[1656]), .B(x[1656]), .Z(n3368) );
  XNOR U5465 ( .A(n3362), .B(n3363), .Z(n3373) );
  XNOR U5466 ( .A(y[1653]), .B(x[1653]), .Z(n3363) );
  XNOR U5467 ( .A(n3364), .B(n3365), .Z(n3362) );
  XNOR U5468 ( .A(y[1654]), .B(x[1654]), .Z(n3365) );
  XNOR U5469 ( .A(y[1655]), .B(x[1655]), .Z(n3364) );
  XOR U5470 ( .A(n3356), .B(n3355), .Z(n3357) );
  XNOR U5471 ( .A(n3351), .B(n3352), .Z(n3355) );
  XNOR U5472 ( .A(y[1650]), .B(x[1650]), .Z(n3352) );
  XNOR U5473 ( .A(n3353), .B(n3354), .Z(n3351) );
  XNOR U5474 ( .A(y[1651]), .B(x[1651]), .Z(n3354) );
  XNOR U5475 ( .A(y[1652]), .B(x[1652]), .Z(n3353) );
  XNOR U5476 ( .A(n3345), .B(n3346), .Z(n3356) );
  XNOR U5477 ( .A(y[1647]), .B(x[1647]), .Z(n3346) );
  XNOR U5478 ( .A(n3347), .B(n3348), .Z(n3345) );
  XNOR U5479 ( .A(y[1648]), .B(x[1648]), .Z(n3348) );
  XNOR U5480 ( .A(y[1649]), .B(x[1649]), .Z(n3347) );
  NAND U5481 ( .A(n3412), .B(n3413), .Z(N13533) );
  NANDN U5482 ( .A(n3414), .B(n3415), .Z(n3413) );
  OR U5483 ( .A(n3416), .B(n3417), .Z(n3415) );
  NAND U5484 ( .A(n3416), .B(n3417), .Z(n3412) );
  XOR U5485 ( .A(n3416), .B(n3418), .Z(N13532) );
  XNOR U5486 ( .A(n3414), .B(n3417), .Z(n3418) );
  AND U5487 ( .A(n3419), .B(n3420), .Z(n3417) );
  NANDN U5488 ( .A(n3421), .B(n3422), .Z(n3420) );
  NANDN U5489 ( .A(n3423), .B(n3424), .Z(n3422) );
  NANDN U5490 ( .A(n3424), .B(n3423), .Z(n3419) );
  NAND U5491 ( .A(n3425), .B(n3426), .Z(n3414) );
  NANDN U5492 ( .A(n3427), .B(n3428), .Z(n3426) );
  OR U5493 ( .A(n3429), .B(n3430), .Z(n3428) );
  NAND U5494 ( .A(n3430), .B(n3429), .Z(n3425) );
  AND U5495 ( .A(n3431), .B(n3432), .Z(n3416) );
  NANDN U5496 ( .A(n3433), .B(n3434), .Z(n3432) );
  NANDN U5497 ( .A(n3435), .B(n3436), .Z(n3434) );
  NANDN U5498 ( .A(n3436), .B(n3435), .Z(n3431) );
  XOR U5499 ( .A(n3430), .B(n3437), .Z(N13531) );
  XOR U5500 ( .A(n3427), .B(n3429), .Z(n3437) );
  XNOR U5501 ( .A(n3423), .B(n3438), .Z(n3429) );
  XNOR U5502 ( .A(n3421), .B(n3424), .Z(n3438) );
  NAND U5503 ( .A(n3439), .B(n3440), .Z(n3424) );
  NAND U5504 ( .A(n3441), .B(n3442), .Z(n3440) );
  OR U5505 ( .A(n3443), .B(n3444), .Z(n3441) );
  NANDN U5506 ( .A(n3445), .B(n3443), .Z(n3439) );
  IV U5507 ( .A(n3444), .Z(n3445) );
  NAND U5508 ( .A(n3446), .B(n3447), .Z(n3421) );
  NAND U5509 ( .A(n3448), .B(n3449), .Z(n3447) );
  NANDN U5510 ( .A(n3450), .B(n3451), .Z(n3448) );
  NANDN U5511 ( .A(n3451), .B(n3450), .Z(n3446) );
  AND U5512 ( .A(n3452), .B(n3453), .Z(n3423) );
  NAND U5513 ( .A(n3454), .B(n3455), .Z(n3453) );
  OR U5514 ( .A(n3456), .B(n3457), .Z(n3454) );
  NANDN U5515 ( .A(n3458), .B(n3456), .Z(n3452) );
  NAND U5516 ( .A(n3459), .B(n3460), .Z(n3427) );
  NANDN U5517 ( .A(n3461), .B(n3462), .Z(n3460) );
  OR U5518 ( .A(n3463), .B(n3464), .Z(n3462) );
  NANDN U5519 ( .A(n3465), .B(n3463), .Z(n3459) );
  IV U5520 ( .A(n3464), .Z(n3465) );
  XNOR U5521 ( .A(n3435), .B(n3466), .Z(n3430) );
  XNOR U5522 ( .A(n3433), .B(n3436), .Z(n3466) );
  NAND U5523 ( .A(n3467), .B(n3468), .Z(n3436) );
  NAND U5524 ( .A(n3469), .B(n3470), .Z(n3468) );
  OR U5525 ( .A(n3471), .B(n3472), .Z(n3469) );
  NANDN U5526 ( .A(n3473), .B(n3471), .Z(n3467) );
  IV U5527 ( .A(n3472), .Z(n3473) );
  NAND U5528 ( .A(n3474), .B(n3475), .Z(n3433) );
  NAND U5529 ( .A(n3476), .B(n3477), .Z(n3475) );
  NANDN U5530 ( .A(n3478), .B(n3479), .Z(n3476) );
  NANDN U5531 ( .A(n3479), .B(n3478), .Z(n3474) );
  AND U5532 ( .A(n3480), .B(n3481), .Z(n3435) );
  NAND U5533 ( .A(n3482), .B(n3483), .Z(n3481) );
  OR U5534 ( .A(n3484), .B(n3485), .Z(n3482) );
  NANDN U5535 ( .A(n3486), .B(n3484), .Z(n3480) );
  XNOR U5536 ( .A(n3461), .B(n3487), .Z(N13530) );
  XOR U5537 ( .A(n3463), .B(n3464), .Z(n3487) );
  XNOR U5538 ( .A(n3477), .B(n3488), .Z(n3464) );
  XOR U5539 ( .A(n3478), .B(n3479), .Z(n3488) );
  XOR U5540 ( .A(n3484), .B(n3489), .Z(n3479) );
  XOR U5541 ( .A(n3483), .B(n3486), .Z(n3489) );
  IV U5542 ( .A(n3485), .Z(n3486) );
  NAND U5543 ( .A(n3490), .B(n3491), .Z(n3485) );
  OR U5544 ( .A(n3492), .B(n3493), .Z(n3491) );
  OR U5545 ( .A(n3494), .B(n3495), .Z(n3490) );
  NAND U5546 ( .A(n3496), .B(n3497), .Z(n3483) );
  OR U5547 ( .A(n3498), .B(n3499), .Z(n3497) );
  OR U5548 ( .A(n3500), .B(n3501), .Z(n3496) );
  NOR U5549 ( .A(n3502), .B(n3503), .Z(n3484) );
  ANDN U5550 ( .B(n3504), .A(n3505), .Z(n3478) );
  XNOR U5551 ( .A(n3471), .B(n3506), .Z(n3477) );
  XNOR U5552 ( .A(n3470), .B(n3472), .Z(n3506) );
  NAND U5553 ( .A(n3507), .B(n3508), .Z(n3472) );
  OR U5554 ( .A(n3509), .B(n3510), .Z(n3508) );
  OR U5555 ( .A(n3511), .B(n3512), .Z(n3507) );
  NAND U5556 ( .A(n3513), .B(n3514), .Z(n3470) );
  OR U5557 ( .A(n3515), .B(n3516), .Z(n3514) );
  OR U5558 ( .A(n3517), .B(n3518), .Z(n3513) );
  ANDN U5559 ( .B(n3519), .A(n3520), .Z(n3471) );
  IV U5560 ( .A(n3521), .Z(n3519) );
  ANDN U5561 ( .B(n3522), .A(n3523), .Z(n3463) );
  XOR U5562 ( .A(n3449), .B(n3524), .Z(n3461) );
  XOR U5563 ( .A(n3450), .B(n3451), .Z(n3524) );
  XOR U5564 ( .A(n3456), .B(n3525), .Z(n3451) );
  XOR U5565 ( .A(n3455), .B(n3458), .Z(n3525) );
  IV U5566 ( .A(n3457), .Z(n3458) );
  NAND U5567 ( .A(n3526), .B(n3527), .Z(n3457) );
  OR U5568 ( .A(n3528), .B(n3529), .Z(n3527) );
  OR U5569 ( .A(n3530), .B(n3531), .Z(n3526) );
  NAND U5570 ( .A(n3532), .B(n3533), .Z(n3455) );
  OR U5571 ( .A(n3534), .B(n3535), .Z(n3533) );
  OR U5572 ( .A(n3536), .B(n3537), .Z(n3532) );
  NOR U5573 ( .A(n3538), .B(n3539), .Z(n3456) );
  ANDN U5574 ( .B(n3540), .A(n3541), .Z(n3450) );
  IV U5575 ( .A(n3542), .Z(n3540) );
  XNOR U5576 ( .A(n3443), .B(n3543), .Z(n3449) );
  XNOR U5577 ( .A(n3442), .B(n3444), .Z(n3543) );
  NAND U5578 ( .A(n3544), .B(n3545), .Z(n3444) );
  OR U5579 ( .A(n3546), .B(n3547), .Z(n3545) );
  OR U5580 ( .A(n3548), .B(n3549), .Z(n3544) );
  NAND U5581 ( .A(n3550), .B(n3551), .Z(n3442) );
  OR U5582 ( .A(n3552), .B(n3553), .Z(n3551) );
  OR U5583 ( .A(n3554), .B(n3555), .Z(n3550) );
  ANDN U5584 ( .B(n3556), .A(n3557), .Z(n3443) );
  IV U5585 ( .A(n3558), .Z(n3556) );
  XNOR U5586 ( .A(n3523), .B(n3522), .Z(N13529) );
  XOR U5587 ( .A(n3542), .B(n3541), .Z(n3522) );
  XNOR U5588 ( .A(n3557), .B(n3558), .Z(n3541) );
  XNOR U5589 ( .A(n3552), .B(n3553), .Z(n3558) );
  XNOR U5590 ( .A(n3554), .B(n3555), .Z(n3553) );
  XNOR U5591 ( .A(y[1645]), .B(x[1645]), .Z(n3555) );
  XNOR U5592 ( .A(y[1646]), .B(x[1646]), .Z(n3554) );
  XNOR U5593 ( .A(y[1644]), .B(x[1644]), .Z(n3552) );
  XNOR U5594 ( .A(n3546), .B(n3547), .Z(n3557) );
  XNOR U5595 ( .A(y[1641]), .B(x[1641]), .Z(n3547) );
  XNOR U5596 ( .A(n3548), .B(n3549), .Z(n3546) );
  XNOR U5597 ( .A(y[1642]), .B(x[1642]), .Z(n3549) );
  XNOR U5598 ( .A(y[1643]), .B(x[1643]), .Z(n3548) );
  XNOR U5599 ( .A(n3539), .B(n3538), .Z(n3542) );
  XNOR U5600 ( .A(n3534), .B(n3535), .Z(n3538) );
  XNOR U5601 ( .A(y[1638]), .B(x[1638]), .Z(n3535) );
  XNOR U5602 ( .A(n3536), .B(n3537), .Z(n3534) );
  XNOR U5603 ( .A(y[1639]), .B(x[1639]), .Z(n3537) );
  XNOR U5604 ( .A(y[1640]), .B(x[1640]), .Z(n3536) );
  XNOR U5605 ( .A(n3528), .B(n3529), .Z(n3539) );
  XNOR U5606 ( .A(y[1635]), .B(x[1635]), .Z(n3529) );
  XNOR U5607 ( .A(n3530), .B(n3531), .Z(n3528) );
  XNOR U5608 ( .A(y[1636]), .B(x[1636]), .Z(n3531) );
  XNOR U5609 ( .A(y[1637]), .B(x[1637]), .Z(n3530) );
  XOR U5610 ( .A(n3504), .B(n3505), .Z(n3523) );
  XNOR U5611 ( .A(n3520), .B(n3521), .Z(n3505) );
  XNOR U5612 ( .A(n3515), .B(n3516), .Z(n3521) );
  XNOR U5613 ( .A(n3517), .B(n3518), .Z(n3516) );
  XNOR U5614 ( .A(y[1633]), .B(x[1633]), .Z(n3518) );
  XNOR U5615 ( .A(y[1634]), .B(x[1634]), .Z(n3517) );
  XNOR U5616 ( .A(y[1632]), .B(x[1632]), .Z(n3515) );
  XNOR U5617 ( .A(n3509), .B(n3510), .Z(n3520) );
  XNOR U5618 ( .A(y[1629]), .B(x[1629]), .Z(n3510) );
  XNOR U5619 ( .A(n3511), .B(n3512), .Z(n3509) );
  XNOR U5620 ( .A(y[1630]), .B(x[1630]), .Z(n3512) );
  XNOR U5621 ( .A(y[1631]), .B(x[1631]), .Z(n3511) );
  XOR U5622 ( .A(n3503), .B(n3502), .Z(n3504) );
  XNOR U5623 ( .A(n3498), .B(n3499), .Z(n3502) );
  XNOR U5624 ( .A(y[1626]), .B(x[1626]), .Z(n3499) );
  XNOR U5625 ( .A(n3500), .B(n3501), .Z(n3498) );
  XNOR U5626 ( .A(y[1627]), .B(x[1627]), .Z(n3501) );
  XNOR U5627 ( .A(y[1628]), .B(x[1628]), .Z(n3500) );
  XNOR U5628 ( .A(n3492), .B(n3493), .Z(n3503) );
  XNOR U5629 ( .A(y[1623]), .B(x[1623]), .Z(n3493) );
  XNOR U5630 ( .A(n3494), .B(n3495), .Z(n3492) );
  XNOR U5631 ( .A(y[1624]), .B(x[1624]), .Z(n3495) );
  XNOR U5632 ( .A(y[1625]), .B(x[1625]), .Z(n3494) );
  NAND U5633 ( .A(n3559), .B(n3560), .Z(N13522) );
  NANDN U5634 ( .A(n3561), .B(n3562), .Z(n3560) );
  OR U5635 ( .A(n3563), .B(n3564), .Z(n3562) );
  NAND U5636 ( .A(n3563), .B(n3564), .Z(n3559) );
  XOR U5637 ( .A(n3563), .B(n3565), .Z(N13521) );
  XNOR U5638 ( .A(n3561), .B(n3564), .Z(n3565) );
  AND U5639 ( .A(n3566), .B(n3567), .Z(n3564) );
  NANDN U5640 ( .A(n3568), .B(n3569), .Z(n3567) );
  NANDN U5641 ( .A(n3570), .B(n3571), .Z(n3569) );
  NANDN U5642 ( .A(n3571), .B(n3570), .Z(n3566) );
  NAND U5643 ( .A(n3572), .B(n3573), .Z(n3561) );
  NANDN U5644 ( .A(n3574), .B(n3575), .Z(n3573) );
  OR U5645 ( .A(n3576), .B(n3577), .Z(n3575) );
  NAND U5646 ( .A(n3577), .B(n3576), .Z(n3572) );
  AND U5647 ( .A(n3578), .B(n3579), .Z(n3563) );
  NANDN U5648 ( .A(n3580), .B(n3581), .Z(n3579) );
  NANDN U5649 ( .A(n3582), .B(n3583), .Z(n3581) );
  NANDN U5650 ( .A(n3583), .B(n3582), .Z(n3578) );
  XOR U5651 ( .A(n3577), .B(n3584), .Z(N13520) );
  XOR U5652 ( .A(n3574), .B(n3576), .Z(n3584) );
  XNOR U5653 ( .A(n3570), .B(n3585), .Z(n3576) );
  XNOR U5654 ( .A(n3568), .B(n3571), .Z(n3585) );
  NAND U5655 ( .A(n3586), .B(n3587), .Z(n3571) );
  NAND U5656 ( .A(n3588), .B(n3589), .Z(n3587) );
  OR U5657 ( .A(n3590), .B(n3591), .Z(n3588) );
  NANDN U5658 ( .A(n3592), .B(n3590), .Z(n3586) );
  IV U5659 ( .A(n3591), .Z(n3592) );
  NAND U5660 ( .A(n3593), .B(n3594), .Z(n3568) );
  NAND U5661 ( .A(n3595), .B(n3596), .Z(n3594) );
  NANDN U5662 ( .A(n3597), .B(n3598), .Z(n3595) );
  NANDN U5663 ( .A(n3598), .B(n3597), .Z(n3593) );
  AND U5664 ( .A(n3599), .B(n3600), .Z(n3570) );
  NAND U5665 ( .A(n3601), .B(n3602), .Z(n3600) );
  OR U5666 ( .A(n3603), .B(n3604), .Z(n3601) );
  NANDN U5667 ( .A(n3605), .B(n3603), .Z(n3599) );
  NAND U5668 ( .A(n3606), .B(n3607), .Z(n3574) );
  NANDN U5669 ( .A(n3608), .B(n3609), .Z(n3607) );
  OR U5670 ( .A(n3610), .B(n3611), .Z(n3609) );
  NANDN U5671 ( .A(n3612), .B(n3610), .Z(n3606) );
  IV U5672 ( .A(n3611), .Z(n3612) );
  XNOR U5673 ( .A(n3582), .B(n3613), .Z(n3577) );
  XNOR U5674 ( .A(n3580), .B(n3583), .Z(n3613) );
  NAND U5675 ( .A(n3614), .B(n3615), .Z(n3583) );
  NAND U5676 ( .A(n3616), .B(n3617), .Z(n3615) );
  OR U5677 ( .A(n3618), .B(n3619), .Z(n3616) );
  NANDN U5678 ( .A(n3620), .B(n3618), .Z(n3614) );
  IV U5679 ( .A(n3619), .Z(n3620) );
  NAND U5680 ( .A(n3621), .B(n3622), .Z(n3580) );
  NAND U5681 ( .A(n3623), .B(n3624), .Z(n3622) );
  NANDN U5682 ( .A(n3625), .B(n3626), .Z(n3623) );
  NANDN U5683 ( .A(n3626), .B(n3625), .Z(n3621) );
  AND U5684 ( .A(n3627), .B(n3628), .Z(n3582) );
  NAND U5685 ( .A(n3629), .B(n3630), .Z(n3628) );
  OR U5686 ( .A(n3631), .B(n3632), .Z(n3629) );
  NANDN U5687 ( .A(n3633), .B(n3631), .Z(n3627) );
  XNOR U5688 ( .A(n3608), .B(n3634), .Z(N13519) );
  XOR U5689 ( .A(n3610), .B(n3611), .Z(n3634) );
  XNOR U5690 ( .A(n3624), .B(n3635), .Z(n3611) );
  XOR U5691 ( .A(n3625), .B(n3626), .Z(n3635) );
  XOR U5692 ( .A(n3631), .B(n3636), .Z(n3626) );
  XOR U5693 ( .A(n3630), .B(n3633), .Z(n3636) );
  IV U5694 ( .A(n3632), .Z(n3633) );
  NAND U5695 ( .A(n3637), .B(n3638), .Z(n3632) );
  OR U5696 ( .A(n3639), .B(n3640), .Z(n3638) );
  OR U5697 ( .A(n3641), .B(n3642), .Z(n3637) );
  NAND U5698 ( .A(n3643), .B(n3644), .Z(n3630) );
  OR U5699 ( .A(n3645), .B(n3646), .Z(n3644) );
  OR U5700 ( .A(n3647), .B(n3648), .Z(n3643) );
  NOR U5701 ( .A(n3649), .B(n3650), .Z(n3631) );
  ANDN U5702 ( .B(n3651), .A(n3652), .Z(n3625) );
  XNOR U5703 ( .A(n3618), .B(n3653), .Z(n3624) );
  XNOR U5704 ( .A(n3617), .B(n3619), .Z(n3653) );
  NAND U5705 ( .A(n3654), .B(n3655), .Z(n3619) );
  OR U5706 ( .A(n3656), .B(n3657), .Z(n3655) );
  OR U5707 ( .A(n3658), .B(n3659), .Z(n3654) );
  NAND U5708 ( .A(n3660), .B(n3661), .Z(n3617) );
  OR U5709 ( .A(n3662), .B(n3663), .Z(n3661) );
  OR U5710 ( .A(n3664), .B(n3665), .Z(n3660) );
  ANDN U5711 ( .B(n3666), .A(n3667), .Z(n3618) );
  IV U5712 ( .A(n3668), .Z(n3666) );
  ANDN U5713 ( .B(n3669), .A(n3670), .Z(n3610) );
  XOR U5714 ( .A(n3596), .B(n3671), .Z(n3608) );
  XOR U5715 ( .A(n3597), .B(n3598), .Z(n3671) );
  XOR U5716 ( .A(n3603), .B(n3672), .Z(n3598) );
  XOR U5717 ( .A(n3602), .B(n3605), .Z(n3672) );
  IV U5718 ( .A(n3604), .Z(n3605) );
  NAND U5719 ( .A(n3673), .B(n3674), .Z(n3604) );
  OR U5720 ( .A(n3675), .B(n3676), .Z(n3674) );
  OR U5721 ( .A(n3677), .B(n3678), .Z(n3673) );
  NAND U5722 ( .A(n3679), .B(n3680), .Z(n3602) );
  OR U5723 ( .A(n3681), .B(n3682), .Z(n3680) );
  OR U5724 ( .A(n3683), .B(n3684), .Z(n3679) );
  NOR U5725 ( .A(n3685), .B(n3686), .Z(n3603) );
  ANDN U5726 ( .B(n3687), .A(n3688), .Z(n3597) );
  IV U5727 ( .A(n3689), .Z(n3687) );
  XNOR U5728 ( .A(n3590), .B(n3690), .Z(n3596) );
  XNOR U5729 ( .A(n3589), .B(n3591), .Z(n3690) );
  NAND U5730 ( .A(n3691), .B(n3692), .Z(n3591) );
  OR U5731 ( .A(n3693), .B(n3694), .Z(n3692) );
  OR U5732 ( .A(n3695), .B(n3696), .Z(n3691) );
  NAND U5733 ( .A(n3697), .B(n3698), .Z(n3589) );
  OR U5734 ( .A(n3699), .B(n3700), .Z(n3698) );
  OR U5735 ( .A(n3701), .B(n3702), .Z(n3697) );
  ANDN U5736 ( .B(n3703), .A(n3704), .Z(n3590) );
  IV U5737 ( .A(n3705), .Z(n3703) );
  XNOR U5738 ( .A(n3670), .B(n3669), .Z(N13518) );
  XOR U5739 ( .A(n3689), .B(n3688), .Z(n3669) );
  XNOR U5740 ( .A(n3704), .B(n3705), .Z(n3688) );
  XNOR U5741 ( .A(n3699), .B(n3700), .Z(n3705) );
  XNOR U5742 ( .A(n3701), .B(n3702), .Z(n3700) );
  XNOR U5743 ( .A(y[1621]), .B(x[1621]), .Z(n3702) );
  XNOR U5744 ( .A(y[1622]), .B(x[1622]), .Z(n3701) );
  XNOR U5745 ( .A(y[1620]), .B(x[1620]), .Z(n3699) );
  XNOR U5746 ( .A(n3693), .B(n3694), .Z(n3704) );
  XNOR U5747 ( .A(y[1617]), .B(x[1617]), .Z(n3694) );
  XNOR U5748 ( .A(n3695), .B(n3696), .Z(n3693) );
  XNOR U5749 ( .A(y[1618]), .B(x[1618]), .Z(n3696) );
  XNOR U5750 ( .A(y[1619]), .B(x[1619]), .Z(n3695) );
  XNOR U5751 ( .A(n3686), .B(n3685), .Z(n3689) );
  XNOR U5752 ( .A(n3681), .B(n3682), .Z(n3685) );
  XNOR U5753 ( .A(y[1614]), .B(x[1614]), .Z(n3682) );
  XNOR U5754 ( .A(n3683), .B(n3684), .Z(n3681) );
  XNOR U5755 ( .A(y[1615]), .B(x[1615]), .Z(n3684) );
  XNOR U5756 ( .A(y[1616]), .B(x[1616]), .Z(n3683) );
  XNOR U5757 ( .A(n3675), .B(n3676), .Z(n3686) );
  XNOR U5758 ( .A(y[1611]), .B(x[1611]), .Z(n3676) );
  XNOR U5759 ( .A(n3677), .B(n3678), .Z(n3675) );
  XNOR U5760 ( .A(y[1612]), .B(x[1612]), .Z(n3678) );
  XNOR U5761 ( .A(y[1613]), .B(x[1613]), .Z(n3677) );
  XOR U5762 ( .A(n3651), .B(n3652), .Z(n3670) );
  XNOR U5763 ( .A(n3667), .B(n3668), .Z(n3652) );
  XNOR U5764 ( .A(n3662), .B(n3663), .Z(n3668) );
  XNOR U5765 ( .A(n3664), .B(n3665), .Z(n3663) );
  XNOR U5766 ( .A(y[1609]), .B(x[1609]), .Z(n3665) );
  XNOR U5767 ( .A(y[1610]), .B(x[1610]), .Z(n3664) );
  XNOR U5768 ( .A(y[1608]), .B(x[1608]), .Z(n3662) );
  XNOR U5769 ( .A(n3656), .B(n3657), .Z(n3667) );
  XNOR U5770 ( .A(y[1605]), .B(x[1605]), .Z(n3657) );
  XNOR U5771 ( .A(n3658), .B(n3659), .Z(n3656) );
  XNOR U5772 ( .A(y[1606]), .B(x[1606]), .Z(n3659) );
  XNOR U5773 ( .A(y[1607]), .B(x[1607]), .Z(n3658) );
  XOR U5774 ( .A(n3650), .B(n3649), .Z(n3651) );
  XNOR U5775 ( .A(n3645), .B(n3646), .Z(n3649) );
  XNOR U5776 ( .A(y[1602]), .B(x[1602]), .Z(n3646) );
  XNOR U5777 ( .A(n3647), .B(n3648), .Z(n3645) );
  XNOR U5778 ( .A(y[1603]), .B(x[1603]), .Z(n3648) );
  XNOR U5779 ( .A(y[1604]), .B(x[1604]), .Z(n3647) );
  XNOR U5780 ( .A(n3639), .B(n3640), .Z(n3650) );
  XNOR U5781 ( .A(y[1599]), .B(x[1599]), .Z(n3640) );
  XNOR U5782 ( .A(n3641), .B(n3642), .Z(n3639) );
  XNOR U5783 ( .A(y[1600]), .B(x[1600]), .Z(n3642) );
  XNOR U5784 ( .A(y[1601]), .B(x[1601]), .Z(n3641) );
  NAND U5785 ( .A(n3706), .B(n3707), .Z(N13511) );
  NANDN U5786 ( .A(n3708), .B(n3709), .Z(n3707) );
  OR U5787 ( .A(n3710), .B(n3711), .Z(n3709) );
  NAND U5788 ( .A(n3710), .B(n3711), .Z(n3706) );
  XOR U5789 ( .A(n3710), .B(n3712), .Z(N13510) );
  XNOR U5790 ( .A(n3708), .B(n3711), .Z(n3712) );
  AND U5791 ( .A(n3713), .B(n3714), .Z(n3711) );
  NANDN U5792 ( .A(n3715), .B(n3716), .Z(n3714) );
  NANDN U5793 ( .A(n3717), .B(n3718), .Z(n3716) );
  NANDN U5794 ( .A(n3718), .B(n3717), .Z(n3713) );
  NAND U5795 ( .A(n3719), .B(n3720), .Z(n3708) );
  NANDN U5796 ( .A(n3721), .B(n3722), .Z(n3720) );
  OR U5797 ( .A(n3723), .B(n3724), .Z(n3722) );
  NAND U5798 ( .A(n3724), .B(n3723), .Z(n3719) );
  AND U5799 ( .A(n3725), .B(n3726), .Z(n3710) );
  NANDN U5800 ( .A(n3727), .B(n3728), .Z(n3726) );
  NANDN U5801 ( .A(n3729), .B(n3730), .Z(n3728) );
  NANDN U5802 ( .A(n3730), .B(n3729), .Z(n3725) );
  XOR U5803 ( .A(n3724), .B(n3731), .Z(N13509) );
  XOR U5804 ( .A(n3721), .B(n3723), .Z(n3731) );
  XNOR U5805 ( .A(n3717), .B(n3732), .Z(n3723) );
  XNOR U5806 ( .A(n3715), .B(n3718), .Z(n3732) );
  NAND U5807 ( .A(n3733), .B(n3734), .Z(n3718) );
  NAND U5808 ( .A(n3735), .B(n3736), .Z(n3734) );
  OR U5809 ( .A(n3737), .B(n3738), .Z(n3735) );
  NANDN U5810 ( .A(n3739), .B(n3737), .Z(n3733) );
  IV U5811 ( .A(n3738), .Z(n3739) );
  NAND U5812 ( .A(n3740), .B(n3741), .Z(n3715) );
  NAND U5813 ( .A(n3742), .B(n3743), .Z(n3741) );
  NANDN U5814 ( .A(n3744), .B(n3745), .Z(n3742) );
  NANDN U5815 ( .A(n3745), .B(n3744), .Z(n3740) );
  AND U5816 ( .A(n3746), .B(n3747), .Z(n3717) );
  NAND U5817 ( .A(n3748), .B(n3749), .Z(n3747) );
  OR U5818 ( .A(n3750), .B(n3751), .Z(n3748) );
  NANDN U5819 ( .A(n3752), .B(n3750), .Z(n3746) );
  NAND U5820 ( .A(n3753), .B(n3754), .Z(n3721) );
  NANDN U5821 ( .A(n3755), .B(n3756), .Z(n3754) );
  OR U5822 ( .A(n3757), .B(n3758), .Z(n3756) );
  NANDN U5823 ( .A(n3759), .B(n3757), .Z(n3753) );
  IV U5824 ( .A(n3758), .Z(n3759) );
  XNOR U5825 ( .A(n3729), .B(n3760), .Z(n3724) );
  XNOR U5826 ( .A(n3727), .B(n3730), .Z(n3760) );
  NAND U5827 ( .A(n3761), .B(n3762), .Z(n3730) );
  NAND U5828 ( .A(n3763), .B(n3764), .Z(n3762) );
  OR U5829 ( .A(n3765), .B(n3766), .Z(n3763) );
  NANDN U5830 ( .A(n3767), .B(n3765), .Z(n3761) );
  IV U5831 ( .A(n3766), .Z(n3767) );
  NAND U5832 ( .A(n3768), .B(n3769), .Z(n3727) );
  NAND U5833 ( .A(n3770), .B(n3771), .Z(n3769) );
  NANDN U5834 ( .A(n3772), .B(n3773), .Z(n3770) );
  NANDN U5835 ( .A(n3773), .B(n3772), .Z(n3768) );
  AND U5836 ( .A(n3774), .B(n3775), .Z(n3729) );
  NAND U5837 ( .A(n3776), .B(n3777), .Z(n3775) );
  OR U5838 ( .A(n3778), .B(n3779), .Z(n3776) );
  NANDN U5839 ( .A(n3780), .B(n3778), .Z(n3774) );
  XNOR U5840 ( .A(n3755), .B(n3781), .Z(N13508) );
  XOR U5841 ( .A(n3757), .B(n3758), .Z(n3781) );
  XNOR U5842 ( .A(n3771), .B(n3782), .Z(n3758) );
  XOR U5843 ( .A(n3772), .B(n3773), .Z(n3782) );
  XOR U5844 ( .A(n3778), .B(n3783), .Z(n3773) );
  XOR U5845 ( .A(n3777), .B(n3780), .Z(n3783) );
  IV U5846 ( .A(n3779), .Z(n3780) );
  NAND U5847 ( .A(n3784), .B(n3785), .Z(n3779) );
  OR U5848 ( .A(n3786), .B(n3787), .Z(n3785) );
  OR U5849 ( .A(n3788), .B(n3789), .Z(n3784) );
  NAND U5850 ( .A(n3790), .B(n3791), .Z(n3777) );
  OR U5851 ( .A(n3792), .B(n3793), .Z(n3791) );
  OR U5852 ( .A(n3794), .B(n3795), .Z(n3790) );
  NOR U5853 ( .A(n3796), .B(n3797), .Z(n3778) );
  ANDN U5854 ( .B(n3798), .A(n3799), .Z(n3772) );
  XNOR U5855 ( .A(n3765), .B(n3800), .Z(n3771) );
  XNOR U5856 ( .A(n3764), .B(n3766), .Z(n3800) );
  NAND U5857 ( .A(n3801), .B(n3802), .Z(n3766) );
  OR U5858 ( .A(n3803), .B(n3804), .Z(n3802) );
  OR U5859 ( .A(n3805), .B(n3806), .Z(n3801) );
  NAND U5860 ( .A(n3807), .B(n3808), .Z(n3764) );
  OR U5861 ( .A(n3809), .B(n3810), .Z(n3808) );
  OR U5862 ( .A(n3811), .B(n3812), .Z(n3807) );
  ANDN U5863 ( .B(n3813), .A(n3814), .Z(n3765) );
  IV U5864 ( .A(n3815), .Z(n3813) );
  ANDN U5865 ( .B(n3816), .A(n3817), .Z(n3757) );
  XOR U5866 ( .A(n3743), .B(n3818), .Z(n3755) );
  XOR U5867 ( .A(n3744), .B(n3745), .Z(n3818) );
  XOR U5868 ( .A(n3750), .B(n3819), .Z(n3745) );
  XOR U5869 ( .A(n3749), .B(n3752), .Z(n3819) );
  IV U5870 ( .A(n3751), .Z(n3752) );
  NAND U5871 ( .A(n3820), .B(n3821), .Z(n3751) );
  OR U5872 ( .A(n3822), .B(n3823), .Z(n3821) );
  OR U5873 ( .A(n3824), .B(n3825), .Z(n3820) );
  NAND U5874 ( .A(n3826), .B(n3827), .Z(n3749) );
  OR U5875 ( .A(n3828), .B(n3829), .Z(n3827) );
  OR U5876 ( .A(n3830), .B(n3831), .Z(n3826) );
  NOR U5877 ( .A(n3832), .B(n3833), .Z(n3750) );
  ANDN U5878 ( .B(n3834), .A(n3835), .Z(n3744) );
  IV U5879 ( .A(n3836), .Z(n3834) );
  XNOR U5880 ( .A(n3737), .B(n3837), .Z(n3743) );
  XNOR U5881 ( .A(n3736), .B(n3738), .Z(n3837) );
  NAND U5882 ( .A(n3838), .B(n3839), .Z(n3738) );
  OR U5883 ( .A(n3840), .B(n3841), .Z(n3839) );
  OR U5884 ( .A(n3842), .B(n3843), .Z(n3838) );
  NAND U5885 ( .A(n3844), .B(n3845), .Z(n3736) );
  OR U5886 ( .A(n3846), .B(n3847), .Z(n3845) );
  OR U5887 ( .A(n3848), .B(n3849), .Z(n3844) );
  ANDN U5888 ( .B(n3850), .A(n3851), .Z(n3737) );
  IV U5889 ( .A(n3852), .Z(n3850) );
  XNOR U5890 ( .A(n3817), .B(n3816), .Z(N13507) );
  XOR U5891 ( .A(n3836), .B(n3835), .Z(n3816) );
  XNOR U5892 ( .A(n3851), .B(n3852), .Z(n3835) );
  XNOR U5893 ( .A(n3846), .B(n3847), .Z(n3852) );
  XNOR U5894 ( .A(n3848), .B(n3849), .Z(n3847) );
  XNOR U5895 ( .A(y[1597]), .B(x[1597]), .Z(n3849) );
  XNOR U5896 ( .A(y[1598]), .B(x[1598]), .Z(n3848) );
  XNOR U5897 ( .A(y[1596]), .B(x[1596]), .Z(n3846) );
  XNOR U5898 ( .A(n3840), .B(n3841), .Z(n3851) );
  XNOR U5899 ( .A(y[1593]), .B(x[1593]), .Z(n3841) );
  XNOR U5900 ( .A(n3842), .B(n3843), .Z(n3840) );
  XNOR U5901 ( .A(y[1594]), .B(x[1594]), .Z(n3843) );
  XNOR U5902 ( .A(y[1595]), .B(x[1595]), .Z(n3842) );
  XNOR U5903 ( .A(n3833), .B(n3832), .Z(n3836) );
  XNOR U5904 ( .A(n3828), .B(n3829), .Z(n3832) );
  XNOR U5905 ( .A(y[1590]), .B(x[1590]), .Z(n3829) );
  XNOR U5906 ( .A(n3830), .B(n3831), .Z(n3828) );
  XNOR U5907 ( .A(y[1591]), .B(x[1591]), .Z(n3831) );
  XNOR U5908 ( .A(y[1592]), .B(x[1592]), .Z(n3830) );
  XNOR U5909 ( .A(n3822), .B(n3823), .Z(n3833) );
  XNOR U5910 ( .A(y[1587]), .B(x[1587]), .Z(n3823) );
  XNOR U5911 ( .A(n3824), .B(n3825), .Z(n3822) );
  XNOR U5912 ( .A(y[1588]), .B(x[1588]), .Z(n3825) );
  XNOR U5913 ( .A(y[1589]), .B(x[1589]), .Z(n3824) );
  XOR U5914 ( .A(n3798), .B(n3799), .Z(n3817) );
  XNOR U5915 ( .A(n3814), .B(n3815), .Z(n3799) );
  XNOR U5916 ( .A(n3809), .B(n3810), .Z(n3815) );
  XNOR U5917 ( .A(n3811), .B(n3812), .Z(n3810) );
  XNOR U5918 ( .A(y[1585]), .B(x[1585]), .Z(n3812) );
  XNOR U5919 ( .A(y[1586]), .B(x[1586]), .Z(n3811) );
  XNOR U5920 ( .A(y[1584]), .B(x[1584]), .Z(n3809) );
  XNOR U5921 ( .A(n3803), .B(n3804), .Z(n3814) );
  XNOR U5922 ( .A(y[1581]), .B(x[1581]), .Z(n3804) );
  XNOR U5923 ( .A(n3805), .B(n3806), .Z(n3803) );
  XNOR U5924 ( .A(y[1582]), .B(x[1582]), .Z(n3806) );
  XNOR U5925 ( .A(y[1583]), .B(x[1583]), .Z(n3805) );
  XOR U5926 ( .A(n3797), .B(n3796), .Z(n3798) );
  XNOR U5927 ( .A(n3792), .B(n3793), .Z(n3796) );
  XNOR U5928 ( .A(y[1578]), .B(x[1578]), .Z(n3793) );
  XNOR U5929 ( .A(n3794), .B(n3795), .Z(n3792) );
  XNOR U5930 ( .A(y[1579]), .B(x[1579]), .Z(n3795) );
  XNOR U5931 ( .A(y[1580]), .B(x[1580]), .Z(n3794) );
  XNOR U5932 ( .A(n3786), .B(n3787), .Z(n3797) );
  XNOR U5933 ( .A(y[1575]), .B(x[1575]), .Z(n3787) );
  XNOR U5934 ( .A(n3788), .B(n3789), .Z(n3786) );
  XNOR U5935 ( .A(y[1576]), .B(x[1576]), .Z(n3789) );
  XNOR U5936 ( .A(y[1577]), .B(x[1577]), .Z(n3788) );
  NAND U5937 ( .A(n3853), .B(n3854), .Z(N13500) );
  NANDN U5938 ( .A(n3855), .B(n3856), .Z(n3854) );
  OR U5939 ( .A(n3857), .B(n3858), .Z(n3856) );
  NAND U5940 ( .A(n3857), .B(n3858), .Z(n3853) );
  XOR U5941 ( .A(n3857), .B(n3859), .Z(N13499) );
  XNOR U5942 ( .A(n3855), .B(n3858), .Z(n3859) );
  AND U5943 ( .A(n3860), .B(n3861), .Z(n3858) );
  NANDN U5944 ( .A(n3862), .B(n3863), .Z(n3861) );
  NANDN U5945 ( .A(n3864), .B(n3865), .Z(n3863) );
  NANDN U5946 ( .A(n3865), .B(n3864), .Z(n3860) );
  NAND U5947 ( .A(n3866), .B(n3867), .Z(n3855) );
  NANDN U5948 ( .A(n3868), .B(n3869), .Z(n3867) );
  OR U5949 ( .A(n3870), .B(n3871), .Z(n3869) );
  NAND U5950 ( .A(n3871), .B(n3870), .Z(n3866) );
  AND U5951 ( .A(n3872), .B(n3873), .Z(n3857) );
  NANDN U5952 ( .A(n3874), .B(n3875), .Z(n3873) );
  NANDN U5953 ( .A(n3876), .B(n3877), .Z(n3875) );
  NANDN U5954 ( .A(n3877), .B(n3876), .Z(n3872) );
  XOR U5955 ( .A(n3871), .B(n3878), .Z(N13498) );
  XOR U5956 ( .A(n3868), .B(n3870), .Z(n3878) );
  XNOR U5957 ( .A(n3864), .B(n3879), .Z(n3870) );
  XNOR U5958 ( .A(n3862), .B(n3865), .Z(n3879) );
  NAND U5959 ( .A(n3880), .B(n3881), .Z(n3865) );
  NAND U5960 ( .A(n3882), .B(n3883), .Z(n3881) );
  OR U5961 ( .A(n3884), .B(n3885), .Z(n3882) );
  NANDN U5962 ( .A(n3886), .B(n3884), .Z(n3880) );
  IV U5963 ( .A(n3885), .Z(n3886) );
  NAND U5964 ( .A(n3887), .B(n3888), .Z(n3862) );
  NAND U5965 ( .A(n3889), .B(n3890), .Z(n3888) );
  NANDN U5966 ( .A(n3891), .B(n3892), .Z(n3889) );
  NANDN U5967 ( .A(n3892), .B(n3891), .Z(n3887) );
  AND U5968 ( .A(n3893), .B(n3894), .Z(n3864) );
  NAND U5969 ( .A(n3895), .B(n3896), .Z(n3894) );
  OR U5970 ( .A(n3897), .B(n3898), .Z(n3895) );
  NANDN U5971 ( .A(n3899), .B(n3897), .Z(n3893) );
  NAND U5972 ( .A(n3900), .B(n3901), .Z(n3868) );
  NANDN U5973 ( .A(n3902), .B(n3903), .Z(n3901) );
  OR U5974 ( .A(n3904), .B(n3905), .Z(n3903) );
  NANDN U5975 ( .A(n3906), .B(n3904), .Z(n3900) );
  IV U5976 ( .A(n3905), .Z(n3906) );
  XNOR U5977 ( .A(n3876), .B(n3907), .Z(n3871) );
  XNOR U5978 ( .A(n3874), .B(n3877), .Z(n3907) );
  NAND U5979 ( .A(n3908), .B(n3909), .Z(n3877) );
  NAND U5980 ( .A(n3910), .B(n3911), .Z(n3909) );
  OR U5981 ( .A(n3912), .B(n3913), .Z(n3910) );
  NANDN U5982 ( .A(n3914), .B(n3912), .Z(n3908) );
  IV U5983 ( .A(n3913), .Z(n3914) );
  NAND U5984 ( .A(n3915), .B(n3916), .Z(n3874) );
  NAND U5985 ( .A(n3917), .B(n3918), .Z(n3916) );
  NANDN U5986 ( .A(n3919), .B(n3920), .Z(n3917) );
  NANDN U5987 ( .A(n3920), .B(n3919), .Z(n3915) );
  AND U5988 ( .A(n3921), .B(n3922), .Z(n3876) );
  NAND U5989 ( .A(n3923), .B(n3924), .Z(n3922) );
  OR U5990 ( .A(n3925), .B(n3926), .Z(n3923) );
  NANDN U5991 ( .A(n3927), .B(n3925), .Z(n3921) );
  XNOR U5992 ( .A(n3902), .B(n3928), .Z(N13497) );
  XOR U5993 ( .A(n3904), .B(n3905), .Z(n3928) );
  XNOR U5994 ( .A(n3918), .B(n3929), .Z(n3905) );
  XOR U5995 ( .A(n3919), .B(n3920), .Z(n3929) );
  XOR U5996 ( .A(n3925), .B(n3930), .Z(n3920) );
  XOR U5997 ( .A(n3924), .B(n3927), .Z(n3930) );
  IV U5998 ( .A(n3926), .Z(n3927) );
  NAND U5999 ( .A(n3931), .B(n3932), .Z(n3926) );
  OR U6000 ( .A(n3933), .B(n3934), .Z(n3932) );
  OR U6001 ( .A(n3935), .B(n3936), .Z(n3931) );
  NAND U6002 ( .A(n3937), .B(n3938), .Z(n3924) );
  OR U6003 ( .A(n3939), .B(n3940), .Z(n3938) );
  OR U6004 ( .A(n3941), .B(n3942), .Z(n3937) );
  NOR U6005 ( .A(n3943), .B(n3944), .Z(n3925) );
  ANDN U6006 ( .B(n3945), .A(n3946), .Z(n3919) );
  XNOR U6007 ( .A(n3912), .B(n3947), .Z(n3918) );
  XNOR U6008 ( .A(n3911), .B(n3913), .Z(n3947) );
  NAND U6009 ( .A(n3948), .B(n3949), .Z(n3913) );
  OR U6010 ( .A(n3950), .B(n3951), .Z(n3949) );
  OR U6011 ( .A(n3952), .B(n3953), .Z(n3948) );
  NAND U6012 ( .A(n3954), .B(n3955), .Z(n3911) );
  OR U6013 ( .A(n3956), .B(n3957), .Z(n3955) );
  OR U6014 ( .A(n3958), .B(n3959), .Z(n3954) );
  ANDN U6015 ( .B(n3960), .A(n3961), .Z(n3912) );
  IV U6016 ( .A(n3962), .Z(n3960) );
  ANDN U6017 ( .B(n3963), .A(n3964), .Z(n3904) );
  XOR U6018 ( .A(n3890), .B(n3965), .Z(n3902) );
  XOR U6019 ( .A(n3891), .B(n3892), .Z(n3965) );
  XOR U6020 ( .A(n3897), .B(n3966), .Z(n3892) );
  XOR U6021 ( .A(n3896), .B(n3899), .Z(n3966) );
  IV U6022 ( .A(n3898), .Z(n3899) );
  NAND U6023 ( .A(n3967), .B(n3968), .Z(n3898) );
  OR U6024 ( .A(n3969), .B(n3970), .Z(n3968) );
  OR U6025 ( .A(n3971), .B(n3972), .Z(n3967) );
  NAND U6026 ( .A(n3973), .B(n3974), .Z(n3896) );
  OR U6027 ( .A(n3975), .B(n3976), .Z(n3974) );
  OR U6028 ( .A(n3977), .B(n3978), .Z(n3973) );
  NOR U6029 ( .A(n3979), .B(n3980), .Z(n3897) );
  ANDN U6030 ( .B(n3981), .A(n3982), .Z(n3891) );
  IV U6031 ( .A(n3983), .Z(n3981) );
  XNOR U6032 ( .A(n3884), .B(n3984), .Z(n3890) );
  XNOR U6033 ( .A(n3883), .B(n3885), .Z(n3984) );
  NAND U6034 ( .A(n3985), .B(n3986), .Z(n3885) );
  OR U6035 ( .A(n3987), .B(n3988), .Z(n3986) );
  OR U6036 ( .A(n3989), .B(n3990), .Z(n3985) );
  NAND U6037 ( .A(n3991), .B(n3992), .Z(n3883) );
  OR U6038 ( .A(n3993), .B(n3994), .Z(n3992) );
  OR U6039 ( .A(n3995), .B(n3996), .Z(n3991) );
  ANDN U6040 ( .B(n3997), .A(n3998), .Z(n3884) );
  IV U6041 ( .A(n3999), .Z(n3997) );
  XNOR U6042 ( .A(n3964), .B(n3963), .Z(N13496) );
  XOR U6043 ( .A(n3983), .B(n3982), .Z(n3963) );
  XNOR U6044 ( .A(n3998), .B(n3999), .Z(n3982) );
  XNOR U6045 ( .A(n3993), .B(n3994), .Z(n3999) );
  XNOR U6046 ( .A(n3995), .B(n3996), .Z(n3994) );
  XNOR U6047 ( .A(y[1573]), .B(x[1573]), .Z(n3996) );
  XNOR U6048 ( .A(y[1574]), .B(x[1574]), .Z(n3995) );
  XNOR U6049 ( .A(y[1572]), .B(x[1572]), .Z(n3993) );
  XNOR U6050 ( .A(n3987), .B(n3988), .Z(n3998) );
  XNOR U6051 ( .A(y[1569]), .B(x[1569]), .Z(n3988) );
  XNOR U6052 ( .A(n3989), .B(n3990), .Z(n3987) );
  XNOR U6053 ( .A(y[1570]), .B(x[1570]), .Z(n3990) );
  XNOR U6054 ( .A(y[1571]), .B(x[1571]), .Z(n3989) );
  XNOR U6055 ( .A(n3980), .B(n3979), .Z(n3983) );
  XNOR U6056 ( .A(n3975), .B(n3976), .Z(n3979) );
  XNOR U6057 ( .A(y[1566]), .B(x[1566]), .Z(n3976) );
  XNOR U6058 ( .A(n3977), .B(n3978), .Z(n3975) );
  XNOR U6059 ( .A(y[1567]), .B(x[1567]), .Z(n3978) );
  XNOR U6060 ( .A(y[1568]), .B(x[1568]), .Z(n3977) );
  XNOR U6061 ( .A(n3969), .B(n3970), .Z(n3980) );
  XNOR U6062 ( .A(y[1563]), .B(x[1563]), .Z(n3970) );
  XNOR U6063 ( .A(n3971), .B(n3972), .Z(n3969) );
  XNOR U6064 ( .A(y[1564]), .B(x[1564]), .Z(n3972) );
  XNOR U6065 ( .A(y[1565]), .B(x[1565]), .Z(n3971) );
  XOR U6066 ( .A(n3945), .B(n3946), .Z(n3964) );
  XNOR U6067 ( .A(n3961), .B(n3962), .Z(n3946) );
  XNOR U6068 ( .A(n3956), .B(n3957), .Z(n3962) );
  XNOR U6069 ( .A(n3958), .B(n3959), .Z(n3957) );
  XNOR U6070 ( .A(y[1561]), .B(x[1561]), .Z(n3959) );
  XNOR U6071 ( .A(y[1562]), .B(x[1562]), .Z(n3958) );
  XNOR U6072 ( .A(y[1560]), .B(x[1560]), .Z(n3956) );
  XNOR U6073 ( .A(n3950), .B(n3951), .Z(n3961) );
  XNOR U6074 ( .A(y[1557]), .B(x[1557]), .Z(n3951) );
  XNOR U6075 ( .A(n3952), .B(n3953), .Z(n3950) );
  XNOR U6076 ( .A(y[1558]), .B(x[1558]), .Z(n3953) );
  XNOR U6077 ( .A(y[1559]), .B(x[1559]), .Z(n3952) );
  XOR U6078 ( .A(n3944), .B(n3943), .Z(n3945) );
  XNOR U6079 ( .A(n3939), .B(n3940), .Z(n3943) );
  XNOR U6080 ( .A(y[1554]), .B(x[1554]), .Z(n3940) );
  XNOR U6081 ( .A(n3941), .B(n3942), .Z(n3939) );
  XNOR U6082 ( .A(y[1555]), .B(x[1555]), .Z(n3942) );
  XNOR U6083 ( .A(y[1556]), .B(x[1556]), .Z(n3941) );
  XNOR U6084 ( .A(n3933), .B(n3934), .Z(n3944) );
  XNOR U6085 ( .A(y[1551]), .B(x[1551]), .Z(n3934) );
  XNOR U6086 ( .A(n3935), .B(n3936), .Z(n3933) );
  XNOR U6087 ( .A(y[1552]), .B(x[1552]), .Z(n3936) );
  XNOR U6088 ( .A(y[1553]), .B(x[1553]), .Z(n3935) );
  NAND U6089 ( .A(n4000), .B(n4001), .Z(N13489) );
  NANDN U6090 ( .A(n4002), .B(n4003), .Z(n4001) );
  OR U6091 ( .A(n4004), .B(n4005), .Z(n4003) );
  NAND U6092 ( .A(n4004), .B(n4005), .Z(n4000) );
  XOR U6093 ( .A(n4004), .B(n4006), .Z(N13488) );
  XNOR U6094 ( .A(n4002), .B(n4005), .Z(n4006) );
  AND U6095 ( .A(n4007), .B(n4008), .Z(n4005) );
  NANDN U6096 ( .A(n4009), .B(n4010), .Z(n4008) );
  NANDN U6097 ( .A(n4011), .B(n4012), .Z(n4010) );
  NANDN U6098 ( .A(n4012), .B(n4011), .Z(n4007) );
  NAND U6099 ( .A(n4013), .B(n4014), .Z(n4002) );
  NANDN U6100 ( .A(n4015), .B(n4016), .Z(n4014) );
  OR U6101 ( .A(n4017), .B(n4018), .Z(n4016) );
  NAND U6102 ( .A(n4018), .B(n4017), .Z(n4013) );
  AND U6103 ( .A(n4019), .B(n4020), .Z(n4004) );
  NANDN U6104 ( .A(n4021), .B(n4022), .Z(n4020) );
  NANDN U6105 ( .A(n4023), .B(n4024), .Z(n4022) );
  NANDN U6106 ( .A(n4024), .B(n4023), .Z(n4019) );
  XOR U6107 ( .A(n4018), .B(n4025), .Z(N13487) );
  XOR U6108 ( .A(n4015), .B(n4017), .Z(n4025) );
  XNOR U6109 ( .A(n4011), .B(n4026), .Z(n4017) );
  XNOR U6110 ( .A(n4009), .B(n4012), .Z(n4026) );
  NAND U6111 ( .A(n4027), .B(n4028), .Z(n4012) );
  NAND U6112 ( .A(n4029), .B(n4030), .Z(n4028) );
  OR U6113 ( .A(n4031), .B(n4032), .Z(n4029) );
  NANDN U6114 ( .A(n4033), .B(n4031), .Z(n4027) );
  IV U6115 ( .A(n4032), .Z(n4033) );
  NAND U6116 ( .A(n4034), .B(n4035), .Z(n4009) );
  NAND U6117 ( .A(n4036), .B(n4037), .Z(n4035) );
  NANDN U6118 ( .A(n4038), .B(n4039), .Z(n4036) );
  NANDN U6119 ( .A(n4039), .B(n4038), .Z(n4034) );
  AND U6120 ( .A(n4040), .B(n4041), .Z(n4011) );
  NAND U6121 ( .A(n4042), .B(n4043), .Z(n4041) );
  OR U6122 ( .A(n4044), .B(n4045), .Z(n4042) );
  NANDN U6123 ( .A(n4046), .B(n4044), .Z(n4040) );
  NAND U6124 ( .A(n4047), .B(n4048), .Z(n4015) );
  NANDN U6125 ( .A(n4049), .B(n4050), .Z(n4048) );
  OR U6126 ( .A(n4051), .B(n4052), .Z(n4050) );
  NANDN U6127 ( .A(n4053), .B(n4051), .Z(n4047) );
  IV U6128 ( .A(n4052), .Z(n4053) );
  XNOR U6129 ( .A(n4023), .B(n4054), .Z(n4018) );
  XNOR U6130 ( .A(n4021), .B(n4024), .Z(n4054) );
  NAND U6131 ( .A(n4055), .B(n4056), .Z(n4024) );
  NAND U6132 ( .A(n4057), .B(n4058), .Z(n4056) );
  OR U6133 ( .A(n4059), .B(n4060), .Z(n4057) );
  NANDN U6134 ( .A(n4061), .B(n4059), .Z(n4055) );
  IV U6135 ( .A(n4060), .Z(n4061) );
  NAND U6136 ( .A(n4062), .B(n4063), .Z(n4021) );
  NAND U6137 ( .A(n4064), .B(n4065), .Z(n4063) );
  NANDN U6138 ( .A(n4066), .B(n4067), .Z(n4064) );
  NANDN U6139 ( .A(n4067), .B(n4066), .Z(n4062) );
  AND U6140 ( .A(n4068), .B(n4069), .Z(n4023) );
  NAND U6141 ( .A(n4070), .B(n4071), .Z(n4069) );
  OR U6142 ( .A(n4072), .B(n4073), .Z(n4070) );
  NANDN U6143 ( .A(n4074), .B(n4072), .Z(n4068) );
  XNOR U6144 ( .A(n4049), .B(n4075), .Z(N13486) );
  XOR U6145 ( .A(n4051), .B(n4052), .Z(n4075) );
  XNOR U6146 ( .A(n4065), .B(n4076), .Z(n4052) );
  XOR U6147 ( .A(n4066), .B(n4067), .Z(n4076) );
  XOR U6148 ( .A(n4072), .B(n4077), .Z(n4067) );
  XOR U6149 ( .A(n4071), .B(n4074), .Z(n4077) );
  IV U6150 ( .A(n4073), .Z(n4074) );
  NAND U6151 ( .A(n4078), .B(n4079), .Z(n4073) );
  OR U6152 ( .A(n4080), .B(n4081), .Z(n4079) );
  OR U6153 ( .A(n4082), .B(n4083), .Z(n4078) );
  NAND U6154 ( .A(n4084), .B(n4085), .Z(n4071) );
  OR U6155 ( .A(n4086), .B(n4087), .Z(n4085) );
  OR U6156 ( .A(n4088), .B(n4089), .Z(n4084) );
  NOR U6157 ( .A(n4090), .B(n4091), .Z(n4072) );
  ANDN U6158 ( .B(n4092), .A(n4093), .Z(n4066) );
  XNOR U6159 ( .A(n4059), .B(n4094), .Z(n4065) );
  XNOR U6160 ( .A(n4058), .B(n4060), .Z(n4094) );
  NAND U6161 ( .A(n4095), .B(n4096), .Z(n4060) );
  OR U6162 ( .A(n4097), .B(n4098), .Z(n4096) );
  OR U6163 ( .A(n4099), .B(n4100), .Z(n4095) );
  NAND U6164 ( .A(n4101), .B(n4102), .Z(n4058) );
  OR U6165 ( .A(n4103), .B(n4104), .Z(n4102) );
  OR U6166 ( .A(n4105), .B(n4106), .Z(n4101) );
  ANDN U6167 ( .B(n4107), .A(n4108), .Z(n4059) );
  IV U6168 ( .A(n4109), .Z(n4107) );
  ANDN U6169 ( .B(n4110), .A(n4111), .Z(n4051) );
  XOR U6170 ( .A(n4037), .B(n4112), .Z(n4049) );
  XOR U6171 ( .A(n4038), .B(n4039), .Z(n4112) );
  XOR U6172 ( .A(n4044), .B(n4113), .Z(n4039) );
  XOR U6173 ( .A(n4043), .B(n4046), .Z(n4113) );
  IV U6174 ( .A(n4045), .Z(n4046) );
  NAND U6175 ( .A(n4114), .B(n4115), .Z(n4045) );
  OR U6176 ( .A(n4116), .B(n4117), .Z(n4115) );
  OR U6177 ( .A(n4118), .B(n4119), .Z(n4114) );
  NAND U6178 ( .A(n4120), .B(n4121), .Z(n4043) );
  OR U6179 ( .A(n4122), .B(n4123), .Z(n4121) );
  OR U6180 ( .A(n4124), .B(n4125), .Z(n4120) );
  NOR U6181 ( .A(n4126), .B(n4127), .Z(n4044) );
  ANDN U6182 ( .B(n4128), .A(n4129), .Z(n4038) );
  IV U6183 ( .A(n4130), .Z(n4128) );
  XNOR U6184 ( .A(n4031), .B(n4131), .Z(n4037) );
  XNOR U6185 ( .A(n4030), .B(n4032), .Z(n4131) );
  NAND U6186 ( .A(n4132), .B(n4133), .Z(n4032) );
  OR U6187 ( .A(n4134), .B(n4135), .Z(n4133) );
  OR U6188 ( .A(n4136), .B(n4137), .Z(n4132) );
  NAND U6189 ( .A(n4138), .B(n4139), .Z(n4030) );
  OR U6190 ( .A(n4140), .B(n4141), .Z(n4139) );
  OR U6191 ( .A(n4142), .B(n4143), .Z(n4138) );
  ANDN U6192 ( .B(n4144), .A(n4145), .Z(n4031) );
  IV U6193 ( .A(n4146), .Z(n4144) );
  XNOR U6194 ( .A(n4111), .B(n4110), .Z(N13485) );
  XOR U6195 ( .A(n4130), .B(n4129), .Z(n4110) );
  XNOR U6196 ( .A(n4145), .B(n4146), .Z(n4129) );
  XNOR U6197 ( .A(n4140), .B(n4141), .Z(n4146) );
  XNOR U6198 ( .A(n4142), .B(n4143), .Z(n4141) );
  XNOR U6199 ( .A(y[1549]), .B(x[1549]), .Z(n4143) );
  XNOR U6200 ( .A(y[1550]), .B(x[1550]), .Z(n4142) );
  XNOR U6201 ( .A(y[1548]), .B(x[1548]), .Z(n4140) );
  XNOR U6202 ( .A(n4134), .B(n4135), .Z(n4145) );
  XNOR U6203 ( .A(y[1545]), .B(x[1545]), .Z(n4135) );
  XNOR U6204 ( .A(n4136), .B(n4137), .Z(n4134) );
  XNOR U6205 ( .A(y[1546]), .B(x[1546]), .Z(n4137) );
  XNOR U6206 ( .A(y[1547]), .B(x[1547]), .Z(n4136) );
  XNOR U6207 ( .A(n4127), .B(n4126), .Z(n4130) );
  XNOR U6208 ( .A(n4122), .B(n4123), .Z(n4126) );
  XNOR U6209 ( .A(y[1542]), .B(x[1542]), .Z(n4123) );
  XNOR U6210 ( .A(n4124), .B(n4125), .Z(n4122) );
  XNOR U6211 ( .A(y[1543]), .B(x[1543]), .Z(n4125) );
  XNOR U6212 ( .A(y[1544]), .B(x[1544]), .Z(n4124) );
  XNOR U6213 ( .A(n4116), .B(n4117), .Z(n4127) );
  XNOR U6214 ( .A(y[1539]), .B(x[1539]), .Z(n4117) );
  XNOR U6215 ( .A(n4118), .B(n4119), .Z(n4116) );
  XNOR U6216 ( .A(y[1540]), .B(x[1540]), .Z(n4119) );
  XNOR U6217 ( .A(y[1541]), .B(x[1541]), .Z(n4118) );
  XOR U6218 ( .A(n4092), .B(n4093), .Z(n4111) );
  XNOR U6219 ( .A(n4108), .B(n4109), .Z(n4093) );
  XNOR U6220 ( .A(n4103), .B(n4104), .Z(n4109) );
  XNOR U6221 ( .A(n4105), .B(n4106), .Z(n4104) );
  XNOR U6222 ( .A(y[1537]), .B(x[1537]), .Z(n4106) );
  XNOR U6223 ( .A(y[1538]), .B(x[1538]), .Z(n4105) );
  XNOR U6224 ( .A(y[1536]), .B(x[1536]), .Z(n4103) );
  XNOR U6225 ( .A(n4097), .B(n4098), .Z(n4108) );
  XNOR U6226 ( .A(y[1533]), .B(x[1533]), .Z(n4098) );
  XNOR U6227 ( .A(n4099), .B(n4100), .Z(n4097) );
  XNOR U6228 ( .A(y[1534]), .B(x[1534]), .Z(n4100) );
  XNOR U6229 ( .A(y[1535]), .B(x[1535]), .Z(n4099) );
  XOR U6230 ( .A(n4091), .B(n4090), .Z(n4092) );
  XNOR U6231 ( .A(n4086), .B(n4087), .Z(n4090) );
  XNOR U6232 ( .A(y[1530]), .B(x[1530]), .Z(n4087) );
  XNOR U6233 ( .A(n4088), .B(n4089), .Z(n4086) );
  XNOR U6234 ( .A(y[1531]), .B(x[1531]), .Z(n4089) );
  XNOR U6235 ( .A(y[1532]), .B(x[1532]), .Z(n4088) );
  XNOR U6236 ( .A(n4080), .B(n4081), .Z(n4091) );
  XNOR U6237 ( .A(y[1527]), .B(x[1527]), .Z(n4081) );
  XNOR U6238 ( .A(n4082), .B(n4083), .Z(n4080) );
  XNOR U6239 ( .A(y[1528]), .B(x[1528]), .Z(n4083) );
  XNOR U6240 ( .A(y[1529]), .B(x[1529]), .Z(n4082) );
  NAND U6241 ( .A(n4147), .B(n4148), .Z(N13478) );
  NANDN U6242 ( .A(n4149), .B(n4150), .Z(n4148) );
  OR U6243 ( .A(n4151), .B(n4152), .Z(n4150) );
  NAND U6244 ( .A(n4151), .B(n4152), .Z(n4147) );
  XOR U6245 ( .A(n4151), .B(n4153), .Z(N13477) );
  XNOR U6246 ( .A(n4149), .B(n4152), .Z(n4153) );
  AND U6247 ( .A(n4154), .B(n4155), .Z(n4152) );
  NANDN U6248 ( .A(n4156), .B(n4157), .Z(n4155) );
  NANDN U6249 ( .A(n4158), .B(n4159), .Z(n4157) );
  NANDN U6250 ( .A(n4159), .B(n4158), .Z(n4154) );
  NAND U6251 ( .A(n4160), .B(n4161), .Z(n4149) );
  NANDN U6252 ( .A(n4162), .B(n4163), .Z(n4161) );
  OR U6253 ( .A(n4164), .B(n4165), .Z(n4163) );
  NAND U6254 ( .A(n4165), .B(n4164), .Z(n4160) );
  AND U6255 ( .A(n4166), .B(n4167), .Z(n4151) );
  NANDN U6256 ( .A(n4168), .B(n4169), .Z(n4167) );
  NANDN U6257 ( .A(n4170), .B(n4171), .Z(n4169) );
  NANDN U6258 ( .A(n4171), .B(n4170), .Z(n4166) );
  XOR U6259 ( .A(n4165), .B(n4172), .Z(N13476) );
  XOR U6260 ( .A(n4162), .B(n4164), .Z(n4172) );
  XNOR U6261 ( .A(n4158), .B(n4173), .Z(n4164) );
  XNOR U6262 ( .A(n4156), .B(n4159), .Z(n4173) );
  NAND U6263 ( .A(n4174), .B(n4175), .Z(n4159) );
  NAND U6264 ( .A(n4176), .B(n4177), .Z(n4175) );
  OR U6265 ( .A(n4178), .B(n4179), .Z(n4176) );
  NANDN U6266 ( .A(n4180), .B(n4178), .Z(n4174) );
  IV U6267 ( .A(n4179), .Z(n4180) );
  NAND U6268 ( .A(n4181), .B(n4182), .Z(n4156) );
  NAND U6269 ( .A(n4183), .B(n4184), .Z(n4182) );
  NANDN U6270 ( .A(n4185), .B(n4186), .Z(n4183) );
  NANDN U6271 ( .A(n4186), .B(n4185), .Z(n4181) );
  AND U6272 ( .A(n4187), .B(n4188), .Z(n4158) );
  NAND U6273 ( .A(n4189), .B(n4190), .Z(n4188) );
  OR U6274 ( .A(n4191), .B(n4192), .Z(n4189) );
  NANDN U6275 ( .A(n4193), .B(n4191), .Z(n4187) );
  NAND U6276 ( .A(n4194), .B(n4195), .Z(n4162) );
  NANDN U6277 ( .A(n4196), .B(n4197), .Z(n4195) );
  OR U6278 ( .A(n4198), .B(n4199), .Z(n4197) );
  NANDN U6279 ( .A(n4200), .B(n4198), .Z(n4194) );
  IV U6280 ( .A(n4199), .Z(n4200) );
  XNOR U6281 ( .A(n4170), .B(n4201), .Z(n4165) );
  XNOR U6282 ( .A(n4168), .B(n4171), .Z(n4201) );
  NAND U6283 ( .A(n4202), .B(n4203), .Z(n4171) );
  NAND U6284 ( .A(n4204), .B(n4205), .Z(n4203) );
  OR U6285 ( .A(n4206), .B(n4207), .Z(n4204) );
  NANDN U6286 ( .A(n4208), .B(n4206), .Z(n4202) );
  IV U6287 ( .A(n4207), .Z(n4208) );
  NAND U6288 ( .A(n4209), .B(n4210), .Z(n4168) );
  NAND U6289 ( .A(n4211), .B(n4212), .Z(n4210) );
  NANDN U6290 ( .A(n4213), .B(n4214), .Z(n4211) );
  NANDN U6291 ( .A(n4214), .B(n4213), .Z(n4209) );
  AND U6292 ( .A(n4215), .B(n4216), .Z(n4170) );
  NAND U6293 ( .A(n4217), .B(n4218), .Z(n4216) );
  OR U6294 ( .A(n4219), .B(n4220), .Z(n4217) );
  NANDN U6295 ( .A(n4221), .B(n4219), .Z(n4215) );
  XNOR U6296 ( .A(n4196), .B(n4222), .Z(N13475) );
  XOR U6297 ( .A(n4198), .B(n4199), .Z(n4222) );
  XNOR U6298 ( .A(n4212), .B(n4223), .Z(n4199) );
  XOR U6299 ( .A(n4213), .B(n4214), .Z(n4223) );
  XOR U6300 ( .A(n4219), .B(n4224), .Z(n4214) );
  XOR U6301 ( .A(n4218), .B(n4221), .Z(n4224) );
  IV U6302 ( .A(n4220), .Z(n4221) );
  NAND U6303 ( .A(n4225), .B(n4226), .Z(n4220) );
  OR U6304 ( .A(n4227), .B(n4228), .Z(n4226) );
  OR U6305 ( .A(n4229), .B(n4230), .Z(n4225) );
  NAND U6306 ( .A(n4231), .B(n4232), .Z(n4218) );
  OR U6307 ( .A(n4233), .B(n4234), .Z(n4232) );
  OR U6308 ( .A(n4235), .B(n4236), .Z(n4231) );
  NOR U6309 ( .A(n4237), .B(n4238), .Z(n4219) );
  ANDN U6310 ( .B(n4239), .A(n4240), .Z(n4213) );
  XNOR U6311 ( .A(n4206), .B(n4241), .Z(n4212) );
  XNOR U6312 ( .A(n4205), .B(n4207), .Z(n4241) );
  NAND U6313 ( .A(n4242), .B(n4243), .Z(n4207) );
  OR U6314 ( .A(n4244), .B(n4245), .Z(n4243) );
  OR U6315 ( .A(n4246), .B(n4247), .Z(n4242) );
  NAND U6316 ( .A(n4248), .B(n4249), .Z(n4205) );
  OR U6317 ( .A(n4250), .B(n4251), .Z(n4249) );
  OR U6318 ( .A(n4252), .B(n4253), .Z(n4248) );
  ANDN U6319 ( .B(n4254), .A(n4255), .Z(n4206) );
  IV U6320 ( .A(n4256), .Z(n4254) );
  ANDN U6321 ( .B(n4257), .A(n4258), .Z(n4198) );
  XOR U6322 ( .A(n4184), .B(n4259), .Z(n4196) );
  XOR U6323 ( .A(n4185), .B(n4186), .Z(n4259) );
  XOR U6324 ( .A(n4191), .B(n4260), .Z(n4186) );
  XOR U6325 ( .A(n4190), .B(n4193), .Z(n4260) );
  IV U6326 ( .A(n4192), .Z(n4193) );
  NAND U6327 ( .A(n4261), .B(n4262), .Z(n4192) );
  OR U6328 ( .A(n4263), .B(n4264), .Z(n4262) );
  OR U6329 ( .A(n4265), .B(n4266), .Z(n4261) );
  NAND U6330 ( .A(n4267), .B(n4268), .Z(n4190) );
  OR U6331 ( .A(n4269), .B(n4270), .Z(n4268) );
  OR U6332 ( .A(n4271), .B(n4272), .Z(n4267) );
  NOR U6333 ( .A(n4273), .B(n4274), .Z(n4191) );
  ANDN U6334 ( .B(n4275), .A(n4276), .Z(n4185) );
  IV U6335 ( .A(n4277), .Z(n4275) );
  XNOR U6336 ( .A(n4178), .B(n4278), .Z(n4184) );
  XNOR U6337 ( .A(n4177), .B(n4179), .Z(n4278) );
  NAND U6338 ( .A(n4279), .B(n4280), .Z(n4179) );
  OR U6339 ( .A(n4281), .B(n4282), .Z(n4280) );
  OR U6340 ( .A(n4283), .B(n4284), .Z(n4279) );
  NAND U6341 ( .A(n4285), .B(n4286), .Z(n4177) );
  OR U6342 ( .A(n4287), .B(n4288), .Z(n4286) );
  OR U6343 ( .A(n4289), .B(n4290), .Z(n4285) );
  ANDN U6344 ( .B(n4291), .A(n4292), .Z(n4178) );
  IV U6345 ( .A(n4293), .Z(n4291) );
  XNOR U6346 ( .A(n4258), .B(n4257), .Z(N13474) );
  XOR U6347 ( .A(n4277), .B(n4276), .Z(n4257) );
  XNOR U6348 ( .A(n4292), .B(n4293), .Z(n4276) );
  XNOR U6349 ( .A(n4287), .B(n4288), .Z(n4293) );
  XNOR U6350 ( .A(n4289), .B(n4290), .Z(n4288) );
  XNOR U6351 ( .A(y[1525]), .B(x[1525]), .Z(n4290) );
  XNOR U6352 ( .A(y[1526]), .B(x[1526]), .Z(n4289) );
  XNOR U6353 ( .A(y[1524]), .B(x[1524]), .Z(n4287) );
  XNOR U6354 ( .A(n4281), .B(n4282), .Z(n4292) );
  XNOR U6355 ( .A(y[1521]), .B(x[1521]), .Z(n4282) );
  XNOR U6356 ( .A(n4283), .B(n4284), .Z(n4281) );
  XNOR U6357 ( .A(y[1522]), .B(x[1522]), .Z(n4284) );
  XNOR U6358 ( .A(y[1523]), .B(x[1523]), .Z(n4283) );
  XNOR U6359 ( .A(n4274), .B(n4273), .Z(n4277) );
  XNOR U6360 ( .A(n4269), .B(n4270), .Z(n4273) );
  XNOR U6361 ( .A(y[1518]), .B(x[1518]), .Z(n4270) );
  XNOR U6362 ( .A(n4271), .B(n4272), .Z(n4269) );
  XNOR U6363 ( .A(y[1519]), .B(x[1519]), .Z(n4272) );
  XNOR U6364 ( .A(y[1520]), .B(x[1520]), .Z(n4271) );
  XNOR U6365 ( .A(n4263), .B(n4264), .Z(n4274) );
  XNOR U6366 ( .A(y[1515]), .B(x[1515]), .Z(n4264) );
  XNOR U6367 ( .A(n4265), .B(n4266), .Z(n4263) );
  XNOR U6368 ( .A(y[1516]), .B(x[1516]), .Z(n4266) );
  XNOR U6369 ( .A(y[1517]), .B(x[1517]), .Z(n4265) );
  XOR U6370 ( .A(n4239), .B(n4240), .Z(n4258) );
  XNOR U6371 ( .A(n4255), .B(n4256), .Z(n4240) );
  XNOR U6372 ( .A(n4250), .B(n4251), .Z(n4256) );
  XNOR U6373 ( .A(n4252), .B(n4253), .Z(n4251) );
  XNOR U6374 ( .A(y[1513]), .B(x[1513]), .Z(n4253) );
  XNOR U6375 ( .A(y[1514]), .B(x[1514]), .Z(n4252) );
  XNOR U6376 ( .A(y[1512]), .B(x[1512]), .Z(n4250) );
  XNOR U6377 ( .A(n4244), .B(n4245), .Z(n4255) );
  XNOR U6378 ( .A(y[1509]), .B(x[1509]), .Z(n4245) );
  XNOR U6379 ( .A(n4246), .B(n4247), .Z(n4244) );
  XNOR U6380 ( .A(y[1510]), .B(x[1510]), .Z(n4247) );
  XNOR U6381 ( .A(y[1511]), .B(x[1511]), .Z(n4246) );
  XOR U6382 ( .A(n4238), .B(n4237), .Z(n4239) );
  XNOR U6383 ( .A(n4233), .B(n4234), .Z(n4237) );
  XNOR U6384 ( .A(y[1506]), .B(x[1506]), .Z(n4234) );
  XNOR U6385 ( .A(n4235), .B(n4236), .Z(n4233) );
  XNOR U6386 ( .A(y[1507]), .B(x[1507]), .Z(n4236) );
  XNOR U6387 ( .A(y[1508]), .B(x[1508]), .Z(n4235) );
  XNOR U6388 ( .A(n4227), .B(n4228), .Z(n4238) );
  XNOR U6389 ( .A(y[1503]), .B(x[1503]), .Z(n4228) );
  XNOR U6390 ( .A(n4229), .B(n4230), .Z(n4227) );
  XNOR U6391 ( .A(y[1504]), .B(x[1504]), .Z(n4230) );
  XNOR U6392 ( .A(y[1505]), .B(x[1505]), .Z(n4229) );
  NAND U6393 ( .A(n4294), .B(n4295), .Z(N13467) );
  NANDN U6394 ( .A(n4296), .B(n4297), .Z(n4295) );
  OR U6395 ( .A(n4298), .B(n4299), .Z(n4297) );
  NAND U6396 ( .A(n4298), .B(n4299), .Z(n4294) );
  XOR U6397 ( .A(n4298), .B(n4300), .Z(N13466) );
  XNOR U6398 ( .A(n4296), .B(n4299), .Z(n4300) );
  AND U6399 ( .A(n4301), .B(n4302), .Z(n4299) );
  NANDN U6400 ( .A(n4303), .B(n4304), .Z(n4302) );
  NANDN U6401 ( .A(n4305), .B(n4306), .Z(n4304) );
  NANDN U6402 ( .A(n4306), .B(n4305), .Z(n4301) );
  NAND U6403 ( .A(n4307), .B(n4308), .Z(n4296) );
  NANDN U6404 ( .A(n4309), .B(n4310), .Z(n4308) );
  OR U6405 ( .A(n4311), .B(n4312), .Z(n4310) );
  NAND U6406 ( .A(n4312), .B(n4311), .Z(n4307) );
  AND U6407 ( .A(n4313), .B(n4314), .Z(n4298) );
  NANDN U6408 ( .A(n4315), .B(n4316), .Z(n4314) );
  NANDN U6409 ( .A(n4317), .B(n4318), .Z(n4316) );
  NANDN U6410 ( .A(n4318), .B(n4317), .Z(n4313) );
  XOR U6411 ( .A(n4312), .B(n4319), .Z(N13465) );
  XOR U6412 ( .A(n4309), .B(n4311), .Z(n4319) );
  XNOR U6413 ( .A(n4305), .B(n4320), .Z(n4311) );
  XNOR U6414 ( .A(n4303), .B(n4306), .Z(n4320) );
  NAND U6415 ( .A(n4321), .B(n4322), .Z(n4306) );
  NAND U6416 ( .A(n4323), .B(n4324), .Z(n4322) );
  OR U6417 ( .A(n4325), .B(n4326), .Z(n4323) );
  NANDN U6418 ( .A(n4327), .B(n4325), .Z(n4321) );
  IV U6419 ( .A(n4326), .Z(n4327) );
  NAND U6420 ( .A(n4328), .B(n4329), .Z(n4303) );
  NAND U6421 ( .A(n4330), .B(n4331), .Z(n4329) );
  NANDN U6422 ( .A(n4332), .B(n4333), .Z(n4330) );
  NANDN U6423 ( .A(n4333), .B(n4332), .Z(n4328) );
  AND U6424 ( .A(n4334), .B(n4335), .Z(n4305) );
  NAND U6425 ( .A(n4336), .B(n4337), .Z(n4335) );
  OR U6426 ( .A(n4338), .B(n4339), .Z(n4336) );
  NANDN U6427 ( .A(n4340), .B(n4338), .Z(n4334) );
  NAND U6428 ( .A(n4341), .B(n4342), .Z(n4309) );
  NANDN U6429 ( .A(n4343), .B(n4344), .Z(n4342) );
  OR U6430 ( .A(n4345), .B(n4346), .Z(n4344) );
  NANDN U6431 ( .A(n4347), .B(n4345), .Z(n4341) );
  IV U6432 ( .A(n4346), .Z(n4347) );
  XNOR U6433 ( .A(n4317), .B(n4348), .Z(n4312) );
  XNOR U6434 ( .A(n4315), .B(n4318), .Z(n4348) );
  NAND U6435 ( .A(n4349), .B(n4350), .Z(n4318) );
  NAND U6436 ( .A(n4351), .B(n4352), .Z(n4350) );
  OR U6437 ( .A(n4353), .B(n4354), .Z(n4351) );
  NANDN U6438 ( .A(n4355), .B(n4353), .Z(n4349) );
  IV U6439 ( .A(n4354), .Z(n4355) );
  NAND U6440 ( .A(n4356), .B(n4357), .Z(n4315) );
  NAND U6441 ( .A(n4358), .B(n4359), .Z(n4357) );
  NANDN U6442 ( .A(n4360), .B(n4361), .Z(n4358) );
  NANDN U6443 ( .A(n4361), .B(n4360), .Z(n4356) );
  AND U6444 ( .A(n4362), .B(n4363), .Z(n4317) );
  NAND U6445 ( .A(n4364), .B(n4365), .Z(n4363) );
  OR U6446 ( .A(n4366), .B(n4367), .Z(n4364) );
  NANDN U6447 ( .A(n4368), .B(n4366), .Z(n4362) );
  XNOR U6448 ( .A(n4343), .B(n4369), .Z(N13464) );
  XOR U6449 ( .A(n4345), .B(n4346), .Z(n4369) );
  XNOR U6450 ( .A(n4359), .B(n4370), .Z(n4346) );
  XOR U6451 ( .A(n4360), .B(n4361), .Z(n4370) );
  XOR U6452 ( .A(n4366), .B(n4371), .Z(n4361) );
  XOR U6453 ( .A(n4365), .B(n4368), .Z(n4371) );
  IV U6454 ( .A(n4367), .Z(n4368) );
  NAND U6455 ( .A(n4372), .B(n4373), .Z(n4367) );
  OR U6456 ( .A(n4374), .B(n4375), .Z(n4373) );
  OR U6457 ( .A(n4376), .B(n4377), .Z(n4372) );
  NAND U6458 ( .A(n4378), .B(n4379), .Z(n4365) );
  OR U6459 ( .A(n4380), .B(n4381), .Z(n4379) );
  OR U6460 ( .A(n4382), .B(n4383), .Z(n4378) );
  NOR U6461 ( .A(n4384), .B(n4385), .Z(n4366) );
  ANDN U6462 ( .B(n4386), .A(n4387), .Z(n4360) );
  XNOR U6463 ( .A(n4353), .B(n4388), .Z(n4359) );
  XNOR U6464 ( .A(n4352), .B(n4354), .Z(n4388) );
  NAND U6465 ( .A(n4389), .B(n4390), .Z(n4354) );
  OR U6466 ( .A(n4391), .B(n4392), .Z(n4390) );
  OR U6467 ( .A(n4393), .B(n4394), .Z(n4389) );
  NAND U6468 ( .A(n4395), .B(n4396), .Z(n4352) );
  OR U6469 ( .A(n4397), .B(n4398), .Z(n4396) );
  OR U6470 ( .A(n4399), .B(n4400), .Z(n4395) );
  ANDN U6471 ( .B(n4401), .A(n4402), .Z(n4353) );
  IV U6472 ( .A(n4403), .Z(n4401) );
  ANDN U6473 ( .B(n4404), .A(n4405), .Z(n4345) );
  XOR U6474 ( .A(n4331), .B(n4406), .Z(n4343) );
  XOR U6475 ( .A(n4332), .B(n4333), .Z(n4406) );
  XOR U6476 ( .A(n4338), .B(n4407), .Z(n4333) );
  XOR U6477 ( .A(n4337), .B(n4340), .Z(n4407) );
  IV U6478 ( .A(n4339), .Z(n4340) );
  NAND U6479 ( .A(n4408), .B(n4409), .Z(n4339) );
  OR U6480 ( .A(n4410), .B(n4411), .Z(n4409) );
  OR U6481 ( .A(n4412), .B(n4413), .Z(n4408) );
  NAND U6482 ( .A(n4414), .B(n4415), .Z(n4337) );
  OR U6483 ( .A(n4416), .B(n4417), .Z(n4415) );
  OR U6484 ( .A(n4418), .B(n4419), .Z(n4414) );
  NOR U6485 ( .A(n4420), .B(n4421), .Z(n4338) );
  ANDN U6486 ( .B(n4422), .A(n4423), .Z(n4332) );
  IV U6487 ( .A(n4424), .Z(n4422) );
  XNOR U6488 ( .A(n4325), .B(n4425), .Z(n4331) );
  XNOR U6489 ( .A(n4324), .B(n4326), .Z(n4425) );
  NAND U6490 ( .A(n4426), .B(n4427), .Z(n4326) );
  OR U6491 ( .A(n4428), .B(n4429), .Z(n4427) );
  OR U6492 ( .A(n4430), .B(n4431), .Z(n4426) );
  NAND U6493 ( .A(n4432), .B(n4433), .Z(n4324) );
  OR U6494 ( .A(n4434), .B(n4435), .Z(n4433) );
  OR U6495 ( .A(n4436), .B(n4437), .Z(n4432) );
  ANDN U6496 ( .B(n4438), .A(n4439), .Z(n4325) );
  IV U6497 ( .A(n4440), .Z(n4438) );
  XNOR U6498 ( .A(n4405), .B(n4404), .Z(N13463) );
  XOR U6499 ( .A(n4424), .B(n4423), .Z(n4404) );
  XNOR U6500 ( .A(n4439), .B(n4440), .Z(n4423) );
  XNOR U6501 ( .A(n4434), .B(n4435), .Z(n4440) );
  XNOR U6502 ( .A(n4436), .B(n4437), .Z(n4435) );
  XNOR U6503 ( .A(y[1501]), .B(x[1501]), .Z(n4437) );
  XNOR U6504 ( .A(y[1502]), .B(x[1502]), .Z(n4436) );
  XNOR U6505 ( .A(y[1500]), .B(x[1500]), .Z(n4434) );
  XNOR U6506 ( .A(n4428), .B(n4429), .Z(n4439) );
  XNOR U6507 ( .A(y[1497]), .B(x[1497]), .Z(n4429) );
  XNOR U6508 ( .A(n4430), .B(n4431), .Z(n4428) );
  XNOR U6509 ( .A(y[1498]), .B(x[1498]), .Z(n4431) );
  XNOR U6510 ( .A(y[1499]), .B(x[1499]), .Z(n4430) );
  XNOR U6511 ( .A(n4421), .B(n4420), .Z(n4424) );
  XNOR U6512 ( .A(n4416), .B(n4417), .Z(n4420) );
  XNOR U6513 ( .A(y[1494]), .B(x[1494]), .Z(n4417) );
  XNOR U6514 ( .A(n4418), .B(n4419), .Z(n4416) );
  XNOR U6515 ( .A(y[1495]), .B(x[1495]), .Z(n4419) );
  XNOR U6516 ( .A(y[1496]), .B(x[1496]), .Z(n4418) );
  XNOR U6517 ( .A(n4410), .B(n4411), .Z(n4421) );
  XNOR U6518 ( .A(y[1491]), .B(x[1491]), .Z(n4411) );
  XNOR U6519 ( .A(n4412), .B(n4413), .Z(n4410) );
  XNOR U6520 ( .A(y[1492]), .B(x[1492]), .Z(n4413) );
  XNOR U6521 ( .A(y[1493]), .B(x[1493]), .Z(n4412) );
  XOR U6522 ( .A(n4386), .B(n4387), .Z(n4405) );
  XNOR U6523 ( .A(n4402), .B(n4403), .Z(n4387) );
  XNOR U6524 ( .A(n4397), .B(n4398), .Z(n4403) );
  XNOR U6525 ( .A(n4399), .B(n4400), .Z(n4398) );
  XNOR U6526 ( .A(y[1489]), .B(x[1489]), .Z(n4400) );
  XNOR U6527 ( .A(y[1490]), .B(x[1490]), .Z(n4399) );
  XNOR U6528 ( .A(y[1488]), .B(x[1488]), .Z(n4397) );
  XNOR U6529 ( .A(n4391), .B(n4392), .Z(n4402) );
  XNOR U6530 ( .A(y[1485]), .B(x[1485]), .Z(n4392) );
  XNOR U6531 ( .A(n4393), .B(n4394), .Z(n4391) );
  XNOR U6532 ( .A(y[1486]), .B(x[1486]), .Z(n4394) );
  XNOR U6533 ( .A(y[1487]), .B(x[1487]), .Z(n4393) );
  XOR U6534 ( .A(n4385), .B(n4384), .Z(n4386) );
  XNOR U6535 ( .A(n4380), .B(n4381), .Z(n4384) );
  XNOR U6536 ( .A(y[1482]), .B(x[1482]), .Z(n4381) );
  XNOR U6537 ( .A(n4382), .B(n4383), .Z(n4380) );
  XNOR U6538 ( .A(y[1483]), .B(x[1483]), .Z(n4383) );
  XNOR U6539 ( .A(y[1484]), .B(x[1484]), .Z(n4382) );
  XNOR U6540 ( .A(n4374), .B(n4375), .Z(n4385) );
  XNOR U6541 ( .A(y[1479]), .B(x[1479]), .Z(n4375) );
  XNOR U6542 ( .A(n4376), .B(n4377), .Z(n4374) );
  XNOR U6543 ( .A(y[1480]), .B(x[1480]), .Z(n4377) );
  XNOR U6544 ( .A(y[1481]), .B(x[1481]), .Z(n4376) );
  NAND U6545 ( .A(n4441), .B(n4442), .Z(N13456) );
  NANDN U6546 ( .A(n4443), .B(n4444), .Z(n4442) );
  OR U6547 ( .A(n4445), .B(n4446), .Z(n4444) );
  NAND U6548 ( .A(n4445), .B(n4446), .Z(n4441) );
  XOR U6549 ( .A(n4445), .B(n4447), .Z(N13455) );
  XNOR U6550 ( .A(n4443), .B(n4446), .Z(n4447) );
  AND U6551 ( .A(n4448), .B(n4449), .Z(n4446) );
  NANDN U6552 ( .A(n4450), .B(n4451), .Z(n4449) );
  NANDN U6553 ( .A(n4452), .B(n4453), .Z(n4451) );
  NANDN U6554 ( .A(n4453), .B(n4452), .Z(n4448) );
  NAND U6555 ( .A(n4454), .B(n4455), .Z(n4443) );
  NANDN U6556 ( .A(n4456), .B(n4457), .Z(n4455) );
  OR U6557 ( .A(n4458), .B(n4459), .Z(n4457) );
  NAND U6558 ( .A(n4459), .B(n4458), .Z(n4454) );
  AND U6559 ( .A(n4460), .B(n4461), .Z(n4445) );
  NANDN U6560 ( .A(n4462), .B(n4463), .Z(n4461) );
  NANDN U6561 ( .A(n4464), .B(n4465), .Z(n4463) );
  NANDN U6562 ( .A(n4465), .B(n4464), .Z(n4460) );
  XOR U6563 ( .A(n4459), .B(n4466), .Z(N13454) );
  XOR U6564 ( .A(n4456), .B(n4458), .Z(n4466) );
  XNOR U6565 ( .A(n4452), .B(n4467), .Z(n4458) );
  XNOR U6566 ( .A(n4450), .B(n4453), .Z(n4467) );
  NAND U6567 ( .A(n4468), .B(n4469), .Z(n4453) );
  NAND U6568 ( .A(n4470), .B(n4471), .Z(n4469) );
  OR U6569 ( .A(n4472), .B(n4473), .Z(n4470) );
  NANDN U6570 ( .A(n4474), .B(n4472), .Z(n4468) );
  IV U6571 ( .A(n4473), .Z(n4474) );
  NAND U6572 ( .A(n4475), .B(n4476), .Z(n4450) );
  NAND U6573 ( .A(n4477), .B(n4478), .Z(n4476) );
  NANDN U6574 ( .A(n4479), .B(n4480), .Z(n4477) );
  NANDN U6575 ( .A(n4480), .B(n4479), .Z(n4475) );
  AND U6576 ( .A(n4481), .B(n4482), .Z(n4452) );
  NAND U6577 ( .A(n4483), .B(n4484), .Z(n4482) );
  OR U6578 ( .A(n4485), .B(n4486), .Z(n4483) );
  NANDN U6579 ( .A(n4487), .B(n4485), .Z(n4481) );
  NAND U6580 ( .A(n4488), .B(n4489), .Z(n4456) );
  NANDN U6581 ( .A(n4490), .B(n4491), .Z(n4489) );
  OR U6582 ( .A(n4492), .B(n4493), .Z(n4491) );
  NANDN U6583 ( .A(n4494), .B(n4492), .Z(n4488) );
  IV U6584 ( .A(n4493), .Z(n4494) );
  XNOR U6585 ( .A(n4464), .B(n4495), .Z(n4459) );
  XNOR U6586 ( .A(n4462), .B(n4465), .Z(n4495) );
  NAND U6587 ( .A(n4496), .B(n4497), .Z(n4465) );
  NAND U6588 ( .A(n4498), .B(n4499), .Z(n4497) );
  OR U6589 ( .A(n4500), .B(n4501), .Z(n4498) );
  NANDN U6590 ( .A(n4502), .B(n4500), .Z(n4496) );
  IV U6591 ( .A(n4501), .Z(n4502) );
  NAND U6592 ( .A(n4503), .B(n4504), .Z(n4462) );
  NAND U6593 ( .A(n4505), .B(n4506), .Z(n4504) );
  NANDN U6594 ( .A(n4507), .B(n4508), .Z(n4505) );
  NANDN U6595 ( .A(n4508), .B(n4507), .Z(n4503) );
  AND U6596 ( .A(n4509), .B(n4510), .Z(n4464) );
  NAND U6597 ( .A(n4511), .B(n4512), .Z(n4510) );
  OR U6598 ( .A(n4513), .B(n4514), .Z(n4511) );
  NANDN U6599 ( .A(n4515), .B(n4513), .Z(n4509) );
  XNOR U6600 ( .A(n4490), .B(n4516), .Z(N13453) );
  XOR U6601 ( .A(n4492), .B(n4493), .Z(n4516) );
  XNOR U6602 ( .A(n4506), .B(n4517), .Z(n4493) );
  XOR U6603 ( .A(n4507), .B(n4508), .Z(n4517) );
  XOR U6604 ( .A(n4513), .B(n4518), .Z(n4508) );
  XOR U6605 ( .A(n4512), .B(n4515), .Z(n4518) );
  IV U6606 ( .A(n4514), .Z(n4515) );
  NAND U6607 ( .A(n4519), .B(n4520), .Z(n4514) );
  OR U6608 ( .A(n4521), .B(n4522), .Z(n4520) );
  OR U6609 ( .A(n4523), .B(n4524), .Z(n4519) );
  NAND U6610 ( .A(n4525), .B(n4526), .Z(n4512) );
  OR U6611 ( .A(n4527), .B(n4528), .Z(n4526) );
  OR U6612 ( .A(n4529), .B(n4530), .Z(n4525) );
  NOR U6613 ( .A(n4531), .B(n4532), .Z(n4513) );
  ANDN U6614 ( .B(n4533), .A(n4534), .Z(n4507) );
  XNOR U6615 ( .A(n4500), .B(n4535), .Z(n4506) );
  XNOR U6616 ( .A(n4499), .B(n4501), .Z(n4535) );
  NAND U6617 ( .A(n4536), .B(n4537), .Z(n4501) );
  OR U6618 ( .A(n4538), .B(n4539), .Z(n4537) );
  OR U6619 ( .A(n4540), .B(n4541), .Z(n4536) );
  NAND U6620 ( .A(n4542), .B(n4543), .Z(n4499) );
  OR U6621 ( .A(n4544), .B(n4545), .Z(n4543) );
  OR U6622 ( .A(n4546), .B(n4547), .Z(n4542) );
  ANDN U6623 ( .B(n4548), .A(n4549), .Z(n4500) );
  IV U6624 ( .A(n4550), .Z(n4548) );
  ANDN U6625 ( .B(n4551), .A(n4552), .Z(n4492) );
  XOR U6626 ( .A(n4478), .B(n4553), .Z(n4490) );
  XOR U6627 ( .A(n4479), .B(n4480), .Z(n4553) );
  XOR U6628 ( .A(n4485), .B(n4554), .Z(n4480) );
  XOR U6629 ( .A(n4484), .B(n4487), .Z(n4554) );
  IV U6630 ( .A(n4486), .Z(n4487) );
  NAND U6631 ( .A(n4555), .B(n4556), .Z(n4486) );
  OR U6632 ( .A(n4557), .B(n4558), .Z(n4556) );
  OR U6633 ( .A(n4559), .B(n4560), .Z(n4555) );
  NAND U6634 ( .A(n4561), .B(n4562), .Z(n4484) );
  OR U6635 ( .A(n4563), .B(n4564), .Z(n4562) );
  OR U6636 ( .A(n4565), .B(n4566), .Z(n4561) );
  NOR U6637 ( .A(n4567), .B(n4568), .Z(n4485) );
  ANDN U6638 ( .B(n4569), .A(n4570), .Z(n4479) );
  IV U6639 ( .A(n4571), .Z(n4569) );
  XNOR U6640 ( .A(n4472), .B(n4572), .Z(n4478) );
  XNOR U6641 ( .A(n4471), .B(n4473), .Z(n4572) );
  NAND U6642 ( .A(n4573), .B(n4574), .Z(n4473) );
  OR U6643 ( .A(n4575), .B(n4576), .Z(n4574) );
  OR U6644 ( .A(n4577), .B(n4578), .Z(n4573) );
  NAND U6645 ( .A(n4579), .B(n4580), .Z(n4471) );
  OR U6646 ( .A(n4581), .B(n4582), .Z(n4580) );
  OR U6647 ( .A(n4583), .B(n4584), .Z(n4579) );
  ANDN U6648 ( .B(n4585), .A(n4586), .Z(n4472) );
  IV U6649 ( .A(n4587), .Z(n4585) );
  XNOR U6650 ( .A(n4552), .B(n4551), .Z(N13452) );
  XOR U6651 ( .A(n4571), .B(n4570), .Z(n4551) );
  XNOR U6652 ( .A(n4586), .B(n4587), .Z(n4570) );
  XNOR U6653 ( .A(n4581), .B(n4582), .Z(n4587) );
  XNOR U6654 ( .A(n4583), .B(n4584), .Z(n4582) );
  XNOR U6655 ( .A(y[1477]), .B(x[1477]), .Z(n4584) );
  XNOR U6656 ( .A(y[1478]), .B(x[1478]), .Z(n4583) );
  XNOR U6657 ( .A(y[1476]), .B(x[1476]), .Z(n4581) );
  XNOR U6658 ( .A(n4575), .B(n4576), .Z(n4586) );
  XNOR U6659 ( .A(y[1473]), .B(x[1473]), .Z(n4576) );
  XNOR U6660 ( .A(n4577), .B(n4578), .Z(n4575) );
  XNOR U6661 ( .A(y[1474]), .B(x[1474]), .Z(n4578) );
  XNOR U6662 ( .A(y[1475]), .B(x[1475]), .Z(n4577) );
  XNOR U6663 ( .A(n4568), .B(n4567), .Z(n4571) );
  XNOR U6664 ( .A(n4563), .B(n4564), .Z(n4567) );
  XNOR U6665 ( .A(y[1470]), .B(x[1470]), .Z(n4564) );
  XNOR U6666 ( .A(n4565), .B(n4566), .Z(n4563) );
  XNOR U6667 ( .A(y[1471]), .B(x[1471]), .Z(n4566) );
  XNOR U6668 ( .A(y[1472]), .B(x[1472]), .Z(n4565) );
  XNOR U6669 ( .A(n4557), .B(n4558), .Z(n4568) );
  XNOR U6670 ( .A(y[1467]), .B(x[1467]), .Z(n4558) );
  XNOR U6671 ( .A(n4559), .B(n4560), .Z(n4557) );
  XNOR U6672 ( .A(y[1468]), .B(x[1468]), .Z(n4560) );
  XNOR U6673 ( .A(y[1469]), .B(x[1469]), .Z(n4559) );
  XOR U6674 ( .A(n4533), .B(n4534), .Z(n4552) );
  XNOR U6675 ( .A(n4549), .B(n4550), .Z(n4534) );
  XNOR U6676 ( .A(n4544), .B(n4545), .Z(n4550) );
  XNOR U6677 ( .A(n4546), .B(n4547), .Z(n4545) );
  XNOR U6678 ( .A(y[1465]), .B(x[1465]), .Z(n4547) );
  XNOR U6679 ( .A(y[1466]), .B(x[1466]), .Z(n4546) );
  XNOR U6680 ( .A(y[1464]), .B(x[1464]), .Z(n4544) );
  XNOR U6681 ( .A(n4538), .B(n4539), .Z(n4549) );
  XNOR U6682 ( .A(y[1461]), .B(x[1461]), .Z(n4539) );
  XNOR U6683 ( .A(n4540), .B(n4541), .Z(n4538) );
  XNOR U6684 ( .A(y[1462]), .B(x[1462]), .Z(n4541) );
  XNOR U6685 ( .A(y[1463]), .B(x[1463]), .Z(n4540) );
  XOR U6686 ( .A(n4532), .B(n4531), .Z(n4533) );
  XNOR U6687 ( .A(n4527), .B(n4528), .Z(n4531) );
  XNOR U6688 ( .A(y[1458]), .B(x[1458]), .Z(n4528) );
  XNOR U6689 ( .A(n4529), .B(n4530), .Z(n4527) );
  XNOR U6690 ( .A(y[1459]), .B(x[1459]), .Z(n4530) );
  XNOR U6691 ( .A(y[1460]), .B(x[1460]), .Z(n4529) );
  XNOR U6692 ( .A(n4521), .B(n4522), .Z(n4532) );
  XNOR U6693 ( .A(y[1455]), .B(x[1455]), .Z(n4522) );
  XNOR U6694 ( .A(n4523), .B(n4524), .Z(n4521) );
  XNOR U6695 ( .A(y[1456]), .B(x[1456]), .Z(n4524) );
  XNOR U6696 ( .A(y[1457]), .B(x[1457]), .Z(n4523) );
  NAND U6697 ( .A(n4588), .B(n4589), .Z(N13445) );
  NANDN U6698 ( .A(n4590), .B(n4591), .Z(n4589) );
  OR U6699 ( .A(n4592), .B(n4593), .Z(n4591) );
  NAND U6700 ( .A(n4592), .B(n4593), .Z(n4588) );
  XOR U6701 ( .A(n4592), .B(n4594), .Z(N13444) );
  XNOR U6702 ( .A(n4590), .B(n4593), .Z(n4594) );
  AND U6703 ( .A(n4595), .B(n4596), .Z(n4593) );
  NANDN U6704 ( .A(n4597), .B(n4598), .Z(n4596) );
  NANDN U6705 ( .A(n4599), .B(n4600), .Z(n4598) );
  NANDN U6706 ( .A(n4600), .B(n4599), .Z(n4595) );
  NAND U6707 ( .A(n4601), .B(n4602), .Z(n4590) );
  NANDN U6708 ( .A(n4603), .B(n4604), .Z(n4602) );
  OR U6709 ( .A(n4605), .B(n4606), .Z(n4604) );
  NAND U6710 ( .A(n4606), .B(n4605), .Z(n4601) );
  AND U6711 ( .A(n4607), .B(n4608), .Z(n4592) );
  NANDN U6712 ( .A(n4609), .B(n4610), .Z(n4608) );
  NANDN U6713 ( .A(n4611), .B(n4612), .Z(n4610) );
  NANDN U6714 ( .A(n4612), .B(n4611), .Z(n4607) );
  XOR U6715 ( .A(n4606), .B(n4613), .Z(N13443) );
  XOR U6716 ( .A(n4603), .B(n4605), .Z(n4613) );
  XNOR U6717 ( .A(n4599), .B(n4614), .Z(n4605) );
  XNOR U6718 ( .A(n4597), .B(n4600), .Z(n4614) );
  NAND U6719 ( .A(n4615), .B(n4616), .Z(n4600) );
  NAND U6720 ( .A(n4617), .B(n4618), .Z(n4616) );
  OR U6721 ( .A(n4619), .B(n4620), .Z(n4617) );
  NANDN U6722 ( .A(n4621), .B(n4619), .Z(n4615) );
  IV U6723 ( .A(n4620), .Z(n4621) );
  NAND U6724 ( .A(n4622), .B(n4623), .Z(n4597) );
  NAND U6725 ( .A(n4624), .B(n4625), .Z(n4623) );
  NANDN U6726 ( .A(n4626), .B(n4627), .Z(n4624) );
  NANDN U6727 ( .A(n4627), .B(n4626), .Z(n4622) );
  AND U6728 ( .A(n4628), .B(n4629), .Z(n4599) );
  NAND U6729 ( .A(n4630), .B(n4631), .Z(n4629) );
  OR U6730 ( .A(n4632), .B(n4633), .Z(n4630) );
  NANDN U6731 ( .A(n4634), .B(n4632), .Z(n4628) );
  NAND U6732 ( .A(n4635), .B(n4636), .Z(n4603) );
  NANDN U6733 ( .A(n4637), .B(n4638), .Z(n4636) );
  OR U6734 ( .A(n4639), .B(n4640), .Z(n4638) );
  NANDN U6735 ( .A(n4641), .B(n4639), .Z(n4635) );
  IV U6736 ( .A(n4640), .Z(n4641) );
  XNOR U6737 ( .A(n4611), .B(n4642), .Z(n4606) );
  XNOR U6738 ( .A(n4609), .B(n4612), .Z(n4642) );
  NAND U6739 ( .A(n4643), .B(n4644), .Z(n4612) );
  NAND U6740 ( .A(n4645), .B(n4646), .Z(n4644) );
  OR U6741 ( .A(n4647), .B(n4648), .Z(n4645) );
  NANDN U6742 ( .A(n4649), .B(n4647), .Z(n4643) );
  IV U6743 ( .A(n4648), .Z(n4649) );
  NAND U6744 ( .A(n4650), .B(n4651), .Z(n4609) );
  NAND U6745 ( .A(n4652), .B(n4653), .Z(n4651) );
  NANDN U6746 ( .A(n4654), .B(n4655), .Z(n4652) );
  NANDN U6747 ( .A(n4655), .B(n4654), .Z(n4650) );
  AND U6748 ( .A(n4656), .B(n4657), .Z(n4611) );
  NAND U6749 ( .A(n4658), .B(n4659), .Z(n4657) );
  OR U6750 ( .A(n4660), .B(n4661), .Z(n4658) );
  NANDN U6751 ( .A(n4662), .B(n4660), .Z(n4656) );
  XNOR U6752 ( .A(n4637), .B(n4663), .Z(N13442) );
  XOR U6753 ( .A(n4639), .B(n4640), .Z(n4663) );
  XNOR U6754 ( .A(n4653), .B(n4664), .Z(n4640) );
  XOR U6755 ( .A(n4654), .B(n4655), .Z(n4664) );
  XOR U6756 ( .A(n4660), .B(n4665), .Z(n4655) );
  XOR U6757 ( .A(n4659), .B(n4662), .Z(n4665) );
  IV U6758 ( .A(n4661), .Z(n4662) );
  NAND U6759 ( .A(n4666), .B(n4667), .Z(n4661) );
  OR U6760 ( .A(n4668), .B(n4669), .Z(n4667) );
  OR U6761 ( .A(n4670), .B(n4671), .Z(n4666) );
  NAND U6762 ( .A(n4672), .B(n4673), .Z(n4659) );
  OR U6763 ( .A(n4674), .B(n4675), .Z(n4673) );
  OR U6764 ( .A(n4676), .B(n4677), .Z(n4672) );
  NOR U6765 ( .A(n4678), .B(n4679), .Z(n4660) );
  ANDN U6766 ( .B(n4680), .A(n4681), .Z(n4654) );
  XNOR U6767 ( .A(n4647), .B(n4682), .Z(n4653) );
  XNOR U6768 ( .A(n4646), .B(n4648), .Z(n4682) );
  NAND U6769 ( .A(n4683), .B(n4684), .Z(n4648) );
  OR U6770 ( .A(n4685), .B(n4686), .Z(n4684) );
  OR U6771 ( .A(n4687), .B(n4688), .Z(n4683) );
  NAND U6772 ( .A(n4689), .B(n4690), .Z(n4646) );
  OR U6773 ( .A(n4691), .B(n4692), .Z(n4690) );
  OR U6774 ( .A(n4693), .B(n4694), .Z(n4689) );
  ANDN U6775 ( .B(n4695), .A(n4696), .Z(n4647) );
  IV U6776 ( .A(n4697), .Z(n4695) );
  ANDN U6777 ( .B(n4698), .A(n4699), .Z(n4639) );
  XOR U6778 ( .A(n4625), .B(n4700), .Z(n4637) );
  XOR U6779 ( .A(n4626), .B(n4627), .Z(n4700) );
  XOR U6780 ( .A(n4632), .B(n4701), .Z(n4627) );
  XOR U6781 ( .A(n4631), .B(n4634), .Z(n4701) );
  IV U6782 ( .A(n4633), .Z(n4634) );
  NAND U6783 ( .A(n4702), .B(n4703), .Z(n4633) );
  OR U6784 ( .A(n4704), .B(n4705), .Z(n4703) );
  OR U6785 ( .A(n4706), .B(n4707), .Z(n4702) );
  NAND U6786 ( .A(n4708), .B(n4709), .Z(n4631) );
  OR U6787 ( .A(n4710), .B(n4711), .Z(n4709) );
  OR U6788 ( .A(n4712), .B(n4713), .Z(n4708) );
  NOR U6789 ( .A(n4714), .B(n4715), .Z(n4632) );
  ANDN U6790 ( .B(n4716), .A(n4717), .Z(n4626) );
  IV U6791 ( .A(n4718), .Z(n4716) );
  XNOR U6792 ( .A(n4619), .B(n4719), .Z(n4625) );
  XNOR U6793 ( .A(n4618), .B(n4620), .Z(n4719) );
  NAND U6794 ( .A(n4720), .B(n4721), .Z(n4620) );
  OR U6795 ( .A(n4722), .B(n4723), .Z(n4721) );
  OR U6796 ( .A(n4724), .B(n4725), .Z(n4720) );
  NAND U6797 ( .A(n4726), .B(n4727), .Z(n4618) );
  OR U6798 ( .A(n4728), .B(n4729), .Z(n4727) );
  OR U6799 ( .A(n4730), .B(n4731), .Z(n4726) );
  ANDN U6800 ( .B(n4732), .A(n4733), .Z(n4619) );
  IV U6801 ( .A(n4734), .Z(n4732) );
  XNOR U6802 ( .A(n4699), .B(n4698), .Z(N13441) );
  XOR U6803 ( .A(n4718), .B(n4717), .Z(n4698) );
  XNOR U6804 ( .A(n4733), .B(n4734), .Z(n4717) );
  XNOR U6805 ( .A(n4728), .B(n4729), .Z(n4734) );
  XNOR U6806 ( .A(n4730), .B(n4731), .Z(n4729) );
  XNOR U6807 ( .A(y[1453]), .B(x[1453]), .Z(n4731) );
  XNOR U6808 ( .A(y[1454]), .B(x[1454]), .Z(n4730) );
  XNOR U6809 ( .A(y[1452]), .B(x[1452]), .Z(n4728) );
  XNOR U6810 ( .A(n4722), .B(n4723), .Z(n4733) );
  XNOR U6811 ( .A(y[1449]), .B(x[1449]), .Z(n4723) );
  XNOR U6812 ( .A(n4724), .B(n4725), .Z(n4722) );
  XNOR U6813 ( .A(y[1450]), .B(x[1450]), .Z(n4725) );
  XNOR U6814 ( .A(y[1451]), .B(x[1451]), .Z(n4724) );
  XNOR U6815 ( .A(n4715), .B(n4714), .Z(n4718) );
  XNOR U6816 ( .A(n4710), .B(n4711), .Z(n4714) );
  XNOR U6817 ( .A(y[1446]), .B(x[1446]), .Z(n4711) );
  XNOR U6818 ( .A(n4712), .B(n4713), .Z(n4710) );
  XNOR U6819 ( .A(y[1447]), .B(x[1447]), .Z(n4713) );
  XNOR U6820 ( .A(y[1448]), .B(x[1448]), .Z(n4712) );
  XNOR U6821 ( .A(n4704), .B(n4705), .Z(n4715) );
  XNOR U6822 ( .A(y[1443]), .B(x[1443]), .Z(n4705) );
  XNOR U6823 ( .A(n4706), .B(n4707), .Z(n4704) );
  XNOR U6824 ( .A(y[1444]), .B(x[1444]), .Z(n4707) );
  XNOR U6825 ( .A(y[1445]), .B(x[1445]), .Z(n4706) );
  XOR U6826 ( .A(n4680), .B(n4681), .Z(n4699) );
  XNOR U6827 ( .A(n4696), .B(n4697), .Z(n4681) );
  XNOR U6828 ( .A(n4691), .B(n4692), .Z(n4697) );
  XNOR U6829 ( .A(n4693), .B(n4694), .Z(n4692) );
  XNOR U6830 ( .A(y[1441]), .B(x[1441]), .Z(n4694) );
  XNOR U6831 ( .A(y[1442]), .B(x[1442]), .Z(n4693) );
  XNOR U6832 ( .A(y[1440]), .B(x[1440]), .Z(n4691) );
  XNOR U6833 ( .A(n4685), .B(n4686), .Z(n4696) );
  XNOR U6834 ( .A(y[1437]), .B(x[1437]), .Z(n4686) );
  XNOR U6835 ( .A(n4687), .B(n4688), .Z(n4685) );
  XNOR U6836 ( .A(y[1438]), .B(x[1438]), .Z(n4688) );
  XNOR U6837 ( .A(y[1439]), .B(x[1439]), .Z(n4687) );
  XOR U6838 ( .A(n4679), .B(n4678), .Z(n4680) );
  XNOR U6839 ( .A(n4674), .B(n4675), .Z(n4678) );
  XNOR U6840 ( .A(y[1434]), .B(x[1434]), .Z(n4675) );
  XNOR U6841 ( .A(n4676), .B(n4677), .Z(n4674) );
  XNOR U6842 ( .A(y[1435]), .B(x[1435]), .Z(n4677) );
  XNOR U6843 ( .A(y[1436]), .B(x[1436]), .Z(n4676) );
  XNOR U6844 ( .A(n4668), .B(n4669), .Z(n4679) );
  XNOR U6845 ( .A(y[1431]), .B(x[1431]), .Z(n4669) );
  XNOR U6846 ( .A(n4670), .B(n4671), .Z(n4668) );
  XNOR U6847 ( .A(y[1432]), .B(x[1432]), .Z(n4671) );
  XNOR U6848 ( .A(y[1433]), .B(x[1433]), .Z(n4670) );
  NAND U6849 ( .A(n4735), .B(n4736), .Z(N13434) );
  NANDN U6850 ( .A(n4737), .B(n4738), .Z(n4736) );
  OR U6851 ( .A(n4739), .B(n4740), .Z(n4738) );
  NAND U6852 ( .A(n4739), .B(n4740), .Z(n4735) );
  XOR U6853 ( .A(n4739), .B(n4741), .Z(N13433) );
  XNOR U6854 ( .A(n4737), .B(n4740), .Z(n4741) );
  AND U6855 ( .A(n4742), .B(n4743), .Z(n4740) );
  NANDN U6856 ( .A(n4744), .B(n4745), .Z(n4743) );
  NANDN U6857 ( .A(n4746), .B(n4747), .Z(n4745) );
  NANDN U6858 ( .A(n4747), .B(n4746), .Z(n4742) );
  NAND U6859 ( .A(n4748), .B(n4749), .Z(n4737) );
  NANDN U6860 ( .A(n4750), .B(n4751), .Z(n4749) );
  OR U6861 ( .A(n4752), .B(n4753), .Z(n4751) );
  NAND U6862 ( .A(n4753), .B(n4752), .Z(n4748) );
  AND U6863 ( .A(n4754), .B(n4755), .Z(n4739) );
  NANDN U6864 ( .A(n4756), .B(n4757), .Z(n4755) );
  NANDN U6865 ( .A(n4758), .B(n4759), .Z(n4757) );
  NANDN U6866 ( .A(n4759), .B(n4758), .Z(n4754) );
  XOR U6867 ( .A(n4753), .B(n4760), .Z(N13432) );
  XOR U6868 ( .A(n4750), .B(n4752), .Z(n4760) );
  XNOR U6869 ( .A(n4746), .B(n4761), .Z(n4752) );
  XNOR U6870 ( .A(n4744), .B(n4747), .Z(n4761) );
  NAND U6871 ( .A(n4762), .B(n4763), .Z(n4747) );
  NAND U6872 ( .A(n4764), .B(n4765), .Z(n4763) );
  OR U6873 ( .A(n4766), .B(n4767), .Z(n4764) );
  NANDN U6874 ( .A(n4768), .B(n4766), .Z(n4762) );
  IV U6875 ( .A(n4767), .Z(n4768) );
  NAND U6876 ( .A(n4769), .B(n4770), .Z(n4744) );
  NAND U6877 ( .A(n4771), .B(n4772), .Z(n4770) );
  NANDN U6878 ( .A(n4773), .B(n4774), .Z(n4771) );
  NANDN U6879 ( .A(n4774), .B(n4773), .Z(n4769) );
  AND U6880 ( .A(n4775), .B(n4776), .Z(n4746) );
  NAND U6881 ( .A(n4777), .B(n4778), .Z(n4776) );
  OR U6882 ( .A(n4779), .B(n4780), .Z(n4777) );
  NANDN U6883 ( .A(n4781), .B(n4779), .Z(n4775) );
  NAND U6884 ( .A(n4782), .B(n4783), .Z(n4750) );
  NANDN U6885 ( .A(n4784), .B(n4785), .Z(n4783) );
  OR U6886 ( .A(n4786), .B(n4787), .Z(n4785) );
  NANDN U6887 ( .A(n4788), .B(n4786), .Z(n4782) );
  IV U6888 ( .A(n4787), .Z(n4788) );
  XNOR U6889 ( .A(n4758), .B(n4789), .Z(n4753) );
  XNOR U6890 ( .A(n4756), .B(n4759), .Z(n4789) );
  NAND U6891 ( .A(n4790), .B(n4791), .Z(n4759) );
  NAND U6892 ( .A(n4792), .B(n4793), .Z(n4791) );
  OR U6893 ( .A(n4794), .B(n4795), .Z(n4792) );
  NANDN U6894 ( .A(n4796), .B(n4794), .Z(n4790) );
  IV U6895 ( .A(n4795), .Z(n4796) );
  NAND U6896 ( .A(n4797), .B(n4798), .Z(n4756) );
  NAND U6897 ( .A(n4799), .B(n4800), .Z(n4798) );
  NANDN U6898 ( .A(n4801), .B(n4802), .Z(n4799) );
  NANDN U6899 ( .A(n4802), .B(n4801), .Z(n4797) );
  AND U6900 ( .A(n4803), .B(n4804), .Z(n4758) );
  NAND U6901 ( .A(n4805), .B(n4806), .Z(n4804) );
  OR U6902 ( .A(n4807), .B(n4808), .Z(n4805) );
  NANDN U6903 ( .A(n4809), .B(n4807), .Z(n4803) );
  XNOR U6904 ( .A(n4784), .B(n4810), .Z(N13431) );
  XOR U6905 ( .A(n4786), .B(n4787), .Z(n4810) );
  XNOR U6906 ( .A(n4800), .B(n4811), .Z(n4787) );
  XOR U6907 ( .A(n4801), .B(n4802), .Z(n4811) );
  XOR U6908 ( .A(n4807), .B(n4812), .Z(n4802) );
  XOR U6909 ( .A(n4806), .B(n4809), .Z(n4812) );
  IV U6910 ( .A(n4808), .Z(n4809) );
  NAND U6911 ( .A(n4813), .B(n4814), .Z(n4808) );
  OR U6912 ( .A(n4815), .B(n4816), .Z(n4814) );
  OR U6913 ( .A(n4817), .B(n4818), .Z(n4813) );
  NAND U6914 ( .A(n4819), .B(n4820), .Z(n4806) );
  OR U6915 ( .A(n4821), .B(n4822), .Z(n4820) );
  OR U6916 ( .A(n4823), .B(n4824), .Z(n4819) );
  NOR U6917 ( .A(n4825), .B(n4826), .Z(n4807) );
  ANDN U6918 ( .B(n4827), .A(n4828), .Z(n4801) );
  XNOR U6919 ( .A(n4794), .B(n4829), .Z(n4800) );
  XNOR U6920 ( .A(n4793), .B(n4795), .Z(n4829) );
  NAND U6921 ( .A(n4830), .B(n4831), .Z(n4795) );
  OR U6922 ( .A(n4832), .B(n4833), .Z(n4831) );
  OR U6923 ( .A(n4834), .B(n4835), .Z(n4830) );
  NAND U6924 ( .A(n4836), .B(n4837), .Z(n4793) );
  OR U6925 ( .A(n4838), .B(n4839), .Z(n4837) );
  OR U6926 ( .A(n4840), .B(n4841), .Z(n4836) );
  ANDN U6927 ( .B(n4842), .A(n4843), .Z(n4794) );
  IV U6928 ( .A(n4844), .Z(n4842) );
  ANDN U6929 ( .B(n4845), .A(n4846), .Z(n4786) );
  XOR U6930 ( .A(n4772), .B(n4847), .Z(n4784) );
  XOR U6931 ( .A(n4773), .B(n4774), .Z(n4847) );
  XOR U6932 ( .A(n4779), .B(n4848), .Z(n4774) );
  XOR U6933 ( .A(n4778), .B(n4781), .Z(n4848) );
  IV U6934 ( .A(n4780), .Z(n4781) );
  NAND U6935 ( .A(n4849), .B(n4850), .Z(n4780) );
  OR U6936 ( .A(n4851), .B(n4852), .Z(n4850) );
  OR U6937 ( .A(n4853), .B(n4854), .Z(n4849) );
  NAND U6938 ( .A(n4855), .B(n4856), .Z(n4778) );
  OR U6939 ( .A(n4857), .B(n4858), .Z(n4856) );
  OR U6940 ( .A(n4859), .B(n4860), .Z(n4855) );
  NOR U6941 ( .A(n4861), .B(n4862), .Z(n4779) );
  ANDN U6942 ( .B(n4863), .A(n4864), .Z(n4773) );
  IV U6943 ( .A(n4865), .Z(n4863) );
  XNOR U6944 ( .A(n4766), .B(n4866), .Z(n4772) );
  XNOR U6945 ( .A(n4765), .B(n4767), .Z(n4866) );
  NAND U6946 ( .A(n4867), .B(n4868), .Z(n4767) );
  OR U6947 ( .A(n4869), .B(n4870), .Z(n4868) );
  OR U6948 ( .A(n4871), .B(n4872), .Z(n4867) );
  NAND U6949 ( .A(n4873), .B(n4874), .Z(n4765) );
  OR U6950 ( .A(n4875), .B(n4876), .Z(n4874) );
  OR U6951 ( .A(n4877), .B(n4878), .Z(n4873) );
  ANDN U6952 ( .B(n4879), .A(n4880), .Z(n4766) );
  IV U6953 ( .A(n4881), .Z(n4879) );
  XNOR U6954 ( .A(n4846), .B(n4845), .Z(N13430) );
  XOR U6955 ( .A(n4865), .B(n4864), .Z(n4845) );
  XNOR U6956 ( .A(n4880), .B(n4881), .Z(n4864) );
  XNOR U6957 ( .A(n4875), .B(n4876), .Z(n4881) );
  XNOR U6958 ( .A(n4877), .B(n4878), .Z(n4876) );
  XNOR U6959 ( .A(y[1429]), .B(x[1429]), .Z(n4878) );
  XNOR U6960 ( .A(y[1430]), .B(x[1430]), .Z(n4877) );
  XNOR U6961 ( .A(y[1428]), .B(x[1428]), .Z(n4875) );
  XNOR U6962 ( .A(n4869), .B(n4870), .Z(n4880) );
  XNOR U6963 ( .A(y[1425]), .B(x[1425]), .Z(n4870) );
  XNOR U6964 ( .A(n4871), .B(n4872), .Z(n4869) );
  XNOR U6965 ( .A(y[1426]), .B(x[1426]), .Z(n4872) );
  XNOR U6966 ( .A(y[1427]), .B(x[1427]), .Z(n4871) );
  XNOR U6967 ( .A(n4862), .B(n4861), .Z(n4865) );
  XNOR U6968 ( .A(n4857), .B(n4858), .Z(n4861) );
  XNOR U6969 ( .A(y[1422]), .B(x[1422]), .Z(n4858) );
  XNOR U6970 ( .A(n4859), .B(n4860), .Z(n4857) );
  XNOR U6971 ( .A(y[1423]), .B(x[1423]), .Z(n4860) );
  XNOR U6972 ( .A(y[1424]), .B(x[1424]), .Z(n4859) );
  XNOR U6973 ( .A(n4851), .B(n4852), .Z(n4862) );
  XNOR U6974 ( .A(y[1419]), .B(x[1419]), .Z(n4852) );
  XNOR U6975 ( .A(n4853), .B(n4854), .Z(n4851) );
  XNOR U6976 ( .A(y[1420]), .B(x[1420]), .Z(n4854) );
  XNOR U6977 ( .A(y[1421]), .B(x[1421]), .Z(n4853) );
  XOR U6978 ( .A(n4827), .B(n4828), .Z(n4846) );
  XNOR U6979 ( .A(n4843), .B(n4844), .Z(n4828) );
  XNOR U6980 ( .A(n4838), .B(n4839), .Z(n4844) );
  XNOR U6981 ( .A(n4840), .B(n4841), .Z(n4839) );
  XNOR U6982 ( .A(y[1417]), .B(x[1417]), .Z(n4841) );
  XNOR U6983 ( .A(y[1418]), .B(x[1418]), .Z(n4840) );
  XNOR U6984 ( .A(y[1416]), .B(x[1416]), .Z(n4838) );
  XNOR U6985 ( .A(n4832), .B(n4833), .Z(n4843) );
  XNOR U6986 ( .A(y[1413]), .B(x[1413]), .Z(n4833) );
  XNOR U6987 ( .A(n4834), .B(n4835), .Z(n4832) );
  XNOR U6988 ( .A(y[1414]), .B(x[1414]), .Z(n4835) );
  XNOR U6989 ( .A(y[1415]), .B(x[1415]), .Z(n4834) );
  XOR U6990 ( .A(n4826), .B(n4825), .Z(n4827) );
  XNOR U6991 ( .A(n4821), .B(n4822), .Z(n4825) );
  XNOR U6992 ( .A(y[1410]), .B(x[1410]), .Z(n4822) );
  XNOR U6993 ( .A(n4823), .B(n4824), .Z(n4821) );
  XNOR U6994 ( .A(y[1411]), .B(x[1411]), .Z(n4824) );
  XNOR U6995 ( .A(y[1412]), .B(x[1412]), .Z(n4823) );
  XNOR U6996 ( .A(n4815), .B(n4816), .Z(n4826) );
  XNOR U6997 ( .A(y[1407]), .B(x[1407]), .Z(n4816) );
  XNOR U6998 ( .A(n4817), .B(n4818), .Z(n4815) );
  XNOR U6999 ( .A(y[1408]), .B(x[1408]), .Z(n4818) );
  XNOR U7000 ( .A(y[1409]), .B(x[1409]), .Z(n4817) );
  NAND U7001 ( .A(n4882), .B(n4883), .Z(N13423) );
  NANDN U7002 ( .A(n4884), .B(n4885), .Z(n4883) );
  OR U7003 ( .A(n4886), .B(n4887), .Z(n4885) );
  NAND U7004 ( .A(n4886), .B(n4887), .Z(n4882) );
  XOR U7005 ( .A(n4886), .B(n4888), .Z(N13422) );
  XNOR U7006 ( .A(n4884), .B(n4887), .Z(n4888) );
  AND U7007 ( .A(n4889), .B(n4890), .Z(n4887) );
  NANDN U7008 ( .A(n4891), .B(n4892), .Z(n4890) );
  NANDN U7009 ( .A(n4893), .B(n4894), .Z(n4892) );
  NANDN U7010 ( .A(n4894), .B(n4893), .Z(n4889) );
  NAND U7011 ( .A(n4895), .B(n4896), .Z(n4884) );
  NANDN U7012 ( .A(n4897), .B(n4898), .Z(n4896) );
  OR U7013 ( .A(n4899), .B(n4900), .Z(n4898) );
  NAND U7014 ( .A(n4900), .B(n4899), .Z(n4895) );
  AND U7015 ( .A(n4901), .B(n4902), .Z(n4886) );
  NANDN U7016 ( .A(n4903), .B(n4904), .Z(n4902) );
  NANDN U7017 ( .A(n4905), .B(n4906), .Z(n4904) );
  NANDN U7018 ( .A(n4906), .B(n4905), .Z(n4901) );
  XOR U7019 ( .A(n4900), .B(n4907), .Z(N13421) );
  XOR U7020 ( .A(n4897), .B(n4899), .Z(n4907) );
  XNOR U7021 ( .A(n4893), .B(n4908), .Z(n4899) );
  XNOR U7022 ( .A(n4891), .B(n4894), .Z(n4908) );
  NAND U7023 ( .A(n4909), .B(n4910), .Z(n4894) );
  NAND U7024 ( .A(n4911), .B(n4912), .Z(n4910) );
  OR U7025 ( .A(n4913), .B(n4914), .Z(n4911) );
  NANDN U7026 ( .A(n4915), .B(n4913), .Z(n4909) );
  IV U7027 ( .A(n4914), .Z(n4915) );
  NAND U7028 ( .A(n4916), .B(n4917), .Z(n4891) );
  NAND U7029 ( .A(n4918), .B(n4919), .Z(n4917) );
  NANDN U7030 ( .A(n4920), .B(n4921), .Z(n4918) );
  NANDN U7031 ( .A(n4921), .B(n4920), .Z(n4916) );
  AND U7032 ( .A(n4922), .B(n4923), .Z(n4893) );
  NAND U7033 ( .A(n4924), .B(n4925), .Z(n4923) );
  OR U7034 ( .A(n4926), .B(n4927), .Z(n4924) );
  NANDN U7035 ( .A(n4928), .B(n4926), .Z(n4922) );
  NAND U7036 ( .A(n4929), .B(n4930), .Z(n4897) );
  NANDN U7037 ( .A(n4931), .B(n4932), .Z(n4930) );
  OR U7038 ( .A(n4933), .B(n4934), .Z(n4932) );
  NANDN U7039 ( .A(n4935), .B(n4933), .Z(n4929) );
  IV U7040 ( .A(n4934), .Z(n4935) );
  XNOR U7041 ( .A(n4905), .B(n4936), .Z(n4900) );
  XNOR U7042 ( .A(n4903), .B(n4906), .Z(n4936) );
  NAND U7043 ( .A(n4937), .B(n4938), .Z(n4906) );
  NAND U7044 ( .A(n4939), .B(n4940), .Z(n4938) );
  OR U7045 ( .A(n4941), .B(n4942), .Z(n4939) );
  NANDN U7046 ( .A(n4943), .B(n4941), .Z(n4937) );
  IV U7047 ( .A(n4942), .Z(n4943) );
  NAND U7048 ( .A(n4944), .B(n4945), .Z(n4903) );
  NAND U7049 ( .A(n4946), .B(n4947), .Z(n4945) );
  NANDN U7050 ( .A(n4948), .B(n4949), .Z(n4946) );
  NANDN U7051 ( .A(n4949), .B(n4948), .Z(n4944) );
  AND U7052 ( .A(n4950), .B(n4951), .Z(n4905) );
  NAND U7053 ( .A(n4952), .B(n4953), .Z(n4951) );
  OR U7054 ( .A(n4954), .B(n4955), .Z(n4952) );
  NANDN U7055 ( .A(n4956), .B(n4954), .Z(n4950) );
  XNOR U7056 ( .A(n4931), .B(n4957), .Z(N13420) );
  XOR U7057 ( .A(n4933), .B(n4934), .Z(n4957) );
  XNOR U7058 ( .A(n4947), .B(n4958), .Z(n4934) );
  XOR U7059 ( .A(n4948), .B(n4949), .Z(n4958) );
  XOR U7060 ( .A(n4954), .B(n4959), .Z(n4949) );
  XOR U7061 ( .A(n4953), .B(n4956), .Z(n4959) );
  IV U7062 ( .A(n4955), .Z(n4956) );
  NAND U7063 ( .A(n4960), .B(n4961), .Z(n4955) );
  OR U7064 ( .A(n4962), .B(n4963), .Z(n4961) );
  OR U7065 ( .A(n4964), .B(n4965), .Z(n4960) );
  NAND U7066 ( .A(n4966), .B(n4967), .Z(n4953) );
  OR U7067 ( .A(n4968), .B(n4969), .Z(n4967) );
  OR U7068 ( .A(n4970), .B(n4971), .Z(n4966) );
  NOR U7069 ( .A(n4972), .B(n4973), .Z(n4954) );
  ANDN U7070 ( .B(n4974), .A(n4975), .Z(n4948) );
  XNOR U7071 ( .A(n4941), .B(n4976), .Z(n4947) );
  XNOR U7072 ( .A(n4940), .B(n4942), .Z(n4976) );
  NAND U7073 ( .A(n4977), .B(n4978), .Z(n4942) );
  OR U7074 ( .A(n4979), .B(n4980), .Z(n4978) );
  OR U7075 ( .A(n4981), .B(n4982), .Z(n4977) );
  NAND U7076 ( .A(n4983), .B(n4984), .Z(n4940) );
  OR U7077 ( .A(n4985), .B(n4986), .Z(n4984) );
  OR U7078 ( .A(n4987), .B(n4988), .Z(n4983) );
  ANDN U7079 ( .B(n4989), .A(n4990), .Z(n4941) );
  IV U7080 ( .A(n4991), .Z(n4989) );
  ANDN U7081 ( .B(n4992), .A(n4993), .Z(n4933) );
  XOR U7082 ( .A(n4919), .B(n4994), .Z(n4931) );
  XOR U7083 ( .A(n4920), .B(n4921), .Z(n4994) );
  XOR U7084 ( .A(n4926), .B(n4995), .Z(n4921) );
  XOR U7085 ( .A(n4925), .B(n4928), .Z(n4995) );
  IV U7086 ( .A(n4927), .Z(n4928) );
  NAND U7087 ( .A(n4996), .B(n4997), .Z(n4927) );
  OR U7088 ( .A(n4998), .B(n4999), .Z(n4997) );
  OR U7089 ( .A(n5000), .B(n5001), .Z(n4996) );
  NAND U7090 ( .A(n5002), .B(n5003), .Z(n4925) );
  OR U7091 ( .A(n5004), .B(n5005), .Z(n5003) );
  OR U7092 ( .A(n5006), .B(n5007), .Z(n5002) );
  NOR U7093 ( .A(n5008), .B(n5009), .Z(n4926) );
  ANDN U7094 ( .B(n5010), .A(n5011), .Z(n4920) );
  IV U7095 ( .A(n5012), .Z(n5010) );
  XNOR U7096 ( .A(n4913), .B(n5013), .Z(n4919) );
  XNOR U7097 ( .A(n4912), .B(n4914), .Z(n5013) );
  NAND U7098 ( .A(n5014), .B(n5015), .Z(n4914) );
  OR U7099 ( .A(n5016), .B(n5017), .Z(n5015) );
  OR U7100 ( .A(n5018), .B(n5019), .Z(n5014) );
  NAND U7101 ( .A(n5020), .B(n5021), .Z(n4912) );
  OR U7102 ( .A(n5022), .B(n5023), .Z(n5021) );
  OR U7103 ( .A(n5024), .B(n5025), .Z(n5020) );
  ANDN U7104 ( .B(n5026), .A(n5027), .Z(n4913) );
  IV U7105 ( .A(n5028), .Z(n5026) );
  XNOR U7106 ( .A(n4993), .B(n4992), .Z(N13419) );
  XOR U7107 ( .A(n5012), .B(n5011), .Z(n4992) );
  XNOR U7108 ( .A(n5027), .B(n5028), .Z(n5011) );
  XNOR U7109 ( .A(n5022), .B(n5023), .Z(n5028) );
  XNOR U7110 ( .A(n5024), .B(n5025), .Z(n5023) );
  XNOR U7111 ( .A(y[1405]), .B(x[1405]), .Z(n5025) );
  XNOR U7112 ( .A(y[1406]), .B(x[1406]), .Z(n5024) );
  XNOR U7113 ( .A(y[1404]), .B(x[1404]), .Z(n5022) );
  XNOR U7114 ( .A(n5016), .B(n5017), .Z(n5027) );
  XNOR U7115 ( .A(y[1401]), .B(x[1401]), .Z(n5017) );
  XNOR U7116 ( .A(n5018), .B(n5019), .Z(n5016) );
  XNOR U7117 ( .A(y[1402]), .B(x[1402]), .Z(n5019) );
  XNOR U7118 ( .A(y[1403]), .B(x[1403]), .Z(n5018) );
  XNOR U7119 ( .A(n5009), .B(n5008), .Z(n5012) );
  XNOR U7120 ( .A(n5004), .B(n5005), .Z(n5008) );
  XNOR U7121 ( .A(y[1398]), .B(x[1398]), .Z(n5005) );
  XNOR U7122 ( .A(n5006), .B(n5007), .Z(n5004) );
  XNOR U7123 ( .A(y[1399]), .B(x[1399]), .Z(n5007) );
  XNOR U7124 ( .A(y[1400]), .B(x[1400]), .Z(n5006) );
  XNOR U7125 ( .A(n4998), .B(n4999), .Z(n5009) );
  XNOR U7126 ( .A(y[1395]), .B(x[1395]), .Z(n4999) );
  XNOR U7127 ( .A(n5000), .B(n5001), .Z(n4998) );
  XNOR U7128 ( .A(y[1396]), .B(x[1396]), .Z(n5001) );
  XNOR U7129 ( .A(y[1397]), .B(x[1397]), .Z(n5000) );
  XOR U7130 ( .A(n4974), .B(n4975), .Z(n4993) );
  XNOR U7131 ( .A(n4990), .B(n4991), .Z(n4975) );
  XNOR U7132 ( .A(n4985), .B(n4986), .Z(n4991) );
  XNOR U7133 ( .A(n4987), .B(n4988), .Z(n4986) );
  XNOR U7134 ( .A(y[1393]), .B(x[1393]), .Z(n4988) );
  XNOR U7135 ( .A(y[1394]), .B(x[1394]), .Z(n4987) );
  XNOR U7136 ( .A(y[1392]), .B(x[1392]), .Z(n4985) );
  XNOR U7137 ( .A(n4979), .B(n4980), .Z(n4990) );
  XNOR U7138 ( .A(y[1389]), .B(x[1389]), .Z(n4980) );
  XNOR U7139 ( .A(n4981), .B(n4982), .Z(n4979) );
  XNOR U7140 ( .A(y[1390]), .B(x[1390]), .Z(n4982) );
  XNOR U7141 ( .A(y[1391]), .B(x[1391]), .Z(n4981) );
  XOR U7142 ( .A(n4973), .B(n4972), .Z(n4974) );
  XNOR U7143 ( .A(n4968), .B(n4969), .Z(n4972) );
  XNOR U7144 ( .A(y[1386]), .B(x[1386]), .Z(n4969) );
  XNOR U7145 ( .A(n4970), .B(n4971), .Z(n4968) );
  XNOR U7146 ( .A(y[1387]), .B(x[1387]), .Z(n4971) );
  XNOR U7147 ( .A(y[1388]), .B(x[1388]), .Z(n4970) );
  XNOR U7148 ( .A(n4962), .B(n4963), .Z(n4973) );
  XNOR U7149 ( .A(y[1383]), .B(x[1383]), .Z(n4963) );
  XNOR U7150 ( .A(n4964), .B(n4965), .Z(n4962) );
  XNOR U7151 ( .A(y[1384]), .B(x[1384]), .Z(n4965) );
  XNOR U7152 ( .A(y[1385]), .B(x[1385]), .Z(n4964) );
  NAND U7153 ( .A(n5029), .B(n5030), .Z(N13412) );
  NANDN U7154 ( .A(n5031), .B(n5032), .Z(n5030) );
  OR U7155 ( .A(n5033), .B(n5034), .Z(n5032) );
  NAND U7156 ( .A(n5033), .B(n5034), .Z(n5029) );
  XOR U7157 ( .A(n5033), .B(n5035), .Z(N13411) );
  XNOR U7158 ( .A(n5031), .B(n5034), .Z(n5035) );
  AND U7159 ( .A(n5036), .B(n5037), .Z(n5034) );
  NANDN U7160 ( .A(n5038), .B(n5039), .Z(n5037) );
  NANDN U7161 ( .A(n5040), .B(n5041), .Z(n5039) );
  NANDN U7162 ( .A(n5041), .B(n5040), .Z(n5036) );
  NAND U7163 ( .A(n5042), .B(n5043), .Z(n5031) );
  NANDN U7164 ( .A(n5044), .B(n5045), .Z(n5043) );
  OR U7165 ( .A(n5046), .B(n5047), .Z(n5045) );
  NAND U7166 ( .A(n5047), .B(n5046), .Z(n5042) );
  AND U7167 ( .A(n5048), .B(n5049), .Z(n5033) );
  NANDN U7168 ( .A(n5050), .B(n5051), .Z(n5049) );
  NANDN U7169 ( .A(n5052), .B(n5053), .Z(n5051) );
  NANDN U7170 ( .A(n5053), .B(n5052), .Z(n5048) );
  XOR U7171 ( .A(n5047), .B(n5054), .Z(N13410) );
  XOR U7172 ( .A(n5044), .B(n5046), .Z(n5054) );
  XNOR U7173 ( .A(n5040), .B(n5055), .Z(n5046) );
  XNOR U7174 ( .A(n5038), .B(n5041), .Z(n5055) );
  NAND U7175 ( .A(n5056), .B(n5057), .Z(n5041) );
  NAND U7176 ( .A(n5058), .B(n5059), .Z(n5057) );
  OR U7177 ( .A(n5060), .B(n5061), .Z(n5058) );
  NANDN U7178 ( .A(n5062), .B(n5060), .Z(n5056) );
  IV U7179 ( .A(n5061), .Z(n5062) );
  NAND U7180 ( .A(n5063), .B(n5064), .Z(n5038) );
  NAND U7181 ( .A(n5065), .B(n5066), .Z(n5064) );
  NANDN U7182 ( .A(n5067), .B(n5068), .Z(n5065) );
  NANDN U7183 ( .A(n5068), .B(n5067), .Z(n5063) );
  AND U7184 ( .A(n5069), .B(n5070), .Z(n5040) );
  NAND U7185 ( .A(n5071), .B(n5072), .Z(n5070) );
  OR U7186 ( .A(n5073), .B(n5074), .Z(n5071) );
  NANDN U7187 ( .A(n5075), .B(n5073), .Z(n5069) );
  NAND U7188 ( .A(n5076), .B(n5077), .Z(n5044) );
  NANDN U7189 ( .A(n5078), .B(n5079), .Z(n5077) );
  OR U7190 ( .A(n5080), .B(n5081), .Z(n5079) );
  NANDN U7191 ( .A(n5082), .B(n5080), .Z(n5076) );
  IV U7192 ( .A(n5081), .Z(n5082) );
  XNOR U7193 ( .A(n5052), .B(n5083), .Z(n5047) );
  XNOR U7194 ( .A(n5050), .B(n5053), .Z(n5083) );
  NAND U7195 ( .A(n5084), .B(n5085), .Z(n5053) );
  NAND U7196 ( .A(n5086), .B(n5087), .Z(n5085) );
  OR U7197 ( .A(n5088), .B(n5089), .Z(n5086) );
  NANDN U7198 ( .A(n5090), .B(n5088), .Z(n5084) );
  IV U7199 ( .A(n5089), .Z(n5090) );
  NAND U7200 ( .A(n5091), .B(n5092), .Z(n5050) );
  NAND U7201 ( .A(n5093), .B(n5094), .Z(n5092) );
  NANDN U7202 ( .A(n5095), .B(n5096), .Z(n5093) );
  NANDN U7203 ( .A(n5096), .B(n5095), .Z(n5091) );
  AND U7204 ( .A(n5097), .B(n5098), .Z(n5052) );
  NAND U7205 ( .A(n5099), .B(n5100), .Z(n5098) );
  OR U7206 ( .A(n5101), .B(n5102), .Z(n5099) );
  NANDN U7207 ( .A(n5103), .B(n5101), .Z(n5097) );
  XNOR U7208 ( .A(n5078), .B(n5104), .Z(N13409) );
  XOR U7209 ( .A(n5080), .B(n5081), .Z(n5104) );
  XNOR U7210 ( .A(n5094), .B(n5105), .Z(n5081) );
  XOR U7211 ( .A(n5095), .B(n5096), .Z(n5105) );
  XOR U7212 ( .A(n5101), .B(n5106), .Z(n5096) );
  XOR U7213 ( .A(n5100), .B(n5103), .Z(n5106) );
  IV U7214 ( .A(n5102), .Z(n5103) );
  NAND U7215 ( .A(n5107), .B(n5108), .Z(n5102) );
  OR U7216 ( .A(n5109), .B(n5110), .Z(n5108) );
  OR U7217 ( .A(n5111), .B(n5112), .Z(n5107) );
  NAND U7218 ( .A(n5113), .B(n5114), .Z(n5100) );
  OR U7219 ( .A(n5115), .B(n5116), .Z(n5114) );
  OR U7220 ( .A(n5117), .B(n5118), .Z(n5113) );
  NOR U7221 ( .A(n5119), .B(n5120), .Z(n5101) );
  ANDN U7222 ( .B(n5121), .A(n5122), .Z(n5095) );
  XNOR U7223 ( .A(n5088), .B(n5123), .Z(n5094) );
  XNOR U7224 ( .A(n5087), .B(n5089), .Z(n5123) );
  NAND U7225 ( .A(n5124), .B(n5125), .Z(n5089) );
  OR U7226 ( .A(n5126), .B(n5127), .Z(n5125) );
  OR U7227 ( .A(n5128), .B(n5129), .Z(n5124) );
  NAND U7228 ( .A(n5130), .B(n5131), .Z(n5087) );
  OR U7229 ( .A(n5132), .B(n5133), .Z(n5131) );
  OR U7230 ( .A(n5134), .B(n5135), .Z(n5130) );
  ANDN U7231 ( .B(n5136), .A(n5137), .Z(n5088) );
  IV U7232 ( .A(n5138), .Z(n5136) );
  ANDN U7233 ( .B(n5139), .A(n5140), .Z(n5080) );
  XOR U7234 ( .A(n5066), .B(n5141), .Z(n5078) );
  XOR U7235 ( .A(n5067), .B(n5068), .Z(n5141) );
  XOR U7236 ( .A(n5073), .B(n5142), .Z(n5068) );
  XOR U7237 ( .A(n5072), .B(n5075), .Z(n5142) );
  IV U7238 ( .A(n5074), .Z(n5075) );
  NAND U7239 ( .A(n5143), .B(n5144), .Z(n5074) );
  OR U7240 ( .A(n5145), .B(n5146), .Z(n5144) );
  OR U7241 ( .A(n5147), .B(n5148), .Z(n5143) );
  NAND U7242 ( .A(n5149), .B(n5150), .Z(n5072) );
  OR U7243 ( .A(n5151), .B(n5152), .Z(n5150) );
  OR U7244 ( .A(n5153), .B(n5154), .Z(n5149) );
  NOR U7245 ( .A(n5155), .B(n5156), .Z(n5073) );
  ANDN U7246 ( .B(n5157), .A(n5158), .Z(n5067) );
  IV U7247 ( .A(n5159), .Z(n5157) );
  XNOR U7248 ( .A(n5060), .B(n5160), .Z(n5066) );
  XNOR U7249 ( .A(n5059), .B(n5061), .Z(n5160) );
  NAND U7250 ( .A(n5161), .B(n5162), .Z(n5061) );
  OR U7251 ( .A(n5163), .B(n5164), .Z(n5162) );
  OR U7252 ( .A(n5165), .B(n5166), .Z(n5161) );
  NAND U7253 ( .A(n5167), .B(n5168), .Z(n5059) );
  OR U7254 ( .A(n5169), .B(n5170), .Z(n5168) );
  OR U7255 ( .A(n5171), .B(n5172), .Z(n5167) );
  ANDN U7256 ( .B(n5173), .A(n5174), .Z(n5060) );
  IV U7257 ( .A(n5175), .Z(n5173) );
  XNOR U7258 ( .A(n5140), .B(n5139), .Z(N13408) );
  XOR U7259 ( .A(n5159), .B(n5158), .Z(n5139) );
  XNOR U7260 ( .A(n5174), .B(n5175), .Z(n5158) );
  XNOR U7261 ( .A(n5169), .B(n5170), .Z(n5175) );
  XNOR U7262 ( .A(n5171), .B(n5172), .Z(n5170) );
  XNOR U7263 ( .A(y[1381]), .B(x[1381]), .Z(n5172) );
  XNOR U7264 ( .A(y[1382]), .B(x[1382]), .Z(n5171) );
  XNOR U7265 ( .A(y[1380]), .B(x[1380]), .Z(n5169) );
  XNOR U7266 ( .A(n5163), .B(n5164), .Z(n5174) );
  XNOR U7267 ( .A(y[1377]), .B(x[1377]), .Z(n5164) );
  XNOR U7268 ( .A(n5165), .B(n5166), .Z(n5163) );
  XNOR U7269 ( .A(y[1378]), .B(x[1378]), .Z(n5166) );
  XNOR U7270 ( .A(y[1379]), .B(x[1379]), .Z(n5165) );
  XNOR U7271 ( .A(n5156), .B(n5155), .Z(n5159) );
  XNOR U7272 ( .A(n5151), .B(n5152), .Z(n5155) );
  XNOR U7273 ( .A(y[1374]), .B(x[1374]), .Z(n5152) );
  XNOR U7274 ( .A(n5153), .B(n5154), .Z(n5151) );
  XNOR U7275 ( .A(y[1375]), .B(x[1375]), .Z(n5154) );
  XNOR U7276 ( .A(y[1376]), .B(x[1376]), .Z(n5153) );
  XNOR U7277 ( .A(n5145), .B(n5146), .Z(n5156) );
  XNOR U7278 ( .A(y[1371]), .B(x[1371]), .Z(n5146) );
  XNOR U7279 ( .A(n5147), .B(n5148), .Z(n5145) );
  XNOR U7280 ( .A(y[1372]), .B(x[1372]), .Z(n5148) );
  XNOR U7281 ( .A(y[1373]), .B(x[1373]), .Z(n5147) );
  XOR U7282 ( .A(n5121), .B(n5122), .Z(n5140) );
  XNOR U7283 ( .A(n5137), .B(n5138), .Z(n5122) );
  XNOR U7284 ( .A(n5132), .B(n5133), .Z(n5138) );
  XNOR U7285 ( .A(n5134), .B(n5135), .Z(n5133) );
  XNOR U7286 ( .A(y[1369]), .B(x[1369]), .Z(n5135) );
  XNOR U7287 ( .A(y[1370]), .B(x[1370]), .Z(n5134) );
  XNOR U7288 ( .A(y[1368]), .B(x[1368]), .Z(n5132) );
  XNOR U7289 ( .A(n5126), .B(n5127), .Z(n5137) );
  XNOR U7290 ( .A(y[1365]), .B(x[1365]), .Z(n5127) );
  XNOR U7291 ( .A(n5128), .B(n5129), .Z(n5126) );
  XNOR U7292 ( .A(y[1366]), .B(x[1366]), .Z(n5129) );
  XNOR U7293 ( .A(y[1367]), .B(x[1367]), .Z(n5128) );
  XOR U7294 ( .A(n5120), .B(n5119), .Z(n5121) );
  XNOR U7295 ( .A(n5115), .B(n5116), .Z(n5119) );
  XNOR U7296 ( .A(y[1362]), .B(x[1362]), .Z(n5116) );
  XNOR U7297 ( .A(n5117), .B(n5118), .Z(n5115) );
  XNOR U7298 ( .A(y[1363]), .B(x[1363]), .Z(n5118) );
  XNOR U7299 ( .A(y[1364]), .B(x[1364]), .Z(n5117) );
  XNOR U7300 ( .A(n5109), .B(n5110), .Z(n5120) );
  XNOR U7301 ( .A(y[1359]), .B(x[1359]), .Z(n5110) );
  XNOR U7302 ( .A(n5111), .B(n5112), .Z(n5109) );
  XNOR U7303 ( .A(y[1360]), .B(x[1360]), .Z(n5112) );
  XNOR U7304 ( .A(y[1361]), .B(x[1361]), .Z(n5111) );
  NAND U7305 ( .A(n5176), .B(n5177), .Z(N13401) );
  NANDN U7306 ( .A(n5178), .B(n5179), .Z(n5177) );
  OR U7307 ( .A(n5180), .B(n5181), .Z(n5179) );
  NAND U7308 ( .A(n5180), .B(n5181), .Z(n5176) );
  XOR U7309 ( .A(n5180), .B(n5182), .Z(N13400) );
  XNOR U7310 ( .A(n5178), .B(n5181), .Z(n5182) );
  AND U7311 ( .A(n5183), .B(n5184), .Z(n5181) );
  NANDN U7312 ( .A(n5185), .B(n5186), .Z(n5184) );
  NANDN U7313 ( .A(n5187), .B(n5188), .Z(n5186) );
  NANDN U7314 ( .A(n5188), .B(n5187), .Z(n5183) );
  NAND U7315 ( .A(n5189), .B(n5190), .Z(n5178) );
  NANDN U7316 ( .A(n5191), .B(n5192), .Z(n5190) );
  OR U7317 ( .A(n5193), .B(n5194), .Z(n5192) );
  NAND U7318 ( .A(n5194), .B(n5193), .Z(n5189) );
  AND U7319 ( .A(n5195), .B(n5196), .Z(n5180) );
  NANDN U7320 ( .A(n5197), .B(n5198), .Z(n5196) );
  NANDN U7321 ( .A(n5199), .B(n5200), .Z(n5198) );
  NANDN U7322 ( .A(n5200), .B(n5199), .Z(n5195) );
  XOR U7323 ( .A(n5194), .B(n5201), .Z(N13399) );
  XOR U7324 ( .A(n5191), .B(n5193), .Z(n5201) );
  XNOR U7325 ( .A(n5187), .B(n5202), .Z(n5193) );
  XNOR U7326 ( .A(n5185), .B(n5188), .Z(n5202) );
  NAND U7327 ( .A(n5203), .B(n5204), .Z(n5188) );
  NAND U7328 ( .A(n5205), .B(n5206), .Z(n5204) );
  OR U7329 ( .A(n5207), .B(n5208), .Z(n5205) );
  NANDN U7330 ( .A(n5209), .B(n5207), .Z(n5203) );
  IV U7331 ( .A(n5208), .Z(n5209) );
  NAND U7332 ( .A(n5210), .B(n5211), .Z(n5185) );
  NAND U7333 ( .A(n5212), .B(n5213), .Z(n5211) );
  NANDN U7334 ( .A(n5214), .B(n5215), .Z(n5212) );
  NANDN U7335 ( .A(n5215), .B(n5214), .Z(n5210) );
  AND U7336 ( .A(n5216), .B(n5217), .Z(n5187) );
  NAND U7337 ( .A(n5218), .B(n5219), .Z(n5217) );
  OR U7338 ( .A(n5220), .B(n5221), .Z(n5218) );
  NANDN U7339 ( .A(n5222), .B(n5220), .Z(n5216) );
  NAND U7340 ( .A(n5223), .B(n5224), .Z(n5191) );
  NANDN U7341 ( .A(n5225), .B(n5226), .Z(n5224) );
  OR U7342 ( .A(n5227), .B(n5228), .Z(n5226) );
  NANDN U7343 ( .A(n5229), .B(n5227), .Z(n5223) );
  IV U7344 ( .A(n5228), .Z(n5229) );
  XNOR U7345 ( .A(n5199), .B(n5230), .Z(n5194) );
  XNOR U7346 ( .A(n5197), .B(n5200), .Z(n5230) );
  NAND U7347 ( .A(n5231), .B(n5232), .Z(n5200) );
  NAND U7348 ( .A(n5233), .B(n5234), .Z(n5232) );
  OR U7349 ( .A(n5235), .B(n5236), .Z(n5233) );
  NANDN U7350 ( .A(n5237), .B(n5235), .Z(n5231) );
  IV U7351 ( .A(n5236), .Z(n5237) );
  NAND U7352 ( .A(n5238), .B(n5239), .Z(n5197) );
  NAND U7353 ( .A(n5240), .B(n5241), .Z(n5239) );
  NANDN U7354 ( .A(n5242), .B(n5243), .Z(n5240) );
  NANDN U7355 ( .A(n5243), .B(n5242), .Z(n5238) );
  AND U7356 ( .A(n5244), .B(n5245), .Z(n5199) );
  NAND U7357 ( .A(n5246), .B(n5247), .Z(n5245) );
  OR U7358 ( .A(n5248), .B(n5249), .Z(n5246) );
  NANDN U7359 ( .A(n5250), .B(n5248), .Z(n5244) );
  XNOR U7360 ( .A(n5225), .B(n5251), .Z(N13398) );
  XOR U7361 ( .A(n5227), .B(n5228), .Z(n5251) );
  XNOR U7362 ( .A(n5241), .B(n5252), .Z(n5228) );
  XOR U7363 ( .A(n5242), .B(n5243), .Z(n5252) );
  XOR U7364 ( .A(n5248), .B(n5253), .Z(n5243) );
  XOR U7365 ( .A(n5247), .B(n5250), .Z(n5253) );
  IV U7366 ( .A(n5249), .Z(n5250) );
  NAND U7367 ( .A(n5254), .B(n5255), .Z(n5249) );
  OR U7368 ( .A(n5256), .B(n5257), .Z(n5255) );
  OR U7369 ( .A(n5258), .B(n5259), .Z(n5254) );
  NAND U7370 ( .A(n5260), .B(n5261), .Z(n5247) );
  OR U7371 ( .A(n5262), .B(n5263), .Z(n5261) );
  OR U7372 ( .A(n5264), .B(n5265), .Z(n5260) );
  NOR U7373 ( .A(n5266), .B(n5267), .Z(n5248) );
  ANDN U7374 ( .B(n5268), .A(n5269), .Z(n5242) );
  XNOR U7375 ( .A(n5235), .B(n5270), .Z(n5241) );
  XNOR U7376 ( .A(n5234), .B(n5236), .Z(n5270) );
  NAND U7377 ( .A(n5271), .B(n5272), .Z(n5236) );
  OR U7378 ( .A(n5273), .B(n5274), .Z(n5272) );
  OR U7379 ( .A(n5275), .B(n5276), .Z(n5271) );
  NAND U7380 ( .A(n5277), .B(n5278), .Z(n5234) );
  OR U7381 ( .A(n5279), .B(n5280), .Z(n5278) );
  OR U7382 ( .A(n5281), .B(n5282), .Z(n5277) );
  ANDN U7383 ( .B(n5283), .A(n5284), .Z(n5235) );
  IV U7384 ( .A(n5285), .Z(n5283) );
  ANDN U7385 ( .B(n5286), .A(n5287), .Z(n5227) );
  XOR U7386 ( .A(n5213), .B(n5288), .Z(n5225) );
  XOR U7387 ( .A(n5214), .B(n5215), .Z(n5288) );
  XOR U7388 ( .A(n5220), .B(n5289), .Z(n5215) );
  XOR U7389 ( .A(n5219), .B(n5222), .Z(n5289) );
  IV U7390 ( .A(n5221), .Z(n5222) );
  NAND U7391 ( .A(n5290), .B(n5291), .Z(n5221) );
  OR U7392 ( .A(n5292), .B(n5293), .Z(n5291) );
  OR U7393 ( .A(n5294), .B(n5295), .Z(n5290) );
  NAND U7394 ( .A(n5296), .B(n5297), .Z(n5219) );
  OR U7395 ( .A(n5298), .B(n5299), .Z(n5297) );
  OR U7396 ( .A(n5300), .B(n5301), .Z(n5296) );
  NOR U7397 ( .A(n5302), .B(n5303), .Z(n5220) );
  ANDN U7398 ( .B(n5304), .A(n5305), .Z(n5214) );
  IV U7399 ( .A(n5306), .Z(n5304) );
  XNOR U7400 ( .A(n5207), .B(n5307), .Z(n5213) );
  XNOR U7401 ( .A(n5206), .B(n5208), .Z(n5307) );
  NAND U7402 ( .A(n5308), .B(n5309), .Z(n5208) );
  OR U7403 ( .A(n5310), .B(n5311), .Z(n5309) );
  OR U7404 ( .A(n5312), .B(n5313), .Z(n5308) );
  NAND U7405 ( .A(n5314), .B(n5315), .Z(n5206) );
  OR U7406 ( .A(n5316), .B(n5317), .Z(n5315) );
  OR U7407 ( .A(n5318), .B(n5319), .Z(n5314) );
  ANDN U7408 ( .B(n5320), .A(n5321), .Z(n5207) );
  IV U7409 ( .A(n5322), .Z(n5320) );
  XNOR U7410 ( .A(n5287), .B(n5286), .Z(N13397) );
  XOR U7411 ( .A(n5306), .B(n5305), .Z(n5286) );
  XNOR U7412 ( .A(n5321), .B(n5322), .Z(n5305) );
  XNOR U7413 ( .A(n5316), .B(n5317), .Z(n5322) );
  XNOR U7414 ( .A(n5318), .B(n5319), .Z(n5317) );
  XNOR U7415 ( .A(y[1357]), .B(x[1357]), .Z(n5319) );
  XNOR U7416 ( .A(y[1358]), .B(x[1358]), .Z(n5318) );
  XNOR U7417 ( .A(y[1356]), .B(x[1356]), .Z(n5316) );
  XNOR U7418 ( .A(n5310), .B(n5311), .Z(n5321) );
  XNOR U7419 ( .A(y[1353]), .B(x[1353]), .Z(n5311) );
  XNOR U7420 ( .A(n5312), .B(n5313), .Z(n5310) );
  XNOR U7421 ( .A(y[1354]), .B(x[1354]), .Z(n5313) );
  XNOR U7422 ( .A(y[1355]), .B(x[1355]), .Z(n5312) );
  XNOR U7423 ( .A(n5303), .B(n5302), .Z(n5306) );
  XNOR U7424 ( .A(n5298), .B(n5299), .Z(n5302) );
  XNOR U7425 ( .A(y[1350]), .B(x[1350]), .Z(n5299) );
  XNOR U7426 ( .A(n5300), .B(n5301), .Z(n5298) );
  XNOR U7427 ( .A(y[1351]), .B(x[1351]), .Z(n5301) );
  XNOR U7428 ( .A(y[1352]), .B(x[1352]), .Z(n5300) );
  XNOR U7429 ( .A(n5292), .B(n5293), .Z(n5303) );
  XNOR U7430 ( .A(y[1347]), .B(x[1347]), .Z(n5293) );
  XNOR U7431 ( .A(n5294), .B(n5295), .Z(n5292) );
  XNOR U7432 ( .A(y[1348]), .B(x[1348]), .Z(n5295) );
  XNOR U7433 ( .A(y[1349]), .B(x[1349]), .Z(n5294) );
  XOR U7434 ( .A(n5268), .B(n5269), .Z(n5287) );
  XNOR U7435 ( .A(n5284), .B(n5285), .Z(n5269) );
  XNOR U7436 ( .A(n5279), .B(n5280), .Z(n5285) );
  XNOR U7437 ( .A(n5281), .B(n5282), .Z(n5280) );
  XNOR U7438 ( .A(y[1345]), .B(x[1345]), .Z(n5282) );
  XNOR U7439 ( .A(y[1346]), .B(x[1346]), .Z(n5281) );
  XNOR U7440 ( .A(y[1344]), .B(x[1344]), .Z(n5279) );
  XNOR U7441 ( .A(n5273), .B(n5274), .Z(n5284) );
  XNOR U7442 ( .A(y[1341]), .B(x[1341]), .Z(n5274) );
  XNOR U7443 ( .A(n5275), .B(n5276), .Z(n5273) );
  XNOR U7444 ( .A(y[1342]), .B(x[1342]), .Z(n5276) );
  XNOR U7445 ( .A(y[1343]), .B(x[1343]), .Z(n5275) );
  XOR U7446 ( .A(n5267), .B(n5266), .Z(n5268) );
  XNOR U7447 ( .A(n5262), .B(n5263), .Z(n5266) );
  XNOR U7448 ( .A(y[1338]), .B(x[1338]), .Z(n5263) );
  XNOR U7449 ( .A(n5264), .B(n5265), .Z(n5262) );
  XNOR U7450 ( .A(y[1339]), .B(x[1339]), .Z(n5265) );
  XNOR U7451 ( .A(y[1340]), .B(x[1340]), .Z(n5264) );
  XNOR U7452 ( .A(n5256), .B(n5257), .Z(n5267) );
  XNOR U7453 ( .A(y[1335]), .B(x[1335]), .Z(n5257) );
  XNOR U7454 ( .A(n5258), .B(n5259), .Z(n5256) );
  XNOR U7455 ( .A(y[1336]), .B(x[1336]), .Z(n5259) );
  XNOR U7456 ( .A(y[1337]), .B(x[1337]), .Z(n5258) );
  NAND U7457 ( .A(n5323), .B(n5324), .Z(N13390) );
  NANDN U7458 ( .A(n5325), .B(n5326), .Z(n5324) );
  OR U7459 ( .A(n5327), .B(n5328), .Z(n5326) );
  NAND U7460 ( .A(n5327), .B(n5328), .Z(n5323) );
  XOR U7461 ( .A(n5327), .B(n5329), .Z(N13389) );
  XNOR U7462 ( .A(n5325), .B(n5328), .Z(n5329) );
  AND U7463 ( .A(n5330), .B(n5331), .Z(n5328) );
  NANDN U7464 ( .A(n5332), .B(n5333), .Z(n5331) );
  NANDN U7465 ( .A(n5334), .B(n5335), .Z(n5333) );
  NANDN U7466 ( .A(n5335), .B(n5334), .Z(n5330) );
  NAND U7467 ( .A(n5336), .B(n5337), .Z(n5325) );
  NANDN U7468 ( .A(n5338), .B(n5339), .Z(n5337) );
  OR U7469 ( .A(n5340), .B(n5341), .Z(n5339) );
  NAND U7470 ( .A(n5341), .B(n5340), .Z(n5336) );
  AND U7471 ( .A(n5342), .B(n5343), .Z(n5327) );
  NANDN U7472 ( .A(n5344), .B(n5345), .Z(n5343) );
  NANDN U7473 ( .A(n5346), .B(n5347), .Z(n5345) );
  NANDN U7474 ( .A(n5347), .B(n5346), .Z(n5342) );
  XOR U7475 ( .A(n5341), .B(n5348), .Z(N13388) );
  XOR U7476 ( .A(n5338), .B(n5340), .Z(n5348) );
  XNOR U7477 ( .A(n5334), .B(n5349), .Z(n5340) );
  XNOR U7478 ( .A(n5332), .B(n5335), .Z(n5349) );
  NAND U7479 ( .A(n5350), .B(n5351), .Z(n5335) );
  NAND U7480 ( .A(n5352), .B(n5353), .Z(n5351) );
  OR U7481 ( .A(n5354), .B(n5355), .Z(n5352) );
  NANDN U7482 ( .A(n5356), .B(n5354), .Z(n5350) );
  IV U7483 ( .A(n5355), .Z(n5356) );
  NAND U7484 ( .A(n5357), .B(n5358), .Z(n5332) );
  NAND U7485 ( .A(n5359), .B(n5360), .Z(n5358) );
  NANDN U7486 ( .A(n5361), .B(n5362), .Z(n5359) );
  NANDN U7487 ( .A(n5362), .B(n5361), .Z(n5357) );
  AND U7488 ( .A(n5363), .B(n5364), .Z(n5334) );
  NAND U7489 ( .A(n5365), .B(n5366), .Z(n5364) );
  OR U7490 ( .A(n5367), .B(n5368), .Z(n5365) );
  NANDN U7491 ( .A(n5369), .B(n5367), .Z(n5363) );
  NAND U7492 ( .A(n5370), .B(n5371), .Z(n5338) );
  NANDN U7493 ( .A(n5372), .B(n5373), .Z(n5371) );
  OR U7494 ( .A(n5374), .B(n5375), .Z(n5373) );
  NANDN U7495 ( .A(n5376), .B(n5374), .Z(n5370) );
  IV U7496 ( .A(n5375), .Z(n5376) );
  XNOR U7497 ( .A(n5346), .B(n5377), .Z(n5341) );
  XNOR U7498 ( .A(n5344), .B(n5347), .Z(n5377) );
  NAND U7499 ( .A(n5378), .B(n5379), .Z(n5347) );
  NAND U7500 ( .A(n5380), .B(n5381), .Z(n5379) );
  OR U7501 ( .A(n5382), .B(n5383), .Z(n5380) );
  NANDN U7502 ( .A(n5384), .B(n5382), .Z(n5378) );
  IV U7503 ( .A(n5383), .Z(n5384) );
  NAND U7504 ( .A(n5385), .B(n5386), .Z(n5344) );
  NAND U7505 ( .A(n5387), .B(n5388), .Z(n5386) );
  NANDN U7506 ( .A(n5389), .B(n5390), .Z(n5387) );
  NANDN U7507 ( .A(n5390), .B(n5389), .Z(n5385) );
  AND U7508 ( .A(n5391), .B(n5392), .Z(n5346) );
  NAND U7509 ( .A(n5393), .B(n5394), .Z(n5392) );
  OR U7510 ( .A(n5395), .B(n5396), .Z(n5393) );
  NANDN U7511 ( .A(n5397), .B(n5395), .Z(n5391) );
  XNOR U7512 ( .A(n5372), .B(n5398), .Z(N13387) );
  XOR U7513 ( .A(n5374), .B(n5375), .Z(n5398) );
  XNOR U7514 ( .A(n5388), .B(n5399), .Z(n5375) );
  XOR U7515 ( .A(n5389), .B(n5390), .Z(n5399) );
  XOR U7516 ( .A(n5395), .B(n5400), .Z(n5390) );
  XOR U7517 ( .A(n5394), .B(n5397), .Z(n5400) );
  IV U7518 ( .A(n5396), .Z(n5397) );
  NAND U7519 ( .A(n5401), .B(n5402), .Z(n5396) );
  OR U7520 ( .A(n5403), .B(n5404), .Z(n5402) );
  OR U7521 ( .A(n5405), .B(n5406), .Z(n5401) );
  NAND U7522 ( .A(n5407), .B(n5408), .Z(n5394) );
  OR U7523 ( .A(n5409), .B(n5410), .Z(n5408) );
  OR U7524 ( .A(n5411), .B(n5412), .Z(n5407) );
  NOR U7525 ( .A(n5413), .B(n5414), .Z(n5395) );
  ANDN U7526 ( .B(n5415), .A(n5416), .Z(n5389) );
  XNOR U7527 ( .A(n5382), .B(n5417), .Z(n5388) );
  XNOR U7528 ( .A(n5381), .B(n5383), .Z(n5417) );
  NAND U7529 ( .A(n5418), .B(n5419), .Z(n5383) );
  OR U7530 ( .A(n5420), .B(n5421), .Z(n5419) );
  OR U7531 ( .A(n5422), .B(n5423), .Z(n5418) );
  NAND U7532 ( .A(n5424), .B(n5425), .Z(n5381) );
  OR U7533 ( .A(n5426), .B(n5427), .Z(n5425) );
  OR U7534 ( .A(n5428), .B(n5429), .Z(n5424) );
  ANDN U7535 ( .B(n5430), .A(n5431), .Z(n5382) );
  IV U7536 ( .A(n5432), .Z(n5430) );
  ANDN U7537 ( .B(n5433), .A(n5434), .Z(n5374) );
  XOR U7538 ( .A(n5360), .B(n5435), .Z(n5372) );
  XOR U7539 ( .A(n5361), .B(n5362), .Z(n5435) );
  XOR U7540 ( .A(n5367), .B(n5436), .Z(n5362) );
  XOR U7541 ( .A(n5366), .B(n5369), .Z(n5436) );
  IV U7542 ( .A(n5368), .Z(n5369) );
  NAND U7543 ( .A(n5437), .B(n5438), .Z(n5368) );
  OR U7544 ( .A(n5439), .B(n5440), .Z(n5438) );
  OR U7545 ( .A(n5441), .B(n5442), .Z(n5437) );
  NAND U7546 ( .A(n5443), .B(n5444), .Z(n5366) );
  OR U7547 ( .A(n5445), .B(n5446), .Z(n5444) );
  OR U7548 ( .A(n5447), .B(n5448), .Z(n5443) );
  NOR U7549 ( .A(n5449), .B(n5450), .Z(n5367) );
  ANDN U7550 ( .B(n5451), .A(n5452), .Z(n5361) );
  IV U7551 ( .A(n5453), .Z(n5451) );
  XNOR U7552 ( .A(n5354), .B(n5454), .Z(n5360) );
  XNOR U7553 ( .A(n5353), .B(n5355), .Z(n5454) );
  NAND U7554 ( .A(n5455), .B(n5456), .Z(n5355) );
  OR U7555 ( .A(n5457), .B(n5458), .Z(n5456) );
  OR U7556 ( .A(n5459), .B(n5460), .Z(n5455) );
  NAND U7557 ( .A(n5461), .B(n5462), .Z(n5353) );
  OR U7558 ( .A(n5463), .B(n5464), .Z(n5462) );
  OR U7559 ( .A(n5465), .B(n5466), .Z(n5461) );
  ANDN U7560 ( .B(n5467), .A(n5468), .Z(n5354) );
  IV U7561 ( .A(n5469), .Z(n5467) );
  XNOR U7562 ( .A(n5434), .B(n5433), .Z(N13386) );
  XOR U7563 ( .A(n5453), .B(n5452), .Z(n5433) );
  XNOR U7564 ( .A(n5468), .B(n5469), .Z(n5452) );
  XNOR U7565 ( .A(n5463), .B(n5464), .Z(n5469) );
  XNOR U7566 ( .A(n5465), .B(n5466), .Z(n5464) );
  XNOR U7567 ( .A(y[1333]), .B(x[1333]), .Z(n5466) );
  XNOR U7568 ( .A(y[1334]), .B(x[1334]), .Z(n5465) );
  XNOR U7569 ( .A(y[1332]), .B(x[1332]), .Z(n5463) );
  XNOR U7570 ( .A(n5457), .B(n5458), .Z(n5468) );
  XNOR U7571 ( .A(y[1329]), .B(x[1329]), .Z(n5458) );
  XNOR U7572 ( .A(n5459), .B(n5460), .Z(n5457) );
  XNOR U7573 ( .A(y[1330]), .B(x[1330]), .Z(n5460) );
  XNOR U7574 ( .A(y[1331]), .B(x[1331]), .Z(n5459) );
  XNOR U7575 ( .A(n5450), .B(n5449), .Z(n5453) );
  XNOR U7576 ( .A(n5445), .B(n5446), .Z(n5449) );
  XNOR U7577 ( .A(y[1326]), .B(x[1326]), .Z(n5446) );
  XNOR U7578 ( .A(n5447), .B(n5448), .Z(n5445) );
  XNOR U7579 ( .A(y[1327]), .B(x[1327]), .Z(n5448) );
  XNOR U7580 ( .A(y[1328]), .B(x[1328]), .Z(n5447) );
  XNOR U7581 ( .A(n5439), .B(n5440), .Z(n5450) );
  XNOR U7582 ( .A(y[1323]), .B(x[1323]), .Z(n5440) );
  XNOR U7583 ( .A(n5441), .B(n5442), .Z(n5439) );
  XNOR U7584 ( .A(y[1324]), .B(x[1324]), .Z(n5442) );
  XNOR U7585 ( .A(y[1325]), .B(x[1325]), .Z(n5441) );
  XOR U7586 ( .A(n5415), .B(n5416), .Z(n5434) );
  XNOR U7587 ( .A(n5431), .B(n5432), .Z(n5416) );
  XNOR U7588 ( .A(n5426), .B(n5427), .Z(n5432) );
  XNOR U7589 ( .A(n5428), .B(n5429), .Z(n5427) );
  XNOR U7590 ( .A(y[1321]), .B(x[1321]), .Z(n5429) );
  XNOR U7591 ( .A(y[1322]), .B(x[1322]), .Z(n5428) );
  XNOR U7592 ( .A(y[1320]), .B(x[1320]), .Z(n5426) );
  XNOR U7593 ( .A(n5420), .B(n5421), .Z(n5431) );
  XNOR U7594 ( .A(y[1317]), .B(x[1317]), .Z(n5421) );
  XNOR U7595 ( .A(n5422), .B(n5423), .Z(n5420) );
  XNOR U7596 ( .A(y[1318]), .B(x[1318]), .Z(n5423) );
  XNOR U7597 ( .A(y[1319]), .B(x[1319]), .Z(n5422) );
  XOR U7598 ( .A(n5414), .B(n5413), .Z(n5415) );
  XNOR U7599 ( .A(n5409), .B(n5410), .Z(n5413) );
  XNOR U7600 ( .A(y[1314]), .B(x[1314]), .Z(n5410) );
  XNOR U7601 ( .A(n5411), .B(n5412), .Z(n5409) );
  XNOR U7602 ( .A(y[1315]), .B(x[1315]), .Z(n5412) );
  XNOR U7603 ( .A(y[1316]), .B(x[1316]), .Z(n5411) );
  XNOR U7604 ( .A(n5403), .B(n5404), .Z(n5414) );
  XNOR U7605 ( .A(y[1311]), .B(x[1311]), .Z(n5404) );
  XNOR U7606 ( .A(n5405), .B(n5406), .Z(n5403) );
  XNOR U7607 ( .A(y[1312]), .B(x[1312]), .Z(n5406) );
  XNOR U7608 ( .A(y[1313]), .B(x[1313]), .Z(n5405) );
  NAND U7609 ( .A(n5470), .B(n5471), .Z(N13379) );
  NANDN U7610 ( .A(n5472), .B(n5473), .Z(n5471) );
  OR U7611 ( .A(n5474), .B(n5475), .Z(n5473) );
  NAND U7612 ( .A(n5474), .B(n5475), .Z(n5470) );
  XOR U7613 ( .A(n5474), .B(n5476), .Z(N13378) );
  XNOR U7614 ( .A(n5472), .B(n5475), .Z(n5476) );
  AND U7615 ( .A(n5477), .B(n5478), .Z(n5475) );
  NANDN U7616 ( .A(n5479), .B(n5480), .Z(n5478) );
  NANDN U7617 ( .A(n5481), .B(n5482), .Z(n5480) );
  NANDN U7618 ( .A(n5482), .B(n5481), .Z(n5477) );
  NAND U7619 ( .A(n5483), .B(n5484), .Z(n5472) );
  NANDN U7620 ( .A(n5485), .B(n5486), .Z(n5484) );
  OR U7621 ( .A(n5487), .B(n5488), .Z(n5486) );
  NAND U7622 ( .A(n5488), .B(n5487), .Z(n5483) );
  AND U7623 ( .A(n5489), .B(n5490), .Z(n5474) );
  NANDN U7624 ( .A(n5491), .B(n5492), .Z(n5490) );
  NANDN U7625 ( .A(n5493), .B(n5494), .Z(n5492) );
  NANDN U7626 ( .A(n5494), .B(n5493), .Z(n5489) );
  XOR U7627 ( .A(n5488), .B(n5495), .Z(N13377) );
  XOR U7628 ( .A(n5485), .B(n5487), .Z(n5495) );
  XNOR U7629 ( .A(n5481), .B(n5496), .Z(n5487) );
  XNOR U7630 ( .A(n5479), .B(n5482), .Z(n5496) );
  NAND U7631 ( .A(n5497), .B(n5498), .Z(n5482) );
  NAND U7632 ( .A(n5499), .B(n5500), .Z(n5498) );
  OR U7633 ( .A(n5501), .B(n5502), .Z(n5499) );
  NANDN U7634 ( .A(n5503), .B(n5501), .Z(n5497) );
  IV U7635 ( .A(n5502), .Z(n5503) );
  NAND U7636 ( .A(n5504), .B(n5505), .Z(n5479) );
  NAND U7637 ( .A(n5506), .B(n5507), .Z(n5505) );
  NANDN U7638 ( .A(n5508), .B(n5509), .Z(n5506) );
  NANDN U7639 ( .A(n5509), .B(n5508), .Z(n5504) );
  AND U7640 ( .A(n5510), .B(n5511), .Z(n5481) );
  NAND U7641 ( .A(n5512), .B(n5513), .Z(n5511) );
  OR U7642 ( .A(n5514), .B(n5515), .Z(n5512) );
  NANDN U7643 ( .A(n5516), .B(n5514), .Z(n5510) );
  NAND U7644 ( .A(n5517), .B(n5518), .Z(n5485) );
  NANDN U7645 ( .A(n5519), .B(n5520), .Z(n5518) );
  OR U7646 ( .A(n5521), .B(n5522), .Z(n5520) );
  NANDN U7647 ( .A(n5523), .B(n5521), .Z(n5517) );
  IV U7648 ( .A(n5522), .Z(n5523) );
  XNOR U7649 ( .A(n5493), .B(n5524), .Z(n5488) );
  XNOR U7650 ( .A(n5491), .B(n5494), .Z(n5524) );
  NAND U7651 ( .A(n5525), .B(n5526), .Z(n5494) );
  NAND U7652 ( .A(n5527), .B(n5528), .Z(n5526) );
  OR U7653 ( .A(n5529), .B(n5530), .Z(n5527) );
  NANDN U7654 ( .A(n5531), .B(n5529), .Z(n5525) );
  IV U7655 ( .A(n5530), .Z(n5531) );
  NAND U7656 ( .A(n5532), .B(n5533), .Z(n5491) );
  NAND U7657 ( .A(n5534), .B(n5535), .Z(n5533) );
  NANDN U7658 ( .A(n5536), .B(n5537), .Z(n5534) );
  NANDN U7659 ( .A(n5537), .B(n5536), .Z(n5532) );
  AND U7660 ( .A(n5538), .B(n5539), .Z(n5493) );
  NAND U7661 ( .A(n5540), .B(n5541), .Z(n5539) );
  OR U7662 ( .A(n5542), .B(n5543), .Z(n5540) );
  NANDN U7663 ( .A(n5544), .B(n5542), .Z(n5538) );
  XNOR U7664 ( .A(n5519), .B(n5545), .Z(N13376) );
  XOR U7665 ( .A(n5521), .B(n5522), .Z(n5545) );
  XNOR U7666 ( .A(n5535), .B(n5546), .Z(n5522) );
  XOR U7667 ( .A(n5536), .B(n5537), .Z(n5546) );
  XOR U7668 ( .A(n5542), .B(n5547), .Z(n5537) );
  XOR U7669 ( .A(n5541), .B(n5544), .Z(n5547) );
  IV U7670 ( .A(n5543), .Z(n5544) );
  NAND U7671 ( .A(n5548), .B(n5549), .Z(n5543) );
  OR U7672 ( .A(n5550), .B(n5551), .Z(n5549) );
  OR U7673 ( .A(n5552), .B(n5553), .Z(n5548) );
  NAND U7674 ( .A(n5554), .B(n5555), .Z(n5541) );
  OR U7675 ( .A(n5556), .B(n5557), .Z(n5555) );
  OR U7676 ( .A(n5558), .B(n5559), .Z(n5554) );
  NOR U7677 ( .A(n5560), .B(n5561), .Z(n5542) );
  ANDN U7678 ( .B(n5562), .A(n5563), .Z(n5536) );
  XNOR U7679 ( .A(n5529), .B(n5564), .Z(n5535) );
  XNOR U7680 ( .A(n5528), .B(n5530), .Z(n5564) );
  NAND U7681 ( .A(n5565), .B(n5566), .Z(n5530) );
  OR U7682 ( .A(n5567), .B(n5568), .Z(n5566) );
  OR U7683 ( .A(n5569), .B(n5570), .Z(n5565) );
  NAND U7684 ( .A(n5571), .B(n5572), .Z(n5528) );
  OR U7685 ( .A(n5573), .B(n5574), .Z(n5572) );
  OR U7686 ( .A(n5575), .B(n5576), .Z(n5571) );
  ANDN U7687 ( .B(n5577), .A(n5578), .Z(n5529) );
  IV U7688 ( .A(n5579), .Z(n5577) );
  ANDN U7689 ( .B(n5580), .A(n5581), .Z(n5521) );
  XOR U7690 ( .A(n5507), .B(n5582), .Z(n5519) );
  XOR U7691 ( .A(n5508), .B(n5509), .Z(n5582) );
  XOR U7692 ( .A(n5514), .B(n5583), .Z(n5509) );
  XOR U7693 ( .A(n5513), .B(n5516), .Z(n5583) );
  IV U7694 ( .A(n5515), .Z(n5516) );
  NAND U7695 ( .A(n5584), .B(n5585), .Z(n5515) );
  OR U7696 ( .A(n5586), .B(n5587), .Z(n5585) );
  OR U7697 ( .A(n5588), .B(n5589), .Z(n5584) );
  NAND U7698 ( .A(n5590), .B(n5591), .Z(n5513) );
  OR U7699 ( .A(n5592), .B(n5593), .Z(n5591) );
  OR U7700 ( .A(n5594), .B(n5595), .Z(n5590) );
  NOR U7701 ( .A(n5596), .B(n5597), .Z(n5514) );
  ANDN U7702 ( .B(n5598), .A(n5599), .Z(n5508) );
  IV U7703 ( .A(n5600), .Z(n5598) );
  XNOR U7704 ( .A(n5501), .B(n5601), .Z(n5507) );
  XNOR U7705 ( .A(n5500), .B(n5502), .Z(n5601) );
  NAND U7706 ( .A(n5602), .B(n5603), .Z(n5502) );
  OR U7707 ( .A(n5604), .B(n5605), .Z(n5603) );
  OR U7708 ( .A(n5606), .B(n5607), .Z(n5602) );
  NAND U7709 ( .A(n5608), .B(n5609), .Z(n5500) );
  OR U7710 ( .A(n5610), .B(n5611), .Z(n5609) );
  OR U7711 ( .A(n5612), .B(n5613), .Z(n5608) );
  ANDN U7712 ( .B(n5614), .A(n5615), .Z(n5501) );
  IV U7713 ( .A(n5616), .Z(n5614) );
  XNOR U7714 ( .A(n5581), .B(n5580), .Z(N13375) );
  XOR U7715 ( .A(n5600), .B(n5599), .Z(n5580) );
  XNOR U7716 ( .A(n5615), .B(n5616), .Z(n5599) );
  XNOR U7717 ( .A(n5610), .B(n5611), .Z(n5616) );
  XNOR U7718 ( .A(n5612), .B(n5613), .Z(n5611) );
  XNOR U7719 ( .A(y[1309]), .B(x[1309]), .Z(n5613) );
  XNOR U7720 ( .A(y[1310]), .B(x[1310]), .Z(n5612) );
  XNOR U7721 ( .A(y[1308]), .B(x[1308]), .Z(n5610) );
  XNOR U7722 ( .A(n5604), .B(n5605), .Z(n5615) );
  XNOR U7723 ( .A(y[1305]), .B(x[1305]), .Z(n5605) );
  XNOR U7724 ( .A(n5606), .B(n5607), .Z(n5604) );
  XNOR U7725 ( .A(y[1306]), .B(x[1306]), .Z(n5607) );
  XNOR U7726 ( .A(y[1307]), .B(x[1307]), .Z(n5606) );
  XNOR U7727 ( .A(n5597), .B(n5596), .Z(n5600) );
  XNOR U7728 ( .A(n5592), .B(n5593), .Z(n5596) );
  XNOR U7729 ( .A(y[1302]), .B(x[1302]), .Z(n5593) );
  XNOR U7730 ( .A(n5594), .B(n5595), .Z(n5592) );
  XNOR U7731 ( .A(y[1303]), .B(x[1303]), .Z(n5595) );
  XNOR U7732 ( .A(y[1304]), .B(x[1304]), .Z(n5594) );
  XNOR U7733 ( .A(n5586), .B(n5587), .Z(n5597) );
  XNOR U7734 ( .A(y[1299]), .B(x[1299]), .Z(n5587) );
  XNOR U7735 ( .A(n5588), .B(n5589), .Z(n5586) );
  XNOR U7736 ( .A(y[1300]), .B(x[1300]), .Z(n5589) );
  XNOR U7737 ( .A(y[1301]), .B(x[1301]), .Z(n5588) );
  XOR U7738 ( .A(n5562), .B(n5563), .Z(n5581) );
  XNOR U7739 ( .A(n5578), .B(n5579), .Z(n5563) );
  XNOR U7740 ( .A(n5573), .B(n5574), .Z(n5579) );
  XNOR U7741 ( .A(n5575), .B(n5576), .Z(n5574) );
  XNOR U7742 ( .A(y[1297]), .B(x[1297]), .Z(n5576) );
  XNOR U7743 ( .A(y[1298]), .B(x[1298]), .Z(n5575) );
  XNOR U7744 ( .A(y[1296]), .B(x[1296]), .Z(n5573) );
  XNOR U7745 ( .A(n5567), .B(n5568), .Z(n5578) );
  XNOR U7746 ( .A(y[1293]), .B(x[1293]), .Z(n5568) );
  XNOR U7747 ( .A(n5569), .B(n5570), .Z(n5567) );
  XNOR U7748 ( .A(y[1294]), .B(x[1294]), .Z(n5570) );
  XNOR U7749 ( .A(y[1295]), .B(x[1295]), .Z(n5569) );
  XOR U7750 ( .A(n5561), .B(n5560), .Z(n5562) );
  XNOR U7751 ( .A(n5556), .B(n5557), .Z(n5560) );
  XNOR U7752 ( .A(y[1290]), .B(x[1290]), .Z(n5557) );
  XNOR U7753 ( .A(n5558), .B(n5559), .Z(n5556) );
  XNOR U7754 ( .A(y[1291]), .B(x[1291]), .Z(n5559) );
  XNOR U7755 ( .A(y[1292]), .B(x[1292]), .Z(n5558) );
  XNOR U7756 ( .A(n5550), .B(n5551), .Z(n5561) );
  XNOR U7757 ( .A(y[1287]), .B(x[1287]), .Z(n5551) );
  XNOR U7758 ( .A(n5552), .B(n5553), .Z(n5550) );
  XNOR U7759 ( .A(y[1288]), .B(x[1288]), .Z(n5553) );
  XNOR U7760 ( .A(y[1289]), .B(x[1289]), .Z(n5552) );
  NAND U7761 ( .A(n5617), .B(n5618), .Z(N13368) );
  NANDN U7762 ( .A(n5619), .B(n5620), .Z(n5618) );
  OR U7763 ( .A(n5621), .B(n5622), .Z(n5620) );
  NAND U7764 ( .A(n5621), .B(n5622), .Z(n5617) );
  XOR U7765 ( .A(n5621), .B(n5623), .Z(N13367) );
  XNOR U7766 ( .A(n5619), .B(n5622), .Z(n5623) );
  AND U7767 ( .A(n5624), .B(n5625), .Z(n5622) );
  NANDN U7768 ( .A(n5626), .B(n5627), .Z(n5625) );
  NANDN U7769 ( .A(n5628), .B(n5629), .Z(n5627) );
  NANDN U7770 ( .A(n5629), .B(n5628), .Z(n5624) );
  NAND U7771 ( .A(n5630), .B(n5631), .Z(n5619) );
  NANDN U7772 ( .A(n5632), .B(n5633), .Z(n5631) );
  OR U7773 ( .A(n5634), .B(n5635), .Z(n5633) );
  NAND U7774 ( .A(n5635), .B(n5634), .Z(n5630) );
  AND U7775 ( .A(n5636), .B(n5637), .Z(n5621) );
  NANDN U7776 ( .A(n5638), .B(n5639), .Z(n5637) );
  NANDN U7777 ( .A(n5640), .B(n5641), .Z(n5639) );
  NANDN U7778 ( .A(n5641), .B(n5640), .Z(n5636) );
  XOR U7779 ( .A(n5635), .B(n5642), .Z(N13366) );
  XOR U7780 ( .A(n5632), .B(n5634), .Z(n5642) );
  XNOR U7781 ( .A(n5628), .B(n5643), .Z(n5634) );
  XNOR U7782 ( .A(n5626), .B(n5629), .Z(n5643) );
  NAND U7783 ( .A(n5644), .B(n5645), .Z(n5629) );
  NAND U7784 ( .A(n5646), .B(n5647), .Z(n5645) );
  OR U7785 ( .A(n5648), .B(n5649), .Z(n5646) );
  NANDN U7786 ( .A(n5650), .B(n5648), .Z(n5644) );
  IV U7787 ( .A(n5649), .Z(n5650) );
  NAND U7788 ( .A(n5651), .B(n5652), .Z(n5626) );
  NAND U7789 ( .A(n5653), .B(n5654), .Z(n5652) );
  NANDN U7790 ( .A(n5655), .B(n5656), .Z(n5653) );
  NANDN U7791 ( .A(n5656), .B(n5655), .Z(n5651) );
  AND U7792 ( .A(n5657), .B(n5658), .Z(n5628) );
  NAND U7793 ( .A(n5659), .B(n5660), .Z(n5658) );
  OR U7794 ( .A(n5661), .B(n5662), .Z(n5659) );
  NANDN U7795 ( .A(n5663), .B(n5661), .Z(n5657) );
  NAND U7796 ( .A(n5664), .B(n5665), .Z(n5632) );
  NANDN U7797 ( .A(n5666), .B(n5667), .Z(n5665) );
  OR U7798 ( .A(n5668), .B(n5669), .Z(n5667) );
  NANDN U7799 ( .A(n5670), .B(n5668), .Z(n5664) );
  IV U7800 ( .A(n5669), .Z(n5670) );
  XNOR U7801 ( .A(n5640), .B(n5671), .Z(n5635) );
  XNOR U7802 ( .A(n5638), .B(n5641), .Z(n5671) );
  NAND U7803 ( .A(n5672), .B(n5673), .Z(n5641) );
  NAND U7804 ( .A(n5674), .B(n5675), .Z(n5673) );
  OR U7805 ( .A(n5676), .B(n5677), .Z(n5674) );
  NANDN U7806 ( .A(n5678), .B(n5676), .Z(n5672) );
  IV U7807 ( .A(n5677), .Z(n5678) );
  NAND U7808 ( .A(n5679), .B(n5680), .Z(n5638) );
  NAND U7809 ( .A(n5681), .B(n5682), .Z(n5680) );
  NANDN U7810 ( .A(n5683), .B(n5684), .Z(n5681) );
  NANDN U7811 ( .A(n5684), .B(n5683), .Z(n5679) );
  AND U7812 ( .A(n5685), .B(n5686), .Z(n5640) );
  NAND U7813 ( .A(n5687), .B(n5688), .Z(n5686) );
  OR U7814 ( .A(n5689), .B(n5690), .Z(n5687) );
  NANDN U7815 ( .A(n5691), .B(n5689), .Z(n5685) );
  XNOR U7816 ( .A(n5666), .B(n5692), .Z(N13365) );
  XOR U7817 ( .A(n5668), .B(n5669), .Z(n5692) );
  XNOR U7818 ( .A(n5682), .B(n5693), .Z(n5669) );
  XOR U7819 ( .A(n5683), .B(n5684), .Z(n5693) );
  XOR U7820 ( .A(n5689), .B(n5694), .Z(n5684) );
  XOR U7821 ( .A(n5688), .B(n5691), .Z(n5694) );
  IV U7822 ( .A(n5690), .Z(n5691) );
  NAND U7823 ( .A(n5695), .B(n5696), .Z(n5690) );
  OR U7824 ( .A(n5697), .B(n5698), .Z(n5696) );
  OR U7825 ( .A(n5699), .B(n5700), .Z(n5695) );
  NAND U7826 ( .A(n5701), .B(n5702), .Z(n5688) );
  OR U7827 ( .A(n5703), .B(n5704), .Z(n5702) );
  OR U7828 ( .A(n5705), .B(n5706), .Z(n5701) );
  NOR U7829 ( .A(n5707), .B(n5708), .Z(n5689) );
  ANDN U7830 ( .B(n5709), .A(n5710), .Z(n5683) );
  XNOR U7831 ( .A(n5676), .B(n5711), .Z(n5682) );
  XNOR U7832 ( .A(n5675), .B(n5677), .Z(n5711) );
  NAND U7833 ( .A(n5712), .B(n5713), .Z(n5677) );
  OR U7834 ( .A(n5714), .B(n5715), .Z(n5713) );
  OR U7835 ( .A(n5716), .B(n5717), .Z(n5712) );
  NAND U7836 ( .A(n5718), .B(n5719), .Z(n5675) );
  OR U7837 ( .A(n5720), .B(n5721), .Z(n5719) );
  OR U7838 ( .A(n5722), .B(n5723), .Z(n5718) );
  ANDN U7839 ( .B(n5724), .A(n5725), .Z(n5676) );
  IV U7840 ( .A(n5726), .Z(n5724) );
  ANDN U7841 ( .B(n5727), .A(n5728), .Z(n5668) );
  XOR U7842 ( .A(n5654), .B(n5729), .Z(n5666) );
  XOR U7843 ( .A(n5655), .B(n5656), .Z(n5729) );
  XOR U7844 ( .A(n5661), .B(n5730), .Z(n5656) );
  XOR U7845 ( .A(n5660), .B(n5663), .Z(n5730) );
  IV U7846 ( .A(n5662), .Z(n5663) );
  NAND U7847 ( .A(n5731), .B(n5732), .Z(n5662) );
  OR U7848 ( .A(n5733), .B(n5734), .Z(n5732) );
  OR U7849 ( .A(n5735), .B(n5736), .Z(n5731) );
  NAND U7850 ( .A(n5737), .B(n5738), .Z(n5660) );
  OR U7851 ( .A(n5739), .B(n5740), .Z(n5738) );
  OR U7852 ( .A(n5741), .B(n5742), .Z(n5737) );
  NOR U7853 ( .A(n5743), .B(n5744), .Z(n5661) );
  ANDN U7854 ( .B(n5745), .A(n5746), .Z(n5655) );
  IV U7855 ( .A(n5747), .Z(n5745) );
  XNOR U7856 ( .A(n5648), .B(n5748), .Z(n5654) );
  XNOR U7857 ( .A(n5647), .B(n5649), .Z(n5748) );
  NAND U7858 ( .A(n5749), .B(n5750), .Z(n5649) );
  OR U7859 ( .A(n5751), .B(n5752), .Z(n5750) );
  OR U7860 ( .A(n5753), .B(n5754), .Z(n5749) );
  NAND U7861 ( .A(n5755), .B(n5756), .Z(n5647) );
  OR U7862 ( .A(n5757), .B(n5758), .Z(n5756) );
  OR U7863 ( .A(n5759), .B(n5760), .Z(n5755) );
  ANDN U7864 ( .B(n5761), .A(n5762), .Z(n5648) );
  IV U7865 ( .A(n5763), .Z(n5761) );
  XNOR U7866 ( .A(n5728), .B(n5727), .Z(N13364) );
  XOR U7867 ( .A(n5747), .B(n5746), .Z(n5727) );
  XNOR U7868 ( .A(n5762), .B(n5763), .Z(n5746) );
  XNOR U7869 ( .A(n5757), .B(n5758), .Z(n5763) );
  XNOR U7870 ( .A(n5759), .B(n5760), .Z(n5758) );
  XNOR U7871 ( .A(y[1285]), .B(x[1285]), .Z(n5760) );
  XNOR U7872 ( .A(y[1286]), .B(x[1286]), .Z(n5759) );
  XNOR U7873 ( .A(y[1284]), .B(x[1284]), .Z(n5757) );
  XNOR U7874 ( .A(n5751), .B(n5752), .Z(n5762) );
  XNOR U7875 ( .A(y[1281]), .B(x[1281]), .Z(n5752) );
  XNOR U7876 ( .A(n5753), .B(n5754), .Z(n5751) );
  XNOR U7877 ( .A(y[1282]), .B(x[1282]), .Z(n5754) );
  XNOR U7878 ( .A(y[1283]), .B(x[1283]), .Z(n5753) );
  XNOR U7879 ( .A(n5744), .B(n5743), .Z(n5747) );
  XNOR U7880 ( .A(n5739), .B(n5740), .Z(n5743) );
  XNOR U7881 ( .A(y[1278]), .B(x[1278]), .Z(n5740) );
  XNOR U7882 ( .A(n5741), .B(n5742), .Z(n5739) );
  XNOR U7883 ( .A(y[1279]), .B(x[1279]), .Z(n5742) );
  XNOR U7884 ( .A(y[1280]), .B(x[1280]), .Z(n5741) );
  XNOR U7885 ( .A(n5733), .B(n5734), .Z(n5744) );
  XNOR U7886 ( .A(y[1275]), .B(x[1275]), .Z(n5734) );
  XNOR U7887 ( .A(n5735), .B(n5736), .Z(n5733) );
  XNOR U7888 ( .A(y[1276]), .B(x[1276]), .Z(n5736) );
  XNOR U7889 ( .A(y[1277]), .B(x[1277]), .Z(n5735) );
  XOR U7890 ( .A(n5709), .B(n5710), .Z(n5728) );
  XNOR U7891 ( .A(n5725), .B(n5726), .Z(n5710) );
  XNOR U7892 ( .A(n5720), .B(n5721), .Z(n5726) );
  XNOR U7893 ( .A(n5722), .B(n5723), .Z(n5721) );
  XNOR U7894 ( .A(y[1273]), .B(x[1273]), .Z(n5723) );
  XNOR U7895 ( .A(y[1274]), .B(x[1274]), .Z(n5722) );
  XNOR U7896 ( .A(y[1272]), .B(x[1272]), .Z(n5720) );
  XNOR U7897 ( .A(n5714), .B(n5715), .Z(n5725) );
  XNOR U7898 ( .A(y[1269]), .B(x[1269]), .Z(n5715) );
  XNOR U7899 ( .A(n5716), .B(n5717), .Z(n5714) );
  XNOR U7900 ( .A(y[1270]), .B(x[1270]), .Z(n5717) );
  XNOR U7901 ( .A(y[1271]), .B(x[1271]), .Z(n5716) );
  XOR U7902 ( .A(n5708), .B(n5707), .Z(n5709) );
  XNOR U7903 ( .A(n5703), .B(n5704), .Z(n5707) );
  XNOR U7904 ( .A(y[1266]), .B(x[1266]), .Z(n5704) );
  XNOR U7905 ( .A(n5705), .B(n5706), .Z(n5703) );
  XNOR U7906 ( .A(y[1267]), .B(x[1267]), .Z(n5706) );
  XNOR U7907 ( .A(y[1268]), .B(x[1268]), .Z(n5705) );
  XNOR U7908 ( .A(n5697), .B(n5698), .Z(n5708) );
  XNOR U7909 ( .A(y[1263]), .B(x[1263]), .Z(n5698) );
  XNOR U7910 ( .A(n5699), .B(n5700), .Z(n5697) );
  XNOR U7911 ( .A(y[1264]), .B(x[1264]), .Z(n5700) );
  XNOR U7912 ( .A(y[1265]), .B(x[1265]), .Z(n5699) );
  NAND U7913 ( .A(n5764), .B(n5765), .Z(N13357) );
  NANDN U7914 ( .A(n5766), .B(n5767), .Z(n5765) );
  OR U7915 ( .A(n5768), .B(n5769), .Z(n5767) );
  NAND U7916 ( .A(n5768), .B(n5769), .Z(n5764) );
  XOR U7917 ( .A(n5768), .B(n5770), .Z(N13356) );
  XNOR U7918 ( .A(n5766), .B(n5769), .Z(n5770) );
  AND U7919 ( .A(n5771), .B(n5772), .Z(n5769) );
  NANDN U7920 ( .A(n5773), .B(n5774), .Z(n5772) );
  NANDN U7921 ( .A(n5775), .B(n5776), .Z(n5774) );
  NANDN U7922 ( .A(n5776), .B(n5775), .Z(n5771) );
  NAND U7923 ( .A(n5777), .B(n5778), .Z(n5766) );
  NANDN U7924 ( .A(n5779), .B(n5780), .Z(n5778) );
  OR U7925 ( .A(n5781), .B(n5782), .Z(n5780) );
  NAND U7926 ( .A(n5782), .B(n5781), .Z(n5777) );
  AND U7927 ( .A(n5783), .B(n5784), .Z(n5768) );
  NANDN U7928 ( .A(n5785), .B(n5786), .Z(n5784) );
  NANDN U7929 ( .A(n5787), .B(n5788), .Z(n5786) );
  NANDN U7930 ( .A(n5788), .B(n5787), .Z(n5783) );
  XOR U7931 ( .A(n5782), .B(n5789), .Z(N13355) );
  XOR U7932 ( .A(n5779), .B(n5781), .Z(n5789) );
  XNOR U7933 ( .A(n5775), .B(n5790), .Z(n5781) );
  XNOR U7934 ( .A(n5773), .B(n5776), .Z(n5790) );
  NAND U7935 ( .A(n5791), .B(n5792), .Z(n5776) );
  NAND U7936 ( .A(n5793), .B(n5794), .Z(n5792) );
  OR U7937 ( .A(n5795), .B(n5796), .Z(n5793) );
  NANDN U7938 ( .A(n5797), .B(n5795), .Z(n5791) );
  IV U7939 ( .A(n5796), .Z(n5797) );
  NAND U7940 ( .A(n5798), .B(n5799), .Z(n5773) );
  NAND U7941 ( .A(n5800), .B(n5801), .Z(n5799) );
  NANDN U7942 ( .A(n5802), .B(n5803), .Z(n5800) );
  NANDN U7943 ( .A(n5803), .B(n5802), .Z(n5798) );
  AND U7944 ( .A(n5804), .B(n5805), .Z(n5775) );
  NAND U7945 ( .A(n5806), .B(n5807), .Z(n5805) );
  OR U7946 ( .A(n5808), .B(n5809), .Z(n5806) );
  NANDN U7947 ( .A(n5810), .B(n5808), .Z(n5804) );
  NAND U7948 ( .A(n5811), .B(n5812), .Z(n5779) );
  NANDN U7949 ( .A(n5813), .B(n5814), .Z(n5812) );
  OR U7950 ( .A(n5815), .B(n5816), .Z(n5814) );
  NANDN U7951 ( .A(n5817), .B(n5815), .Z(n5811) );
  IV U7952 ( .A(n5816), .Z(n5817) );
  XNOR U7953 ( .A(n5787), .B(n5818), .Z(n5782) );
  XNOR U7954 ( .A(n5785), .B(n5788), .Z(n5818) );
  NAND U7955 ( .A(n5819), .B(n5820), .Z(n5788) );
  NAND U7956 ( .A(n5821), .B(n5822), .Z(n5820) );
  OR U7957 ( .A(n5823), .B(n5824), .Z(n5821) );
  NANDN U7958 ( .A(n5825), .B(n5823), .Z(n5819) );
  IV U7959 ( .A(n5824), .Z(n5825) );
  NAND U7960 ( .A(n5826), .B(n5827), .Z(n5785) );
  NAND U7961 ( .A(n5828), .B(n5829), .Z(n5827) );
  NANDN U7962 ( .A(n5830), .B(n5831), .Z(n5828) );
  NANDN U7963 ( .A(n5831), .B(n5830), .Z(n5826) );
  AND U7964 ( .A(n5832), .B(n5833), .Z(n5787) );
  NAND U7965 ( .A(n5834), .B(n5835), .Z(n5833) );
  OR U7966 ( .A(n5836), .B(n5837), .Z(n5834) );
  NANDN U7967 ( .A(n5838), .B(n5836), .Z(n5832) );
  XNOR U7968 ( .A(n5813), .B(n5839), .Z(N13354) );
  XOR U7969 ( .A(n5815), .B(n5816), .Z(n5839) );
  XNOR U7970 ( .A(n5829), .B(n5840), .Z(n5816) );
  XOR U7971 ( .A(n5830), .B(n5831), .Z(n5840) );
  XOR U7972 ( .A(n5836), .B(n5841), .Z(n5831) );
  XOR U7973 ( .A(n5835), .B(n5838), .Z(n5841) );
  IV U7974 ( .A(n5837), .Z(n5838) );
  NAND U7975 ( .A(n5842), .B(n5843), .Z(n5837) );
  OR U7976 ( .A(n5844), .B(n5845), .Z(n5843) );
  OR U7977 ( .A(n5846), .B(n5847), .Z(n5842) );
  NAND U7978 ( .A(n5848), .B(n5849), .Z(n5835) );
  OR U7979 ( .A(n5850), .B(n5851), .Z(n5849) );
  OR U7980 ( .A(n5852), .B(n5853), .Z(n5848) );
  NOR U7981 ( .A(n5854), .B(n5855), .Z(n5836) );
  ANDN U7982 ( .B(n5856), .A(n5857), .Z(n5830) );
  XNOR U7983 ( .A(n5823), .B(n5858), .Z(n5829) );
  XNOR U7984 ( .A(n5822), .B(n5824), .Z(n5858) );
  NAND U7985 ( .A(n5859), .B(n5860), .Z(n5824) );
  OR U7986 ( .A(n5861), .B(n5862), .Z(n5860) );
  OR U7987 ( .A(n5863), .B(n5864), .Z(n5859) );
  NAND U7988 ( .A(n5865), .B(n5866), .Z(n5822) );
  OR U7989 ( .A(n5867), .B(n5868), .Z(n5866) );
  OR U7990 ( .A(n5869), .B(n5870), .Z(n5865) );
  ANDN U7991 ( .B(n5871), .A(n5872), .Z(n5823) );
  IV U7992 ( .A(n5873), .Z(n5871) );
  ANDN U7993 ( .B(n5874), .A(n5875), .Z(n5815) );
  XOR U7994 ( .A(n5801), .B(n5876), .Z(n5813) );
  XOR U7995 ( .A(n5802), .B(n5803), .Z(n5876) );
  XOR U7996 ( .A(n5808), .B(n5877), .Z(n5803) );
  XOR U7997 ( .A(n5807), .B(n5810), .Z(n5877) );
  IV U7998 ( .A(n5809), .Z(n5810) );
  NAND U7999 ( .A(n5878), .B(n5879), .Z(n5809) );
  OR U8000 ( .A(n5880), .B(n5881), .Z(n5879) );
  OR U8001 ( .A(n5882), .B(n5883), .Z(n5878) );
  NAND U8002 ( .A(n5884), .B(n5885), .Z(n5807) );
  OR U8003 ( .A(n5886), .B(n5887), .Z(n5885) );
  OR U8004 ( .A(n5888), .B(n5889), .Z(n5884) );
  NOR U8005 ( .A(n5890), .B(n5891), .Z(n5808) );
  ANDN U8006 ( .B(n5892), .A(n5893), .Z(n5802) );
  IV U8007 ( .A(n5894), .Z(n5892) );
  XNOR U8008 ( .A(n5795), .B(n5895), .Z(n5801) );
  XNOR U8009 ( .A(n5794), .B(n5796), .Z(n5895) );
  NAND U8010 ( .A(n5896), .B(n5897), .Z(n5796) );
  OR U8011 ( .A(n5898), .B(n5899), .Z(n5897) );
  OR U8012 ( .A(n5900), .B(n5901), .Z(n5896) );
  NAND U8013 ( .A(n5902), .B(n5903), .Z(n5794) );
  OR U8014 ( .A(n5904), .B(n5905), .Z(n5903) );
  OR U8015 ( .A(n5906), .B(n5907), .Z(n5902) );
  ANDN U8016 ( .B(n5908), .A(n5909), .Z(n5795) );
  IV U8017 ( .A(n5910), .Z(n5908) );
  XNOR U8018 ( .A(n5875), .B(n5874), .Z(N13353) );
  XOR U8019 ( .A(n5894), .B(n5893), .Z(n5874) );
  XNOR U8020 ( .A(n5909), .B(n5910), .Z(n5893) );
  XNOR U8021 ( .A(n5904), .B(n5905), .Z(n5910) );
  XNOR U8022 ( .A(n5906), .B(n5907), .Z(n5905) );
  XNOR U8023 ( .A(y[1261]), .B(x[1261]), .Z(n5907) );
  XNOR U8024 ( .A(y[1262]), .B(x[1262]), .Z(n5906) );
  XNOR U8025 ( .A(y[1260]), .B(x[1260]), .Z(n5904) );
  XNOR U8026 ( .A(n5898), .B(n5899), .Z(n5909) );
  XNOR U8027 ( .A(y[1257]), .B(x[1257]), .Z(n5899) );
  XNOR U8028 ( .A(n5900), .B(n5901), .Z(n5898) );
  XNOR U8029 ( .A(y[1258]), .B(x[1258]), .Z(n5901) );
  XNOR U8030 ( .A(y[1259]), .B(x[1259]), .Z(n5900) );
  XNOR U8031 ( .A(n5891), .B(n5890), .Z(n5894) );
  XNOR U8032 ( .A(n5886), .B(n5887), .Z(n5890) );
  XNOR U8033 ( .A(y[1254]), .B(x[1254]), .Z(n5887) );
  XNOR U8034 ( .A(n5888), .B(n5889), .Z(n5886) );
  XNOR U8035 ( .A(y[1255]), .B(x[1255]), .Z(n5889) );
  XNOR U8036 ( .A(y[1256]), .B(x[1256]), .Z(n5888) );
  XNOR U8037 ( .A(n5880), .B(n5881), .Z(n5891) );
  XNOR U8038 ( .A(y[1251]), .B(x[1251]), .Z(n5881) );
  XNOR U8039 ( .A(n5882), .B(n5883), .Z(n5880) );
  XNOR U8040 ( .A(y[1252]), .B(x[1252]), .Z(n5883) );
  XNOR U8041 ( .A(y[1253]), .B(x[1253]), .Z(n5882) );
  XOR U8042 ( .A(n5856), .B(n5857), .Z(n5875) );
  XNOR U8043 ( .A(n5872), .B(n5873), .Z(n5857) );
  XNOR U8044 ( .A(n5867), .B(n5868), .Z(n5873) );
  XNOR U8045 ( .A(n5869), .B(n5870), .Z(n5868) );
  XNOR U8046 ( .A(y[1249]), .B(x[1249]), .Z(n5870) );
  XNOR U8047 ( .A(y[1250]), .B(x[1250]), .Z(n5869) );
  XNOR U8048 ( .A(y[1248]), .B(x[1248]), .Z(n5867) );
  XNOR U8049 ( .A(n5861), .B(n5862), .Z(n5872) );
  XNOR U8050 ( .A(y[1245]), .B(x[1245]), .Z(n5862) );
  XNOR U8051 ( .A(n5863), .B(n5864), .Z(n5861) );
  XNOR U8052 ( .A(y[1246]), .B(x[1246]), .Z(n5864) );
  XNOR U8053 ( .A(y[1247]), .B(x[1247]), .Z(n5863) );
  XOR U8054 ( .A(n5855), .B(n5854), .Z(n5856) );
  XNOR U8055 ( .A(n5850), .B(n5851), .Z(n5854) );
  XNOR U8056 ( .A(y[1242]), .B(x[1242]), .Z(n5851) );
  XNOR U8057 ( .A(n5852), .B(n5853), .Z(n5850) );
  XNOR U8058 ( .A(y[1243]), .B(x[1243]), .Z(n5853) );
  XNOR U8059 ( .A(y[1244]), .B(x[1244]), .Z(n5852) );
  XNOR U8060 ( .A(n5844), .B(n5845), .Z(n5855) );
  XNOR U8061 ( .A(y[1239]), .B(x[1239]), .Z(n5845) );
  XNOR U8062 ( .A(n5846), .B(n5847), .Z(n5844) );
  XNOR U8063 ( .A(y[1240]), .B(x[1240]), .Z(n5847) );
  XNOR U8064 ( .A(y[1241]), .B(x[1241]), .Z(n5846) );
  NAND U8065 ( .A(n5911), .B(n5912), .Z(N13346) );
  NANDN U8066 ( .A(n5913), .B(n5914), .Z(n5912) );
  OR U8067 ( .A(n5915), .B(n5916), .Z(n5914) );
  NAND U8068 ( .A(n5915), .B(n5916), .Z(n5911) );
  XOR U8069 ( .A(n5915), .B(n5917), .Z(N13345) );
  XNOR U8070 ( .A(n5913), .B(n5916), .Z(n5917) );
  AND U8071 ( .A(n5918), .B(n5919), .Z(n5916) );
  NANDN U8072 ( .A(n5920), .B(n5921), .Z(n5919) );
  NANDN U8073 ( .A(n5922), .B(n5923), .Z(n5921) );
  NANDN U8074 ( .A(n5923), .B(n5922), .Z(n5918) );
  NAND U8075 ( .A(n5924), .B(n5925), .Z(n5913) );
  NANDN U8076 ( .A(n5926), .B(n5927), .Z(n5925) );
  OR U8077 ( .A(n5928), .B(n5929), .Z(n5927) );
  NAND U8078 ( .A(n5929), .B(n5928), .Z(n5924) );
  AND U8079 ( .A(n5930), .B(n5931), .Z(n5915) );
  NANDN U8080 ( .A(n5932), .B(n5933), .Z(n5931) );
  NANDN U8081 ( .A(n5934), .B(n5935), .Z(n5933) );
  NANDN U8082 ( .A(n5935), .B(n5934), .Z(n5930) );
  XOR U8083 ( .A(n5929), .B(n5936), .Z(N13344) );
  XOR U8084 ( .A(n5926), .B(n5928), .Z(n5936) );
  XNOR U8085 ( .A(n5922), .B(n5937), .Z(n5928) );
  XNOR U8086 ( .A(n5920), .B(n5923), .Z(n5937) );
  NAND U8087 ( .A(n5938), .B(n5939), .Z(n5923) );
  NAND U8088 ( .A(n5940), .B(n5941), .Z(n5939) );
  OR U8089 ( .A(n5942), .B(n5943), .Z(n5940) );
  NANDN U8090 ( .A(n5944), .B(n5942), .Z(n5938) );
  IV U8091 ( .A(n5943), .Z(n5944) );
  NAND U8092 ( .A(n5945), .B(n5946), .Z(n5920) );
  NAND U8093 ( .A(n5947), .B(n5948), .Z(n5946) );
  NANDN U8094 ( .A(n5949), .B(n5950), .Z(n5947) );
  NANDN U8095 ( .A(n5950), .B(n5949), .Z(n5945) );
  AND U8096 ( .A(n5951), .B(n5952), .Z(n5922) );
  NAND U8097 ( .A(n5953), .B(n5954), .Z(n5952) );
  OR U8098 ( .A(n5955), .B(n5956), .Z(n5953) );
  NANDN U8099 ( .A(n5957), .B(n5955), .Z(n5951) );
  NAND U8100 ( .A(n5958), .B(n5959), .Z(n5926) );
  NANDN U8101 ( .A(n5960), .B(n5961), .Z(n5959) );
  OR U8102 ( .A(n5962), .B(n5963), .Z(n5961) );
  NANDN U8103 ( .A(n5964), .B(n5962), .Z(n5958) );
  IV U8104 ( .A(n5963), .Z(n5964) );
  XNOR U8105 ( .A(n5934), .B(n5965), .Z(n5929) );
  XNOR U8106 ( .A(n5932), .B(n5935), .Z(n5965) );
  NAND U8107 ( .A(n5966), .B(n5967), .Z(n5935) );
  NAND U8108 ( .A(n5968), .B(n5969), .Z(n5967) );
  OR U8109 ( .A(n5970), .B(n5971), .Z(n5968) );
  NANDN U8110 ( .A(n5972), .B(n5970), .Z(n5966) );
  IV U8111 ( .A(n5971), .Z(n5972) );
  NAND U8112 ( .A(n5973), .B(n5974), .Z(n5932) );
  NAND U8113 ( .A(n5975), .B(n5976), .Z(n5974) );
  NANDN U8114 ( .A(n5977), .B(n5978), .Z(n5975) );
  NANDN U8115 ( .A(n5978), .B(n5977), .Z(n5973) );
  AND U8116 ( .A(n5979), .B(n5980), .Z(n5934) );
  NAND U8117 ( .A(n5981), .B(n5982), .Z(n5980) );
  OR U8118 ( .A(n5983), .B(n5984), .Z(n5981) );
  NANDN U8119 ( .A(n5985), .B(n5983), .Z(n5979) );
  XNOR U8120 ( .A(n5960), .B(n5986), .Z(N13343) );
  XOR U8121 ( .A(n5962), .B(n5963), .Z(n5986) );
  XNOR U8122 ( .A(n5976), .B(n5987), .Z(n5963) );
  XOR U8123 ( .A(n5977), .B(n5978), .Z(n5987) );
  XOR U8124 ( .A(n5983), .B(n5988), .Z(n5978) );
  XOR U8125 ( .A(n5982), .B(n5985), .Z(n5988) );
  IV U8126 ( .A(n5984), .Z(n5985) );
  NAND U8127 ( .A(n5989), .B(n5990), .Z(n5984) );
  OR U8128 ( .A(n5991), .B(n5992), .Z(n5990) );
  OR U8129 ( .A(n5993), .B(n5994), .Z(n5989) );
  NAND U8130 ( .A(n5995), .B(n5996), .Z(n5982) );
  OR U8131 ( .A(n5997), .B(n5998), .Z(n5996) );
  OR U8132 ( .A(n5999), .B(n6000), .Z(n5995) );
  NOR U8133 ( .A(n6001), .B(n6002), .Z(n5983) );
  ANDN U8134 ( .B(n6003), .A(n6004), .Z(n5977) );
  XNOR U8135 ( .A(n5970), .B(n6005), .Z(n5976) );
  XNOR U8136 ( .A(n5969), .B(n5971), .Z(n6005) );
  NAND U8137 ( .A(n6006), .B(n6007), .Z(n5971) );
  OR U8138 ( .A(n6008), .B(n6009), .Z(n6007) );
  OR U8139 ( .A(n6010), .B(n6011), .Z(n6006) );
  NAND U8140 ( .A(n6012), .B(n6013), .Z(n5969) );
  OR U8141 ( .A(n6014), .B(n6015), .Z(n6013) );
  OR U8142 ( .A(n6016), .B(n6017), .Z(n6012) );
  ANDN U8143 ( .B(n6018), .A(n6019), .Z(n5970) );
  IV U8144 ( .A(n6020), .Z(n6018) );
  ANDN U8145 ( .B(n6021), .A(n6022), .Z(n5962) );
  XOR U8146 ( .A(n5948), .B(n6023), .Z(n5960) );
  XOR U8147 ( .A(n5949), .B(n5950), .Z(n6023) );
  XOR U8148 ( .A(n5955), .B(n6024), .Z(n5950) );
  XOR U8149 ( .A(n5954), .B(n5957), .Z(n6024) );
  IV U8150 ( .A(n5956), .Z(n5957) );
  NAND U8151 ( .A(n6025), .B(n6026), .Z(n5956) );
  OR U8152 ( .A(n6027), .B(n6028), .Z(n6026) );
  OR U8153 ( .A(n6029), .B(n6030), .Z(n6025) );
  NAND U8154 ( .A(n6031), .B(n6032), .Z(n5954) );
  OR U8155 ( .A(n6033), .B(n6034), .Z(n6032) );
  OR U8156 ( .A(n6035), .B(n6036), .Z(n6031) );
  NOR U8157 ( .A(n6037), .B(n6038), .Z(n5955) );
  ANDN U8158 ( .B(n6039), .A(n6040), .Z(n5949) );
  IV U8159 ( .A(n6041), .Z(n6039) );
  XNOR U8160 ( .A(n5942), .B(n6042), .Z(n5948) );
  XNOR U8161 ( .A(n5941), .B(n5943), .Z(n6042) );
  NAND U8162 ( .A(n6043), .B(n6044), .Z(n5943) );
  OR U8163 ( .A(n6045), .B(n6046), .Z(n6044) );
  OR U8164 ( .A(n6047), .B(n6048), .Z(n6043) );
  NAND U8165 ( .A(n6049), .B(n6050), .Z(n5941) );
  OR U8166 ( .A(n6051), .B(n6052), .Z(n6050) );
  OR U8167 ( .A(n6053), .B(n6054), .Z(n6049) );
  ANDN U8168 ( .B(n6055), .A(n6056), .Z(n5942) );
  IV U8169 ( .A(n6057), .Z(n6055) );
  XNOR U8170 ( .A(n6022), .B(n6021), .Z(N13342) );
  XOR U8171 ( .A(n6041), .B(n6040), .Z(n6021) );
  XNOR U8172 ( .A(n6056), .B(n6057), .Z(n6040) );
  XNOR U8173 ( .A(n6051), .B(n6052), .Z(n6057) );
  XNOR U8174 ( .A(n6053), .B(n6054), .Z(n6052) );
  XNOR U8175 ( .A(y[1237]), .B(x[1237]), .Z(n6054) );
  XNOR U8176 ( .A(y[1238]), .B(x[1238]), .Z(n6053) );
  XNOR U8177 ( .A(y[1236]), .B(x[1236]), .Z(n6051) );
  XNOR U8178 ( .A(n6045), .B(n6046), .Z(n6056) );
  XNOR U8179 ( .A(y[1233]), .B(x[1233]), .Z(n6046) );
  XNOR U8180 ( .A(n6047), .B(n6048), .Z(n6045) );
  XNOR U8181 ( .A(y[1234]), .B(x[1234]), .Z(n6048) );
  XNOR U8182 ( .A(y[1235]), .B(x[1235]), .Z(n6047) );
  XNOR U8183 ( .A(n6038), .B(n6037), .Z(n6041) );
  XNOR U8184 ( .A(n6033), .B(n6034), .Z(n6037) );
  XNOR U8185 ( .A(y[1230]), .B(x[1230]), .Z(n6034) );
  XNOR U8186 ( .A(n6035), .B(n6036), .Z(n6033) );
  XNOR U8187 ( .A(y[1231]), .B(x[1231]), .Z(n6036) );
  XNOR U8188 ( .A(y[1232]), .B(x[1232]), .Z(n6035) );
  XNOR U8189 ( .A(n6027), .B(n6028), .Z(n6038) );
  XNOR U8190 ( .A(y[1227]), .B(x[1227]), .Z(n6028) );
  XNOR U8191 ( .A(n6029), .B(n6030), .Z(n6027) );
  XNOR U8192 ( .A(y[1228]), .B(x[1228]), .Z(n6030) );
  XNOR U8193 ( .A(y[1229]), .B(x[1229]), .Z(n6029) );
  XOR U8194 ( .A(n6003), .B(n6004), .Z(n6022) );
  XNOR U8195 ( .A(n6019), .B(n6020), .Z(n6004) );
  XNOR U8196 ( .A(n6014), .B(n6015), .Z(n6020) );
  XNOR U8197 ( .A(n6016), .B(n6017), .Z(n6015) );
  XNOR U8198 ( .A(y[1225]), .B(x[1225]), .Z(n6017) );
  XNOR U8199 ( .A(y[1226]), .B(x[1226]), .Z(n6016) );
  XNOR U8200 ( .A(y[1224]), .B(x[1224]), .Z(n6014) );
  XNOR U8201 ( .A(n6008), .B(n6009), .Z(n6019) );
  XNOR U8202 ( .A(y[1221]), .B(x[1221]), .Z(n6009) );
  XNOR U8203 ( .A(n6010), .B(n6011), .Z(n6008) );
  XNOR U8204 ( .A(y[1222]), .B(x[1222]), .Z(n6011) );
  XNOR U8205 ( .A(y[1223]), .B(x[1223]), .Z(n6010) );
  XOR U8206 ( .A(n6002), .B(n6001), .Z(n6003) );
  XNOR U8207 ( .A(n5997), .B(n5998), .Z(n6001) );
  XNOR U8208 ( .A(y[1218]), .B(x[1218]), .Z(n5998) );
  XNOR U8209 ( .A(n5999), .B(n6000), .Z(n5997) );
  XNOR U8210 ( .A(y[1219]), .B(x[1219]), .Z(n6000) );
  XNOR U8211 ( .A(y[1220]), .B(x[1220]), .Z(n5999) );
  XNOR U8212 ( .A(n5991), .B(n5992), .Z(n6002) );
  XNOR U8213 ( .A(y[1215]), .B(x[1215]), .Z(n5992) );
  XNOR U8214 ( .A(n5993), .B(n5994), .Z(n5991) );
  XNOR U8215 ( .A(y[1216]), .B(x[1216]), .Z(n5994) );
  XNOR U8216 ( .A(y[1217]), .B(x[1217]), .Z(n5993) );
  NAND U8217 ( .A(n6058), .B(n6059), .Z(N13335) );
  NANDN U8218 ( .A(n6060), .B(n6061), .Z(n6059) );
  OR U8219 ( .A(n6062), .B(n6063), .Z(n6061) );
  NAND U8220 ( .A(n6062), .B(n6063), .Z(n6058) );
  XOR U8221 ( .A(n6062), .B(n6064), .Z(N13334) );
  XNOR U8222 ( .A(n6060), .B(n6063), .Z(n6064) );
  AND U8223 ( .A(n6065), .B(n6066), .Z(n6063) );
  NANDN U8224 ( .A(n6067), .B(n6068), .Z(n6066) );
  NANDN U8225 ( .A(n6069), .B(n6070), .Z(n6068) );
  NANDN U8226 ( .A(n6070), .B(n6069), .Z(n6065) );
  NAND U8227 ( .A(n6071), .B(n6072), .Z(n6060) );
  NANDN U8228 ( .A(n6073), .B(n6074), .Z(n6072) );
  OR U8229 ( .A(n6075), .B(n6076), .Z(n6074) );
  NAND U8230 ( .A(n6076), .B(n6075), .Z(n6071) );
  AND U8231 ( .A(n6077), .B(n6078), .Z(n6062) );
  NANDN U8232 ( .A(n6079), .B(n6080), .Z(n6078) );
  NANDN U8233 ( .A(n6081), .B(n6082), .Z(n6080) );
  NANDN U8234 ( .A(n6082), .B(n6081), .Z(n6077) );
  XOR U8235 ( .A(n6076), .B(n6083), .Z(N13333) );
  XOR U8236 ( .A(n6073), .B(n6075), .Z(n6083) );
  XNOR U8237 ( .A(n6069), .B(n6084), .Z(n6075) );
  XNOR U8238 ( .A(n6067), .B(n6070), .Z(n6084) );
  NAND U8239 ( .A(n6085), .B(n6086), .Z(n6070) );
  NAND U8240 ( .A(n6087), .B(n6088), .Z(n6086) );
  OR U8241 ( .A(n6089), .B(n6090), .Z(n6087) );
  NANDN U8242 ( .A(n6091), .B(n6089), .Z(n6085) );
  IV U8243 ( .A(n6090), .Z(n6091) );
  NAND U8244 ( .A(n6092), .B(n6093), .Z(n6067) );
  NAND U8245 ( .A(n6094), .B(n6095), .Z(n6093) );
  NANDN U8246 ( .A(n6096), .B(n6097), .Z(n6094) );
  NANDN U8247 ( .A(n6097), .B(n6096), .Z(n6092) );
  AND U8248 ( .A(n6098), .B(n6099), .Z(n6069) );
  NAND U8249 ( .A(n6100), .B(n6101), .Z(n6099) );
  OR U8250 ( .A(n6102), .B(n6103), .Z(n6100) );
  NANDN U8251 ( .A(n6104), .B(n6102), .Z(n6098) );
  NAND U8252 ( .A(n6105), .B(n6106), .Z(n6073) );
  NANDN U8253 ( .A(n6107), .B(n6108), .Z(n6106) );
  OR U8254 ( .A(n6109), .B(n6110), .Z(n6108) );
  NANDN U8255 ( .A(n6111), .B(n6109), .Z(n6105) );
  IV U8256 ( .A(n6110), .Z(n6111) );
  XNOR U8257 ( .A(n6081), .B(n6112), .Z(n6076) );
  XNOR U8258 ( .A(n6079), .B(n6082), .Z(n6112) );
  NAND U8259 ( .A(n6113), .B(n6114), .Z(n6082) );
  NAND U8260 ( .A(n6115), .B(n6116), .Z(n6114) );
  OR U8261 ( .A(n6117), .B(n6118), .Z(n6115) );
  NANDN U8262 ( .A(n6119), .B(n6117), .Z(n6113) );
  IV U8263 ( .A(n6118), .Z(n6119) );
  NAND U8264 ( .A(n6120), .B(n6121), .Z(n6079) );
  NAND U8265 ( .A(n6122), .B(n6123), .Z(n6121) );
  NANDN U8266 ( .A(n6124), .B(n6125), .Z(n6122) );
  NANDN U8267 ( .A(n6125), .B(n6124), .Z(n6120) );
  AND U8268 ( .A(n6126), .B(n6127), .Z(n6081) );
  NAND U8269 ( .A(n6128), .B(n6129), .Z(n6127) );
  OR U8270 ( .A(n6130), .B(n6131), .Z(n6128) );
  NANDN U8271 ( .A(n6132), .B(n6130), .Z(n6126) );
  XNOR U8272 ( .A(n6107), .B(n6133), .Z(N13332) );
  XOR U8273 ( .A(n6109), .B(n6110), .Z(n6133) );
  XNOR U8274 ( .A(n6123), .B(n6134), .Z(n6110) );
  XOR U8275 ( .A(n6124), .B(n6125), .Z(n6134) );
  XOR U8276 ( .A(n6130), .B(n6135), .Z(n6125) );
  XOR U8277 ( .A(n6129), .B(n6132), .Z(n6135) );
  IV U8278 ( .A(n6131), .Z(n6132) );
  NAND U8279 ( .A(n6136), .B(n6137), .Z(n6131) );
  OR U8280 ( .A(n6138), .B(n6139), .Z(n6137) );
  OR U8281 ( .A(n6140), .B(n6141), .Z(n6136) );
  NAND U8282 ( .A(n6142), .B(n6143), .Z(n6129) );
  OR U8283 ( .A(n6144), .B(n6145), .Z(n6143) );
  OR U8284 ( .A(n6146), .B(n6147), .Z(n6142) );
  NOR U8285 ( .A(n6148), .B(n6149), .Z(n6130) );
  ANDN U8286 ( .B(n6150), .A(n6151), .Z(n6124) );
  XNOR U8287 ( .A(n6117), .B(n6152), .Z(n6123) );
  XNOR U8288 ( .A(n6116), .B(n6118), .Z(n6152) );
  NAND U8289 ( .A(n6153), .B(n6154), .Z(n6118) );
  OR U8290 ( .A(n6155), .B(n6156), .Z(n6154) );
  OR U8291 ( .A(n6157), .B(n6158), .Z(n6153) );
  NAND U8292 ( .A(n6159), .B(n6160), .Z(n6116) );
  OR U8293 ( .A(n6161), .B(n6162), .Z(n6160) );
  OR U8294 ( .A(n6163), .B(n6164), .Z(n6159) );
  ANDN U8295 ( .B(n6165), .A(n6166), .Z(n6117) );
  IV U8296 ( .A(n6167), .Z(n6165) );
  ANDN U8297 ( .B(n6168), .A(n6169), .Z(n6109) );
  XOR U8298 ( .A(n6095), .B(n6170), .Z(n6107) );
  XOR U8299 ( .A(n6096), .B(n6097), .Z(n6170) );
  XOR U8300 ( .A(n6102), .B(n6171), .Z(n6097) );
  XOR U8301 ( .A(n6101), .B(n6104), .Z(n6171) );
  IV U8302 ( .A(n6103), .Z(n6104) );
  NAND U8303 ( .A(n6172), .B(n6173), .Z(n6103) );
  OR U8304 ( .A(n6174), .B(n6175), .Z(n6173) );
  OR U8305 ( .A(n6176), .B(n6177), .Z(n6172) );
  NAND U8306 ( .A(n6178), .B(n6179), .Z(n6101) );
  OR U8307 ( .A(n6180), .B(n6181), .Z(n6179) );
  OR U8308 ( .A(n6182), .B(n6183), .Z(n6178) );
  NOR U8309 ( .A(n6184), .B(n6185), .Z(n6102) );
  ANDN U8310 ( .B(n6186), .A(n6187), .Z(n6096) );
  IV U8311 ( .A(n6188), .Z(n6186) );
  XNOR U8312 ( .A(n6089), .B(n6189), .Z(n6095) );
  XNOR U8313 ( .A(n6088), .B(n6090), .Z(n6189) );
  NAND U8314 ( .A(n6190), .B(n6191), .Z(n6090) );
  OR U8315 ( .A(n6192), .B(n6193), .Z(n6191) );
  OR U8316 ( .A(n6194), .B(n6195), .Z(n6190) );
  NAND U8317 ( .A(n6196), .B(n6197), .Z(n6088) );
  OR U8318 ( .A(n6198), .B(n6199), .Z(n6197) );
  OR U8319 ( .A(n6200), .B(n6201), .Z(n6196) );
  ANDN U8320 ( .B(n6202), .A(n6203), .Z(n6089) );
  IV U8321 ( .A(n6204), .Z(n6202) );
  XNOR U8322 ( .A(n6169), .B(n6168), .Z(N13331) );
  XOR U8323 ( .A(n6188), .B(n6187), .Z(n6168) );
  XNOR U8324 ( .A(n6203), .B(n6204), .Z(n6187) );
  XNOR U8325 ( .A(n6198), .B(n6199), .Z(n6204) );
  XNOR U8326 ( .A(n6200), .B(n6201), .Z(n6199) );
  XNOR U8327 ( .A(y[1213]), .B(x[1213]), .Z(n6201) );
  XNOR U8328 ( .A(y[1214]), .B(x[1214]), .Z(n6200) );
  XNOR U8329 ( .A(y[1212]), .B(x[1212]), .Z(n6198) );
  XNOR U8330 ( .A(n6192), .B(n6193), .Z(n6203) );
  XNOR U8331 ( .A(y[1209]), .B(x[1209]), .Z(n6193) );
  XNOR U8332 ( .A(n6194), .B(n6195), .Z(n6192) );
  XNOR U8333 ( .A(y[1210]), .B(x[1210]), .Z(n6195) );
  XNOR U8334 ( .A(y[1211]), .B(x[1211]), .Z(n6194) );
  XNOR U8335 ( .A(n6185), .B(n6184), .Z(n6188) );
  XNOR U8336 ( .A(n6180), .B(n6181), .Z(n6184) );
  XNOR U8337 ( .A(y[1206]), .B(x[1206]), .Z(n6181) );
  XNOR U8338 ( .A(n6182), .B(n6183), .Z(n6180) );
  XNOR U8339 ( .A(y[1207]), .B(x[1207]), .Z(n6183) );
  XNOR U8340 ( .A(y[1208]), .B(x[1208]), .Z(n6182) );
  XNOR U8341 ( .A(n6174), .B(n6175), .Z(n6185) );
  XNOR U8342 ( .A(y[1203]), .B(x[1203]), .Z(n6175) );
  XNOR U8343 ( .A(n6176), .B(n6177), .Z(n6174) );
  XNOR U8344 ( .A(y[1204]), .B(x[1204]), .Z(n6177) );
  XNOR U8345 ( .A(y[1205]), .B(x[1205]), .Z(n6176) );
  XOR U8346 ( .A(n6150), .B(n6151), .Z(n6169) );
  XNOR U8347 ( .A(n6166), .B(n6167), .Z(n6151) );
  XNOR U8348 ( .A(n6161), .B(n6162), .Z(n6167) );
  XNOR U8349 ( .A(n6163), .B(n6164), .Z(n6162) );
  XNOR U8350 ( .A(y[1201]), .B(x[1201]), .Z(n6164) );
  XNOR U8351 ( .A(y[1202]), .B(x[1202]), .Z(n6163) );
  XNOR U8352 ( .A(y[1200]), .B(x[1200]), .Z(n6161) );
  XNOR U8353 ( .A(n6155), .B(n6156), .Z(n6166) );
  XNOR U8354 ( .A(y[1197]), .B(x[1197]), .Z(n6156) );
  XNOR U8355 ( .A(n6157), .B(n6158), .Z(n6155) );
  XNOR U8356 ( .A(y[1198]), .B(x[1198]), .Z(n6158) );
  XNOR U8357 ( .A(y[1199]), .B(x[1199]), .Z(n6157) );
  XOR U8358 ( .A(n6149), .B(n6148), .Z(n6150) );
  XNOR U8359 ( .A(n6144), .B(n6145), .Z(n6148) );
  XNOR U8360 ( .A(y[1194]), .B(x[1194]), .Z(n6145) );
  XNOR U8361 ( .A(n6146), .B(n6147), .Z(n6144) );
  XNOR U8362 ( .A(y[1195]), .B(x[1195]), .Z(n6147) );
  XNOR U8363 ( .A(y[1196]), .B(x[1196]), .Z(n6146) );
  XNOR U8364 ( .A(n6138), .B(n6139), .Z(n6149) );
  XNOR U8365 ( .A(y[1191]), .B(x[1191]), .Z(n6139) );
  XNOR U8366 ( .A(n6140), .B(n6141), .Z(n6138) );
  XNOR U8367 ( .A(y[1192]), .B(x[1192]), .Z(n6141) );
  XNOR U8368 ( .A(y[1193]), .B(x[1193]), .Z(n6140) );
  NAND U8369 ( .A(n6205), .B(n6206), .Z(N13324) );
  NANDN U8370 ( .A(n6207), .B(n6208), .Z(n6206) );
  OR U8371 ( .A(n6209), .B(n6210), .Z(n6208) );
  NAND U8372 ( .A(n6209), .B(n6210), .Z(n6205) );
  XOR U8373 ( .A(n6209), .B(n6211), .Z(N13323) );
  XNOR U8374 ( .A(n6207), .B(n6210), .Z(n6211) );
  AND U8375 ( .A(n6212), .B(n6213), .Z(n6210) );
  NANDN U8376 ( .A(n6214), .B(n6215), .Z(n6213) );
  NANDN U8377 ( .A(n6216), .B(n6217), .Z(n6215) );
  NANDN U8378 ( .A(n6217), .B(n6216), .Z(n6212) );
  NAND U8379 ( .A(n6218), .B(n6219), .Z(n6207) );
  NANDN U8380 ( .A(n6220), .B(n6221), .Z(n6219) );
  OR U8381 ( .A(n6222), .B(n6223), .Z(n6221) );
  NAND U8382 ( .A(n6223), .B(n6222), .Z(n6218) );
  AND U8383 ( .A(n6224), .B(n6225), .Z(n6209) );
  NANDN U8384 ( .A(n6226), .B(n6227), .Z(n6225) );
  NANDN U8385 ( .A(n6228), .B(n6229), .Z(n6227) );
  NANDN U8386 ( .A(n6229), .B(n6228), .Z(n6224) );
  XOR U8387 ( .A(n6223), .B(n6230), .Z(N13322) );
  XOR U8388 ( .A(n6220), .B(n6222), .Z(n6230) );
  XNOR U8389 ( .A(n6216), .B(n6231), .Z(n6222) );
  XNOR U8390 ( .A(n6214), .B(n6217), .Z(n6231) );
  NAND U8391 ( .A(n6232), .B(n6233), .Z(n6217) );
  NAND U8392 ( .A(n6234), .B(n6235), .Z(n6233) );
  OR U8393 ( .A(n6236), .B(n6237), .Z(n6234) );
  NANDN U8394 ( .A(n6238), .B(n6236), .Z(n6232) );
  IV U8395 ( .A(n6237), .Z(n6238) );
  NAND U8396 ( .A(n6239), .B(n6240), .Z(n6214) );
  NAND U8397 ( .A(n6241), .B(n6242), .Z(n6240) );
  NANDN U8398 ( .A(n6243), .B(n6244), .Z(n6241) );
  NANDN U8399 ( .A(n6244), .B(n6243), .Z(n6239) );
  AND U8400 ( .A(n6245), .B(n6246), .Z(n6216) );
  NAND U8401 ( .A(n6247), .B(n6248), .Z(n6246) );
  OR U8402 ( .A(n6249), .B(n6250), .Z(n6247) );
  NANDN U8403 ( .A(n6251), .B(n6249), .Z(n6245) );
  NAND U8404 ( .A(n6252), .B(n6253), .Z(n6220) );
  NANDN U8405 ( .A(n6254), .B(n6255), .Z(n6253) );
  OR U8406 ( .A(n6256), .B(n6257), .Z(n6255) );
  NANDN U8407 ( .A(n6258), .B(n6256), .Z(n6252) );
  IV U8408 ( .A(n6257), .Z(n6258) );
  XNOR U8409 ( .A(n6228), .B(n6259), .Z(n6223) );
  XNOR U8410 ( .A(n6226), .B(n6229), .Z(n6259) );
  NAND U8411 ( .A(n6260), .B(n6261), .Z(n6229) );
  NAND U8412 ( .A(n6262), .B(n6263), .Z(n6261) );
  OR U8413 ( .A(n6264), .B(n6265), .Z(n6262) );
  NANDN U8414 ( .A(n6266), .B(n6264), .Z(n6260) );
  IV U8415 ( .A(n6265), .Z(n6266) );
  NAND U8416 ( .A(n6267), .B(n6268), .Z(n6226) );
  NAND U8417 ( .A(n6269), .B(n6270), .Z(n6268) );
  NANDN U8418 ( .A(n6271), .B(n6272), .Z(n6269) );
  NANDN U8419 ( .A(n6272), .B(n6271), .Z(n6267) );
  AND U8420 ( .A(n6273), .B(n6274), .Z(n6228) );
  NAND U8421 ( .A(n6275), .B(n6276), .Z(n6274) );
  OR U8422 ( .A(n6277), .B(n6278), .Z(n6275) );
  NANDN U8423 ( .A(n6279), .B(n6277), .Z(n6273) );
  XNOR U8424 ( .A(n6254), .B(n6280), .Z(N13321) );
  XOR U8425 ( .A(n6256), .B(n6257), .Z(n6280) );
  XNOR U8426 ( .A(n6270), .B(n6281), .Z(n6257) );
  XOR U8427 ( .A(n6271), .B(n6272), .Z(n6281) );
  XOR U8428 ( .A(n6277), .B(n6282), .Z(n6272) );
  XOR U8429 ( .A(n6276), .B(n6279), .Z(n6282) );
  IV U8430 ( .A(n6278), .Z(n6279) );
  NAND U8431 ( .A(n6283), .B(n6284), .Z(n6278) );
  OR U8432 ( .A(n6285), .B(n6286), .Z(n6284) );
  OR U8433 ( .A(n6287), .B(n6288), .Z(n6283) );
  NAND U8434 ( .A(n6289), .B(n6290), .Z(n6276) );
  OR U8435 ( .A(n6291), .B(n6292), .Z(n6290) );
  OR U8436 ( .A(n6293), .B(n6294), .Z(n6289) );
  NOR U8437 ( .A(n6295), .B(n6296), .Z(n6277) );
  ANDN U8438 ( .B(n6297), .A(n6298), .Z(n6271) );
  XNOR U8439 ( .A(n6264), .B(n6299), .Z(n6270) );
  XNOR U8440 ( .A(n6263), .B(n6265), .Z(n6299) );
  NAND U8441 ( .A(n6300), .B(n6301), .Z(n6265) );
  OR U8442 ( .A(n6302), .B(n6303), .Z(n6301) );
  OR U8443 ( .A(n6304), .B(n6305), .Z(n6300) );
  NAND U8444 ( .A(n6306), .B(n6307), .Z(n6263) );
  OR U8445 ( .A(n6308), .B(n6309), .Z(n6307) );
  OR U8446 ( .A(n6310), .B(n6311), .Z(n6306) );
  ANDN U8447 ( .B(n6312), .A(n6313), .Z(n6264) );
  IV U8448 ( .A(n6314), .Z(n6312) );
  ANDN U8449 ( .B(n6315), .A(n6316), .Z(n6256) );
  XOR U8450 ( .A(n6242), .B(n6317), .Z(n6254) );
  XOR U8451 ( .A(n6243), .B(n6244), .Z(n6317) );
  XOR U8452 ( .A(n6249), .B(n6318), .Z(n6244) );
  XOR U8453 ( .A(n6248), .B(n6251), .Z(n6318) );
  IV U8454 ( .A(n6250), .Z(n6251) );
  NAND U8455 ( .A(n6319), .B(n6320), .Z(n6250) );
  OR U8456 ( .A(n6321), .B(n6322), .Z(n6320) );
  OR U8457 ( .A(n6323), .B(n6324), .Z(n6319) );
  NAND U8458 ( .A(n6325), .B(n6326), .Z(n6248) );
  OR U8459 ( .A(n6327), .B(n6328), .Z(n6326) );
  OR U8460 ( .A(n6329), .B(n6330), .Z(n6325) );
  NOR U8461 ( .A(n6331), .B(n6332), .Z(n6249) );
  ANDN U8462 ( .B(n6333), .A(n6334), .Z(n6243) );
  IV U8463 ( .A(n6335), .Z(n6333) );
  XNOR U8464 ( .A(n6236), .B(n6336), .Z(n6242) );
  XNOR U8465 ( .A(n6235), .B(n6237), .Z(n6336) );
  NAND U8466 ( .A(n6337), .B(n6338), .Z(n6237) );
  OR U8467 ( .A(n6339), .B(n6340), .Z(n6338) );
  OR U8468 ( .A(n6341), .B(n6342), .Z(n6337) );
  NAND U8469 ( .A(n6343), .B(n6344), .Z(n6235) );
  OR U8470 ( .A(n6345), .B(n6346), .Z(n6344) );
  OR U8471 ( .A(n6347), .B(n6348), .Z(n6343) );
  ANDN U8472 ( .B(n6349), .A(n6350), .Z(n6236) );
  IV U8473 ( .A(n6351), .Z(n6349) );
  XNOR U8474 ( .A(n6316), .B(n6315), .Z(N13320) );
  XOR U8475 ( .A(n6335), .B(n6334), .Z(n6315) );
  XNOR U8476 ( .A(n6350), .B(n6351), .Z(n6334) );
  XNOR U8477 ( .A(n6345), .B(n6346), .Z(n6351) );
  XNOR U8478 ( .A(n6347), .B(n6348), .Z(n6346) );
  XNOR U8479 ( .A(y[1189]), .B(x[1189]), .Z(n6348) );
  XNOR U8480 ( .A(y[1190]), .B(x[1190]), .Z(n6347) );
  XNOR U8481 ( .A(y[1188]), .B(x[1188]), .Z(n6345) );
  XNOR U8482 ( .A(n6339), .B(n6340), .Z(n6350) );
  XNOR U8483 ( .A(y[1185]), .B(x[1185]), .Z(n6340) );
  XNOR U8484 ( .A(n6341), .B(n6342), .Z(n6339) );
  XNOR U8485 ( .A(y[1186]), .B(x[1186]), .Z(n6342) );
  XNOR U8486 ( .A(y[1187]), .B(x[1187]), .Z(n6341) );
  XNOR U8487 ( .A(n6332), .B(n6331), .Z(n6335) );
  XNOR U8488 ( .A(n6327), .B(n6328), .Z(n6331) );
  XNOR U8489 ( .A(y[1182]), .B(x[1182]), .Z(n6328) );
  XNOR U8490 ( .A(n6329), .B(n6330), .Z(n6327) );
  XNOR U8491 ( .A(y[1183]), .B(x[1183]), .Z(n6330) );
  XNOR U8492 ( .A(y[1184]), .B(x[1184]), .Z(n6329) );
  XNOR U8493 ( .A(n6321), .B(n6322), .Z(n6332) );
  XNOR U8494 ( .A(y[1179]), .B(x[1179]), .Z(n6322) );
  XNOR U8495 ( .A(n6323), .B(n6324), .Z(n6321) );
  XNOR U8496 ( .A(y[1180]), .B(x[1180]), .Z(n6324) );
  XNOR U8497 ( .A(y[1181]), .B(x[1181]), .Z(n6323) );
  XOR U8498 ( .A(n6297), .B(n6298), .Z(n6316) );
  XNOR U8499 ( .A(n6313), .B(n6314), .Z(n6298) );
  XNOR U8500 ( .A(n6308), .B(n6309), .Z(n6314) );
  XNOR U8501 ( .A(n6310), .B(n6311), .Z(n6309) );
  XNOR U8502 ( .A(y[1177]), .B(x[1177]), .Z(n6311) );
  XNOR U8503 ( .A(y[1178]), .B(x[1178]), .Z(n6310) );
  XNOR U8504 ( .A(y[1176]), .B(x[1176]), .Z(n6308) );
  XNOR U8505 ( .A(n6302), .B(n6303), .Z(n6313) );
  XNOR U8506 ( .A(y[1173]), .B(x[1173]), .Z(n6303) );
  XNOR U8507 ( .A(n6304), .B(n6305), .Z(n6302) );
  XNOR U8508 ( .A(y[1174]), .B(x[1174]), .Z(n6305) );
  XNOR U8509 ( .A(y[1175]), .B(x[1175]), .Z(n6304) );
  XOR U8510 ( .A(n6296), .B(n6295), .Z(n6297) );
  XNOR U8511 ( .A(n6291), .B(n6292), .Z(n6295) );
  XNOR U8512 ( .A(y[1170]), .B(x[1170]), .Z(n6292) );
  XNOR U8513 ( .A(n6293), .B(n6294), .Z(n6291) );
  XNOR U8514 ( .A(y[1171]), .B(x[1171]), .Z(n6294) );
  XNOR U8515 ( .A(y[1172]), .B(x[1172]), .Z(n6293) );
  XNOR U8516 ( .A(n6285), .B(n6286), .Z(n6296) );
  XNOR U8517 ( .A(y[1167]), .B(x[1167]), .Z(n6286) );
  XNOR U8518 ( .A(n6287), .B(n6288), .Z(n6285) );
  XNOR U8519 ( .A(y[1168]), .B(x[1168]), .Z(n6288) );
  XNOR U8520 ( .A(y[1169]), .B(x[1169]), .Z(n6287) );
  NAND U8521 ( .A(n6352), .B(n6353), .Z(N13313) );
  NANDN U8522 ( .A(n6354), .B(n6355), .Z(n6353) );
  OR U8523 ( .A(n6356), .B(n6357), .Z(n6355) );
  NAND U8524 ( .A(n6356), .B(n6357), .Z(n6352) );
  XOR U8525 ( .A(n6356), .B(n6358), .Z(N13312) );
  XNOR U8526 ( .A(n6354), .B(n6357), .Z(n6358) );
  AND U8527 ( .A(n6359), .B(n6360), .Z(n6357) );
  NANDN U8528 ( .A(n6361), .B(n6362), .Z(n6360) );
  NANDN U8529 ( .A(n6363), .B(n6364), .Z(n6362) );
  NANDN U8530 ( .A(n6364), .B(n6363), .Z(n6359) );
  NAND U8531 ( .A(n6365), .B(n6366), .Z(n6354) );
  NANDN U8532 ( .A(n6367), .B(n6368), .Z(n6366) );
  OR U8533 ( .A(n6369), .B(n6370), .Z(n6368) );
  NAND U8534 ( .A(n6370), .B(n6369), .Z(n6365) );
  AND U8535 ( .A(n6371), .B(n6372), .Z(n6356) );
  NANDN U8536 ( .A(n6373), .B(n6374), .Z(n6372) );
  NANDN U8537 ( .A(n6375), .B(n6376), .Z(n6374) );
  NANDN U8538 ( .A(n6376), .B(n6375), .Z(n6371) );
  XOR U8539 ( .A(n6370), .B(n6377), .Z(N13311) );
  XOR U8540 ( .A(n6367), .B(n6369), .Z(n6377) );
  XNOR U8541 ( .A(n6363), .B(n6378), .Z(n6369) );
  XNOR U8542 ( .A(n6361), .B(n6364), .Z(n6378) );
  NAND U8543 ( .A(n6379), .B(n6380), .Z(n6364) );
  NAND U8544 ( .A(n6381), .B(n6382), .Z(n6380) );
  OR U8545 ( .A(n6383), .B(n6384), .Z(n6381) );
  NANDN U8546 ( .A(n6385), .B(n6383), .Z(n6379) );
  IV U8547 ( .A(n6384), .Z(n6385) );
  NAND U8548 ( .A(n6386), .B(n6387), .Z(n6361) );
  NAND U8549 ( .A(n6388), .B(n6389), .Z(n6387) );
  NANDN U8550 ( .A(n6390), .B(n6391), .Z(n6388) );
  NANDN U8551 ( .A(n6391), .B(n6390), .Z(n6386) );
  AND U8552 ( .A(n6392), .B(n6393), .Z(n6363) );
  NAND U8553 ( .A(n6394), .B(n6395), .Z(n6393) );
  OR U8554 ( .A(n6396), .B(n6397), .Z(n6394) );
  NANDN U8555 ( .A(n6398), .B(n6396), .Z(n6392) );
  NAND U8556 ( .A(n6399), .B(n6400), .Z(n6367) );
  NANDN U8557 ( .A(n6401), .B(n6402), .Z(n6400) );
  OR U8558 ( .A(n6403), .B(n6404), .Z(n6402) );
  NANDN U8559 ( .A(n6405), .B(n6403), .Z(n6399) );
  IV U8560 ( .A(n6404), .Z(n6405) );
  XNOR U8561 ( .A(n6375), .B(n6406), .Z(n6370) );
  XNOR U8562 ( .A(n6373), .B(n6376), .Z(n6406) );
  NAND U8563 ( .A(n6407), .B(n6408), .Z(n6376) );
  NAND U8564 ( .A(n6409), .B(n6410), .Z(n6408) );
  OR U8565 ( .A(n6411), .B(n6412), .Z(n6409) );
  NANDN U8566 ( .A(n6413), .B(n6411), .Z(n6407) );
  IV U8567 ( .A(n6412), .Z(n6413) );
  NAND U8568 ( .A(n6414), .B(n6415), .Z(n6373) );
  NAND U8569 ( .A(n6416), .B(n6417), .Z(n6415) );
  NANDN U8570 ( .A(n6418), .B(n6419), .Z(n6416) );
  NANDN U8571 ( .A(n6419), .B(n6418), .Z(n6414) );
  AND U8572 ( .A(n6420), .B(n6421), .Z(n6375) );
  NAND U8573 ( .A(n6422), .B(n6423), .Z(n6421) );
  OR U8574 ( .A(n6424), .B(n6425), .Z(n6422) );
  NANDN U8575 ( .A(n6426), .B(n6424), .Z(n6420) );
  XNOR U8576 ( .A(n6401), .B(n6427), .Z(N13310) );
  XOR U8577 ( .A(n6403), .B(n6404), .Z(n6427) );
  XNOR U8578 ( .A(n6417), .B(n6428), .Z(n6404) );
  XOR U8579 ( .A(n6418), .B(n6419), .Z(n6428) );
  XOR U8580 ( .A(n6424), .B(n6429), .Z(n6419) );
  XOR U8581 ( .A(n6423), .B(n6426), .Z(n6429) );
  IV U8582 ( .A(n6425), .Z(n6426) );
  NAND U8583 ( .A(n6430), .B(n6431), .Z(n6425) );
  OR U8584 ( .A(n6432), .B(n6433), .Z(n6431) );
  OR U8585 ( .A(n6434), .B(n6435), .Z(n6430) );
  NAND U8586 ( .A(n6436), .B(n6437), .Z(n6423) );
  OR U8587 ( .A(n6438), .B(n6439), .Z(n6437) );
  OR U8588 ( .A(n6440), .B(n6441), .Z(n6436) );
  NOR U8589 ( .A(n6442), .B(n6443), .Z(n6424) );
  ANDN U8590 ( .B(n6444), .A(n6445), .Z(n6418) );
  XNOR U8591 ( .A(n6411), .B(n6446), .Z(n6417) );
  XNOR U8592 ( .A(n6410), .B(n6412), .Z(n6446) );
  NAND U8593 ( .A(n6447), .B(n6448), .Z(n6412) );
  OR U8594 ( .A(n6449), .B(n6450), .Z(n6448) );
  OR U8595 ( .A(n6451), .B(n6452), .Z(n6447) );
  NAND U8596 ( .A(n6453), .B(n6454), .Z(n6410) );
  OR U8597 ( .A(n6455), .B(n6456), .Z(n6454) );
  OR U8598 ( .A(n6457), .B(n6458), .Z(n6453) );
  ANDN U8599 ( .B(n6459), .A(n6460), .Z(n6411) );
  IV U8600 ( .A(n6461), .Z(n6459) );
  ANDN U8601 ( .B(n6462), .A(n6463), .Z(n6403) );
  XOR U8602 ( .A(n6389), .B(n6464), .Z(n6401) );
  XOR U8603 ( .A(n6390), .B(n6391), .Z(n6464) );
  XOR U8604 ( .A(n6396), .B(n6465), .Z(n6391) );
  XOR U8605 ( .A(n6395), .B(n6398), .Z(n6465) );
  IV U8606 ( .A(n6397), .Z(n6398) );
  NAND U8607 ( .A(n6466), .B(n6467), .Z(n6397) );
  OR U8608 ( .A(n6468), .B(n6469), .Z(n6467) );
  OR U8609 ( .A(n6470), .B(n6471), .Z(n6466) );
  NAND U8610 ( .A(n6472), .B(n6473), .Z(n6395) );
  OR U8611 ( .A(n6474), .B(n6475), .Z(n6473) );
  OR U8612 ( .A(n6476), .B(n6477), .Z(n6472) );
  NOR U8613 ( .A(n6478), .B(n6479), .Z(n6396) );
  ANDN U8614 ( .B(n6480), .A(n6481), .Z(n6390) );
  IV U8615 ( .A(n6482), .Z(n6480) );
  XNOR U8616 ( .A(n6383), .B(n6483), .Z(n6389) );
  XNOR U8617 ( .A(n6382), .B(n6384), .Z(n6483) );
  NAND U8618 ( .A(n6484), .B(n6485), .Z(n6384) );
  OR U8619 ( .A(n6486), .B(n6487), .Z(n6485) );
  OR U8620 ( .A(n6488), .B(n6489), .Z(n6484) );
  NAND U8621 ( .A(n6490), .B(n6491), .Z(n6382) );
  OR U8622 ( .A(n6492), .B(n6493), .Z(n6491) );
  OR U8623 ( .A(n6494), .B(n6495), .Z(n6490) );
  ANDN U8624 ( .B(n6496), .A(n6497), .Z(n6383) );
  IV U8625 ( .A(n6498), .Z(n6496) );
  XNOR U8626 ( .A(n6463), .B(n6462), .Z(N13309) );
  XOR U8627 ( .A(n6482), .B(n6481), .Z(n6462) );
  XNOR U8628 ( .A(n6497), .B(n6498), .Z(n6481) );
  XNOR U8629 ( .A(n6492), .B(n6493), .Z(n6498) );
  XNOR U8630 ( .A(n6494), .B(n6495), .Z(n6493) );
  XNOR U8631 ( .A(y[1165]), .B(x[1165]), .Z(n6495) );
  XNOR U8632 ( .A(y[1166]), .B(x[1166]), .Z(n6494) );
  XNOR U8633 ( .A(y[1164]), .B(x[1164]), .Z(n6492) );
  XNOR U8634 ( .A(n6486), .B(n6487), .Z(n6497) );
  XNOR U8635 ( .A(y[1161]), .B(x[1161]), .Z(n6487) );
  XNOR U8636 ( .A(n6488), .B(n6489), .Z(n6486) );
  XNOR U8637 ( .A(y[1162]), .B(x[1162]), .Z(n6489) );
  XNOR U8638 ( .A(y[1163]), .B(x[1163]), .Z(n6488) );
  XNOR U8639 ( .A(n6479), .B(n6478), .Z(n6482) );
  XNOR U8640 ( .A(n6474), .B(n6475), .Z(n6478) );
  XNOR U8641 ( .A(y[1158]), .B(x[1158]), .Z(n6475) );
  XNOR U8642 ( .A(n6476), .B(n6477), .Z(n6474) );
  XNOR U8643 ( .A(y[1159]), .B(x[1159]), .Z(n6477) );
  XNOR U8644 ( .A(y[1160]), .B(x[1160]), .Z(n6476) );
  XNOR U8645 ( .A(n6468), .B(n6469), .Z(n6479) );
  XNOR U8646 ( .A(y[1155]), .B(x[1155]), .Z(n6469) );
  XNOR U8647 ( .A(n6470), .B(n6471), .Z(n6468) );
  XNOR U8648 ( .A(y[1156]), .B(x[1156]), .Z(n6471) );
  XNOR U8649 ( .A(y[1157]), .B(x[1157]), .Z(n6470) );
  XOR U8650 ( .A(n6444), .B(n6445), .Z(n6463) );
  XNOR U8651 ( .A(n6460), .B(n6461), .Z(n6445) );
  XNOR U8652 ( .A(n6455), .B(n6456), .Z(n6461) );
  XNOR U8653 ( .A(n6457), .B(n6458), .Z(n6456) );
  XNOR U8654 ( .A(y[1153]), .B(x[1153]), .Z(n6458) );
  XNOR U8655 ( .A(y[1154]), .B(x[1154]), .Z(n6457) );
  XNOR U8656 ( .A(y[1152]), .B(x[1152]), .Z(n6455) );
  XNOR U8657 ( .A(n6449), .B(n6450), .Z(n6460) );
  XNOR U8658 ( .A(y[1149]), .B(x[1149]), .Z(n6450) );
  XNOR U8659 ( .A(n6451), .B(n6452), .Z(n6449) );
  XNOR U8660 ( .A(y[1150]), .B(x[1150]), .Z(n6452) );
  XNOR U8661 ( .A(y[1151]), .B(x[1151]), .Z(n6451) );
  XOR U8662 ( .A(n6443), .B(n6442), .Z(n6444) );
  XNOR U8663 ( .A(n6438), .B(n6439), .Z(n6442) );
  XNOR U8664 ( .A(y[1146]), .B(x[1146]), .Z(n6439) );
  XNOR U8665 ( .A(n6440), .B(n6441), .Z(n6438) );
  XNOR U8666 ( .A(y[1147]), .B(x[1147]), .Z(n6441) );
  XNOR U8667 ( .A(y[1148]), .B(x[1148]), .Z(n6440) );
  XNOR U8668 ( .A(n6432), .B(n6433), .Z(n6443) );
  XNOR U8669 ( .A(y[1143]), .B(x[1143]), .Z(n6433) );
  XNOR U8670 ( .A(n6434), .B(n6435), .Z(n6432) );
  XNOR U8671 ( .A(y[1144]), .B(x[1144]), .Z(n6435) );
  XNOR U8672 ( .A(y[1145]), .B(x[1145]), .Z(n6434) );
  NAND U8673 ( .A(n6499), .B(n6500), .Z(N13302) );
  NANDN U8674 ( .A(n6501), .B(n6502), .Z(n6500) );
  OR U8675 ( .A(n6503), .B(n6504), .Z(n6502) );
  NAND U8676 ( .A(n6503), .B(n6504), .Z(n6499) );
  XOR U8677 ( .A(n6503), .B(n6505), .Z(N13301) );
  XNOR U8678 ( .A(n6501), .B(n6504), .Z(n6505) );
  AND U8679 ( .A(n6506), .B(n6507), .Z(n6504) );
  NANDN U8680 ( .A(n6508), .B(n6509), .Z(n6507) );
  NANDN U8681 ( .A(n6510), .B(n6511), .Z(n6509) );
  NANDN U8682 ( .A(n6511), .B(n6510), .Z(n6506) );
  NAND U8683 ( .A(n6512), .B(n6513), .Z(n6501) );
  NANDN U8684 ( .A(n6514), .B(n6515), .Z(n6513) );
  OR U8685 ( .A(n6516), .B(n6517), .Z(n6515) );
  NAND U8686 ( .A(n6517), .B(n6516), .Z(n6512) );
  AND U8687 ( .A(n6518), .B(n6519), .Z(n6503) );
  NANDN U8688 ( .A(n6520), .B(n6521), .Z(n6519) );
  NANDN U8689 ( .A(n6522), .B(n6523), .Z(n6521) );
  NANDN U8690 ( .A(n6523), .B(n6522), .Z(n6518) );
  XOR U8691 ( .A(n6517), .B(n6524), .Z(N13300) );
  XOR U8692 ( .A(n6514), .B(n6516), .Z(n6524) );
  XNOR U8693 ( .A(n6510), .B(n6525), .Z(n6516) );
  XNOR U8694 ( .A(n6508), .B(n6511), .Z(n6525) );
  NAND U8695 ( .A(n6526), .B(n6527), .Z(n6511) );
  NAND U8696 ( .A(n6528), .B(n6529), .Z(n6527) );
  OR U8697 ( .A(n6530), .B(n6531), .Z(n6528) );
  NANDN U8698 ( .A(n6532), .B(n6530), .Z(n6526) );
  IV U8699 ( .A(n6531), .Z(n6532) );
  NAND U8700 ( .A(n6533), .B(n6534), .Z(n6508) );
  NAND U8701 ( .A(n6535), .B(n6536), .Z(n6534) );
  NANDN U8702 ( .A(n6537), .B(n6538), .Z(n6535) );
  NANDN U8703 ( .A(n6538), .B(n6537), .Z(n6533) );
  AND U8704 ( .A(n6539), .B(n6540), .Z(n6510) );
  NAND U8705 ( .A(n6541), .B(n6542), .Z(n6540) );
  OR U8706 ( .A(n6543), .B(n6544), .Z(n6541) );
  NANDN U8707 ( .A(n6545), .B(n6543), .Z(n6539) );
  NAND U8708 ( .A(n6546), .B(n6547), .Z(n6514) );
  NANDN U8709 ( .A(n6548), .B(n6549), .Z(n6547) );
  OR U8710 ( .A(n6550), .B(n6551), .Z(n6549) );
  NANDN U8711 ( .A(n6552), .B(n6550), .Z(n6546) );
  IV U8712 ( .A(n6551), .Z(n6552) );
  XNOR U8713 ( .A(n6522), .B(n6553), .Z(n6517) );
  XNOR U8714 ( .A(n6520), .B(n6523), .Z(n6553) );
  NAND U8715 ( .A(n6554), .B(n6555), .Z(n6523) );
  NAND U8716 ( .A(n6556), .B(n6557), .Z(n6555) );
  OR U8717 ( .A(n6558), .B(n6559), .Z(n6556) );
  NANDN U8718 ( .A(n6560), .B(n6558), .Z(n6554) );
  IV U8719 ( .A(n6559), .Z(n6560) );
  NAND U8720 ( .A(n6561), .B(n6562), .Z(n6520) );
  NAND U8721 ( .A(n6563), .B(n6564), .Z(n6562) );
  NANDN U8722 ( .A(n6565), .B(n6566), .Z(n6563) );
  NANDN U8723 ( .A(n6566), .B(n6565), .Z(n6561) );
  AND U8724 ( .A(n6567), .B(n6568), .Z(n6522) );
  NAND U8725 ( .A(n6569), .B(n6570), .Z(n6568) );
  OR U8726 ( .A(n6571), .B(n6572), .Z(n6569) );
  NANDN U8727 ( .A(n6573), .B(n6571), .Z(n6567) );
  XNOR U8728 ( .A(n6548), .B(n6574), .Z(N13299) );
  XOR U8729 ( .A(n6550), .B(n6551), .Z(n6574) );
  XNOR U8730 ( .A(n6564), .B(n6575), .Z(n6551) );
  XOR U8731 ( .A(n6565), .B(n6566), .Z(n6575) );
  XOR U8732 ( .A(n6571), .B(n6576), .Z(n6566) );
  XOR U8733 ( .A(n6570), .B(n6573), .Z(n6576) );
  IV U8734 ( .A(n6572), .Z(n6573) );
  NAND U8735 ( .A(n6577), .B(n6578), .Z(n6572) );
  OR U8736 ( .A(n6579), .B(n6580), .Z(n6578) );
  OR U8737 ( .A(n6581), .B(n6582), .Z(n6577) );
  NAND U8738 ( .A(n6583), .B(n6584), .Z(n6570) );
  OR U8739 ( .A(n6585), .B(n6586), .Z(n6584) );
  OR U8740 ( .A(n6587), .B(n6588), .Z(n6583) );
  NOR U8741 ( .A(n6589), .B(n6590), .Z(n6571) );
  ANDN U8742 ( .B(n6591), .A(n6592), .Z(n6565) );
  XNOR U8743 ( .A(n6558), .B(n6593), .Z(n6564) );
  XNOR U8744 ( .A(n6557), .B(n6559), .Z(n6593) );
  NAND U8745 ( .A(n6594), .B(n6595), .Z(n6559) );
  OR U8746 ( .A(n6596), .B(n6597), .Z(n6595) );
  OR U8747 ( .A(n6598), .B(n6599), .Z(n6594) );
  NAND U8748 ( .A(n6600), .B(n6601), .Z(n6557) );
  OR U8749 ( .A(n6602), .B(n6603), .Z(n6601) );
  OR U8750 ( .A(n6604), .B(n6605), .Z(n6600) );
  ANDN U8751 ( .B(n6606), .A(n6607), .Z(n6558) );
  IV U8752 ( .A(n6608), .Z(n6606) );
  ANDN U8753 ( .B(n6609), .A(n6610), .Z(n6550) );
  XOR U8754 ( .A(n6536), .B(n6611), .Z(n6548) );
  XOR U8755 ( .A(n6537), .B(n6538), .Z(n6611) );
  XOR U8756 ( .A(n6543), .B(n6612), .Z(n6538) );
  XOR U8757 ( .A(n6542), .B(n6545), .Z(n6612) );
  IV U8758 ( .A(n6544), .Z(n6545) );
  NAND U8759 ( .A(n6613), .B(n6614), .Z(n6544) );
  OR U8760 ( .A(n6615), .B(n6616), .Z(n6614) );
  OR U8761 ( .A(n6617), .B(n6618), .Z(n6613) );
  NAND U8762 ( .A(n6619), .B(n6620), .Z(n6542) );
  OR U8763 ( .A(n6621), .B(n6622), .Z(n6620) );
  OR U8764 ( .A(n6623), .B(n6624), .Z(n6619) );
  NOR U8765 ( .A(n6625), .B(n6626), .Z(n6543) );
  ANDN U8766 ( .B(n6627), .A(n6628), .Z(n6537) );
  IV U8767 ( .A(n6629), .Z(n6627) );
  XNOR U8768 ( .A(n6530), .B(n6630), .Z(n6536) );
  XNOR U8769 ( .A(n6529), .B(n6531), .Z(n6630) );
  NAND U8770 ( .A(n6631), .B(n6632), .Z(n6531) );
  OR U8771 ( .A(n6633), .B(n6634), .Z(n6632) );
  OR U8772 ( .A(n6635), .B(n6636), .Z(n6631) );
  NAND U8773 ( .A(n6637), .B(n6638), .Z(n6529) );
  OR U8774 ( .A(n6639), .B(n6640), .Z(n6638) );
  OR U8775 ( .A(n6641), .B(n6642), .Z(n6637) );
  ANDN U8776 ( .B(n6643), .A(n6644), .Z(n6530) );
  IV U8777 ( .A(n6645), .Z(n6643) );
  XNOR U8778 ( .A(n6610), .B(n6609), .Z(N13298) );
  XOR U8779 ( .A(n6629), .B(n6628), .Z(n6609) );
  XNOR U8780 ( .A(n6644), .B(n6645), .Z(n6628) );
  XNOR U8781 ( .A(n6639), .B(n6640), .Z(n6645) );
  XNOR U8782 ( .A(n6641), .B(n6642), .Z(n6640) );
  XNOR U8783 ( .A(y[1141]), .B(x[1141]), .Z(n6642) );
  XNOR U8784 ( .A(y[1142]), .B(x[1142]), .Z(n6641) );
  XNOR U8785 ( .A(y[1140]), .B(x[1140]), .Z(n6639) );
  XNOR U8786 ( .A(n6633), .B(n6634), .Z(n6644) );
  XNOR U8787 ( .A(y[1137]), .B(x[1137]), .Z(n6634) );
  XNOR U8788 ( .A(n6635), .B(n6636), .Z(n6633) );
  XNOR U8789 ( .A(y[1138]), .B(x[1138]), .Z(n6636) );
  XNOR U8790 ( .A(y[1139]), .B(x[1139]), .Z(n6635) );
  XNOR U8791 ( .A(n6626), .B(n6625), .Z(n6629) );
  XNOR U8792 ( .A(n6621), .B(n6622), .Z(n6625) );
  XNOR U8793 ( .A(y[1134]), .B(x[1134]), .Z(n6622) );
  XNOR U8794 ( .A(n6623), .B(n6624), .Z(n6621) );
  XNOR U8795 ( .A(y[1135]), .B(x[1135]), .Z(n6624) );
  XNOR U8796 ( .A(y[1136]), .B(x[1136]), .Z(n6623) );
  XNOR U8797 ( .A(n6615), .B(n6616), .Z(n6626) );
  XNOR U8798 ( .A(y[1131]), .B(x[1131]), .Z(n6616) );
  XNOR U8799 ( .A(n6617), .B(n6618), .Z(n6615) );
  XNOR U8800 ( .A(y[1132]), .B(x[1132]), .Z(n6618) );
  XNOR U8801 ( .A(y[1133]), .B(x[1133]), .Z(n6617) );
  XOR U8802 ( .A(n6591), .B(n6592), .Z(n6610) );
  XNOR U8803 ( .A(n6607), .B(n6608), .Z(n6592) );
  XNOR U8804 ( .A(n6602), .B(n6603), .Z(n6608) );
  XNOR U8805 ( .A(n6604), .B(n6605), .Z(n6603) );
  XNOR U8806 ( .A(y[1129]), .B(x[1129]), .Z(n6605) );
  XNOR U8807 ( .A(y[1130]), .B(x[1130]), .Z(n6604) );
  XNOR U8808 ( .A(y[1128]), .B(x[1128]), .Z(n6602) );
  XNOR U8809 ( .A(n6596), .B(n6597), .Z(n6607) );
  XNOR U8810 ( .A(y[1125]), .B(x[1125]), .Z(n6597) );
  XNOR U8811 ( .A(n6598), .B(n6599), .Z(n6596) );
  XNOR U8812 ( .A(y[1126]), .B(x[1126]), .Z(n6599) );
  XNOR U8813 ( .A(y[1127]), .B(x[1127]), .Z(n6598) );
  XOR U8814 ( .A(n6590), .B(n6589), .Z(n6591) );
  XNOR U8815 ( .A(n6585), .B(n6586), .Z(n6589) );
  XNOR U8816 ( .A(y[1122]), .B(x[1122]), .Z(n6586) );
  XNOR U8817 ( .A(n6587), .B(n6588), .Z(n6585) );
  XNOR U8818 ( .A(y[1123]), .B(x[1123]), .Z(n6588) );
  XNOR U8819 ( .A(y[1124]), .B(x[1124]), .Z(n6587) );
  XNOR U8820 ( .A(n6579), .B(n6580), .Z(n6590) );
  XNOR U8821 ( .A(y[1119]), .B(x[1119]), .Z(n6580) );
  XNOR U8822 ( .A(n6581), .B(n6582), .Z(n6579) );
  XNOR U8823 ( .A(y[1120]), .B(x[1120]), .Z(n6582) );
  XNOR U8824 ( .A(y[1121]), .B(x[1121]), .Z(n6581) );
  NAND U8825 ( .A(n6646), .B(n6647), .Z(N13291) );
  NANDN U8826 ( .A(n6648), .B(n6649), .Z(n6647) );
  OR U8827 ( .A(n6650), .B(n6651), .Z(n6649) );
  NAND U8828 ( .A(n6650), .B(n6651), .Z(n6646) );
  XOR U8829 ( .A(n6650), .B(n6652), .Z(N13290) );
  XNOR U8830 ( .A(n6648), .B(n6651), .Z(n6652) );
  AND U8831 ( .A(n6653), .B(n6654), .Z(n6651) );
  NANDN U8832 ( .A(n6655), .B(n6656), .Z(n6654) );
  NANDN U8833 ( .A(n6657), .B(n6658), .Z(n6656) );
  NANDN U8834 ( .A(n6658), .B(n6657), .Z(n6653) );
  NAND U8835 ( .A(n6659), .B(n6660), .Z(n6648) );
  NANDN U8836 ( .A(n6661), .B(n6662), .Z(n6660) );
  OR U8837 ( .A(n6663), .B(n6664), .Z(n6662) );
  NAND U8838 ( .A(n6664), .B(n6663), .Z(n6659) );
  AND U8839 ( .A(n6665), .B(n6666), .Z(n6650) );
  NANDN U8840 ( .A(n6667), .B(n6668), .Z(n6666) );
  NANDN U8841 ( .A(n6669), .B(n6670), .Z(n6668) );
  NANDN U8842 ( .A(n6670), .B(n6669), .Z(n6665) );
  XOR U8843 ( .A(n6664), .B(n6671), .Z(N13289) );
  XOR U8844 ( .A(n6661), .B(n6663), .Z(n6671) );
  XNOR U8845 ( .A(n6657), .B(n6672), .Z(n6663) );
  XNOR U8846 ( .A(n6655), .B(n6658), .Z(n6672) );
  NAND U8847 ( .A(n6673), .B(n6674), .Z(n6658) );
  NAND U8848 ( .A(n6675), .B(n6676), .Z(n6674) );
  OR U8849 ( .A(n6677), .B(n6678), .Z(n6675) );
  NANDN U8850 ( .A(n6679), .B(n6677), .Z(n6673) );
  IV U8851 ( .A(n6678), .Z(n6679) );
  NAND U8852 ( .A(n6680), .B(n6681), .Z(n6655) );
  NAND U8853 ( .A(n6682), .B(n6683), .Z(n6681) );
  NANDN U8854 ( .A(n6684), .B(n6685), .Z(n6682) );
  NANDN U8855 ( .A(n6685), .B(n6684), .Z(n6680) );
  AND U8856 ( .A(n6686), .B(n6687), .Z(n6657) );
  NAND U8857 ( .A(n6688), .B(n6689), .Z(n6687) );
  OR U8858 ( .A(n6690), .B(n6691), .Z(n6688) );
  NANDN U8859 ( .A(n6692), .B(n6690), .Z(n6686) );
  NAND U8860 ( .A(n6693), .B(n6694), .Z(n6661) );
  NANDN U8861 ( .A(n6695), .B(n6696), .Z(n6694) );
  OR U8862 ( .A(n6697), .B(n6698), .Z(n6696) );
  NANDN U8863 ( .A(n6699), .B(n6697), .Z(n6693) );
  IV U8864 ( .A(n6698), .Z(n6699) );
  XNOR U8865 ( .A(n6669), .B(n6700), .Z(n6664) );
  XNOR U8866 ( .A(n6667), .B(n6670), .Z(n6700) );
  NAND U8867 ( .A(n6701), .B(n6702), .Z(n6670) );
  NAND U8868 ( .A(n6703), .B(n6704), .Z(n6702) );
  OR U8869 ( .A(n6705), .B(n6706), .Z(n6703) );
  NANDN U8870 ( .A(n6707), .B(n6705), .Z(n6701) );
  IV U8871 ( .A(n6706), .Z(n6707) );
  NAND U8872 ( .A(n6708), .B(n6709), .Z(n6667) );
  NAND U8873 ( .A(n6710), .B(n6711), .Z(n6709) );
  NANDN U8874 ( .A(n6712), .B(n6713), .Z(n6710) );
  NANDN U8875 ( .A(n6713), .B(n6712), .Z(n6708) );
  AND U8876 ( .A(n6714), .B(n6715), .Z(n6669) );
  NAND U8877 ( .A(n6716), .B(n6717), .Z(n6715) );
  OR U8878 ( .A(n6718), .B(n6719), .Z(n6716) );
  NANDN U8879 ( .A(n6720), .B(n6718), .Z(n6714) );
  XNOR U8880 ( .A(n6695), .B(n6721), .Z(N13288) );
  XOR U8881 ( .A(n6697), .B(n6698), .Z(n6721) );
  XNOR U8882 ( .A(n6711), .B(n6722), .Z(n6698) );
  XOR U8883 ( .A(n6712), .B(n6713), .Z(n6722) );
  XOR U8884 ( .A(n6718), .B(n6723), .Z(n6713) );
  XOR U8885 ( .A(n6717), .B(n6720), .Z(n6723) );
  IV U8886 ( .A(n6719), .Z(n6720) );
  NAND U8887 ( .A(n6724), .B(n6725), .Z(n6719) );
  OR U8888 ( .A(n6726), .B(n6727), .Z(n6725) );
  OR U8889 ( .A(n6728), .B(n6729), .Z(n6724) );
  NAND U8890 ( .A(n6730), .B(n6731), .Z(n6717) );
  OR U8891 ( .A(n6732), .B(n6733), .Z(n6731) );
  OR U8892 ( .A(n6734), .B(n6735), .Z(n6730) );
  NOR U8893 ( .A(n6736), .B(n6737), .Z(n6718) );
  ANDN U8894 ( .B(n6738), .A(n6739), .Z(n6712) );
  XNOR U8895 ( .A(n6705), .B(n6740), .Z(n6711) );
  XNOR U8896 ( .A(n6704), .B(n6706), .Z(n6740) );
  NAND U8897 ( .A(n6741), .B(n6742), .Z(n6706) );
  OR U8898 ( .A(n6743), .B(n6744), .Z(n6742) );
  OR U8899 ( .A(n6745), .B(n6746), .Z(n6741) );
  NAND U8900 ( .A(n6747), .B(n6748), .Z(n6704) );
  OR U8901 ( .A(n6749), .B(n6750), .Z(n6748) );
  OR U8902 ( .A(n6751), .B(n6752), .Z(n6747) );
  ANDN U8903 ( .B(n6753), .A(n6754), .Z(n6705) );
  IV U8904 ( .A(n6755), .Z(n6753) );
  ANDN U8905 ( .B(n6756), .A(n6757), .Z(n6697) );
  XOR U8906 ( .A(n6683), .B(n6758), .Z(n6695) );
  XOR U8907 ( .A(n6684), .B(n6685), .Z(n6758) );
  XOR U8908 ( .A(n6690), .B(n6759), .Z(n6685) );
  XOR U8909 ( .A(n6689), .B(n6692), .Z(n6759) );
  IV U8910 ( .A(n6691), .Z(n6692) );
  NAND U8911 ( .A(n6760), .B(n6761), .Z(n6691) );
  OR U8912 ( .A(n6762), .B(n6763), .Z(n6761) );
  OR U8913 ( .A(n6764), .B(n6765), .Z(n6760) );
  NAND U8914 ( .A(n6766), .B(n6767), .Z(n6689) );
  OR U8915 ( .A(n6768), .B(n6769), .Z(n6767) );
  OR U8916 ( .A(n6770), .B(n6771), .Z(n6766) );
  NOR U8917 ( .A(n6772), .B(n6773), .Z(n6690) );
  ANDN U8918 ( .B(n6774), .A(n6775), .Z(n6684) );
  IV U8919 ( .A(n6776), .Z(n6774) );
  XNOR U8920 ( .A(n6677), .B(n6777), .Z(n6683) );
  XNOR U8921 ( .A(n6676), .B(n6678), .Z(n6777) );
  NAND U8922 ( .A(n6778), .B(n6779), .Z(n6678) );
  OR U8923 ( .A(n6780), .B(n6781), .Z(n6779) );
  OR U8924 ( .A(n6782), .B(n6783), .Z(n6778) );
  NAND U8925 ( .A(n6784), .B(n6785), .Z(n6676) );
  OR U8926 ( .A(n6786), .B(n6787), .Z(n6785) );
  OR U8927 ( .A(n6788), .B(n6789), .Z(n6784) );
  ANDN U8928 ( .B(n6790), .A(n6791), .Z(n6677) );
  IV U8929 ( .A(n6792), .Z(n6790) );
  XNOR U8930 ( .A(n6757), .B(n6756), .Z(N13287) );
  XOR U8931 ( .A(n6776), .B(n6775), .Z(n6756) );
  XNOR U8932 ( .A(n6791), .B(n6792), .Z(n6775) );
  XNOR U8933 ( .A(n6786), .B(n6787), .Z(n6792) );
  XNOR U8934 ( .A(n6788), .B(n6789), .Z(n6787) );
  XNOR U8935 ( .A(y[1117]), .B(x[1117]), .Z(n6789) );
  XNOR U8936 ( .A(y[1118]), .B(x[1118]), .Z(n6788) );
  XNOR U8937 ( .A(y[1116]), .B(x[1116]), .Z(n6786) );
  XNOR U8938 ( .A(n6780), .B(n6781), .Z(n6791) );
  XNOR U8939 ( .A(y[1113]), .B(x[1113]), .Z(n6781) );
  XNOR U8940 ( .A(n6782), .B(n6783), .Z(n6780) );
  XNOR U8941 ( .A(y[1114]), .B(x[1114]), .Z(n6783) );
  XNOR U8942 ( .A(y[1115]), .B(x[1115]), .Z(n6782) );
  XNOR U8943 ( .A(n6773), .B(n6772), .Z(n6776) );
  XNOR U8944 ( .A(n6768), .B(n6769), .Z(n6772) );
  XNOR U8945 ( .A(y[1110]), .B(x[1110]), .Z(n6769) );
  XNOR U8946 ( .A(n6770), .B(n6771), .Z(n6768) );
  XNOR U8947 ( .A(y[1111]), .B(x[1111]), .Z(n6771) );
  XNOR U8948 ( .A(y[1112]), .B(x[1112]), .Z(n6770) );
  XNOR U8949 ( .A(n6762), .B(n6763), .Z(n6773) );
  XNOR U8950 ( .A(y[1107]), .B(x[1107]), .Z(n6763) );
  XNOR U8951 ( .A(n6764), .B(n6765), .Z(n6762) );
  XNOR U8952 ( .A(y[1108]), .B(x[1108]), .Z(n6765) );
  XNOR U8953 ( .A(y[1109]), .B(x[1109]), .Z(n6764) );
  XOR U8954 ( .A(n6738), .B(n6739), .Z(n6757) );
  XNOR U8955 ( .A(n6754), .B(n6755), .Z(n6739) );
  XNOR U8956 ( .A(n6749), .B(n6750), .Z(n6755) );
  XNOR U8957 ( .A(n6751), .B(n6752), .Z(n6750) );
  XNOR U8958 ( .A(y[1105]), .B(x[1105]), .Z(n6752) );
  XNOR U8959 ( .A(y[1106]), .B(x[1106]), .Z(n6751) );
  XNOR U8960 ( .A(y[1104]), .B(x[1104]), .Z(n6749) );
  XNOR U8961 ( .A(n6743), .B(n6744), .Z(n6754) );
  XNOR U8962 ( .A(y[1101]), .B(x[1101]), .Z(n6744) );
  XNOR U8963 ( .A(n6745), .B(n6746), .Z(n6743) );
  XNOR U8964 ( .A(y[1102]), .B(x[1102]), .Z(n6746) );
  XNOR U8965 ( .A(y[1103]), .B(x[1103]), .Z(n6745) );
  XOR U8966 ( .A(n6737), .B(n6736), .Z(n6738) );
  XNOR U8967 ( .A(n6732), .B(n6733), .Z(n6736) );
  XNOR U8968 ( .A(y[1098]), .B(x[1098]), .Z(n6733) );
  XNOR U8969 ( .A(n6734), .B(n6735), .Z(n6732) );
  XNOR U8970 ( .A(y[1099]), .B(x[1099]), .Z(n6735) );
  XNOR U8971 ( .A(y[1100]), .B(x[1100]), .Z(n6734) );
  XNOR U8972 ( .A(n6726), .B(n6727), .Z(n6737) );
  XNOR U8973 ( .A(y[1095]), .B(x[1095]), .Z(n6727) );
  XNOR U8974 ( .A(n6728), .B(n6729), .Z(n6726) );
  XNOR U8975 ( .A(y[1096]), .B(x[1096]), .Z(n6729) );
  XNOR U8976 ( .A(y[1097]), .B(x[1097]), .Z(n6728) );
  NAND U8977 ( .A(n6793), .B(n6794), .Z(N13280) );
  NANDN U8978 ( .A(n6795), .B(n6796), .Z(n6794) );
  OR U8979 ( .A(n6797), .B(n6798), .Z(n6796) );
  NAND U8980 ( .A(n6797), .B(n6798), .Z(n6793) );
  XOR U8981 ( .A(n6797), .B(n6799), .Z(N13279) );
  XNOR U8982 ( .A(n6795), .B(n6798), .Z(n6799) );
  AND U8983 ( .A(n6800), .B(n6801), .Z(n6798) );
  NANDN U8984 ( .A(n6802), .B(n6803), .Z(n6801) );
  NANDN U8985 ( .A(n6804), .B(n6805), .Z(n6803) );
  NANDN U8986 ( .A(n6805), .B(n6804), .Z(n6800) );
  NAND U8987 ( .A(n6806), .B(n6807), .Z(n6795) );
  NANDN U8988 ( .A(n6808), .B(n6809), .Z(n6807) );
  OR U8989 ( .A(n6810), .B(n6811), .Z(n6809) );
  NAND U8990 ( .A(n6811), .B(n6810), .Z(n6806) );
  AND U8991 ( .A(n6812), .B(n6813), .Z(n6797) );
  NANDN U8992 ( .A(n6814), .B(n6815), .Z(n6813) );
  NANDN U8993 ( .A(n6816), .B(n6817), .Z(n6815) );
  NANDN U8994 ( .A(n6817), .B(n6816), .Z(n6812) );
  XOR U8995 ( .A(n6811), .B(n6818), .Z(N13278) );
  XOR U8996 ( .A(n6808), .B(n6810), .Z(n6818) );
  XNOR U8997 ( .A(n6804), .B(n6819), .Z(n6810) );
  XNOR U8998 ( .A(n6802), .B(n6805), .Z(n6819) );
  NAND U8999 ( .A(n6820), .B(n6821), .Z(n6805) );
  NAND U9000 ( .A(n6822), .B(n6823), .Z(n6821) );
  OR U9001 ( .A(n6824), .B(n6825), .Z(n6822) );
  NANDN U9002 ( .A(n6826), .B(n6824), .Z(n6820) );
  IV U9003 ( .A(n6825), .Z(n6826) );
  NAND U9004 ( .A(n6827), .B(n6828), .Z(n6802) );
  NAND U9005 ( .A(n6829), .B(n6830), .Z(n6828) );
  NANDN U9006 ( .A(n6831), .B(n6832), .Z(n6829) );
  NANDN U9007 ( .A(n6832), .B(n6831), .Z(n6827) );
  AND U9008 ( .A(n6833), .B(n6834), .Z(n6804) );
  NAND U9009 ( .A(n6835), .B(n6836), .Z(n6834) );
  OR U9010 ( .A(n6837), .B(n6838), .Z(n6835) );
  NANDN U9011 ( .A(n6839), .B(n6837), .Z(n6833) );
  NAND U9012 ( .A(n6840), .B(n6841), .Z(n6808) );
  NANDN U9013 ( .A(n6842), .B(n6843), .Z(n6841) );
  OR U9014 ( .A(n6844), .B(n6845), .Z(n6843) );
  NANDN U9015 ( .A(n6846), .B(n6844), .Z(n6840) );
  IV U9016 ( .A(n6845), .Z(n6846) );
  XNOR U9017 ( .A(n6816), .B(n6847), .Z(n6811) );
  XNOR U9018 ( .A(n6814), .B(n6817), .Z(n6847) );
  NAND U9019 ( .A(n6848), .B(n6849), .Z(n6817) );
  NAND U9020 ( .A(n6850), .B(n6851), .Z(n6849) );
  OR U9021 ( .A(n6852), .B(n6853), .Z(n6850) );
  NANDN U9022 ( .A(n6854), .B(n6852), .Z(n6848) );
  IV U9023 ( .A(n6853), .Z(n6854) );
  NAND U9024 ( .A(n6855), .B(n6856), .Z(n6814) );
  NAND U9025 ( .A(n6857), .B(n6858), .Z(n6856) );
  NANDN U9026 ( .A(n6859), .B(n6860), .Z(n6857) );
  NANDN U9027 ( .A(n6860), .B(n6859), .Z(n6855) );
  AND U9028 ( .A(n6861), .B(n6862), .Z(n6816) );
  NAND U9029 ( .A(n6863), .B(n6864), .Z(n6862) );
  OR U9030 ( .A(n6865), .B(n6866), .Z(n6863) );
  NANDN U9031 ( .A(n6867), .B(n6865), .Z(n6861) );
  XNOR U9032 ( .A(n6842), .B(n6868), .Z(N13277) );
  XOR U9033 ( .A(n6844), .B(n6845), .Z(n6868) );
  XNOR U9034 ( .A(n6858), .B(n6869), .Z(n6845) );
  XOR U9035 ( .A(n6859), .B(n6860), .Z(n6869) );
  XOR U9036 ( .A(n6865), .B(n6870), .Z(n6860) );
  XOR U9037 ( .A(n6864), .B(n6867), .Z(n6870) );
  IV U9038 ( .A(n6866), .Z(n6867) );
  NAND U9039 ( .A(n6871), .B(n6872), .Z(n6866) );
  OR U9040 ( .A(n6873), .B(n6874), .Z(n6872) );
  OR U9041 ( .A(n6875), .B(n6876), .Z(n6871) );
  NAND U9042 ( .A(n6877), .B(n6878), .Z(n6864) );
  OR U9043 ( .A(n6879), .B(n6880), .Z(n6878) );
  OR U9044 ( .A(n6881), .B(n6882), .Z(n6877) );
  NOR U9045 ( .A(n6883), .B(n6884), .Z(n6865) );
  ANDN U9046 ( .B(n6885), .A(n6886), .Z(n6859) );
  XNOR U9047 ( .A(n6852), .B(n6887), .Z(n6858) );
  XNOR U9048 ( .A(n6851), .B(n6853), .Z(n6887) );
  NAND U9049 ( .A(n6888), .B(n6889), .Z(n6853) );
  OR U9050 ( .A(n6890), .B(n6891), .Z(n6889) );
  OR U9051 ( .A(n6892), .B(n6893), .Z(n6888) );
  NAND U9052 ( .A(n6894), .B(n6895), .Z(n6851) );
  OR U9053 ( .A(n6896), .B(n6897), .Z(n6895) );
  OR U9054 ( .A(n6898), .B(n6899), .Z(n6894) );
  ANDN U9055 ( .B(n6900), .A(n6901), .Z(n6852) );
  IV U9056 ( .A(n6902), .Z(n6900) );
  ANDN U9057 ( .B(n6903), .A(n6904), .Z(n6844) );
  XOR U9058 ( .A(n6830), .B(n6905), .Z(n6842) );
  XOR U9059 ( .A(n6831), .B(n6832), .Z(n6905) );
  XOR U9060 ( .A(n6837), .B(n6906), .Z(n6832) );
  XOR U9061 ( .A(n6836), .B(n6839), .Z(n6906) );
  IV U9062 ( .A(n6838), .Z(n6839) );
  NAND U9063 ( .A(n6907), .B(n6908), .Z(n6838) );
  OR U9064 ( .A(n6909), .B(n6910), .Z(n6908) );
  OR U9065 ( .A(n6911), .B(n6912), .Z(n6907) );
  NAND U9066 ( .A(n6913), .B(n6914), .Z(n6836) );
  OR U9067 ( .A(n6915), .B(n6916), .Z(n6914) );
  OR U9068 ( .A(n6917), .B(n6918), .Z(n6913) );
  NOR U9069 ( .A(n6919), .B(n6920), .Z(n6837) );
  ANDN U9070 ( .B(n6921), .A(n6922), .Z(n6831) );
  IV U9071 ( .A(n6923), .Z(n6921) );
  XNOR U9072 ( .A(n6824), .B(n6924), .Z(n6830) );
  XNOR U9073 ( .A(n6823), .B(n6825), .Z(n6924) );
  NAND U9074 ( .A(n6925), .B(n6926), .Z(n6825) );
  OR U9075 ( .A(n6927), .B(n6928), .Z(n6926) );
  OR U9076 ( .A(n6929), .B(n6930), .Z(n6925) );
  NAND U9077 ( .A(n6931), .B(n6932), .Z(n6823) );
  OR U9078 ( .A(n6933), .B(n6934), .Z(n6932) );
  OR U9079 ( .A(n6935), .B(n6936), .Z(n6931) );
  ANDN U9080 ( .B(n6937), .A(n6938), .Z(n6824) );
  IV U9081 ( .A(n6939), .Z(n6937) );
  XNOR U9082 ( .A(n6904), .B(n6903), .Z(N13276) );
  XOR U9083 ( .A(n6923), .B(n6922), .Z(n6903) );
  XNOR U9084 ( .A(n6938), .B(n6939), .Z(n6922) );
  XNOR U9085 ( .A(n6933), .B(n6934), .Z(n6939) );
  XNOR U9086 ( .A(n6935), .B(n6936), .Z(n6934) );
  XNOR U9087 ( .A(y[1093]), .B(x[1093]), .Z(n6936) );
  XNOR U9088 ( .A(y[1094]), .B(x[1094]), .Z(n6935) );
  XNOR U9089 ( .A(y[1092]), .B(x[1092]), .Z(n6933) );
  XNOR U9090 ( .A(n6927), .B(n6928), .Z(n6938) );
  XNOR U9091 ( .A(y[1089]), .B(x[1089]), .Z(n6928) );
  XNOR U9092 ( .A(n6929), .B(n6930), .Z(n6927) );
  XNOR U9093 ( .A(y[1090]), .B(x[1090]), .Z(n6930) );
  XNOR U9094 ( .A(y[1091]), .B(x[1091]), .Z(n6929) );
  XNOR U9095 ( .A(n6920), .B(n6919), .Z(n6923) );
  XNOR U9096 ( .A(n6915), .B(n6916), .Z(n6919) );
  XNOR U9097 ( .A(y[1086]), .B(x[1086]), .Z(n6916) );
  XNOR U9098 ( .A(n6917), .B(n6918), .Z(n6915) );
  XNOR U9099 ( .A(y[1087]), .B(x[1087]), .Z(n6918) );
  XNOR U9100 ( .A(y[1088]), .B(x[1088]), .Z(n6917) );
  XNOR U9101 ( .A(n6909), .B(n6910), .Z(n6920) );
  XNOR U9102 ( .A(y[1083]), .B(x[1083]), .Z(n6910) );
  XNOR U9103 ( .A(n6911), .B(n6912), .Z(n6909) );
  XNOR U9104 ( .A(y[1084]), .B(x[1084]), .Z(n6912) );
  XNOR U9105 ( .A(y[1085]), .B(x[1085]), .Z(n6911) );
  XOR U9106 ( .A(n6885), .B(n6886), .Z(n6904) );
  XNOR U9107 ( .A(n6901), .B(n6902), .Z(n6886) );
  XNOR U9108 ( .A(n6896), .B(n6897), .Z(n6902) );
  XNOR U9109 ( .A(n6898), .B(n6899), .Z(n6897) );
  XNOR U9110 ( .A(y[1081]), .B(x[1081]), .Z(n6899) );
  XNOR U9111 ( .A(y[1082]), .B(x[1082]), .Z(n6898) );
  XNOR U9112 ( .A(y[1080]), .B(x[1080]), .Z(n6896) );
  XNOR U9113 ( .A(n6890), .B(n6891), .Z(n6901) );
  XNOR U9114 ( .A(y[1077]), .B(x[1077]), .Z(n6891) );
  XNOR U9115 ( .A(n6892), .B(n6893), .Z(n6890) );
  XNOR U9116 ( .A(y[1078]), .B(x[1078]), .Z(n6893) );
  XNOR U9117 ( .A(y[1079]), .B(x[1079]), .Z(n6892) );
  XOR U9118 ( .A(n6884), .B(n6883), .Z(n6885) );
  XNOR U9119 ( .A(n6879), .B(n6880), .Z(n6883) );
  XNOR U9120 ( .A(y[1074]), .B(x[1074]), .Z(n6880) );
  XNOR U9121 ( .A(n6881), .B(n6882), .Z(n6879) );
  XNOR U9122 ( .A(y[1075]), .B(x[1075]), .Z(n6882) );
  XNOR U9123 ( .A(y[1076]), .B(x[1076]), .Z(n6881) );
  XNOR U9124 ( .A(n6873), .B(n6874), .Z(n6884) );
  XNOR U9125 ( .A(y[1071]), .B(x[1071]), .Z(n6874) );
  XNOR U9126 ( .A(n6875), .B(n6876), .Z(n6873) );
  XNOR U9127 ( .A(y[1072]), .B(x[1072]), .Z(n6876) );
  XNOR U9128 ( .A(y[1073]), .B(x[1073]), .Z(n6875) );
  NAND U9129 ( .A(n6940), .B(n6941), .Z(N13269) );
  NANDN U9130 ( .A(n6942), .B(n6943), .Z(n6941) );
  OR U9131 ( .A(n6944), .B(n6945), .Z(n6943) );
  NAND U9132 ( .A(n6944), .B(n6945), .Z(n6940) );
  XOR U9133 ( .A(n6944), .B(n6946), .Z(N13268) );
  XNOR U9134 ( .A(n6942), .B(n6945), .Z(n6946) );
  AND U9135 ( .A(n6947), .B(n6948), .Z(n6945) );
  NANDN U9136 ( .A(n6949), .B(n6950), .Z(n6948) );
  NANDN U9137 ( .A(n6951), .B(n6952), .Z(n6950) );
  NANDN U9138 ( .A(n6952), .B(n6951), .Z(n6947) );
  NAND U9139 ( .A(n6953), .B(n6954), .Z(n6942) );
  NANDN U9140 ( .A(n6955), .B(n6956), .Z(n6954) );
  OR U9141 ( .A(n6957), .B(n6958), .Z(n6956) );
  NAND U9142 ( .A(n6958), .B(n6957), .Z(n6953) );
  AND U9143 ( .A(n6959), .B(n6960), .Z(n6944) );
  NANDN U9144 ( .A(n6961), .B(n6962), .Z(n6960) );
  NANDN U9145 ( .A(n6963), .B(n6964), .Z(n6962) );
  NANDN U9146 ( .A(n6964), .B(n6963), .Z(n6959) );
  XOR U9147 ( .A(n6958), .B(n6965), .Z(N13267) );
  XOR U9148 ( .A(n6955), .B(n6957), .Z(n6965) );
  XNOR U9149 ( .A(n6951), .B(n6966), .Z(n6957) );
  XNOR U9150 ( .A(n6949), .B(n6952), .Z(n6966) );
  NAND U9151 ( .A(n6967), .B(n6968), .Z(n6952) );
  NAND U9152 ( .A(n6969), .B(n6970), .Z(n6968) );
  OR U9153 ( .A(n6971), .B(n6972), .Z(n6969) );
  NANDN U9154 ( .A(n6973), .B(n6971), .Z(n6967) );
  IV U9155 ( .A(n6972), .Z(n6973) );
  NAND U9156 ( .A(n6974), .B(n6975), .Z(n6949) );
  NAND U9157 ( .A(n6976), .B(n6977), .Z(n6975) );
  NANDN U9158 ( .A(n6978), .B(n6979), .Z(n6976) );
  NANDN U9159 ( .A(n6979), .B(n6978), .Z(n6974) );
  AND U9160 ( .A(n6980), .B(n6981), .Z(n6951) );
  NAND U9161 ( .A(n6982), .B(n6983), .Z(n6981) );
  OR U9162 ( .A(n6984), .B(n6985), .Z(n6982) );
  NANDN U9163 ( .A(n6986), .B(n6984), .Z(n6980) );
  NAND U9164 ( .A(n6987), .B(n6988), .Z(n6955) );
  NANDN U9165 ( .A(n6989), .B(n6990), .Z(n6988) );
  OR U9166 ( .A(n6991), .B(n6992), .Z(n6990) );
  NANDN U9167 ( .A(n6993), .B(n6991), .Z(n6987) );
  IV U9168 ( .A(n6992), .Z(n6993) );
  XNOR U9169 ( .A(n6963), .B(n6994), .Z(n6958) );
  XNOR U9170 ( .A(n6961), .B(n6964), .Z(n6994) );
  NAND U9171 ( .A(n6995), .B(n6996), .Z(n6964) );
  NAND U9172 ( .A(n6997), .B(n6998), .Z(n6996) );
  OR U9173 ( .A(n6999), .B(n7000), .Z(n6997) );
  NANDN U9174 ( .A(n7001), .B(n6999), .Z(n6995) );
  IV U9175 ( .A(n7000), .Z(n7001) );
  NAND U9176 ( .A(n7002), .B(n7003), .Z(n6961) );
  NAND U9177 ( .A(n7004), .B(n7005), .Z(n7003) );
  NANDN U9178 ( .A(n7006), .B(n7007), .Z(n7004) );
  NANDN U9179 ( .A(n7007), .B(n7006), .Z(n7002) );
  AND U9180 ( .A(n7008), .B(n7009), .Z(n6963) );
  NAND U9181 ( .A(n7010), .B(n7011), .Z(n7009) );
  OR U9182 ( .A(n7012), .B(n7013), .Z(n7010) );
  NANDN U9183 ( .A(n7014), .B(n7012), .Z(n7008) );
  XNOR U9184 ( .A(n6989), .B(n7015), .Z(N13266) );
  XOR U9185 ( .A(n6991), .B(n6992), .Z(n7015) );
  XNOR U9186 ( .A(n7005), .B(n7016), .Z(n6992) );
  XOR U9187 ( .A(n7006), .B(n7007), .Z(n7016) );
  XOR U9188 ( .A(n7012), .B(n7017), .Z(n7007) );
  XOR U9189 ( .A(n7011), .B(n7014), .Z(n7017) );
  IV U9190 ( .A(n7013), .Z(n7014) );
  NAND U9191 ( .A(n7018), .B(n7019), .Z(n7013) );
  OR U9192 ( .A(n7020), .B(n7021), .Z(n7019) );
  OR U9193 ( .A(n7022), .B(n7023), .Z(n7018) );
  NAND U9194 ( .A(n7024), .B(n7025), .Z(n7011) );
  OR U9195 ( .A(n7026), .B(n7027), .Z(n7025) );
  OR U9196 ( .A(n7028), .B(n7029), .Z(n7024) );
  NOR U9197 ( .A(n7030), .B(n7031), .Z(n7012) );
  ANDN U9198 ( .B(n7032), .A(n7033), .Z(n7006) );
  XNOR U9199 ( .A(n6999), .B(n7034), .Z(n7005) );
  XNOR U9200 ( .A(n6998), .B(n7000), .Z(n7034) );
  NAND U9201 ( .A(n7035), .B(n7036), .Z(n7000) );
  OR U9202 ( .A(n7037), .B(n7038), .Z(n7036) );
  OR U9203 ( .A(n7039), .B(n7040), .Z(n7035) );
  NAND U9204 ( .A(n7041), .B(n7042), .Z(n6998) );
  OR U9205 ( .A(n7043), .B(n7044), .Z(n7042) );
  OR U9206 ( .A(n7045), .B(n7046), .Z(n7041) );
  ANDN U9207 ( .B(n7047), .A(n7048), .Z(n6999) );
  IV U9208 ( .A(n7049), .Z(n7047) );
  ANDN U9209 ( .B(n7050), .A(n7051), .Z(n6991) );
  XOR U9210 ( .A(n6977), .B(n7052), .Z(n6989) );
  XOR U9211 ( .A(n6978), .B(n6979), .Z(n7052) );
  XOR U9212 ( .A(n6984), .B(n7053), .Z(n6979) );
  XOR U9213 ( .A(n6983), .B(n6986), .Z(n7053) );
  IV U9214 ( .A(n6985), .Z(n6986) );
  NAND U9215 ( .A(n7054), .B(n7055), .Z(n6985) );
  OR U9216 ( .A(n7056), .B(n7057), .Z(n7055) );
  OR U9217 ( .A(n7058), .B(n7059), .Z(n7054) );
  NAND U9218 ( .A(n7060), .B(n7061), .Z(n6983) );
  OR U9219 ( .A(n7062), .B(n7063), .Z(n7061) );
  OR U9220 ( .A(n7064), .B(n7065), .Z(n7060) );
  NOR U9221 ( .A(n7066), .B(n7067), .Z(n6984) );
  ANDN U9222 ( .B(n7068), .A(n7069), .Z(n6978) );
  IV U9223 ( .A(n7070), .Z(n7068) );
  XNOR U9224 ( .A(n6971), .B(n7071), .Z(n6977) );
  XNOR U9225 ( .A(n6970), .B(n6972), .Z(n7071) );
  NAND U9226 ( .A(n7072), .B(n7073), .Z(n6972) );
  OR U9227 ( .A(n7074), .B(n7075), .Z(n7073) );
  OR U9228 ( .A(n7076), .B(n7077), .Z(n7072) );
  NAND U9229 ( .A(n7078), .B(n7079), .Z(n6970) );
  OR U9230 ( .A(n7080), .B(n7081), .Z(n7079) );
  OR U9231 ( .A(n7082), .B(n7083), .Z(n7078) );
  ANDN U9232 ( .B(n7084), .A(n7085), .Z(n6971) );
  IV U9233 ( .A(n7086), .Z(n7084) );
  XNOR U9234 ( .A(n7051), .B(n7050), .Z(N13265) );
  XOR U9235 ( .A(n7070), .B(n7069), .Z(n7050) );
  XNOR U9236 ( .A(n7085), .B(n7086), .Z(n7069) );
  XNOR U9237 ( .A(n7080), .B(n7081), .Z(n7086) );
  XNOR U9238 ( .A(n7082), .B(n7083), .Z(n7081) );
  XNOR U9239 ( .A(y[1069]), .B(x[1069]), .Z(n7083) );
  XNOR U9240 ( .A(y[1070]), .B(x[1070]), .Z(n7082) );
  XNOR U9241 ( .A(y[1068]), .B(x[1068]), .Z(n7080) );
  XNOR U9242 ( .A(n7074), .B(n7075), .Z(n7085) );
  XNOR U9243 ( .A(y[1065]), .B(x[1065]), .Z(n7075) );
  XNOR U9244 ( .A(n7076), .B(n7077), .Z(n7074) );
  XNOR U9245 ( .A(y[1066]), .B(x[1066]), .Z(n7077) );
  XNOR U9246 ( .A(y[1067]), .B(x[1067]), .Z(n7076) );
  XNOR U9247 ( .A(n7067), .B(n7066), .Z(n7070) );
  XNOR U9248 ( .A(n7062), .B(n7063), .Z(n7066) );
  XNOR U9249 ( .A(y[1062]), .B(x[1062]), .Z(n7063) );
  XNOR U9250 ( .A(n7064), .B(n7065), .Z(n7062) );
  XNOR U9251 ( .A(y[1063]), .B(x[1063]), .Z(n7065) );
  XNOR U9252 ( .A(y[1064]), .B(x[1064]), .Z(n7064) );
  XNOR U9253 ( .A(n7056), .B(n7057), .Z(n7067) );
  XNOR U9254 ( .A(y[1059]), .B(x[1059]), .Z(n7057) );
  XNOR U9255 ( .A(n7058), .B(n7059), .Z(n7056) );
  XNOR U9256 ( .A(y[1060]), .B(x[1060]), .Z(n7059) );
  XNOR U9257 ( .A(y[1061]), .B(x[1061]), .Z(n7058) );
  XOR U9258 ( .A(n7032), .B(n7033), .Z(n7051) );
  XNOR U9259 ( .A(n7048), .B(n7049), .Z(n7033) );
  XNOR U9260 ( .A(n7043), .B(n7044), .Z(n7049) );
  XNOR U9261 ( .A(n7045), .B(n7046), .Z(n7044) );
  XNOR U9262 ( .A(y[1057]), .B(x[1057]), .Z(n7046) );
  XNOR U9263 ( .A(y[1058]), .B(x[1058]), .Z(n7045) );
  XNOR U9264 ( .A(y[1056]), .B(x[1056]), .Z(n7043) );
  XNOR U9265 ( .A(n7037), .B(n7038), .Z(n7048) );
  XNOR U9266 ( .A(y[1053]), .B(x[1053]), .Z(n7038) );
  XNOR U9267 ( .A(n7039), .B(n7040), .Z(n7037) );
  XNOR U9268 ( .A(y[1054]), .B(x[1054]), .Z(n7040) );
  XNOR U9269 ( .A(y[1055]), .B(x[1055]), .Z(n7039) );
  XOR U9270 ( .A(n7031), .B(n7030), .Z(n7032) );
  XNOR U9271 ( .A(n7026), .B(n7027), .Z(n7030) );
  XNOR U9272 ( .A(y[1050]), .B(x[1050]), .Z(n7027) );
  XNOR U9273 ( .A(n7028), .B(n7029), .Z(n7026) );
  XNOR U9274 ( .A(y[1051]), .B(x[1051]), .Z(n7029) );
  XNOR U9275 ( .A(y[1052]), .B(x[1052]), .Z(n7028) );
  XNOR U9276 ( .A(n7020), .B(n7021), .Z(n7031) );
  XNOR U9277 ( .A(y[1047]), .B(x[1047]), .Z(n7021) );
  XNOR U9278 ( .A(n7022), .B(n7023), .Z(n7020) );
  XNOR U9279 ( .A(y[1048]), .B(x[1048]), .Z(n7023) );
  XNOR U9280 ( .A(y[1049]), .B(x[1049]), .Z(n7022) );
  NAND U9281 ( .A(n7087), .B(n7088), .Z(N13258) );
  NANDN U9282 ( .A(n7089), .B(n7090), .Z(n7088) );
  OR U9283 ( .A(n7091), .B(n7092), .Z(n7090) );
  NAND U9284 ( .A(n7091), .B(n7092), .Z(n7087) );
  XOR U9285 ( .A(n7091), .B(n7093), .Z(N13257) );
  XNOR U9286 ( .A(n7089), .B(n7092), .Z(n7093) );
  AND U9287 ( .A(n7094), .B(n7095), .Z(n7092) );
  NANDN U9288 ( .A(n7096), .B(n7097), .Z(n7095) );
  NANDN U9289 ( .A(n7098), .B(n7099), .Z(n7097) );
  NANDN U9290 ( .A(n7099), .B(n7098), .Z(n7094) );
  NAND U9291 ( .A(n7100), .B(n7101), .Z(n7089) );
  NANDN U9292 ( .A(n7102), .B(n7103), .Z(n7101) );
  OR U9293 ( .A(n7104), .B(n7105), .Z(n7103) );
  NAND U9294 ( .A(n7105), .B(n7104), .Z(n7100) );
  AND U9295 ( .A(n7106), .B(n7107), .Z(n7091) );
  NANDN U9296 ( .A(n7108), .B(n7109), .Z(n7107) );
  NANDN U9297 ( .A(n7110), .B(n7111), .Z(n7109) );
  NANDN U9298 ( .A(n7111), .B(n7110), .Z(n7106) );
  XOR U9299 ( .A(n7105), .B(n7112), .Z(N13256) );
  XOR U9300 ( .A(n7102), .B(n7104), .Z(n7112) );
  XNOR U9301 ( .A(n7098), .B(n7113), .Z(n7104) );
  XNOR U9302 ( .A(n7096), .B(n7099), .Z(n7113) );
  NAND U9303 ( .A(n7114), .B(n7115), .Z(n7099) );
  NAND U9304 ( .A(n7116), .B(n7117), .Z(n7115) );
  OR U9305 ( .A(n7118), .B(n7119), .Z(n7116) );
  NANDN U9306 ( .A(n7120), .B(n7118), .Z(n7114) );
  IV U9307 ( .A(n7119), .Z(n7120) );
  NAND U9308 ( .A(n7121), .B(n7122), .Z(n7096) );
  NAND U9309 ( .A(n7123), .B(n7124), .Z(n7122) );
  NANDN U9310 ( .A(n7125), .B(n7126), .Z(n7123) );
  NANDN U9311 ( .A(n7126), .B(n7125), .Z(n7121) );
  AND U9312 ( .A(n7127), .B(n7128), .Z(n7098) );
  NAND U9313 ( .A(n7129), .B(n7130), .Z(n7128) );
  OR U9314 ( .A(n7131), .B(n7132), .Z(n7129) );
  NANDN U9315 ( .A(n7133), .B(n7131), .Z(n7127) );
  NAND U9316 ( .A(n7134), .B(n7135), .Z(n7102) );
  NANDN U9317 ( .A(n7136), .B(n7137), .Z(n7135) );
  OR U9318 ( .A(n7138), .B(n7139), .Z(n7137) );
  NANDN U9319 ( .A(n7140), .B(n7138), .Z(n7134) );
  IV U9320 ( .A(n7139), .Z(n7140) );
  XNOR U9321 ( .A(n7110), .B(n7141), .Z(n7105) );
  XNOR U9322 ( .A(n7108), .B(n7111), .Z(n7141) );
  NAND U9323 ( .A(n7142), .B(n7143), .Z(n7111) );
  NAND U9324 ( .A(n7144), .B(n7145), .Z(n7143) );
  OR U9325 ( .A(n7146), .B(n7147), .Z(n7144) );
  NANDN U9326 ( .A(n7148), .B(n7146), .Z(n7142) );
  IV U9327 ( .A(n7147), .Z(n7148) );
  NAND U9328 ( .A(n7149), .B(n7150), .Z(n7108) );
  NAND U9329 ( .A(n7151), .B(n7152), .Z(n7150) );
  NANDN U9330 ( .A(n7153), .B(n7154), .Z(n7151) );
  NANDN U9331 ( .A(n7154), .B(n7153), .Z(n7149) );
  AND U9332 ( .A(n7155), .B(n7156), .Z(n7110) );
  NAND U9333 ( .A(n7157), .B(n7158), .Z(n7156) );
  OR U9334 ( .A(n7159), .B(n7160), .Z(n7157) );
  NANDN U9335 ( .A(n7161), .B(n7159), .Z(n7155) );
  XNOR U9336 ( .A(n7136), .B(n7162), .Z(N13255) );
  XOR U9337 ( .A(n7138), .B(n7139), .Z(n7162) );
  XNOR U9338 ( .A(n7152), .B(n7163), .Z(n7139) );
  XOR U9339 ( .A(n7153), .B(n7154), .Z(n7163) );
  XOR U9340 ( .A(n7159), .B(n7164), .Z(n7154) );
  XOR U9341 ( .A(n7158), .B(n7161), .Z(n7164) );
  IV U9342 ( .A(n7160), .Z(n7161) );
  NAND U9343 ( .A(n7165), .B(n7166), .Z(n7160) );
  OR U9344 ( .A(n7167), .B(n7168), .Z(n7166) );
  OR U9345 ( .A(n7169), .B(n7170), .Z(n7165) );
  NAND U9346 ( .A(n7171), .B(n7172), .Z(n7158) );
  OR U9347 ( .A(n7173), .B(n7174), .Z(n7172) );
  OR U9348 ( .A(n7175), .B(n7176), .Z(n7171) );
  NOR U9349 ( .A(n7177), .B(n7178), .Z(n7159) );
  ANDN U9350 ( .B(n7179), .A(n7180), .Z(n7153) );
  XNOR U9351 ( .A(n7146), .B(n7181), .Z(n7152) );
  XNOR U9352 ( .A(n7145), .B(n7147), .Z(n7181) );
  NAND U9353 ( .A(n7182), .B(n7183), .Z(n7147) );
  OR U9354 ( .A(n7184), .B(n7185), .Z(n7183) );
  OR U9355 ( .A(n7186), .B(n7187), .Z(n7182) );
  NAND U9356 ( .A(n7188), .B(n7189), .Z(n7145) );
  OR U9357 ( .A(n7190), .B(n7191), .Z(n7189) );
  OR U9358 ( .A(n7192), .B(n7193), .Z(n7188) );
  ANDN U9359 ( .B(n7194), .A(n7195), .Z(n7146) );
  IV U9360 ( .A(n7196), .Z(n7194) );
  ANDN U9361 ( .B(n7197), .A(n7198), .Z(n7138) );
  XOR U9362 ( .A(n7124), .B(n7199), .Z(n7136) );
  XOR U9363 ( .A(n7125), .B(n7126), .Z(n7199) );
  XOR U9364 ( .A(n7131), .B(n7200), .Z(n7126) );
  XOR U9365 ( .A(n7130), .B(n7133), .Z(n7200) );
  IV U9366 ( .A(n7132), .Z(n7133) );
  NAND U9367 ( .A(n7201), .B(n7202), .Z(n7132) );
  OR U9368 ( .A(n7203), .B(n7204), .Z(n7202) );
  OR U9369 ( .A(n7205), .B(n7206), .Z(n7201) );
  NAND U9370 ( .A(n7207), .B(n7208), .Z(n7130) );
  OR U9371 ( .A(n7209), .B(n7210), .Z(n7208) );
  OR U9372 ( .A(n7211), .B(n7212), .Z(n7207) );
  NOR U9373 ( .A(n7213), .B(n7214), .Z(n7131) );
  ANDN U9374 ( .B(n7215), .A(n7216), .Z(n7125) );
  IV U9375 ( .A(n7217), .Z(n7215) );
  XNOR U9376 ( .A(n7118), .B(n7218), .Z(n7124) );
  XNOR U9377 ( .A(n7117), .B(n7119), .Z(n7218) );
  NAND U9378 ( .A(n7219), .B(n7220), .Z(n7119) );
  OR U9379 ( .A(n7221), .B(n7222), .Z(n7220) );
  OR U9380 ( .A(n7223), .B(n7224), .Z(n7219) );
  NAND U9381 ( .A(n7225), .B(n7226), .Z(n7117) );
  OR U9382 ( .A(n7227), .B(n7228), .Z(n7226) );
  OR U9383 ( .A(n7229), .B(n7230), .Z(n7225) );
  ANDN U9384 ( .B(n7231), .A(n7232), .Z(n7118) );
  IV U9385 ( .A(n7233), .Z(n7231) );
  XNOR U9386 ( .A(n7198), .B(n7197), .Z(N13254) );
  XOR U9387 ( .A(n7217), .B(n7216), .Z(n7197) );
  XNOR U9388 ( .A(n7232), .B(n7233), .Z(n7216) );
  XNOR U9389 ( .A(n7227), .B(n7228), .Z(n7233) );
  XNOR U9390 ( .A(n7229), .B(n7230), .Z(n7228) );
  XNOR U9391 ( .A(y[1045]), .B(x[1045]), .Z(n7230) );
  XNOR U9392 ( .A(y[1046]), .B(x[1046]), .Z(n7229) );
  XNOR U9393 ( .A(y[1044]), .B(x[1044]), .Z(n7227) );
  XNOR U9394 ( .A(n7221), .B(n7222), .Z(n7232) );
  XNOR U9395 ( .A(y[1041]), .B(x[1041]), .Z(n7222) );
  XNOR U9396 ( .A(n7223), .B(n7224), .Z(n7221) );
  XNOR U9397 ( .A(y[1042]), .B(x[1042]), .Z(n7224) );
  XNOR U9398 ( .A(y[1043]), .B(x[1043]), .Z(n7223) );
  XNOR U9399 ( .A(n7214), .B(n7213), .Z(n7217) );
  XNOR U9400 ( .A(n7209), .B(n7210), .Z(n7213) );
  XNOR U9401 ( .A(y[1038]), .B(x[1038]), .Z(n7210) );
  XNOR U9402 ( .A(n7211), .B(n7212), .Z(n7209) );
  XNOR U9403 ( .A(y[1039]), .B(x[1039]), .Z(n7212) );
  XNOR U9404 ( .A(y[1040]), .B(x[1040]), .Z(n7211) );
  XNOR U9405 ( .A(n7203), .B(n7204), .Z(n7214) );
  XNOR U9406 ( .A(y[1035]), .B(x[1035]), .Z(n7204) );
  XNOR U9407 ( .A(n7205), .B(n7206), .Z(n7203) );
  XNOR U9408 ( .A(y[1036]), .B(x[1036]), .Z(n7206) );
  XNOR U9409 ( .A(y[1037]), .B(x[1037]), .Z(n7205) );
  XOR U9410 ( .A(n7179), .B(n7180), .Z(n7198) );
  XNOR U9411 ( .A(n7195), .B(n7196), .Z(n7180) );
  XNOR U9412 ( .A(n7190), .B(n7191), .Z(n7196) );
  XNOR U9413 ( .A(n7192), .B(n7193), .Z(n7191) );
  XNOR U9414 ( .A(y[1033]), .B(x[1033]), .Z(n7193) );
  XNOR U9415 ( .A(y[1034]), .B(x[1034]), .Z(n7192) );
  XNOR U9416 ( .A(y[1032]), .B(x[1032]), .Z(n7190) );
  XNOR U9417 ( .A(n7184), .B(n7185), .Z(n7195) );
  XNOR U9418 ( .A(y[1029]), .B(x[1029]), .Z(n7185) );
  XNOR U9419 ( .A(n7186), .B(n7187), .Z(n7184) );
  XNOR U9420 ( .A(y[1030]), .B(x[1030]), .Z(n7187) );
  XNOR U9421 ( .A(y[1031]), .B(x[1031]), .Z(n7186) );
  XOR U9422 ( .A(n7178), .B(n7177), .Z(n7179) );
  XNOR U9423 ( .A(n7173), .B(n7174), .Z(n7177) );
  XNOR U9424 ( .A(y[1026]), .B(x[1026]), .Z(n7174) );
  XNOR U9425 ( .A(n7175), .B(n7176), .Z(n7173) );
  XNOR U9426 ( .A(y[1027]), .B(x[1027]), .Z(n7176) );
  XNOR U9427 ( .A(y[1028]), .B(x[1028]), .Z(n7175) );
  XNOR U9428 ( .A(n7167), .B(n7168), .Z(n7178) );
  XNOR U9429 ( .A(y[1023]), .B(x[1023]), .Z(n7168) );
  XNOR U9430 ( .A(n7169), .B(n7170), .Z(n7167) );
  XNOR U9431 ( .A(y[1024]), .B(x[1024]), .Z(n7170) );
  XNOR U9432 ( .A(y[1025]), .B(x[1025]), .Z(n7169) );
  NAND U9433 ( .A(n7234), .B(n7235), .Z(N13247) );
  NANDN U9434 ( .A(n7236), .B(n7237), .Z(n7235) );
  OR U9435 ( .A(n7238), .B(n7239), .Z(n7237) );
  NAND U9436 ( .A(n7238), .B(n7239), .Z(n7234) );
  XOR U9437 ( .A(n7238), .B(n7240), .Z(N13246) );
  XNOR U9438 ( .A(n7236), .B(n7239), .Z(n7240) );
  AND U9439 ( .A(n7241), .B(n7242), .Z(n7239) );
  NANDN U9440 ( .A(n7243), .B(n7244), .Z(n7242) );
  NANDN U9441 ( .A(n7245), .B(n7246), .Z(n7244) );
  NANDN U9442 ( .A(n7246), .B(n7245), .Z(n7241) );
  NAND U9443 ( .A(n7247), .B(n7248), .Z(n7236) );
  NANDN U9444 ( .A(n7249), .B(n7250), .Z(n7248) );
  OR U9445 ( .A(n7251), .B(n7252), .Z(n7250) );
  NAND U9446 ( .A(n7252), .B(n7251), .Z(n7247) );
  AND U9447 ( .A(n7253), .B(n7254), .Z(n7238) );
  NANDN U9448 ( .A(n7255), .B(n7256), .Z(n7254) );
  NANDN U9449 ( .A(n7257), .B(n7258), .Z(n7256) );
  NANDN U9450 ( .A(n7258), .B(n7257), .Z(n7253) );
  XOR U9451 ( .A(n7252), .B(n7259), .Z(N13245) );
  XOR U9452 ( .A(n7249), .B(n7251), .Z(n7259) );
  XNOR U9453 ( .A(n7245), .B(n7260), .Z(n7251) );
  XNOR U9454 ( .A(n7243), .B(n7246), .Z(n7260) );
  NAND U9455 ( .A(n7261), .B(n7262), .Z(n7246) );
  NAND U9456 ( .A(n7263), .B(n7264), .Z(n7262) );
  OR U9457 ( .A(n7265), .B(n7266), .Z(n7263) );
  NANDN U9458 ( .A(n7267), .B(n7265), .Z(n7261) );
  IV U9459 ( .A(n7266), .Z(n7267) );
  NAND U9460 ( .A(n7268), .B(n7269), .Z(n7243) );
  NAND U9461 ( .A(n7270), .B(n7271), .Z(n7269) );
  NANDN U9462 ( .A(n7272), .B(n7273), .Z(n7270) );
  NANDN U9463 ( .A(n7273), .B(n7272), .Z(n7268) );
  AND U9464 ( .A(n7274), .B(n7275), .Z(n7245) );
  NAND U9465 ( .A(n7276), .B(n7277), .Z(n7275) );
  OR U9466 ( .A(n7278), .B(n7279), .Z(n7276) );
  NANDN U9467 ( .A(n7280), .B(n7278), .Z(n7274) );
  NAND U9468 ( .A(n7281), .B(n7282), .Z(n7249) );
  NANDN U9469 ( .A(n7283), .B(n7284), .Z(n7282) );
  OR U9470 ( .A(n7285), .B(n7286), .Z(n7284) );
  NANDN U9471 ( .A(n7287), .B(n7285), .Z(n7281) );
  IV U9472 ( .A(n7286), .Z(n7287) );
  XNOR U9473 ( .A(n7257), .B(n7288), .Z(n7252) );
  XNOR U9474 ( .A(n7255), .B(n7258), .Z(n7288) );
  NAND U9475 ( .A(n7289), .B(n7290), .Z(n7258) );
  NAND U9476 ( .A(n7291), .B(n7292), .Z(n7290) );
  OR U9477 ( .A(n7293), .B(n7294), .Z(n7291) );
  NANDN U9478 ( .A(n7295), .B(n7293), .Z(n7289) );
  IV U9479 ( .A(n7294), .Z(n7295) );
  NAND U9480 ( .A(n7296), .B(n7297), .Z(n7255) );
  NAND U9481 ( .A(n7298), .B(n7299), .Z(n7297) );
  NANDN U9482 ( .A(n7300), .B(n7301), .Z(n7298) );
  NANDN U9483 ( .A(n7301), .B(n7300), .Z(n7296) );
  AND U9484 ( .A(n7302), .B(n7303), .Z(n7257) );
  NAND U9485 ( .A(n7304), .B(n7305), .Z(n7303) );
  OR U9486 ( .A(n7306), .B(n7307), .Z(n7304) );
  NANDN U9487 ( .A(n7308), .B(n7306), .Z(n7302) );
  XNOR U9488 ( .A(n7283), .B(n7309), .Z(N13244) );
  XOR U9489 ( .A(n7285), .B(n7286), .Z(n7309) );
  XNOR U9490 ( .A(n7299), .B(n7310), .Z(n7286) );
  XOR U9491 ( .A(n7300), .B(n7301), .Z(n7310) );
  XOR U9492 ( .A(n7306), .B(n7311), .Z(n7301) );
  XOR U9493 ( .A(n7305), .B(n7308), .Z(n7311) );
  IV U9494 ( .A(n7307), .Z(n7308) );
  NAND U9495 ( .A(n7312), .B(n7313), .Z(n7307) );
  OR U9496 ( .A(n7314), .B(n7315), .Z(n7313) );
  OR U9497 ( .A(n7316), .B(n7317), .Z(n7312) );
  NAND U9498 ( .A(n7318), .B(n7319), .Z(n7305) );
  OR U9499 ( .A(n7320), .B(n7321), .Z(n7319) );
  OR U9500 ( .A(n7322), .B(n7323), .Z(n7318) );
  NOR U9501 ( .A(n7324), .B(n7325), .Z(n7306) );
  ANDN U9502 ( .B(n7326), .A(n7327), .Z(n7300) );
  XNOR U9503 ( .A(n7293), .B(n7328), .Z(n7299) );
  XNOR U9504 ( .A(n7292), .B(n7294), .Z(n7328) );
  NAND U9505 ( .A(n7329), .B(n7330), .Z(n7294) );
  OR U9506 ( .A(n7331), .B(n7332), .Z(n7330) );
  OR U9507 ( .A(n7333), .B(n7334), .Z(n7329) );
  NAND U9508 ( .A(n7335), .B(n7336), .Z(n7292) );
  OR U9509 ( .A(n7337), .B(n7338), .Z(n7336) );
  OR U9510 ( .A(n7339), .B(n7340), .Z(n7335) );
  ANDN U9511 ( .B(n7341), .A(n7342), .Z(n7293) );
  IV U9512 ( .A(n7343), .Z(n7341) );
  ANDN U9513 ( .B(n7344), .A(n7345), .Z(n7285) );
  XOR U9514 ( .A(n7271), .B(n7346), .Z(n7283) );
  XOR U9515 ( .A(n7272), .B(n7273), .Z(n7346) );
  XOR U9516 ( .A(n7278), .B(n7347), .Z(n7273) );
  XOR U9517 ( .A(n7277), .B(n7280), .Z(n7347) );
  IV U9518 ( .A(n7279), .Z(n7280) );
  NAND U9519 ( .A(n7348), .B(n7349), .Z(n7279) );
  OR U9520 ( .A(n7350), .B(n7351), .Z(n7349) );
  OR U9521 ( .A(n7352), .B(n7353), .Z(n7348) );
  NAND U9522 ( .A(n7354), .B(n7355), .Z(n7277) );
  OR U9523 ( .A(n7356), .B(n7357), .Z(n7355) );
  OR U9524 ( .A(n7358), .B(n7359), .Z(n7354) );
  NOR U9525 ( .A(n7360), .B(n7361), .Z(n7278) );
  ANDN U9526 ( .B(n7362), .A(n7363), .Z(n7272) );
  IV U9527 ( .A(n7364), .Z(n7362) );
  XNOR U9528 ( .A(n7265), .B(n7365), .Z(n7271) );
  XNOR U9529 ( .A(n7264), .B(n7266), .Z(n7365) );
  NAND U9530 ( .A(n7366), .B(n7367), .Z(n7266) );
  OR U9531 ( .A(n7368), .B(n7369), .Z(n7367) );
  OR U9532 ( .A(n7370), .B(n7371), .Z(n7366) );
  NAND U9533 ( .A(n7372), .B(n7373), .Z(n7264) );
  OR U9534 ( .A(n7374), .B(n7375), .Z(n7373) );
  OR U9535 ( .A(n7376), .B(n7377), .Z(n7372) );
  ANDN U9536 ( .B(n7378), .A(n7379), .Z(n7265) );
  IV U9537 ( .A(n7380), .Z(n7378) );
  XNOR U9538 ( .A(n7345), .B(n7344), .Z(N13243) );
  XOR U9539 ( .A(n7364), .B(n7363), .Z(n7344) );
  XNOR U9540 ( .A(n7379), .B(n7380), .Z(n7363) );
  XNOR U9541 ( .A(n7374), .B(n7375), .Z(n7380) );
  XNOR U9542 ( .A(n7376), .B(n7377), .Z(n7375) );
  XNOR U9543 ( .A(y[1021]), .B(x[1021]), .Z(n7377) );
  XNOR U9544 ( .A(y[1022]), .B(x[1022]), .Z(n7376) );
  XNOR U9545 ( .A(y[1020]), .B(x[1020]), .Z(n7374) );
  XNOR U9546 ( .A(n7368), .B(n7369), .Z(n7379) );
  XNOR U9547 ( .A(y[1017]), .B(x[1017]), .Z(n7369) );
  XNOR U9548 ( .A(n7370), .B(n7371), .Z(n7368) );
  XNOR U9549 ( .A(y[1018]), .B(x[1018]), .Z(n7371) );
  XNOR U9550 ( .A(y[1019]), .B(x[1019]), .Z(n7370) );
  XNOR U9551 ( .A(n7361), .B(n7360), .Z(n7364) );
  XNOR U9552 ( .A(n7356), .B(n7357), .Z(n7360) );
  XNOR U9553 ( .A(y[1014]), .B(x[1014]), .Z(n7357) );
  XNOR U9554 ( .A(n7358), .B(n7359), .Z(n7356) );
  XNOR U9555 ( .A(y[1015]), .B(x[1015]), .Z(n7359) );
  XNOR U9556 ( .A(y[1016]), .B(x[1016]), .Z(n7358) );
  XNOR U9557 ( .A(n7350), .B(n7351), .Z(n7361) );
  XNOR U9558 ( .A(y[1011]), .B(x[1011]), .Z(n7351) );
  XNOR U9559 ( .A(n7352), .B(n7353), .Z(n7350) );
  XNOR U9560 ( .A(y[1012]), .B(x[1012]), .Z(n7353) );
  XNOR U9561 ( .A(y[1013]), .B(x[1013]), .Z(n7352) );
  XOR U9562 ( .A(n7326), .B(n7327), .Z(n7345) );
  XNOR U9563 ( .A(n7342), .B(n7343), .Z(n7327) );
  XNOR U9564 ( .A(n7337), .B(n7338), .Z(n7343) );
  XNOR U9565 ( .A(n7339), .B(n7340), .Z(n7338) );
  XNOR U9566 ( .A(y[1009]), .B(x[1009]), .Z(n7340) );
  XNOR U9567 ( .A(y[1010]), .B(x[1010]), .Z(n7339) );
  XNOR U9568 ( .A(y[1008]), .B(x[1008]), .Z(n7337) );
  XNOR U9569 ( .A(n7331), .B(n7332), .Z(n7342) );
  XNOR U9570 ( .A(y[1005]), .B(x[1005]), .Z(n7332) );
  XNOR U9571 ( .A(n7333), .B(n7334), .Z(n7331) );
  XNOR U9572 ( .A(y[1006]), .B(x[1006]), .Z(n7334) );
  XNOR U9573 ( .A(y[1007]), .B(x[1007]), .Z(n7333) );
  XOR U9574 ( .A(n7325), .B(n7324), .Z(n7326) );
  XNOR U9575 ( .A(n7320), .B(n7321), .Z(n7324) );
  XNOR U9576 ( .A(y[1002]), .B(x[1002]), .Z(n7321) );
  XNOR U9577 ( .A(n7322), .B(n7323), .Z(n7320) );
  XNOR U9578 ( .A(y[1003]), .B(x[1003]), .Z(n7323) );
  XNOR U9579 ( .A(y[1004]), .B(x[1004]), .Z(n7322) );
  XNOR U9580 ( .A(n7314), .B(n7315), .Z(n7325) );
  XNOR U9581 ( .A(y[999]), .B(x[999]), .Z(n7315) );
  XNOR U9582 ( .A(n7316), .B(n7317), .Z(n7314) );
  XNOR U9583 ( .A(y[1000]), .B(x[1000]), .Z(n7317) );
  XNOR U9584 ( .A(y[1001]), .B(x[1001]), .Z(n7316) );
  NAND U9585 ( .A(n7381), .B(n7382), .Z(N13236) );
  NANDN U9586 ( .A(n7383), .B(n7384), .Z(n7382) );
  OR U9587 ( .A(n7385), .B(n7386), .Z(n7384) );
  NAND U9588 ( .A(n7385), .B(n7386), .Z(n7381) );
  XOR U9589 ( .A(n7385), .B(n7387), .Z(N13235) );
  XNOR U9590 ( .A(n7383), .B(n7386), .Z(n7387) );
  AND U9591 ( .A(n7388), .B(n7389), .Z(n7386) );
  NANDN U9592 ( .A(n7390), .B(n7391), .Z(n7389) );
  NANDN U9593 ( .A(n7392), .B(n7393), .Z(n7391) );
  NANDN U9594 ( .A(n7393), .B(n7392), .Z(n7388) );
  NAND U9595 ( .A(n7394), .B(n7395), .Z(n7383) );
  NANDN U9596 ( .A(n7396), .B(n7397), .Z(n7395) );
  OR U9597 ( .A(n7398), .B(n7399), .Z(n7397) );
  NAND U9598 ( .A(n7399), .B(n7398), .Z(n7394) );
  AND U9599 ( .A(n7400), .B(n7401), .Z(n7385) );
  NANDN U9600 ( .A(n7402), .B(n7403), .Z(n7401) );
  NANDN U9601 ( .A(n7404), .B(n7405), .Z(n7403) );
  NANDN U9602 ( .A(n7405), .B(n7404), .Z(n7400) );
  XOR U9603 ( .A(n7399), .B(n7406), .Z(N13234) );
  XOR U9604 ( .A(n7396), .B(n7398), .Z(n7406) );
  XNOR U9605 ( .A(n7392), .B(n7407), .Z(n7398) );
  XNOR U9606 ( .A(n7390), .B(n7393), .Z(n7407) );
  NAND U9607 ( .A(n7408), .B(n7409), .Z(n7393) );
  NAND U9608 ( .A(n7410), .B(n7411), .Z(n7409) );
  OR U9609 ( .A(n7412), .B(n7413), .Z(n7410) );
  NANDN U9610 ( .A(n7414), .B(n7412), .Z(n7408) );
  IV U9611 ( .A(n7413), .Z(n7414) );
  NAND U9612 ( .A(n7415), .B(n7416), .Z(n7390) );
  NAND U9613 ( .A(n7417), .B(n7418), .Z(n7416) );
  NANDN U9614 ( .A(n7419), .B(n7420), .Z(n7417) );
  NANDN U9615 ( .A(n7420), .B(n7419), .Z(n7415) );
  AND U9616 ( .A(n7421), .B(n7422), .Z(n7392) );
  NAND U9617 ( .A(n7423), .B(n7424), .Z(n7422) );
  OR U9618 ( .A(n7425), .B(n7426), .Z(n7423) );
  NANDN U9619 ( .A(n7427), .B(n7425), .Z(n7421) );
  NAND U9620 ( .A(n7428), .B(n7429), .Z(n7396) );
  NANDN U9621 ( .A(n7430), .B(n7431), .Z(n7429) );
  OR U9622 ( .A(n7432), .B(n7433), .Z(n7431) );
  NANDN U9623 ( .A(n7434), .B(n7432), .Z(n7428) );
  IV U9624 ( .A(n7433), .Z(n7434) );
  XNOR U9625 ( .A(n7404), .B(n7435), .Z(n7399) );
  XNOR U9626 ( .A(n7402), .B(n7405), .Z(n7435) );
  NAND U9627 ( .A(n7436), .B(n7437), .Z(n7405) );
  NAND U9628 ( .A(n7438), .B(n7439), .Z(n7437) );
  OR U9629 ( .A(n7440), .B(n7441), .Z(n7438) );
  NANDN U9630 ( .A(n7442), .B(n7440), .Z(n7436) );
  IV U9631 ( .A(n7441), .Z(n7442) );
  NAND U9632 ( .A(n7443), .B(n7444), .Z(n7402) );
  NAND U9633 ( .A(n7445), .B(n7446), .Z(n7444) );
  NANDN U9634 ( .A(n7447), .B(n7448), .Z(n7445) );
  NANDN U9635 ( .A(n7448), .B(n7447), .Z(n7443) );
  AND U9636 ( .A(n7449), .B(n7450), .Z(n7404) );
  NAND U9637 ( .A(n7451), .B(n7452), .Z(n7450) );
  OR U9638 ( .A(n7453), .B(n7454), .Z(n7451) );
  NANDN U9639 ( .A(n7455), .B(n7453), .Z(n7449) );
  XNOR U9640 ( .A(n7430), .B(n7456), .Z(N13233) );
  XOR U9641 ( .A(n7432), .B(n7433), .Z(n7456) );
  XNOR U9642 ( .A(n7446), .B(n7457), .Z(n7433) );
  XOR U9643 ( .A(n7447), .B(n7448), .Z(n7457) );
  XOR U9644 ( .A(n7453), .B(n7458), .Z(n7448) );
  XOR U9645 ( .A(n7452), .B(n7455), .Z(n7458) );
  IV U9646 ( .A(n7454), .Z(n7455) );
  NAND U9647 ( .A(n7459), .B(n7460), .Z(n7454) );
  OR U9648 ( .A(n7461), .B(n7462), .Z(n7460) );
  OR U9649 ( .A(n7463), .B(n7464), .Z(n7459) );
  NAND U9650 ( .A(n7465), .B(n7466), .Z(n7452) );
  OR U9651 ( .A(n7467), .B(n7468), .Z(n7466) );
  OR U9652 ( .A(n7469), .B(n7470), .Z(n7465) );
  NOR U9653 ( .A(n7471), .B(n7472), .Z(n7453) );
  ANDN U9654 ( .B(n7473), .A(n7474), .Z(n7447) );
  XNOR U9655 ( .A(n7440), .B(n7475), .Z(n7446) );
  XNOR U9656 ( .A(n7439), .B(n7441), .Z(n7475) );
  NAND U9657 ( .A(n7476), .B(n7477), .Z(n7441) );
  OR U9658 ( .A(n7478), .B(n7479), .Z(n7477) );
  OR U9659 ( .A(n7480), .B(n7481), .Z(n7476) );
  NAND U9660 ( .A(n7482), .B(n7483), .Z(n7439) );
  OR U9661 ( .A(n7484), .B(n7485), .Z(n7483) );
  OR U9662 ( .A(n7486), .B(n7487), .Z(n7482) );
  ANDN U9663 ( .B(n7488), .A(n7489), .Z(n7440) );
  IV U9664 ( .A(n7490), .Z(n7488) );
  ANDN U9665 ( .B(n7491), .A(n7492), .Z(n7432) );
  XOR U9666 ( .A(n7418), .B(n7493), .Z(n7430) );
  XOR U9667 ( .A(n7419), .B(n7420), .Z(n7493) );
  XOR U9668 ( .A(n7425), .B(n7494), .Z(n7420) );
  XOR U9669 ( .A(n7424), .B(n7427), .Z(n7494) );
  IV U9670 ( .A(n7426), .Z(n7427) );
  NAND U9671 ( .A(n7495), .B(n7496), .Z(n7426) );
  OR U9672 ( .A(n7497), .B(n7498), .Z(n7496) );
  OR U9673 ( .A(n7499), .B(n7500), .Z(n7495) );
  NAND U9674 ( .A(n7501), .B(n7502), .Z(n7424) );
  OR U9675 ( .A(n7503), .B(n7504), .Z(n7502) );
  OR U9676 ( .A(n7505), .B(n7506), .Z(n7501) );
  NOR U9677 ( .A(n7507), .B(n7508), .Z(n7425) );
  ANDN U9678 ( .B(n7509), .A(n7510), .Z(n7419) );
  IV U9679 ( .A(n7511), .Z(n7509) );
  XNOR U9680 ( .A(n7412), .B(n7512), .Z(n7418) );
  XNOR U9681 ( .A(n7411), .B(n7413), .Z(n7512) );
  NAND U9682 ( .A(n7513), .B(n7514), .Z(n7413) );
  OR U9683 ( .A(n7515), .B(n7516), .Z(n7514) );
  OR U9684 ( .A(n7517), .B(n7518), .Z(n7513) );
  NAND U9685 ( .A(n7519), .B(n7520), .Z(n7411) );
  OR U9686 ( .A(n7521), .B(n7522), .Z(n7520) );
  OR U9687 ( .A(n7523), .B(n7524), .Z(n7519) );
  ANDN U9688 ( .B(n7525), .A(n7526), .Z(n7412) );
  IV U9689 ( .A(n7527), .Z(n7525) );
  XNOR U9690 ( .A(n7492), .B(n7491), .Z(N13232) );
  XOR U9691 ( .A(n7511), .B(n7510), .Z(n7491) );
  XNOR U9692 ( .A(n7526), .B(n7527), .Z(n7510) );
  XNOR U9693 ( .A(n7521), .B(n7522), .Z(n7527) );
  XNOR U9694 ( .A(n7523), .B(n7524), .Z(n7522) );
  XNOR U9695 ( .A(y[997]), .B(x[997]), .Z(n7524) );
  XNOR U9696 ( .A(y[998]), .B(x[998]), .Z(n7523) );
  XNOR U9697 ( .A(y[996]), .B(x[996]), .Z(n7521) );
  XNOR U9698 ( .A(n7515), .B(n7516), .Z(n7526) );
  XNOR U9699 ( .A(y[993]), .B(x[993]), .Z(n7516) );
  XNOR U9700 ( .A(n7517), .B(n7518), .Z(n7515) );
  XNOR U9701 ( .A(y[994]), .B(x[994]), .Z(n7518) );
  XNOR U9702 ( .A(y[995]), .B(x[995]), .Z(n7517) );
  XNOR U9703 ( .A(n7508), .B(n7507), .Z(n7511) );
  XNOR U9704 ( .A(n7503), .B(n7504), .Z(n7507) );
  XNOR U9705 ( .A(y[990]), .B(x[990]), .Z(n7504) );
  XNOR U9706 ( .A(n7505), .B(n7506), .Z(n7503) );
  XNOR U9707 ( .A(y[991]), .B(x[991]), .Z(n7506) );
  XNOR U9708 ( .A(y[992]), .B(x[992]), .Z(n7505) );
  XNOR U9709 ( .A(n7497), .B(n7498), .Z(n7508) );
  XNOR U9710 ( .A(y[987]), .B(x[987]), .Z(n7498) );
  XNOR U9711 ( .A(n7499), .B(n7500), .Z(n7497) );
  XNOR U9712 ( .A(y[988]), .B(x[988]), .Z(n7500) );
  XNOR U9713 ( .A(y[989]), .B(x[989]), .Z(n7499) );
  XOR U9714 ( .A(n7473), .B(n7474), .Z(n7492) );
  XNOR U9715 ( .A(n7489), .B(n7490), .Z(n7474) );
  XNOR U9716 ( .A(n7484), .B(n7485), .Z(n7490) );
  XNOR U9717 ( .A(n7486), .B(n7487), .Z(n7485) );
  XNOR U9718 ( .A(y[985]), .B(x[985]), .Z(n7487) );
  XNOR U9719 ( .A(y[986]), .B(x[986]), .Z(n7486) );
  XNOR U9720 ( .A(y[984]), .B(x[984]), .Z(n7484) );
  XNOR U9721 ( .A(n7478), .B(n7479), .Z(n7489) );
  XNOR U9722 ( .A(y[981]), .B(x[981]), .Z(n7479) );
  XNOR U9723 ( .A(n7480), .B(n7481), .Z(n7478) );
  XNOR U9724 ( .A(y[982]), .B(x[982]), .Z(n7481) );
  XNOR U9725 ( .A(y[983]), .B(x[983]), .Z(n7480) );
  XOR U9726 ( .A(n7472), .B(n7471), .Z(n7473) );
  XNOR U9727 ( .A(n7467), .B(n7468), .Z(n7471) );
  XNOR U9728 ( .A(y[978]), .B(x[978]), .Z(n7468) );
  XNOR U9729 ( .A(n7469), .B(n7470), .Z(n7467) );
  XNOR U9730 ( .A(y[979]), .B(x[979]), .Z(n7470) );
  XNOR U9731 ( .A(y[980]), .B(x[980]), .Z(n7469) );
  XNOR U9732 ( .A(n7461), .B(n7462), .Z(n7472) );
  XNOR U9733 ( .A(y[975]), .B(x[975]), .Z(n7462) );
  XNOR U9734 ( .A(n7463), .B(n7464), .Z(n7461) );
  XNOR U9735 ( .A(y[976]), .B(x[976]), .Z(n7464) );
  XNOR U9736 ( .A(y[977]), .B(x[977]), .Z(n7463) );
  NAND U9737 ( .A(n7528), .B(n7529), .Z(N13225) );
  NANDN U9738 ( .A(n7530), .B(n7531), .Z(n7529) );
  OR U9739 ( .A(n7532), .B(n7533), .Z(n7531) );
  NAND U9740 ( .A(n7532), .B(n7533), .Z(n7528) );
  XOR U9741 ( .A(n7532), .B(n7534), .Z(N13224) );
  XNOR U9742 ( .A(n7530), .B(n7533), .Z(n7534) );
  AND U9743 ( .A(n7535), .B(n7536), .Z(n7533) );
  NANDN U9744 ( .A(n7537), .B(n7538), .Z(n7536) );
  NANDN U9745 ( .A(n7539), .B(n7540), .Z(n7538) );
  NANDN U9746 ( .A(n7540), .B(n7539), .Z(n7535) );
  NAND U9747 ( .A(n7541), .B(n7542), .Z(n7530) );
  NANDN U9748 ( .A(n7543), .B(n7544), .Z(n7542) );
  OR U9749 ( .A(n7545), .B(n7546), .Z(n7544) );
  NAND U9750 ( .A(n7546), .B(n7545), .Z(n7541) );
  AND U9751 ( .A(n7547), .B(n7548), .Z(n7532) );
  NANDN U9752 ( .A(n7549), .B(n7550), .Z(n7548) );
  NANDN U9753 ( .A(n7551), .B(n7552), .Z(n7550) );
  NANDN U9754 ( .A(n7552), .B(n7551), .Z(n7547) );
  XOR U9755 ( .A(n7546), .B(n7553), .Z(N13223) );
  XOR U9756 ( .A(n7543), .B(n7545), .Z(n7553) );
  XNOR U9757 ( .A(n7539), .B(n7554), .Z(n7545) );
  XNOR U9758 ( .A(n7537), .B(n7540), .Z(n7554) );
  NAND U9759 ( .A(n7555), .B(n7556), .Z(n7540) );
  NAND U9760 ( .A(n7557), .B(n7558), .Z(n7556) );
  OR U9761 ( .A(n7559), .B(n7560), .Z(n7557) );
  NANDN U9762 ( .A(n7561), .B(n7559), .Z(n7555) );
  IV U9763 ( .A(n7560), .Z(n7561) );
  NAND U9764 ( .A(n7562), .B(n7563), .Z(n7537) );
  NAND U9765 ( .A(n7564), .B(n7565), .Z(n7563) );
  NANDN U9766 ( .A(n7566), .B(n7567), .Z(n7564) );
  NANDN U9767 ( .A(n7567), .B(n7566), .Z(n7562) );
  AND U9768 ( .A(n7568), .B(n7569), .Z(n7539) );
  NAND U9769 ( .A(n7570), .B(n7571), .Z(n7569) );
  OR U9770 ( .A(n7572), .B(n7573), .Z(n7570) );
  NANDN U9771 ( .A(n7574), .B(n7572), .Z(n7568) );
  NAND U9772 ( .A(n7575), .B(n7576), .Z(n7543) );
  NANDN U9773 ( .A(n7577), .B(n7578), .Z(n7576) );
  OR U9774 ( .A(n7579), .B(n7580), .Z(n7578) );
  NANDN U9775 ( .A(n7581), .B(n7579), .Z(n7575) );
  IV U9776 ( .A(n7580), .Z(n7581) );
  XNOR U9777 ( .A(n7551), .B(n7582), .Z(n7546) );
  XNOR U9778 ( .A(n7549), .B(n7552), .Z(n7582) );
  NAND U9779 ( .A(n7583), .B(n7584), .Z(n7552) );
  NAND U9780 ( .A(n7585), .B(n7586), .Z(n7584) );
  OR U9781 ( .A(n7587), .B(n7588), .Z(n7585) );
  NANDN U9782 ( .A(n7589), .B(n7587), .Z(n7583) );
  IV U9783 ( .A(n7588), .Z(n7589) );
  NAND U9784 ( .A(n7590), .B(n7591), .Z(n7549) );
  NAND U9785 ( .A(n7592), .B(n7593), .Z(n7591) );
  NANDN U9786 ( .A(n7594), .B(n7595), .Z(n7592) );
  NANDN U9787 ( .A(n7595), .B(n7594), .Z(n7590) );
  AND U9788 ( .A(n7596), .B(n7597), .Z(n7551) );
  NAND U9789 ( .A(n7598), .B(n7599), .Z(n7597) );
  OR U9790 ( .A(n7600), .B(n7601), .Z(n7598) );
  NANDN U9791 ( .A(n7602), .B(n7600), .Z(n7596) );
  XNOR U9792 ( .A(n7577), .B(n7603), .Z(N13222) );
  XOR U9793 ( .A(n7579), .B(n7580), .Z(n7603) );
  XNOR U9794 ( .A(n7593), .B(n7604), .Z(n7580) );
  XOR U9795 ( .A(n7594), .B(n7595), .Z(n7604) );
  XOR U9796 ( .A(n7600), .B(n7605), .Z(n7595) );
  XOR U9797 ( .A(n7599), .B(n7602), .Z(n7605) );
  IV U9798 ( .A(n7601), .Z(n7602) );
  NAND U9799 ( .A(n7606), .B(n7607), .Z(n7601) );
  OR U9800 ( .A(n7608), .B(n7609), .Z(n7607) );
  OR U9801 ( .A(n7610), .B(n7611), .Z(n7606) );
  NAND U9802 ( .A(n7612), .B(n7613), .Z(n7599) );
  OR U9803 ( .A(n7614), .B(n7615), .Z(n7613) );
  OR U9804 ( .A(n7616), .B(n7617), .Z(n7612) );
  NOR U9805 ( .A(n7618), .B(n7619), .Z(n7600) );
  ANDN U9806 ( .B(n7620), .A(n7621), .Z(n7594) );
  XNOR U9807 ( .A(n7587), .B(n7622), .Z(n7593) );
  XNOR U9808 ( .A(n7586), .B(n7588), .Z(n7622) );
  NAND U9809 ( .A(n7623), .B(n7624), .Z(n7588) );
  OR U9810 ( .A(n7625), .B(n7626), .Z(n7624) );
  OR U9811 ( .A(n7627), .B(n7628), .Z(n7623) );
  NAND U9812 ( .A(n7629), .B(n7630), .Z(n7586) );
  OR U9813 ( .A(n7631), .B(n7632), .Z(n7630) );
  OR U9814 ( .A(n7633), .B(n7634), .Z(n7629) );
  ANDN U9815 ( .B(n7635), .A(n7636), .Z(n7587) );
  IV U9816 ( .A(n7637), .Z(n7635) );
  ANDN U9817 ( .B(n7638), .A(n7639), .Z(n7579) );
  XOR U9818 ( .A(n7565), .B(n7640), .Z(n7577) );
  XOR U9819 ( .A(n7566), .B(n7567), .Z(n7640) );
  XOR U9820 ( .A(n7572), .B(n7641), .Z(n7567) );
  XOR U9821 ( .A(n7571), .B(n7574), .Z(n7641) );
  IV U9822 ( .A(n7573), .Z(n7574) );
  NAND U9823 ( .A(n7642), .B(n7643), .Z(n7573) );
  OR U9824 ( .A(n7644), .B(n7645), .Z(n7643) );
  OR U9825 ( .A(n7646), .B(n7647), .Z(n7642) );
  NAND U9826 ( .A(n7648), .B(n7649), .Z(n7571) );
  OR U9827 ( .A(n7650), .B(n7651), .Z(n7649) );
  OR U9828 ( .A(n7652), .B(n7653), .Z(n7648) );
  NOR U9829 ( .A(n7654), .B(n7655), .Z(n7572) );
  ANDN U9830 ( .B(n7656), .A(n7657), .Z(n7566) );
  IV U9831 ( .A(n7658), .Z(n7656) );
  XNOR U9832 ( .A(n7559), .B(n7659), .Z(n7565) );
  XNOR U9833 ( .A(n7558), .B(n7560), .Z(n7659) );
  NAND U9834 ( .A(n7660), .B(n7661), .Z(n7560) );
  OR U9835 ( .A(n7662), .B(n7663), .Z(n7661) );
  OR U9836 ( .A(n7664), .B(n7665), .Z(n7660) );
  NAND U9837 ( .A(n7666), .B(n7667), .Z(n7558) );
  OR U9838 ( .A(n7668), .B(n7669), .Z(n7667) );
  OR U9839 ( .A(n7670), .B(n7671), .Z(n7666) );
  ANDN U9840 ( .B(n7672), .A(n7673), .Z(n7559) );
  IV U9841 ( .A(n7674), .Z(n7672) );
  XNOR U9842 ( .A(n7639), .B(n7638), .Z(N13221) );
  XOR U9843 ( .A(n7658), .B(n7657), .Z(n7638) );
  XNOR U9844 ( .A(n7673), .B(n7674), .Z(n7657) );
  XNOR U9845 ( .A(n7668), .B(n7669), .Z(n7674) );
  XNOR U9846 ( .A(n7670), .B(n7671), .Z(n7669) );
  XNOR U9847 ( .A(y[973]), .B(x[973]), .Z(n7671) );
  XNOR U9848 ( .A(y[974]), .B(x[974]), .Z(n7670) );
  XNOR U9849 ( .A(y[972]), .B(x[972]), .Z(n7668) );
  XNOR U9850 ( .A(n7662), .B(n7663), .Z(n7673) );
  XNOR U9851 ( .A(y[969]), .B(x[969]), .Z(n7663) );
  XNOR U9852 ( .A(n7664), .B(n7665), .Z(n7662) );
  XNOR U9853 ( .A(y[970]), .B(x[970]), .Z(n7665) );
  XNOR U9854 ( .A(y[971]), .B(x[971]), .Z(n7664) );
  XNOR U9855 ( .A(n7655), .B(n7654), .Z(n7658) );
  XNOR U9856 ( .A(n7650), .B(n7651), .Z(n7654) );
  XNOR U9857 ( .A(y[966]), .B(x[966]), .Z(n7651) );
  XNOR U9858 ( .A(n7652), .B(n7653), .Z(n7650) );
  XNOR U9859 ( .A(y[967]), .B(x[967]), .Z(n7653) );
  XNOR U9860 ( .A(y[968]), .B(x[968]), .Z(n7652) );
  XNOR U9861 ( .A(n7644), .B(n7645), .Z(n7655) );
  XNOR U9862 ( .A(y[963]), .B(x[963]), .Z(n7645) );
  XNOR U9863 ( .A(n7646), .B(n7647), .Z(n7644) );
  XNOR U9864 ( .A(y[964]), .B(x[964]), .Z(n7647) );
  XNOR U9865 ( .A(y[965]), .B(x[965]), .Z(n7646) );
  XOR U9866 ( .A(n7620), .B(n7621), .Z(n7639) );
  XNOR U9867 ( .A(n7636), .B(n7637), .Z(n7621) );
  XNOR U9868 ( .A(n7631), .B(n7632), .Z(n7637) );
  XNOR U9869 ( .A(n7633), .B(n7634), .Z(n7632) );
  XNOR U9870 ( .A(y[961]), .B(x[961]), .Z(n7634) );
  XNOR U9871 ( .A(y[962]), .B(x[962]), .Z(n7633) );
  XNOR U9872 ( .A(y[960]), .B(x[960]), .Z(n7631) );
  XNOR U9873 ( .A(n7625), .B(n7626), .Z(n7636) );
  XNOR U9874 ( .A(y[957]), .B(x[957]), .Z(n7626) );
  XNOR U9875 ( .A(n7627), .B(n7628), .Z(n7625) );
  XNOR U9876 ( .A(y[958]), .B(x[958]), .Z(n7628) );
  XNOR U9877 ( .A(y[959]), .B(x[959]), .Z(n7627) );
  XOR U9878 ( .A(n7619), .B(n7618), .Z(n7620) );
  XNOR U9879 ( .A(n7614), .B(n7615), .Z(n7618) );
  XNOR U9880 ( .A(y[954]), .B(x[954]), .Z(n7615) );
  XNOR U9881 ( .A(n7616), .B(n7617), .Z(n7614) );
  XNOR U9882 ( .A(y[955]), .B(x[955]), .Z(n7617) );
  XNOR U9883 ( .A(y[956]), .B(x[956]), .Z(n7616) );
  XNOR U9884 ( .A(n7608), .B(n7609), .Z(n7619) );
  XNOR U9885 ( .A(y[951]), .B(x[951]), .Z(n7609) );
  XNOR U9886 ( .A(n7610), .B(n7611), .Z(n7608) );
  XNOR U9887 ( .A(y[952]), .B(x[952]), .Z(n7611) );
  XNOR U9888 ( .A(y[953]), .B(x[953]), .Z(n7610) );
  NAND U9889 ( .A(n7675), .B(n7676), .Z(N13214) );
  NANDN U9890 ( .A(n7677), .B(n7678), .Z(n7676) );
  OR U9891 ( .A(n7679), .B(n7680), .Z(n7678) );
  NAND U9892 ( .A(n7679), .B(n7680), .Z(n7675) );
  XOR U9893 ( .A(n7679), .B(n7681), .Z(N13213) );
  XNOR U9894 ( .A(n7677), .B(n7680), .Z(n7681) );
  AND U9895 ( .A(n7682), .B(n7683), .Z(n7680) );
  NANDN U9896 ( .A(n7684), .B(n7685), .Z(n7683) );
  NANDN U9897 ( .A(n7686), .B(n7687), .Z(n7685) );
  NANDN U9898 ( .A(n7687), .B(n7686), .Z(n7682) );
  NAND U9899 ( .A(n7688), .B(n7689), .Z(n7677) );
  NANDN U9900 ( .A(n7690), .B(n7691), .Z(n7689) );
  OR U9901 ( .A(n7692), .B(n7693), .Z(n7691) );
  NAND U9902 ( .A(n7693), .B(n7692), .Z(n7688) );
  AND U9903 ( .A(n7694), .B(n7695), .Z(n7679) );
  NANDN U9904 ( .A(n7696), .B(n7697), .Z(n7695) );
  NANDN U9905 ( .A(n7698), .B(n7699), .Z(n7697) );
  NANDN U9906 ( .A(n7699), .B(n7698), .Z(n7694) );
  XOR U9907 ( .A(n7693), .B(n7700), .Z(N13212) );
  XOR U9908 ( .A(n7690), .B(n7692), .Z(n7700) );
  XNOR U9909 ( .A(n7686), .B(n7701), .Z(n7692) );
  XNOR U9910 ( .A(n7684), .B(n7687), .Z(n7701) );
  NAND U9911 ( .A(n7702), .B(n7703), .Z(n7687) );
  NAND U9912 ( .A(n7704), .B(n7705), .Z(n7703) );
  OR U9913 ( .A(n7706), .B(n7707), .Z(n7704) );
  NANDN U9914 ( .A(n7708), .B(n7706), .Z(n7702) );
  IV U9915 ( .A(n7707), .Z(n7708) );
  NAND U9916 ( .A(n7709), .B(n7710), .Z(n7684) );
  NAND U9917 ( .A(n7711), .B(n7712), .Z(n7710) );
  NANDN U9918 ( .A(n7713), .B(n7714), .Z(n7711) );
  NANDN U9919 ( .A(n7714), .B(n7713), .Z(n7709) );
  AND U9920 ( .A(n7715), .B(n7716), .Z(n7686) );
  NAND U9921 ( .A(n7717), .B(n7718), .Z(n7716) );
  OR U9922 ( .A(n7719), .B(n7720), .Z(n7717) );
  NANDN U9923 ( .A(n7721), .B(n7719), .Z(n7715) );
  NAND U9924 ( .A(n7722), .B(n7723), .Z(n7690) );
  NANDN U9925 ( .A(n7724), .B(n7725), .Z(n7723) );
  OR U9926 ( .A(n7726), .B(n7727), .Z(n7725) );
  NANDN U9927 ( .A(n7728), .B(n7726), .Z(n7722) );
  IV U9928 ( .A(n7727), .Z(n7728) );
  XNOR U9929 ( .A(n7698), .B(n7729), .Z(n7693) );
  XNOR U9930 ( .A(n7696), .B(n7699), .Z(n7729) );
  NAND U9931 ( .A(n7730), .B(n7731), .Z(n7699) );
  NAND U9932 ( .A(n7732), .B(n7733), .Z(n7731) );
  OR U9933 ( .A(n7734), .B(n7735), .Z(n7732) );
  NANDN U9934 ( .A(n7736), .B(n7734), .Z(n7730) );
  IV U9935 ( .A(n7735), .Z(n7736) );
  NAND U9936 ( .A(n7737), .B(n7738), .Z(n7696) );
  NAND U9937 ( .A(n7739), .B(n7740), .Z(n7738) );
  NANDN U9938 ( .A(n7741), .B(n7742), .Z(n7739) );
  NANDN U9939 ( .A(n7742), .B(n7741), .Z(n7737) );
  AND U9940 ( .A(n7743), .B(n7744), .Z(n7698) );
  NAND U9941 ( .A(n7745), .B(n7746), .Z(n7744) );
  OR U9942 ( .A(n7747), .B(n7748), .Z(n7745) );
  NANDN U9943 ( .A(n7749), .B(n7747), .Z(n7743) );
  XNOR U9944 ( .A(n7724), .B(n7750), .Z(N13211) );
  XOR U9945 ( .A(n7726), .B(n7727), .Z(n7750) );
  XNOR U9946 ( .A(n7740), .B(n7751), .Z(n7727) );
  XOR U9947 ( .A(n7741), .B(n7742), .Z(n7751) );
  XOR U9948 ( .A(n7747), .B(n7752), .Z(n7742) );
  XOR U9949 ( .A(n7746), .B(n7749), .Z(n7752) );
  IV U9950 ( .A(n7748), .Z(n7749) );
  NAND U9951 ( .A(n7753), .B(n7754), .Z(n7748) );
  OR U9952 ( .A(n7755), .B(n7756), .Z(n7754) );
  OR U9953 ( .A(n7757), .B(n7758), .Z(n7753) );
  NAND U9954 ( .A(n7759), .B(n7760), .Z(n7746) );
  OR U9955 ( .A(n7761), .B(n7762), .Z(n7760) );
  OR U9956 ( .A(n7763), .B(n7764), .Z(n7759) );
  NOR U9957 ( .A(n7765), .B(n7766), .Z(n7747) );
  ANDN U9958 ( .B(n7767), .A(n7768), .Z(n7741) );
  XNOR U9959 ( .A(n7734), .B(n7769), .Z(n7740) );
  XNOR U9960 ( .A(n7733), .B(n7735), .Z(n7769) );
  NAND U9961 ( .A(n7770), .B(n7771), .Z(n7735) );
  OR U9962 ( .A(n7772), .B(n7773), .Z(n7771) );
  OR U9963 ( .A(n7774), .B(n7775), .Z(n7770) );
  NAND U9964 ( .A(n7776), .B(n7777), .Z(n7733) );
  OR U9965 ( .A(n7778), .B(n7779), .Z(n7777) );
  OR U9966 ( .A(n7780), .B(n7781), .Z(n7776) );
  ANDN U9967 ( .B(n7782), .A(n7783), .Z(n7734) );
  IV U9968 ( .A(n7784), .Z(n7782) );
  ANDN U9969 ( .B(n7785), .A(n7786), .Z(n7726) );
  XOR U9970 ( .A(n7712), .B(n7787), .Z(n7724) );
  XOR U9971 ( .A(n7713), .B(n7714), .Z(n7787) );
  XOR U9972 ( .A(n7719), .B(n7788), .Z(n7714) );
  XOR U9973 ( .A(n7718), .B(n7721), .Z(n7788) );
  IV U9974 ( .A(n7720), .Z(n7721) );
  NAND U9975 ( .A(n7789), .B(n7790), .Z(n7720) );
  OR U9976 ( .A(n7791), .B(n7792), .Z(n7790) );
  OR U9977 ( .A(n7793), .B(n7794), .Z(n7789) );
  NAND U9978 ( .A(n7795), .B(n7796), .Z(n7718) );
  OR U9979 ( .A(n7797), .B(n7798), .Z(n7796) );
  OR U9980 ( .A(n7799), .B(n7800), .Z(n7795) );
  NOR U9981 ( .A(n7801), .B(n7802), .Z(n7719) );
  ANDN U9982 ( .B(n7803), .A(n7804), .Z(n7713) );
  IV U9983 ( .A(n7805), .Z(n7803) );
  XNOR U9984 ( .A(n7706), .B(n7806), .Z(n7712) );
  XNOR U9985 ( .A(n7705), .B(n7707), .Z(n7806) );
  NAND U9986 ( .A(n7807), .B(n7808), .Z(n7707) );
  OR U9987 ( .A(n7809), .B(n7810), .Z(n7808) );
  OR U9988 ( .A(n7811), .B(n7812), .Z(n7807) );
  NAND U9989 ( .A(n7813), .B(n7814), .Z(n7705) );
  OR U9990 ( .A(n7815), .B(n7816), .Z(n7814) );
  OR U9991 ( .A(n7817), .B(n7818), .Z(n7813) );
  ANDN U9992 ( .B(n7819), .A(n7820), .Z(n7706) );
  IV U9993 ( .A(n7821), .Z(n7819) );
  XNOR U9994 ( .A(n7786), .B(n7785), .Z(N13210) );
  XOR U9995 ( .A(n7805), .B(n7804), .Z(n7785) );
  XNOR U9996 ( .A(n7820), .B(n7821), .Z(n7804) );
  XNOR U9997 ( .A(n7815), .B(n7816), .Z(n7821) );
  XNOR U9998 ( .A(n7817), .B(n7818), .Z(n7816) );
  XNOR U9999 ( .A(y[949]), .B(x[949]), .Z(n7818) );
  XNOR U10000 ( .A(y[950]), .B(x[950]), .Z(n7817) );
  XNOR U10001 ( .A(y[948]), .B(x[948]), .Z(n7815) );
  XNOR U10002 ( .A(n7809), .B(n7810), .Z(n7820) );
  XNOR U10003 ( .A(y[945]), .B(x[945]), .Z(n7810) );
  XNOR U10004 ( .A(n7811), .B(n7812), .Z(n7809) );
  XNOR U10005 ( .A(y[946]), .B(x[946]), .Z(n7812) );
  XNOR U10006 ( .A(y[947]), .B(x[947]), .Z(n7811) );
  XNOR U10007 ( .A(n7802), .B(n7801), .Z(n7805) );
  XNOR U10008 ( .A(n7797), .B(n7798), .Z(n7801) );
  XNOR U10009 ( .A(y[942]), .B(x[942]), .Z(n7798) );
  XNOR U10010 ( .A(n7799), .B(n7800), .Z(n7797) );
  XNOR U10011 ( .A(y[943]), .B(x[943]), .Z(n7800) );
  XNOR U10012 ( .A(y[944]), .B(x[944]), .Z(n7799) );
  XNOR U10013 ( .A(n7791), .B(n7792), .Z(n7802) );
  XNOR U10014 ( .A(y[939]), .B(x[939]), .Z(n7792) );
  XNOR U10015 ( .A(n7793), .B(n7794), .Z(n7791) );
  XNOR U10016 ( .A(y[940]), .B(x[940]), .Z(n7794) );
  XNOR U10017 ( .A(y[941]), .B(x[941]), .Z(n7793) );
  XOR U10018 ( .A(n7767), .B(n7768), .Z(n7786) );
  XNOR U10019 ( .A(n7783), .B(n7784), .Z(n7768) );
  XNOR U10020 ( .A(n7778), .B(n7779), .Z(n7784) );
  XNOR U10021 ( .A(n7780), .B(n7781), .Z(n7779) );
  XNOR U10022 ( .A(y[937]), .B(x[937]), .Z(n7781) );
  XNOR U10023 ( .A(y[938]), .B(x[938]), .Z(n7780) );
  XNOR U10024 ( .A(y[936]), .B(x[936]), .Z(n7778) );
  XNOR U10025 ( .A(n7772), .B(n7773), .Z(n7783) );
  XNOR U10026 ( .A(y[933]), .B(x[933]), .Z(n7773) );
  XNOR U10027 ( .A(n7774), .B(n7775), .Z(n7772) );
  XNOR U10028 ( .A(y[934]), .B(x[934]), .Z(n7775) );
  XNOR U10029 ( .A(y[935]), .B(x[935]), .Z(n7774) );
  XOR U10030 ( .A(n7766), .B(n7765), .Z(n7767) );
  XNOR U10031 ( .A(n7761), .B(n7762), .Z(n7765) );
  XNOR U10032 ( .A(y[930]), .B(x[930]), .Z(n7762) );
  XNOR U10033 ( .A(n7763), .B(n7764), .Z(n7761) );
  XNOR U10034 ( .A(y[931]), .B(x[931]), .Z(n7764) );
  XNOR U10035 ( .A(y[932]), .B(x[932]), .Z(n7763) );
  XNOR U10036 ( .A(n7755), .B(n7756), .Z(n7766) );
  XNOR U10037 ( .A(y[927]), .B(x[927]), .Z(n7756) );
  XNOR U10038 ( .A(n7757), .B(n7758), .Z(n7755) );
  XNOR U10039 ( .A(y[928]), .B(x[928]), .Z(n7758) );
  XNOR U10040 ( .A(y[929]), .B(x[929]), .Z(n7757) );
  NAND U10041 ( .A(n7822), .B(n7823), .Z(N13203) );
  NANDN U10042 ( .A(n7824), .B(n7825), .Z(n7823) );
  OR U10043 ( .A(n7826), .B(n7827), .Z(n7825) );
  NAND U10044 ( .A(n7826), .B(n7827), .Z(n7822) );
  XOR U10045 ( .A(n7826), .B(n7828), .Z(N13202) );
  XNOR U10046 ( .A(n7824), .B(n7827), .Z(n7828) );
  AND U10047 ( .A(n7829), .B(n7830), .Z(n7827) );
  NANDN U10048 ( .A(n7831), .B(n7832), .Z(n7830) );
  NANDN U10049 ( .A(n7833), .B(n7834), .Z(n7832) );
  NANDN U10050 ( .A(n7834), .B(n7833), .Z(n7829) );
  NAND U10051 ( .A(n7835), .B(n7836), .Z(n7824) );
  NANDN U10052 ( .A(n7837), .B(n7838), .Z(n7836) );
  OR U10053 ( .A(n7839), .B(n7840), .Z(n7838) );
  NAND U10054 ( .A(n7840), .B(n7839), .Z(n7835) );
  AND U10055 ( .A(n7841), .B(n7842), .Z(n7826) );
  NANDN U10056 ( .A(n7843), .B(n7844), .Z(n7842) );
  NANDN U10057 ( .A(n7845), .B(n7846), .Z(n7844) );
  NANDN U10058 ( .A(n7846), .B(n7845), .Z(n7841) );
  XOR U10059 ( .A(n7840), .B(n7847), .Z(N13201) );
  XOR U10060 ( .A(n7837), .B(n7839), .Z(n7847) );
  XNOR U10061 ( .A(n7833), .B(n7848), .Z(n7839) );
  XNOR U10062 ( .A(n7831), .B(n7834), .Z(n7848) );
  NAND U10063 ( .A(n7849), .B(n7850), .Z(n7834) );
  NAND U10064 ( .A(n7851), .B(n7852), .Z(n7850) );
  OR U10065 ( .A(n7853), .B(n7854), .Z(n7851) );
  NANDN U10066 ( .A(n7855), .B(n7853), .Z(n7849) );
  IV U10067 ( .A(n7854), .Z(n7855) );
  NAND U10068 ( .A(n7856), .B(n7857), .Z(n7831) );
  NAND U10069 ( .A(n7858), .B(n7859), .Z(n7857) );
  NANDN U10070 ( .A(n7860), .B(n7861), .Z(n7858) );
  NANDN U10071 ( .A(n7861), .B(n7860), .Z(n7856) );
  AND U10072 ( .A(n7862), .B(n7863), .Z(n7833) );
  NAND U10073 ( .A(n7864), .B(n7865), .Z(n7863) );
  OR U10074 ( .A(n7866), .B(n7867), .Z(n7864) );
  NANDN U10075 ( .A(n7868), .B(n7866), .Z(n7862) );
  NAND U10076 ( .A(n7869), .B(n7870), .Z(n7837) );
  NANDN U10077 ( .A(n7871), .B(n7872), .Z(n7870) );
  OR U10078 ( .A(n7873), .B(n7874), .Z(n7872) );
  NANDN U10079 ( .A(n7875), .B(n7873), .Z(n7869) );
  IV U10080 ( .A(n7874), .Z(n7875) );
  XNOR U10081 ( .A(n7845), .B(n7876), .Z(n7840) );
  XNOR U10082 ( .A(n7843), .B(n7846), .Z(n7876) );
  NAND U10083 ( .A(n7877), .B(n7878), .Z(n7846) );
  NAND U10084 ( .A(n7879), .B(n7880), .Z(n7878) );
  OR U10085 ( .A(n7881), .B(n7882), .Z(n7879) );
  NANDN U10086 ( .A(n7883), .B(n7881), .Z(n7877) );
  IV U10087 ( .A(n7882), .Z(n7883) );
  NAND U10088 ( .A(n7884), .B(n7885), .Z(n7843) );
  NAND U10089 ( .A(n7886), .B(n7887), .Z(n7885) );
  NANDN U10090 ( .A(n7888), .B(n7889), .Z(n7886) );
  NANDN U10091 ( .A(n7889), .B(n7888), .Z(n7884) );
  AND U10092 ( .A(n7890), .B(n7891), .Z(n7845) );
  NAND U10093 ( .A(n7892), .B(n7893), .Z(n7891) );
  OR U10094 ( .A(n7894), .B(n7895), .Z(n7892) );
  NANDN U10095 ( .A(n7896), .B(n7894), .Z(n7890) );
  XNOR U10096 ( .A(n7871), .B(n7897), .Z(N13200) );
  XOR U10097 ( .A(n7873), .B(n7874), .Z(n7897) );
  XNOR U10098 ( .A(n7887), .B(n7898), .Z(n7874) );
  XOR U10099 ( .A(n7888), .B(n7889), .Z(n7898) );
  XOR U10100 ( .A(n7894), .B(n7899), .Z(n7889) );
  XOR U10101 ( .A(n7893), .B(n7896), .Z(n7899) );
  IV U10102 ( .A(n7895), .Z(n7896) );
  NAND U10103 ( .A(n7900), .B(n7901), .Z(n7895) );
  OR U10104 ( .A(n7902), .B(n7903), .Z(n7901) );
  OR U10105 ( .A(n7904), .B(n7905), .Z(n7900) );
  NAND U10106 ( .A(n7906), .B(n7907), .Z(n7893) );
  OR U10107 ( .A(n7908), .B(n7909), .Z(n7907) );
  OR U10108 ( .A(n7910), .B(n7911), .Z(n7906) );
  NOR U10109 ( .A(n7912), .B(n7913), .Z(n7894) );
  ANDN U10110 ( .B(n7914), .A(n7915), .Z(n7888) );
  XNOR U10111 ( .A(n7881), .B(n7916), .Z(n7887) );
  XNOR U10112 ( .A(n7880), .B(n7882), .Z(n7916) );
  NAND U10113 ( .A(n7917), .B(n7918), .Z(n7882) );
  OR U10114 ( .A(n7919), .B(n7920), .Z(n7918) );
  OR U10115 ( .A(n7921), .B(n7922), .Z(n7917) );
  NAND U10116 ( .A(n7923), .B(n7924), .Z(n7880) );
  OR U10117 ( .A(n7925), .B(n7926), .Z(n7924) );
  OR U10118 ( .A(n7927), .B(n7928), .Z(n7923) );
  ANDN U10119 ( .B(n7929), .A(n7930), .Z(n7881) );
  IV U10120 ( .A(n7931), .Z(n7929) );
  ANDN U10121 ( .B(n7932), .A(n7933), .Z(n7873) );
  XOR U10122 ( .A(n7859), .B(n7934), .Z(n7871) );
  XOR U10123 ( .A(n7860), .B(n7861), .Z(n7934) );
  XOR U10124 ( .A(n7866), .B(n7935), .Z(n7861) );
  XOR U10125 ( .A(n7865), .B(n7868), .Z(n7935) );
  IV U10126 ( .A(n7867), .Z(n7868) );
  NAND U10127 ( .A(n7936), .B(n7937), .Z(n7867) );
  OR U10128 ( .A(n7938), .B(n7939), .Z(n7937) );
  OR U10129 ( .A(n7940), .B(n7941), .Z(n7936) );
  NAND U10130 ( .A(n7942), .B(n7943), .Z(n7865) );
  OR U10131 ( .A(n7944), .B(n7945), .Z(n7943) );
  OR U10132 ( .A(n7946), .B(n7947), .Z(n7942) );
  NOR U10133 ( .A(n7948), .B(n7949), .Z(n7866) );
  ANDN U10134 ( .B(n7950), .A(n7951), .Z(n7860) );
  IV U10135 ( .A(n7952), .Z(n7950) );
  XNOR U10136 ( .A(n7853), .B(n7953), .Z(n7859) );
  XNOR U10137 ( .A(n7852), .B(n7854), .Z(n7953) );
  NAND U10138 ( .A(n7954), .B(n7955), .Z(n7854) );
  OR U10139 ( .A(n7956), .B(n7957), .Z(n7955) );
  OR U10140 ( .A(n7958), .B(n7959), .Z(n7954) );
  NAND U10141 ( .A(n7960), .B(n7961), .Z(n7852) );
  OR U10142 ( .A(n7962), .B(n7963), .Z(n7961) );
  OR U10143 ( .A(n7964), .B(n7965), .Z(n7960) );
  ANDN U10144 ( .B(n7966), .A(n7967), .Z(n7853) );
  IV U10145 ( .A(n7968), .Z(n7966) );
  XNOR U10146 ( .A(n7933), .B(n7932), .Z(N13199) );
  XOR U10147 ( .A(n7952), .B(n7951), .Z(n7932) );
  XNOR U10148 ( .A(n7967), .B(n7968), .Z(n7951) );
  XNOR U10149 ( .A(n7962), .B(n7963), .Z(n7968) );
  XNOR U10150 ( .A(n7964), .B(n7965), .Z(n7963) );
  XNOR U10151 ( .A(y[925]), .B(x[925]), .Z(n7965) );
  XNOR U10152 ( .A(y[926]), .B(x[926]), .Z(n7964) );
  XNOR U10153 ( .A(y[924]), .B(x[924]), .Z(n7962) );
  XNOR U10154 ( .A(n7956), .B(n7957), .Z(n7967) );
  XNOR U10155 ( .A(y[921]), .B(x[921]), .Z(n7957) );
  XNOR U10156 ( .A(n7958), .B(n7959), .Z(n7956) );
  XNOR U10157 ( .A(y[922]), .B(x[922]), .Z(n7959) );
  XNOR U10158 ( .A(y[923]), .B(x[923]), .Z(n7958) );
  XNOR U10159 ( .A(n7949), .B(n7948), .Z(n7952) );
  XNOR U10160 ( .A(n7944), .B(n7945), .Z(n7948) );
  XNOR U10161 ( .A(y[918]), .B(x[918]), .Z(n7945) );
  XNOR U10162 ( .A(n7946), .B(n7947), .Z(n7944) );
  XNOR U10163 ( .A(y[919]), .B(x[919]), .Z(n7947) );
  XNOR U10164 ( .A(y[920]), .B(x[920]), .Z(n7946) );
  XNOR U10165 ( .A(n7938), .B(n7939), .Z(n7949) );
  XNOR U10166 ( .A(y[915]), .B(x[915]), .Z(n7939) );
  XNOR U10167 ( .A(n7940), .B(n7941), .Z(n7938) );
  XNOR U10168 ( .A(y[916]), .B(x[916]), .Z(n7941) );
  XNOR U10169 ( .A(y[917]), .B(x[917]), .Z(n7940) );
  XOR U10170 ( .A(n7914), .B(n7915), .Z(n7933) );
  XNOR U10171 ( .A(n7930), .B(n7931), .Z(n7915) );
  XNOR U10172 ( .A(n7925), .B(n7926), .Z(n7931) );
  XNOR U10173 ( .A(n7927), .B(n7928), .Z(n7926) );
  XNOR U10174 ( .A(y[913]), .B(x[913]), .Z(n7928) );
  XNOR U10175 ( .A(y[914]), .B(x[914]), .Z(n7927) );
  XNOR U10176 ( .A(y[912]), .B(x[912]), .Z(n7925) );
  XNOR U10177 ( .A(n7919), .B(n7920), .Z(n7930) );
  XNOR U10178 ( .A(y[909]), .B(x[909]), .Z(n7920) );
  XNOR U10179 ( .A(n7921), .B(n7922), .Z(n7919) );
  XNOR U10180 ( .A(y[910]), .B(x[910]), .Z(n7922) );
  XNOR U10181 ( .A(y[911]), .B(x[911]), .Z(n7921) );
  XOR U10182 ( .A(n7913), .B(n7912), .Z(n7914) );
  XNOR U10183 ( .A(n7908), .B(n7909), .Z(n7912) );
  XNOR U10184 ( .A(y[906]), .B(x[906]), .Z(n7909) );
  XNOR U10185 ( .A(n7910), .B(n7911), .Z(n7908) );
  XNOR U10186 ( .A(y[907]), .B(x[907]), .Z(n7911) );
  XNOR U10187 ( .A(y[908]), .B(x[908]), .Z(n7910) );
  XNOR U10188 ( .A(n7902), .B(n7903), .Z(n7913) );
  XNOR U10189 ( .A(y[903]), .B(x[903]), .Z(n7903) );
  XNOR U10190 ( .A(n7904), .B(n7905), .Z(n7902) );
  XNOR U10191 ( .A(y[904]), .B(x[904]), .Z(n7905) );
  XNOR U10192 ( .A(y[905]), .B(x[905]), .Z(n7904) );
  NAND U10193 ( .A(n7969), .B(n7970), .Z(N13192) );
  NANDN U10194 ( .A(n7971), .B(n7972), .Z(n7970) );
  OR U10195 ( .A(n7973), .B(n7974), .Z(n7972) );
  NAND U10196 ( .A(n7973), .B(n7974), .Z(n7969) );
  XOR U10197 ( .A(n7973), .B(n7975), .Z(N13191) );
  XNOR U10198 ( .A(n7971), .B(n7974), .Z(n7975) );
  AND U10199 ( .A(n7976), .B(n7977), .Z(n7974) );
  NANDN U10200 ( .A(n7978), .B(n7979), .Z(n7977) );
  NANDN U10201 ( .A(n7980), .B(n7981), .Z(n7979) );
  NANDN U10202 ( .A(n7981), .B(n7980), .Z(n7976) );
  NAND U10203 ( .A(n7982), .B(n7983), .Z(n7971) );
  NANDN U10204 ( .A(n7984), .B(n7985), .Z(n7983) );
  OR U10205 ( .A(n7986), .B(n7987), .Z(n7985) );
  NAND U10206 ( .A(n7987), .B(n7986), .Z(n7982) );
  AND U10207 ( .A(n7988), .B(n7989), .Z(n7973) );
  NANDN U10208 ( .A(n7990), .B(n7991), .Z(n7989) );
  NANDN U10209 ( .A(n7992), .B(n7993), .Z(n7991) );
  NANDN U10210 ( .A(n7993), .B(n7992), .Z(n7988) );
  XOR U10211 ( .A(n7987), .B(n7994), .Z(N13190) );
  XOR U10212 ( .A(n7984), .B(n7986), .Z(n7994) );
  XNOR U10213 ( .A(n7980), .B(n7995), .Z(n7986) );
  XNOR U10214 ( .A(n7978), .B(n7981), .Z(n7995) );
  NAND U10215 ( .A(n7996), .B(n7997), .Z(n7981) );
  NAND U10216 ( .A(n7998), .B(n7999), .Z(n7997) );
  OR U10217 ( .A(n8000), .B(n8001), .Z(n7998) );
  NANDN U10218 ( .A(n8002), .B(n8000), .Z(n7996) );
  IV U10219 ( .A(n8001), .Z(n8002) );
  NAND U10220 ( .A(n8003), .B(n8004), .Z(n7978) );
  NAND U10221 ( .A(n8005), .B(n8006), .Z(n8004) );
  NANDN U10222 ( .A(n8007), .B(n8008), .Z(n8005) );
  NANDN U10223 ( .A(n8008), .B(n8007), .Z(n8003) );
  AND U10224 ( .A(n8009), .B(n8010), .Z(n7980) );
  NAND U10225 ( .A(n8011), .B(n8012), .Z(n8010) );
  OR U10226 ( .A(n8013), .B(n8014), .Z(n8011) );
  NANDN U10227 ( .A(n8015), .B(n8013), .Z(n8009) );
  NAND U10228 ( .A(n8016), .B(n8017), .Z(n7984) );
  NANDN U10229 ( .A(n8018), .B(n8019), .Z(n8017) );
  OR U10230 ( .A(n8020), .B(n8021), .Z(n8019) );
  NANDN U10231 ( .A(n8022), .B(n8020), .Z(n8016) );
  IV U10232 ( .A(n8021), .Z(n8022) );
  XNOR U10233 ( .A(n7992), .B(n8023), .Z(n7987) );
  XNOR U10234 ( .A(n7990), .B(n7993), .Z(n8023) );
  NAND U10235 ( .A(n8024), .B(n8025), .Z(n7993) );
  NAND U10236 ( .A(n8026), .B(n8027), .Z(n8025) );
  OR U10237 ( .A(n8028), .B(n8029), .Z(n8026) );
  NANDN U10238 ( .A(n8030), .B(n8028), .Z(n8024) );
  IV U10239 ( .A(n8029), .Z(n8030) );
  NAND U10240 ( .A(n8031), .B(n8032), .Z(n7990) );
  NAND U10241 ( .A(n8033), .B(n8034), .Z(n8032) );
  NANDN U10242 ( .A(n8035), .B(n8036), .Z(n8033) );
  NANDN U10243 ( .A(n8036), .B(n8035), .Z(n8031) );
  AND U10244 ( .A(n8037), .B(n8038), .Z(n7992) );
  NAND U10245 ( .A(n8039), .B(n8040), .Z(n8038) );
  OR U10246 ( .A(n8041), .B(n8042), .Z(n8039) );
  NANDN U10247 ( .A(n8043), .B(n8041), .Z(n8037) );
  XNOR U10248 ( .A(n8018), .B(n8044), .Z(N13189) );
  XOR U10249 ( .A(n8020), .B(n8021), .Z(n8044) );
  XNOR U10250 ( .A(n8034), .B(n8045), .Z(n8021) );
  XOR U10251 ( .A(n8035), .B(n8036), .Z(n8045) );
  XOR U10252 ( .A(n8041), .B(n8046), .Z(n8036) );
  XOR U10253 ( .A(n8040), .B(n8043), .Z(n8046) );
  IV U10254 ( .A(n8042), .Z(n8043) );
  NAND U10255 ( .A(n8047), .B(n8048), .Z(n8042) );
  OR U10256 ( .A(n8049), .B(n8050), .Z(n8048) );
  OR U10257 ( .A(n8051), .B(n8052), .Z(n8047) );
  NAND U10258 ( .A(n8053), .B(n8054), .Z(n8040) );
  OR U10259 ( .A(n8055), .B(n8056), .Z(n8054) );
  OR U10260 ( .A(n8057), .B(n8058), .Z(n8053) );
  NOR U10261 ( .A(n8059), .B(n8060), .Z(n8041) );
  ANDN U10262 ( .B(n8061), .A(n8062), .Z(n8035) );
  XNOR U10263 ( .A(n8028), .B(n8063), .Z(n8034) );
  XNOR U10264 ( .A(n8027), .B(n8029), .Z(n8063) );
  NAND U10265 ( .A(n8064), .B(n8065), .Z(n8029) );
  OR U10266 ( .A(n8066), .B(n8067), .Z(n8065) );
  OR U10267 ( .A(n8068), .B(n8069), .Z(n8064) );
  NAND U10268 ( .A(n8070), .B(n8071), .Z(n8027) );
  OR U10269 ( .A(n8072), .B(n8073), .Z(n8071) );
  OR U10270 ( .A(n8074), .B(n8075), .Z(n8070) );
  ANDN U10271 ( .B(n8076), .A(n8077), .Z(n8028) );
  IV U10272 ( .A(n8078), .Z(n8076) );
  ANDN U10273 ( .B(n8079), .A(n8080), .Z(n8020) );
  XOR U10274 ( .A(n8006), .B(n8081), .Z(n8018) );
  XOR U10275 ( .A(n8007), .B(n8008), .Z(n8081) );
  XOR U10276 ( .A(n8013), .B(n8082), .Z(n8008) );
  XOR U10277 ( .A(n8012), .B(n8015), .Z(n8082) );
  IV U10278 ( .A(n8014), .Z(n8015) );
  NAND U10279 ( .A(n8083), .B(n8084), .Z(n8014) );
  OR U10280 ( .A(n8085), .B(n8086), .Z(n8084) );
  OR U10281 ( .A(n8087), .B(n8088), .Z(n8083) );
  NAND U10282 ( .A(n8089), .B(n8090), .Z(n8012) );
  OR U10283 ( .A(n8091), .B(n8092), .Z(n8090) );
  OR U10284 ( .A(n8093), .B(n8094), .Z(n8089) );
  NOR U10285 ( .A(n8095), .B(n8096), .Z(n8013) );
  ANDN U10286 ( .B(n8097), .A(n8098), .Z(n8007) );
  IV U10287 ( .A(n8099), .Z(n8097) );
  XNOR U10288 ( .A(n8000), .B(n8100), .Z(n8006) );
  XNOR U10289 ( .A(n7999), .B(n8001), .Z(n8100) );
  NAND U10290 ( .A(n8101), .B(n8102), .Z(n8001) );
  OR U10291 ( .A(n8103), .B(n8104), .Z(n8102) );
  OR U10292 ( .A(n8105), .B(n8106), .Z(n8101) );
  NAND U10293 ( .A(n8107), .B(n8108), .Z(n7999) );
  OR U10294 ( .A(n8109), .B(n8110), .Z(n8108) );
  OR U10295 ( .A(n8111), .B(n8112), .Z(n8107) );
  ANDN U10296 ( .B(n8113), .A(n8114), .Z(n8000) );
  IV U10297 ( .A(n8115), .Z(n8113) );
  XNOR U10298 ( .A(n8080), .B(n8079), .Z(N13188) );
  XOR U10299 ( .A(n8099), .B(n8098), .Z(n8079) );
  XNOR U10300 ( .A(n8114), .B(n8115), .Z(n8098) );
  XNOR U10301 ( .A(n8109), .B(n8110), .Z(n8115) );
  XNOR U10302 ( .A(n8111), .B(n8112), .Z(n8110) );
  XNOR U10303 ( .A(y[901]), .B(x[901]), .Z(n8112) );
  XNOR U10304 ( .A(y[902]), .B(x[902]), .Z(n8111) );
  XNOR U10305 ( .A(y[900]), .B(x[900]), .Z(n8109) );
  XNOR U10306 ( .A(n8103), .B(n8104), .Z(n8114) );
  XNOR U10307 ( .A(y[897]), .B(x[897]), .Z(n8104) );
  XNOR U10308 ( .A(n8105), .B(n8106), .Z(n8103) );
  XNOR U10309 ( .A(y[898]), .B(x[898]), .Z(n8106) );
  XNOR U10310 ( .A(y[899]), .B(x[899]), .Z(n8105) );
  XNOR U10311 ( .A(n8096), .B(n8095), .Z(n8099) );
  XNOR U10312 ( .A(n8091), .B(n8092), .Z(n8095) );
  XNOR U10313 ( .A(y[894]), .B(x[894]), .Z(n8092) );
  XNOR U10314 ( .A(n8093), .B(n8094), .Z(n8091) );
  XNOR U10315 ( .A(y[895]), .B(x[895]), .Z(n8094) );
  XNOR U10316 ( .A(y[896]), .B(x[896]), .Z(n8093) );
  XNOR U10317 ( .A(n8085), .B(n8086), .Z(n8096) );
  XNOR U10318 ( .A(y[891]), .B(x[891]), .Z(n8086) );
  XNOR U10319 ( .A(n8087), .B(n8088), .Z(n8085) );
  XNOR U10320 ( .A(y[892]), .B(x[892]), .Z(n8088) );
  XNOR U10321 ( .A(y[893]), .B(x[893]), .Z(n8087) );
  XOR U10322 ( .A(n8061), .B(n8062), .Z(n8080) );
  XNOR U10323 ( .A(n8077), .B(n8078), .Z(n8062) );
  XNOR U10324 ( .A(n8072), .B(n8073), .Z(n8078) );
  XNOR U10325 ( .A(n8074), .B(n8075), .Z(n8073) );
  XNOR U10326 ( .A(y[889]), .B(x[889]), .Z(n8075) );
  XNOR U10327 ( .A(y[890]), .B(x[890]), .Z(n8074) );
  XNOR U10328 ( .A(y[888]), .B(x[888]), .Z(n8072) );
  XNOR U10329 ( .A(n8066), .B(n8067), .Z(n8077) );
  XNOR U10330 ( .A(y[885]), .B(x[885]), .Z(n8067) );
  XNOR U10331 ( .A(n8068), .B(n8069), .Z(n8066) );
  XNOR U10332 ( .A(y[886]), .B(x[886]), .Z(n8069) );
  XNOR U10333 ( .A(y[887]), .B(x[887]), .Z(n8068) );
  XOR U10334 ( .A(n8060), .B(n8059), .Z(n8061) );
  XNOR U10335 ( .A(n8055), .B(n8056), .Z(n8059) );
  XNOR U10336 ( .A(y[882]), .B(x[882]), .Z(n8056) );
  XNOR U10337 ( .A(n8057), .B(n8058), .Z(n8055) );
  XNOR U10338 ( .A(y[883]), .B(x[883]), .Z(n8058) );
  XNOR U10339 ( .A(y[884]), .B(x[884]), .Z(n8057) );
  XNOR U10340 ( .A(n8049), .B(n8050), .Z(n8060) );
  XNOR U10341 ( .A(y[879]), .B(x[879]), .Z(n8050) );
  XNOR U10342 ( .A(n8051), .B(n8052), .Z(n8049) );
  XNOR U10343 ( .A(y[880]), .B(x[880]), .Z(n8052) );
  XNOR U10344 ( .A(y[881]), .B(x[881]), .Z(n8051) );
  NAND U10345 ( .A(n8116), .B(n8117), .Z(N13181) );
  NANDN U10346 ( .A(n8118), .B(n8119), .Z(n8117) );
  OR U10347 ( .A(n8120), .B(n8121), .Z(n8119) );
  NAND U10348 ( .A(n8120), .B(n8121), .Z(n8116) );
  XOR U10349 ( .A(n8120), .B(n8122), .Z(N13180) );
  XNOR U10350 ( .A(n8118), .B(n8121), .Z(n8122) );
  AND U10351 ( .A(n8123), .B(n8124), .Z(n8121) );
  NANDN U10352 ( .A(n8125), .B(n8126), .Z(n8124) );
  NANDN U10353 ( .A(n8127), .B(n8128), .Z(n8126) );
  NANDN U10354 ( .A(n8128), .B(n8127), .Z(n8123) );
  NAND U10355 ( .A(n8129), .B(n8130), .Z(n8118) );
  NANDN U10356 ( .A(n8131), .B(n8132), .Z(n8130) );
  OR U10357 ( .A(n8133), .B(n8134), .Z(n8132) );
  NAND U10358 ( .A(n8134), .B(n8133), .Z(n8129) );
  AND U10359 ( .A(n8135), .B(n8136), .Z(n8120) );
  NANDN U10360 ( .A(n8137), .B(n8138), .Z(n8136) );
  NANDN U10361 ( .A(n8139), .B(n8140), .Z(n8138) );
  NANDN U10362 ( .A(n8140), .B(n8139), .Z(n8135) );
  XOR U10363 ( .A(n8134), .B(n8141), .Z(N13179) );
  XOR U10364 ( .A(n8131), .B(n8133), .Z(n8141) );
  XNOR U10365 ( .A(n8127), .B(n8142), .Z(n8133) );
  XNOR U10366 ( .A(n8125), .B(n8128), .Z(n8142) );
  NAND U10367 ( .A(n8143), .B(n8144), .Z(n8128) );
  NAND U10368 ( .A(n8145), .B(n8146), .Z(n8144) );
  OR U10369 ( .A(n8147), .B(n8148), .Z(n8145) );
  NANDN U10370 ( .A(n8149), .B(n8147), .Z(n8143) );
  IV U10371 ( .A(n8148), .Z(n8149) );
  NAND U10372 ( .A(n8150), .B(n8151), .Z(n8125) );
  NAND U10373 ( .A(n8152), .B(n8153), .Z(n8151) );
  NANDN U10374 ( .A(n8154), .B(n8155), .Z(n8152) );
  NANDN U10375 ( .A(n8155), .B(n8154), .Z(n8150) );
  AND U10376 ( .A(n8156), .B(n8157), .Z(n8127) );
  NAND U10377 ( .A(n8158), .B(n8159), .Z(n8157) );
  OR U10378 ( .A(n8160), .B(n8161), .Z(n8158) );
  NANDN U10379 ( .A(n8162), .B(n8160), .Z(n8156) );
  NAND U10380 ( .A(n8163), .B(n8164), .Z(n8131) );
  NANDN U10381 ( .A(n8165), .B(n8166), .Z(n8164) );
  OR U10382 ( .A(n8167), .B(n8168), .Z(n8166) );
  NANDN U10383 ( .A(n8169), .B(n8167), .Z(n8163) );
  IV U10384 ( .A(n8168), .Z(n8169) );
  XNOR U10385 ( .A(n8139), .B(n8170), .Z(n8134) );
  XNOR U10386 ( .A(n8137), .B(n8140), .Z(n8170) );
  NAND U10387 ( .A(n8171), .B(n8172), .Z(n8140) );
  NAND U10388 ( .A(n8173), .B(n8174), .Z(n8172) );
  OR U10389 ( .A(n8175), .B(n8176), .Z(n8173) );
  NANDN U10390 ( .A(n8177), .B(n8175), .Z(n8171) );
  IV U10391 ( .A(n8176), .Z(n8177) );
  NAND U10392 ( .A(n8178), .B(n8179), .Z(n8137) );
  NAND U10393 ( .A(n8180), .B(n8181), .Z(n8179) );
  NANDN U10394 ( .A(n8182), .B(n8183), .Z(n8180) );
  NANDN U10395 ( .A(n8183), .B(n8182), .Z(n8178) );
  AND U10396 ( .A(n8184), .B(n8185), .Z(n8139) );
  NAND U10397 ( .A(n8186), .B(n8187), .Z(n8185) );
  OR U10398 ( .A(n8188), .B(n8189), .Z(n8186) );
  NANDN U10399 ( .A(n8190), .B(n8188), .Z(n8184) );
  XNOR U10400 ( .A(n8165), .B(n8191), .Z(N13178) );
  XOR U10401 ( .A(n8167), .B(n8168), .Z(n8191) );
  XNOR U10402 ( .A(n8181), .B(n8192), .Z(n8168) );
  XOR U10403 ( .A(n8182), .B(n8183), .Z(n8192) );
  XOR U10404 ( .A(n8188), .B(n8193), .Z(n8183) );
  XOR U10405 ( .A(n8187), .B(n8190), .Z(n8193) );
  IV U10406 ( .A(n8189), .Z(n8190) );
  NAND U10407 ( .A(n8194), .B(n8195), .Z(n8189) );
  OR U10408 ( .A(n8196), .B(n8197), .Z(n8195) );
  OR U10409 ( .A(n8198), .B(n8199), .Z(n8194) );
  NAND U10410 ( .A(n8200), .B(n8201), .Z(n8187) );
  OR U10411 ( .A(n8202), .B(n8203), .Z(n8201) );
  OR U10412 ( .A(n8204), .B(n8205), .Z(n8200) );
  NOR U10413 ( .A(n8206), .B(n8207), .Z(n8188) );
  ANDN U10414 ( .B(n8208), .A(n8209), .Z(n8182) );
  XNOR U10415 ( .A(n8175), .B(n8210), .Z(n8181) );
  XNOR U10416 ( .A(n8174), .B(n8176), .Z(n8210) );
  NAND U10417 ( .A(n8211), .B(n8212), .Z(n8176) );
  OR U10418 ( .A(n8213), .B(n8214), .Z(n8212) );
  OR U10419 ( .A(n8215), .B(n8216), .Z(n8211) );
  NAND U10420 ( .A(n8217), .B(n8218), .Z(n8174) );
  OR U10421 ( .A(n8219), .B(n8220), .Z(n8218) );
  OR U10422 ( .A(n8221), .B(n8222), .Z(n8217) );
  ANDN U10423 ( .B(n8223), .A(n8224), .Z(n8175) );
  IV U10424 ( .A(n8225), .Z(n8223) );
  ANDN U10425 ( .B(n8226), .A(n8227), .Z(n8167) );
  XOR U10426 ( .A(n8153), .B(n8228), .Z(n8165) );
  XOR U10427 ( .A(n8154), .B(n8155), .Z(n8228) );
  XOR U10428 ( .A(n8160), .B(n8229), .Z(n8155) );
  XOR U10429 ( .A(n8159), .B(n8162), .Z(n8229) );
  IV U10430 ( .A(n8161), .Z(n8162) );
  NAND U10431 ( .A(n8230), .B(n8231), .Z(n8161) );
  OR U10432 ( .A(n8232), .B(n8233), .Z(n8231) );
  OR U10433 ( .A(n8234), .B(n8235), .Z(n8230) );
  NAND U10434 ( .A(n8236), .B(n8237), .Z(n8159) );
  OR U10435 ( .A(n8238), .B(n8239), .Z(n8237) );
  OR U10436 ( .A(n8240), .B(n8241), .Z(n8236) );
  NOR U10437 ( .A(n8242), .B(n8243), .Z(n8160) );
  ANDN U10438 ( .B(n8244), .A(n8245), .Z(n8154) );
  IV U10439 ( .A(n8246), .Z(n8244) );
  XNOR U10440 ( .A(n8147), .B(n8247), .Z(n8153) );
  XNOR U10441 ( .A(n8146), .B(n8148), .Z(n8247) );
  NAND U10442 ( .A(n8248), .B(n8249), .Z(n8148) );
  OR U10443 ( .A(n8250), .B(n8251), .Z(n8249) );
  OR U10444 ( .A(n8252), .B(n8253), .Z(n8248) );
  NAND U10445 ( .A(n8254), .B(n8255), .Z(n8146) );
  OR U10446 ( .A(n8256), .B(n8257), .Z(n8255) );
  OR U10447 ( .A(n8258), .B(n8259), .Z(n8254) );
  ANDN U10448 ( .B(n8260), .A(n8261), .Z(n8147) );
  IV U10449 ( .A(n8262), .Z(n8260) );
  XNOR U10450 ( .A(n8227), .B(n8226), .Z(N13177) );
  XOR U10451 ( .A(n8246), .B(n8245), .Z(n8226) );
  XNOR U10452 ( .A(n8261), .B(n8262), .Z(n8245) );
  XNOR U10453 ( .A(n8256), .B(n8257), .Z(n8262) );
  XNOR U10454 ( .A(n8258), .B(n8259), .Z(n8257) );
  XNOR U10455 ( .A(y[877]), .B(x[877]), .Z(n8259) );
  XNOR U10456 ( .A(y[878]), .B(x[878]), .Z(n8258) );
  XNOR U10457 ( .A(y[876]), .B(x[876]), .Z(n8256) );
  XNOR U10458 ( .A(n8250), .B(n8251), .Z(n8261) );
  XNOR U10459 ( .A(y[873]), .B(x[873]), .Z(n8251) );
  XNOR U10460 ( .A(n8252), .B(n8253), .Z(n8250) );
  XNOR U10461 ( .A(y[874]), .B(x[874]), .Z(n8253) );
  XNOR U10462 ( .A(y[875]), .B(x[875]), .Z(n8252) );
  XNOR U10463 ( .A(n8243), .B(n8242), .Z(n8246) );
  XNOR U10464 ( .A(n8238), .B(n8239), .Z(n8242) );
  XNOR U10465 ( .A(y[870]), .B(x[870]), .Z(n8239) );
  XNOR U10466 ( .A(n8240), .B(n8241), .Z(n8238) );
  XNOR U10467 ( .A(y[871]), .B(x[871]), .Z(n8241) );
  XNOR U10468 ( .A(y[872]), .B(x[872]), .Z(n8240) );
  XNOR U10469 ( .A(n8232), .B(n8233), .Z(n8243) );
  XNOR U10470 ( .A(y[867]), .B(x[867]), .Z(n8233) );
  XNOR U10471 ( .A(n8234), .B(n8235), .Z(n8232) );
  XNOR U10472 ( .A(y[868]), .B(x[868]), .Z(n8235) );
  XNOR U10473 ( .A(y[869]), .B(x[869]), .Z(n8234) );
  XOR U10474 ( .A(n8208), .B(n8209), .Z(n8227) );
  XNOR U10475 ( .A(n8224), .B(n8225), .Z(n8209) );
  XNOR U10476 ( .A(n8219), .B(n8220), .Z(n8225) );
  XNOR U10477 ( .A(n8221), .B(n8222), .Z(n8220) );
  XNOR U10478 ( .A(y[865]), .B(x[865]), .Z(n8222) );
  XNOR U10479 ( .A(y[866]), .B(x[866]), .Z(n8221) );
  XNOR U10480 ( .A(y[864]), .B(x[864]), .Z(n8219) );
  XNOR U10481 ( .A(n8213), .B(n8214), .Z(n8224) );
  XNOR U10482 ( .A(y[861]), .B(x[861]), .Z(n8214) );
  XNOR U10483 ( .A(n8215), .B(n8216), .Z(n8213) );
  XNOR U10484 ( .A(y[862]), .B(x[862]), .Z(n8216) );
  XNOR U10485 ( .A(y[863]), .B(x[863]), .Z(n8215) );
  XOR U10486 ( .A(n8207), .B(n8206), .Z(n8208) );
  XNOR U10487 ( .A(n8202), .B(n8203), .Z(n8206) );
  XNOR U10488 ( .A(y[858]), .B(x[858]), .Z(n8203) );
  XNOR U10489 ( .A(n8204), .B(n8205), .Z(n8202) );
  XNOR U10490 ( .A(y[859]), .B(x[859]), .Z(n8205) );
  XNOR U10491 ( .A(y[860]), .B(x[860]), .Z(n8204) );
  XNOR U10492 ( .A(n8196), .B(n8197), .Z(n8207) );
  XNOR U10493 ( .A(y[855]), .B(x[855]), .Z(n8197) );
  XNOR U10494 ( .A(n8198), .B(n8199), .Z(n8196) );
  XNOR U10495 ( .A(y[856]), .B(x[856]), .Z(n8199) );
  XNOR U10496 ( .A(y[857]), .B(x[857]), .Z(n8198) );
  NAND U10497 ( .A(n8263), .B(n8264), .Z(N13170) );
  NANDN U10498 ( .A(n8265), .B(n8266), .Z(n8264) );
  OR U10499 ( .A(n8267), .B(n8268), .Z(n8266) );
  NAND U10500 ( .A(n8267), .B(n8268), .Z(n8263) );
  XOR U10501 ( .A(n8267), .B(n8269), .Z(N13169) );
  XNOR U10502 ( .A(n8265), .B(n8268), .Z(n8269) );
  AND U10503 ( .A(n8270), .B(n8271), .Z(n8268) );
  NANDN U10504 ( .A(n8272), .B(n8273), .Z(n8271) );
  NANDN U10505 ( .A(n8274), .B(n8275), .Z(n8273) );
  NANDN U10506 ( .A(n8275), .B(n8274), .Z(n8270) );
  NAND U10507 ( .A(n8276), .B(n8277), .Z(n8265) );
  NANDN U10508 ( .A(n8278), .B(n8279), .Z(n8277) );
  OR U10509 ( .A(n8280), .B(n8281), .Z(n8279) );
  NAND U10510 ( .A(n8281), .B(n8280), .Z(n8276) );
  AND U10511 ( .A(n8282), .B(n8283), .Z(n8267) );
  NANDN U10512 ( .A(n8284), .B(n8285), .Z(n8283) );
  NANDN U10513 ( .A(n8286), .B(n8287), .Z(n8285) );
  NANDN U10514 ( .A(n8287), .B(n8286), .Z(n8282) );
  XOR U10515 ( .A(n8281), .B(n8288), .Z(N13168) );
  XOR U10516 ( .A(n8278), .B(n8280), .Z(n8288) );
  XNOR U10517 ( .A(n8274), .B(n8289), .Z(n8280) );
  XNOR U10518 ( .A(n8272), .B(n8275), .Z(n8289) );
  NAND U10519 ( .A(n8290), .B(n8291), .Z(n8275) );
  NAND U10520 ( .A(n8292), .B(n8293), .Z(n8291) );
  OR U10521 ( .A(n8294), .B(n8295), .Z(n8292) );
  NANDN U10522 ( .A(n8296), .B(n8294), .Z(n8290) );
  IV U10523 ( .A(n8295), .Z(n8296) );
  NAND U10524 ( .A(n8297), .B(n8298), .Z(n8272) );
  NAND U10525 ( .A(n8299), .B(n8300), .Z(n8298) );
  NANDN U10526 ( .A(n8301), .B(n8302), .Z(n8299) );
  NANDN U10527 ( .A(n8302), .B(n8301), .Z(n8297) );
  AND U10528 ( .A(n8303), .B(n8304), .Z(n8274) );
  NAND U10529 ( .A(n8305), .B(n8306), .Z(n8304) );
  OR U10530 ( .A(n8307), .B(n8308), .Z(n8305) );
  NANDN U10531 ( .A(n8309), .B(n8307), .Z(n8303) );
  NAND U10532 ( .A(n8310), .B(n8311), .Z(n8278) );
  NANDN U10533 ( .A(n8312), .B(n8313), .Z(n8311) );
  OR U10534 ( .A(n8314), .B(n8315), .Z(n8313) );
  NANDN U10535 ( .A(n8316), .B(n8314), .Z(n8310) );
  IV U10536 ( .A(n8315), .Z(n8316) );
  XNOR U10537 ( .A(n8286), .B(n8317), .Z(n8281) );
  XNOR U10538 ( .A(n8284), .B(n8287), .Z(n8317) );
  NAND U10539 ( .A(n8318), .B(n8319), .Z(n8287) );
  NAND U10540 ( .A(n8320), .B(n8321), .Z(n8319) );
  OR U10541 ( .A(n8322), .B(n8323), .Z(n8320) );
  NANDN U10542 ( .A(n8324), .B(n8322), .Z(n8318) );
  IV U10543 ( .A(n8323), .Z(n8324) );
  NAND U10544 ( .A(n8325), .B(n8326), .Z(n8284) );
  NAND U10545 ( .A(n8327), .B(n8328), .Z(n8326) );
  NANDN U10546 ( .A(n8329), .B(n8330), .Z(n8327) );
  NANDN U10547 ( .A(n8330), .B(n8329), .Z(n8325) );
  AND U10548 ( .A(n8331), .B(n8332), .Z(n8286) );
  NAND U10549 ( .A(n8333), .B(n8334), .Z(n8332) );
  OR U10550 ( .A(n8335), .B(n8336), .Z(n8333) );
  NANDN U10551 ( .A(n8337), .B(n8335), .Z(n8331) );
  XNOR U10552 ( .A(n8312), .B(n8338), .Z(N13167) );
  XOR U10553 ( .A(n8314), .B(n8315), .Z(n8338) );
  XNOR U10554 ( .A(n8328), .B(n8339), .Z(n8315) );
  XOR U10555 ( .A(n8329), .B(n8330), .Z(n8339) );
  XOR U10556 ( .A(n8335), .B(n8340), .Z(n8330) );
  XOR U10557 ( .A(n8334), .B(n8337), .Z(n8340) );
  IV U10558 ( .A(n8336), .Z(n8337) );
  NAND U10559 ( .A(n8341), .B(n8342), .Z(n8336) );
  OR U10560 ( .A(n8343), .B(n8344), .Z(n8342) );
  OR U10561 ( .A(n8345), .B(n8346), .Z(n8341) );
  NAND U10562 ( .A(n8347), .B(n8348), .Z(n8334) );
  OR U10563 ( .A(n8349), .B(n8350), .Z(n8348) );
  OR U10564 ( .A(n8351), .B(n8352), .Z(n8347) );
  NOR U10565 ( .A(n8353), .B(n8354), .Z(n8335) );
  ANDN U10566 ( .B(n8355), .A(n8356), .Z(n8329) );
  XNOR U10567 ( .A(n8322), .B(n8357), .Z(n8328) );
  XNOR U10568 ( .A(n8321), .B(n8323), .Z(n8357) );
  NAND U10569 ( .A(n8358), .B(n8359), .Z(n8323) );
  OR U10570 ( .A(n8360), .B(n8361), .Z(n8359) );
  OR U10571 ( .A(n8362), .B(n8363), .Z(n8358) );
  NAND U10572 ( .A(n8364), .B(n8365), .Z(n8321) );
  OR U10573 ( .A(n8366), .B(n8367), .Z(n8365) );
  OR U10574 ( .A(n8368), .B(n8369), .Z(n8364) );
  ANDN U10575 ( .B(n8370), .A(n8371), .Z(n8322) );
  IV U10576 ( .A(n8372), .Z(n8370) );
  ANDN U10577 ( .B(n8373), .A(n8374), .Z(n8314) );
  XOR U10578 ( .A(n8300), .B(n8375), .Z(n8312) );
  XOR U10579 ( .A(n8301), .B(n8302), .Z(n8375) );
  XOR U10580 ( .A(n8307), .B(n8376), .Z(n8302) );
  XOR U10581 ( .A(n8306), .B(n8309), .Z(n8376) );
  IV U10582 ( .A(n8308), .Z(n8309) );
  NAND U10583 ( .A(n8377), .B(n8378), .Z(n8308) );
  OR U10584 ( .A(n8379), .B(n8380), .Z(n8378) );
  OR U10585 ( .A(n8381), .B(n8382), .Z(n8377) );
  NAND U10586 ( .A(n8383), .B(n8384), .Z(n8306) );
  OR U10587 ( .A(n8385), .B(n8386), .Z(n8384) );
  OR U10588 ( .A(n8387), .B(n8388), .Z(n8383) );
  NOR U10589 ( .A(n8389), .B(n8390), .Z(n8307) );
  ANDN U10590 ( .B(n8391), .A(n8392), .Z(n8301) );
  IV U10591 ( .A(n8393), .Z(n8391) );
  XNOR U10592 ( .A(n8294), .B(n8394), .Z(n8300) );
  XNOR U10593 ( .A(n8293), .B(n8295), .Z(n8394) );
  NAND U10594 ( .A(n8395), .B(n8396), .Z(n8295) );
  OR U10595 ( .A(n8397), .B(n8398), .Z(n8396) );
  OR U10596 ( .A(n8399), .B(n8400), .Z(n8395) );
  NAND U10597 ( .A(n8401), .B(n8402), .Z(n8293) );
  OR U10598 ( .A(n8403), .B(n8404), .Z(n8402) );
  OR U10599 ( .A(n8405), .B(n8406), .Z(n8401) );
  ANDN U10600 ( .B(n8407), .A(n8408), .Z(n8294) );
  IV U10601 ( .A(n8409), .Z(n8407) );
  XNOR U10602 ( .A(n8374), .B(n8373), .Z(N13166) );
  XOR U10603 ( .A(n8393), .B(n8392), .Z(n8373) );
  XNOR U10604 ( .A(n8408), .B(n8409), .Z(n8392) );
  XNOR U10605 ( .A(n8403), .B(n8404), .Z(n8409) );
  XNOR U10606 ( .A(n8405), .B(n8406), .Z(n8404) );
  XNOR U10607 ( .A(y[853]), .B(x[853]), .Z(n8406) );
  XNOR U10608 ( .A(y[854]), .B(x[854]), .Z(n8405) );
  XNOR U10609 ( .A(y[852]), .B(x[852]), .Z(n8403) );
  XNOR U10610 ( .A(n8397), .B(n8398), .Z(n8408) );
  XNOR U10611 ( .A(y[849]), .B(x[849]), .Z(n8398) );
  XNOR U10612 ( .A(n8399), .B(n8400), .Z(n8397) );
  XNOR U10613 ( .A(y[850]), .B(x[850]), .Z(n8400) );
  XNOR U10614 ( .A(y[851]), .B(x[851]), .Z(n8399) );
  XNOR U10615 ( .A(n8390), .B(n8389), .Z(n8393) );
  XNOR U10616 ( .A(n8385), .B(n8386), .Z(n8389) );
  XNOR U10617 ( .A(y[846]), .B(x[846]), .Z(n8386) );
  XNOR U10618 ( .A(n8387), .B(n8388), .Z(n8385) );
  XNOR U10619 ( .A(y[847]), .B(x[847]), .Z(n8388) );
  XNOR U10620 ( .A(y[848]), .B(x[848]), .Z(n8387) );
  XNOR U10621 ( .A(n8379), .B(n8380), .Z(n8390) );
  XNOR U10622 ( .A(y[843]), .B(x[843]), .Z(n8380) );
  XNOR U10623 ( .A(n8381), .B(n8382), .Z(n8379) );
  XNOR U10624 ( .A(y[844]), .B(x[844]), .Z(n8382) );
  XNOR U10625 ( .A(y[845]), .B(x[845]), .Z(n8381) );
  XOR U10626 ( .A(n8355), .B(n8356), .Z(n8374) );
  XNOR U10627 ( .A(n8371), .B(n8372), .Z(n8356) );
  XNOR U10628 ( .A(n8366), .B(n8367), .Z(n8372) );
  XNOR U10629 ( .A(n8368), .B(n8369), .Z(n8367) );
  XNOR U10630 ( .A(y[841]), .B(x[841]), .Z(n8369) );
  XNOR U10631 ( .A(y[842]), .B(x[842]), .Z(n8368) );
  XNOR U10632 ( .A(y[840]), .B(x[840]), .Z(n8366) );
  XNOR U10633 ( .A(n8360), .B(n8361), .Z(n8371) );
  XNOR U10634 ( .A(y[837]), .B(x[837]), .Z(n8361) );
  XNOR U10635 ( .A(n8362), .B(n8363), .Z(n8360) );
  XNOR U10636 ( .A(y[838]), .B(x[838]), .Z(n8363) );
  XNOR U10637 ( .A(y[839]), .B(x[839]), .Z(n8362) );
  XOR U10638 ( .A(n8354), .B(n8353), .Z(n8355) );
  XNOR U10639 ( .A(n8349), .B(n8350), .Z(n8353) );
  XNOR U10640 ( .A(y[834]), .B(x[834]), .Z(n8350) );
  XNOR U10641 ( .A(n8351), .B(n8352), .Z(n8349) );
  XNOR U10642 ( .A(y[835]), .B(x[835]), .Z(n8352) );
  XNOR U10643 ( .A(y[836]), .B(x[836]), .Z(n8351) );
  XNOR U10644 ( .A(n8343), .B(n8344), .Z(n8354) );
  XNOR U10645 ( .A(y[831]), .B(x[831]), .Z(n8344) );
  XNOR U10646 ( .A(n8345), .B(n8346), .Z(n8343) );
  XNOR U10647 ( .A(y[832]), .B(x[832]), .Z(n8346) );
  XNOR U10648 ( .A(y[833]), .B(x[833]), .Z(n8345) );
  NAND U10649 ( .A(n8410), .B(n8411), .Z(N13159) );
  NANDN U10650 ( .A(n8412), .B(n8413), .Z(n8411) );
  OR U10651 ( .A(n8414), .B(n8415), .Z(n8413) );
  NAND U10652 ( .A(n8414), .B(n8415), .Z(n8410) );
  XOR U10653 ( .A(n8414), .B(n8416), .Z(N13158) );
  XNOR U10654 ( .A(n8412), .B(n8415), .Z(n8416) );
  AND U10655 ( .A(n8417), .B(n8418), .Z(n8415) );
  NANDN U10656 ( .A(n8419), .B(n8420), .Z(n8418) );
  NANDN U10657 ( .A(n8421), .B(n8422), .Z(n8420) );
  NANDN U10658 ( .A(n8422), .B(n8421), .Z(n8417) );
  NAND U10659 ( .A(n8423), .B(n8424), .Z(n8412) );
  NANDN U10660 ( .A(n8425), .B(n8426), .Z(n8424) );
  OR U10661 ( .A(n8427), .B(n8428), .Z(n8426) );
  NAND U10662 ( .A(n8428), .B(n8427), .Z(n8423) );
  AND U10663 ( .A(n8429), .B(n8430), .Z(n8414) );
  NANDN U10664 ( .A(n8431), .B(n8432), .Z(n8430) );
  NANDN U10665 ( .A(n8433), .B(n8434), .Z(n8432) );
  NANDN U10666 ( .A(n8434), .B(n8433), .Z(n8429) );
  XOR U10667 ( .A(n8428), .B(n8435), .Z(N13157) );
  XOR U10668 ( .A(n8425), .B(n8427), .Z(n8435) );
  XNOR U10669 ( .A(n8421), .B(n8436), .Z(n8427) );
  XNOR U10670 ( .A(n8419), .B(n8422), .Z(n8436) );
  NAND U10671 ( .A(n8437), .B(n8438), .Z(n8422) );
  NAND U10672 ( .A(n8439), .B(n8440), .Z(n8438) );
  OR U10673 ( .A(n8441), .B(n8442), .Z(n8439) );
  NANDN U10674 ( .A(n8443), .B(n8441), .Z(n8437) );
  IV U10675 ( .A(n8442), .Z(n8443) );
  NAND U10676 ( .A(n8444), .B(n8445), .Z(n8419) );
  NAND U10677 ( .A(n8446), .B(n8447), .Z(n8445) );
  NANDN U10678 ( .A(n8448), .B(n8449), .Z(n8446) );
  NANDN U10679 ( .A(n8449), .B(n8448), .Z(n8444) );
  AND U10680 ( .A(n8450), .B(n8451), .Z(n8421) );
  NAND U10681 ( .A(n8452), .B(n8453), .Z(n8451) );
  OR U10682 ( .A(n8454), .B(n8455), .Z(n8452) );
  NANDN U10683 ( .A(n8456), .B(n8454), .Z(n8450) );
  NAND U10684 ( .A(n8457), .B(n8458), .Z(n8425) );
  NANDN U10685 ( .A(n8459), .B(n8460), .Z(n8458) );
  OR U10686 ( .A(n8461), .B(n8462), .Z(n8460) );
  NANDN U10687 ( .A(n8463), .B(n8461), .Z(n8457) );
  IV U10688 ( .A(n8462), .Z(n8463) );
  XNOR U10689 ( .A(n8433), .B(n8464), .Z(n8428) );
  XNOR U10690 ( .A(n8431), .B(n8434), .Z(n8464) );
  NAND U10691 ( .A(n8465), .B(n8466), .Z(n8434) );
  NAND U10692 ( .A(n8467), .B(n8468), .Z(n8466) );
  OR U10693 ( .A(n8469), .B(n8470), .Z(n8467) );
  NANDN U10694 ( .A(n8471), .B(n8469), .Z(n8465) );
  IV U10695 ( .A(n8470), .Z(n8471) );
  NAND U10696 ( .A(n8472), .B(n8473), .Z(n8431) );
  NAND U10697 ( .A(n8474), .B(n8475), .Z(n8473) );
  NANDN U10698 ( .A(n8476), .B(n8477), .Z(n8474) );
  NANDN U10699 ( .A(n8477), .B(n8476), .Z(n8472) );
  AND U10700 ( .A(n8478), .B(n8479), .Z(n8433) );
  NAND U10701 ( .A(n8480), .B(n8481), .Z(n8479) );
  OR U10702 ( .A(n8482), .B(n8483), .Z(n8480) );
  NANDN U10703 ( .A(n8484), .B(n8482), .Z(n8478) );
  XNOR U10704 ( .A(n8459), .B(n8485), .Z(N13156) );
  XOR U10705 ( .A(n8461), .B(n8462), .Z(n8485) );
  XNOR U10706 ( .A(n8475), .B(n8486), .Z(n8462) );
  XOR U10707 ( .A(n8476), .B(n8477), .Z(n8486) );
  XOR U10708 ( .A(n8482), .B(n8487), .Z(n8477) );
  XOR U10709 ( .A(n8481), .B(n8484), .Z(n8487) );
  IV U10710 ( .A(n8483), .Z(n8484) );
  NAND U10711 ( .A(n8488), .B(n8489), .Z(n8483) );
  OR U10712 ( .A(n8490), .B(n8491), .Z(n8489) );
  OR U10713 ( .A(n8492), .B(n8493), .Z(n8488) );
  NAND U10714 ( .A(n8494), .B(n8495), .Z(n8481) );
  OR U10715 ( .A(n8496), .B(n8497), .Z(n8495) );
  OR U10716 ( .A(n8498), .B(n8499), .Z(n8494) );
  NOR U10717 ( .A(n8500), .B(n8501), .Z(n8482) );
  ANDN U10718 ( .B(n8502), .A(n8503), .Z(n8476) );
  XNOR U10719 ( .A(n8469), .B(n8504), .Z(n8475) );
  XNOR U10720 ( .A(n8468), .B(n8470), .Z(n8504) );
  NAND U10721 ( .A(n8505), .B(n8506), .Z(n8470) );
  OR U10722 ( .A(n8507), .B(n8508), .Z(n8506) );
  OR U10723 ( .A(n8509), .B(n8510), .Z(n8505) );
  NAND U10724 ( .A(n8511), .B(n8512), .Z(n8468) );
  OR U10725 ( .A(n8513), .B(n8514), .Z(n8512) );
  OR U10726 ( .A(n8515), .B(n8516), .Z(n8511) );
  ANDN U10727 ( .B(n8517), .A(n8518), .Z(n8469) );
  IV U10728 ( .A(n8519), .Z(n8517) );
  ANDN U10729 ( .B(n8520), .A(n8521), .Z(n8461) );
  XOR U10730 ( .A(n8447), .B(n8522), .Z(n8459) );
  XOR U10731 ( .A(n8448), .B(n8449), .Z(n8522) );
  XOR U10732 ( .A(n8454), .B(n8523), .Z(n8449) );
  XOR U10733 ( .A(n8453), .B(n8456), .Z(n8523) );
  IV U10734 ( .A(n8455), .Z(n8456) );
  NAND U10735 ( .A(n8524), .B(n8525), .Z(n8455) );
  OR U10736 ( .A(n8526), .B(n8527), .Z(n8525) );
  OR U10737 ( .A(n8528), .B(n8529), .Z(n8524) );
  NAND U10738 ( .A(n8530), .B(n8531), .Z(n8453) );
  OR U10739 ( .A(n8532), .B(n8533), .Z(n8531) );
  OR U10740 ( .A(n8534), .B(n8535), .Z(n8530) );
  NOR U10741 ( .A(n8536), .B(n8537), .Z(n8454) );
  ANDN U10742 ( .B(n8538), .A(n8539), .Z(n8448) );
  IV U10743 ( .A(n8540), .Z(n8538) );
  XNOR U10744 ( .A(n8441), .B(n8541), .Z(n8447) );
  XNOR U10745 ( .A(n8440), .B(n8442), .Z(n8541) );
  NAND U10746 ( .A(n8542), .B(n8543), .Z(n8442) );
  OR U10747 ( .A(n8544), .B(n8545), .Z(n8543) );
  OR U10748 ( .A(n8546), .B(n8547), .Z(n8542) );
  NAND U10749 ( .A(n8548), .B(n8549), .Z(n8440) );
  OR U10750 ( .A(n8550), .B(n8551), .Z(n8549) );
  OR U10751 ( .A(n8552), .B(n8553), .Z(n8548) );
  ANDN U10752 ( .B(n8554), .A(n8555), .Z(n8441) );
  IV U10753 ( .A(n8556), .Z(n8554) );
  XNOR U10754 ( .A(n8521), .B(n8520), .Z(N13155) );
  XOR U10755 ( .A(n8540), .B(n8539), .Z(n8520) );
  XNOR U10756 ( .A(n8555), .B(n8556), .Z(n8539) );
  XNOR U10757 ( .A(n8550), .B(n8551), .Z(n8556) );
  XNOR U10758 ( .A(n8552), .B(n8553), .Z(n8551) );
  XNOR U10759 ( .A(y[829]), .B(x[829]), .Z(n8553) );
  XNOR U10760 ( .A(y[830]), .B(x[830]), .Z(n8552) );
  XNOR U10761 ( .A(y[828]), .B(x[828]), .Z(n8550) );
  XNOR U10762 ( .A(n8544), .B(n8545), .Z(n8555) );
  XNOR U10763 ( .A(y[825]), .B(x[825]), .Z(n8545) );
  XNOR U10764 ( .A(n8546), .B(n8547), .Z(n8544) );
  XNOR U10765 ( .A(y[826]), .B(x[826]), .Z(n8547) );
  XNOR U10766 ( .A(y[827]), .B(x[827]), .Z(n8546) );
  XNOR U10767 ( .A(n8537), .B(n8536), .Z(n8540) );
  XNOR U10768 ( .A(n8532), .B(n8533), .Z(n8536) );
  XNOR U10769 ( .A(y[822]), .B(x[822]), .Z(n8533) );
  XNOR U10770 ( .A(n8534), .B(n8535), .Z(n8532) );
  XNOR U10771 ( .A(y[823]), .B(x[823]), .Z(n8535) );
  XNOR U10772 ( .A(y[824]), .B(x[824]), .Z(n8534) );
  XNOR U10773 ( .A(n8526), .B(n8527), .Z(n8537) );
  XNOR U10774 ( .A(y[819]), .B(x[819]), .Z(n8527) );
  XNOR U10775 ( .A(n8528), .B(n8529), .Z(n8526) );
  XNOR U10776 ( .A(y[820]), .B(x[820]), .Z(n8529) );
  XNOR U10777 ( .A(y[821]), .B(x[821]), .Z(n8528) );
  XOR U10778 ( .A(n8502), .B(n8503), .Z(n8521) );
  XNOR U10779 ( .A(n8518), .B(n8519), .Z(n8503) );
  XNOR U10780 ( .A(n8513), .B(n8514), .Z(n8519) );
  XNOR U10781 ( .A(n8515), .B(n8516), .Z(n8514) );
  XNOR U10782 ( .A(y[817]), .B(x[817]), .Z(n8516) );
  XNOR U10783 ( .A(y[818]), .B(x[818]), .Z(n8515) );
  XNOR U10784 ( .A(y[816]), .B(x[816]), .Z(n8513) );
  XNOR U10785 ( .A(n8507), .B(n8508), .Z(n8518) );
  XNOR U10786 ( .A(y[813]), .B(x[813]), .Z(n8508) );
  XNOR U10787 ( .A(n8509), .B(n8510), .Z(n8507) );
  XNOR U10788 ( .A(y[814]), .B(x[814]), .Z(n8510) );
  XNOR U10789 ( .A(y[815]), .B(x[815]), .Z(n8509) );
  XOR U10790 ( .A(n8501), .B(n8500), .Z(n8502) );
  XNOR U10791 ( .A(n8496), .B(n8497), .Z(n8500) );
  XNOR U10792 ( .A(y[810]), .B(x[810]), .Z(n8497) );
  XNOR U10793 ( .A(n8498), .B(n8499), .Z(n8496) );
  XNOR U10794 ( .A(y[811]), .B(x[811]), .Z(n8499) );
  XNOR U10795 ( .A(y[812]), .B(x[812]), .Z(n8498) );
  XNOR U10796 ( .A(n8490), .B(n8491), .Z(n8501) );
  XNOR U10797 ( .A(y[807]), .B(x[807]), .Z(n8491) );
  XNOR U10798 ( .A(n8492), .B(n8493), .Z(n8490) );
  XNOR U10799 ( .A(y[808]), .B(x[808]), .Z(n8493) );
  XNOR U10800 ( .A(y[809]), .B(x[809]), .Z(n8492) );
  NAND U10801 ( .A(n8557), .B(n8558), .Z(N13148) );
  NANDN U10802 ( .A(n8559), .B(n8560), .Z(n8558) );
  OR U10803 ( .A(n8561), .B(n8562), .Z(n8560) );
  NAND U10804 ( .A(n8561), .B(n8562), .Z(n8557) );
  XOR U10805 ( .A(n8561), .B(n8563), .Z(N13147) );
  XNOR U10806 ( .A(n8559), .B(n8562), .Z(n8563) );
  AND U10807 ( .A(n8564), .B(n8565), .Z(n8562) );
  NANDN U10808 ( .A(n8566), .B(n8567), .Z(n8565) );
  NANDN U10809 ( .A(n8568), .B(n8569), .Z(n8567) );
  NANDN U10810 ( .A(n8569), .B(n8568), .Z(n8564) );
  NAND U10811 ( .A(n8570), .B(n8571), .Z(n8559) );
  NANDN U10812 ( .A(n8572), .B(n8573), .Z(n8571) );
  OR U10813 ( .A(n8574), .B(n8575), .Z(n8573) );
  NAND U10814 ( .A(n8575), .B(n8574), .Z(n8570) );
  AND U10815 ( .A(n8576), .B(n8577), .Z(n8561) );
  NANDN U10816 ( .A(n8578), .B(n8579), .Z(n8577) );
  NANDN U10817 ( .A(n8580), .B(n8581), .Z(n8579) );
  NANDN U10818 ( .A(n8581), .B(n8580), .Z(n8576) );
  XOR U10819 ( .A(n8575), .B(n8582), .Z(N13146) );
  XOR U10820 ( .A(n8572), .B(n8574), .Z(n8582) );
  XNOR U10821 ( .A(n8568), .B(n8583), .Z(n8574) );
  XNOR U10822 ( .A(n8566), .B(n8569), .Z(n8583) );
  NAND U10823 ( .A(n8584), .B(n8585), .Z(n8569) );
  NAND U10824 ( .A(n8586), .B(n8587), .Z(n8585) );
  OR U10825 ( .A(n8588), .B(n8589), .Z(n8586) );
  NANDN U10826 ( .A(n8590), .B(n8588), .Z(n8584) );
  IV U10827 ( .A(n8589), .Z(n8590) );
  NAND U10828 ( .A(n8591), .B(n8592), .Z(n8566) );
  NAND U10829 ( .A(n8593), .B(n8594), .Z(n8592) );
  NANDN U10830 ( .A(n8595), .B(n8596), .Z(n8593) );
  NANDN U10831 ( .A(n8596), .B(n8595), .Z(n8591) );
  AND U10832 ( .A(n8597), .B(n8598), .Z(n8568) );
  NAND U10833 ( .A(n8599), .B(n8600), .Z(n8598) );
  OR U10834 ( .A(n8601), .B(n8602), .Z(n8599) );
  NANDN U10835 ( .A(n8603), .B(n8601), .Z(n8597) );
  NAND U10836 ( .A(n8604), .B(n8605), .Z(n8572) );
  NANDN U10837 ( .A(n8606), .B(n8607), .Z(n8605) );
  OR U10838 ( .A(n8608), .B(n8609), .Z(n8607) );
  NANDN U10839 ( .A(n8610), .B(n8608), .Z(n8604) );
  IV U10840 ( .A(n8609), .Z(n8610) );
  XNOR U10841 ( .A(n8580), .B(n8611), .Z(n8575) );
  XNOR U10842 ( .A(n8578), .B(n8581), .Z(n8611) );
  NAND U10843 ( .A(n8612), .B(n8613), .Z(n8581) );
  NAND U10844 ( .A(n8614), .B(n8615), .Z(n8613) );
  OR U10845 ( .A(n8616), .B(n8617), .Z(n8614) );
  NANDN U10846 ( .A(n8618), .B(n8616), .Z(n8612) );
  IV U10847 ( .A(n8617), .Z(n8618) );
  NAND U10848 ( .A(n8619), .B(n8620), .Z(n8578) );
  NAND U10849 ( .A(n8621), .B(n8622), .Z(n8620) );
  NANDN U10850 ( .A(n8623), .B(n8624), .Z(n8621) );
  NANDN U10851 ( .A(n8624), .B(n8623), .Z(n8619) );
  AND U10852 ( .A(n8625), .B(n8626), .Z(n8580) );
  NAND U10853 ( .A(n8627), .B(n8628), .Z(n8626) );
  OR U10854 ( .A(n8629), .B(n8630), .Z(n8627) );
  NANDN U10855 ( .A(n8631), .B(n8629), .Z(n8625) );
  XNOR U10856 ( .A(n8606), .B(n8632), .Z(N13145) );
  XOR U10857 ( .A(n8608), .B(n8609), .Z(n8632) );
  XNOR U10858 ( .A(n8622), .B(n8633), .Z(n8609) );
  XOR U10859 ( .A(n8623), .B(n8624), .Z(n8633) );
  XOR U10860 ( .A(n8629), .B(n8634), .Z(n8624) );
  XOR U10861 ( .A(n8628), .B(n8631), .Z(n8634) );
  IV U10862 ( .A(n8630), .Z(n8631) );
  NAND U10863 ( .A(n8635), .B(n8636), .Z(n8630) );
  OR U10864 ( .A(n8637), .B(n8638), .Z(n8636) );
  OR U10865 ( .A(n8639), .B(n8640), .Z(n8635) );
  NAND U10866 ( .A(n8641), .B(n8642), .Z(n8628) );
  OR U10867 ( .A(n8643), .B(n8644), .Z(n8642) );
  OR U10868 ( .A(n8645), .B(n8646), .Z(n8641) );
  NOR U10869 ( .A(n8647), .B(n8648), .Z(n8629) );
  ANDN U10870 ( .B(n8649), .A(n8650), .Z(n8623) );
  XNOR U10871 ( .A(n8616), .B(n8651), .Z(n8622) );
  XNOR U10872 ( .A(n8615), .B(n8617), .Z(n8651) );
  NAND U10873 ( .A(n8652), .B(n8653), .Z(n8617) );
  OR U10874 ( .A(n8654), .B(n8655), .Z(n8653) );
  OR U10875 ( .A(n8656), .B(n8657), .Z(n8652) );
  NAND U10876 ( .A(n8658), .B(n8659), .Z(n8615) );
  OR U10877 ( .A(n8660), .B(n8661), .Z(n8659) );
  OR U10878 ( .A(n8662), .B(n8663), .Z(n8658) );
  ANDN U10879 ( .B(n8664), .A(n8665), .Z(n8616) );
  IV U10880 ( .A(n8666), .Z(n8664) );
  ANDN U10881 ( .B(n8667), .A(n8668), .Z(n8608) );
  XOR U10882 ( .A(n8594), .B(n8669), .Z(n8606) );
  XOR U10883 ( .A(n8595), .B(n8596), .Z(n8669) );
  XOR U10884 ( .A(n8601), .B(n8670), .Z(n8596) );
  XOR U10885 ( .A(n8600), .B(n8603), .Z(n8670) );
  IV U10886 ( .A(n8602), .Z(n8603) );
  NAND U10887 ( .A(n8671), .B(n8672), .Z(n8602) );
  OR U10888 ( .A(n8673), .B(n8674), .Z(n8672) );
  OR U10889 ( .A(n8675), .B(n8676), .Z(n8671) );
  NAND U10890 ( .A(n8677), .B(n8678), .Z(n8600) );
  OR U10891 ( .A(n8679), .B(n8680), .Z(n8678) );
  OR U10892 ( .A(n8681), .B(n8682), .Z(n8677) );
  NOR U10893 ( .A(n8683), .B(n8684), .Z(n8601) );
  ANDN U10894 ( .B(n8685), .A(n8686), .Z(n8595) );
  IV U10895 ( .A(n8687), .Z(n8685) );
  XNOR U10896 ( .A(n8588), .B(n8688), .Z(n8594) );
  XNOR U10897 ( .A(n8587), .B(n8589), .Z(n8688) );
  NAND U10898 ( .A(n8689), .B(n8690), .Z(n8589) );
  OR U10899 ( .A(n8691), .B(n8692), .Z(n8690) );
  OR U10900 ( .A(n8693), .B(n8694), .Z(n8689) );
  NAND U10901 ( .A(n8695), .B(n8696), .Z(n8587) );
  OR U10902 ( .A(n8697), .B(n8698), .Z(n8696) );
  OR U10903 ( .A(n8699), .B(n8700), .Z(n8695) );
  ANDN U10904 ( .B(n8701), .A(n8702), .Z(n8588) );
  IV U10905 ( .A(n8703), .Z(n8701) );
  XNOR U10906 ( .A(n8668), .B(n8667), .Z(N13144) );
  XOR U10907 ( .A(n8687), .B(n8686), .Z(n8667) );
  XNOR U10908 ( .A(n8702), .B(n8703), .Z(n8686) );
  XNOR U10909 ( .A(n8697), .B(n8698), .Z(n8703) );
  XNOR U10910 ( .A(n8699), .B(n8700), .Z(n8698) );
  XNOR U10911 ( .A(y[805]), .B(x[805]), .Z(n8700) );
  XNOR U10912 ( .A(y[806]), .B(x[806]), .Z(n8699) );
  XNOR U10913 ( .A(y[804]), .B(x[804]), .Z(n8697) );
  XNOR U10914 ( .A(n8691), .B(n8692), .Z(n8702) );
  XNOR U10915 ( .A(y[801]), .B(x[801]), .Z(n8692) );
  XNOR U10916 ( .A(n8693), .B(n8694), .Z(n8691) );
  XNOR U10917 ( .A(y[802]), .B(x[802]), .Z(n8694) );
  XNOR U10918 ( .A(y[803]), .B(x[803]), .Z(n8693) );
  XNOR U10919 ( .A(n8684), .B(n8683), .Z(n8687) );
  XNOR U10920 ( .A(n8679), .B(n8680), .Z(n8683) );
  XNOR U10921 ( .A(y[798]), .B(x[798]), .Z(n8680) );
  XNOR U10922 ( .A(n8681), .B(n8682), .Z(n8679) );
  XNOR U10923 ( .A(y[799]), .B(x[799]), .Z(n8682) );
  XNOR U10924 ( .A(y[800]), .B(x[800]), .Z(n8681) );
  XNOR U10925 ( .A(n8673), .B(n8674), .Z(n8684) );
  XNOR U10926 ( .A(y[795]), .B(x[795]), .Z(n8674) );
  XNOR U10927 ( .A(n8675), .B(n8676), .Z(n8673) );
  XNOR U10928 ( .A(y[796]), .B(x[796]), .Z(n8676) );
  XNOR U10929 ( .A(y[797]), .B(x[797]), .Z(n8675) );
  XOR U10930 ( .A(n8649), .B(n8650), .Z(n8668) );
  XNOR U10931 ( .A(n8665), .B(n8666), .Z(n8650) );
  XNOR U10932 ( .A(n8660), .B(n8661), .Z(n8666) );
  XNOR U10933 ( .A(n8662), .B(n8663), .Z(n8661) );
  XNOR U10934 ( .A(y[793]), .B(x[793]), .Z(n8663) );
  XNOR U10935 ( .A(y[794]), .B(x[794]), .Z(n8662) );
  XNOR U10936 ( .A(y[792]), .B(x[792]), .Z(n8660) );
  XNOR U10937 ( .A(n8654), .B(n8655), .Z(n8665) );
  XNOR U10938 ( .A(y[789]), .B(x[789]), .Z(n8655) );
  XNOR U10939 ( .A(n8656), .B(n8657), .Z(n8654) );
  XNOR U10940 ( .A(y[790]), .B(x[790]), .Z(n8657) );
  XNOR U10941 ( .A(y[791]), .B(x[791]), .Z(n8656) );
  XOR U10942 ( .A(n8648), .B(n8647), .Z(n8649) );
  XNOR U10943 ( .A(n8643), .B(n8644), .Z(n8647) );
  XNOR U10944 ( .A(y[786]), .B(x[786]), .Z(n8644) );
  XNOR U10945 ( .A(n8645), .B(n8646), .Z(n8643) );
  XNOR U10946 ( .A(y[787]), .B(x[787]), .Z(n8646) );
  XNOR U10947 ( .A(y[788]), .B(x[788]), .Z(n8645) );
  XNOR U10948 ( .A(n8637), .B(n8638), .Z(n8648) );
  XNOR U10949 ( .A(y[783]), .B(x[783]), .Z(n8638) );
  XNOR U10950 ( .A(n8639), .B(n8640), .Z(n8637) );
  XNOR U10951 ( .A(y[784]), .B(x[784]), .Z(n8640) );
  XNOR U10952 ( .A(y[785]), .B(x[785]), .Z(n8639) );
  NAND U10953 ( .A(n8704), .B(n8705), .Z(N13137) );
  NANDN U10954 ( .A(n8706), .B(n8707), .Z(n8705) );
  OR U10955 ( .A(n8708), .B(n8709), .Z(n8707) );
  NAND U10956 ( .A(n8708), .B(n8709), .Z(n8704) );
  XOR U10957 ( .A(n8708), .B(n8710), .Z(N13136) );
  XNOR U10958 ( .A(n8706), .B(n8709), .Z(n8710) );
  AND U10959 ( .A(n8711), .B(n8712), .Z(n8709) );
  NANDN U10960 ( .A(n8713), .B(n8714), .Z(n8712) );
  NANDN U10961 ( .A(n8715), .B(n8716), .Z(n8714) );
  NANDN U10962 ( .A(n8716), .B(n8715), .Z(n8711) );
  NAND U10963 ( .A(n8717), .B(n8718), .Z(n8706) );
  NANDN U10964 ( .A(n8719), .B(n8720), .Z(n8718) );
  OR U10965 ( .A(n8721), .B(n8722), .Z(n8720) );
  NAND U10966 ( .A(n8722), .B(n8721), .Z(n8717) );
  AND U10967 ( .A(n8723), .B(n8724), .Z(n8708) );
  NANDN U10968 ( .A(n8725), .B(n8726), .Z(n8724) );
  NANDN U10969 ( .A(n8727), .B(n8728), .Z(n8726) );
  NANDN U10970 ( .A(n8728), .B(n8727), .Z(n8723) );
  XOR U10971 ( .A(n8722), .B(n8729), .Z(N13135) );
  XOR U10972 ( .A(n8719), .B(n8721), .Z(n8729) );
  XNOR U10973 ( .A(n8715), .B(n8730), .Z(n8721) );
  XNOR U10974 ( .A(n8713), .B(n8716), .Z(n8730) );
  NAND U10975 ( .A(n8731), .B(n8732), .Z(n8716) );
  NAND U10976 ( .A(n8733), .B(n8734), .Z(n8732) );
  OR U10977 ( .A(n8735), .B(n8736), .Z(n8733) );
  NANDN U10978 ( .A(n8737), .B(n8735), .Z(n8731) );
  IV U10979 ( .A(n8736), .Z(n8737) );
  NAND U10980 ( .A(n8738), .B(n8739), .Z(n8713) );
  NAND U10981 ( .A(n8740), .B(n8741), .Z(n8739) );
  NANDN U10982 ( .A(n8742), .B(n8743), .Z(n8740) );
  NANDN U10983 ( .A(n8743), .B(n8742), .Z(n8738) );
  AND U10984 ( .A(n8744), .B(n8745), .Z(n8715) );
  NAND U10985 ( .A(n8746), .B(n8747), .Z(n8745) );
  OR U10986 ( .A(n8748), .B(n8749), .Z(n8746) );
  NANDN U10987 ( .A(n8750), .B(n8748), .Z(n8744) );
  NAND U10988 ( .A(n8751), .B(n8752), .Z(n8719) );
  NANDN U10989 ( .A(n8753), .B(n8754), .Z(n8752) );
  OR U10990 ( .A(n8755), .B(n8756), .Z(n8754) );
  NANDN U10991 ( .A(n8757), .B(n8755), .Z(n8751) );
  IV U10992 ( .A(n8756), .Z(n8757) );
  XNOR U10993 ( .A(n8727), .B(n8758), .Z(n8722) );
  XNOR U10994 ( .A(n8725), .B(n8728), .Z(n8758) );
  NAND U10995 ( .A(n8759), .B(n8760), .Z(n8728) );
  NAND U10996 ( .A(n8761), .B(n8762), .Z(n8760) );
  OR U10997 ( .A(n8763), .B(n8764), .Z(n8761) );
  NANDN U10998 ( .A(n8765), .B(n8763), .Z(n8759) );
  IV U10999 ( .A(n8764), .Z(n8765) );
  NAND U11000 ( .A(n8766), .B(n8767), .Z(n8725) );
  NAND U11001 ( .A(n8768), .B(n8769), .Z(n8767) );
  NANDN U11002 ( .A(n8770), .B(n8771), .Z(n8768) );
  NANDN U11003 ( .A(n8771), .B(n8770), .Z(n8766) );
  AND U11004 ( .A(n8772), .B(n8773), .Z(n8727) );
  NAND U11005 ( .A(n8774), .B(n8775), .Z(n8773) );
  OR U11006 ( .A(n8776), .B(n8777), .Z(n8774) );
  NANDN U11007 ( .A(n8778), .B(n8776), .Z(n8772) );
  XNOR U11008 ( .A(n8753), .B(n8779), .Z(N13134) );
  XOR U11009 ( .A(n8755), .B(n8756), .Z(n8779) );
  XNOR U11010 ( .A(n8769), .B(n8780), .Z(n8756) );
  XOR U11011 ( .A(n8770), .B(n8771), .Z(n8780) );
  XOR U11012 ( .A(n8776), .B(n8781), .Z(n8771) );
  XOR U11013 ( .A(n8775), .B(n8778), .Z(n8781) );
  IV U11014 ( .A(n8777), .Z(n8778) );
  NAND U11015 ( .A(n8782), .B(n8783), .Z(n8777) );
  OR U11016 ( .A(n8784), .B(n8785), .Z(n8783) );
  OR U11017 ( .A(n8786), .B(n8787), .Z(n8782) );
  NAND U11018 ( .A(n8788), .B(n8789), .Z(n8775) );
  OR U11019 ( .A(n8790), .B(n8791), .Z(n8789) );
  OR U11020 ( .A(n8792), .B(n8793), .Z(n8788) );
  NOR U11021 ( .A(n8794), .B(n8795), .Z(n8776) );
  ANDN U11022 ( .B(n8796), .A(n8797), .Z(n8770) );
  XNOR U11023 ( .A(n8763), .B(n8798), .Z(n8769) );
  XNOR U11024 ( .A(n8762), .B(n8764), .Z(n8798) );
  NAND U11025 ( .A(n8799), .B(n8800), .Z(n8764) );
  OR U11026 ( .A(n8801), .B(n8802), .Z(n8800) );
  OR U11027 ( .A(n8803), .B(n8804), .Z(n8799) );
  NAND U11028 ( .A(n8805), .B(n8806), .Z(n8762) );
  OR U11029 ( .A(n8807), .B(n8808), .Z(n8806) );
  OR U11030 ( .A(n8809), .B(n8810), .Z(n8805) );
  ANDN U11031 ( .B(n8811), .A(n8812), .Z(n8763) );
  IV U11032 ( .A(n8813), .Z(n8811) );
  ANDN U11033 ( .B(n8814), .A(n8815), .Z(n8755) );
  XOR U11034 ( .A(n8741), .B(n8816), .Z(n8753) );
  XOR U11035 ( .A(n8742), .B(n8743), .Z(n8816) );
  XOR U11036 ( .A(n8748), .B(n8817), .Z(n8743) );
  XOR U11037 ( .A(n8747), .B(n8750), .Z(n8817) );
  IV U11038 ( .A(n8749), .Z(n8750) );
  NAND U11039 ( .A(n8818), .B(n8819), .Z(n8749) );
  OR U11040 ( .A(n8820), .B(n8821), .Z(n8819) );
  OR U11041 ( .A(n8822), .B(n8823), .Z(n8818) );
  NAND U11042 ( .A(n8824), .B(n8825), .Z(n8747) );
  OR U11043 ( .A(n8826), .B(n8827), .Z(n8825) );
  OR U11044 ( .A(n8828), .B(n8829), .Z(n8824) );
  NOR U11045 ( .A(n8830), .B(n8831), .Z(n8748) );
  ANDN U11046 ( .B(n8832), .A(n8833), .Z(n8742) );
  IV U11047 ( .A(n8834), .Z(n8832) );
  XNOR U11048 ( .A(n8735), .B(n8835), .Z(n8741) );
  XNOR U11049 ( .A(n8734), .B(n8736), .Z(n8835) );
  NAND U11050 ( .A(n8836), .B(n8837), .Z(n8736) );
  OR U11051 ( .A(n8838), .B(n8839), .Z(n8837) );
  OR U11052 ( .A(n8840), .B(n8841), .Z(n8836) );
  NAND U11053 ( .A(n8842), .B(n8843), .Z(n8734) );
  OR U11054 ( .A(n8844), .B(n8845), .Z(n8843) );
  OR U11055 ( .A(n8846), .B(n8847), .Z(n8842) );
  ANDN U11056 ( .B(n8848), .A(n8849), .Z(n8735) );
  IV U11057 ( .A(n8850), .Z(n8848) );
  XNOR U11058 ( .A(n8815), .B(n8814), .Z(N13133) );
  XOR U11059 ( .A(n8834), .B(n8833), .Z(n8814) );
  XNOR U11060 ( .A(n8849), .B(n8850), .Z(n8833) );
  XNOR U11061 ( .A(n8844), .B(n8845), .Z(n8850) );
  XNOR U11062 ( .A(n8846), .B(n8847), .Z(n8845) );
  XNOR U11063 ( .A(y[781]), .B(x[781]), .Z(n8847) );
  XNOR U11064 ( .A(y[782]), .B(x[782]), .Z(n8846) );
  XNOR U11065 ( .A(y[780]), .B(x[780]), .Z(n8844) );
  XNOR U11066 ( .A(n8838), .B(n8839), .Z(n8849) );
  XNOR U11067 ( .A(y[777]), .B(x[777]), .Z(n8839) );
  XNOR U11068 ( .A(n8840), .B(n8841), .Z(n8838) );
  XNOR U11069 ( .A(y[778]), .B(x[778]), .Z(n8841) );
  XNOR U11070 ( .A(y[779]), .B(x[779]), .Z(n8840) );
  XNOR U11071 ( .A(n8831), .B(n8830), .Z(n8834) );
  XNOR U11072 ( .A(n8826), .B(n8827), .Z(n8830) );
  XNOR U11073 ( .A(y[774]), .B(x[774]), .Z(n8827) );
  XNOR U11074 ( .A(n8828), .B(n8829), .Z(n8826) );
  XNOR U11075 ( .A(y[775]), .B(x[775]), .Z(n8829) );
  XNOR U11076 ( .A(y[776]), .B(x[776]), .Z(n8828) );
  XNOR U11077 ( .A(n8820), .B(n8821), .Z(n8831) );
  XNOR U11078 ( .A(y[771]), .B(x[771]), .Z(n8821) );
  XNOR U11079 ( .A(n8822), .B(n8823), .Z(n8820) );
  XNOR U11080 ( .A(y[772]), .B(x[772]), .Z(n8823) );
  XNOR U11081 ( .A(y[773]), .B(x[773]), .Z(n8822) );
  XOR U11082 ( .A(n8796), .B(n8797), .Z(n8815) );
  XNOR U11083 ( .A(n8812), .B(n8813), .Z(n8797) );
  XNOR U11084 ( .A(n8807), .B(n8808), .Z(n8813) );
  XNOR U11085 ( .A(n8809), .B(n8810), .Z(n8808) );
  XNOR U11086 ( .A(y[769]), .B(x[769]), .Z(n8810) );
  XNOR U11087 ( .A(y[770]), .B(x[770]), .Z(n8809) );
  XNOR U11088 ( .A(y[768]), .B(x[768]), .Z(n8807) );
  XNOR U11089 ( .A(n8801), .B(n8802), .Z(n8812) );
  XNOR U11090 ( .A(y[765]), .B(x[765]), .Z(n8802) );
  XNOR U11091 ( .A(n8803), .B(n8804), .Z(n8801) );
  XNOR U11092 ( .A(y[766]), .B(x[766]), .Z(n8804) );
  XNOR U11093 ( .A(y[767]), .B(x[767]), .Z(n8803) );
  XOR U11094 ( .A(n8795), .B(n8794), .Z(n8796) );
  XNOR U11095 ( .A(n8790), .B(n8791), .Z(n8794) );
  XNOR U11096 ( .A(y[762]), .B(x[762]), .Z(n8791) );
  XNOR U11097 ( .A(n8792), .B(n8793), .Z(n8790) );
  XNOR U11098 ( .A(y[763]), .B(x[763]), .Z(n8793) );
  XNOR U11099 ( .A(y[764]), .B(x[764]), .Z(n8792) );
  XNOR U11100 ( .A(n8784), .B(n8785), .Z(n8795) );
  XNOR U11101 ( .A(y[759]), .B(x[759]), .Z(n8785) );
  XNOR U11102 ( .A(n8786), .B(n8787), .Z(n8784) );
  XNOR U11103 ( .A(y[760]), .B(x[760]), .Z(n8787) );
  XNOR U11104 ( .A(y[761]), .B(x[761]), .Z(n8786) );
  NAND U11105 ( .A(n8851), .B(n8852), .Z(N13126) );
  NANDN U11106 ( .A(n8853), .B(n8854), .Z(n8852) );
  OR U11107 ( .A(n8855), .B(n8856), .Z(n8854) );
  NAND U11108 ( .A(n8855), .B(n8856), .Z(n8851) );
  XOR U11109 ( .A(n8855), .B(n8857), .Z(N13125) );
  XNOR U11110 ( .A(n8853), .B(n8856), .Z(n8857) );
  AND U11111 ( .A(n8858), .B(n8859), .Z(n8856) );
  NANDN U11112 ( .A(n8860), .B(n8861), .Z(n8859) );
  NANDN U11113 ( .A(n8862), .B(n8863), .Z(n8861) );
  NANDN U11114 ( .A(n8863), .B(n8862), .Z(n8858) );
  NAND U11115 ( .A(n8864), .B(n8865), .Z(n8853) );
  NANDN U11116 ( .A(n8866), .B(n8867), .Z(n8865) );
  OR U11117 ( .A(n8868), .B(n8869), .Z(n8867) );
  NAND U11118 ( .A(n8869), .B(n8868), .Z(n8864) );
  AND U11119 ( .A(n8870), .B(n8871), .Z(n8855) );
  NANDN U11120 ( .A(n8872), .B(n8873), .Z(n8871) );
  NANDN U11121 ( .A(n8874), .B(n8875), .Z(n8873) );
  NANDN U11122 ( .A(n8875), .B(n8874), .Z(n8870) );
  XOR U11123 ( .A(n8869), .B(n8876), .Z(N13124) );
  XOR U11124 ( .A(n8866), .B(n8868), .Z(n8876) );
  XNOR U11125 ( .A(n8862), .B(n8877), .Z(n8868) );
  XNOR U11126 ( .A(n8860), .B(n8863), .Z(n8877) );
  NAND U11127 ( .A(n8878), .B(n8879), .Z(n8863) );
  NAND U11128 ( .A(n8880), .B(n8881), .Z(n8879) );
  OR U11129 ( .A(n8882), .B(n8883), .Z(n8880) );
  NANDN U11130 ( .A(n8884), .B(n8882), .Z(n8878) );
  IV U11131 ( .A(n8883), .Z(n8884) );
  NAND U11132 ( .A(n8885), .B(n8886), .Z(n8860) );
  NAND U11133 ( .A(n8887), .B(n8888), .Z(n8886) );
  NANDN U11134 ( .A(n8889), .B(n8890), .Z(n8887) );
  NANDN U11135 ( .A(n8890), .B(n8889), .Z(n8885) );
  AND U11136 ( .A(n8891), .B(n8892), .Z(n8862) );
  NAND U11137 ( .A(n8893), .B(n8894), .Z(n8892) );
  OR U11138 ( .A(n8895), .B(n8896), .Z(n8893) );
  NANDN U11139 ( .A(n8897), .B(n8895), .Z(n8891) );
  NAND U11140 ( .A(n8898), .B(n8899), .Z(n8866) );
  NANDN U11141 ( .A(n8900), .B(n8901), .Z(n8899) );
  OR U11142 ( .A(n8902), .B(n8903), .Z(n8901) );
  NANDN U11143 ( .A(n8904), .B(n8902), .Z(n8898) );
  IV U11144 ( .A(n8903), .Z(n8904) );
  XNOR U11145 ( .A(n8874), .B(n8905), .Z(n8869) );
  XNOR U11146 ( .A(n8872), .B(n8875), .Z(n8905) );
  NAND U11147 ( .A(n8906), .B(n8907), .Z(n8875) );
  NAND U11148 ( .A(n8908), .B(n8909), .Z(n8907) );
  OR U11149 ( .A(n8910), .B(n8911), .Z(n8908) );
  NANDN U11150 ( .A(n8912), .B(n8910), .Z(n8906) );
  IV U11151 ( .A(n8911), .Z(n8912) );
  NAND U11152 ( .A(n8913), .B(n8914), .Z(n8872) );
  NAND U11153 ( .A(n8915), .B(n8916), .Z(n8914) );
  NANDN U11154 ( .A(n8917), .B(n8918), .Z(n8915) );
  NANDN U11155 ( .A(n8918), .B(n8917), .Z(n8913) );
  AND U11156 ( .A(n8919), .B(n8920), .Z(n8874) );
  NAND U11157 ( .A(n8921), .B(n8922), .Z(n8920) );
  OR U11158 ( .A(n8923), .B(n8924), .Z(n8921) );
  NANDN U11159 ( .A(n8925), .B(n8923), .Z(n8919) );
  XNOR U11160 ( .A(n8900), .B(n8926), .Z(N13123) );
  XOR U11161 ( .A(n8902), .B(n8903), .Z(n8926) );
  XNOR U11162 ( .A(n8916), .B(n8927), .Z(n8903) );
  XOR U11163 ( .A(n8917), .B(n8918), .Z(n8927) );
  XOR U11164 ( .A(n8923), .B(n8928), .Z(n8918) );
  XOR U11165 ( .A(n8922), .B(n8925), .Z(n8928) );
  IV U11166 ( .A(n8924), .Z(n8925) );
  NAND U11167 ( .A(n8929), .B(n8930), .Z(n8924) );
  OR U11168 ( .A(n8931), .B(n8932), .Z(n8930) );
  OR U11169 ( .A(n8933), .B(n8934), .Z(n8929) );
  NAND U11170 ( .A(n8935), .B(n8936), .Z(n8922) );
  OR U11171 ( .A(n8937), .B(n8938), .Z(n8936) );
  OR U11172 ( .A(n8939), .B(n8940), .Z(n8935) );
  NOR U11173 ( .A(n8941), .B(n8942), .Z(n8923) );
  ANDN U11174 ( .B(n8943), .A(n8944), .Z(n8917) );
  XNOR U11175 ( .A(n8910), .B(n8945), .Z(n8916) );
  XNOR U11176 ( .A(n8909), .B(n8911), .Z(n8945) );
  NAND U11177 ( .A(n8946), .B(n8947), .Z(n8911) );
  OR U11178 ( .A(n8948), .B(n8949), .Z(n8947) );
  OR U11179 ( .A(n8950), .B(n8951), .Z(n8946) );
  NAND U11180 ( .A(n8952), .B(n8953), .Z(n8909) );
  OR U11181 ( .A(n8954), .B(n8955), .Z(n8953) );
  OR U11182 ( .A(n8956), .B(n8957), .Z(n8952) );
  ANDN U11183 ( .B(n8958), .A(n8959), .Z(n8910) );
  IV U11184 ( .A(n8960), .Z(n8958) );
  ANDN U11185 ( .B(n8961), .A(n8962), .Z(n8902) );
  XOR U11186 ( .A(n8888), .B(n8963), .Z(n8900) );
  XOR U11187 ( .A(n8889), .B(n8890), .Z(n8963) );
  XOR U11188 ( .A(n8895), .B(n8964), .Z(n8890) );
  XOR U11189 ( .A(n8894), .B(n8897), .Z(n8964) );
  IV U11190 ( .A(n8896), .Z(n8897) );
  NAND U11191 ( .A(n8965), .B(n8966), .Z(n8896) );
  OR U11192 ( .A(n8967), .B(n8968), .Z(n8966) );
  OR U11193 ( .A(n8969), .B(n8970), .Z(n8965) );
  NAND U11194 ( .A(n8971), .B(n8972), .Z(n8894) );
  OR U11195 ( .A(n8973), .B(n8974), .Z(n8972) );
  OR U11196 ( .A(n8975), .B(n8976), .Z(n8971) );
  NOR U11197 ( .A(n8977), .B(n8978), .Z(n8895) );
  ANDN U11198 ( .B(n8979), .A(n8980), .Z(n8889) );
  IV U11199 ( .A(n8981), .Z(n8979) );
  XNOR U11200 ( .A(n8882), .B(n8982), .Z(n8888) );
  XNOR U11201 ( .A(n8881), .B(n8883), .Z(n8982) );
  NAND U11202 ( .A(n8983), .B(n8984), .Z(n8883) );
  OR U11203 ( .A(n8985), .B(n8986), .Z(n8984) );
  OR U11204 ( .A(n8987), .B(n8988), .Z(n8983) );
  NAND U11205 ( .A(n8989), .B(n8990), .Z(n8881) );
  OR U11206 ( .A(n8991), .B(n8992), .Z(n8990) );
  OR U11207 ( .A(n8993), .B(n8994), .Z(n8989) );
  ANDN U11208 ( .B(n8995), .A(n8996), .Z(n8882) );
  IV U11209 ( .A(n8997), .Z(n8995) );
  XNOR U11210 ( .A(n8962), .B(n8961), .Z(N13122) );
  XOR U11211 ( .A(n8981), .B(n8980), .Z(n8961) );
  XNOR U11212 ( .A(n8996), .B(n8997), .Z(n8980) );
  XNOR U11213 ( .A(n8991), .B(n8992), .Z(n8997) );
  XNOR U11214 ( .A(n8993), .B(n8994), .Z(n8992) );
  XNOR U11215 ( .A(y[757]), .B(x[757]), .Z(n8994) );
  XNOR U11216 ( .A(y[758]), .B(x[758]), .Z(n8993) );
  XNOR U11217 ( .A(y[756]), .B(x[756]), .Z(n8991) );
  XNOR U11218 ( .A(n8985), .B(n8986), .Z(n8996) );
  XNOR U11219 ( .A(y[753]), .B(x[753]), .Z(n8986) );
  XNOR U11220 ( .A(n8987), .B(n8988), .Z(n8985) );
  XNOR U11221 ( .A(y[754]), .B(x[754]), .Z(n8988) );
  XNOR U11222 ( .A(y[755]), .B(x[755]), .Z(n8987) );
  XNOR U11223 ( .A(n8978), .B(n8977), .Z(n8981) );
  XNOR U11224 ( .A(n8973), .B(n8974), .Z(n8977) );
  XNOR U11225 ( .A(y[750]), .B(x[750]), .Z(n8974) );
  XNOR U11226 ( .A(n8975), .B(n8976), .Z(n8973) );
  XNOR U11227 ( .A(y[751]), .B(x[751]), .Z(n8976) );
  XNOR U11228 ( .A(y[752]), .B(x[752]), .Z(n8975) );
  XNOR U11229 ( .A(n8967), .B(n8968), .Z(n8978) );
  XNOR U11230 ( .A(y[747]), .B(x[747]), .Z(n8968) );
  XNOR U11231 ( .A(n8969), .B(n8970), .Z(n8967) );
  XNOR U11232 ( .A(y[748]), .B(x[748]), .Z(n8970) );
  XNOR U11233 ( .A(y[749]), .B(x[749]), .Z(n8969) );
  XOR U11234 ( .A(n8943), .B(n8944), .Z(n8962) );
  XNOR U11235 ( .A(n8959), .B(n8960), .Z(n8944) );
  XNOR U11236 ( .A(n8954), .B(n8955), .Z(n8960) );
  XNOR U11237 ( .A(n8956), .B(n8957), .Z(n8955) );
  XNOR U11238 ( .A(y[745]), .B(x[745]), .Z(n8957) );
  XNOR U11239 ( .A(y[746]), .B(x[746]), .Z(n8956) );
  XNOR U11240 ( .A(y[744]), .B(x[744]), .Z(n8954) );
  XNOR U11241 ( .A(n8948), .B(n8949), .Z(n8959) );
  XNOR U11242 ( .A(y[741]), .B(x[741]), .Z(n8949) );
  XNOR U11243 ( .A(n8950), .B(n8951), .Z(n8948) );
  XNOR U11244 ( .A(y[742]), .B(x[742]), .Z(n8951) );
  XNOR U11245 ( .A(y[743]), .B(x[743]), .Z(n8950) );
  XOR U11246 ( .A(n8942), .B(n8941), .Z(n8943) );
  XNOR U11247 ( .A(n8937), .B(n8938), .Z(n8941) );
  XNOR U11248 ( .A(y[738]), .B(x[738]), .Z(n8938) );
  XNOR U11249 ( .A(n8939), .B(n8940), .Z(n8937) );
  XNOR U11250 ( .A(y[739]), .B(x[739]), .Z(n8940) );
  XNOR U11251 ( .A(y[740]), .B(x[740]), .Z(n8939) );
  XNOR U11252 ( .A(n8931), .B(n8932), .Z(n8942) );
  XNOR U11253 ( .A(y[735]), .B(x[735]), .Z(n8932) );
  XNOR U11254 ( .A(n8933), .B(n8934), .Z(n8931) );
  XNOR U11255 ( .A(y[736]), .B(x[736]), .Z(n8934) );
  XNOR U11256 ( .A(y[737]), .B(x[737]), .Z(n8933) );
  NAND U11257 ( .A(n8998), .B(n8999), .Z(N13115) );
  NANDN U11258 ( .A(n9000), .B(n9001), .Z(n8999) );
  OR U11259 ( .A(n9002), .B(n9003), .Z(n9001) );
  NAND U11260 ( .A(n9002), .B(n9003), .Z(n8998) );
  XOR U11261 ( .A(n9002), .B(n9004), .Z(N13114) );
  XNOR U11262 ( .A(n9000), .B(n9003), .Z(n9004) );
  AND U11263 ( .A(n9005), .B(n9006), .Z(n9003) );
  NANDN U11264 ( .A(n9007), .B(n9008), .Z(n9006) );
  NANDN U11265 ( .A(n9009), .B(n9010), .Z(n9008) );
  NANDN U11266 ( .A(n9010), .B(n9009), .Z(n9005) );
  NAND U11267 ( .A(n9011), .B(n9012), .Z(n9000) );
  NANDN U11268 ( .A(n9013), .B(n9014), .Z(n9012) );
  OR U11269 ( .A(n9015), .B(n9016), .Z(n9014) );
  NAND U11270 ( .A(n9016), .B(n9015), .Z(n9011) );
  AND U11271 ( .A(n9017), .B(n9018), .Z(n9002) );
  NANDN U11272 ( .A(n9019), .B(n9020), .Z(n9018) );
  NANDN U11273 ( .A(n9021), .B(n9022), .Z(n9020) );
  NANDN U11274 ( .A(n9022), .B(n9021), .Z(n9017) );
  XOR U11275 ( .A(n9016), .B(n9023), .Z(N13113) );
  XOR U11276 ( .A(n9013), .B(n9015), .Z(n9023) );
  XNOR U11277 ( .A(n9009), .B(n9024), .Z(n9015) );
  XNOR U11278 ( .A(n9007), .B(n9010), .Z(n9024) );
  NAND U11279 ( .A(n9025), .B(n9026), .Z(n9010) );
  NAND U11280 ( .A(n9027), .B(n9028), .Z(n9026) );
  OR U11281 ( .A(n9029), .B(n9030), .Z(n9027) );
  NANDN U11282 ( .A(n9031), .B(n9029), .Z(n9025) );
  IV U11283 ( .A(n9030), .Z(n9031) );
  NAND U11284 ( .A(n9032), .B(n9033), .Z(n9007) );
  NAND U11285 ( .A(n9034), .B(n9035), .Z(n9033) );
  NANDN U11286 ( .A(n9036), .B(n9037), .Z(n9034) );
  NANDN U11287 ( .A(n9037), .B(n9036), .Z(n9032) );
  AND U11288 ( .A(n9038), .B(n9039), .Z(n9009) );
  NAND U11289 ( .A(n9040), .B(n9041), .Z(n9039) );
  OR U11290 ( .A(n9042), .B(n9043), .Z(n9040) );
  NANDN U11291 ( .A(n9044), .B(n9042), .Z(n9038) );
  NAND U11292 ( .A(n9045), .B(n9046), .Z(n9013) );
  NANDN U11293 ( .A(n9047), .B(n9048), .Z(n9046) );
  OR U11294 ( .A(n9049), .B(n9050), .Z(n9048) );
  NANDN U11295 ( .A(n9051), .B(n9049), .Z(n9045) );
  IV U11296 ( .A(n9050), .Z(n9051) );
  XNOR U11297 ( .A(n9021), .B(n9052), .Z(n9016) );
  XNOR U11298 ( .A(n9019), .B(n9022), .Z(n9052) );
  NAND U11299 ( .A(n9053), .B(n9054), .Z(n9022) );
  NAND U11300 ( .A(n9055), .B(n9056), .Z(n9054) );
  OR U11301 ( .A(n9057), .B(n9058), .Z(n9055) );
  NANDN U11302 ( .A(n9059), .B(n9057), .Z(n9053) );
  IV U11303 ( .A(n9058), .Z(n9059) );
  NAND U11304 ( .A(n9060), .B(n9061), .Z(n9019) );
  NAND U11305 ( .A(n9062), .B(n9063), .Z(n9061) );
  NANDN U11306 ( .A(n9064), .B(n9065), .Z(n9062) );
  NANDN U11307 ( .A(n9065), .B(n9064), .Z(n9060) );
  AND U11308 ( .A(n9066), .B(n9067), .Z(n9021) );
  NAND U11309 ( .A(n9068), .B(n9069), .Z(n9067) );
  OR U11310 ( .A(n9070), .B(n9071), .Z(n9068) );
  NANDN U11311 ( .A(n9072), .B(n9070), .Z(n9066) );
  XNOR U11312 ( .A(n9047), .B(n9073), .Z(N13112) );
  XOR U11313 ( .A(n9049), .B(n9050), .Z(n9073) );
  XNOR U11314 ( .A(n9063), .B(n9074), .Z(n9050) );
  XOR U11315 ( .A(n9064), .B(n9065), .Z(n9074) );
  XOR U11316 ( .A(n9070), .B(n9075), .Z(n9065) );
  XOR U11317 ( .A(n9069), .B(n9072), .Z(n9075) );
  IV U11318 ( .A(n9071), .Z(n9072) );
  NAND U11319 ( .A(n9076), .B(n9077), .Z(n9071) );
  OR U11320 ( .A(n9078), .B(n9079), .Z(n9077) );
  OR U11321 ( .A(n9080), .B(n9081), .Z(n9076) );
  NAND U11322 ( .A(n9082), .B(n9083), .Z(n9069) );
  OR U11323 ( .A(n9084), .B(n9085), .Z(n9083) );
  OR U11324 ( .A(n9086), .B(n9087), .Z(n9082) );
  NOR U11325 ( .A(n9088), .B(n9089), .Z(n9070) );
  ANDN U11326 ( .B(n9090), .A(n9091), .Z(n9064) );
  XNOR U11327 ( .A(n9057), .B(n9092), .Z(n9063) );
  XNOR U11328 ( .A(n9056), .B(n9058), .Z(n9092) );
  NAND U11329 ( .A(n9093), .B(n9094), .Z(n9058) );
  OR U11330 ( .A(n9095), .B(n9096), .Z(n9094) );
  OR U11331 ( .A(n9097), .B(n9098), .Z(n9093) );
  NAND U11332 ( .A(n9099), .B(n9100), .Z(n9056) );
  OR U11333 ( .A(n9101), .B(n9102), .Z(n9100) );
  OR U11334 ( .A(n9103), .B(n9104), .Z(n9099) );
  ANDN U11335 ( .B(n9105), .A(n9106), .Z(n9057) );
  IV U11336 ( .A(n9107), .Z(n9105) );
  ANDN U11337 ( .B(n9108), .A(n9109), .Z(n9049) );
  XOR U11338 ( .A(n9035), .B(n9110), .Z(n9047) );
  XOR U11339 ( .A(n9036), .B(n9037), .Z(n9110) );
  XOR U11340 ( .A(n9042), .B(n9111), .Z(n9037) );
  XOR U11341 ( .A(n9041), .B(n9044), .Z(n9111) );
  IV U11342 ( .A(n9043), .Z(n9044) );
  NAND U11343 ( .A(n9112), .B(n9113), .Z(n9043) );
  OR U11344 ( .A(n9114), .B(n9115), .Z(n9113) );
  OR U11345 ( .A(n9116), .B(n9117), .Z(n9112) );
  NAND U11346 ( .A(n9118), .B(n9119), .Z(n9041) );
  OR U11347 ( .A(n9120), .B(n9121), .Z(n9119) );
  OR U11348 ( .A(n9122), .B(n9123), .Z(n9118) );
  NOR U11349 ( .A(n9124), .B(n9125), .Z(n9042) );
  ANDN U11350 ( .B(n9126), .A(n9127), .Z(n9036) );
  IV U11351 ( .A(n9128), .Z(n9126) );
  XNOR U11352 ( .A(n9029), .B(n9129), .Z(n9035) );
  XNOR U11353 ( .A(n9028), .B(n9030), .Z(n9129) );
  NAND U11354 ( .A(n9130), .B(n9131), .Z(n9030) );
  OR U11355 ( .A(n9132), .B(n9133), .Z(n9131) );
  OR U11356 ( .A(n9134), .B(n9135), .Z(n9130) );
  NAND U11357 ( .A(n9136), .B(n9137), .Z(n9028) );
  OR U11358 ( .A(n9138), .B(n9139), .Z(n9137) );
  OR U11359 ( .A(n9140), .B(n9141), .Z(n9136) );
  ANDN U11360 ( .B(n9142), .A(n9143), .Z(n9029) );
  IV U11361 ( .A(n9144), .Z(n9142) );
  XNOR U11362 ( .A(n9109), .B(n9108), .Z(N13111) );
  XOR U11363 ( .A(n9128), .B(n9127), .Z(n9108) );
  XNOR U11364 ( .A(n9143), .B(n9144), .Z(n9127) );
  XNOR U11365 ( .A(n9138), .B(n9139), .Z(n9144) );
  XNOR U11366 ( .A(n9140), .B(n9141), .Z(n9139) );
  XNOR U11367 ( .A(y[733]), .B(x[733]), .Z(n9141) );
  XNOR U11368 ( .A(y[734]), .B(x[734]), .Z(n9140) );
  XNOR U11369 ( .A(y[732]), .B(x[732]), .Z(n9138) );
  XNOR U11370 ( .A(n9132), .B(n9133), .Z(n9143) );
  XNOR U11371 ( .A(y[729]), .B(x[729]), .Z(n9133) );
  XNOR U11372 ( .A(n9134), .B(n9135), .Z(n9132) );
  XNOR U11373 ( .A(y[730]), .B(x[730]), .Z(n9135) );
  XNOR U11374 ( .A(y[731]), .B(x[731]), .Z(n9134) );
  XNOR U11375 ( .A(n9125), .B(n9124), .Z(n9128) );
  XNOR U11376 ( .A(n9120), .B(n9121), .Z(n9124) );
  XNOR U11377 ( .A(y[726]), .B(x[726]), .Z(n9121) );
  XNOR U11378 ( .A(n9122), .B(n9123), .Z(n9120) );
  XNOR U11379 ( .A(y[727]), .B(x[727]), .Z(n9123) );
  XNOR U11380 ( .A(y[728]), .B(x[728]), .Z(n9122) );
  XNOR U11381 ( .A(n9114), .B(n9115), .Z(n9125) );
  XNOR U11382 ( .A(y[723]), .B(x[723]), .Z(n9115) );
  XNOR U11383 ( .A(n9116), .B(n9117), .Z(n9114) );
  XNOR U11384 ( .A(y[724]), .B(x[724]), .Z(n9117) );
  XNOR U11385 ( .A(y[725]), .B(x[725]), .Z(n9116) );
  XOR U11386 ( .A(n9090), .B(n9091), .Z(n9109) );
  XNOR U11387 ( .A(n9106), .B(n9107), .Z(n9091) );
  XNOR U11388 ( .A(n9101), .B(n9102), .Z(n9107) );
  XNOR U11389 ( .A(n9103), .B(n9104), .Z(n9102) );
  XNOR U11390 ( .A(y[721]), .B(x[721]), .Z(n9104) );
  XNOR U11391 ( .A(y[722]), .B(x[722]), .Z(n9103) );
  XNOR U11392 ( .A(y[720]), .B(x[720]), .Z(n9101) );
  XNOR U11393 ( .A(n9095), .B(n9096), .Z(n9106) );
  XNOR U11394 ( .A(y[717]), .B(x[717]), .Z(n9096) );
  XNOR U11395 ( .A(n9097), .B(n9098), .Z(n9095) );
  XNOR U11396 ( .A(y[718]), .B(x[718]), .Z(n9098) );
  XNOR U11397 ( .A(y[719]), .B(x[719]), .Z(n9097) );
  XOR U11398 ( .A(n9089), .B(n9088), .Z(n9090) );
  XNOR U11399 ( .A(n9084), .B(n9085), .Z(n9088) );
  XNOR U11400 ( .A(y[714]), .B(x[714]), .Z(n9085) );
  XNOR U11401 ( .A(n9086), .B(n9087), .Z(n9084) );
  XNOR U11402 ( .A(y[715]), .B(x[715]), .Z(n9087) );
  XNOR U11403 ( .A(y[716]), .B(x[716]), .Z(n9086) );
  XNOR U11404 ( .A(n9078), .B(n9079), .Z(n9089) );
  XNOR U11405 ( .A(y[711]), .B(x[711]), .Z(n9079) );
  XNOR U11406 ( .A(n9080), .B(n9081), .Z(n9078) );
  XNOR U11407 ( .A(y[712]), .B(x[712]), .Z(n9081) );
  XNOR U11408 ( .A(y[713]), .B(x[713]), .Z(n9080) );
  NAND U11409 ( .A(n9145), .B(n9146), .Z(N13104) );
  NANDN U11410 ( .A(n9147), .B(n9148), .Z(n9146) );
  OR U11411 ( .A(n9149), .B(n9150), .Z(n9148) );
  NAND U11412 ( .A(n9149), .B(n9150), .Z(n9145) );
  XOR U11413 ( .A(n9149), .B(n9151), .Z(N13103) );
  XNOR U11414 ( .A(n9147), .B(n9150), .Z(n9151) );
  AND U11415 ( .A(n9152), .B(n9153), .Z(n9150) );
  NANDN U11416 ( .A(n9154), .B(n9155), .Z(n9153) );
  NANDN U11417 ( .A(n9156), .B(n9157), .Z(n9155) );
  NANDN U11418 ( .A(n9157), .B(n9156), .Z(n9152) );
  NAND U11419 ( .A(n9158), .B(n9159), .Z(n9147) );
  NANDN U11420 ( .A(n9160), .B(n9161), .Z(n9159) );
  OR U11421 ( .A(n9162), .B(n9163), .Z(n9161) );
  NAND U11422 ( .A(n9163), .B(n9162), .Z(n9158) );
  AND U11423 ( .A(n9164), .B(n9165), .Z(n9149) );
  NANDN U11424 ( .A(n9166), .B(n9167), .Z(n9165) );
  NANDN U11425 ( .A(n9168), .B(n9169), .Z(n9167) );
  NANDN U11426 ( .A(n9169), .B(n9168), .Z(n9164) );
  XOR U11427 ( .A(n9163), .B(n9170), .Z(N13102) );
  XOR U11428 ( .A(n9160), .B(n9162), .Z(n9170) );
  XNOR U11429 ( .A(n9156), .B(n9171), .Z(n9162) );
  XNOR U11430 ( .A(n9154), .B(n9157), .Z(n9171) );
  NAND U11431 ( .A(n9172), .B(n9173), .Z(n9157) );
  NAND U11432 ( .A(n9174), .B(n9175), .Z(n9173) );
  OR U11433 ( .A(n9176), .B(n9177), .Z(n9174) );
  NANDN U11434 ( .A(n9178), .B(n9176), .Z(n9172) );
  IV U11435 ( .A(n9177), .Z(n9178) );
  NAND U11436 ( .A(n9179), .B(n9180), .Z(n9154) );
  NAND U11437 ( .A(n9181), .B(n9182), .Z(n9180) );
  NANDN U11438 ( .A(n9183), .B(n9184), .Z(n9181) );
  NANDN U11439 ( .A(n9184), .B(n9183), .Z(n9179) );
  AND U11440 ( .A(n9185), .B(n9186), .Z(n9156) );
  NAND U11441 ( .A(n9187), .B(n9188), .Z(n9186) );
  OR U11442 ( .A(n9189), .B(n9190), .Z(n9187) );
  NANDN U11443 ( .A(n9191), .B(n9189), .Z(n9185) );
  NAND U11444 ( .A(n9192), .B(n9193), .Z(n9160) );
  NANDN U11445 ( .A(n9194), .B(n9195), .Z(n9193) );
  OR U11446 ( .A(n9196), .B(n9197), .Z(n9195) );
  NANDN U11447 ( .A(n9198), .B(n9196), .Z(n9192) );
  IV U11448 ( .A(n9197), .Z(n9198) );
  XNOR U11449 ( .A(n9168), .B(n9199), .Z(n9163) );
  XNOR U11450 ( .A(n9166), .B(n9169), .Z(n9199) );
  NAND U11451 ( .A(n9200), .B(n9201), .Z(n9169) );
  NAND U11452 ( .A(n9202), .B(n9203), .Z(n9201) );
  OR U11453 ( .A(n9204), .B(n9205), .Z(n9202) );
  NANDN U11454 ( .A(n9206), .B(n9204), .Z(n9200) );
  IV U11455 ( .A(n9205), .Z(n9206) );
  NAND U11456 ( .A(n9207), .B(n9208), .Z(n9166) );
  NAND U11457 ( .A(n9209), .B(n9210), .Z(n9208) );
  NANDN U11458 ( .A(n9211), .B(n9212), .Z(n9209) );
  NANDN U11459 ( .A(n9212), .B(n9211), .Z(n9207) );
  AND U11460 ( .A(n9213), .B(n9214), .Z(n9168) );
  NAND U11461 ( .A(n9215), .B(n9216), .Z(n9214) );
  OR U11462 ( .A(n9217), .B(n9218), .Z(n9215) );
  NANDN U11463 ( .A(n9219), .B(n9217), .Z(n9213) );
  XNOR U11464 ( .A(n9194), .B(n9220), .Z(N13101) );
  XOR U11465 ( .A(n9196), .B(n9197), .Z(n9220) );
  XNOR U11466 ( .A(n9210), .B(n9221), .Z(n9197) );
  XOR U11467 ( .A(n9211), .B(n9212), .Z(n9221) );
  XOR U11468 ( .A(n9217), .B(n9222), .Z(n9212) );
  XOR U11469 ( .A(n9216), .B(n9219), .Z(n9222) );
  IV U11470 ( .A(n9218), .Z(n9219) );
  NAND U11471 ( .A(n9223), .B(n9224), .Z(n9218) );
  OR U11472 ( .A(n9225), .B(n9226), .Z(n9224) );
  OR U11473 ( .A(n9227), .B(n9228), .Z(n9223) );
  NAND U11474 ( .A(n9229), .B(n9230), .Z(n9216) );
  OR U11475 ( .A(n9231), .B(n9232), .Z(n9230) );
  OR U11476 ( .A(n9233), .B(n9234), .Z(n9229) );
  NOR U11477 ( .A(n9235), .B(n9236), .Z(n9217) );
  ANDN U11478 ( .B(n9237), .A(n9238), .Z(n9211) );
  XNOR U11479 ( .A(n9204), .B(n9239), .Z(n9210) );
  XNOR U11480 ( .A(n9203), .B(n9205), .Z(n9239) );
  NAND U11481 ( .A(n9240), .B(n9241), .Z(n9205) );
  OR U11482 ( .A(n9242), .B(n9243), .Z(n9241) );
  OR U11483 ( .A(n9244), .B(n9245), .Z(n9240) );
  NAND U11484 ( .A(n9246), .B(n9247), .Z(n9203) );
  OR U11485 ( .A(n9248), .B(n9249), .Z(n9247) );
  OR U11486 ( .A(n9250), .B(n9251), .Z(n9246) );
  ANDN U11487 ( .B(n9252), .A(n9253), .Z(n9204) );
  IV U11488 ( .A(n9254), .Z(n9252) );
  ANDN U11489 ( .B(n9255), .A(n9256), .Z(n9196) );
  XOR U11490 ( .A(n9182), .B(n9257), .Z(n9194) );
  XOR U11491 ( .A(n9183), .B(n9184), .Z(n9257) );
  XOR U11492 ( .A(n9189), .B(n9258), .Z(n9184) );
  XOR U11493 ( .A(n9188), .B(n9191), .Z(n9258) );
  IV U11494 ( .A(n9190), .Z(n9191) );
  NAND U11495 ( .A(n9259), .B(n9260), .Z(n9190) );
  OR U11496 ( .A(n9261), .B(n9262), .Z(n9260) );
  OR U11497 ( .A(n9263), .B(n9264), .Z(n9259) );
  NAND U11498 ( .A(n9265), .B(n9266), .Z(n9188) );
  OR U11499 ( .A(n9267), .B(n9268), .Z(n9266) );
  OR U11500 ( .A(n9269), .B(n9270), .Z(n9265) );
  NOR U11501 ( .A(n9271), .B(n9272), .Z(n9189) );
  ANDN U11502 ( .B(n9273), .A(n9274), .Z(n9183) );
  IV U11503 ( .A(n9275), .Z(n9273) );
  XNOR U11504 ( .A(n9176), .B(n9276), .Z(n9182) );
  XNOR U11505 ( .A(n9175), .B(n9177), .Z(n9276) );
  NAND U11506 ( .A(n9277), .B(n9278), .Z(n9177) );
  OR U11507 ( .A(n9279), .B(n9280), .Z(n9278) );
  OR U11508 ( .A(n9281), .B(n9282), .Z(n9277) );
  NAND U11509 ( .A(n9283), .B(n9284), .Z(n9175) );
  OR U11510 ( .A(n9285), .B(n9286), .Z(n9284) );
  OR U11511 ( .A(n9287), .B(n9288), .Z(n9283) );
  ANDN U11512 ( .B(n9289), .A(n9290), .Z(n9176) );
  IV U11513 ( .A(n9291), .Z(n9289) );
  XNOR U11514 ( .A(n9256), .B(n9255), .Z(N13100) );
  XOR U11515 ( .A(n9275), .B(n9274), .Z(n9255) );
  XNOR U11516 ( .A(n9290), .B(n9291), .Z(n9274) );
  XNOR U11517 ( .A(n9285), .B(n9286), .Z(n9291) );
  XNOR U11518 ( .A(n9287), .B(n9288), .Z(n9286) );
  XNOR U11519 ( .A(y[709]), .B(x[709]), .Z(n9288) );
  XNOR U11520 ( .A(y[710]), .B(x[710]), .Z(n9287) );
  XNOR U11521 ( .A(y[708]), .B(x[708]), .Z(n9285) );
  XNOR U11522 ( .A(n9279), .B(n9280), .Z(n9290) );
  XNOR U11523 ( .A(y[705]), .B(x[705]), .Z(n9280) );
  XNOR U11524 ( .A(n9281), .B(n9282), .Z(n9279) );
  XNOR U11525 ( .A(y[706]), .B(x[706]), .Z(n9282) );
  XNOR U11526 ( .A(y[707]), .B(x[707]), .Z(n9281) );
  XNOR U11527 ( .A(n9272), .B(n9271), .Z(n9275) );
  XNOR U11528 ( .A(n9267), .B(n9268), .Z(n9271) );
  XNOR U11529 ( .A(y[702]), .B(x[702]), .Z(n9268) );
  XNOR U11530 ( .A(n9269), .B(n9270), .Z(n9267) );
  XNOR U11531 ( .A(y[703]), .B(x[703]), .Z(n9270) );
  XNOR U11532 ( .A(y[704]), .B(x[704]), .Z(n9269) );
  XNOR U11533 ( .A(n9261), .B(n9262), .Z(n9272) );
  XNOR U11534 ( .A(y[699]), .B(x[699]), .Z(n9262) );
  XNOR U11535 ( .A(n9263), .B(n9264), .Z(n9261) );
  XNOR U11536 ( .A(y[700]), .B(x[700]), .Z(n9264) );
  XNOR U11537 ( .A(y[701]), .B(x[701]), .Z(n9263) );
  XOR U11538 ( .A(n9237), .B(n9238), .Z(n9256) );
  XNOR U11539 ( .A(n9253), .B(n9254), .Z(n9238) );
  XNOR U11540 ( .A(n9248), .B(n9249), .Z(n9254) );
  XNOR U11541 ( .A(n9250), .B(n9251), .Z(n9249) );
  XNOR U11542 ( .A(y[697]), .B(x[697]), .Z(n9251) );
  XNOR U11543 ( .A(y[698]), .B(x[698]), .Z(n9250) );
  XNOR U11544 ( .A(y[696]), .B(x[696]), .Z(n9248) );
  XNOR U11545 ( .A(n9242), .B(n9243), .Z(n9253) );
  XNOR U11546 ( .A(y[693]), .B(x[693]), .Z(n9243) );
  XNOR U11547 ( .A(n9244), .B(n9245), .Z(n9242) );
  XNOR U11548 ( .A(y[694]), .B(x[694]), .Z(n9245) );
  XNOR U11549 ( .A(y[695]), .B(x[695]), .Z(n9244) );
  XOR U11550 ( .A(n9236), .B(n9235), .Z(n9237) );
  XNOR U11551 ( .A(n9231), .B(n9232), .Z(n9235) );
  XNOR U11552 ( .A(y[690]), .B(x[690]), .Z(n9232) );
  XNOR U11553 ( .A(n9233), .B(n9234), .Z(n9231) );
  XNOR U11554 ( .A(y[691]), .B(x[691]), .Z(n9234) );
  XNOR U11555 ( .A(y[692]), .B(x[692]), .Z(n9233) );
  XNOR U11556 ( .A(n9225), .B(n9226), .Z(n9236) );
  XNOR U11557 ( .A(y[687]), .B(x[687]), .Z(n9226) );
  XNOR U11558 ( .A(n9227), .B(n9228), .Z(n9225) );
  XNOR U11559 ( .A(y[688]), .B(x[688]), .Z(n9228) );
  XNOR U11560 ( .A(y[689]), .B(x[689]), .Z(n9227) );
  NAND U11561 ( .A(n9292), .B(n9293), .Z(N13093) );
  NANDN U11562 ( .A(n9294), .B(n9295), .Z(n9293) );
  OR U11563 ( .A(n9296), .B(n9297), .Z(n9295) );
  NAND U11564 ( .A(n9296), .B(n9297), .Z(n9292) );
  XOR U11565 ( .A(n9296), .B(n9298), .Z(N13092) );
  XNOR U11566 ( .A(n9294), .B(n9297), .Z(n9298) );
  AND U11567 ( .A(n9299), .B(n9300), .Z(n9297) );
  NANDN U11568 ( .A(n9301), .B(n9302), .Z(n9300) );
  NANDN U11569 ( .A(n9303), .B(n9304), .Z(n9302) );
  NANDN U11570 ( .A(n9304), .B(n9303), .Z(n9299) );
  NAND U11571 ( .A(n9305), .B(n9306), .Z(n9294) );
  NANDN U11572 ( .A(n9307), .B(n9308), .Z(n9306) );
  OR U11573 ( .A(n9309), .B(n9310), .Z(n9308) );
  NAND U11574 ( .A(n9310), .B(n9309), .Z(n9305) );
  AND U11575 ( .A(n9311), .B(n9312), .Z(n9296) );
  NANDN U11576 ( .A(n9313), .B(n9314), .Z(n9312) );
  NANDN U11577 ( .A(n9315), .B(n9316), .Z(n9314) );
  NANDN U11578 ( .A(n9316), .B(n9315), .Z(n9311) );
  XOR U11579 ( .A(n9310), .B(n9317), .Z(N13091) );
  XOR U11580 ( .A(n9307), .B(n9309), .Z(n9317) );
  XNOR U11581 ( .A(n9303), .B(n9318), .Z(n9309) );
  XNOR U11582 ( .A(n9301), .B(n9304), .Z(n9318) );
  NAND U11583 ( .A(n9319), .B(n9320), .Z(n9304) );
  NAND U11584 ( .A(n9321), .B(n9322), .Z(n9320) );
  OR U11585 ( .A(n9323), .B(n9324), .Z(n9321) );
  NANDN U11586 ( .A(n9325), .B(n9323), .Z(n9319) );
  IV U11587 ( .A(n9324), .Z(n9325) );
  NAND U11588 ( .A(n9326), .B(n9327), .Z(n9301) );
  NAND U11589 ( .A(n9328), .B(n9329), .Z(n9327) );
  NANDN U11590 ( .A(n9330), .B(n9331), .Z(n9328) );
  NANDN U11591 ( .A(n9331), .B(n9330), .Z(n9326) );
  AND U11592 ( .A(n9332), .B(n9333), .Z(n9303) );
  NAND U11593 ( .A(n9334), .B(n9335), .Z(n9333) );
  OR U11594 ( .A(n9336), .B(n9337), .Z(n9334) );
  NANDN U11595 ( .A(n9338), .B(n9336), .Z(n9332) );
  NAND U11596 ( .A(n9339), .B(n9340), .Z(n9307) );
  NANDN U11597 ( .A(n9341), .B(n9342), .Z(n9340) );
  OR U11598 ( .A(n9343), .B(n9344), .Z(n9342) );
  NANDN U11599 ( .A(n9345), .B(n9343), .Z(n9339) );
  IV U11600 ( .A(n9344), .Z(n9345) );
  XNOR U11601 ( .A(n9315), .B(n9346), .Z(n9310) );
  XNOR U11602 ( .A(n9313), .B(n9316), .Z(n9346) );
  NAND U11603 ( .A(n9347), .B(n9348), .Z(n9316) );
  NAND U11604 ( .A(n9349), .B(n9350), .Z(n9348) );
  OR U11605 ( .A(n9351), .B(n9352), .Z(n9349) );
  NANDN U11606 ( .A(n9353), .B(n9351), .Z(n9347) );
  IV U11607 ( .A(n9352), .Z(n9353) );
  NAND U11608 ( .A(n9354), .B(n9355), .Z(n9313) );
  NAND U11609 ( .A(n9356), .B(n9357), .Z(n9355) );
  NANDN U11610 ( .A(n9358), .B(n9359), .Z(n9356) );
  NANDN U11611 ( .A(n9359), .B(n9358), .Z(n9354) );
  AND U11612 ( .A(n9360), .B(n9361), .Z(n9315) );
  NAND U11613 ( .A(n9362), .B(n9363), .Z(n9361) );
  OR U11614 ( .A(n9364), .B(n9365), .Z(n9362) );
  NANDN U11615 ( .A(n9366), .B(n9364), .Z(n9360) );
  XNOR U11616 ( .A(n9341), .B(n9367), .Z(N13090) );
  XOR U11617 ( .A(n9343), .B(n9344), .Z(n9367) );
  XNOR U11618 ( .A(n9357), .B(n9368), .Z(n9344) );
  XOR U11619 ( .A(n9358), .B(n9359), .Z(n9368) );
  XOR U11620 ( .A(n9364), .B(n9369), .Z(n9359) );
  XOR U11621 ( .A(n9363), .B(n9366), .Z(n9369) );
  IV U11622 ( .A(n9365), .Z(n9366) );
  NAND U11623 ( .A(n9370), .B(n9371), .Z(n9365) );
  OR U11624 ( .A(n9372), .B(n9373), .Z(n9371) );
  OR U11625 ( .A(n9374), .B(n9375), .Z(n9370) );
  NAND U11626 ( .A(n9376), .B(n9377), .Z(n9363) );
  OR U11627 ( .A(n9378), .B(n9379), .Z(n9377) );
  OR U11628 ( .A(n9380), .B(n9381), .Z(n9376) );
  NOR U11629 ( .A(n9382), .B(n9383), .Z(n9364) );
  ANDN U11630 ( .B(n9384), .A(n9385), .Z(n9358) );
  XNOR U11631 ( .A(n9351), .B(n9386), .Z(n9357) );
  XNOR U11632 ( .A(n9350), .B(n9352), .Z(n9386) );
  NAND U11633 ( .A(n9387), .B(n9388), .Z(n9352) );
  OR U11634 ( .A(n9389), .B(n9390), .Z(n9388) );
  OR U11635 ( .A(n9391), .B(n9392), .Z(n9387) );
  NAND U11636 ( .A(n9393), .B(n9394), .Z(n9350) );
  OR U11637 ( .A(n9395), .B(n9396), .Z(n9394) );
  OR U11638 ( .A(n9397), .B(n9398), .Z(n9393) );
  ANDN U11639 ( .B(n9399), .A(n9400), .Z(n9351) );
  IV U11640 ( .A(n9401), .Z(n9399) );
  ANDN U11641 ( .B(n9402), .A(n9403), .Z(n9343) );
  XOR U11642 ( .A(n9329), .B(n9404), .Z(n9341) );
  XOR U11643 ( .A(n9330), .B(n9331), .Z(n9404) );
  XOR U11644 ( .A(n9336), .B(n9405), .Z(n9331) );
  XOR U11645 ( .A(n9335), .B(n9338), .Z(n9405) );
  IV U11646 ( .A(n9337), .Z(n9338) );
  NAND U11647 ( .A(n9406), .B(n9407), .Z(n9337) );
  OR U11648 ( .A(n9408), .B(n9409), .Z(n9407) );
  OR U11649 ( .A(n9410), .B(n9411), .Z(n9406) );
  NAND U11650 ( .A(n9412), .B(n9413), .Z(n9335) );
  OR U11651 ( .A(n9414), .B(n9415), .Z(n9413) );
  OR U11652 ( .A(n9416), .B(n9417), .Z(n9412) );
  NOR U11653 ( .A(n9418), .B(n9419), .Z(n9336) );
  ANDN U11654 ( .B(n9420), .A(n9421), .Z(n9330) );
  IV U11655 ( .A(n9422), .Z(n9420) );
  XNOR U11656 ( .A(n9323), .B(n9423), .Z(n9329) );
  XNOR U11657 ( .A(n9322), .B(n9324), .Z(n9423) );
  NAND U11658 ( .A(n9424), .B(n9425), .Z(n9324) );
  OR U11659 ( .A(n9426), .B(n9427), .Z(n9425) );
  OR U11660 ( .A(n9428), .B(n9429), .Z(n9424) );
  NAND U11661 ( .A(n9430), .B(n9431), .Z(n9322) );
  OR U11662 ( .A(n9432), .B(n9433), .Z(n9431) );
  OR U11663 ( .A(n9434), .B(n9435), .Z(n9430) );
  ANDN U11664 ( .B(n9436), .A(n9437), .Z(n9323) );
  IV U11665 ( .A(n9438), .Z(n9436) );
  XNOR U11666 ( .A(n9403), .B(n9402), .Z(N13089) );
  XOR U11667 ( .A(n9422), .B(n9421), .Z(n9402) );
  XNOR U11668 ( .A(n9437), .B(n9438), .Z(n9421) );
  XNOR U11669 ( .A(n9432), .B(n9433), .Z(n9438) );
  XNOR U11670 ( .A(n9434), .B(n9435), .Z(n9433) );
  XNOR U11671 ( .A(y[685]), .B(x[685]), .Z(n9435) );
  XNOR U11672 ( .A(y[686]), .B(x[686]), .Z(n9434) );
  XNOR U11673 ( .A(y[684]), .B(x[684]), .Z(n9432) );
  XNOR U11674 ( .A(n9426), .B(n9427), .Z(n9437) );
  XNOR U11675 ( .A(y[681]), .B(x[681]), .Z(n9427) );
  XNOR U11676 ( .A(n9428), .B(n9429), .Z(n9426) );
  XNOR U11677 ( .A(y[682]), .B(x[682]), .Z(n9429) );
  XNOR U11678 ( .A(y[683]), .B(x[683]), .Z(n9428) );
  XNOR U11679 ( .A(n9419), .B(n9418), .Z(n9422) );
  XNOR U11680 ( .A(n9414), .B(n9415), .Z(n9418) );
  XNOR U11681 ( .A(y[678]), .B(x[678]), .Z(n9415) );
  XNOR U11682 ( .A(n9416), .B(n9417), .Z(n9414) );
  XNOR U11683 ( .A(y[679]), .B(x[679]), .Z(n9417) );
  XNOR U11684 ( .A(y[680]), .B(x[680]), .Z(n9416) );
  XNOR U11685 ( .A(n9408), .B(n9409), .Z(n9419) );
  XNOR U11686 ( .A(y[675]), .B(x[675]), .Z(n9409) );
  XNOR U11687 ( .A(n9410), .B(n9411), .Z(n9408) );
  XNOR U11688 ( .A(y[676]), .B(x[676]), .Z(n9411) );
  XNOR U11689 ( .A(y[677]), .B(x[677]), .Z(n9410) );
  XOR U11690 ( .A(n9384), .B(n9385), .Z(n9403) );
  XNOR U11691 ( .A(n9400), .B(n9401), .Z(n9385) );
  XNOR U11692 ( .A(n9395), .B(n9396), .Z(n9401) );
  XNOR U11693 ( .A(n9397), .B(n9398), .Z(n9396) );
  XNOR U11694 ( .A(y[673]), .B(x[673]), .Z(n9398) );
  XNOR U11695 ( .A(y[674]), .B(x[674]), .Z(n9397) );
  XNOR U11696 ( .A(y[672]), .B(x[672]), .Z(n9395) );
  XNOR U11697 ( .A(n9389), .B(n9390), .Z(n9400) );
  XNOR U11698 ( .A(y[669]), .B(x[669]), .Z(n9390) );
  XNOR U11699 ( .A(n9391), .B(n9392), .Z(n9389) );
  XNOR U11700 ( .A(y[670]), .B(x[670]), .Z(n9392) );
  XNOR U11701 ( .A(y[671]), .B(x[671]), .Z(n9391) );
  XOR U11702 ( .A(n9383), .B(n9382), .Z(n9384) );
  XNOR U11703 ( .A(n9378), .B(n9379), .Z(n9382) );
  XNOR U11704 ( .A(y[666]), .B(x[666]), .Z(n9379) );
  XNOR U11705 ( .A(n9380), .B(n9381), .Z(n9378) );
  XNOR U11706 ( .A(y[667]), .B(x[667]), .Z(n9381) );
  XNOR U11707 ( .A(y[668]), .B(x[668]), .Z(n9380) );
  XNOR U11708 ( .A(n9372), .B(n9373), .Z(n9383) );
  XNOR U11709 ( .A(y[663]), .B(x[663]), .Z(n9373) );
  XNOR U11710 ( .A(n9374), .B(n9375), .Z(n9372) );
  XNOR U11711 ( .A(y[664]), .B(x[664]), .Z(n9375) );
  XNOR U11712 ( .A(y[665]), .B(x[665]), .Z(n9374) );
  NAND U11713 ( .A(n9439), .B(n9440), .Z(N13082) );
  NANDN U11714 ( .A(n9441), .B(n9442), .Z(n9440) );
  OR U11715 ( .A(n9443), .B(n9444), .Z(n9442) );
  NAND U11716 ( .A(n9443), .B(n9444), .Z(n9439) );
  XOR U11717 ( .A(n9443), .B(n9445), .Z(N13081) );
  XNOR U11718 ( .A(n9441), .B(n9444), .Z(n9445) );
  AND U11719 ( .A(n9446), .B(n9447), .Z(n9444) );
  NANDN U11720 ( .A(n9448), .B(n9449), .Z(n9447) );
  NANDN U11721 ( .A(n9450), .B(n9451), .Z(n9449) );
  NANDN U11722 ( .A(n9451), .B(n9450), .Z(n9446) );
  NAND U11723 ( .A(n9452), .B(n9453), .Z(n9441) );
  NANDN U11724 ( .A(n9454), .B(n9455), .Z(n9453) );
  OR U11725 ( .A(n9456), .B(n9457), .Z(n9455) );
  NAND U11726 ( .A(n9457), .B(n9456), .Z(n9452) );
  AND U11727 ( .A(n9458), .B(n9459), .Z(n9443) );
  NANDN U11728 ( .A(n9460), .B(n9461), .Z(n9459) );
  NANDN U11729 ( .A(n9462), .B(n9463), .Z(n9461) );
  NANDN U11730 ( .A(n9463), .B(n9462), .Z(n9458) );
  XOR U11731 ( .A(n9457), .B(n9464), .Z(N13080) );
  XOR U11732 ( .A(n9454), .B(n9456), .Z(n9464) );
  XNOR U11733 ( .A(n9450), .B(n9465), .Z(n9456) );
  XNOR U11734 ( .A(n9448), .B(n9451), .Z(n9465) );
  NAND U11735 ( .A(n9466), .B(n9467), .Z(n9451) );
  NAND U11736 ( .A(n9468), .B(n9469), .Z(n9467) );
  OR U11737 ( .A(n9470), .B(n9471), .Z(n9468) );
  NANDN U11738 ( .A(n9472), .B(n9470), .Z(n9466) );
  IV U11739 ( .A(n9471), .Z(n9472) );
  NAND U11740 ( .A(n9473), .B(n9474), .Z(n9448) );
  NAND U11741 ( .A(n9475), .B(n9476), .Z(n9474) );
  NANDN U11742 ( .A(n9477), .B(n9478), .Z(n9475) );
  NANDN U11743 ( .A(n9478), .B(n9477), .Z(n9473) );
  AND U11744 ( .A(n9479), .B(n9480), .Z(n9450) );
  NAND U11745 ( .A(n9481), .B(n9482), .Z(n9480) );
  OR U11746 ( .A(n9483), .B(n9484), .Z(n9481) );
  NANDN U11747 ( .A(n9485), .B(n9483), .Z(n9479) );
  NAND U11748 ( .A(n9486), .B(n9487), .Z(n9454) );
  NANDN U11749 ( .A(n9488), .B(n9489), .Z(n9487) );
  OR U11750 ( .A(n9490), .B(n9491), .Z(n9489) );
  NANDN U11751 ( .A(n9492), .B(n9490), .Z(n9486) );
  IV U11752 ( .A(n9491), .Z(n9492) );
  XNOR U11753 ( .A(n9462), .B(n9493), .Z(n9457) );
  XNOR U11754 ( .A(n9460), .B(n9463), .Z(n9493) );
  NAND U11755 ( .A(n9494), .B(n9495), .Z(n9463) );
  NAND U11756 ( .A(n9496), .B(n9497), .Z(n9495) );
  OR U11757 ( .A(n9498), .B(n9499), .Z(n9496) );
  NANDN U11758 ( .A(n9500), .B(n9498), .Z(n9494) );
  IV U11759 ( .A(n9499), .Z(n9500) );
  NAND U11760 ( .A(n9501), .B(n9502), .Z(n9460) );
  NAND U11761 ( .A(n9503), .B(n9504), .Z(n9502) );
  NANDN U11762 ( .A(n9505), .B(n9506), .Z(n9503) );
  NANDN U11763 ( .A(n9506), .B(n9505), .Z(n9501) );
  AND U11764 ( .A(n9507), .B(n9508), .Z(n9462) );
  NAND U11765 ( .A(n9509), .B(n9510), .Z(n9508) );
  OR U11766 ( .A(n9511), .B(n9512), .Z(n9509) );
  NANDN U11767 ( .A(n9513), .B(n9511), .Z(n9507) );
  XNOR U11768 ( .A(n9488), .B(n9514), .Z(N13079) );
  XOR U11769 ( .A(n9490), .B(n9491), .Z(n9514) );
  XNOR U11770 ( .A(n9504), .B(n9515), .Z(n9491) );
  XOR U11771 ( .A(n9505), .B(n9506), .Z(n9515) );
  XOR U11772 ( .A(n9511), .B(n9516), .Z(n9506) );
  XOR U11773 ( .A(n9510), .B(n9513), .Z(n9516) );
  IV U11774 ( .A(n9512), .Z(n9513) );
  NAND U11775 ( .A(n9517), .B(n9518), .Z(n9512) );
  OR U11776 ( .A(n9519), .B(n9520), .Z(n9518) );
  OR U11777 ( .A(n9521), .B(n9522), .Z(n9517) );
  NAND U11778 ( .A(n9523), .B(n9524), .Z(n9510) );
  OR U11779 ( .A(n9525), .B(n9526), .Z(n9524) );
  OR U11780 ( .A(n9527), .B(n9528), .Z(n9523) );
  NOR U11781 ( .A(n9529), .B(n9530), .Z(n9511) );
  ANDN U11782 ( .B(n9531), .A(n9532), .Z(n9505) );
  XNOR U11783 ( .A(n9498), .B(n9533), .Z(n9504) );
  XNOR U11784 ( .A(n9497), .B(n9499), .Z(n9533) );
  NAND U11785 ( .A(n9534), .B(n9535), .Z(n9499) );
  OR U11786 ( .A(n9536), .B(n9537), .Z(n9535) );
  OR U11787 ( .A(n9538), .B(n9539), .Z(n9534) );
  NAND U11788 ( .A(n9540), .B(n9541), .Z(n9497) );
  OR U11789 ( .A(n9542), .B(n9543), .Z(n9541) );
  OR U11790 ( .A(n9544), .B(n9545), .Z(n9540) );
  ANDN U11791 ( .B(n9546), .A(n9547), .Z(n9498) );
  IV U11792 ( .A(n9548), .Z(n9546) );
  ANDN U11793 ( .B(n9549), .A(n9550), .Z(n9490) );
  XOR U11794 ( .A(n9476), .B(n9551), .Z(n9488) );
  XOR U11795 ( .A(n9477), .B(n9478), .Z(n9551) );
  XOR U11796 ( .A(n9483), .B(n9552), .Z(n9478) );
  XOR U11797 ( .A(n9482), .B(n9485), .Z(n9552) );
  IV U11798 ( .A(n9484), .Z(n9485) );
  NAND U11799 ( .A(n9553), .B(n9554), .Z(n9484) );
  OR U11800 ( .A(n9555), .B(n9556), .Z(n9554) );
  OR U11801 ( .A(n9557), .B(n9558), .Z(n9553) );
  NAND U11802 ( .A(n9559), .B(n9560), .Z(n9482) );
  OR U11803 ( .A(n9561), .B(n9562), .Z(n9560) );
  OR U11804 ( .A(n9563), .B(n9564), .Z(n9559) );
  NOR U11805 ( .A(n9565), .B(n9566), .Z(n9483) );
  ANDN U11806 ( .B(n9567), .A(n9568), .Z(n9477) );
  IV U11807 ( .A(n9569), .Z(n9567) );
  XNOR U11808 ( .A(n9470), .B(n9570), .Z(n9476) );
  XNOR U11809 ( .A(n9469), .B(n9471), .Z(n9570) );
  NAND U11810 ( .A(n9571), .B(n9572), .Z(n9471) );
  OR U11811 ( .A(n9573), .B(n9574), .Z(n9572) );
  OR U11812 ( .A(n9575), .B(n9576), .Z(n9571) );
  NAND U11813 ( .A(n9577), .B(n9578), .Z(n9469) );
  OR U11814 ( .A(n9579), .B(n9580), .Z(n9578) );
  OR U11815 ( .A(n9581), .B(n9582), .Z(n9577) );
  ANDN U11816 ( .B(n9583), .A(n9584), .Z(n9470) );
  IV U11817 ( .A(n9585), .Z(n9583) );
  XNOR U11818 ( .A(n9550), .B(n9549), .Z(N13078) );
  XOR U11819 ( .A(n9569), .B(n9568), .Z(n9549) );
  XNOR U11820 ( .A(n9584), .B(n9585), .Z(n9568) );
  XNOR U11821 ( .A(n9579), .B(n9580), .Z(n9585) );
  XNOR U11822 ( .A(n9581), .B(n9582), .Z(n9580) );
  XNOR U11823 ( .A(y[661]), .B(x[661]), .Z(n9582) );
  XNOR U11824 ( .A(y[662]), .B(x[662]), .Z(n9581) );
  XNOR U11825 ( .A(y[660]), .B(x[660]), .Z(n9579) );
  XNOR U11826 ( .A(n9573), .B(n9574), .Z(n9584) );
  XNOR U11827 ( .A(y[657]), .B(x[657]), .Z(n9574) );
  XNOR U11828 ( .A(n9575), .B(n9576), .Z(n9573) );
  XNOR U11829 ( .A(y[658]), .B(x[658]), .Z(n9576) );
  XNOR U11830 ( .A(y[659]), .B(x[659]), .Z(n9575) );
  XNOR U11831 ( .A(n9566), .B(n9565), .Z(n9569) );
  XNOR U11832 ( .A(n9561), .B(n9562), .Z(n9565) );
  XNOR U11833 ( .A(y[654]), .B(x[654]), .Z(n9562) );
  XNOR U11834 ( .A(n9563), .B(n9564), .Z(n9561) );
  XNOR U11835 ( .A(y[655]), .B(x[655]), .Z(n9564) );
  XNOR U11836 ( .A(y[656]), .B(x[656]), .Z(n9563) );
  XNOR U11837 ( .A(n9555), .B(n9556), .Z(n9566) );
  XNOR U11838 ( .A(y[651]), .B(x[651]), .Z(n9556) );
  XNOR U11839 ( .A(n9557), .B(n9558), .Z(n9555) );
  XNOR U11840 ( .A(y[652]), .B(x[652]), .Z(n9558) );
  XNOR U11841 ( .A(y[653]), .B(x[653]), .Z(n9557) );
  XOR U11842 ( .A(n9531), .B(n9532), .Z(n9550) );
  XNOR U11843 ( .A(n9547), .B(n9548), .Z(n9532) );
  XNOR U11844 ( .A(n9542), .B(n9543), .Z(n9548) );
  XNOR U11845 ( .A(n9544), .B(n9545), .Z(n9543) );
  XNOR U11846 ( .A(y[649]), .B(x[649]), .Z(n9545) );
  XNOR U11847 ( .A(y[650]), .B(x[650]), .Z(n9544) );
  XNOR U11848 ( .A(y[648]), .B(x[648]), .Z(n9542) );
  XNOR U11849 ( .A(n9536), .B(n9537), .Z(n9547) );
  XNOR U11850 ( .A(y[645]), .B(x[645]), .Z(n9537) );
  XNOR U11851 ( .A(n9538), .B(n9539), .Z(n9536) );
  XNOR U11852 ( .A(y[646]), .B(x[646]), .Z(n9539) );
  XNOR U11853 ( .A(y[647]), .B(x[647]), .Z(n9538) );
  XOR U11854 ( .A(n9530), .B(n9529), .Z(n9531) );
  XNOR U11855 ( .A(n9525), .B(n9526), .Z(n9529) );
  XNOR U11856 ( .A(y[642]), .B(x[642]), .Z(n9526) );
  XNOR U11857 ( .A(n9527), .B(n9528), .Z(n9525) );
  XNOR U11858 ( .A(y[643]), .B(x[643]), .Z(n9528) );
  XNOR U11859 ( .A(y[644]), .B(x[644]), .Z(n9527) );
  XNOR U11860 ( .A(n9519), .B(n9520), .Z(n9530) );
  XNOR U11861 ( .A(y[639]), .B(x[639]), .Z(n9520) );
  XNOR U11862 ( .A(n9521), .B(n9522), .Z(n9519) );
  XNOR U11863 ( .A(y[640]), .B(x[640]), .Z(n9522) );
  XNOR U11864 ( .A(y[641]), .B(x[641]), .Z(n9521) );
  NAND U11865 ( .A(n9586), .B(n9587), .Z(N13071) );
  NANDN U11866 ( .A(n9588), .B(n9589), .Z(n9587) );
  OR U11867 ( .A(n9590), .B(n9591), .Z(n9589) );
  NAND U11868 ( .A(n9590), .B(n9591), .Z(n9586) );
  XOR U11869 ( .A(n9590), .B(n9592), .Z(N13070) );
  XNOR U11870 ( .A(n9588), .B(n9591), .Z(n9592) );
  AND U11871 ( .A(n9593), .B(n9594), .Z(n9591) );
  NANDN U11872 ( .A(n9595), .B(n9596), .Z(n9594) );
  NANDN U11873 ( .A(n9597), .B(n9598), .Z(n9596) );
  NANDN U11874 ( .A(n9598), .B(n9597), .Z(n9593) );
  NAND U11875 ( .A(n9599), .B(n9600), .Z(n9588) );
  NANDN U11876 ( .A(n9601), .B(n9602), .Z(n9600) );
  OR U11877 ( .A(n9603), .B(n9604), .Z(n9602) );
  NAND U11878 ( .A(n9604), .B(n9603), .Z(n9599) );
  AND U11879 ( .A(n9605), .B(n9606), .Z(n9590) );
  NANDN U11880 ( .A(n9607), .B(n9608), .Z(n9606) );
  NANDN U11881 ( .A(n9609), .B(n9610), .Z(n9608) );
  NANDN U11882 ( .A(n9610), .B(n9609), .Z(n9605) );
  XOR U11883 ( .A(n9604), .B(n9611), .Z(N13069) );
  XOR U11884 ( .A(n9601), .B(n9603), .Z(n9611) );
  XNOR U11885 ( .A(n9597), .B(n9612), .Z(n9603) );
  XNOR U11886 ( .A(n9595), .B(n9598), .Z(n9612) );
  NAND U11887 ( .A(n9613), .B(n9614), .Z(n9598) );
  NAND U11888 ( .A(n9615), .B(n9616), .Z(n9614) );
  OR U11889 ( .A(n9617), .B(n9618), .Z(n9615) );
  NANDN U11890 ( .A(n9619), .B(n9617), .Z(n9613) );
  IV U11891 ( .A(n9618), .Z(n9619) );
  NAND U11892 ( .A(n9620), .B(n9621), .Z(n9595) );
  NAND U11893 ( .A(n9622), .B(n9623), .Z(n9621) );
  NANDN U11894 ( .A(n9624), .B(n9625), .Z(n9622) );
  NANDN U11895 ( .A(n9625), .B(n9624), .Z(n9620) );
  AND U11896 ( .A(n9626), .B(n9627), .Z(n9597) );
  NAND U11897 ( .A(n9628), .B(n9629), .Z(n9627) );
  OR U11898 ( .A(n9630), .B(n9631), .Z(n9628) );
  NANDN U11899 ( .A(n9632), .B(n9630), .Z(n9626) );
  NAND U11900 ( .A(n9633), .B(n9634), .Z(n9601) );
  NANDN U11901 ( .A(n9635), .B(n9636), .Z(n9634) );
  OR U11902 ( .A(n9637), .B(n9638), .Z(n9636) );
  NANDN U11903 ( .A(n9639), .B(n9637), .Z(n9633) );
  IV U11904 ( .A(n9638), .Z(n9639) );
  XNOR U11905 ( .A(n9609), .B(n9640), .Z(n9604) );
  XNOR U11906 ( .A(n9607), .B(n9610), .Z(n9640) );
  NAND U11907 ( .A(n9641), .B(n9642), .Z(n9610) );
  NAND U11908 ( .A(n9643), .B(n9644), .Z(n9642) );
  OR U11909 ( .A(n9645), .B(n9646), .Z(n9643) );
  NANDN U11910 ( .A(n9647), .B(n9645), .Z(n9641) );
  IV U11911 ( .A(n9646), .Z(n9647) );
  NAND U11912 ( .A(n9648), .B(n9649), .Z(n9607) );
  NAND U11913 ( .A(n9650), .B(n9651), .Z(n9649) );
  NANDN U11914 ( .A(n9652), .B(n9653), .Z(n9650) );
  NANDN U11915 ( .A(n9653), .B(n9652), .Z(n9648) );
  AND U11916 ( .A(n9654), .B(n9655), .Z(n9609) );
  NAND U11917 ( .A(n9656), .B(n9657), .Z(n9655) );
  OR U11918 ( .A(n9658), .B(n9659), .Z(n9656) );
  NANDN U11919 ( .A(n9660), .B(n9658), .Z(n9654) );
  XNOR U11920 ( .A(n9635), .B(n9661), .Z(N13068) );
  XOR U11921 ( .A(n9637), .B(n9638), .Z(n9661) );
  XNOR U11922 ( .A(n9651), .B(n9662), .Z(n9638) );
  XOR U11923 ( .A(n9652), .B(n9653), .Z(n9662) );
  XOR U11924 ( .A(n9658), .B(n9663), .Z(n9653) );
  XOR U11925 ( .A(n9657), .B(n9660), .Z(n9663) );
  IV U11926 ( .A(n9659), .Z(n9660) );
  NAND U11927 ( .A(n9664), .B(n9665), .Z(n9659) );
  OR U11928 ( .A(n9666), .B(n9667), .Z(n9665) );
  OR U11929 ( .A(n9668), .B(n9669), .Z(n9664) );
  NAND U11930 ( .A(n9670), .B(n9671), .Z(n9657) );
  OR U11931 ( .A(n9672), .B(n9673), .Z(n9671) );
  OR U11932 ( .A(n9674), .B(n9675), .Z(n9670) );
  NOR U11933 ( .A(n9676), .B(n9677), .Z(n9658) );
  ANDN U11934 ( .B(n9678), .A(n9679), .Z(n9652) );
  XNOR U11935 ( .A(n9645), .B(n9680), .Z(n9651) );
  XNOR U11936 ( .A(n9644), .B(n9646), .Z(n9680) );
  NAND U11937 ( .A(n9681), .B(n9682), .Z(n9646) );
  OR U11938 ( .A(n9683), .B(n9684), .Z(n9682) );
  OR U11939 ( .A(n9685), .B(n9686), .Z(n9681) );
  NAND U11940 ( .A(n9687), .B(n9688), .Z(n9644) );
  OR U11941 ( .A(n9689), .B(n9690), .Z(n9688) );
  OR U11942 ( .A(n9691), .B(n9692), .Z(n9687) );
  ANDN U11943 ( .B(n9693), .A(n9694), .Z(n9645) );
  IV U11944 ( .A(n9695), .Z(n9693) );
  ANDN U11945 ( .B(n9696), .A(n9697), .Z(n9637) );
  XOR U11946 ( .A(n9623), .B(n9698), .Z(n9635) );
  XOR U11947 ( .A(n9624), .B(n9625), .Z(n9698) );
  XOR U11948 ( .A(n9630), .B(n9699), .Z(n9625) );
  XOR U11949 ( .A(n9629), .B(n9632), .Z(n9699) );
  IV U11950 ( .A(n9631), .Z(n9632) );
  NAND U11951 ( .A(n9700), .B(n9701), .Z(n9631) );
  OR U11952 ( .A(n9702), .B(n9703), .Z(n9701) );
  OR U11953 ( .A(n9704), .B(n9705), .Z(n9700) );
  NAND U11954 ( .A(n9706), .B(n9707), .Z(n9629) );
  OR U11955 ( .A(n9708), .B(n9709), .Z(n9707) );
  OR U11956 ( .A(n9710), .B(n9711), .Z(n9706) );
  NOR U11957 ( .A(n9712), .B(n9713), .Z(n9630) );
  ANDN U11958 ( .B(n9714), .A(n9715), .Z(n9624) );
  IV U11959 ( .A(n9716), .Z(n9714) );
  XNOR U11960 ( .A(n9617), .B(n9717), .Z(n9623) );
  XNOR U11961 ( .A(n9616), .B(n9618), .Z(n9717) );
  NAND U11962 ( .A(n9718), .B(n9719), .Z(n9618) );
  OR U11963 ( .A(n9720), .B(n9721), .Z(n9719) );
  OR U11964 ( .A(n9722), .B(n9723), .Z(n9718) );
  NAND U11965 ( .A(n9724), .B(n9725), .Z(n9616) );
  OR U11966 ( .A(n9726), .B(n9727), .Z(n9725) );
  OR U11967 ( .A(n9728), .B(n9729), .Z(n9724) );
  ANDN U11968 ( .B(n9730), .A(n9731), .Z(n9617) );
  IV U11969 ( .A(n9732), .Z(n9730) );
  XNOR U11970 ( .A(n9697), .B(n9696), .Z(N13067) );
  XOR U11971 ( .A(n9716), .B(n9715), .Z(n9696) );
  XNOR U11972 ( .A(n9731), .B(n9732), .Z(n9715) );
  XNOR U11973 ( .A(n9726), .B(n9727), .Z(n9732) );
  XNOR U11974 ( .A(n9728), .B(n9729), .Z(n9727) );
  XNOR U11975 ( .A(y[637]), .B(x[637]), .Z(n9729) );
  XNOR U11976 ( .A(y[638]), .B(x[638]), .Z(n9728) );
  XNOR U11977 ( .A(y[636]), .B(x[636]), .Z(n9726) );
  XNOR U11978 ( .A(n9720), .B(n9721), .Z(n9731) );
  XNOR U11979 ( .A(y[633]), .B(x[633]), .Z(n9721) );
  XNOR U11980 ( .A(n9722), .B(n9723), .Z(n9720) );
  XNOR U11981 ( .A(y[634]), .B(x[634]), .Z(n9723) );
  XNOR U11982 ( .A(y[635]), .B(x[635]), .Z(n9722) );
  XNOR U11983 ( .A(n9713), .B(n9712), .Z(n9716) );
  XNOR U11984 ( .A(n9708), .B(n9709), .Z(n9712) );
  XNOR U11985 ( .A(y[630]), .B(x[630]), .Z(n9709) );
  XNOR U11986 ( .A(n9710), .B(n9711), .Z(n9708) );
  XNOR U11987 ( .A(y[631]), .B(x[631]), .Z(n9711) );
  XNOR U11988 ( .A(y[632]), .B(x[632]), .Z(n9710) );
  XNOR U11989 ( .A(n9702), .B(n9703), .Z(n9713) );
  XNOR U11990 ( .A(y[627]), .B(x[627]), .Z(n9703) );
  XNOR U11991 ( .A(n9704), .B(n9705), .Z(n9702) );
  XNOR U11992 ( .A(y[628]), .B(x[628]), .Z(n9705) );
  XNOR U11993 ( .A(y[629]), .B(x[629]), .Z(n9704) );
  XOR U11994 ( .A(n9678), .B(n9679), .Z(n9697) );
  XNOR U11995 ( .A(n9694), .B(n9695), .Z(n9679) );
  XNOR U11996 ( .A(n9689), .B(n9690), .Z(n9695) );
  XNOR U11997 ( .A(n9691), .B(n9692), .Z(n9690) );
  XNOR U11998 ( .A(y[625]), .B(x[625]), .Z(n9692) );
  XNOR U11999 ( .A(y[626]), .B(x[626]), .Z(n9691) );
  XNOR U12000 ( .A(y[624]), .B(x[624]), .Z(n9689) );
  XNOR U12001 ( .A(n9683), .B(n9684), .Z(n9694) );
  XNOR U12002 ( .A(y[621]), .B(x[621]), .Z(n9684) );
  XNOR U12003 ( .A(n9685), .B(n9686), .Z(n9683) );
  XNOR U12004 ( .A(y[622]), .B(x[622]), .Z(n9686) );
  XNOR U12005 ( .A(y[623]), .B(x[623]), .Z(n9685) );
  XOR U12006 ( .A(n9677), .B(n9676), .Z(n9678) );
  XNOR U12007 ( .A(n9672), .B(n9673), .Z(n9676) );
  XNOR U12008 ( .A(y[618]), .B(x[618]), .Z(n9673) );
  XNOR U12009 ( .A(n9674), .B(n9675), .Z(n9672) );
  XNOR U12010 ( .A(y[619]), .B(x[619]), .Z(n9675) );
  XNOR U12011 ( .A(y[620]), .B(x[620]), .Z(n9674) );
  XNOR U12012 ( .A(n9666), .B(n9667), .Z(n9677) );
  XNOR U12013 ( .A(y[615]), .B(x[615]), .Z(n9667) );
  XNOR U12014 ( .A(n9668), .B(n9669), .Z(n9666) );
  XNOR U12015 ( .A(y[616]), .B(x[616]), .Z(n9669) );
  XNOR U12016 ( .A(y[617]), .B(x[617]), .Z(n9668) );
  NAND U12017 ( .A(n9733), .B(n9734), .Z(N13060) );
  NANDN U12018 ( .A(n9735), .B(n9736), .Z(n9734) );
  OR U12019 ( .A(n9737), .B(n9738), .Z(n9736) );
  NAND U12020 ( .A(n9737), .B(n9738), .Z(n9733) );
  XOR U12021 ( .A(n9737), .B(n9739), .Z(N13059) );
  XNOR U12022 ( .A(n9735), .B(n9738), .Z(n9739) );
  AND U12023 ( .A(n9740), .B(n9741), .Z(n9738) );
  NANDN U12024 ( .A(n9742), .B(n9743), .Z(n9741) );
  NANDN U12025 ( .A(n9744), .B(n9745), .Z(n9743) );
  NANDN U12026 ( .A(n9745), .B(n9744), .Z(n9740) );
  NAND U12027 ( .A(n9746), .B(n9747), .Z(n9735) );
  NANDN U12028 ( .A(n9748), .B(n9749), .Z(n9747) );
  OR U12029 ( .A(n9750), .B(n9751), .Z(n9749) );
  NAND U12030 ( .A(n9751), .B(n9750), .Z(n9746) );
  AND U12031 ( .A(n9752), .B(n9753), .Z(n9737) );
  NANDN U12032 ( .A(n9754), .B(n9755), .Z(n9753) );
  NANDN U12033 ( .A(n9756), .B(n9757), .Z(n9755) );
  NANDN U12034 ( .A(n9757), .B(n9756), .Z(n9752) );
  XOR U12035 ( .A(n9751), .B(n9758), .Z(N13058) );
  XOR U12036 ( .A(n9748), .B(n9750), .Z(n9758) );
  XNOR U12037 ( .A(n9744), .B(n9759), .Z(n9750) );
  XNOR U12038 ( .A(n9742), .B(n9745), .Z(n9759) );
  NAND U12039 ( .A(n9760), .B(n9761), .Z(n9745) );
  NAND U12040 ( .A(n9762), .B(n9763), .Z(n9761) );
  OR U12041 ( .A(n9764), .B(n9765), .Z(n9762) );
  NANDN U12042 ( .A(n9766), .B(n9764), .Z(n9760) );
  IV U12043 ( .A(n9765), .Z(n9766) );
  NAND U12044 ( .A(n9767), .B(n9768), .Z(n9742) );
  NAND U12045 ( .A(n9769), .B(n9770), .Z(n9768) );
  NANDN U12046 ( .A(n9771), .B(n9772), .Z(n9769) );
  NANDN U12047 ( .A(n9772), .B(n9771), .Z(n9767) );
  AND U12048 ( .A(n9773), .B(n9774), .Z(n9744) );
  NAND U12049 ( .A(n9775), .B(n9776), .Z(n9774) );
  OR U12050 ( .A(n9777), .B(n9778), .Z(n9775) );
  NANDN U12051 ( .A(n9779), .B(n9777), .Z(n9773) );
  NAND U12052 ( .A(n9780), .B(n9781), .Z(n9748) );
  NANDN U12053 ( .A(n9782), .B(n9783), .Z(n9781) );
  OR U12054 ( .A(n9784), .B(n9785), .Z(n9783) );
  NANDN U12055 ( .A(n9786), .B(n9784), .Z(n9780) );
  IV U12056 ( .A(n9785), .Z(n9786) );
  XNOR U12057 ( .A(n9756), .B(n9787), .Z(n9751) );
  XNOR U12058 ( .A(n9754), .B(n9757), .Z(n9787) );
  NAND U12059 ( .A(n9788), .B(n9789), .Z(n9757) );
  NAND U12060 ( .A(n9790), .B(n9791), .Z(n9789) );
  OR U12061 ( .A(n9792), .B(n9793), .Z(n9790) );
  NANDN U12062 ( .A(n9794), .B(n9792), .Z(n9788) );
  IV U12063 ( .A(n9793), .Z(n9794) );
  NAND U12064 ( .A(n9795), .B(n9796), .Z(n9754) );
  NAND U12065 ( .A(n9797), .B(n9798), .Z(n9796) );
  NANDN U12066 ( .A(n9799), .B(n9800), .Z(n9797) );
  NANDN U12067 ( .A(n9800), .B(n9799), .Z(n9795) );
  AND U12068 ( .A(n9801), .B(n9802), .Z(n9756) );
  NAND U12069 ( .A(n9803), .B(n9804), .Z(n9802) );
  OR U12070 ( .A(n9805), .B(n9806), .Z(n9803) );
  NANDN U12071 ( .A(n9807), .B(n9805), .Z(n9801) );
  XNOR U12072 ( .A(n9782), .B(n9808), .Z(N13057) );
  XOR U12073 ( .A(n9784), .B(n9785), .Z(n9808) );
  XNOR U12074 ( .A(n9798), .B(n9809), .Z(n9785) );
  XOR U12075 ( .A(n9799), .B(n9800), .Z(n9809) );
  XOR U12076 ( .A(n9805), .B(n9810), .Z(n9800) );
  XOR U12077 ( .A(n9804), .B(n9807), .Z(n9810) );
  IV U12078 ( .A(n9806), .Z(n9807) );
  NAND U12079 ( .A(n9811), .B(n9812), .Z(n9806) );
  OR U12080 ( .A(n9813), .B(n9814), .Z(n9812) );
  OR U12081 ( .A(n9815), .B(n9816), .Z(n9811) );
  NAND U12082 ( .A(n9817), .B(n9818), .Z(n9804) );
  OR U12083 ( .A(n9819), .B(n9820), .Z(n9818) );
  OR U12084 ( .A(n9821), .B(n9822), .Z(n9817) );
  NOR U12085 ( .A(n9823), .B(n9824), .Z(n9805) );
  ANDN U12086 ( .B(n9825), .A(n9826), .Z(n9799) );
  XNOR U12087 ( .A(n9792), .B(n9827), .Z(n9798) );
  XNOR U12088 ( .A(n9791), .B(n9793), .Z(n9827) );
  NAND U12089 ( .A(n9828), .B(n9829), .Z(n9793) );
  OR U12090 ( .A(n9830), .B(n9831), .Z(n9829) );
  OR U12091 ( .A(n9832), .B(n9833), .Z(n9828) );
  NAND U12092 ( .A(n9834), .B(n9835), .Z(n9791) );
  OR U12093 ( .A(n9836), .B(n9837), .Z(n9835) );
  OR U12094 ( .A(n9838), .B(n9839), .Z(n9834) );
  ANDN U12095 ( .B(n9840), .A(n9841), .Z(n9792) );
  IV U12096 ( .A(n9842), .Z(n9840) );
  ANDN U12097 ( .B(n9843), .A(n9844), .Z(n9784) );
  XOR U12098 ( .A(n9770), .B(n9845), .Z(n9782) );
  XOR U12099 ( .A(n9771), .B(n9772), .Z(n9845) );
  XOR U12100 ( .A(n9777), .B(n9846), .Z(n9772) );
  XOR U12101 ( .A(n9776), .B(n9779), .Z(n9846) );
  IV U12102 ( .A(n9778), .Z(n9779) );
  NAND U12103 ( .A(n9847), .B(n9848), .Z(n9778) );
  OR U12104 ( .A(n9849), .B(n9850), .Z(n9848) );
  OR U12105 ( .A(n9851), .B(n9852), .Z(n9847) );
  NAND U12106 ( .A(n9853), .B(n9854), .Z(n9776) );
  OR U12107 ( .A(n9855), .B(n9856), .Z(n9854) );
  OR U12108 ( .A(n9857), .B(n9858), .Z(n9853) );
  NOR U12109 ( .A(n9859), .B(n9860), .Z(n9777) );
  ANDN U12110 ( .B(n9861), .A(n9862), .Z(n9771) );
  IV U12111 ( .A(n9863), .Z(n9861) );
  XNOR U12112 ( .A(n9764), .B(n9864), .Z(n9770) );
  XNOR U12113 ( .A(n9763), .B(n9765), .Z(n9864) );
  NAND U12114 ( .A(n9865), .B(n9866), .Z(n9765) );
  OR U12115 ( .A(n9867), .B(n9868), .Z(n9866) );
  OR U12116 ( .A(n9869), .B(n9870), .Z(n9865) );
  NAND U12117 ( .A(n9871), .B(n9872), .Z(n9763) );
  OR U12118 ( .A(n9873), .B(n9874), .Z(n9872) );
  OR U12119 ( .A(n9875), .B(n9876), .Z(n9871) );
  ANDN U12120 ( .B(n9877), .A(n9878), .Z(n9764) );
  IV U12121 ( .A(n9879), .Z(n9877) );
  XNOR U12122 ( .A(n9844), .B(n9843), .Z(N13056) );
  XOR U12123 ( .A(n9863), .B(n9862), .Z(n9843) );
  XNOR U12124 ( .A(n9878), .B(n9879), .Z(n9862) );
  XNOR U12125 ( .A(n9873), .B(n9874), .Z(n9879) );
  XNOR U12126 ( .A(n9875), .B(n9876), .Z(n9874) );
  XNOR U12127 ( .A(y[613]), .B(x[613]), .Z(n9876) );
  XNOR U12128 ( .A(y[614]), .B(x[614]), .Z(n9875) );
  XNOR U12129 ( .A(y[612]), .B(x[612]), .Z(n9873) );
  XNOR U12130 ( .A(n9867), .B(n9868), .Z(n9878) );
  XNOR U12131 ( .A(y[609]), .B(x[609]), .Z(n9868) );
  XNOR U12132 ( .A(n9869), .B(n9870), .Z(n9867) );
  XNOR U12133 ( .A(y[610]), .B(x[610]), .Z(n9870) );
  XNOR U12134 ( .A(y[611]), .B(x[611]), .Z(n9869) );
  XNOR U12135 ( .A(n9860), .B(n9859), .Z(n9863) );
  XNOR U12136 ( .A(n9855), .B(n9856), .Z(n9859) );
  XNOR U12137 ( .A(y[606]), .B(x[606]), .Z(n9856) );
  XNOR U12138 ( .A(n9857), .B(n9858), .Z(n9855) );
  XNOR U12139 ( .A(y[607]), .B(x[607]), .Z(n9858) );
  XNOR U12140 ( .A(y[608]), .B(x[608]), .Z(n9857) );
  XNOR U12141 ( .A(n9849), .B(n9850), .Z(n9860) );
  XNOR U12142 ( .A(y[603]), .B(x[603]), .Z(n9850) );
  XNOR U12143 ( .A(n9851), .B(n9852), .Z(n9849) );
  XNOR U12144 ( .A(y[604]), .B(x[604]), .Z(n9852) );
  XNOR U12145 ( .A(y[605]), .B(x[605]), .Z(n9851) );
  XOR U12146 ( .A(n9825), .B(n9826), .Z(n9844) );
  XNOR U12147 ( .A(n9841), .B(n9842), .Z(n9826) );
  XNOR U12148 ( .A(n9836), .B(n9837), .Z(n9842) );
  XNOR U12149 ( .A(n9838), .B(n9839), .Z(n9837) );
  XNOR U12150 ( .A(y[601]), .B(x[601]), .Z(n9839) );
  XNOR U12151 ( .A(y[602]), .B(x[602]), .Z(n9838) );
  XNOR U12152 ( .A(y[600]), .B(x[600]), .Z(n9836) );
  XNOR U12153 ( .A(n9830), .B(n9831), .Z(n9841) );
  XNOR U12154 ( .A(y[597]), .B(x[597]), .Z(n9831) );
  XNOR U12155 ( .A(n9832), .B(n9833), .Z(n9830) );
  XNOR U12156 ( .A(y[598]), .B(x[598]), .Z(n9833) );
  XNOR U12157 ( .A(y[599]), .B(x[599]), .Z(n9832) );
  XOR U12158 ( .A(n9824), .B(n9823), .Z(n9825) );
  XNOR U12159 ( .A(n9819), .B(n9820), .Z(n9823) );
  XNOR U12160 ( .A(y[594]), .B(x[594]), .Z(n9820) );
  XNOR U12161 ( .A(n9821), .B(n9822), .Z(n9819) );
  XNOR U12162 ( .A(y[595]), .B(x[595]), .Z(n9822) );
  XNOR U12163 ( .A(y[596]), .B(x[596]), .Z(n9821) );
  XNOR U12164 ( .A(n9813), .B(n9814), .Z(n9824) );
  XNOR U12165 ( .A(y[591]), .B(x[591]), .Z(n9814) );
  XNOR U12166 ( .A(n9815), .B(n9816), .Z(n9813) );
  XNOR U12167 ( .A(y[592]), .B(x[592]), .Z(n9816) );
  XNOR U12168 ( .A(y[593]), .B(x[593]), .Z(n9815) );
  NAND U12169 ( .A(n9880), .B(n9881), .Z(N13049) );
  NANDN U12170 ( .A(n9882), .B(n9883), .Z(n9881) );
  OR U12171 ( .A(n9884), .B(n9885), .Z(n9883) );
  NAND U12172 ( .A(n9884), .B(n9885), .Z(n9880) );
  XOR U12173 ( .A(n9884), .B(n9886), .Z(N13048) );
  XNOR U12174 ( .A(n9882), .B(n9885), .Z(n9886) );
  AND U12175 ( .A(n9887), .B(n9888), .Z(n9885) );
  NANDN U12176 ( .A(n9889), .B(n9890), .Z(n9888) );
  NANDN U12177 ( .A(n9891), .B(n9892), .Z(n9890) );
  NANDN U12178 ( .A(n9892), .B(n9891), .Z(n9887) );
  NAND U12179 ( .A(n9893), .B(n9894), .Z(n9882) );
  NANDN U12180 ( .A(n9895), .B(n9896), .Z(n9894) );
  OR U12181 ( .A(n9897), .B(n9898), .Z(n9896) );
  NAND U12182 ( .A(n9898), .B(n9897), .Z(n9893) );
  AND U12183 ( .A(n9899), .B(n9900), .Z(n9884) );
  NANDN U12184 ( .A(n9901), .B(n9902), .Z(n9900) );
  NANDN U12185 ( .A(n9903), .B(n9904), .Z(n9902) );
  NANDN U12186 ( .A(n9904), .B(n9903), .Z(n9899) );
  XOR U12187 ( .A(n9898), .B(n9905), .Z(N13047) );
  XOR U12188 ( .A(n9895), .B(n9897), .Z(n9905) );
  XNOR U12189 ( .A(n9891), .B(n9906), .Z(n9897) );
  XNOR U12190 ( .A(n9889), .B(n9892), .Z(n9906) );
  NAND U12191 ( .A(n9907), .B(n9908), .Z(n9892) );
  NAND U12192 ( .A(n9909), .B(n9910), .Z(n9908) );
  OR U12193 ( .A(n9911), .B(n9912), .Z(n9909) );
  NANDN U12194 ( .A(n9913), .B(n9911), .Z(n9907) );
  IV U12195 ( .A(n9912), .Z(n9913) );
  NAND U12196 ( .A(n9914), .B(n9915), .Z(n9889) );
  NAND U12197 ( .A(n9916), .B(n9917), .Z(n9915) );
  NANDN U12198 ( .A(n9918), .B(n9919), .Z(n9916) );
  NANDN U12199 ( .A(n9919), .B(n9918), .Z(n9914) );
  AND U12200 ( .A(n9920), .B(n9921), .Z(n9891) );
  NAND U12201 ( .A(n9922), .B(n9923), .Z(n9921) );
  OR U12202 ( .A(n9924), .B(n9925), .Z(n9922) );
  NANDN U12203 ( .A(n9926), .B(n9924), .Z(n9920) );
  NAND U12204 ( .A(n9927), .B(n9928), .Z(n9895) );
  NANDN U12205 ( .A(n9929), .B(n9930), .Z(n9928) );
  OR U12206 ( .A(n9931), .B(n9932), .Z(n9930) );
  NANDN U12207 ( .A(n9933), .B(n9931), .Z(n9927) );
  IV U12208 ( .A(n9932), .Z(n9933) );
  XNOR U12209 ( .A(n9903), .B(n9934), .Z(n9898) );
  XNOR U12210 ( .A(n9901), .B(n9904), .Z(n9934) );
  NAND U12211 ( .A(n9935), .B(n9936), .Z(n9904) );
  NAND U12212 ( .A(n9937), .B(n9938), .Z(n9936) );
  OR U12213 ( .A(n9939), .B(n9940), .Z(n9937) );
  NANDN U12214 ( .A(n9941), .B(n9939), .Z(n9935) );
  IV U12215 ( .A(n9940), .Z(n9941) );
  NAND U12216 ( .A(n9942), .B(n9943), .Z(n9901) );
  NAND U12217 ( .A(n9944), .B(n9945), .Z(n9943) );
  NANDN U12218 ( .A(n9946), .B(n9947), .Z(n9944) );
  NANDN U12219 ( .A(n9947), .B(n9946), .Z(n9942) );
  AND U12220 ( .A(n9948), .B(n9949), .Z(n9903) );
  NAND U12221 ( .A(n9950), .B(n9951), .Z(n9949) );
  OR U12222 ( .A(n9952), .B(n9953), .Z(n9950) );
  NANDN U12223 ( .A(n9954), .B(n9952), .Z(n9948) );
  XNOR U12224 ( .A(n9929), .B(n9955), .Z(N13046) );
  XOR U12225 ( .A(n9931), .B(n9932), .Z(n9955) );
  XNOR U12226 ( .A(n9945), .B(n9956), .Z(n9932) );
  XOR U12227 ( .A(n9946), .B(n9947), .Z(n9956) );
  XOR U12228 ( .A(n9952), .B(n9957), .Z(n9947) );
  XOR U12229 ( .A(n9951), .B(n9954), .Z(n9957) );
  IV U12230 ( .A(n9953), .Z(n9954) );
  NAND U12231 ( .A(n9958), .B(n9959), .Z(n9953) );
  OR U12232 ( .A(n9960), .B(n9961), .Z(n9959) );
  OR U12233 ( .A(n9962), .B(n9963), .Z(n9958) );
  NAND U12234 ( .A(n9964), .B(n9965), .Z(n9951) );
  OR U12235 ( .A(n9966), .B(n9967), .Z(n9965) );
  OR U12236 ( .A(n9968), .B(n9969), .Z(n9964) );
  NOR U12237 ( .A(n9970), .B(n9971), .Z(n9952) );
  ANDN U12238 ( .B(n9972), .A(n9973), .Z(n9946) );
  XNOR U12239 ( .A(n9939), .B(n9974), .Z(n9945) );
  XNOR U12240 ( .A(n9938), .B(n9940), .Z(n9974) );
  NAND U12241 ( .A(n9975), .B(n9976), .Z(n9940) );
  OR U12242 ( .A(n9977), .B(n9978), .Z(n9976) );
  OR U12243 ( .A(n9979), .B(n9980), .Z(n9975) );
  NAND U12244 ( .A(n9981), .B(n9982), .Z(n9938) );
  OR U12245 ( .A(n9983), .B(n9984), .Z(n9982) );
  OR U12246 ( .A(n9985), .B(n9986), .Z(n9981) );
  ANDN U12247 ( .B(n9987), .A(n9988), .Z(n9939) );
  IV U12248 ( .A(n9989), .Z(n9987) );
  ANDN U12249 ( .B(n9990), .A(n9991), .Z(n9931) );
  XOR U12250 ( .A(n9917), .B(n9992), .Z(n9929) );
  XOR U12251 ( .A(n9918), .B(n9919), .Z(n9992) );
  XOR U12252 ( .A(n9924), .B(n9993), .Z(n9919) );
  XOR U12253 ( .A(n9923), .B(n9926), .Z(n9993) );
  IV U12254 ( .A(n9925), .Z(n9926) );
  NAND U12255 ( .A(n9994), .B(n9995), .Z(n9925) );
  OR U12256 ( .A(n9996), .B(n9997), .Z(n9995) );
  OR U12257 ( .A(n9998), .B(n9999), .Z(n9994) );
  NAND U12258 ( .A(n10000), .B(n10001), .Z(n9923) );
  OR U12259 ( .A(n10002), .B(n10003), .Z(n10001) );
  OR U12260 ( .A(n10004), .B(n10005), .Z(n10000) );
  NOR U12261 ( .A(n10006), .B(n10007), .Z(n9924) );
  ANDN U12262 ( .B(n10008), .A(n10009), .Z(n9918) );
  IV U12263 ( .A(n10010), .Z(n10008) );
  XNOR U12264 ( .A(n9911), .B(n10011), .Z(n9917) );
  XNOR U12265 ( .A(n9910), .B(n9912), .Z(n10011) );
  NAND U12266 ( .A(n10012), .B(n10013), .Z(n9912) );
  OR U12267 ( .A(n10014), .B(n10015), .Z(n10013) );
  OR U12268 ( .A(n10016), .B(n10017), .Z(n10012) );
  NAND U12269 ( .A(n10018), .B(n10019), .Z(n9910) );
  OR U12270 ( .A(n10020), .B(n10021), .Z(n10019) );
  OR U12271 ( .A(n10022), .B(n10023), .Z(n10018) );
  ANDN U12272 ( .B(n10024), .A(n10025), .Z(n9911) );
  IV U12273 ( .A(n10026), .Z(n10024) );
  XNOR U12274 ( .A(n9991), .B(n9990), .Z(N13045) );
  XOR U12275 ( .A(n10010), .B(n10009), .Z(n9990) );
  XNOR U12276 ( .A(n10025), .B(n10026), .Z(n10009) );
  XNOR U12277 ( .A(n10020), .B(n10021), .Z(n10026) );
  XNOR U12278 ( .A(n10022), .B(n10023), .Z(n10021) );
  XNOR U12279 ( .A(y[589]), .B(x[589]), .Z(n10023) );
  XNOR U12280 ( .A(y[590]), .B(x[590]), .Z(n10022) );
  XNOR U12281 ( .A(y[588]), .B(x[588]), .Z(n10020) );
  XNOR U12282 ( .A(n10014), .B(n10015), .Z(n10025) );
  XNOR U12283 ( .A(y[585]), .B(x[585]), .Z(n10015) );
  XNOR U12284 ( .A(n10016), .B(n10017), .Z(n10014) );
  XNOR U12285 ( .A(y[586]), .B(x[586]), .Z(n10017) );
  XNOR U12286 ( .A(y[587]), .B(x[587]), .Z(n10016) );
  XNOR U12287 ( .A(n10007), .B(n10006), .Z(n10010) );
  XNOR U12288 ( .A(n10002), .B(n10003), .Z(n10006) );
  XNOR U12289 ( .A(y[582]), .B(x[582]), .Z(n10003) );
  XNOR U12290 ( .A(n10004), .B(n10005), .Z(n10002) );
  XNOR U12291 ( .A(y[583]), .B(x[583]), .Z(n10005) );
  XNOR U12292 ( .A(y[584]), .B(x[584]), .Z(n10004) );
  XNOR U12293 ( .A(n9996), .B(n9997), .Z(n10007) );
  XNOR U12294 ( .A(y[579]), .B(x[579]), .Z(n9997) );
  XNOR U12295 ( .A(n9998), .B(n9999), .Z(n9996) );
  XNOR U12296 ( .A(y[580]), .B(x[580]), .Z(n9999) );
  XNOR U12297 ( .A(y[581]), .B(x[581]), .Z(n9998) );
  XOR U12298 ( .A(n9972), .B(n9973), .Z(n9991) );
  XNOR U12299 ( .A(n9988), .B(n9989), .Z(n9973) );
  XNOR U12300 ( .A(n9983), .B(n9984), .Z(n9989) );
  XNOR U12301 ( .A(n9985), .B(n9986), .Z(n9984) );
  XNOR U12302 ( .A(y[577]), .B(x[577]), .Z(n9986) );
  XNOR U12303 ( .A(y[578]), .B(x[578]), .Z(n9985) );
  XNOR U12304 ( .A(y[576]), .B(x[576]), .Z(n9983) );
  XNOR U12305 ( .A(n9977), .B(n9978), .Z(n9988) );
  XNOR U12306 ( .A(y[573]), .B(x[573]), .Z(n9978) );
  XNOR U12307 ( .A(n9979), .B(n9980), .Z(n9977) );
  XNOR U12308 ( .A(y[574]), .B(x[574]), .Z(n9980) );
  XNOR U12309 ( .A(y[575]), .B(x[575]), .Z(n9979) );
  XOR U12310 ( .A(n9971), .B(n9970), .Z(n9972) );
  XNOR U12311 ( .A(n9966), .B(n9967), .Z(n9970) );
  XNOR U12312 ( .A(y[570]), .B(x[570]), .Z(n9967) );
  XNOR U12313 ( .A(n9968), .B(n9969), .Z(n9966) );
  XNOR U12314 ( .A(y[571]), .B(x[571]), .Z(n9969) );
  XNOR U12315 ( .A(y[572]), .B(x[572]), .Z(n9968) );
  XNOR U12316 ( .A(n9960), .B(n9961), .Z(n9971) );
  XNOR U12317 ( .A(y[567]), .B(x[567]), .Z(n9961) );
  XNOR U12318 ( .A(n9962), .B(n9963), .Z(n9960) );
  XNOR U12319 ( .A(y[568]), .B(x[568]), .Z(n9963) );
  XNOR U12320 ( .A(y[569]), .B(x[569]), .Z(n9962) );
  NAND U12321 ( .A(n10027), .B(n10028), .Z(N13038) );
  NANDN U12322 ( .A(n10029), .B(n10030), .Z(n10028) );
  OR U12323 ( .A(n10031), .B(n10032), .Z(n10030) );
  NAND U12324 ( .A(n10031), .B(n10032), .Z(n10027) );
  XOR U12325 ( .A(n10031), .B(n10033), .Z(N13037) );
  XNOR U12326 ( .A(n10029), .B(n10032), .Z(n10033) );
  AND U12327 ( .A(n10034), .B(n10035), .Z(n10032) );
  NANDN U12328 ( .A(n10036), .B(n10037), .Z(n10035) );
  NANDN U12329 ( .A(n10038), .B(n10039), .Z(n10037) );
  NANDN U12330 ( .A(n10039), .B(n10038), .Z(n10034) );
  NAND U12331 ( .A(n10040), .B(n10041), .Z(n10029) );
  NANDN U12332 ( .A(n10042), .B(n10043), .Z(n10041) );
  OR U12333 ( .A(n10044), .B(n10045), .Z(n10043) );
  NAND U12334 ( .A(n10045), .B(n10044), .Z(n10040) );
  AND U12335 ( .A(n10046), .B(n10047), .Z(n10031) );
  NANDN U12336 ( .A(n10048), .B(n10049), .Z(n10047) );
  NANDN U12337 ( .A(n10050), .B(n10051), .Z(n10049) );
  NANDN U12338 ( .A(n10051), .B(n10050), .Z(n10046) );
  XOR U12339 ( .A(n10045), .B(n10052), .Z(N13036) );
  XOR U12340 ( .A(n10042), .B(n10044), .Z(n10052) );
  XNOR U12341 ( .A(n10038), .B(n10053), .Z(n10044) );
  XNOR U12342 ( .A(n10036), .B(n10039), .Z(n10053) );
  NAND U12343 ( .A(n10054), .B(n10055), .Z(n10039) );
  NAND U12344 ( .A(n10056), .B(n10057), .Z(n10055) );
  OR U12345 ( .A(n10058), .B(n10059), .Z(n10056) );
  NANDN U12346 ( .A(n10060), .B(n10058), .Z(n10054) );
  IV U12347 ( .A(n10059), .Z(n10060) );
  NAND U12348 ( .A(n10061), .B(n10062), .Z(n10036) );
  NAND U12349 ( .A(n10063), .B(n10064), .Z(n10062) );
  NANDN U12350 ( .A(n10065), .B(n10066), .Z(n10063) );
  NANDN U12351 ( .A(n10066), .B(n10065), .Z(n10061) );
  AND U12352 ( .A(n10067), .B(n10068), .Z(n10038) );
  NAND U12353 ( .A(n10069), .B(n10070), .Z(n10068) );
  OR U12354 ( .A(n10071), .B(n10072), .Z(n10069) );
  NANDN U12355 ( .A(n10073), .B(n10071), .Z(n10067) );
  NAND U12356 ( .A(n10074), .B(n10075), .Z(n10042) );
  NANDN U12357 ( .A(n10076), .B(n10077), .Z(n10075) );
  OR U12358 ( .A(n10078), .B(n10079), .Z(n10077) );
  NANDN U12359 ( .A(n10080), .B(n10078), .Z(n10074) );
  IV U12360 ( .A(n10079), .Z(n10080) );
  XNOR U12361 ( .A(n10050), .B(n10081), .Z(n10045) );
  XNOR U12362 ( .A(n10048), .B(n10051), .Z(n10081) );
  NAND U12363 ( .A(n10082), .B(n10083), .Z(n10051) );
  NAND U12364 ( .A(n10084), .B(n10085), .Z(n10083) );
  OR U12365 ( .A(n10086), .B(n10087), .Z(n10084) );
  NANDN U12366 ( .A(n10088), .B(n10086), .Z(n10082) );
  IV U12367 ( .A(n10087), .Z(n10088) );
  NAND U12368 ( .A(n10089), .B(n10090), .Z(n10048) );
  NAND U12369 ( .A(n10091), .B(n10092), .Z(n10090) );
  NANDN U12370 ( .A(n10093), .B(n10094), .Z(n10091) );
  NANDN U12371 ( .A(n10094), .B(n10093), .Z(n10089) );
  AND U12372 ( .A(n10095), .B(n10096), .Z(n10050) );
  NAND U12373 ( .A(n10097), .B(n10098), .Z(n10096) );
  OR U12374 ( .A(n10099), .B(n10100), .Z(n10097) );
  NANDN U12375 ( .A(n10101), .B(n10099), .Z(n10095) );
  XNOR U12376 ( .A(n10076), .B(n10102), .Z(N13035) );
  XOR U12377 ( .A(n10078), .B(n10079), .Z(n10102) );
  XNOR U12378 ( .A(n10092), .B(n10103), .Z(n10079) );
  XOR U12379 ( .A(n10093), .B(n10094), .Z(n10103) );
  XOR U12380 ( .A(n10099), .B(n10104), .Z(n10094) );
  XOR U12381 ( .A(n10098), .B(n10101), .Z(n10104) );
  IV U12382 ( .A(n10100), .Z(n10101) );
  NAND U12383 ( .A(n10105), .B(n10106), .Z(n10100) );
  OR U12384 ( .A(n10107), .B(n10108), .Z(n10106) );
  OR U12385 ( .A(n10109), .B(n10110), .Z(n10105) );
  NAND U12386 ( .A(n10111), .B(n10112), .Z(n10098) );
  OR U12387 ( .A(n10113), .B(n10114), .Z(n10112) );
  OR U12388 ( .A(n10115), .B(n10116), .Z(n10111) );
  NOR U12389 ( .A(n10117), .B(n10118), .Z(n10099) );
  ANDN U12390 ( .B(n10119), .A(n10120), .Z(n10093) );
  XNOR U12391 ( .A(n10086), .B(n10121), .Z(n10092) );
  XNOR U12392 ( .A(n10085), .B(n10087), .Z(n10121) );
  NAND U12393 ( .A(n10122), .B(n10123), .Z(n10087) );
  OR U12394 ( .A(n10124), .B(n10125), .Z(n10123) );
  OR U12395 ( .A(n10126), .B(n10127), .Z(n10122) );
  NAND U12396 ( .A(n10128), .B(n10129), .Z(n10085) );
  OR U12397 ( .A(n10130), .B(n10131), .Z(n10129) );
  OR U12398 ( .A(n10132), .B(n10133), .Z(n10128) );
  ANDN U12399 ( .B(n10134), .A(n10135), .Z(n10086) );
  IV U12400 ( .A(n10136), .Z(n10134) );
  ANDN U12401 ( .B(n10137), .A(n10138), .Z(n10078) );
  XOR U12402 ( .A(n10064), .B(n10139), .Z(n10076) );
  XOR U12403 ( .A(n10065), .B(n10066), .Z(n10139) );
  XOR U12404 ( .A(n10071), .B(n10140), .Z(n10066) );
  XOR U12405 ( .A(n10070), .B(n10073), .Z(n10140) );
  IV U12406 ( .A(n10072), .Z(n10073) );
  NAND U12407 ( .A(n10141), .B(n10142), .Z(n10072) );
  OR U12408 ( .A(n10143), .B(n10144), .Z(n10142) );
  OR U12409 ( .A(n10145), .B(n10146), .Z(n10141) );
  NAND U12410 ( .A(n10147), .B(n10148), .Z(n10070) );
  OR U12411 ( .A(n10149), .B(n10150), .Z(n10148) );
  OR U12412 ( .A(n10151), .B(n10152), .Z(n10147) );
  NOR U12413 ( .A(n10153), .B(n10154), .Z(n10071) );
  ANDN U12414 ( .B(n10155), .A(n10156), .Z(n10065) );
  IV U12415 ( .A(n10157), .Z(n10155) );
  XNOR U12416 ( .A(n10058), .B(n10158), .Z(n10064) );
  XNOR U12417 ( .A(n10057), .B(n10059), .Z(n10158) );
  NAND U12418 ( .A(n10159), .B(n10160), .Z(n10059) );
  OR U12419 ( .A(n10161), .B(n10162), .Z(n10160) );
  OR U12420 ( .A(n10163), .B(n10164), .Z(n10159) );
  NAND U12421 ( .A(n10165), .B(n10166), .Z(n10057) );
  OR U12422 ( .A(n10167), .B(n10168), .Z(n10166) );
  OR U12423 ( .A(n10169), .B(n10170), .Z(n10165) );
  ANDN U12424 ( .B(n10171), .A(n10172), .Z(n10058) );
  IV U12425 ( .A(n10173), .Z(n10171) );
  XNOR U12426 ( .A(n10138), .B(n10137), .Z(N13034) );
  XOR U12427 ( .A(n10157), .B(n10156), .Z(n10137) );
  XNOR U12428 ( .A(n10172), .B(n10173), .Z(n10156) );
  XNOR U12429 ( .A(n10167), .B(n10168), .Z(n10173) );
  XNOR U12430 ( .A(n10169), .B(n10170), .Z(n10168) );
  XNOR U12431 ( .A(y[565]), .B(x[565]), .Z(n10170) );
  XNOR U12432 ( .A(y[566]), .B(x[566]), .Z(n10169) );
  XNOR U12433 ( .A(y[564]), .B(x[564]), .Z(n10167) );
  XNOR U12434 ( .A(n10161), .B(n10162), .Z(n10172) );
  XNOR U12435 ( .A(y[561]), .B(x[561]), .Z(n10162) );
  XNOR U12436 ( .A(n10163), .B(n10164), .Z(n10161) );
  XNOR U12437 ( .A(y[562]), .B(x[562]), .Z(n10164) );
  XNOR U12438 ( .A(y[563]), .B(x[563]), .Z(n10163) );
  XNOR U12439 ( .A(n10154), .B(n10153), .Z(n10157) );
  XNOR U12440 ( .A(n10149), .B(n10150), .Z(n10153) );
  XNOR U12441 ( .A(y[558]), .B(x[558]), .Z(n10150) );
  XNOR U12442 ( .A(n10151), .B(n10152), .Z(n10149) );
  XNOR U12443 ( .A(y[559]), .B(x[559]), .Z(n10152) );
  XNOR U12444 ( .A(y[560]), .B(x[560]), .Z(n10151) );
  XNOR U12445 ( .A(n10143), .B(n10144), .Z(n10154) );
  XNOR U12446 ( .A(y[555]), .B(x[555]), .Z(n10144) );
  XNOR U12447 ( .A(n10145), .B(n10146), .Z(n10143) );
  XNOR U12448 ( .A(y[556]), .B(x[556]), .Z(n10146) );
  XNOR U12449 ( .A(y[557]), .B(x[557]), .Z(n10145) );
  XOR U12450 ( .A(n10119), .B(n10120), .Z(n10138) );
  XNOR U12451 ( .A(n10135), .B(n10136), .Z(n10120) );
  XNOR U12452 ( .A(n10130), .B(n10131), .Z(n10136) );
  XNOR U12453 ( .A(n10132), .B(n10133), .Z(n10131) );
  XNOR U12454 ( .A(y[553]), .B(x[553]), .Z(n10133) );
  XNOR U12455 ( .A(y[554]), .B(x[554]), .Z(n10132) );
  XNOR U12456 ( .A(y[552]), .B(x[552]), .Z(n10130) );
  XNOR U12457 ( .A(n10124), .B(n10125), .Z(n10135) );
  XNOR U12458 ( .A(y[549]), .B(x[549]), .Z(n10125) );
  XNOR U12459 ( .A(n10126), .B(n10127), .Z(n10124) );
  XNOR U12460 ( .A(y[550]), .B(x[550]), .Z(n10127) );
  XNOR U12461 ( .A(y[551]), .B(x[551]), .Z(n10126) );
  XOR U12462 ( .A(n10118), .B(n10117), .Z(n10119) );
  XNOR U12463 ( .A(n10113), .B(n10114), .Z(n10117) );
  XNOR U12464 ( .A(y[546]), .B(x[546]), .Z(n10114) );
  XNOR U12465 ( .A(n10115), .B(n10116), .Z(n10113) );
  XNOR U12466 ( .A(y[547]), .B(x[547]), .Z(n10116) );
  XNOR U12467 ( .A(y[548]), .B(x[548]), .Z(n10115) );
  XNOR U12468 ( .A(n10107), .B(n10108), .Z(n10118) );
  XNOR U12469 ( .A(y[543]), .B(x[543]), .Z(n10108) );
  XNOR U12470 ( .A(n10109), .B(n10110), .Z(n10107) );
  XNOR U12471 ( .A(y[544]), .B(x[544]), .Z(n10110) );
  XNOR U12472 ( .A(y[545]), .B(x[545]), .Z(n10109) );
  NAND U12473 ( .A(n10174), .B(n10175), .Z(N13027) );
  NANDN U12474 ( .A(n10176), .B(n10177), .Z(n10175) );
  OR U12475 ( .A(n10178), .B(n10179), .Z(n10177) );
  NAND U12476 ( .A(n10178), .B(n10179), .Z(n10174) );
  XOR U12477 ( .A(n10178), .B(n10180), .Z(N13026) );
  XNOR U12478 ( .A(n10176), .B(n10179), .Z(n10180) );
  AND U12479 ( .A(n10181), .B(n10182), .Z(n10179) );
  NANDN U12480 ( .A(n10183), .B(n10184), .Z(n10182) );
  NANDN U12481 ( .A(n10185), .B(n10186), .Z(n10184) );
  NANDN U12482 ( .A(n10186), .B(n10185), .Z(n10181) );
  NAND U12483 ( .A(n10187), .B(n10188), .Z(n10176) );
  NANDN U12484 ( .A(n10189), .B(n10190), .Z(n10188) );
  OR U12485 ( .A(n10191), .B(n10192), .Z(n10190) );
  NAND U12486 ( .A(n10192), .B(n10191), .Z(n10187) );
  AND U12487 ( .A(n10193), .B(n10194), .Z(n10178) );
  NANDN U12488 ( .A(n10195), .B(n10196), .Z(n10194) );
  NANDN U12489 ( .A(n10197), .B(n10198), .Z(n10196) );
  NANDN U12490 ( .A(n10198), .B(n10197), .Z(n10193) );
  XOR U12491 ( .A(n10192), .B(n10199), .Z(N13025) );
  XOR U12492 ( .A(n10189), .B(n10191), .Z(n10199) );
  XNOR U12493 ( .A(n10185), .B(n10200), .Z(n10191) );
  XNOR U12494 ( .A(n10183), .B(n10186), .Z(n10200) );
  NAND U12495 ( .A(n10201), .B(n10202), .Z(n10186) );
  NAND U12496 ( .A(n10203), .B(n10204), .Z(n10202) );
  OR U12497 ( .A(n10205), .B(n10206), .Z(n10203) );
  NANDN U12498 ( .A(n10207), .B(n10205), .Z(n10201) );
  IV U12499 ( .A(n10206), .Z(n10207) );
  NAND U12500 ( .A(n10208), .B(n10209), .Z(n10183) );
  NAND U12501 ( .A(n10210), .B(n10211), .Z(n10209) );
  NANDN U12502 ( .A(n10212), .B(n10213), .Z(n10210) );
  NANDN U12503 ( .A(n10213), .B(n10212), .Z(n10208) );
  AND U12504 ( .A(n10214), .B(n10215), .Z(n10185) );
  NAND U12505 ( .A(n10216), .B(n10217), .Z(n10215) );
  OR U12506 ( .A(n10218), .B(n10219), .Z(n10216) );
  NANDN U12507 ( .A(n10220), .B(n10218), .Z(n10214) );
  NAND U12508 ( .A(n10221), .B(n10222), .Z(n10189) );
  NANDN U12509 ( .A(n10223), .B(n10224), .Z(n10222) );
  OR U12510 ( .A(n10225), .B(n10226), .Z(n10224) );
  NANDN U12511 ( .A(n10227), .B(n10225), .Z(n10221) );
  IV U12512 ( .A(n10226), .Z(n10227) );
  XNOR U12513 ( .A(n10197), .B(n10228), .Z(n10192) );
  XNOR U12514 ( .A(n10195), .B(n10198), .Z(n10228) );
  NAND U12515 ( .A(n10229), .B(n10230), .Z(n10198) );
  NAND U12516 ( .A(n10231), .B(n10232), .Z(n10230) );
  OR U12517 ( .A(n10233), .B(n10234), .Z(n10231) );
  NANDN U12518 ( .A(n10235), .B(n10233), .Z(n10229) );
  IV U12519 ( .A(n10234), .Z(n10235) );
  NAND U12520 ( .A(n10236), .B(n10237), .Z(n10195) );
  NAND U12521 ( .A(n10238), .B(n10239), .Z(n10237) );
  NANDN U12522 ( .A(n10240), .B(n10241), .Z(n10238) );
  NANDN U12523 ( .A(n10241), .B(n10240), .Z(n10236) );
  AND U12524 ( .A(n10242), .B(n10243), .Z(n10197) );
  NAND U12525 ( .A(n10244), .B(n10245), .Z(n10243) );
  OR U12526 ( .A(n10246), .B(n10247), .Z(n10244) );
  NANDN U12527 ( .A(n10248), .B(n10246), .Z(n10242) );
  XNOR U12528 ( .A(n10223), .B(n10249), .Z(N13024) );
  XOR U12529 ( .A(n10225), .B(n10226), .Z(n10249) );
  XNOR U12530 ( .A(n10239), .B(n10250), .Z(n10226) );
  XOR U12531 ( .A(n10240), .B(n10241), .Z(n10250) );
  XOR U12532 ( .A(n10246), .B(n10251), .Z(n10241) );
  XOR U12533 ( .A(n10245), .B(n10248), .Z(n10251) );
  IV U12534 ( .A(n10247), .Z(n10248) );
  NAND U12535 ( .A(n10252), .B(n10253), .Z(n10247) );
  OR U12536 ( .A(n10254), .B(n10255), .Z(n10253) );
  OR U12537 ( .A(n10256), .B(n10257), .Z(n10252) );
  NAND U12538 ( .A(n10258), .B(n10259), .Z(n10245) );
  OR U12539 ( .A(n10260), .B(n10261), .Z(n10259) );
  OR U12540 ( .A(n10262), .B(n10263), .Z(n10258) );
  NOR U12541 ( .A(n10264), .B(n10265), .Z(n10246) );
  ANDN U12542 ( .B(n10266), .A(n10267), .Z(n10240) );
  XNOR U12543 ( .A(n10233), .B(n10268), .Z(n10239) );
  XNOR U12544 ( .A(n10232), .B(n10234), .Z(n10268) );
  NAND U12545 ( .A(n10269), .B(n10270), .Z(n10234) );
  OR U12546 ( .A(n10271), .B(n10272), .Z(n10270) );
  OR U12547 ( .A(n10273), .B(n10274), .Z(n10269) );
  NAND U12548 ( .A(n10275), .B(n10276), .Z(n10232) );
  OR U12549 ( .A(n10277), .B(n10278), .Z(n10276) );
  OR U12550 ( .A(n10279), .B(n10280), .Z(n10275) );
  ANDN U12551 ( .B(n10281), .A(n10282), .Z(n10233) );
  IV U12552 ( .A(n10283), .Z(n10281) );
  ANDN U12553 ( .B(n10284), .A(n10285), .Z(n10225) );
  XOR U12554 ( .A(n10211), .B(n10286), .Z(n10223) );
  XOR U12555 ( .A(n10212), .B(n10213), .Z(n10286) );
  XOR U12556 ( .A(n10218), .B(n10287), .Z(n10213) );
  XOR U12557 ( .A(n10217), .B(n10220), .Z(n10287) );
  IV U12558 ( .A(n10219), .Z(n10220) );
  NAND U12559 ( .A(n10288), .B(n10289), .Z(n10219) );
  OR U12560 ( .A(n10290), .B(n10291), .Z(n10289) );
  OR U12561 ( .A(n10292), .B(n10293), .Z(n10288) );
  NAND U12562 ( .A(n10294), .B(n10295), .Z(n10217) );
  OR U12563 ( .A(n10296), .B(n10297), .Z(n10295) );
  OR U12564 ( .A(n10298), .B(n10299), .Z(n10294) );
  NOR U12565 ( .A(n10300), .B(n10301), .Z(n10218) );
  ANDN U12566 ( .B(n10302), .A(n10303), .Z(n10212) );
  IV U12567 ( .A(n10304), .Z(n10302) );
  XNOR U12568 ( .A(n10205), .B(n10305), .Z(n10211) );
  XNOR U12569 ( .A(n10204), .B(n10206), .Z(n10305) );
  NAND U12570 ( .A(n10306), .B(n10307), .Z(n10206) );
  OR U12571 ( .A(n10308), .B(n10309), .Z(n10307) );
  OR U12572 ( .A(n10310), .B(n10311), .Z(n10306) );
  NAND U12573 ( .A(n10312), .B(n10313), .Z(n10204) );
  OR U12574 ( .A(n10314), .B(n10315), .Z(n10313) );
  OR U12575 ( .A(n10316), .B(n10317), .Z(n10312) );
  ANDN U12576 ( .B(n10318), .A(n10319), .Z(n10205) );
  IV U12577 ( .A(n10320), .Z(n10318) );
  XNOR U12578 ( .A(n10285), .B(n10284), .Z(N13023) );
  XOR U12579 ( .A(n10304), .B(n10303), .Z(n10284) );
  XNOR U12580 ( .A(n10319), .B(n10320), .Z(n10303) );
  XNOR U12581 ( .A(n10314), .B(n10315), .Z(n10320) );
  XNOR U12582 ( .A(n10316), .B(n10317), .Z(n10315) );
  XNOR U12583 ( .A(y[541]), .B(x[541]), .Z(n10317) );
  XNOR U12584 ( .A(y[542]), .B(x[542]), .Z(n10316) );
  XNOR U12585 ( .A(y[540]), .B(x[540]), .Z(n10314) );
  XNOR U12586 ( .A(n10308), .B(n10309), .Z(n10319) );
  XNOR U12587 ( .A(y[537]), .B(x[537]), .Z(n10309) );
  XNOR U12588 ( .A(n10310), .B(n10311), .Z(n10308) );
  XNOR U12589 ( .A(y[538]), .B(x[538]), .Z(n10311) );
  XNOR U12590 ( .A(y[539]), .B(x[539]), .Z(n10310) );
  XNOR U12591 ( .A(n10301), .B(n10300), .Z(n10304) );
  XNOR U12592 ( .A(n10296), .B(n10297), .Z(n10300) );
  XNOR U12593 ( .A(y[534]), .B(x[534]), .Z(n10297) );
  XNOR U12594 ( .A(n10298), .B(n10299), .Z(n10296) );
  XNOR U12595 ( .A(y[535]), .B(x[535]), .Z(n10299) );
  XNOR U12596 ( .A(y[536]), .B(x[536]), .Z(n10298) );
  XNOR U12597 ( .A(n10290), .B(n10291), .Z(n10301) );
  XNOR U12598 ( .A(y[531]), .B(x[531]), .Z(n10291) );
  XNOR U12599 ( .A(n10292), .B(n10293), .Z(n10290) );
  XNOR U12600 ( .A(y[532]), .B(x[532]), .Z(n10293) );
  XNOR U12601 ( .A(y[533]), .B(x[533]), .Z(n10292) );
  XOR U12602 ( .A(n10266), .B(n10267), .Z(n10285) );
  XNOR U12603 ( .A(n10282), .B(n10283), .Z(n10267) );
  XNOR U12604 ( .A(n10277), .B(n10278), .Z(n10283) );
  XNOR U12605 ( .A(n10279), .B(n10280), .Z(n10278) );
  XNOR U12606 ( .A(y[529]), .B(x[529]), .Z(n10280) );
  XNOR U12607 ( .A(y[530]), .B(x[530]), .Z(n10279) );
  XNOR U12608 ( .A(y[528]), .B(x[528]), .Z(n10277) );
  XNOR U12609 ( .A(n10271), .B(n10272), .Z(n10282) );
  XNOR U12610 ( .A(y[525]), .B(x[525]), .Z(n10272) );
  XNOR U12611 ( .A(n10273), .B(n10274), .Z(n10271) );
  XNOR U12612 ( .A(y[526]), .B(x[526]), .Z(n10274) );
  XNOR U12613 ( .A(y[527]), .B(x[527]), .Z(n10273) );
  XOR U12614 ( .A(n10265), .B(n10264), .Z(n10266) );
  XNOR U12615 ( .A(n10260), .B(n10261), .Z(n10264) );
  XNOR U12616 ( .A(y[522]), .B(x[522]), .Z(n10261) );
  XNOR U12617 ( .A(n10262), .B(n10263), .Z(n10260) );
  XNOR U12618 ( .A(y[523]), .B(x[523]), .Z(n10263) );
  XNOR U12619 ( .A(y[524]), .B(x[524]), .Z(n10262) );
  XNOR U12620 ( .A(n10254), .B(n10255), .Z(n10265) );
  XNOR U12621 ( .A(y[519]), .B(x[519]), .Z(n10255) );
  XNOR U12622 ( .A(n10256), .B(n10257), .Z(n10254) );
  XNOR U12623 ( .A(y[520]), .B(x[520]), .Z(n10257) );
  XNOR U12624 ( .A(y[521]), .B(x[521]), .Z(n10256) );
  NAND U12625 ( .A(n10321), .B(n10322), .Z(N13016) );
  NANDN U12626 ( .A(n10323), .B(n10324), .Z(n10322) );
  OR U12627 ( .A(n10325), .B(n10326), .Z(n10324) );
  NAND U12628 ( .A(n10325), .B(n10326), .Z(n10321) );
  XOR U12629 ( .A(n10325), .B(n10327), .Z(N13015) );
  XNOR U12630 ( .A(n10323), .B(n10326), .Z(n10327) );
  AND U12631 ( .A(n10328), .B(n10329), .Z(n10326) );
  NANDN U12632 ( .A(n10330), .B(n10331), .Z(n10329) );
  NANDN U12633 ( .A(n10332), .B(n10333), .Z(n10331) );
  NANDN U12634 ( .A(n10333), .B(n10332), .Z(n10328) );
  NAND U12635 ( .A(n10334), .B(n10335), .Z(n10323) );
  NANDN U12636 ( .A(n10336), .B(n10337), .Z(n10335) );
  OR U12637 ( .A(n10338), .B(n10339), .Z(n10337) );
  NAND U12638 ( .A(n10339), .B(n10338), .Z(n10334) );
  AND U12639 ( .A(n10340), .B(n10341), .Z(n10325) );
  NANDN U12640 ( .A(n10342), .B(n10343), .Z(n10341) );
  NANDN U12641 ( .A(n10344), .B(n10345), .Z(n10343) );
  NANDN U12642 ( .A(n10345), .B(n10344), .Z(n10340) );
  XOR U12643 ( .A(n10339), .B(n10346), .Z(N13014) );
  XOR U12644 ( .A(n10336), .B(n10338), .Z(n10346) );
  XNOR U12645 ( .A(n10332), .B(n10347), .Z(n10338) );
  XNOR U12646 ( .A(n10330), .B(n10333), .Z(n10347) );
  NAND U12647 ( .A(n10348), .B(n10349), .Z(n10333) );
  NAND U12648 ( .A(n10350), .B(n10351), .Z(n10349) );
  OR U12649 ( .A(n10352), .B(n10353), .Z(n10350) );
  NANDN U12650 ( .A(n10354), .B(n10352), .Z(n10348) );
  IV U12651 ( .A(n10353), .Z(n10354) );
  NAND U12652 ( .A(n10355), .B(n10356), .Z(n10330) );
  NAND U12653 ( .A(n10357), .B(n10358), .Z(n10356) );
  NANDN U12654 ( .A(n10359), .B(n10360), .Z(n10357) );
  NANDN U12655 ( .A(n10360), .B(n10359), .Z(n10355) );
  AND U12656 ( .A(n10361), .B(n10362), .Z(n10332) );
  NAND U12657 ( .A(n10363), .B(n10364), .Z(n10362) );
  OR U12658 ( .A(n10365), .B(n10366), .Z(n10363) );
  NANDN U12659 ( .A(n10367), .B(n10365), .Z(n10361) );
  NAND U12660 ( .A(n10368), .B(n10369), .Z(n10336) );
  NANDN U12661 ( .A(n10370), .B(n10371), .Z(n10369) );
  OR U12662 ( .A(n10372), .B(n10373), .Z(n10371) );
  NANDN U12663 ( .A(n10374), .B(n10372), .Z(n10368) );
  IV U12664 ( .A(n10373), .Z(n10374) );
  XNOR U12665 ( .A(n10344), .B(n10375), .Z(n10339) );
  XNOR U12666 ( .A(n10342), .B(n10345), .Z(n10375) );
  NAND U12667 ( .A(n10376), .B(n10377), .Z(n10345) );
  NAND U12668 ( .A(n10378), .B(n10379), .Z(n10377) );
  OR U12669 ( .A(n10380), .B(n10381), .Z(n10378) );
  NANDN U12670 ( .A(n10382), .B(n10380), .Z(n10376) );
  IV U12671 ( .A(n10381), .Z(n10382) );
  NAND U12672 ( .A(n10383), .B(n10384), .Z(n10342) );
  NAND U12673 ( .A(n10385), .B(n10386), .Z(n10384) );
  NANDN U12674 ( .A(n10387), .B(n10388), .Z(n10385) );
  NANDN U12675 ( .A(n10388), .B(n10387), .Z(n10383) );
  AND U12676 ( .A(n10389), .B(n10390), .Z(n10344) );
  NAND U12677 ( .A(n10391), .B(n10392), .Z(n10390) );
  OR U12678 ( .A(n10393), .B(n10394), .Z(n10391) );
  NANDN U12679 ( .A(n10395), .B(n10393), .Z(n10389) );
  XNOR U12680 ( .A(n10370), .B(n10396), .Z(N13013) );
  XOR U12681 ( .A(n10372), .B(n10373), .Z(n10396) );
  XNOR U12682 ( .A(n10386), .B(n10397), .Z(n10373) );
  XOR U12683 ( .A(n10387), .B(n10388), .Z(n10397) );
  XOR U12684 ( .A(n10393), .B(n10398), .Z(n10388) );
  XOR U12685 ( .A(n10392), .B(n10395), .Z(n10398) );
  IV U12686 ( .A(n10394), .Z(n10395) );
  NAND U12687 ( .A(n10399), .B(n10400), .Z(n10394) );
  OR U12688 ( .A(n10401), .B(n10402), .Z(n10400) );
  OR U12689 ( .A(n10403), .B(n10404), .Z(n10399) );
  NAND U12690 ( .A(n10405), .B(n10406), .Z(n10392) );
  OR U12691 ( .A(n10407), .B(n10408), .Z(n10406) );
  OR U12692 ( .A(n10409), .B(n10410), .Z(n10405) );
  NOR U12693 ( .A(n10411), .B(n10412), .Z(n10393) );
  ANDN U12694 ( .B(n10413), .A(n10414), .Z(n10387) );
  XNOR U12695 ( .A(n10380), .B(n10415), .Z(n10386) );
  XNOR U12696 ( .A(n10379), .B(n10381), .Z(n10415) );
  NAND U12697 ( .A(n10416), .B(n10417), .Z(n10381) );
  OR U12698 ( .A(n10418), .B(n10419), .Z(n10417) );
  OR U12699 ( .A(n10420), .B(n10421), .Z(n10416) );
  NAND U12700 ( .A(n10422), .B(n10423), .Z(n10379) );
  OR U12701 ( .A(n10424), .B(n10425), .Z(n10423) );
  OR U12702 ( .A(n10426), .B(n10427), .Z(n10422) );
  ANDN U12703 ( .B(n10428), .A(n10429), .Z(n10380) );
  IV U12704 ( .A(n10430), .Z(n10428) );
  ANDN U12705 ( .B(n10431), .A(n10432), .Z(n10372) );
  XOR U12706 ( .A(n10358), .B(n10433), .Z(n10370) );
  XOR U12707 ( .A(n10359), .B(n10360), .Z(n10433) );
  XOR U12708 ( .A(n10365), .B(n10434), .Z(n10360) );
  XOR U12709 ( .A(n10364), .B(n10367), .Z(n10434) );
  IV U12710 ( .A(n10366), .Z(n10367) );
  NAND U12711 ( .A(n10435), .B(n10436), .Z(n10366) );
  OR U12712 ( .A(n10437), .B(n10438), .Z(n10436) );
  OR U12713 ( .A(n10439), .B(n10440), .Z(n10435) );
  NAND U12714 ( .A(n10441), .B(n10442), .Z(n10364) );
  OR U12715 ( .A(n10443), .B(n10444), .Z(n10442) );
  OR U12716 ( .A(n10445), .B(n10446), .Z(n10441) );
  NOR U12717 ( .A(n10447), .B(n10448), .Z(n10365) );
  ANDN U12718 ( .B(n10449), .A(n10450), .Z(n10359) );
  IV U12719 ( .A(n10451), .Z(n10449) );
  XNOR U12720 ( .A(n10352), .B(n10452), .Z(n10358) );
  XNOR U12721 ( .A(n10351), .B(n10353), .Z(n10452) );
  NAND U12722 ( .A(n10453), .B(n10454), .Z(n10353) );
  OR U12723 ( .A(n10455), .B(n10456), .Z(n10454) );
  OR U12724 ( .A(n10457), .B(n10458), .Z(n10453) );
  NAND U12725 ( .A(n10459), .B(n10460), .Z(n10351) );
  OR U12726 ( .A(n10461), .B(n10462), .Z(n10460) );
  OR U12727 ( .A(n10463), .B(n10464), .Z(n10459) );
  ANDN U12728 ( .B(n10465), .A(n10466), .Z(n10352) );
  IV U12729 ( .A(n10467), .Z(n10465) );
  XNOR U12730 ( .A(n10432), .B(n10431), .Z(N13012) );
  XOR U12731 ( .A(n10451), .B(n10450), .Z(n10431) );
  XNOR U12732 ( .A(n10466), .B(n10467), .Z(n10450) );
  XNOR U12733 ( .A(n10461), .B(n10462), .Z(n10467) );
  XNOR U12734 ( .A(n10463), .B(n10464), .Z(n10462) );
  XNOR U12735 ( .A(y[517]), .B(x[517]), .Z(n10464) );
  XNOR U12736 ( .A(y[518]), .B(x[518]), .Z(n10463) );
  XNOR U12737 ( .A(y[516]), .B(x[516]), .Z(n10461) );
  XNOR U12738 ( .A(n10455), .B(n10456), .Z(n10466) );
  XNOR U12739 ( .A(y[513]), .B(x[513]), .Z(n10456) );
  XNOR U12740 ( .A(n10457), .B(n10458), .Z(n10455) );
  XNOR U12741 ( .A(y[514]), .B(x[514]), .Z(n10458) );
  XNOR U12742 ( .A(y[515]), .B(x[515]), .Z(n10457) );
  XNOR U12743 ( .A(n10448), .B(n10447), .Z(n10451) );
  XNOR U12744 ( .A(n10443), .B(n10444), .Z(n10447) );
  XNOR U12745 ( .A(y[510]), .B(x[510]), .Z(n10444) );
  XNOR U12746 ( .A(n10445), .B(n10446), .Z(n10443) );
  XNOR U12747 ( .A(y[511]), .B(x[511]), .Z(n10446) );
  XNOR U12748 ( .A(y[512]), .B(x[512]), .Z(n10445) );
  XNOR U12749 ( .A(n10437), .B(n10438), .Z(n10448) );
  XNOR U12750 ( .A(y[507]), .B(x[507]), .Z(n10438) );
  XNOR U12751 ( .A(n10439), .B(n10440), .Z(n10437) );
  XNOR U12752 ( .A(y[508]), .B(x[508]), .Z(n10440) );
  XNOR U12753 ( .A(y[509]), .B(x[509]), .Z(n10439) );
  XOR U12754 ( .A(n10413), .B(n10414), .Z(n10432) );
  XNOR U12755 ( .A(n10429), .B(n10430), .Z(n10414) );
  XNOR U12756 ( .A(n10424), .B(n10425), .Z(n10430) );
  XNOR U12757 ( .A(n10426), .B(n10427), .Z(n10425) );
  XNOR U12758 ( .A(y[505]), .B(x[505]), .Z(n10427) );
  XNOR U12759 ( .A(y[506]), .B(x[506]), .Z(n10426) );
  XNOR U12760 ( .A(y[504]), .B(x[504]), .Z(n10424) );
  XNOR U12761 ( .A(n10418), .B(n10419), .Z(n10429) );
  XNOR U12762 ( .A(y[501]), .B(x[501]), .Z(n10419) );
  XNOR U12763 ( .A(n10420), .B(n10421), .Z(n10418) );
  XNOR U12764 ( .A(y[502]), .B(x[502]), .Z(n10421) );
  XNOR U12765 ( .A(y[503]), .B(x[503]), .Z(n10420) );
  XOR U12766 ( .A(n10412), .B(n10411), .Z(n10413) );
  XNOR U12767 ( .A(n10407), .B(n10408), .Z(n10411) );
  XNOR U12768 ( .A(y[498]), .B(x[498]), .Z(n10408) );
  XNOR U12769 ( .A(n10409), .B(n10410), .Z(n10407) );
  XNOR U12770 ( .A(y[499]), .B(x[499]), .Z(n10410) );
  XNOR U12771 ( .A(y[500]), .B(x[500]), .Z(n10409) );
  XNOR U12772 ( .A(n10401), .B(n10402), .Z(n10412) );
  XNOR U12773 ( .A(y[495]), .B(x[495]), .Z(n10402) );
  XNOR U12774 ( .A(n10403), .B(n10404), .Z(n10401) );
  XNOR U12775 ( .A(y[496]), .B(x[496]), .Z(n10404) );
  XNOR U12776 ( .A(y[497]), .B(x[497]), .Z(n10403) );
  NAND U12777 ( .A(n10468), .B(n10469), .Z(N13005) );
  NANDN U12778 ( .A(n10470), .B(n10471), .Z(n10469) );
  OR U12779 ( .A(n10472), .B(n10473), .Z(n10471) );
  NAND U12780 ( .A(n10472), .B(n10473), .Z(n10468) );
  XOR U12781 ( .A(n10472), .B(n10474), .Z(N13004) );
  XNOR U12782 ( .A(n10470), .B(n10473), .Z(n10474) );
  AND U12783 ( .A(n10475), .B(n10476), .Z(n10473) );
  NANDN U12784 ( .A(n10477), .B(n10478), .Z(n10476) );
  NANDN U12785 ( .A(n10479), .B(n10480), .Z(n10478) );
  NANDN U12786 ( .A(n10480), .B(n10479), .Z(n10475) );
  NAND U12787 ( .A(n10481), .B(n10482), .Z(n10470) );
  NANDN U12788 ( .A(n10483), .B(n10484), .Z(n10482) );
  OR U12789 ( .A(n10485), .B(n10486), .Z(n10484) );
  NAND U12790 ( .A(n10486), .B(n10485), .Z(n10481) );
  AND U12791 ( .A(n10487), .B(n10488), .Z(n10472) );
  NANDN U12792 ( .A(n10489), .B(n10490), .Z(n10488) );
  NANDN U12793 ( .A(n10491), .B(n10492), .Z(n10490) );
  NANDN U12794 ( .A(n10492), .B(n10491), .Z(n10487) );
  XOR U12795 ( .A(n10486), .B(n10493), .Z(N13003) );
  XOR U12796 ( .A(n10483), .B(n10485), .Z(n10493) );
  XNOR U12797 ( .A(n10479), .B(n10494), .Z(n10485) );
  XNOR U12798 ( .A(n10477), .B(n10480), .Z(n10494) );
  NAND U12799 ( .A(n10495), .B(n10496), .Z(n10480) );
  NAND U12800 ( .A(n10497), .B(n10498), .Z(n10496) );
  OR U12801 ( .A(n10499), .B(n10500), .Z(n10497) );
  NANDN U12802 ( .A(n10501), .B(n10499), .Z(n10495) );
  IV U12803 ( .A(n10500), .Z(n10501) );
  NAND U12804 ( .A(n10502), .B(n10503), .Z(n10477) );
  NAND U12805 ( .A(n10504), .B(n10505), .Z(n10503) );
  NANDN U12806 ( .A(n10506), .B(n10507), .Z(n10504) );
  NANDN U12807 ( .A(n10507), .B(n10506), .Z(n10502) );
  AND U12808 ( .A(n10508), .B(n10509), .Z(n10479) );
  NAND U12809 ( .A(n10510), .B(n10511), .Z(n10509) );
  OR U12810 ( .A(n10512), .B(n10513), .Z(n10510) );
  NANDN U12811 ( .A(n10514), .B(n10512), .Z(n10508) );
  NAND U12812 ( .A(n10515), .B(n10516), .Z(n10483) );
  NANDN U12813 ( .A(n10517), .B(n10518), .Z(n10516) );
  OR U12814 ( .A(n10519), .B(n10520), .Z(n10518) );
  NANDN U12815 ( .A(n10521), .B(n10519), .Z(n10515) );
  IV U12816 ( .A(n10520), .Z(n10521) );
  XNOR U12817 ( .A(n10491), .B(n10522), .Z(n10486) );
  XNOR U12818 ( .A(n10489), .B(n10492), .Z(n10522) );
  NAND U12819 ( .A(n10523), .B(n10524), .Z(n10492) );
  NAND U12820 ( .A(n10525), .B(n10526), .Z(n10524) );
  OR U12821 ( .A(n10527), .B(n10528), .Z(n10525) );
  NANDN U12822 ( .A(n10529), .B(n10527), .Z(n10523) );
  IV U12823 ( .A(n10528), .Z(n10529) );
  NAND U12824 ( .A(n10530), .B(n10531), .Z(n10489) );
  NAND U12825 ( .A(n10532), .B(n10533), .Z(n10531) );
  NANDN U12826 ( .A(n10534), .B(n10535), .Z(n10532) );
  NANDN U12827 ( .A(n10535), .B(n10534), .Z(n10530) );
  AND U12828 ( .A(n10536), .B(n10537), .Z(n10491) );
  NAND U12829 ( .A(n10538), .B(n10539), .Z(n10537) );
  OR U12830 ( .A(n10540), .B(n10541), .Z(n10538) );
  NANDN U12831 ( .A(n10542), .B(n10540), .Z(n10536) );
  XNOR U12832 ( .A(n10517), .B(n10543), .Z(N13002) );
  XOR U12833 ( .A(n10519), .B(n10520), .Z(n10543) );
  XNOR U12834 ( .A(n10533), .B(n10544), .Z(n10520) );
  XOR U12835 ( .A(n10534), .B(n10535), .Z(n10544) );
  XOR U12836 ( .A(n10540), .B(n10545), .Z(n10535) );
  XOR U12837 ( .A(n10539), .B(n10542), .Z(n10545) );
  IV U12838 ( .A(n10541), .Z(n10542) );
  NAND U12839 ( .A(n10546), .B(n10547), .Z(n10541) );
  OR U12840 ( .A(n10548), .B(n10549), .Z(n10547) );
  OR U12841 ( .A(n10550), .B(n10551), .Z(n10546) );
  NAND U12842 ( .A(n10552), .B(n10553), .Z(n10539) );
  OR U12843 ( .A(n10554), .B(n10555), .Z(n10553) );
  OR U12844 ( .A(n10556), .B(n10557), .Z(n10552) );
  NOR U12845 ( .A(n10558), .B(n10559), .Z(n10540) );
  ANDN U12846 ( .B(n10560), .A(n10561), .Z(n10534) );
  XNOR U12847 ( .A(n10527), .B(n10562), .Z(n10533) );
  XNOR U12848 ( .A(n10526), .B(n10528), .Z(n10562) );
  NAND U12849 ( .A(n10563), .B(n10564), .Z(n10528) );
  OR U12850 ( .A(n10565), .B(n10566), .Z(n10564) );
  OR U12851 ( .A(n10567), .B(n10568), .Z(n10563) );
  NAND U12852 ( .A(n10569), .B(n10570), .Z(n10526) );
  OR U12853 ( .A(n10571), .B(n10572), .Z(n10570) );
  OR U12854 ( .A(n10573), .B(n10574), .Z(n10569) );
  ANDN U12855 ( .B(n10575), .A(n10576), .Z(n10527) );
  IV U12856 ( .A(n10577), .Z(n10575) );
  ANDN U12857 ( .B(n10578), .A(n10579), .Z(n10519) );
  XOR U12858 ( .A(n10505), .B(n10580), .Z(n10517) );
  XOR U12859 ( .A(n10506), .B(n10507), .Z(n10580) );
  XOR U12860 ( .A(n10512), .B(n10581), .Z(n10507) );
  XOR U12861 ( .A(n10511), .B(n10514), .Z(n10581) );
  IV U12862 ( .A(n10513), .Z(n10514) );
  NAND U12863 ( .A(n10582), .B(n10583), .Z(n10513) );
  OR U12864 ( .A(n10584), .B(n10585), .Z(n10583) );
  OR U12865 ( .A(n10586), .B(n10587), .Z(n10582) );
  NAND U12866 ( .A(n10588), .B(n10589), .Z(n10511) );
  OR U12867 ( .A(n10590), .B(n10591), .Z(n10589) );
  OR U12868 ( .A(n10592), .B(n10593), .Z(n10588) );
  NOR U12869 ( .A(n10594), .B(n10595), .Z(n10512) );
  ANDN U12870 ( .B(n10596), .A(n10597), .Z(n10506) );
  IV U12871 ( .A(n10598), .Z(n10596) );
  XNOR U12872 ( .A(n10499), .B(n10599), .Z(n10505) );
  XNOR U12873 ( .A(n10498), .B(n10500), .Z(n10599) );
  NAND U12874 ( .A(n10600), .B(n10601), .Z(n10500) );
  OR U12875 ( .A(n10602), .B(n10603), .Z(n10601) );
  OR U12876 ( .A(n10604), .B(n10605), .Z(n10600) );
  NAND U12877 ( .A(n10606), .B(n10607), .Z(n10498) );
  OR U12878 ( .A(n10608), .B(n10609), .Z(n10607) );
  OR U12879 ( .A(n10610), .B(n10611), .Z(n10606) );
  ANDN U12880 ( .B(n10612), .A(n10613), .Z(n10499) );
  IV U12881 ( .A(n10614), .Z(n10612) );
  XNOR U12882 ( .A(n10579), .B(n10578), .Z(N13001) );
  XOR U12883 ( .A(n10598), .B(n10597), .Z(n10578) );
  XNOR U12884 ( .A(n10613), .B(n10614), .Z(n10597) );
  XNOR U12885 ( .A(n10608), .B(n10609), .Z(n10614) );
  XNOR U12886 ( .A(n10610), .B(n10611), .Z(n10609) );
  XNOR U12887 ( .A(y[493]), .B(x[493]), .Z(n10611) );
  XNOR U12888 ( .A(y[494]), .B(x[494]), .Z(n10610) );
  XNOR U12889 ( .A(y[492]), .B(x[492]), .Z(n10608) );
  XNOR U12890 ( .A(n10602), .B(n10603), .Z(n10613) );
  XNOR U12891 ( .A(y[489]), .B(x[489]), .Z(n10603) );
  XNOR U12892 ( .A(n10604), .B(n10605), .Z(n10602) );
  XNOR U12893 ( .A(y[490]), .B(x[490]), .Z(n10605) );
  XNOR U12894 ( .A(y[491]), .B(x[491]), .Z(n10604) );
  XNOR U12895 ( .A(n10595), .B(n10594), .Z(n10598) );
  XNOR U12896 ( .A(n10590), .B(n10591), .Z(n10594) );
  XNOR U12897 ( .A(y[486]), .B(x[486]), .Z(n10591) );
  XNOR U12898 ( .A(n10592), .B(n10593), .Z(n10590) );
  XNOR U12899 ( .A(y[487]), .B(x[487]), .Z(n10593) );
  XNOR U12900 ( .A(y[488]), .B(x[488]), .Z(n10592) );
  XNOR U12901 ( .A(n10584), .B(n10585), .Z(n10595) );
  XNOR U12902 ( .A(y[483]), .B(x[483]), .Z(n10585) );
  XNOR U12903 ( .A(n10586), .B(n10587), .Z(n10584) );
  XNOR U12904 ( .A(y[484]), .B(x[484]), .Z(n10587) );
  XNOR U12905 ( .A(y[485]), .B(x[485]), .Z(n10586) );
  XOR U12906 ( .A(n10560), .B(n10561), .Z(n10579) );
  XNOR U12907 ( .A(n10576), .B(n10577), .Z(n10561) );
  XNOR U12908 ( .A(n10571), .B(n10572), .Z(n10577) );
  XNOR U12909 ( .A(n10573), .B(n10574), .Z(n10572) );
  XNOR U12910 ( .A(y[481]), .B(x[481]), .Z(n10574) );
  XNOR U12911 ( .A(y[482]), .B(x[482]), .Z(n10573) );
  XNOR U12912 ( .A(y[480]), .B(x[480]), .Z(n10571) );
  XNOR U12913 ( .A(n10565), .B(n10566), .Z(n10576) );
  XNOR U12914 ( .A(y[477]), .B(x[477]), .Z(n10566) );
  XNOR U12915 ( .A(n10567), .B(n10568), .Z(n10565) );
  XNOR U12916 ( .A(y[478]), .B(x[478]), .Z(n10568) );
  XNOR U12917 ( .A(y[479]), .B(x[479]), .Z(n10567) );
  XOR U12918 ( .A(n10559), .B(n10558), .Z(n10560) );
  XNOR U12919 ( .A(n10554), .B(n10555), .Z(n10558) );
  XNOR U12920 ( .A(y[474]), .B(x[474]), .Z(n10555) );
  XNOR U12921 ( .A(n10556), .B(n10557), .Z(n10554) );
  XNOR U12922 ( .A(y[475]), .B(x[475]), .Z(n10557) );
  XNOR U12923 ( .A(y[476]), .B(x[476]), .Z(n10556) );
  XNOR U12924 ( .A(n10548), .B(n10549), .Z(n10559) );
  XNOR U12925 ( .A(y[471]), .B(x[471]), .Z(n10549) );
  XNOR U12926 ( .A(n10550), .B(n10551), .Z(n10548) );
  XNOR U12927 ( .A(y[472]), .B(x[472]), .Z(n10551) );
  XNOR U12928 ( .A(y[473]), .B(x[473]), .Z(n10550) );
  NAND U12929 ( .A(n10615), .B(n10616), .Z(N12994) );
  NANDN U12930 ( .A(n10617), .B(n10618), .Z(n10616) );
  OR U12931 ( .A(n10619), .B(n10620), .Z(n10618) );
  NAND U12932 ( .A(n10619), .B(n10620), .Z(n10615) );
  XOR U12933 ( .A(n10619), .B(n10621), .Z(N12993) );
  XNOR U12934 ( .A(n10617), .B(n10620), .Z(n10621) );
  AND U12935 ( .A(n10622), .B(n10623), .Z(n10620) );
  NANDN U12936 ( .A(n10624), .B(n10625), .Z(n10623) );
  NANDN U12937 ( .A(n10626), .B(n10627), .Z(n10625) );
  NANDN U12938 ( .A(n10627), .B(n10626), .Z(n10622) );
  NAND U12939 ( .A(n10628), .B(n10629), .Z(n10617) );
  NANDN U12940 ( .A(n10630), .B(n10631), .Z(n10629) );
  OR U12941 ( .A(n10632), .B(n10633), .Z(n10631) );
  NAND U12942 ( .A(n10633), .B(n10632), .Z(n10628) );
  AND U12943 ( .A(n10634), .B(n10635), .Z(n10619) );
  NANDN U12944 ( .A(n10636), .B(n10637), .Z(n10635) );
  NANDN U12945 ( .A(n10638), .B(n10639), .Z(n10637) );
  NANDN U12946 ( .A(n10639), .B(n10638), .Z(n10634) );
  XOR U12947 ( .A(n10633), .B(n10640), .Z(N12992) );
  XOR U12948 ( .A(n10630), .B(n10632), .Z(n10640) );
  XNOR U12949 ( .A(n10626), .B(n10641), .Z(n10632) );
  XNOR U12950 ( .A(n10624), .B(n10627), .Z(n10641) );
  NAND U12951 ( .A(n10642), .B(n10643), .Z(n10627) );
  NAND U12952 ( .A(n10644), .B(n10645), .Z(n10643) );
  OR U12953 ( .A(n10646), .B(n10647), .Z(n10644) );
  NANDN U12954 ( .A(n10648), .B(n10646), .Z(n10642) );
  IV U12955 ( .A(n10647), .Z(n10648) );
  NAND U12956 ( .A(n10649), .B(n10650), .Z(n10624) );
  NAND U12957 ( .A(n10651), .B(n10652), .Z(n10650) );
  NANDN U12958 ( .A(n10653), .B(n10654), .Z(n10651) );
  NANDN U12959 ( .A(n10654), .B(n10653), .Z(n10649) );
  AND U12960 ( .A(n10655), .B(n10656), .Z(n10626) );
  NAND U12961 ( .A(n10657), .B(n10658), .Z(n10656) );
  OR U12962 ( .A(n10659), .B(n10660), .Z(n10657) );
  NANDN U12963 ( .A(n10661), .B(n10659), .Z(n10655) );
  NAND U12964 ( .A(n10662), .B(n10663), .Z(n10630) );
  NANDN U12965 ( .A(n10664), .B(n10665), .Z(n10663) );
  OR U12966 ( .A(n10666), .B(n10667), .Z(n10665) );
  NANDN U12967 ( .A(n10668), .B(n10666), .Z(n10662) );
  IV U12968 ( .A(n10667), .Z(n10668) );
  XNOR U12969 ( .A(n10638), .B(n10669), .Z(n10633) );
  XNOR U12970 ( .A(n10636), .B(n10639), .Z(n10669) );
  NAND U12971 ( .A(n10670), .B(n10671), .Z(n10639) );
  NAND U12972 ( .A(n10672), .B(n10673), .Z(n10671) );
  OR U12973 ( .A(n10674), .B(n10675), .Z(n10672) );
  NANDN U12974 ( .A(n10676), .B(n10674), .Z(n10670) );
  IV U12975 ( .A(n10675), .Z(n10676) );
  NAND U12976 ( .A(n10677), .B(n10678), .Z(n10636) );
  NAND U12977 ( .A(n10679), .B(n10680), .Z(n10678) );
  NANDN U12978 ( .A(n10681), .B(n10682), .Z(n10679) );
  NANDN U12979 ( .A(n10682), .B(n10681), .Z(n10677) );
  AND U12980 ( .A(n10683), .B(n10684), .Z(n10638) );
  NAND U12981 ( .A(n10685), .B(n10686), .Z(n10684) );
  OR U12982 ( .A(n10687), .B(n10688), .Z(n10685) );
  NANDN U12983 ( .A(n10689), .B(n10687), .Z(n10683) );
  XNOR U12984 ( .A(n10664), .B(n10690), .Z(N12991) );
  XOR U12985 ( .A(n10666), .B(n10667), .Z(n10690) );
  XNOR U12986 ( .A(n10680), .B(n10691), .Z(n10667) );
  XOR U12987 ( .A(n10681), .B(n10682), .Z(n10691) );
  XOR U12988 ( .A(n10687), .B(n10692), .Z(n10682) );
  XOR U12989 ( .A(n10686), .B(n10689), .Z(n10692) );
  IV U12990 ( .A(n10688), .Z(n10689) );
  NAND U12991 ( .A(n10693), .B(n10694), .Z(n10688) );
  OR U12992 ( .A(n10695), .B(n10696), .Z(n10694) );
  OR U12993 ( .A(n10697), .B(n10698), .Z(n10693) );
  NAND U12994 ( .A(n10699), .B(n10700), .Z(n10686) );
  OR U12995 ( .A(n10701), .B(n10702), .Z(n10700) );
  OR U12996 ( .A(n10703), .B(n10704), .Z(n10699) );
  NOR U12997 ( .A(n10705), .B(n10706), .Z(n10687) );
  ANDN U12998 ( .B(n10707), .A(n10708), .Z(n10681) );
  XNOR U12999 ( .A(n10674), .B(n10709), .Z(n10680) );
  XNOR U13000 ( .A(n10673), .B(n10675), .Z(n10709) );
  NAND U13001 ( .A(n10710), .B(n10711), .Z(n10675) );
  OR U13002 ( .A(n10712), .B(n10713), .Z(n10711) );
  OR U13003 ( .A(n10714), .B(n10715), .Z(n10710) );
  NAND U13004 ( .A(n10716), .B(n10717), .Z(n10673) );
  OR U13005 ( .A(n10718), .B(n10719), .Z(n10717) );
  OR U13006 ( .A(n10720), .B(n10721), .Z(n10716) );
  ANDN U13007 ( .B(n10722), .A(n10723), .Z(n10674) );
  IV U13008 ( .A(n10724), .Z(n10722) );
  ANDN U13009 ( .B(n10725), .A(n10726), .Z(n10666) );
  XOR U13010 ( .A(n10652), .B(n10727), .Z(n10664) );
  XOR U13011 ( .A(n10653), .B(n10654), .Z(n10727) );
  XOR U13012 ( .A(n10659), .B(n10728), .Z(n10654) );
  XOR U13013 ( .A(n10658), .B(n10661), .Z(n10728) );
  IV U13014 ( .A(n10660), .Z(n10661) );
  NAND U13015 ( .A(n10729), .B(n10730), .Z(n10660) );
  OR U13016 ( .A(n10731), .B(n10732), .Z(n10730) );
  OR U13017 ( .A(n10733), .B(n10734), .Z(n10729) );
  NAND U13018 ( .A(n10735), .B(n10736), .Z(n10658) );
  OR U13019 ( .A(n10737), .B(n10738), .Z(n10736) );
  OR U13020 ( .A(n10739), .B(n10740), .Z(n10735) );
  NOR U13021 ( .A(n10741), .B(n10742), .Z(n10659) );
  ANDN U13022 ( .B(n10743), .A(n10744), .Z(n10653) );
  IV U13023 ( .A(n10745), .Z(n10743) );
  XNOR U13024 ( .A(n10646), .B(n10746), .Z(n10652) );
  XNOR U13025 ( .A(n10645), .B(n10647), .Z(n10746) );
  NAND U13026 ( .A(n10747), .B(n10748), .Z(n10647) );
  OR U13027 ( .A(n10749), .B(n10750), .Z(n10748) );
  OR U13028 ( .A(n10751), .B(n10752), .Z(n10747) );
  NAND U13029 ( .A(n10753), .B(n10754), .Z(n10645) );
  OR U13030 ( .A(n10755), .B(n10756), .Z(n10754) );
  OR U13031 ( .A(n10757), .B(n10758), .Z(n10753) );
  ANDN U13032 ( .B(n10759), .A(n10760), .Z(n10646) );
  IV U13033 ( .A(n10761), .Z(n10759) );
  XNOR U13034 ( .A(n10726), .B(n10725), .Z(N12990) );
  XOR U13035 ( .A(n10745), .B(n10744), .Z(n10725) );
  XNOR U13036 ( .A(n10760), .B(n10761), .Z(n10744) );
  XNOR U13037 ( .A(n10755), .B(n10756), .Z(n10761) );
  XNOR U13038 ( .A(n10757), .B(n10758), .Z(n10756) );
  XNOR U13039 ( .A(y[469]), .B(x[469]), .Z(n10758) );
  XNOR U13040 ( .A(y[470]), .B(x[470]), .Z(n10757) );
  XNOR U13041 ( .A(y[468]), .B(x[468]), .Z(n10755) );
  XNOR U13042 ( .A(n10749), .B(n10750), .Z(n10760) );
  XNOR U13043 ( .A(y[465]), .B(x[465]), .Z(n10750) );
  XNOR U13044 ( .A(n10751), .B(n10752), .Z(n10749) );
  XNOR U13045 ( .A(y[466]), .B(x[466]), .Z(n10752) );
  XNOR U13046 ( .A(y[467]), .B(x[467]), .Z(n10751) );
  XNOR U13047 ( .A(n10742), .B(n10741), .Z(n10745) );
  XNOR U13048 ( .A(n10737), .B(n10738), .Z(n10741) );
  XNOR U13049 ( .A(y[462]), .B(x[462]), .Z(n10738) );
  XNOR U13050 ( .A(n10739), .B(n10740), .Z(n10737) );
  XNOR U13051 ( .A(y[463]), .B(x[463]), .Z(n10740) );
  XNOR U13052 ( .A(y[464]), .B(x[464]), .Z(n10739) );
  XNOR U13053 ( .A(n10731), .B(n10732), .Z(n10742) );
  XNOR U13054 ( .A(y[459]), .B(x[459]), .Z(n10732) );
  XNOR U13055 ( .A(n10733), .B(n10734), .Z(n10731) );
  XNOR U13056 ( .A(y[460]), .B(x[460]), .Z(n10734) );
  XNOR U13057 ( .A(y[461]), .B(x[461]), .Z(n10733) );
  XOR U13058 ( .A(n10707), .B(n10708), .Z(n10726) );
  XNOR U13059 ( .A(n10723), .B(n10724), .Z(n10708) );
  XNOR U13060 ( .A(n10718), .B(n10719), .Z(n10724) );
  XNOR U13061 ( .A(n10720), .B(n10721), .Z(n10719) );
  XNOR U13062 ( .A(y[457]), .B(x[457]), .Z(n10721) );
  XNOR U13063 ( .A(y[458]), .B(x[458]), .Z(n10720) );
  XNOR U13064 ( .A(y[456]), .B(x[456]), .Z(n10718) );
  XNOR U13065 ( .A(n10712), .B(n10713), .Z(n10723) );
  XNOR U13066 ( .A(y[453]), .B(x[453]), .Z(n10713) );
  XNOR U13067 ( .A(n10714), .B(n10715), .Z(n10712) );
  XNOR U13068 ( .A(y[454]), .B(x[454]), .Z(n10715) );
  XNOR U13069 ( .A(y[455]), .B(x[455]), .Z(n10714) );
  XOR U13070 ( .A(n10706), .B(n10705), .Z(n10707) );
  XNOR U13071 ( .A(n10701), .B(n10702), .Z(n10705) );
  XNOR U13072 ( .A(y[450]), .B(x[450]), .Z(n10702) );
  XNOR U13073 ( .A(n10703), .B(n10704), .Z(n10701) );
  XNOR U13074 ( .A(y[451]), .B(x[451]), .Z(n10704) );
  XNOR U13075 ( .A(y[452]), .B(x[452]), .Z(n10703) );
  XNOR U13076 ( .A(n10695), .B(n10696), .Z(n10706) );
  XNOR U13077 ( .A(y[447]), .B(x[447]), .Z(n10696) );
  XNOR U13078 ( .A(n10697), .B(n10698), .Z(n10695) );
  XNOR U13079 ( .A(y[448]), .B(x[448]), .Z(n10698) );
  XNOR U13080 ( .A(y[449]), .B(x[449]), .Z(n10697) );
  NAND U13081 ( .A(n10762), .B(n10763), .Z(N12983) );
  NANDN U13082 ( .A(n10764), .B(n10765), .Z(n10763) );
  OR U13083 ( .A(n10766), .B(n10767), .Z(n10765) );
  NAND U13084 ( .A(n10766), .B(n10767), .Z(n10762) );
  XOR U13085 ( .A(n10766), .B(n10768), .Z(N12982) );
  XNOR U13086 ( .A(n10764), .B(n10767), .Z(n10768) );
  AND U13087 ( .A(n10769), .B(n10770), .Z(n10767) );
  NANDN U13088 ( .A(n10771), .B(n10772), .Z(n10770) );
  NANDN U13089 ( .A(n10773), .B(n10774), .Z(n10772) );
  NANDN U13090 ( .A(n10774), .B(n10773), .Z(n10769) );
  NAND U13091 ( .A(n10775), .B(n10776), .Z(n10764) );
  NANDN U13092 ( .A(n10777), .B(n10778), .Z(n10776) );
  OR U13093 ( .A(n10779), .B(n10780), .Z(n10778) );
  NAND U13094 ( .A(n10780), .B(n10779), .Z(n10775) );
  AND U13095 ( .A(n10781), .B(n10782), .Z(n10766) );
  NANDN U13096 ( .A(n10783), .B(n10784), .Z(n10782) );
  NANDN U13097 ( .A(n10785), .B(n10786), .Z(n10784) );
  NANDN U13098 ( .A(n10786), .B(n10785), .Z(n10781) );
  XOR U13099 ( .A(n10780), .B(n10787), .Z(N12981) );
  XOR U13100 ( .A(n10777), .B(n10779), .Z(n10787) );
  XNOR U13101 ( .A(n10773), .B(n10788), .Z(n10779) );
  XNOR U13102 ( .A(n10771), .B(n10774), .Z(n10788) );
  NAND U13103 ( .A(n10789), .B(n10790), .Z(n10774) );
  NAND U13104 ( .A(n10791), .B(n10792), .Z(n10790) );
  OR U13105 ( .A(n10793), .B(n10794), .Z(n10791) );
  NANDN U13106 ( .A(n10795), .B(n10793), .Z(n10789) );
  IV U13107 ( .A(n10794), .Z(n10795) );
  NAND U13108 ( .A(n10796), .B(n10797), .Z(n10771) );
  NAND U13109 ( .A(n10798), .B(n10799), .Z(n10797) );
  NANDN U13110 ( .A(n10800), .B(n10801), .Z(n10798) );
  NANDN U13111 ( .A(n10801), .B(n10800), .Z(n10796) );
  AND U13112 ( .A(n10802), .B(n10803), .Z(n10773) );
  NAND U13113 ( .A(n10804), .B(n10805), .Z(n10803) );
  OR U13114 ( .A(n10806), .B(n10807), .Z(n10804) );
  NANDN U13115 ( .A(n10808), .B(n10806), .Z(n10802) );
  NAND U13116 ( .A(n10809), .B(n10810), .Z(n10777) );
  NANDN U13117 ( .A(n10811), .B(n10812), .Z(n10810) );
  OR U13118 ( .A(n10813), .B(n10814), .Z(n10812) );
  NANDN U13119 ( .A(n10815), .B(n10813), .Z(n10809) );
  IV U13120 ( .A(n10814), .Z(n10815) );
  XNOR U13121 ( .A(n10785), .B(n10816), .Z(n10780) );
  XNOR U13122 ( .A(n10783), .B(n10786), .Z(n10816) );
  NAND U13123 ( .A(n10817), .B(n10818), .Z(n10786) );
  NAND U13124 ( .A(n10819), .B(n10820), .Z(n10818) );
  OR U13125 ( .A(n10821), .B(n10822), .Z(n10819) );
  NANDN U13126 ( .A(n10823), .B(n10821), .Z(n10817) );
  IV U13127 ( .A(n10822), .Z(n10823) );
  NAND U13128 ( .A(n10824), .B(n10825), .Z(n10783) );
  NAND U13129 ( .A(n10826), .B(n10827), .Z(n10825) );
  NANDN U13130 ( .A(n10828), .B(n10829), .Z(n10826) );
  NANDN U13131 ( .A(n10829), .B(n10828), .Z(n10824) );
  AND U13132 ( .A(n10830), .B(n10831), .Z(n10785) );
  NAND U13133 ( .A(n10832), .B(n10833), .Z(n10831) );
  OR U13134 ( .A(n10834), .B(n10835), .Z(n10832) );
  NANDN U13135 ( .A(n10836), .B(n10834), .Z(n10830) );
  XNOR U13136 ( .A(n10811), .B(n10837), .Z(N12980) );
  XOR U13137 ( .A(n10813), .B(n10814), .Z(n10837) );
  XNOR U13138 ( .A(n10827), .B(n10838), .Z(n10814) );
  XOR U13139 ( .A(n10828), .B(n10829), .Z(n10838) );
  XOR U13140 ( .A(n10834), .B(n10839), .Z(n10829) );
  XOR U13141 ( .A(n10833), .B(n10836), .Z(n10839) );
  IV U13142 ( .A(n10835), .Z(n10836) );
  NAND U13143 ( .A(n10840), .B(n10841), .Z(n10835) );
  OR U13144 ( .A(n10842), .B(n10843), .Z(n10841) );
  OR U13145 ( .A(n10844), .B(n10845), .Z(n10840) );
  NAND U13146 ( .A(n10846), .B(n10847), .Z(n10833) );
  OR U13147 ( .A(n10848), .B(n10849), .Z(n10847) );
  OR U13148 ( .A(n10850), .B(n10851), .Z(n10846) );
  NOR U13149 ( .A(n10852), .B(n10853), .Z(n10834) );
  ANDN U13150 ( .B(n10854), .A(n10855), .Z(n10828) );
  XNOR U13151 ( .A(n10821), .B(n10856), .Z(n10827) );
  XNOR U13152 ( .A(n10820), .B(n10822), .Z(n10856) );
  NAND U13153 ( .A(n10857), .B(n10858), .Z(n10822) );
  OR U13154 ( .A(n10859), .B(n10860), .Z(n10858) );
  OR U13155 ( .A(n10861), .B(n10862), .Z(n10857) );
  NAND U13156 ( .A(n10863), .B(n10864), .Z(n10820) );
  OR U13157 ( .A(n10865), .B(n10866), .Z(n10864) );
  OR U13158 ( .A(n10867), .B(n10868), .Z(n10863) );
  ANDN U13159 ( .B(n10869), .A(n10870), .Z(n10821) );
  IV U13160 ( .A(n10871), .Z(n10869) );
  ANDN U13161 ( .B(n10872), .A(n10873), .Z(n10813) );
  XOR U13162 ( .A(n10799), .B(n10874), .Z(n10811) );
  XOR U13163 ( .A(n10800), .B(n10801), .Z(n10874) );
  XOR U13164 ( .A(n10806), .B(n10875), .Z(n10801) );
  XOR U13165 ( .A(n10805), .B(n10808), .Z(n10875) );
  IV U13166 ( .A(n10807), .Z(n10808) );
  NAND U13167 ( .A(n10876), .B(n10877), .Z(n10807) );
  OR U13168 ( .A(n10878), .B(n10879), .Z(n10877) );
  OR U13169 ( .A(n10880), .B(n10881), .Z(n10876) );
  NAND U13170 ( .A(n10882), .B(n10883), .Z(n10805) );
  OR U13171 ( .A(n10884), .B(n10885), .Z(n10883) );
  OR U13172 ( .A(n10886), .B(n10887), .Z(n10882) );
  NOR U13173 ( .A(n10888), .B(n10889), .Z(n10806) );
  ANDN U13174 ( .B(n10890), .A(n10891), .Z(n10800) );
  IV U13175 ( .A(n10892), .Z(n10890) );
  XNOR U13176 ( .A(n10793), .B(n10893), .Z(n10799) );
  XNOR U13177 ( .A(n10792), .B(n10794), .Z(n10893) );
  NAND U13178 ( .A(n10894), .B(n10895), .Z(n10794) );
  OR U13179 ( .A(n10896), .B(n10897), .Z(n10895) );
  OR U13180 ( .A(n10898), .B(n10899), .Z(n10894) );
  NAND U13181 ( .A(n10900), .B(n10901), .Z(n10792) );
  OR U13182 ( .A(n10902), .B(n10903), .Z(n10901) );
  OR U13183 ( .A(n10904), .B(n10905), .Z(n10900) );
  ANDN U13184 ( .B(n10906), .A(n10907), .Z(n10793) );
  IV U13185 ( .A(n10908), .Z(n10906) );
  XNOR U13186 ( .A(n10873), .B(n10872), .Z(N12979) );
  XOR U13187 ( .A(n10892), .B(n10891), .Z(n10872) );
  XNOR U13188 ( .A(n10907), .B(n10908), .Z(n10891) );
  XNOR U13189 ( .A(n10902), .B(n10903), .Z(n10908) );
  XNOR U13190 ( .A(n10904), .B(n10905), .Z(n10903) );
  XNOR U13191 ( .A(y[445]), .B(x[445]), .Z(n10905) );
  XNOR U13192 ( .A(y[446]), .B(x[446]), .Z(n10904) );
  XNOR U13193 ( .A(y[444]), .B(x[444]), .Z(n10902) );
  XNOR U13194 ( .A(n10896), .B(n10897), .Z(n10907) );
  XNOR U13195 ( .A(y[441]), .B(x[441]), .Z(n10897) );
  XNOR U13196 ( .A(n10898), .B(n10899), .Z(n10896) );
  XNOR U13197 ( .A(y[442]), .B(x[442]), .Z(n10899) );
  XNOR U13198 ( .A(y[443]), .B(x[443]), .Z(n10898) );
  XNOR U13199 ( .A(n10889), .B(n10888), .Z(n10892) );
  XNOR U13200 ( .A(n10884), .B(n10885), .Z(n10888) );
  XNOR U13201 ( .A(y[438]), .B(x[438]), .Z(n10885) );
  XNOR U13202 ( .A(n10886), .B(n10887), .Z(n10884) );
  XNOR U13203 ( .A(y[439]), .B(x[439]), .Z(n10887) );
  XNOR U13204 ( .A(y[440]), .B(x[440]), .Z(n10886) );
  XNOR U13205 ( .A(n10878), .B(n10879), .Z(n10889) );
  XNOR U13206 ( .A(y[435]), .B(x[435]), .Z(n10879) );
  XNOR U13207 ( .A(n10880), .B(n10881), .Z(n10878) );
  XNOR U13208 ( .A(y[436]), .B(x[436]), .Z(n10881) );
  XNOR U13209 ( .A(y[437]), .B(x[437]), .Z(n10880) );
  XOR U13210 ( .A(n10854), .B(n10855), .Z(n10873) );
  XNOR U13211 ( .A(n10870), .B(n10871), .Z(n10855) );
  XNOR U13212 ( .A(n10865), .B(n10866), .Z(n10871) );
  XNOR U13213 ( .A(n10867), .B(n10868), .Z(n10866) );
  XNOR U13214 ( .A(y[433]), .B(x[433]), .Z(n10868) );
  XNOR U13215 ( .A(y[434]), .B(x[434]), .Z(n10867) );
  XNOR U13216 ( .A(y[432]), .B(x[432]), .Z(n10865) );
  XNOR U13217 ( .A(n10859), .B(n10860), .Z(n10870) );
  XNOR U13218 ( .A(y[429]), .B(x[429]), .Z(n10860) );
  XNOR U13219 ( .A(n10861), .B(n10862), .Z(n10859) );
  XNOR U13220 ( .A(y[430]), .B(x[430]), .Z(n10862) );
  XNOR U13221 ( .A(y[431]), .B(x[431]), .Z(n10861) );
  XOR U13222 ( .A(n10853), .B(n10852), .Z(n10854) );
  XNOR U13223 ( .A(n10848), .B(n10849), .Z(n10852) );
  XNOR U13224 ( .A(y[426]), .B(x[426]), .Z(n10849) );
  XNOR U13225 ( .A(n10850), .B(n10851), .Z(n10848) );
  XNOR U13226 ( .A(y[427]), .B(x[427]), .Z(n10851) );
  XNOR U13227 ( .A(y[428]), .B(x[428]), .Z(n10850) );
  XNOR U13228 ( .A(n10842), .B(n10843), .Z(n10853) );
  XNOR U13229 ( .A(y[423]), .B(x[423]), .Z(n10843) );
  XNOR U13230 ( .A(n10844), .B(n10845), .Z(n10842) );
  XNOR U13231 ( .A(y[424]), .B(x[424]), .Z(n10845) );
  XNOR U13232 ( .A(y[425]), .B(x[425]), .Z(n10844) );
  NAND U13233 ( .A(n10909), .B(n10910), .Z(N12972) );
  NANDN U13234 ( .A(n10911), .B(n10912), .Z(n10910) );
  OR U13235 ( .A(n10913), .B(n10914), .Z(n10912) );
  NAND U13236 ( .A(n10913), .B(n10914), .Z(n10909) );
  XOR U13237 ( .A(n10913), .B(n10915), .Z(N12971) );
  XNOR U13238 ( .A(n10911), .B(n10914), .Z(n10915) );
  AND U13239 ( .A(n10916), .B(n10917), .Z(n10914) );
  NANDN U13240 ( .A(n10918), .B(n10919), .Z(n10917) );
  NANDN U13241 ( .A(n10920), .B(n10921), .Z(n10919) );
  NANDN U13242 ( .A(n10921), .B(n10920), .Z(n10916) );
  NAND U13243 ( .A(n10922), .B(n10923), .Z(n10911) );
  NANDN U13244 ( .A(n10924), .B(n10925), .Z(n10923) );
  OR U13245 ( .A(n10926), .B(n10927), .Z(n10925) );
  NAND U13246 ( .A(n10927), .B(n10926), .Z(n10922) );
  AND U13247 ( .A(n10928), .B(n10929), .Z(n10913) );
  NANDN U13248 ( .A(n10930), .B(n10931), .Z(n10929) );
  NANDN U13249 ( .A(n10932), .B(n10933), .Z(n10931) );
  NANDN U13250 ( .A(n10933), .B(n10932), .Z(n10928) );
  XOR U13251 ( .A(n10927), .B(n10934), .Z(N12970) );
  XOR U13252 ( .A(n10924), .B(n10926), .Z(n10934) );
  XNOR U13253 ( .A(n10920), .B(n10935), .Z(n10926) );
  XNOR U13254 ( .A(n10918), .B(n10921), .Z(n10935) );
  NAND U13255 ( .A(n10936), .B(n10937), .Z(n10921) );
  NAND U13256 ( .A(n10938), .B(n10939), .Z(n10937) );
  OR U13257 ( .A(n10940), .B(n10941), .Z(n10938) );
  NANDN U13258 ( .A(n10942), .B(n10940), .Z(n10936) );
  IV U13259 ( .A(n10941), .Z(n10942) );
  NAND U13260 ( .A(n10943), .B(n10944), .Z(n10918) );
  NAND U13261 ( .A(n10945), .B(n10946), .Z(n10944) );
  NANDN U13262 ( .A(n10947), .B(n10948), .Z(n10945) );
  NANDN U13263 ( .A(n10948), .B(n10947), .Z(n10943) );
  AND U13264 ( .A(n10949), .B(n10950), .Z(n10920) );
  NAND U13265 ( .A(n10951), .B(n10952), .Z(n10950) );
  OR U13266 ( .A(n10953), .B(n10954), .Z(n10951) );
  NANDN U13267 ( .A(n10955), .B(n10953), .Z(n10949) );
  NAND U13268 ( .A(n10956), .B(n10957), .Z(n10924) );
  NANDN U13269 ( .A(n10958), .B(n10959), .Z(n10957) );
  OR U13270 ( .A(n10960), .B(n10961), .Z(n10959) );
  NANDN U13271 ( .A(n10962), .B(n10960), .Z(n10956) );
  IV U13272 ( .A(n10961), .Z(n10962) );
  XNOR U13273 ( .A(n10932), .B(n10963), .Z(n10927) );
  XNOR U13274 ( .A(n10930), .B(n10933), .Z(n10963) );
  NAND U13275 ( .A(n10964), .B(n10965), .Z(n10933) );
  NAND U13276 ( .A(n10966), .B(n10967), .Z(n10965) );
  OR U13277 ( .A(n10968), .B(n10969), .Z(n10966) );
  NANDN U13278 ( .A(n10970), .B(n10968), .Z(n10964) );
  IV U13279 ( .A(n10969), .Z(n10970) );
  NAND U13280 ( .A(n10971), .B(n10972), .Z(n10930) );
  NAND U13281 ( .A(n10973), .B(n10974), .Z(n10972) );
  NANDN U13282 ( .A(n10975), .B(n10976), .Z(n10973) );
  NANDN U13283 ( .A(n10976), .B(n10975), .Z(n10971) );
  AND U13284 ( .A(n10977), .B(n10978), .Z(n10932) );
  NAND U13285 ( .A(n10979), .B(n10980), .Z(n10978) );
  OR U13286 ( .A(n10981), .B(n10982), .Z(n10979) );
  NANDN U13287 ( .A(n10983), .B(n10981), .Z(n10977) );
  XNOR U13288 ( .A(n10958), .B(n10984), .Z(N12969) );
  XOR U13289 ( .A(n10960), .B(n10961), .Z(n10984) );
  XNOR U13290 ( .A(n10974), .B(n10985), .Z(n10961) );
  XOR U13291 ( .A(n10975), .B(n10976), .Z(n10985) );
  XOR U13292 ( .A(n10981), .B(n10986), .Z(n10976) );
  XOR U13293 ( .A(n10980), .B(n10983), .Z(n10986) );
  IV U13294 ( .A(n10982), .Z(n10983) );
  NAND U13295 ( .A(n10987), .B(n10988), .Z(n10982) );
  OR U13296 ( .A(n10989), .B(n10990), .Z(n10988) );
  OR U13297 ( .A(n10991), .B(n10992), .Z(n10987) );
  NAND U13298 ( .A(n10993), .B(n10994), .Z(n10980) );
  OR U13299 ( .A(n10995), .B(n10996), .Z(n10994) );
  OR U13300 ( .A(n10997), .B(n10998), .Z(n10993) );
  NOR U13301 ( .A(n10999), .B(n11000), .Z(n10981) );
  ANDN U13302 ( .B(n11001), .A(n11002), .Z(n10975) );
  XNOR U13303 ( .A(n10968), .B(n11003), .Z(n10974) );
  XNOR U13304 ( .A(n10967), .B(n10969), .Z(n11003) );
  NAND U13305 ( .A(n11004), .B(n11005), .Z(n10969) );
  OR U13306 ( .A(n11006), .B(n11007), .Z(n11005) );
  OR U13307 ( .A(n11008), .B(n11009), .Z(n11004) );
  NAND U13308 ( .A(n11010), .B(n11011), .Z(n10967) );
  OR U13309 ( .A(n11012), .B(n11013), .Z(n11011) );
  OR U13310 ( .A(n11014), .B(n11015), .Z(n11010) );
  ANDN U13311 ( .B(n11016), .A(n11017), .Z(n10968) );
  IV U13312 ( .A(n11018), .Z(n11016) );
  ANDN U13313 ( .B(n11019), .A(n11020), .Z(n10960) );
  XOR U13314 ( .A(n10946), .B(n11021), .Z(n10958) );
  XOR U13315 ( .A(n10947), .B(n10948), .Z(n11021) );
  XOR U13316 ( .A(n10953), .B(n11022), .Z(n10948) );
  XOR U13317 ( .A(n10952), .B(n10955), .Z(n11022) );
  IV U13318 ( .A(n10954), .Z(n10955) );
  NAND U13319 ( .A(n11023), .B(n11024), .Z(n10954) );
  OR U13320 ( .A(n11025), .B(n11026), .Z(n11024) );
  OR U13321 ( .A(n11027), .B(n11028), .Z(n11023) );
  NAND U13322 ( .A(n11029), .B(n11030), .Z(n10952) );
  OR U13323 ( .A(n11031), .B(n11032), .Z(n11030) );
  OR U13324 ( .A(n11033), .B(n11034), .Z(n11029) );
  NOR U13325 ( .A(n11035), .B(n11036), .Z(n10953) );
  ANDN U13326 ( .B(n11037), .A(n11038), .Z(n10947) );
  IV U13327 ( .A(n11039), .Z(n11037) );
  XNOR U13328 ( .A(n10940), .B(n11040), .Z(n10946) );
  XNOR U13329 ( .A(n10939), .B(n10941), .Z(n11040) );
  NAND U13330 ( .A(n11041), .B(n11042), .Z(n10941) );
  OR U13331 ( .A(n11043), .B(n11044), .Z(n11042) );
  OR U13332 ( .A(n11045), .B(n11046), .Z(n11041) );
  NAND U13333 ( .A(n11047), .B(n11048), .Z(n10939) );
  OR U13334 ( .A(n11049), .B(n11050), .Z(n11048) );
  OR U13335 ( .A(n11051), .B(n11052), .Z(n11047) );
  ANDN U13336 ( .B(n11053), .A(n11054), .Z(n10940) );
  IV U13337 ( .A(n11055), .Z(n11053) );
  XNOR U13338 ( .A(n11020), .B(n11019), .Z(N12968) );
  XOR U13339 ( .A(n11039), .B(n11038), .Z(n11019) );
  XNOR U13340 ( .A(n11054), .B(n11055), .Z(n11038) );
  XNOR U13341 ( .A(n11049), .B(n11050), .Z(n11055) );
  XNOR U13342 ( .A(n11051), .B(n11052), .Z(n11050) );
  XNOR U13343 ( .A(y[421]), .B(x[421]), .Z(n11052) );
  XNOR U13344 ( .A(y[422]), .B(x[422]), .Z(n11051) );
  XNOR U13345 ( .A(y[420]), .B(x[420]), .Z(n11049) );
  XNOR U13346 ( .A(n11043), .B(n11044), .Z(n11054) );
  XNOR U13347 ( .A(y[417]), .B(x[417]), .Z(n11044) );
  XNOR U13348 ( .A(n11045), .B(n11046), .Z(n11043) );
  XNOR U13349 ( .A(y[418]), .B(x[418]), .Z(n11046) );
  XNOR U13350 ( .A(y[419]), .B(x[419]), .Z(n11045) );
  XNOR U13351 ( .A(n11036), .B(n11035), .Z(n11039) );
  XNOR U13352 ( .A(n11031), .B(n11032), .Z(n11035) );
  XNOR U13353 ( .A(y[414]), .B(x[414]), .Z(n11032) );
  XNOR U13354 ( .A(n11033), .B(n11034), .Z(n11031) );
  XNOR U13355 ( .A(y[415]), .B(x[415]), .Z(n11034) );
  XNOR U13356 ( .A(y[416]), .B(x[416]), .Z(n11033) );
  XNOR U13357 ( .A(n11025), .B(n11026), .Z(n11036) );
  XNOR U13358 ( .A(y[411]), .B(x[411]), .Z(n11026) );
  XNOR U13359 ( .A(n11027), .B(n11028), .Z(n11025) );
  XNOR U13360 ( .A(y[412]), .B(x[412]), .Z(n11028) );
  XNOR U13361 ( .A(y[413]), .B(x[413]), .Z(n11027) );
  XOR U13362 ( .A(n11001), .B(n11002), .Z(n11020) );
  XNOR U13363 ( .A(n11017), .B(n11018), .Z(n11002) );
  XNOR U13364 ( .A(n11012), .B(n11013), .Z(n11018) );
  XNOR U13365 ( .A(n11014), .B(n11015), .Z(n11013) );
  XNOR U13366 ( .A(y[409]), .B(x[409]), .Z(n11015) );
  XNOR U13367 ( .A(y[410]), .B(x[410]), .Z(n11014) );
  XNOR U13368 ( .A(y[408]), .B(x[408]), .Z(n11012) );
  XNOR U13369 ( .A(n11006), .B(n11007), .Z(n11017) );
  XNOR U13370 ( .A(y[405]), .B(x[405]), .Z(n11007) );
  XNOR U13371 ( .A(n11008), .B(n11009), .Z(n11006) );
  XNOR U13372 ( .A(y[406]), .B(x[406]), .Z(n11009) );
  XNOR U13373 ( .A(y[407]), .B(x[407]), .Z(n11008) );
  XOR U13374 ( .A(n11000), .B(n10999), .Z(n11001) );
  XNOR U13375 ( .A(n10995), .B(n10996), .Z(n10999) );
  XNOR U13376 ( .A(y[402]), .B(x[402]), .Z(n10996) );
  XNOR U13377 ( .A(n10997), .B(n10998), .Z(n10995) );
  XNOR U13378 ( .A(y[403]), .B(x[403]), .Z(n10998) );
  XNOR U13379 ( .A(y[404]), .B(x[404]), .Z(n10997) );
  XNOR U13380 ( .A(n10989), .B(n10990), .Z(n11000) );
  XNOR U13381 ( .A(y[399]), .B(x[399]), .Z(n10990) );
  XNOR U13382 ( .A(n10991), .B(n10992), .Z(n10989) );
  XNOR U13383 ( .A(y[400]), .B(x[400]), .Z(n10992) );
  XNOR U13384 ( .A(y[401]), .B(x[401]), .Z(n10991) );
  NAND U13385 ( .A(n11056), .B(n11057), .Z(N12961) );
  NANDN U13386 ( .A(n11058), .B(n11059), .Z(n11057) );
  OR U13387 ( .A(n11060), .B(n11061), .Z(n11059) );
  NAND U13388 ( .A(n11060), .B(n11061), .Z(n11056) );
  XOR U13389 ( .A(n11060), .B(n11062), .Z(N12960) );
  XNOR U13390 ( .A(n11058), .B(n11061), .Z(n11062) );
  AND U13391 ( .A(n11063), .B(n11064), .Z(n11061) );
  NANDN U13392 ( .A(n11065), .B(n11066), .Z(n11064) );
  NANDN U13393 ( .A(n11067), .B(n11068), .Z(n11066) );
  NANDN U13394 ( .A(n11068), .B(n11067), .Z(n11063) );
  NAND U13395 ( .A(n11069), .B(n11070), .Z(n11058) );
  NANDN U13396 ( .A(n11071), .B(n11072), .Z(n11070) );
  OR U13397 ( .A(n11073), .B(n11074), .Z(n11072) );
  NAND U13398 ( .A(n11074), .B(n11073), .Z(n11069) );
  AND U13399 ( .A(n11075), .B(n11076), .Z(n11060) );
  NANDN U13400 ( .A(n11077), .B(n11078), .Z(n11076) );
  NANDN U13401 ( .A(n11079), .B(n11080), .Z(n11078) );
  NANDN U13402 ( .A(n11080), .B(n11079), .Z(n11075) );
  XOR U13403 ( .A(n11074), .B(n11081), .Z(N12959) );
  XOR U13404 ( .A(n11071), .B(n11073), .Z(n11081) );
  XNOR U13405 ( .A(n11067), .B(n11082), .Z(n11073) );
  XNOR U13406 ( .A(n11065), .B(n11068), .Z(n11082) );
  NAND U13407 ( .A(n11083), .B(n11084), .Z(n11068) );
  NAND U13408 ( .A(n11085), .B(n11086), .Z(n11084) );
  OR U13409 ( .A(n11087), .B(n11088), .Z(n11085) );
  NANDN U13410 ( .A(n11089), .B(n11087), .Z(n11083) );
  IV U13411 ( .A(n11088), .Z(n11089) );
  NAND U13412 ( .A(n11090), .B(n11091), .Z(n11065) );
  NAND U13413 ( .A(n11092), .B(n11093), .Z(n11091) );
  NANDN U13414 ( .A(n11094), .B(n11095), .Z(n11092) );
  NANDN U13415 ( .A(n11095), .B(n11094), .Z(n11090) );
  AND U13416 ( .A(n11096), .B(n11097), .Z(n11067) );
  NAND U13417 ( .A(n11098), .B(n11099), .Z(n11097) );
  OR U13418 ( .A(n11100), .B(n11101), .Z(n11098) );
  NANDN U13419 ( .A(n11102), .B(n11100), .Z(n11096) );
  NAND U13420 ( .A(n11103), .B(n11104), .Z(n11071) );
  NANDN U13421 ( .A(n11105), .B(n11106), .Z(n11104) );
  OR U13422 ( .A(n11107), .B(n11108), .Z(n11106) );
  NANDN U13423 ( .A(n11109), .B(n11107), .Z(n11103) );
  IV U13424 ( .A(n11108), .Z(n11109) );
  XNOR U13425 ( .A(n11079), .B(n11110), .Z(n11074) );
  XNOR U13426 ( .A(n11077), .B(n11080), .Z(n11110) );
  NAND U13427 ( .A(n11111), .B(n11112), .Z(n11080) );
  NAND U13428 ( .A(n11113), .B(n11114), .Z(n11112) );
  OR U13429 ( .A(n11115), .B(n11116), .Z(n11113) );
  NANDN U13430 ( .A(n11117), .B(n11115), .Z(n11111) );
  IV U13431 ( .A(n11116), .Z(n11117) );
  NAND U13432 ( .A(n11118), .B(n11119), .Z(n11077) );
  NAND U13433 ( .A(n11120), .B(n11121), .Z(n11119) );
  NANDN U13434 ( .A(n11122), .B(n11123), .Z(n11120) );
  NANDN U13435 ( .A(n11123), .B(n11122), .Z(n11118) );
  AND U13436 ( .A(n11124), .B(n11125), .Z(n11079) );
  NAND U13437 ( .A(n11126), .B(n11127), .Z(n11125) );
  OR U13438 ( .A(n11128), .B(n11129), .Z(n11126) );
  NANDN U13439 ( .A(n11130), .B(n11128), .Z(n11124) );
  XNOR U13440 ( .A(n11105), .B(n11131), .Z(N12958) );
  XOR U13441 ( .A(n11107), .B(n11108), .Z(n11131) );
  XNOR U13442 ( .A(n11121), .B(n11132), .Z(n11108) );
  XOR U13443 ( .A(n11122), .B(n11123), .Z(n11132) );
  XOR U13444 ( .A(n11128), .B(n11133), .Z(n11123) );
  XOR U13445 ( .A(n11127), .B(n11130), .Z(n11133) );
  IV U13446 ( .A(n11129), .Z(n11130) );
  NAND U13447 ( .A(n11134), .B(n11135), .Z(n11129) );
  OR U13448 ( .A(n11136), .B(n11137), .Z(n11135) );
  OR U13449 ( .A(n11138), .B(n11139), .Z(n11134) );
  NAND U13450 ( .A(n11140), .B(n11141), .Z(n11127) );
  OR U13451 ( .A(n11142), .B(n11143), .Z(n11141) );
  OR U13452 ( .A(n11144), .B(n11145), .Z(n11140) );
  NOR U13453 ( .A(n11146), .B(n11147), .Z(n11128) );
  ANDN U13454 ( .B(n11148), .A(n11149), .Z(n11122) );
  XNOR U13455 ( .A(n11115), .B(n11150), .Z(n11121) );
  XNOR U13456 ( .A(n11114), .B(n11116), .Z(n11150) );
  NAND U13457 ( .A(n11151), .B(n11152), .Z(n11116) );
  OR U13458 ( .A(n11153), .B(n11154), .Z(n11152) );
  OR U13459 ( .A(n11155), .B(n11156), .Z(n11151) );
  NAND U13460 ( .A(n11157), .B(n11158), .Z(n11114) );
  OR U13461 ( .A(n11159), .B(n11160), .Z(n11158) );
  OR U13462 ( .A(n11161), .B(n11162), .Z(n11157) );
  ANDN U13463 ( .B(n11163), .A(n11164), .Z(n11115) );
  IV U13464 ( .A(n11165), .Z(n11163) );
  ANDN U13465 ( .B(n11166), .A(n11167), .Z(n11107) );
  XOR U13466 ( .A(n11093), .B(n11168), .Z(n11105) );
  XOR U13467 ( .A(n11094), .B(n11095), .Z(n11168) );
  XOR U13468 ( .A(n11100), .B(n11169), .Z(n11095) );
  XOR U13469 ( .A(n11099), .B(n11102), .Z(n11169) );
  IV U13470 ( .A(n11101), .Z(n11102) );
  NAND U13471 ( .A(n11170), .B(n11171), .Z(n11101) );
  OR U13472 ( .A(n11172), .B(n11173), .Z(n11171) );
  OR U13473 ( .A(n11174), .B(n11175), .Z(n11170) );
  NAND U13474 ( .A(n11176), .B(n11177), .Z(n11099) );
  OR U13475 ( .A(n11178), .B(n11179), .Z(n11177) );
  OR U13476 ( .A(n11180), .B(n11181), .Z(n11176) );
  NOR U13477 ( .A(n11182), .B(n11183), .Z(n11100) );
  ANDN U13478 ( .B(n11184), .A(n11185), .Z(n11094) );
  IV U13479 ( .A(n11186), .Z(n11184) );
  XNOR U13480 ( .A(n11087), .B(n11187), .Z(n11093) );
  XNOR U13481 ( .A(n11086), .B(n11088), .Z(n11187) );
  NAND U13482 ( .A(n11188), .B(n11189), .Z(n11088) );
  OR U13483 ( .A(n11190), .B(n11191), .Z(n11189) );
  OR U13484 ( .A(n11192), .B(n11193), .Z(n11188) );
  NAND U13485 ( .A(n11194), .B(n11195), .Z(n11086) );
  OR U13486 ( .A(n11196), .B(n11197), .Z(n11195) );
  OR U13487 ( .A(n11198), .B(n11199), .Z(n11194) );
  ANDN U13488 ( .B(n11200), .A(n11201), .Z(n11087) );
  IV U13489 ( .A(n11202), .Z(n11200) );
  XNOR U13490 ( .A(n11167), .B(n11166), .Z(N12957) );
  XOR U13491 ( .A(n11186), .B(n11185), .Z(n11166) );
  XNOR U13492 ( .A(n11201), .B(n11202), .Z(n11185) );
  XNOR U13493 ( .A(n11196), .B(n11197), .Z(n11202) );
  XNOR U13494 ( .A(n11198), .B(n11199), .Z(n11197) );
  XNOR U13495 ( .A(y[397]), .B(x[397]), .Z(n11199) );
  XNOR U13496 ( .A(y[398]), .B(x[398]), .Z(n11198) );
  XNOR U13497 ( .A(y[396]), .B(x[396]), .Z(n11196) );
  XNOR U13498 ( .A(n11190), .B(n11191), .Z(n11201) );
  XNOR U13499 ( .A(y[393]), .B(x[393]), .Z(n11191) );
  XNOR U13500 ( .A(n11192), .B(n11193), .Z(n11190) );
  XNOR U13501 ( .A(y[394]), .B(x[394]), .Z(n11193) );
  XNOR U13502 ( .A(y[395]), .B(x[395]), .Z(n11192) );
  XNOR U13503 ( .A(n11183), .B(n11182), .Z(n11186) );
  XNOR U13504 ( .A(n11178), .B(n11179), .Z(n11182) );
  XNOR U13505 ( .A(y[390]), .B(x[390]), .Z(n11179) );
  XNOR U13506 ( .A(n11180), .B(n11181), .Z(n11178) );
  XNOR U13507 ( .A(y[391]), .B(x[391]), .Z(n11181) );
  XNOR U13508 ( .A(y[392]), .B(x[392]), .Z(n11180) );
  XNOR U13509 ( .A(n11172), .B(n11173), .Z(n11183) );
  XNOR U13510 ( .A(y[387]), .B(x[387]), .Z(n11173) );
  XNOR U13511 ( .A(n11174), .B(n11175), .Z(n11172) );
  XNOR U13512 ( .A(y[388]), .B(x[388]), .Z(n11175) );
  XNOR U13513 ( .A(y[389]), .B(x[389]), .Z(n11174) );
  XOR U13514 ( .A(n11148), .B(n11149), .Z(n11167) );
  XNOR U13515 ( .A(n11164), .B(n11165), .Z(n11149) );
  XNOR U13516 ( .A(n11159), .B(n11160), .Z(n11165) );
  XNOR U13517 ( .A(n11161), .B(n11162), .Z(n11160) );
  XNOR U13518 ( .A(y[385]), .B(x[385]), .Z(n11162) );
  XNOR U13519 ( .A(y[386]), .B(x[386]), .Z(n11161) );
  XNOR U13520 ( .A(y[384]), .B(x[384]), .Z(n11159) );
  XNOR U13521 ( .A(n11153), .B(n11154), .Z(n11164) );
  XNOR U13522 ( .A(y[381]), .B(x[381]), .Z(n11154) );
  XNOR U13523 ( .A(n11155), .B(n11156), .Z(n11153) );
  XNOR U13524 ( .A(y[382]), .B(x[382]), .Z(n11156) );
  XNOR U13525 ( .A(y[383]), .B(x[383]), .Z(n11155) );
  XOR U13526 ( .A(n11147), .B(n11146), .Z(n11148) );
  XNOR U13527 ( .A(n11142), .B(n11143), .Z(n11146) );
  XNOR U13528 ( .A(y[378]), .B(x[378]), .Z(n11143) );
  XNOR U13529 ( .A(n11144), .B(n11145), .Z(n11142) );
  XNOR U13530 ( .A(y[379]), .B(x[379]), .Z(n11145) );
  XNOR U13531 ( .A(y[380]), .B(x[380]), .Z(n11144) );
  XNOR U13532 ( .A(n11136), .B(n11137), .Z(n11147) );
  XNOR U13533 ( .A(y[375]), .B(x[375]), .Z(n11137) );
  XNOR U13534 ( .A(n11138), .B(n11139), .Z(n11136) );
  XNOR U13535 ( .A(y[376]), .B(x[376]), .Z(n11139) );
  XNOR U13536 ( .A(y[377]), .B(x[377]), .Z(n11138) );
  NAND U13537 ( .A(n11203), .B(n11204), .Z(N12950) );
  NANDN U13538 ( .A(n11205), .B(n11206), .Z(n11204) );
  OR U13539 ( .A(n11207), .B(n11208), .Z(n11206) );
  NAND U13540 ( .A(n11207), .B(n11208), .Z(n11203) );
  XOR U13541 ( .A(n11207), .B(n11209), .Z(N12949) );
  XNOR U13542 ( .A(n11205), .B(n11208), .Z(n11209) );
  AND U13543 ( .A(n11210), .B(n11211), .Z(n11208) );
  NANDN U13544 ( .A(n11212), .B(n11213), .Z(n11211) );
  NANDN U13545 ( .A(n11214), .B(n11215), .Z(n11213) );
  NANDN U13546 ( .A(n11215), .B(n11214), .Z(n11210) );
  NAND U13547 ( .A(n11216), .B(n11217), .Z(n11205) );
  NANDN U13548 ( .A(n11218), .B(n11219), .Z(n11217) );
  OR U13549 ( .A(n11220), .B(n11221), .Z(n11219) );
  NAND U13550 ( .A(n11221), .B(n11220), .Z(n11216) );
  AND U13551 ( .A(n11222), .B(n11223), .Z(n11207) );
  NANDN U13552 ( .A(n11224), .B(n11225), .Z(n11223) );
  NANDN U13553 ( .A(n11226), .B(n11227), .Z(n11225) );
  NANDN U13554 ( .A(n11227), .B(n11226), .Z(n11222) );
  XOR U13555 ( .A(n11221), .B(n11228), .Z(N12948) );
  XOR U13556 ( .A(n11218), .B(n11220), .Z(n11228) );
  XNOR U13557 ( .A(n11214), .B(n11229), .Z(n11220) );
  XNOR U13558 ( .A(n11212), .B(n11215), .Z(n11229) );
  NAND U13559 ( .A(n11230), .B(n11231), .Z(n11215) );
  NAND U13560 ( .A(n11232), .B(n11233), .Z(n11231) );
  OR U13561 ( .A(n11234), .B(n11235), .Z(n11232) );
  NANDN U13562 ( .A(n11236), .B(n11234), .Z(n11230) );
  IV U13563 ( .A(n11235), .Z(n11236) );
  NAND U13564 ( .A(n11237), .B(n11238), .Z(n11212) );
  NAND U13565 ( .A(n11239), .B(n11240), .Z(n11238) );
  NANDN U13566 ( .A(n11241), .B(n11242), .Z(n11239) );
  NANDN U13567 ( .A(n11242), .B(n11241), .Z(n11237) );
  AND U13568 ( .A(n11243), .B(n11244), .Z(n11214) );
  NAND U13569 ( .A(n11245), .B(n11246), .Z(n11244) );
  OR U13570 ( .A(n11247), .B(n11248), .Z(n11245) );
  NANDN U13571 ( .A(n11249), .B(n11247), .Z(n11243) );
  NAND U13572 ( .A(n11250), .B(n11251), .Z(n11218) );
  NANDN U13573 ( .A(n11252), .B(n11253), .Z(n11251) );
  OR U13574 ( .A(n11254), .B(n11255), .Z(n11253) );
  NANDN U13575 ( .A(n11256), .B(n11254), .Z(n11250) );
  IV U13576 ( .A(n11255), .Z(n11256) );
  XNOR U13577 ( .A(n11226), .B(n11257), .Z(n11221) );
  XNOR U13578 ( .A(n11224), .B(n11227), .Z(n11257) );
  NAND U13579 ( .A(n11258), .B(n11259), .Z(n11227) );
  NAND U13580 ( .A(n11260), .B(n11261), .Z(n11259) );
  OR U13581 ( .A(n11262), .B(n11263), .Z(n11260) );
  NANDN U13582 ( .A(n11264), .B(n11262), .Z(n11258) );
  IV U13583 ( .A(n11263), .Z(n11264) );
  NAND U13584 ( .A(n11265), .B(n11266), .Z(n11224) );
  NAND U13585 ( .A(n11267), .B(n11268), .Z(n11266) );
  NANDN U13586 ( .A(n11269), .B(n11270), .Z(n11267) );
  NANDN U13587 ( .A(n11270), .B(n11269), .Z(n11265) );
  AND U13588 ( .A(n11271), .B(n11272), .Z(n11226) );
  NAND U13589 ( .A(n11273), .B(n11274), .Z(n11272) );
  OR U13590 ( .A(n11275), .B(n11276), .Z(n11273) );
  NANDN U13591 ( .A(n11277), .B(n11275), .Z(n11271) );
  XNOR U13592 ( .A(n11252), .B(n11278), .Z(N12947) );
  XOR U13593 ( .A(n11254), .B(n11255), .Z(n11278) );
  XNOR U13594 ( .A(n11268), .B(n11279), .Z(n11255) );
  XOR U13595 ( .A(n11269), .B(n11270), .Z(n11279) );
  XOR U13596 ( .A(n11275), .B(n11280), .Z(n11270) );
  XOR U13597 ( .A(n11274), .B(n11277), .Z(n11280) );
  IV U13598 ( .A(n11276), .Z(n11277) );
  NAND U13599 ( .A(n11281), .B(n11282), .Z(n11276) );
  OR U13600 ( .A(n11283), .B(n11284), .Z(n11282) );
  OR U13601 ( .A(n11285), .B(n11286), .Z(n11281) );
  NAND U13602 ( .A(n11287), .B(n11288), .Z(n11274) );
  OR U13603 ( .A(n11289), .B(n11290), .Z(n11288) );
  OR U13604 ( .A(n11291), .B(n11292), .Z(n11287) );
  NOR U13605 ( .A(n11293), .B(n11294), .Z(n11275) );
  ANDN U13606 ( .B(n11295), .A(n11296), .Z(n11269) );
  XNOR U13607 ( .A(n11262), .B(n11297), .Z(n11268) );
  XNOR U13608 ( .A(n11261), .B(n11263), .Z(n11297) );
  NAND U13609 ( .A(n11298), .B(n11299), .Z(n11263) );
  OR U13610 ( .A(n11300), .B(n11301), .Z(n11299) );
  OR U13611 ( .A(n11302), .B(n11303), .Z(n11298) );
  NAND U13612 ( .A(n11304), .B(n11305), .Z(n11261) );
  OR U13613 ( .A(n11306), .B(n11307), .Z(n11305) );
  OR U13614 ( .A(n11308), .B(n11309), .Z(n11304) );
  ANDN U13615 ( .B(n11310), .A(n11311), .Z(n11262) );
  IV U13616 ( .A(n11312), .Z(n11310) );
  ANDN U13617 ( .B(n11313), .A(n11314), .Z(n11254) );
  XOR U13618 ( .A(n11240), .B(n11315), .Z(n11252) );
  XOR U13619 ( .A(n11241), .B(n11242), .Z(n11315) );
  XOR U13620 ( .A(n11247), .B(n11316), .Z(n11242) );
  XOR U13621 ( .A(n11246), .B(n11249), .Z(n11316) );
  IV U13622 ( .A(n11248), .Z(n11249) );
  NAND U13623 ( .A(n11317), .B(n11318), .Z(n11248) );
  OR U13624 ( .A(n11319), .B(n11320), .Z(n11318) );
  OR U13625 ( .A(n11321), .B(n11322), .Z(n11317) );
  NAND U13626 ( .A(n11323), .B(n11324), .Z(n11246) );
  OR U13627 ( .A(n11325), .B(n11326), .Z(n11324) );
  OR U13628 ( .A(n11327), .B(n11328), .Z(n11323) );
  NOR U13629 ( .A(n11329), .B(n11330), .Z(n11247) );
  ANDN U13630 ( .B(n11331), .A(n11332), .Z(n11241) );
  IV U13631 ( .A(n11333), .Z(n11331) );
  XNOR U13632 ( .A(n11234), .B(n11334), .Z(n11240) );
  XNOR U13633 ( .A(n11233), .B(n11235), .Z(n11334) );
  NAND U13634 ( .A(n11335), .B(n11336), .Z(n11235) );
  OR U13635 ( .A(n11337), .B(n11338), .Z(n11336) );
  OR U13636 ( .A(n11339), .B(n11340), .Z(n11335) );
  NAND U13637 ( .A(n11341), .B(n11342), .Z(n11233) );
  OR U13638 ( .A(n11343), .B(n11344), .Z(n11342) );
  OR U13639 ( .A(n11345), .B(n11346), .Z(n11341) );
  ANDN U13640 ( .B(n11347), .A(n11348), .Z(n11234) );
  IV U13641 ( .A(n11349), .Z(n11347) );
  XNOR U13642 ( .A(n11314), .B(n11313), .Z(N12946) );
  XOR U13643 ( .A(n11333), .B(n11332), .Z(n11313) );
  XNOR U13644 ( .A(n11348), .B(n11349), .Z(n11332) );
  XNOR U13645 ( .A(n11343), .B(n11344), .Z(n11349) );
  XNOR U13646 ( .A(n11345), .B(n11346), .Z(n11344) );
  XNOR U13647 ( .A(y[373]), .B(x[373]), .Z(n11346) );
  XNOR U13648 ( .A(y[374]), .B(x[374]), .Z(n11345) );
  XNOR U13649 ( .A(y[372]), .B(x[372]), .Z(n11343) );
  XNOR U13650 ( .A(n11337), .B(n11338), .Z(n11348) );
  XNOR U13651 ( .A(y[369]), .B(x[369]), .Z(n11338) );
  XNOR U13652 ( .A(n11339), .B(n11340), .Z(n11337) );
  XNOR U13653 ( .A(y[370]), .B(x[370]), .Z(n11340) );
  XNOR U13654 ( .A(y[371]), .B(x[371]), .Z(n11339) );
  XNOR U13655 ( .A(n11330), .B(n11329), .Z(n11333) );
  XNOR U13656 ( .A(n11325), .B(n11326), .Z(n11329) );
  XNOR U13657 ( .A(y[366]), .B(x[366]), .Z(n11326) );
  XNOR U13658 ( .A(n11327), .B(n11328), .Z(n11325) );
  XNOR U13659 ( .A(y[367]), .B(x[367]), .Z(n11328) );
  XNOR U13660 ( .A(y[368]), .B(x[368]), .Z(n11327) );
  XNOR U13661 ( .A(n11319), .B(n11320), .Z(n11330) );
  XNOR U13662 ( .A(y[363]), .B(x[363]), .Z(n11320) );
  XNOR U13663 ( .A(n11321), .B(n11322), .Z(n11319) );
  XNOR U13664 ( .A(y[364]), .B(x[364]), .Z(n11322) );
  XNOR U13665 ( .A(y[365]), .B(x[365]), .Z(n11321) );
  XOR U13666 ( .A(n11295), .B(n11296), .Z(n11314) );
  XNOR U13667 ( .A(n11311), .B(n11312), .Z(n11296) );
  XNOR U13668 ( .A(n11306), .B(n11307), .Z(n11312) );
  XNOR U13669 ( .A(n11308), .B(n11309), .Z(n11307) );
  XNOR U13670 ( .A(y[361]), .B(x[361]), .Z(n11309) );
  XNOR U13671 ( .A(y[362]), .B(x[362]), .Z(n11308) );
  XNOR U13672 ( .A(y[360]), .B(x[360]), .Z(n11306) );
  XNOR U13673 ( .A(n11300), .B(n11301), .Z(n11311) );
  XNOR U13674 ( .A(y[357]), .B(x[357]), .Z(n11301) );
  XNOR U13675 ( .A(n11302), .B(n11303), .Z(n11300) );
  XNOR U13676 ( .A(y[358]), .B(x[358]), .Z(n11303) );
  XNOR U13677 ( .A(y[359]), .B(x[359]), .Z(n11302) );
  XOR U13678 ( .A(n11294), .B(n11293), .Z(n11295) );
  XNOR U13679 ( .A(n11289), .B(n11290), .Z(n11293) );
  XNOR U13680 ( .A(y[354]), .B(x[354]), .Z(n11290) );
  XNOR U13681 ( .A(n11291), .B(n11292), .Z(n11289) );
  XNOR U13682 ( .A(y[355]), .B(x[355]), .Z(n11292) );
  XNOR U13683 ( .A(y[356]), .B(x[356]), .Z(n11291) );
  XNOR U13684 ( .A(n11283), .B(n11284), .Z(n11294) );
  XNOR U13685 ( .A(y[351]), .B(x[351]), .Z(n11284) );
  XNOR U13686 ( .A(n11285), .B(n11286), .Z(n11283) );
  XNOR U13687 ( .A(y[352]), .B(x[352]), .Z(n11286) );
  XNOR U13688 ( .A(y[353]), .B(x[353]), .Z(n11285) );
  NAND U13689 ( .A(n11350), .B(n11351), .Z(N12939) );
  NANDN U13690 ( .A(n11352), .B(n11353), .Z(n11351) );
  OR U13691 ( .A(n11354), .B(n11355), .Z(n11353) );
  NAND U13692 ( .A(n11354), .B(n11355), .Z(n11350) );
  XOR U13693 ( .A(n11354), .B(n11356), .Z(N12938) );
  XNOR U13694 ( .A(n11352), .B(n11355), .Z(n11356) );
  AND U13695 ( .A(n11357), .B(n11358), .Z(n11355) );
  NANDN U13696 ( .A(n11359), .B(n11360), .Z(n11358) );
  NANDN U13697 ( .A(n11361), .B(n11362), .Z(n11360) );
  NANDN U13698 ( .A(n11362), .B(n11361), .Z(n11357) );
  NAND U13699 ( .A(n11363), .B(n11364), .Z(n11352) );
  NANDN U13700 ( .A(n11365), .B(n11366), .Z(n11364) );
  OR U13701 ( .A(n11367), .B(n11368), .Z(n11366) );
  NAND U13702 ( .A(n11368), .B(n11367), .Z(n11363) );
  AND U13703 ( .A(n11369), .B(n11370), .Z(n11354) );
  NANDN U13704 ( .A(n11371), .B(n11372), .Z(n11370) );
  NANDN U13705 ( .A(n11373), .B(n11374), .Z(n11372) );
  NANDN U13706 ( .A(n11374), .B(n11373), .Z(n11369) );
  XOR U13707 ( .A(n11368), .B(n11375), .Z(N12937) );
  XOR U13708 ( .A(n11365), .B(n11367), .Z(n11375) );
  XNOR U13709 ( .A(n11361), .B(n11376), .Z(n11367) );
  XNOR U13710 ( .A(n11359), .B(n11362), .Z(n11376) );
  NAND U13711 ( .A(n11377), .B(n11378), .Z(n11362) );
  NAND U13712 ( .A(n11379), .B(n11380), .Z(n11378) );
  OR U13713 ( .A(n11381), .B(n11382), .Z(n11379) );
  NANDN U13714 ( .A(n11383), .B(n11381), .Z(n11377) );
  IV U13715 ( .A(n11382), .Z(n11383) );
  NAND U13716 ( .A(n11384), .B(n11385), .Z(n11359) );
  NAND U13717 ( .A(n11386), .B(n11387), .Z(n11385) );
  NANDN U13718 ( .A(n11388), .B(n11389), .Z(n11386) );
  NANDN U13719 ( .A(n11389), .B(n11388), .Z(n11384) );
  AND U13720 ( .A(n11390), .B(n11391), .Z(n11361) );
  NAND U13721 ( .A(n11392), .B(n11393), .Z(n11391) );
  OR U13722 ( .A(n11394), .B(n11395), .Z(n11392) );
  NANDN U13723 ( .A(n11396), .B(n11394), .Z(n11390) );
  NAND U13724 ( .A(n11397), .B(n11398), .Z(n11365) );
  NANDN U13725 ( .A(n11399), .B(n11400), .Z(n11398) );
  OR U13726 ( .A(n11401), .B(n11402), .Z(n11400) );
  NANDN U13727 ( .A(n11403), .B(n11401), .Z(n11397) );
  IV U13728 ( .A(n11402), .Z(n11403) );
  XNOR U13729 ( .A(n11373), .B(n11404), .Z(n11368) );
  XNOR U13730 ( .A(n11371), .B(n11374), .Z(n11404) );
  NAND U13731 ( .A(n11405), .B(n11406), .Z(n11374) );
  NAND U13732 ( .A(n11407), .B(n11408), .Z(n11406) );
  OR U13733 ( .A(n11409), .B(n11410), .Z(n11407) );
  NANDN U13734 ( .A(n11411), .B(n11409), .Z(n11405) );
  IV U13735 ( .A(n11410), .Z(n11411) );
  NAND U13736 ( .A(n11412), .B(n11413), .Z(n11371) );
  NAND U13737 ( .A(n11414), .B(n11415), .Z(n11413) );
  NANDN U13738 ( .A(n11416), .B(n11417), .Z(n11414) );
  NANDN U13739 ( .A(n11417), .B(n11416), .Z(n11412) );
  AND U13740 ( .A(n11418), .B(n11419), .Z(n11373) );
  NAND U13741 ( .A(n11420), .B(n11421), .Z(n11419) );
  OR U13742 ( .A(n11422), .B(n11423), .Z(n11420) );
  NANDN U13743 ( .A(n11424), .B(n11422), .Z(n11418) );
  XNOR U13744 ( .A(n11399), .B(n11425), .Z(N12936) );
  XOR U13745 ( .A(n11401), .B(n11402), .Z(n11425) );
  XNOR U13746 ( .A(n11415), .B(n11426), .Z(n11402) );
  XOR U13747 ( .A(n11416), .B(n11417), .Z(n11426) );
  XOR U13748 ( .A(n11422), .B(n11427), .Z(n11417) );
  XOR U13749 ( .A(n11421), .B(n11424), .Z(n11427) );
  IV U13750 ( .A(n11423), .Z(n11424) );
  NAND U13751 ( .A(n11428), .B(n11429), .Z(n11423) );
  OR U13752 ( .A(n11430), .B(n11431), .Z(n11429) );
  OR U13753 ( .A(n11432), .B(n11433), .Z(n11428) );
  NAND U13754 ( .A(n11434), .B(n11435), .Z(n11421) );
  OR U13755 ( .A(n11436), .B(n11437), .Z(n11435) );
  OR U13756 ( .A(n11438), .B(n11439), .Z(n11434) );
  NOR U13757 ( .A(n11440), .B(n11441), .Z(n11422) );
  ANDN U13758 ( .B(n11442), .A(n11443), .Z(n11416) );
  XNOR U13759 ( .A(n11409), .B(n11444), .Z(n11415) );
  XNOR U13760 ( .A(n11408), .B(n11410), .Z(n11444) );
  NAND U13761 ( .A(n11445), .B(n11446), .Z(n11410) );
  OR U13762 ( .A(n11447), .B(n11448), .Z(n11446) );
  OR U13763 ( .A(n11449), .B(n11450), .Z(n11445) );
  NAND U13764 ( .A(n11451), .B(n11452), .Z(n11408) );
  OR U13765 ( .A(n11453), .B(n11454), .Z(n11452) );
  OR U13766 ( .A(n11455), .B(n11456), .Z(n11451) );
  ANDN U13767 ( .B(n11457), .A(n11458), .Z(n11409) );
  IV U13768 ( .A(n11459), .Z(n11457) );
  ANDN U13769 ( .B(n11460), .A(n11461), .Z(n11401) );
  XOR U13770 ( .A(n11387), .B(n11462), .Z(n11399) );
  XOR U13771 ( .A(n11388), .B(n11389), .Z(n11462) );
  XOR U13772 ( .A(n11394), .B(n11463), .Z(n11389) );
  XOR U13773 ( .A(n11393), .B(n11396), .Z(n11463) );
  IV U13774 ( .A(n11395), .Z(n11396) );
  NAND U13775 ( .A(n11464), .B(n11465), .Z(n11395) );
  OR U13776 ( .A(n11466), .B(n11467), .Z(n11465) );
  OR U13777 ( .A(n11468), .B(n11469), .Z(n11464) );
  NAND U13778 ( .A(n11470), .B(n11471), .Z(n11393) );
  OR U13779 ( .A(n11472), .B(n11473), .Z(n11471) );
  OR U13780 ( .A(n11474), .B(n11475), .Z(n11470) );
  NOR U13781 ( .A(n11476), .B(n11477), .Z(n11394) );
  ANDN U13782 ( .B(n11478), .A(n11479), .Z(n11388) );
  IV U13783 ( .A(n11480), .Z(n11478) );
  XNOR U13784 ( .A(n11381), .B(n11481), .Z(n11387) );
  XNOR U13785 ( .A(n11380), .B(n11382), .Z(n11481) );
  NAND U13786 ( .A(n11482), .B(n11483), .Z(n11382) );
  OR U13787 ( .A(n11484), .B(n11485), .Z(n11483) );
  OR U13788 ( .A(n11486), .B(n11487), .Z(n11482) );
  NAND U13789 ( .A(n11488), .B(n11489), .Z(n11380) );
  OR U13790 ( .A(n11490), .B(n11491), .Z(n11489) );
  OR U13791 ( .A(n11492), .B(n11493), .Z(n11488) );
  ANDN U13792 ( .B(n11494), .A(n11495), .Z(n11381) );
  IV U13793 ( .A(n11496), .Z(n11494) );
  XNOR U13794 ( .A(n11461), .B(n11460), .Z(N12935) );
  XOR U13795 ( .A(n11480), .B(n11479), .Z(n11460) );
  XNOR U13796 ( .A(n11495), .B(n11496), .Z(n11479) );
  XNOR U13797 ( .A(n11490), .B(n11491), .Z(n11496) );
  XNOR U13798 ( .A(n11492), .B(n11493), .Z(n11491) );
  XNOR U13799 ( .A(y[349]), .B(x[349]), .Z(n11493) );
  XNOR U13800 ( .A(y[350]), .B(x[350]), .Z(n11492) );
  XNOR U13801 ( .A(y[348]), .B(x[348]), .Z(n11490) );
  XNOR U13802 ( .A(n11484), .B(n11485), .Z(n11495) );
  XNOR U13803 ( .A(y[345]), .B(x[345]), .Z(n11485) );
  XNOR U13804 ( .A(n11486), .B(n11487), .Z(n11484) );
  XNOR U13805 ( .A(y[346]), .B(x[346]), .Z(n11487) );
  XNOR U13806 ( .A(y[347]), .B(x[347]), .Z(n11486) );
  XNOR U13807 ( .A(n11477), .B(n11476), .Z(n11480) );
  XNOR U13808 ( .A(n11472), .B(n11473), .Z(n11476) );
  XNOR U13809 ( .A(y[342]), .B(x[342]), .Z(n11473) );
  XNOR U13810 ( .A(n11474), .B(n11475), .Z(n11472) );
  XNOR U13811 ( .A(y[343]), .B(x[343]), .Z(n11475) );
  XNOR U13812 ( .A(y[344]), .B(x[344]), .Z(n11474) );
  XNOR U13813 ( .A(n11466), .B(n11467), .Z(n11477) );
  XNOR U13814 ( .A(y[339]), .B(x[339]), .Z(n11467) );
  XNOR U13815 ( .A(n11468), .B(n11469), .Z(n11466) );
  XNOR U13816 ( .A(y[340]), .B(x[340]), .Z(n11469) );
  XNOR U13817 ( .A(y[341]), .B(x[341]), .Z(n11468) );
  XOR U13818 ( .A(n11442), .B(n11443), .Z(n11461) );
  XNOR U13819 ( .A(n11458), .B(n11459), .Z(n11443) );
  XNOR U13820 ( .A(n11453), .B(n11454), .Z(n11459) );
  XNOR U13821 ( .A(n11455), .B(n11456), .Z(n11454) );
  XNOR U13822 ( .A(y[337]), .B(x[337]), .Z(n11456) );
  XNOR U13823 ( .A(y[338]), .B(x[338]), .Z(n11455) );
  XNOR U13824 ( .A(y[336]), .B(x[336]), .Z(n11453) );
  XNOR U13825 ( .A(n11447), .B(n11448), .Z(n11458) );
  XNOR U13826 ( .A(y[333]), .B(x[333]), .Z(n11448) );
  XNOR U13827 ( .A(n11449), .B(n11450), .Z(n11447) );
  XNOR U13828 ( .A(y[334]), .B(x[334]), .Z(n11450) );
  XNOR U13829 ( .A(y[335]), .B(x[335]), .Z(n11449) );
  XOR U13830 ( .A(n11441), .B(n11440), .Z(n11442) );
  XNOR U13831 ( .A(n11436), .B(n11437), .Z(n11440) );
  XNOR U13832 ( .A(y[330]), .B(x[330]), .Z(n11437) );
  XNOR U13833 ( .A(n11438), .B(n11439), .Z(n11436) );
  XNOR U13834 ( .A(y[331]), .B(x[331]), .Z(n11439) );
  XNOR U13835 ( .A(y[332]), .B(x[332]), .Z(n11438) );
  XNOR U13836 ( .A(n11430), .B(n11431), .Z(n11441) );
  XNOR U13837 ( .A(y[327]), .B(x[327]), .Z(n11431) );
  XNOR U13838 ( .A(n11432), .B(n11433), .Z(n11430) );
  XNOR U13839 ( .A(y[328]), .B(x[328]), .Z(n11433) );
  XNOR U13840 ( .A(y[329]), .B(x[329]), .Z(n11432) );
  NAND U13841 ( .A(n11497), .B(n11498), .Z(N12928) );
  NANDN U13842 ( .A(n11499), .B(n11500), .Z(n11498) );
  OR U13843 ( .A(n11501), .B(n11502), .Z(n11500) );
  NAND U13844 ( .A(n11501), .B(n11502), .Z(n11497) );
  XOR U13845 ( .A(n11501), .B(n11503), .Z(N12927) );
  XNOR U13846 ( .A(n11499), .B(n11502), .Z(n11503) );
  AND U13847 ( .A(n11504), .B(n11505), .Z(n11502) );
  NANDN U13848 ( .A(n11506), .B(n11507), .Z(n11505) );
  NANDN U13849 ( .A(n11508), .B(n11509), .Z(n11507) );
  NANDN U13850 ( .A(n11509), .B(n11508), .Z(n11504) );
  NAND U13851 ( .A(n11510), .B(n11511), .Z(n11499) );
  NANDN U13852 ( .A(n11512), .B(n11513), .Z(n11511) );
  OR U13853 ( .A(n11514), .B(n11515), .Z(n11513) );
  NAND U13854 ( .A(n11515), .B(n11514), .Z(n11510) );
  AND U13855 ( .A(n11516), .B(n11517), .Z(n11501) );
  NANDN U13856 ( .A(n11518), .B(n11519), .Z(n11517) );
  NANDN U13857 ( .A(n11520), .B(n11521), .Z(n11519) );
  NANDN U13858 ( .A(n11521), .B(n11520), .Z(n11516) );
  XOR U13859 ( .A(n11515), .B(n11522), .Z(N12926) );
  XOR U13860 ( .A(n11512), .B(n11514), .Z(n11522) );
  XNOR U13861 ( .A(n11508), .B(n11523), .Z(n11514) );
  XNOR U13862 ( .A(n11506), .B(n11509), .Z(n11523) );
  NAND U13863 ( .A(n11524), .B(n11525), .Z(n11509) );
  NAND U13864 ( .A(n11526), .B(n11527), .Z(n11525) );
  OR U13865 ( .A(n11528), .B(n11529), .Z(n11526) );
  NANDN U13866 ( .A(n11530), .B(n11528), .Z(n11524) );
  IV U13867 ( .A(n11529), .Z(n11530) );
  NAND U13868 ( .A(n11531), .B(n11532), .Z(n11506) );
  NAND U13869 ( .A(n11533), .B(n11534), .Z(n11532) );
  NANDN U13870 ( .A(n11535), .B(n11536), .Z(n11533) );
  NANDN U13871 ( .A(n11536), .B(n11535), .Z(n11531) );
  AND U13872 ( .A(n11537), .B(n11538), .Z(n11508) );
  NAND U13873 ( .A(n11539), .B(n11540), .Z(n11538) );
  OR U13874 ( .A(n11541), .B(n11542), .Z(n11539) );
  NANDN U13875 ( .A(n11543), .B(n11541), .Z(n11537) );
  NAND U13876 ( .A(n11544), .B(n11545), .Z(n11512) );
  NANDN U13877 ( .A(n11546), .B(n11547), .Z(n11545) );
  OR U13878 ( .A(n11548), .B(n11549), .Z(n11547) );
  NANDN U13879 ( .A(n11550), .B(n11548), .Z(n11544) );
  IV U13880 ( .A(n11549), .Z(n11550) );
  XNOR U13881 ( .A(n11520), .B(n11551), .Z(n11515) );
  XNOR U13882 ( .A(n11518), .B(n11521), .Z(n11551) );
  NAND U13883 ( .A(n11552), .B(n11553), .Z(n11521) );
  NAND U13884 ( .A(n11554), .B(n11555), .Z(n11553) );
  OR U13885 ( .A(n11556), .B(n11557), .Z(n11554) );
  NANDN U13886 ( .A(n11558), .B(n11556), .Z(n11552) );
  IV U13887 ( .A(n11557), .Z(n11558) );
  NAND U13888 ( .A(n11559), .B(n11560), .Z(n11518) );
  NAND U13889 ( .A(n11561), .B(n11562), .Z(n11560) );
  NANDN U13890 ( .A(n11563), .B(n11564), .Z(n11561) );
  NANDN U13891 ( .A(n11564), .B(n11563), .Z(n11559) );
  AND U13892 ( .A(n11565), .B(n11566), .Z(n11520) );
  NAND U13893 ( .A(n11567), .B(n11568), .Z(n11566) );
  OR U13894 ( .A(n11569), .B(n11570), .Z(n11567) );
  NANDN U13895 ( .A(n11571), .B(n11569), .Z(n11565) );
  XNOR U13896 ( .A(n11546), .B(n11572), .Z(N12925) );
  XOR U13897 ( .A(n11548), .B(n11549), .Z(n11572) );
  XNOR U13898 ( .A(n11562), .B(n11573), .Z(n11549) );
  XOR U13899 ( .A(n11563), .B(n11564), .Z(n11573) );
  XOR U13900 ( .A(n11569), .B(n11574), .Z(n11564) );
  XOR U13901 ( .A(n11568), .B(n11571), .Z(n11574) );
  IV U13902 ( .A(n11570), .Z(n11571) );
  NAND U13903 ( .A(n11575), .B(n11576), .Z(n11570) );
  OR U13904 ( .A(n11577), .B(n11578), .Z(n11576) );
  OR U13905 ( .A(n11579), .B(n11580), .Z(n11575) );
  NAND U13906 ( .A(n11581), .B(n11582), .Z(n11568) );
  OR U13907 ( .A(n11583), .B(n11584), .Z(n11582) );
  OR U13908 ( .A(n11585), .B(n11586), .Z(n11581) );
  NOR U13909 ( .A(n11587), .B(n11588), .Z(n11569) );
  ANDN U13910 ( .B(n11589), .A(n11590), .Z(n11563) );
  XNOR U13911 ( .A(n11556), .B(n11591), .Z(n11562) );
  XNOR U13912 ( .A(n11555), .B(n11557), .Z(n11591) );
  NAND U13913 ( .A(n11592), .B(n11593), .Z(n11557) );
  OR U13914 ( .A(n11594), .B(n11595), .Z(n11593) );
  OR U13915 ( .A(n11596), .B(n11597), .Z(n11592) );
  NAND U13916 ( .A(n11598), .B(n11599), .Z(n11555) );
  OR U13917 ( .A(n11600), .B(n11601), .Z(n11599) );
  OR U13918 ( .A(n11602), .B(n11603), .Z(n11598) );
  ANDN U13919 ( .B(n11604), .A(n11605), .Z(n11556) );
  IV U13920 ( .A(n11606), .Z(n11604) );
  ANDN U13921 ( .B(n11607), .A(n11608), .Z(n11548) );
  XOR U13922 ( .A(n11534), .B(n11609), .Z(n11546) );
  XOR U13923 ( .A(n11535), .B(n11536), .Z(n11609) );
  XOR U13924 ( .A(n11541), .B(n11610), .Z(n11536) );
  XOR U13925 ( .A(n11540), .B(n11543), .Z(n11610) );
  IV U13926 ( .A(n11542), .Z(n11543) );
  NAND U13927 ( .A(n11611), .B(n11612), .Z(n11542) );
  OR U13928 ( .A(n11613), .B(n11614), .Z(n11612) );
  OR U13929 ( .A(n11615), .B(n11616), .Z(n11611) );
  NAND U13930 ( .A(n11617), .B(n11618), .Z(n11540) );
  OR U13931 ( .A(n11619), .B(n11620), .Z(n11618) );
  OR U13932 ( .A(n11621), .B(n11622), .Z(n11617) );
  NOR U13933 ( .A(n11623), .B(n11624), .Z(n11541) );
  ANDN U13934 ( .B(n11625), .A(n11626), .Z(n11535) );
  IV U13935 ( .A(n11627), .Z(n11625) );
  XNOR U13936 ( .A(n11528), .B(n11628), .Z(n11534) );
  XNOR U13937 ( .A(n11527), .B(n11529), .Z(n11628) );
  NAND U13938 ( .A(n11629), .B(n11630), .Z(n11529) );
  OR U13939 ( .A(n11631), .B(n11632), .Z(n11630) );
  OR U13940 ( .A(n11633), .B(n11634), .Z(n11629) );
  NAND U13941 ( .A(n11635), .B(n11636), .Z(n11527) );
  OR U13942 ( .A(n11637), .B(n11638), .Z(n11636) );
  OR U13943 ( .A(n11639), .B(n11640), .Z(n11635) );
  ANDN U13944 ( .B(n11641), .A(n11642), .Z(n11528) );
  IV U13945 ( .A(n11643), .Z(n11641) );
  XNOR U13946 ( .A(n11608), .B(n11607), .Z(N12924) );
  XOR U13947 ( .A(n11627), .B(n11626), .Z(n11607) );
  XNOR U13948 ( .A(n11642), .B(n11643), .Z(n11626) );
  XNOR U13949 ( .A(n11637), .B(n11638), .Z(n11643) );
  XNOR U13950 ( .A(n11639), .B(n11640), .Z(n11638) );
  XNOR U13951 ( .A(y[325]), .B(x[325]), .Z(n11640) );
  XNOR U13952 ( .A(y[326]), .B(x[326]), .Z(n11639) );
  XNOR U13953 ( .A(y[324]), .B(x[324]), .Z(n11637) );
  XNOR U13954 ( .A(n11631), .B(n11632), .Z(n11642) );
  XNOR U13955 ( .A(y[321]), .B(x[321]), .Z(n11632) );
  XNOR U13956 ( .A(n11633), .B(n11634), .Z(n11631) );
  XNOR U13957 ( .A(y[322]), .B(x[322]), .Z(n11634) );
  XNOR U13958 ( .A(y[323]), .B(x[323]), .Z(n11633) );
  XNOR U13959 ( .A(n11624), .B(n11623), .Z(n11627) );
  XNOR U13960 ( .A(n11619), .B(n11620), .Z(n11623) );
  XNOR U13961 ( .A(y[318]), .B(x[318]), .Z(n11620) );
  XNOR U13962 ( .A(n11621), .B(n11622), .Z(n11619) );
  XNOR U13963 ( .A(y[319]), .B(x[319]), .Z(n11622) );
  XNOR U13964 ( .A(y[320]), .B(x[320]), .Z(n11621) );
  XNOR U13965 ( .A(n11613), .B(n11614), .Z(n11624) );
  XNOR U13966 ( .A(y[315]), .B(x[315]), .Z(n11614) );
  XNOR U13967 ( .A(n11615), .B(n11616), .Z(n11613) );
  XNOR U13968 ( .A(y[316]), .B(x[316]), .Z(n11616) );
  XNOR U13969 ( .A(y[317]), .B(x[317]), .Z(n11615) );
  XOR U13970 ( .A(n11589), .B(n11590), .Z(n11608) );
  XNOR U13971 ( .A(n11605), .B(n11606), .Z(n11590) );
  XNOR U13972 ( .A(n11600), .B(n11601), .Z(n11606) );
  XNOR U13973 ( .A(n11602), .B(n11603), .Z(n11601) );
  XNOR U13974 ( .A(y[313]), .B(x[313]), .Z(n11603) );
  XNOR U13975 ( .A(y[314]), .B(x[314]), .Z(n11602) );
  XNOR U13976 ( .A(y[312]), .B(x[312]), .Z(n11600) );
  XNOR U13977 ( .A(n11594), .B(n11595), .Z(n11605) );
  XNOR U13978 ( .A(y[309]), .B(x[309]), .Z(n11595) );
  XNOR U13979 ( .A(n11596), .B(n11597), .Z(n11594) );
  XNOR U13980 ( .A(y[310]), .B(x[310]), .Z(n11597) );
  XNOR U13981 ( .A(y[311]), .B(x[311]), .Z(n11596) );
  XOR U13982 ( .A(n11588), .B(n11587), .Z(n11589) );
  XNOR U13983 ( .A(n11583), .B(n11584), .Z(n11587) );
  XNOR U13984 ( .A(y[306]), .B(x[306]), .Z(n11584) );
  XNOR U13985 ( .A(n11585), .B(n11586), .Z(n11583) );
  XNOR U13986 ( .A(y[307]), .B(x[307]), .Z(n11586) );
  XNOR U13987 ( .A(y[308]), .B(x[308]), .Z(n11585) );
  XNOR U13988 ( .A(n11577), .B(n11578), .Z(n11588) );
  XNOR U13989 ( .A(y[303]), .B(x[303]), .Z(n11578) );
  XNOR U13990 ( .A(n11579), .B(n11580), .Z(n11577) );
  XNOR U13991 ( .A(y[304]), .B(x[304]), .Z(n11580) );
  XNOR U13992 ( .A(y[305]), .B(x[305]), .Z(n11579) );
  NAND U13993 ( .A(n11644), .B(n11645), .Z(N12917) );
  NANDN U13994 ( .A(n11646), .B(n11647), .Z(n11645) );
  OR U13995 ( .A(n11648), .B(n11649), .Z(n11647) );
  NAND U13996 ( .A(n11648), .B(n11649), .Z(n11644) );
  XOR U13997 ( .A(n11648), .B(n11650), .Z(N12916) );
  XNOR U13998 ( .A(n11646), .B(n11649), .Z(n11650) );
  AND U13999 ( .A(n11651), .B(n11652), .Z(n11649) );
  NANDN U14000 ( .A(n11653), .B(n11654), .Z(n11652) );
  NANDN U14001 ( .A(n11655), .B(n11656), .Z(n11654) );
  NANDN U14002 ( .A(n11656), .B(n11655), .Z(n11651) );
  NAND U14003 ( .A(n11657), .B(n11658), .Z(n11646) );
  NANDN U14004 ( .A(n11659), .B(n11660), .Z(n11658) );
  OR U14005 ( .A(n11661), .B(n11662), .Z(n11660) );
  NAND U14006 ( .A(n11662), .B(n11661), .Z(n11657) );
  AND U14007 ( .A(n11663), .B(n11664), .Z(n11648) );
  NANDN U14008 ( .A(n11665), .B(n11666), .Z(n11664) );
  NANDN U14009 ( .A(n11667), .B(n11668), .Z(n11666) );
  NANDN U14010 ( .A(n11668), .B(n11667), .Z(n11663) );
  XOR U14011 ( .A(n11662), .B(n11669), .Z(N12915) );
  XOR U14012 ( .A(n11659), .B(n11661), .Z(n11669) );
  XNOR U14013 ( .A(n11655), .B(n11670), .Z(n11661) );
  XNOR U14014 ( .A(n11653), .B(n11656), .Z(n11670) );
  NAND U14015 ( .A(n11671), .B(n11672), .Z(n11656) );
  NAND U14016 ( .A(n11673), .B(n11674), .Z(n11672) );
  OR U14017 ( .A(n11675), .B(n11676), .Z(n11673) );
  NANDN U14018 ( .A(n11677), .B(n11675), .Z(n11671) );
  IV U14019 ( .A(n11676), .Z(n11677) );
  NAND U14020 ( .A(n11678), .B(n11679), .Z(n11653) );
  NAND U14021 ( .A(n11680), .B(n11681), .Z(n11679) );
  NANDN U14022 ( .A(n11682), .B(n11683), .Z(n11680) );
  NANDN U14023 ( .A(n11683), .B(n11682), .Z(n11678) );
  AND U14024 ( .A(n11684), .B(n11685), .Z(n11655) );
  NAND U14025 ( .A(n11686), .B(n11687), .Z(n11685) );
  OR U14026 ( .A(n11688), .B(n11689), .Z(n11686) );
  NANDN U14027 ( .A(n11690), .B(n11688), .Z(n11684) );
  NAND U14028 ( .A(n11691), .B(n11692), .Z(n11659) );
  NANDN U14029 ( .A(n11693), .B(n11694), .Z(n11692) );
  OR U14030 ( .A(n11695), .B(n11696), .Z(n11694) );
  NANDN U14031 ( .A(n11697), .B(n11695), .Z(n11691) );
  IV U14032 ( .A(n11696), .Z(n11697) );
  XNOR U14033 ( .A(n11667), .B(n11698), .Z(n11662) );
  XNOR U14034 ( .A(n11665), .B(n11668), .Z(n11698) );
  NAND U14035 ( .A(n11699), .B(n11700), .Z(n11668) );
  NAND U14036 ( .A(n11701), .B(n11702), .Z(n11700) );
  OR U14037 ( .A(n11703), .B(n11704), .Z(n11701) );
  NANDN U14038 ( .A(n11705), .B(n11703), .Z(n11699) );
  IV U14039 ( .A(n11704), .Z(n11705) );
  NAND U14040 ( .A(n11706), .B(n11707), .Z(n11665) );
  NAND U14041 ( .A(n11708), .B(n11709), .Z(n11707) );
  NANDN U14042 ( .A(n11710), .B(n11711), .Z(n11708) );
  NANDN U14043 ( .A(n11711), .B(n11710), .Z(n11706) );
  AND U14044 ( .A(n11712), .B(n11713), .Z(n11667) );
  NAND U14045 ( .A(n11714), .B(n11715), .Z(n11713) );
  OR U14046 ( .A(n11716), .B(n11717), .Z(n11714) );
  NANDN U14047 ( .A(n11718), .B(n11716), .Z(n11712) );
  XNOR U14048 ( .A(n11693), .B(n11719), .Z(N12914) );
  XOR U14049 ( .A(n11695), .B(n11696), .Z(n11719) );
  XNOR U14050 ( .A(n11709), .B(n11720), .Z(n11696) );
  XOR U14051 ( .A(n11710), .B(n11711), .Z(n11720) );
  XOR U14052 ( .A(n11716), .B(n11721), .Z(n11711) );
  XOR U14053 ( .A(n11715), .B(n11718), .Z(n11721) );
  IV U14054 ( .A(n11717), .Z(n11718) );
  NAND U14055 ( .A(n11722), .B(n11723), .Z(n11717) );
  OR U14056 ( .A(n11724), .B(n11725), .Z(n11723) );
  OR U14057 ( .A(n11726), .B(n11727), .Z(n11722) );
  NAND U14058 ( .A(n11728), .B(n11729), .Z(n11715) );
  OR U14059 ( .A(n11730), .B(n11731), .Z(n11729) );
  OR U14060 ( .A(n11732), .B(n11733), .Z(n11728) );
  NOR U14061 ( .A(n11734), .B(n11735), .Z(n11716) );
  ANDN U14062 ( .B(n11736), .A(n11737), .Z(n11710) );
  XNOR U14063 ( .A(n11703), .B(n11738), .Z(n11709) );
  XNOR U14064 ( .A(n11702), .B(n11704), .Z(n11738) );
  NAND U14065 ( .A(n11739), .B(n11740), .Z(n11704) );
  OR U14066 ( .A(n11741), .B(n11742), .Z(n11740) );
  OR U14067 ( .A(n11743), .B(n11744), .Z(n11739) );
  NAND U14068 ( .A(n11745), .B(n11746), .Z(n11702) );
  OR U14069 ( .A(n11747), .B(n11748), .Z(n11746) );
  OR U14070 ( .A(n11749), .B(n11750), .Z(n11745) );
  ANDN U14071 ( .B(n11751), .A(n11752), .Z(n11703) );
  IV U14072 ( .A(n11753), .Z(n11751) );
  ANDN U14073 ( .B(n11754), .A(n11755), .Z(n11695) );
  XOR U14074 ( .A(n11681), .B(n11756), .Z(n11693) );
  XOR U14075 ( .A(n11682), .B(n11683), .Z(n11756) );
  XOR U14076 ( .A(n11688), .B(n11757), .Z(n11683) );
  XOR U14077 ( .A(n11687), .B(n11690), .Z(n11757) );
  IV U14078 ( .A(n11689), .Z(n11690) );
  NAND U14079 ( .A(n11758), .B(n11759), .Z(n11689) );
  OR U14080 ( .A(n11760), .B(n11761), .Z(n11759) );
  OR U14081 ( .A(n11762), .B(n11763), .Z(n11758) );
  NAND U14082 ( .A(n11764), .B(n11765), .Z(n11687) );
  OR U14083 ( .A(n11766), .B(n11767), .Z(n11765) );
  OR U14084 ( .A(n11768), .B(n11769), .Z(n11764) );
  NOR U14085 ( .A(n11770), .B(n11771), .Z(n11688) );
  ANDN U14086 ( .B(n11772), .A(n11773), .Z(n11682) );
  IV U14087 ( .A(n11774), .Z(n11772) );
  XNOR U14088 ( .A(n11675), .B(n11775), .Z(n11681) );
  XNOR U14089 ( .A(n11674), .B(n11676), .Z(n11775) );
  NAND U14090 ( .A(n11776), .B(n11777), .Z(n11676) );
  OR U14091 ( .A(n11778), .B(n11779), .Z(n11777) );
  OR U14092 ( .A(n11780), .B(n11781), .Z(n11776) );
  NAND U14093 ( .A(n11782), .B(n11783), .Z(n11674) );
  OR U14094 ( .A(n11784), .B(n11785), .Z(n11783) );
  OR U14095 ( .A(n11786), .B(n11787), .Z(n11782) );
  ANDN U14096 ( .B(n11788), .A(n11789), .Z(n11675) );
  IV U14097 ( .A(n11790), .Z(n11788) );
  XNOR U14098 ( .A(n11755), .B(n11754), .Z(N12913) );
  XOR U14099 ( .A(n11774), .B(n11773), .Z(n11754) );
  XNOR U14100 ( .A(n11789), .B(n11790), .Z(n11773) );
  XNOR U14101 ( .A(n11784), .B(n11785), .Z(n11790) );
  XNOR U14102 ( .A(n11786), .B(n11787), .Z(n11785) );
  XNOR U14103 ( .A(y[301]), .B(x[301]), .Z(n11787) );
  XNOR U14104 ( .A(y[302]), .B(x[302]), .Z(n11786) );
  XNOR U14105 ( .A(y[300]), .B(x[300]), .Z(n11784) );
  XNOR U14106 ( .A(n11778), .B(n11779), .Z(n11789) );
  XNOR U14107 ( .A(y[297]), .B(x[297]), .Z(n11779) );
  XNOR U14108 ( .A(n11780), .B(n11781), .Z(n11778) );
  XNOR U14109 ( .A(y[298]), .B(x[298]), .Z(n11781) );
  XNOR U14110 ( .A(y[299]), .B(x[299]), .Z(n11780) );
  XNOR U14111 ( .A(n11771), .B(n11770), .Z(n11774) );
  XNOR U14112 ( .A(n11766), .B(n11767), .Z(n11770) );
  XNOR U14113 ( .A(y[294]), .B(x[294]), .Z(n11767) );
  XNOR U14114 ( .A(n11768), .B(n11769), .Z(n11766) );
  XNOR U14115 ( .A(y[295]), .B(x[295]), .Z(n11769) );
  XNOR U14116 ( .A(y[296]), .B(x[296]), .Z(n11768) );
  XNOR U14117 ( .A(n11760), .B(n11761), .Z(n11771) );
  XNOR U14118 ( .A(y[291]), .B(x[291]), .Z(n11761) );
  XNOR U14119 ( .A(n11762), .B(n11763), .Z(n11760) );
  XNOR U14120 ( .A(y[292]), .B(x[292]), .Z(n11763) );
  XNOR U14121 ( .A(y[293]), .B(x[293]), .Z(n11762) );
  XOR U14122 ( .A(n11736), .B(n11737), .Z(n11755) );
  XNOR U14123 ( .A(n11752), .B(n11753), .Z(n11737) );
  XNOR U14124 ( .A(n11747), .B(n11748), .Z(n11753) );
  XNOR U14125 ( .A(n11749), .B(n11750), .Z(n11748) );
  XNOR U14126 ( .A(y[289]), .B(x[289]), .Z(n11750) );
  XNOR U14127 ( .A(y[290]), .B(x[290]), .Z(n11749) );
  XNOR U14128 ( .A(y[288]), .B(x[288]), .Z(n11747) );
  XNOR U14129 ( .A(n11741), .B(n11742), .Z(n11752) );
  XNOR U14130 ( .A(y[285]), .B(x[285]), .Z(n11742) );
  XNOR U14131 ( .A(n11743), .B(n11744), .Z(n11741) );
  XNOR U14132 ( .A(y[286]), .B(x[286]), .Z(n11744) );
  XNOR U14133 ( .A(y[287]), .B(x[287]), .Z(n11743) );
  XOR U14134 ( .A(n11735), .B(n11734), .Z(n11736) );
  XNOR U14135 ( .A(n11730), .B(n11731), .Z(n11734) );
  XNOR U14136 ( .A(y[282]), .B(x[282]), .Z(n11731) );
  XNOR U14137 ( .A(n11732), .B(n11733), .Z(n11730) );
  XNOR U14138 ( .A(y[283]), .B(x[283]), .Z(n11733) );
  XNOR U14139 ( .A(y[284]), .B(x[284]), .Z(n11732) );
  XNOR U14140 ( .A(n11724), .B(n11725), .Z(n11735) );
  XNOR U14141 ( .A(y[279]), .B(x[279]), .Z(n11725) );
  XNOR U14142 ( .A(n11726), .B(n11727), .Z(n11724) );
  XNOR U14143 ( .A(y[280]), .B(x[280]), .Z(n11727) );
  XNOR U14144 ( .A(y[281]), .B(x[281]), .Z(n11726) );
  NAND U14145 ( .A(n11791), .B(n11792), .Z(N12906) );
  NANDN U14146 ( .A(n11793), .B(n11794), .Z(n11792) );
  OR U14147 ( .A(n11795), .B(n11796), .Z(n11794) );
  NAND U14148 ( .A(n11795), .B(n11796), .Z(n11791) );
  XOR U14149 ( .A(n11795), .B(n11797), .Z(N12905) );
  XNOR U14150 ( .A(n11793), .B(n11796), .Z(n11797) );
  AND U14151 ( .A(n11798), .B(n11799), .Z(n11796) );
  NANDN U14152 ( .A(n11800), .B(n11801), .Z(n11799) );
  NANDN U14153 ( .A(n11802), .B(n11803), .Z(n11801) );
  NANDN U14154 ( .A(n11803), .B(n11802), .Z(n11798) );
  NAND U14155 ( .A(n11804), .B(n11805), .Z(n11793) );
  NANDN U14156 ( .A(n11806), .B(n11807), .Z(n11805) );
  OR U14157 ( .A(n11808), .B(n11809), .Z(n11807) );
  NAND U14158 ( .A(n11809), .B(n11808), .Z(n11804) );
  AND U14159 ( .A(n11810), .B(n11811), .Z(n11795) );
  NANDN U14160 ( .A(n11812), .B(n11813), .Z(n11811) );
  NANDN U14161 ( .A(n11814), .B(n11815), .Z(n11813) );
  NANDN U14162 ( .A(n11815), .B(n11814), .Z(n11810) );
  XOR U14163 ( .A(n11809), .B(n11816), .Z(N12904) );
  XOR U14164 ( .A(n11806), .B(n11808), .Z(n11816) );
  XNOR U14165 ( .A(n11802), .B(n11817), .Z(n11808) );
  XNOR U14166 ( .A(n11800), .B(n11803), .Z(n11817) );
  NAND U14167 ( .A(n11818), .B(n11819), .Z(n11803) );
  NAND U14168 ( .A(n11820), .B(n11821), .Z(n11819) );
  OR U14169 ( .A(n11822), .B(n11823), .Z(n11820) );
  NANDN U14170 ( .A(n11824), .B(n11822), .Z(n11818) );
  IV U14171 ( .A(n11823), .Z(n11824) );
  NAND U14172 ( .A(n11825), .B(n11826), .Z(n11800) );
  NAND U14173 ( .A(n11827), .B(n11828), .Z(n11826) );
  NANDN U14174 ( .A(n11829), .B(n11830), .Z(n11827) );
  NANDN U14175 ( .A(n11830), .B(n11829), .Z(n11825) );
  AND U14176 ( .A(n11831), .B(n11832), .Z(n11802) );
  NAND U14177 ( .A(n11833), .B(n11834), .Z(n11832) );
  OR U14178 ( .A(n11835), .B(n11836), .Z(n11833) );
  NANDN U14179 ( .A(n11837), .B(n11835), .Z(n11831) );
  NAND U14180 ( .A(n11838), .B(n11839), .Z(n11806) );
  NANDN U14181 ( .A(n11840), .B(n11841), .Z(n11839) );
  OR U14182 ( .A(n11842), .B(n11843), .Z(n11841) );
  NANDN U14183 ( .A(n11844), .B(n11842), .Z(n11838) );
  IV U14184 ( .A(n11843), .Z(n11844) );
  XNOR U14185 ( .A(n11814), .B(n11845), .Z(n11809) );
  XNOR U14186 ( .A(n11812), .B(n11815), .Z(n11845) );
  NAND U14187 ( .A(n11846), .B(n11847), .Z(n11815) );
  NAND U14188 ( .A(n11848), .B(n11849), .Z(n11847) );
  OR U14189 ( .A(n11850), .B(n11851), .Z(n11848) );
  NANDN U14190 ( .A(n11852), .B(n11850), .Z(n11846) );
  IV U14191 ( .A(n11851), .Z(n11852) );
  NAND U14192 ( .A(n11853), .B(n11854), .Z(n11812) );
  NAND U14193 ( .A(n11855), .B(n11856), .Z(n11854) );
  NANDN U14194 ( .A(n11857), .B(n11858), .Z(n11855) );
  NANDN U14195 ( .A(n11858), .B(n11857), .Z(n11853) );
  AND U14196 ( .A(n11859), .B(n11860), .Z(n11814) );
  NAND U14197 ( .A(n11861), .B(n11862), .Z(n11860) );
  OR U14198 ( .A(n11863), .B(n11864), .Z(n11861) );
  NANDN U14199 ( .A(n11865), .B(n11863), .Z(n11859) );
  XNOR U14200 ( .A(n11840), .B(n11866), .Z(N12903) );
  XOR U14201 ( .A(n11842), .B(n11843), .Z(n11866) );
  XNOR U14202 ( .A(n11856), .B(n11867), .Z(n11843) );
  XOR U14203 ( .A(n11857), .B(n11858), .Z(n11867) );
  XOR U14204 ( .A(n11863), .B(n11868), .Z(n11858) );
  XOR U14205 ( .A(n11862), .B(n11865), .Z(n11868) );
  IV U14206 ( .A(n11864), .Z(n11865) );
  NAND U14207 ( .A(n11869), .B(n11870), .Z(n11864) );
  OR U14208 ( .A(n11871), .B(n11872), .Z(n11870) );
  OR U14209 ( .A(n11873), .B(n11874), .Z(n11869) );
  NAND U14210 ( .A(n11875), .B(n11876), .Z(n11862) );
  OR U14211 ( .A(n11877), .B(n11878), .Z(n11876) );
  OR U14212 ( .A(n11879), .B(n11880), .Z(n11875) );
  NOR U14213 ( .A(n11881), .B(n11882), .Z(n11863) );
  ANDN U14214 ( .B(n11883), .A(n11884), .Z(n11857) );
  XNOR U14215 ( .A(n11850), .B(n11885), .Z(n11856) );
  XNOR U14216 ( .A(n11849), .B(n11851), .Z(n11885) );
  NAND U14217 ( .A(n11886), .B(n11887), .Z(n11851) );
  OR U14218 ( .A(n11888), .B(n11889), .Z(n11887) );
  OR U14219 ( .A(n11890), .B(n11891), .Z(n11886) );
  NAND U14220 ( .A(n11892), .B(n11893), .Z(n11849) );
  OR U14221 ( .A(n11894), .B(n11895), .Z(n11893) );
  OR U14222 ( .A(n11896), .B(n11897), .Z(n11892) );
  ANDN U14223 ( .B(n11898), .A(n11899), .Z(n11850) );
  IV U14224 ( .A(n11900), .Z(n11898) );
  ANDN U14225 ( .B(n11901), .A(n11902), .Z(n11842) );
  XOR U14226 ( .A(n11828), .B(n11903), .Z(n11840) );
  XOR U14227 ( .A(n11829), .B(n11830), .Z(n11903) );
  XOR U14228 ( .A(n11835), .B(n11904), .Z(n11830) );
  XOR U14229 ( .A(n11834), .B(n11837), .Z(n11904) );
  IV U14230 ( .A(n11836), .Z(n11837) );
  NAND U14231 ( .A(n11905), .B(n11906), .Z(n11836) );
  OR U14232 ( .A(n11907), .B(n11908), .Z(n11906) );
  OR U14233 ( .A(n11909), .B(n11910), .Z(n11905) );
  NAND U14234 ( .A(n11911), .B(n11912), .Z(n11834) );
  OR U14235 ( .A(n11913), .B(n11914), .Z(n11912) );
  OR U14236 ( .A(n11915), .B(n11916), .Z(n11911) );
  NOR U14237 ( .A(n11917), .B(n11918), .Z(n11835) );
  ANDN U14238 ( .B(n11919), .A(n11920), .Z(n11829) );
  IV U14239 ( .A(n11921), .Z(n11919) );
  XNOR U14240 ( .A(n11822), .B(n11922), .Z(n11828) );
  XNOR U14241 ( .A(n11821), .B(n11823), .Z(n11922) );
  NAND U14242 ( .A(n11923), .B(n11924), .Z(n11823) );
  OR U14243 ( .A(n11925), .B(n11926), .Z(n11924) );
  OR U14244 ( .A(n11927), .B(n11928), .Z(n11923) );
  NAND U14245 ( .A(n11929), .B(n11930), .Z(n11821) );
  OR U14246 ( .A(n11931), .B(n11932), .Z(n11930) );
  OR U14247 ( .A(n11933), .B(n11934), .Z(n11929) );
  ANDN U14248 ( .B(n11935), .A(n11936), .Z(n11822) );
  IV U14249 ( .A(n11937), .Z(n11935) );
  XNOR U14250 ( .A(n11902), .B(n11901), .Z(N12902) );
  XOR U14251 ( .A(n11921), .B(n11920), .Z(n11901) );
  XNOR U14252 ( .A(n11936), .B(n11937), .Z(n11920) );
  XNOR U14253 ( .A(n11931), .B(n11932), .Z(n11937) );
  XNOR U14254 ( .A(n11933), .B(n11934), .Z(n11932) );
  XNOR U14255 ( .A(y[277]), .B(x[277]), .Z(n11934) );
  XNOR U14256 ( .A(y[278]), .B(x[278]), .Z(n11933) );
  XNOR U14257 ( .A(y[276]), .B(x[276]), .Z(n11931) );
  XNOR U14258 ( .A(n11925), .B(n11926), .Z(n11936) );
  XNOR U14259 ( .A(y[273]), .B(x[273]), .Z(n11926) );
  XNOR U14260 ( .A(n11927), .B(n11928), .Z(n11925) );
  XNOR U14261 ( .A(y[274]), .B(x[274]), .Z(n11928) );
  XNOR U14262 ( .A(y[275]), .B(x[275]), .Z(n11927) );
  XNOR U14263 ( .A(n11918), .B(n11917), .Z(n11921) );
  XNOR U14264 ( .A(n11913), .B(n11914), .Z(n11917) );
  XNOR U14265 ( .A(y[270]), .B(x[270]), .Z(n11914) );
  XNOR U14266 ( .A(n11915), .B(n11916), .Z(n11913) );
  XNOR U14267 ( .A(y[271]), .B(x[271]), .Z(n11916) );
  XNOR U14268 ( .A(y[272]), .B(x[272]), .Z(n11915) );
  XNOR U14269 ( .A(n11907), .B(n11908), .Z(n11918) );
  XNOR U14270 ( .A(y[267]), .B(x[267]), .Z(n11908) );
  XNOR U14271 ( .A(n11909), .B(n11910), .Z(n11907) );
  XNOR U14272 ( .A(y[268]), .B(x[268]), .Z(n11910) );
  XNOR U14273 ( .A(y[269]), .B(x[269]), .Z(n11909) );
  XOR U14274 ( .A(n11883), .B(n11884), .Z(n11902) );
  XNOR U14275 ( .A(n11899), .B(n11900), .Z(n11884) );
  XNOR U14276 ( .A(n11894), .B(n11895), .Z(n11900) );
  XNOR U14277 ( .A(n11896), .B(n11897), .Z(n11895) );
  XNOR U14278 ( .A(y[265]), .B(x[265]), .Z(n11897) );
  XNOR U14279 ( .A(y[266]), .B(x[266]), .Z(n11896) );
  XNOR U14280 ( .A(y[264]), .B(x[264]), .Z(n11894) );
  XNOR U14281 ( .A(n11888), .B(n11889), .Z(n11899) );
  XNOR U14282 ( .A(y[261]), .B(x[261]), .Z(n11889) );
  XNOR U14283 ( .A(n11890), .B(n11891), .Z(n11888) );
  XNOR U14284 ( .A(y[262]), .B(x[262]), .Z(n11891) );
  XNOR U14285 ( .A(y[263]), .B(x[263]), .Z(n11890) );
  XOR U14286 ( .A(n11882), .B(n11881), .Z(n11883) );
  XNOR U14287 ( .A(n11877), .B(n11878), .Z(n11881) );
  XNOR U14288 ( .A(y[258]), .B(x[258]), .Z(n11878) );
  XNOR U14289 ( .A(n11879), .B(n11880), .Z(n11877) );
  XNOR U14290 ( .A(y[259]), .B(x[259]), .Z(n11880) );
  XNOR U14291 ( .A(y[260]), .B(x[260]), .Z(n11879) );
  XNOR U14292 ( .A(n11871), .B(n11872), .Z(n11882) );
  XNOR U14293 ( .A(y[255]), .B(x[255]), .Z(n11872) );
  XNOR U14294 ( .A(n11873), .B(n11874), .Z(n11871) );
  XNOR U14295 ( .A(y[256]), .B(x[256]), .Z(n11874) );
  XNOR U14296 ( .A(y[257]), .B(x[257]), .Z(n11873) );
  NAND U14297 ( .A(n11938), .B(n11939), .Z(N12895) );
  NANDN U14298 ( .A(n11940), .B(n11941), .Z(n11939) );
  OR U14299 ( .A(n11942), .B(n11943), .Z(n11941) );
  NAND U14300 ( .A(n11942), .B(n11943), .Z(n11938) );
  XOR U14301 ( .A(n11942), .B(n11944), .Z(N12894) );
  XNOR U14302 ( .A(n11940), .B(n11943), .Z(n11944) );
  AND U14303 ( .A(n11945), .B(n11946), .Z(n11943) );
  NANDN U14304 ( .A(n11947), .B(n11948), .Z(n11946) );
  NANDN U14305 ( .A(n11949), .B(n11950), .Z(n11948) );
  NANDN U14306 ( .A(n11950), .B(n11949), .Z(n11945) );
  NAND U14307 ( .A(n11951), .B(n11952), .Z(n11940) );
  NANDN U14308 ( .A(n11953), .B(n11954), .Z(n11952) );
  OR U14309 ( .A(n11955), .B(n11956), .Z(n11954) );
  NAND U14310 ( .A(n11956), .B(n11955), .Z(n11951) );
  AND U14311 ( .A(n11957), .B(n11958), .Z(n11942) );
  NANDN U14312 ( .A(n11959), .B(n11960), .Z(n11958) );
  NANDN U14313 ( .A(n11961), .B(n11962), .Z(n11960) );
  NANDN U14314 ( .A(n11962), .B(n11961), .Z(n11957) );
  XOR U14315 ( .A(n11956), .B(n11963), .Z(N12893) );
  XOR U14316 ( .A(n11953), .B(n11955), .Z(n11963) );
  XNOR U14317 ( .A(n11949), .B(n11964), .Z(n11955) );
  XNOR U14318 ( .A(n11947), .B(n11950), .Z(n11964) );
  NAND U14319 ( .A(n11965), .B(n11966), .Z(n11950) );
  NAND U14320 ( .A(n11967), .B(n11968), .Z(n11966) );
  OR U14321 ( .A(n11969), .B(n11970), .Z(n11967) );
  NANDN U14322 ( .A(n11971), .B(n11969), .Z(n11965) );
  IV U14323 ( .A(n11970), .Z(n11971) );
  NAND U14324 ( .A(n11972), .B(n11973), .Z(n11947) );
  NAND U14325 ( .A(n11974), .B(n11975), .Z(n11973) );
  NANDN U14326 ( .A(n11976), .B(n11977), .Z(n11974) );
  NANDN U14327 ( .A(n11977), .B(n11976), .Z(n11972) );
  AND U14328 ( .A(n11978), .B(n11979), .Z(n11949) );
  NAND U14329 ( .A(n11980), .B(n11981), .Z(n11979) );
  OR U14330 ( .A(n11982), .B(n11983), .Z(n11980) );
  NANDN U14331 ( .A(n11984), .B(n11982), .Z(n11978) );
  NAND U14332 ( .A(n11985), .B(n11986), .Z(n11953) );
  NANDN U14333 ( .A(n11987), .B(n11988), .Z(n11986) );
  OR U14334 ( .A(n11989), .B(n11990), .Z(n11988) );
  NANDN U14335 ( .A(n11991), .B(n11989), .Z(n11985) );
  IV U14336 ( .A(n11990), .Z(n11991) );
  XNOR U14337 ( .A(n11961), .B(n11992), .Z(n11956) );
  XNOR U14338 ( .A(n11959), .B(n11962), .Z(n11992) );
  NAND U14339 ( .A(n11993), .B(n11994), .Z(n11962) );
  NAND U14340 ( .A(n11995), .B(n11996), .Z(n11994) );
  OR U14341 ( .A(n11997), .B(n11998), .Z(n11995) );
  NANDN U14342 ( .A(n11999), .B(n11997), .Z(n11993) );
  IV U14343 ( .A(n11998), .Z(n11999) );
  NAND U14344 ( .A(n12000), .B(n12001), .Z(n11959) );
  NAND U14345 ( .A(n12002), .B(n12003), .Z(n12001) );
  NANDN U14346 ( .A(n12004), .B(n12005), .Z(n12002) );
  NANDN U14347 ( .A(n12005), .B(n12004), .Z(n12000) );
  AND U14348 ( .A(n12006), .B(n12007), .Z(n11961) );
  NAND U14349 ( .A(n12008), .B(n12009), .Z(n12007) );
  OR U14350 ( .A(n12010), .B(n12011), .Z(n12008) );
  NANDN U14351 ( .A(n12012), .B(n12010), .Z(n12006) );
  XNOR U14352 ( .A(n11987), .B(n12013), .Z(N12892) );
  XOR U14353 ( .A(n11989), .B(n11990), .Z(n12013) );
  XNOR U14354 ( .A(n12003), .B(n12014), .Z(n11990) );
  XOR U14355 ( .A(n12004), .B(n12005), .Z(n12014) );
  XOR U14356 ( .A(n12010), .B(n12015), .Z(n12005) );
  XOR U14357 ( .A(n12009), .B(n12012), .Z(n12015) );
  IV U14358 ( .A(n12011), .Z(n12012) );
  NAND U14359 ( .A(n12016), .B(n12017), .Z(n12011) );
  OR U14360 ( .A(n12018), .B(n12019), .Z(n12017) );
  OR U14361 ( .A(n12020), .B(n12021), .Z(n12016) );
  NAND U14362 ( .A(n12022), .B(n12023), .Z(n12009) );
  OR U14363 ( .A(n12024), .B(n12025), .Z(n12023) );
  OR U14364 ( .A(n12026), .B(n12027), .Z(n12022) );
  NOR U14365 ( .A(n12028), .B(n12029), .Z(n12010) );
  ANDN U14366 ( .B(n12030), .A(n12031), .Z(n12004) );
  XNOR U14367 ( .A(n11997), .B(n12032), .Z(n12003) );
  XNOR U14368 ( .A(n11996), .B(n11998), .Z(n12032) );
  NAND U14369 ( .A(n12033), .B(n12034), .Z(n11998) );
  OR U14370 ( .A(n12035), .B(n12036), .Z(n12034) );
  OR U14371 ( .A(n12037), .B(n12038), .Z(n12033) );
  NAND U14372 ( .A(n12039), .B(n12040), .Z(n11996) );
  OR U14373 ( .A(n12041), .B(n12042), .Z(n12040) );
  OR U14374 ( .A(n12043), .B(n12044), .Z(n12039) );
  ANDN U14375 ( .B(n12045), .A(n12046), .Z(n11997) );
  IV U14376 ( .A(n12047), .Z(n12045) );
  ANDN U14377 ( .B(n12048), .A(n12049), .Z(n11989) );
  XOR U14378 ( .A(n11975), .B(n12050), .Z(n11987) );
  XOR U14379 ( .A(n11976), .B(n11977), .Z(n12050) );
  XOR U14380 ( .A(n11982), .B(n12051), .Z(n11977) );
  XOR U14381 ( .A(n11981), .B(n11984), .Z(n12051) );
  IV U14382 ( .A(n11983), .Z(n11984) );
  NAND U14383 ( .A(n12052), .B(n12053), .Z(n11983) );
  OR U14384 ( .A(n12054), .B(n12055), .Z(n12053) );
  OR U14385 ( .A(n12056), .B(n12057), .Z(n12052) );
  NAND U14386 ( .A(n12058), .B(n12059), .Z(n11981) );
  OR U14387 ( .A(n12060), .B(n12061), .Z(n12059) );
  OR U14388 ( .A(n12062), .B(n12063), .Z(n12058) );
  NOR U14389 ( .A(n12064), .B(n12065), .Z(n11982) );
  ANDN U14390 ( .B(n12066), .A(n12067), .Z(n11976) );
  IV U14391 ( .A(n12068), .Z(n12066) );
  XNOR U14392 ( .A(n11969), .B(n12069), .Z(n11975) );
  XNOR U14393 ( .A(n11968), .B(n11970), .Z(n12069) );
  NAND U14394 ( .A(n12070), .B(n12071), .Z(n11970) );
  OR U14395 ( .A(n12072), .B(n12073), .Z(n12071) );
  OR U14396 ( .A(n12074), .B(n12075), .Z(n12070) );
  NAND U14397 ( .A(n12076), .B(n12077), .Z(n11968) );
  OR U14398 ( .A(n12078), .B(n12079), .Z(n12077) );
  OR U14399 ( .A(n12080), .B(n12081), .Z(n12076) );
  ANDN U14400 ( .B(n12082), .A(n12083), .Z(n11969) );
  IV U14401 ( .A(n12084), .Z(n12082) );
  XNOR U14402 ( .A(n12049), .B(n12048), .Z(N12891) );
  XOR U14403 ( .A(n12068), .B(n12067), .Z(n12048) );
  XNOR U14404 ( .A(n12083), .B(n12084), .Z(n12067) );
  XNOR U14405 ( .A(n12078), .B(n12079), .Z(n12084) );
  XNOR U14406 ( .A(n12080), .B(n12081), .Z(n12079) );
  XNOR U14407 ( .A(y[253]), .B(x[253]), .Z(n12081) );
  XNOR U14408 ( .A(y[254]), .B(x[254]), .Z(n12080) );
  XNOR U14409 ( .A(y[252]), .B(x[252]), .Z(n12078) );
  XNOR U14410 ( .A(n12072), .B(n12073), .Z(n12083) );
  XNOR U14411 ( .A(y[249]), .B(x[249]), .Z(n12073) );
  XNOR U14412 ( .A(n12074), .B(n12075), .Z(n12072) );
  XNOR U14413 ( .A(y[250]), .B(x[250]), .Z(n12075) );
  XNOR U14414 ( .A(y[251]), .B(x[251]), .Z(n12074) );
  XNOR U14415 ( .A(n12065), .B(n12064), .Z(n12068) );
  XNOR U14416 ( .A(n12060), .B(n12061), .Z(n12064) );
  XNOR U14417 ( .A(y[246]), .B(x[246]), .Z(n12061) );
  XNOR U14418 ( .A(n12062), .B(n12063), .Z(n12060) );
  XNOR U14419 ( .A(y[247]), .B(x[247]), .Z(n12063) );
  XNOR U14420 ( .A(y[248]), .B(x[248]), .Z(n12062) );
  XNOR U14421 ( .A(n12054), .B(n12055), .Z(n12065) );
  XNOR U14422 ( .A(y[243]), .B(x[243]), .Z(n12055) );
  XNOR U14423 ( .A(n12056), .B(n12057), .Z(n12054) );
  XNOR U14424 ( .A(y[244]), .B(x[244]), .Z(n12057) );
  XNOR U14425 ( .A(y[245]), .B(x[245]), .Z(n12056) );
  XOR U14426 ( .A(n12030), .B(n12031), .Z(n12049) );
  XNOR U14427 ( .A(n12046), .B(n12047), .Z(n12031) );
  XNOR U14428 ( .A(n12041), .B(n12042), .Z(n12047) );
  XNOR U14429 ( .A(n12043), .B(n12044), .Z(n12042) );
  XNOR U14430 ( .A(y[241]), .B(x[241]), .Z(n12044) );
  XNOR U14431 ( .A(y[242]), .B(x[242]), .Z(n12043) );
  XNOR U14432 ( .A(y[240]), .B(x[240]), .Z(n12041) );
  XNOR U14433 ( .A(n12035), .B(n12036), .Z(n12046) );
  XNOR U14434 ( .A(y[237]), .B(x[237]), .Z(n12036) );
  XNOR U14435 ( .A(n12037), .B(n12038), .Z(n12035) );
  XNOR U14436 ( .A(y[238]), .B(x[238]), .Z(n12038) );
  XNOR U14437 ( .A(y[239]), .B(x[239]), .Z(n12037) );
  XOR U14438 ( .A(n12029), .B(n12028), .Z(n12030) );
  XNOR U14439 ( .A(n12024), .B(n12025), .Z(n12028) );
  XNOR U14440 ( .A(y[234]), .B(x[234]), .Z(n12025) );
  XNOR U14441 ( .A(n12026), .B(n12027), .Z(n12024) );
  XNOR U14442 ( .A(y[235]), .B(x[235]), .Z(n12027) );
  XNOR U14443 ( .A(y[236]), .B(x[236]), .Z(n12026) );
  XNOR U14444 ( .A(n12018), .B(n12019), .Z(n12029) );
  XNOR U14445 ( .A(y[231]), .B(x[231]), .Z(n12019) );
  XNOR U14446 ( .A(n12020), .B(n12021), .Z(n12018) );
  XNOR U14447 ( .A(y[232]), .B(x[232]), .Z(n12021) );
  XNOR U14448 ( .A(y[233]), .B(x[233]), .Z(n12020) );
  NAND U14449 ( .A(n12085), .B(n12086), .Z(N12884) );
  NANDN U14450 ( .A(n12087), .B(n12088), .Z(n12086) );
  OR U14451 ( .A(n12089), .B(n12090), .Z(n12088) );
  NAND U14452 ( .A(n12089), .B(n12090), .Z(n12085) );
  XOR U14453 ( .A(n12089), .B(n12091), .Z(N12883) );
  XNOR U14454 ( .A(n12087), .B(n12090), .Z(n12091) );
  AND U14455 ( .A(n12092), .B(n12093), .Z(n12090) );
  NANDN U14456 ( .A(n12094), .B(n12095), .Z(n12093) );
  NANDN U14457 ( .A(n12096), .B(n12097), .Z(n12095) );
  NANDN U14458 ( .A(n12097), .B(n12096), .Z(n12092) );
  NAND U14459 ( .A(n12098), .B(n12099), .Z(n12087) );
  NANDN U14460 ( .A(n12100), .B(n12101), .Z(n12099) );
  OR U14461 ( .A(n12102), .B(n12103), .Z(n12101) );
  NAND U14462 ( .A(n12103), .B(n12102), .Z(n12098) );
  AND U14463 ( .A(n12104), .B(n12105), .Z(n12089) );
  NANDN U14464 ( .A(n12106), .B(n12107), .Z(n12105) );
  NANDN U14465 ( .A(n12108), .B(n12109), .Z(n12107) );
  NANDN U14466 ( .A(n12109), .B(n12108), .Z(n12104) );
  XOR U14467 ( .A(n12103), .B(n12110), .Z(N12882) );
  XOR U14468 ( .A(n12100), .B(n12102), .Z(n12110) );
  XNOR U14469 ( .A(n12096), .B(n12111), .Z(n12102) );
  XNOR U14470 ( .A(n12094), .B(n12097), .Z(n12111) );
  NAND U14471 ( .A(n12112), .B(n12113), .Z(n12097) );
  NAND U14472 ( .A(n12114), .B(n12115), .Z(n12113) );
  OR U14473 ( .A(n12116), .B(n12117), .Z(n12114) );
  NANDN U14474 ( .A(n12118), .B(n12116), .Z(n12112) );
  IV U14475 ( .A(n12117), .Z(n12118) );
  NAND U14476 ( .A(n12119), .B(n12120), .Z(n12094) );
  NAND U14477 ( .A(n12121), .B(n12122), .Z(n12120) );
  NANDN U14478 ( .A(n12123), .B(n12124), .Z(n12121) );
  NANDN U14479 ( .A(n12124), .B(n12123), .Z(n12119) );
  AND U14480 ( .A(n12125), .B(n12126), .Z(n12096) );
  NAND U14481 ( .A(n12127), .B(n12128), .Z(n12126) );
  OR U14482 ( .A(n12129), .B(n12130), .Z(n12127) );
  NANDN U14483 ( .A(n12131), .B(n12129), .Z(n12125) );
  NAND U14484 ( .A(n12132), .B(n12133), .Z(n12100) );
  NANDN U14485 ( .A(n12134), .B(n12135), .Z(n12133) );
  OR U14486 ( .A(n12136), .B(n12137), .Z(n12135) );
  NANDN U14487 ( .A(n12138), .B(n12136), .Z(n12132) );
  IV U14488 ( .A(n12137), .Z(n12138) );
  XNOR U14489 ( .A(n12108), .B(n12139), .Z(n12103) );
  XNOR U14490 ( .A(n12106), .B(n12109), .Z(n12139) );
  NAND U14491 ( .A(n12140), .B(n12141), .Z(n12109) );
  NAND U14492 ( .A(n12142), .B(n12143), .Z(n12141) );
  OR U14493 ( .A(n12144), .B(n12145), .Z(n12142) );
  NANDN U14494 ( .A(n12146), .B(n12144), .Z(n12140) );
  IV U14495 ( .A(n12145), .Z(n12146) );
  NAND U14496 ( .A(n12147), .B(n12148), .Z(n12106) );
  NAND U14497 ( .A(n12149), .B(n12150), .Z(n12148) );
  NANDN U14498 ( .A(n12151), .B(n12152), .Z(n12149) );
  NANDN U14499 ( .A(n12152), .B(n12151), .Z(n12147) );
  AND U14500 ( .A(n12153), .B(n12154), .Z(n12108) );
  NAND U14501 ( .A(n12155), .B(n12156), .Z(n12154) );
  OR U14502 ( .A(n12157), .B(n12158), .Z(n12155) );
  NANDN U14503 ( .A(n12159), .B(n12157), .Z(n12153) );
  XNOR U14504 ( .A(n12134), .B(n12160), .Z(N12881) );
  XOR U14505 ( .A(n12136), .B(n12137), .Z(n12160) );
  XNOR U14506 ( .A(n12150), .B(n12161), .Z(n12137) );
  XOR U14507 ( .A(n12151), .B(n12152), .Z(n12161) );
  XOR U14508 ( .A(n12157), .B(n12162), .Z(n12152) );
  XOR U14509 ( .A(n12156), .B(n12159), .Z(n12162) );
  IV U14510 ( .A(n12158), .Z(n12159) );
  NAND U14511 ( .A(n12163), .B(n12164), .Z(n12158) );
  OR U14512 ( .A(n12165), .B(n12166), .Z(n12164) );
  OR U14513 ( .A(n12167), .B(n12168), .Z(n12163) );
  NAND U14514 ( .A(n12169), .B(n12170), .Z(n12156) );
  OR U14515 ( .A(n12171), .B(n12172), .Z(n12170) );
  OR U14516 ( .A(n12173), .B(n12174), .Z(n12169) );
  NOR U14517 ( .A(n12175), .B(n12176), .Z(n12157) );
  ANDN U14518 ( .B(n12177), .A(n12178), .Z(n12151) );
  XNOR U14519 ( .A(n12144), .B(n12179), .Z(n12150) );
  XNOR U14520 ( .A(n12143), .B(n12145), .Z(n12179) );
  NAND U14521 ( .A(n12180), .B(n12181), .Z(n12145) );
  OR U14522 ( .A(n12182), .B(n12183), .Z(n12181) );
  OR U14523 ( .A(n12184), .B(n12185), .Z(n12180) );
  NAND U14524 ( .A(n12186), .B(n12187), .Z(n12143) );
  OR U14525 ( .A(n12188), .B(n12189), .Z(n12187) );
  OR U14526 ( .A(n12190), .B(n12191), .Z(n12186) );
  ANDN U14527 ( .B(n12192), .A(n12193), .Z(n12144) );
  IV U14528 ( .A(n12194), .Z(n12192) );
  ANDN U14529 ( .B(n12195), .A(n12196), .Z(n12136) );
  XOR U14530 ( .A(n12122), .B(n12197), .Z(n12134) );
  XOR U14531 ( .A(n12123), .B(n12124), .Z(n12197) );
  XOR U14532 ( .A(n12129), .B(n12198), .Z(n12124) );
  XOR U14533 ( .A(n12128), .B(n12131), .Z(n12198) );
  IV U14534 ( .A(n12130), .Z(n12131) );
  NAND U14535 ( .A(n12199), .B(n12200), .Z(n12130) );
  OR U14536 ( .A(n12201), .B(n12202), .Z(n12200) );
  OR U14537 ( .A(n12203), .B(n12204), .Z(n12199) );
  NAND U14538 ( .A(n12205), .B(n12206), .Z(n12128) );
  OR U14539 ( .A(n12207), .B(n12208), .Z(n12206) );
  OR U14540 ( .A(n12209), .B(n12210), .Z(n12205) );
  NOR U14541 ( .A(n12211), .B(n12212), .Z(n12129) );
  ANDN U14542 ( .B(n12213), .A(n12214), .Z(n12123) );
  IV U14543 ( .A(n12215), .Z(n12213) );
  XNOR U14544 ( .A(n12116), .B(n12216), .Z(n12122) );
  XNOR U14545 ( .A(n12115), .B(n12117), .Z(n12216) );
  NAND U14546 ( .A(n12217), .B(n12218), .Z(n12117) );
  OR U14547 ( .A(n12219), .B(n12220), .Z(n12218) );
  OR U14548 ( .A(n12221), .B(n12222), .Z(n12217) );
  NAND U14549 ( .A(n12223), .B(n12224), .Z(n12115) );
  OR U14550 ( .A(n12225), .B(n12226), .Z(n12224) );
  OR U14551 ( .A(n12227), .B(n12228), .Z(n12223) );
  ANDN U14552 ( .B(n12229), .A(n12230), .Z(n12116) );
  IV U14553 ( .A(n12231), .Z(n12229) );
  XNOR U14554 ( .A(n12196), .B(n12195), .Z(N12880) );
  XOR U14555 ( .A(n12215), .B(n12214), .Z(n12195) );
  XNOR U14556 ( .A(n12230), .B(n12231), .Z(n12214) );
  XNOR U14557 ( .A(n12225), .B(n12226), .Z(n12231) );
  XNOR U14558 ( .A(n12227), .B(n12228), .Z(n12226) );
  XNOR U14559 ( .A(y[229]), .B(x[229]), .Z(n12228) );
  XNOR U14560 ( .A(y[230]), .B(x[230]), .Z(n12227) );
  XNOR U14561 ( .A(y[228]), .B(x[228]), .Z(n12225) );
  XNOR U14562 ( .A(n12219), .B(n12220), .Z(n12230) );
  XNOR U14563 ( .A(y[225]), .B(x[225]), .Z(n12220) );
  XNOR U14564 ( .A(n12221), .B(n12222), .Z(n12219) );
  XNOR U14565 ( .A(y[226]), .B(x[226]), .Z(n12222) );
  XNOR U14566 ( .A(y[227]), .B(x[227]), .Z(n12221) );
  XNOR U14567 ( .A(n12212), .B(n12211), .Z(n12215) );
  XNOR U14568 ( .A(n12207), .B(n12208), .Z(n12211) );
  XNOR U14569 ( .A(y[222]), .B(x[222]), .Z(n12208) );
  XNOR U14570 ( .A(n12209), .B(n12210), .Z(n12207) );
  XNOR U14571 ( .A(y[223]), .B(x[223]), .Z(n12210) );
  XNOR U14572 ( .A(y[224]), .B(x[224]), .Z(n12209) );
  XNOR U14573 ( .A(n12201), .B(n12202), .Z(n12212) );
  XNOR U14574 ( .A(y[219]), .B(x[219]), .Z(n12202) );
  XNOR U14575 ( .A(n12203), .B(n12204), .Z(n12201) );
  XNOR U14576 ( .A(y[220]), .B(x[220]), .Z(n12204) );
  XNOR U14577 ( .A(y[221]), .B(x[221]), .Z(n12203) );
  XOR U14578 ( .A(n12177), .B(n12178), .Z(n12196) );
  XNOR U14579 ( .A(n12193), .B(n12194), .Z(n12178) );
  XNOR U14580 ( .A(n12188), .B(n12189), .Z(n12194) );
  XNOR U14581 ( .A(n12190), .B(n12191), .Z(n12189) );
  XNOR U14582 ( .A(y[217]), .B(x[217]), .Z(n12191) );
  XNOR U14583 ( .A(y[218]), .B(x[218]), .Z(n12190) );
  XNOR U14584 ( .A(y[216]), .B(x[216]), .Z(n12188) );
  XNOR U14585 ( .A(n12182), .B(n12183), .Z(n12193) );
  XNOR U14586 ( .A(y[213]), .B(x[213]), .Z(n12183) );
  XNOR U14587 ( .A(n12184), .B(n12185), .Z(n12182) );
  XNOR U14588 ( .A(y[214]), .B(x[214]), .Z(n12185) );
  XNOR U14589 ( .A(y[215]), .B(x[215]), .Z(n12184) );
  XOR U14590 ( .A(n12176), .B(n12175), .Z(n12177) );
  XNOR U14591 ( .A(n12171), .B(n12172), .Z(n12175) );
  XNOR U14592 ( .A(y[210]), .B(x[210]), .Z(n12172) );
  XNOR U14593 ( .A(n12173), .B(n12174), .Z(n12171) );
  XNOR U14594 ( .A(y[211]), .B(x[211]), .Z(n12174) );
  XNOR U14595 ( .A(y[212]), .B(x[212]), .Z(n12173) );
  XNOR U14596 ( .A(n12165), .B(n12166), .Z(n12176) );
  XNOR U14597 ( .A(y[207]), .B(x[207]), .Z(n12166) );
  XNOR U14598 ( .A(n12167), .B(n12168), .Z(n12165) );
  XNOR U14599 ( .A(y[208]), .B(x[208]), .Z(n12168) );
  XNOR U14600 ( .A(y[209]), .B(x[209]), .Z(n12167) );
  NAND U14601 ( .A(n12232), .B(n12233), .Z(N12873) );
  NANDN U14602 ( .A(n12234), .B(n12235), .Z(n12233) );
  OR U14603 ( .A(n12236), .B(n12237), .Z(n12235) );
  NAND U14604 ( .A(n12236), .B(n12237), .Z(n12232) );
  XOR U14605 ( .A(n12236), .B(n12238), .Z(N12872) );
  XNOR U14606 ( .A(n12234), .B(n12237), .Z(n12238) );
  AND U14607 ( .A(n12239), .B(n12240), .Z(n12237) );
  NANDN U14608 ( .A(n12241), .B(n12242), .Z(n12240) );
  NANDN U14609 ( .A(n12243), .B(n12244), .Z(n12242) );
  NANDN U14610 ( .A(n12244), .B(n12243), .Z(n12239) );
  NAND U14611 ( .A(n12245), .B(n12246), .Z(n12234) );
  NANDN U14612 ( .A(n12247), .B(n12248), .Z(n12246) );
  OR U14613 ( .A(n12249), .B(n12250), .Z(n12248) );
  NAND U14614 ( .A(n12250), .B(n12249), .Z(n12245) );
  AND U14615 ( .A(n12251), .B(n12252), .Z(n12236) );
  NANDN U14616 ( .A(n12253), .B(n12254), .Z(n12252) );
  NANDN U14617 ( .A(n12255), .B(n12256), .Z(n12254) );
  NANDN U14618 ( .A(n12256), .B(n12255), .Z(n12251) );
  XOR U14619 ( .A(n12250), .B(n12257), .Z(N12871) );
  XOR U14620 ( .A(n12247), .B(n12249), .Z(n12257) );
  XNOR U14621 ( .A(n12243), .B(n12258), .Z(n12249) );
  XNOR U14622 ( .A(n12241), .B(n12244), .Z(n12258) );
  NAND U14623 ( .A(n12259), .B(n12260), .Z(n12244) );
  NAND U14624 ( .A(n12261), .B(n12262), .Z(n12260) );
  OR U14625 ( .A(n12263), .B(n12264), .Z(n12261) );
  NANDN U14626 ( .A(n12265), .B(n12263), .Z(n12259) );
  IV U14627 ( .A(n12264), .Z(n12265) );
  NAND U14628 ( .A(n12266), .B(n12267), .Z(n12241) );
  NAND U14629 ( .A(n12268), .B(n12269), .Z(n12267) );
  NANDN U14630 ( .A(n12270), .B(n12271), .Z(n12268) );
  NANDN U14631 ( .A(n12271), .B(n12270), .Z(n12266) );
  AND U14632 ( .A(n12272), .B(n12273), .Z(n12243) );
  NAND U14633 ( .A(n12274), .B(n12275), .Z(n12273) );
  OR U14634 ( .A(n12276), .B(n12277), .Z(n12274) );
  NANDN U14635 ( .A(n12278), .B(n12276), .Z(n12272) );
  NAND U14636 ( .A(n12279), .B(n12280), .Z(n12247) );
  NANDN U14637 ( .A(n12281), .B(n12282), .Z(n12280) );
  OR U14638 ( .A(n12283), .B(n12284), .Z(n12282) );
  NANDN U14639 ( .A(n12285), .B(n12283), .Z(n12279) );
  IV U14640 ( .A(n12284), .Z(n12285) );
  XNOR U14641 ( .A(n12255), .B(n12286), .Z(n12250) );
  XNOR U14642 ( .A(n12253), .B(n12256), .Z(n12286) );
  NAND U14643 ( .A(n12287), .B(n12288), .Z(n12256) );
  NAND U14644 ( .A(n12289), .B(n12290), .Z(n12288) );
  OR U14645 ( .A(n12291), .B(n12292), .Z(n12289) );
  NANDN U14646 ( .A(n12293), .B(n12291), .Z(n12287) );
  IV U14647 ( .A(n12292), .Z(n12293) );
  NAND U14648 ( .A(n12294), .B(n12295), .Z(n12253) );
  NAND U14649 ( .A(n12296), .B(n12297), .Z(n12295) );
  NANDN U14650 ( .A(n12298), .B(n12299), .Z(n12296) );
  NANDN U14651 ( .A(n12299), .B(n12298), .Z(n12294) );
  AND U14652 ( .A(n12300), .B(n12301), .Z(n12255) );
  NAND U14653 ( .A(n12302), .B(n12303), .Z(n12301) );
  OR U14654 ( .A(n12304), .B(n12305), .Z(n12302) );
  NANDN U14655 ( .A(n12306), .B(n12304), .Z(n12300) );
  XNOR U14656 ( .A(n12281), .B(n12307), .Z(N12870) );
  XOR U14657 ( .A(n12283), .B(n12284), .Z(n12307) );
  XNOR U14658 ( .A(n12297), .B(n12308), .Z(n12284) );
  XOR U14659 ( .A(n12298), .B(n12299), .Z(n12308) );
  XOR U14660 ( .A(n12304), .B(n12309), .Z(n12299) );
  XOR U14661 ( .A(n12303), .B(n12306), .Z(n12309) );
  IV U14662 ( .A(n12305), .Z(n12306) );
  NAND U14663 ( .A(n12310), .B(n12311), .Z(n12305) );
  OR U14664 ( .A(n12312), .B(n12313), .Z(n12311) );
  OR U14665 ( .A(n12314), .B(n12315), .Z(n12310) );
  NAND U14666 ( .A(n12316), .B(n12317), .Z(n12303) );
  OR U14667 ( .A(n12318), .B(n12319), .Z(n12317) );
  OR U14668 ( .A(n12320), .B(n12321), .Z(n12316) );
  NOR U14669 ( .A(n12322), .B(n12323), .Z(n12304) );
  ANDN U14670 ( .B(n12324), .A(n12325), .Z(n12298) );
  XNOR U14671 ( .A(n12291), .B(n12326), .Z(n12297) );
  XNOR U14672 ( .A(n12290), .B(n12292), .Z(n12326) );
  NAND U14673 ( .A(n12327), .B(n12328), .Z(n12292) );
  OR U14674 ( .A(n12329), .B(n12330), .Z(n12328) );
  OR U14675 ( .A(n12331), .B(n12332), .Z(n12327) );
  NAND U14676 ( .A(n12333), .B(n12334), .Z(n12290) );
  OR U14677 ( .A(n12335), .B(n12336), .Z(n12334) );
  OR U14678 ( .A(n12337), .B(n12338), .Z(n12333) );
  ANDN U14679 ( .B(n12339), .A(n12340), .Z(n12291) );
  IV U14680 ( .A(n12341), .Z(n12339) );
  ANDN U14681 ( .B(n12342), .A(n12343), .Z(n12283) );
  XOR U14682 ( .A(n12269), .B(n12344), .Z(n12281) );
  XOR U14683 ( .A(n12270), .B(n12271), .Z(n12344) );
  XOR U14684 ( .A(n12276), .B(n12345), .Z(n12271) );
  XOR U14685 ( .A(n12275), .B(n12278), .Z(n12345) );
  IV U14686 ( .A(n12277), .Z(n12278) );
  NAND U14687 ( .A(n12346), .B(n12347), .Z(n12277) );
  OR U14688 ( .A(n12348), .B(n12349), .Z(n12347) );
  OR U14689 ( .A(n12350), .B(n12351), .Z(n12346) );
  NAND U14690 ( .A(n12352), .B(n12353), .Z(n12275) );
  OR U14691 ( .A(n12354), .B(n12355), .Z(n12353) );
  OR U14692 ( .A(n12356), .B(n12357), .Z(n12352) );
  NOR U14693 ( .A(n12358), .B(n12359), .Z(n12276) );
  ANDN U14694 ( .B(n12360), .A(n12361), .Z(n12270) );
  IV U14695 ( .A(n12362), .Z(n12360) );
  XNOR U14696 ( .A(n12263), .B(n12363), .Z(n12269) );
  XNOR U14697 ( .A(n12262), .B(n12264), .Z(n12363) );
  NAND U14698 ( .A(n12364), .B(n12365), .Z(n12264) );
  OR U14699 ( .A(n12366), .B(n12367), .Z(n12365) );
  OR U14700 ( .A(n12368), .B(n12369), .Z(n12364) );
  NAND U14701 ( .A(n12370), .B(n12371), .Z(n12262) );
  OR U14702 ( .A(n12372), .B(n12373), .Z(n12371) );
  OR U14703 ( .A(n12374), .B(n12375), .Z(n12370) );
  ANDN U14704 ( .B(n12376), .A(n12377), .Z(n12263) );
  IV U14705 ( .A(n12378), .Z(n12376) );
  XNOR U14706 ( .A(n12343), .B(n12342), .Z(N12869) );
  XOR U14707 ( .A(n12362), .B(n12361), .Z(n12342) );
  XNOR U14708 ( .A(n12377), .B(n12378), .Z(n12361) );
  XNOR U14709 ( .A(n12372), .B(n12373), .Z(n12378) );
  XNOR U14710 ( .A(n12374), .B(n12375), .Z(n12373) );
  XNOR U14711 ( .A(y[205]), .B(x[205]), .Z(n12375) );
  XNOR U14712 ( .A(y[206]), .B(x[206]), .Z(n12374) );
  XNOR U14713 ( .A(y[204]), .B(x[204]), .Z(n12372) );
  XNOR U14714 ( .A(n12366), .B(n12367), .Z(n12377) );
  XNOR U14715 ( .A(y[201]), .B(x[201]), .Z(n12367) );
  XNOR U14716 ( .A(n12368), .B(n12369), .Z(n12366) );
  XNOR U14717 ( .A(y[202]), .B(x[202]), .Z(n12369) );
  XNOR U14718 ( .A(y[203]), .B(x[203]), .Z(n12368) );
  XNOR U14719 ( .A(n12359), .B(n12358), .Z(n12362) );
  XNOR U14720 ( .A(n12354), .B(n12355), .Z(n12358) );
  XNOR U14721 ( .A(y[198]), .B(x[198]), .Z(n12355) );
  XNOR U14722 ( .A(n12356), .B(n12357), .Z(n12354) );
  XNOR U14723 ( .A(y[199]), .B(x[199]), .Z(n12357) );
  XNOR U14724 ( .A(y[200]), .B(x[200]), .Z(n12356) );
  XNOR U14725 ( .A(n12348), .B(n12349), .Z(n12359) );
  XNOR U14726 ( .A(y[195]), .B(x[195]), .Z(n12349) );
  XNOR U14727 ( .A(n12350), .B(n12351), .Z(n12348) );
  XNOR U14728 ( .A(y[196]), .B(x[196]), .Z(n12351) );
  XNOR U14729 ( .A(y[197]), .B(x[197]), .Z(n12350) );
  XOR U14730 ( .A(n12324), .B(n12325), .Z(n12343) );
  XNOR U14731 ( .A(n12340), .B(n12341), .Z(n12325) );
  XNOR U14732 ( .A(n12335), .B(n12336), .Z(n12341) );
  XNOR U14733 ( .A(n12337), .B(n12338), .Z(n12336) );
  XNOR U14734 ( .A(y[193]), .B(x[193]), .Z(n12338) );
  XNOR U14735 ( .A(y[194]), .B(x[194]), .Z(n12337) );
  XNOR U14736 ( .A(y[192]), .B(x[192]), .Z(n12335) );
  XNOR U14737 ( .A(n12329), .B(n12330), .Z(n12340) );
  XNOR U14738 ( .A(y[189]), .B(x[189]), .Z(n12330) );
  XNOR U14739 ( .A(n12331), .B(n12332), .Z(n12329) );
  XNOR U14740 ( .A(y[190]), .B(x[190]), .Z(n12332) );
  XNOR U14741 ( .A(y[191]), .B(x[191]), .Z(n12331) );
  XOR U14742 ( .A(n12323), .B(n12322), .Z(n12324) );
  XNOR U14743 ( .A(n12318), .B(n12319), .Z(n12322) );
  XNOR U14744 ( .A(y[186]), .B(x[186]), .Z(n12319) );
  XNOR U14745 ( .A(n12320), .B(n12321), .Z(n12318) );
  XNOR U14746 ( .A(y[187]), .B(x[187]), .Z(n12321) );
  XNOR U14747 ( .A(y[188]), .B(x[188]), .Z(n12320) );
  XNOR U14748 ( .A(n12312), .B(n12313), .Z(n12323) );
  XNOR U14749 ( .A(y[183]), .B(x[183]), .Z(n12313) );
  XNOR U14750 ( .A(n12314), .B(n12315), .Z(n12312) );
  XNOR U14751 ( .A(y[184]), .B(x[184]), .Z(n12315) );
  XNOR U14752 ( .A(y[185]), .B(x[185]), .Z(n12314) );
  NAND U14753 ( .A(n12379), .B(n12380), .Z(N12862) );
  NANDN U14754 ( .A(n12381), .B(n12382), .Z(n12380) );
  OR U14755 ( .A(n12383), .B(n12384), .Z(n12382) );
  NAND U14756 ( .A(n12383), .B(n12384), .Z(n12379) );
  XOR U14757 ( .A(n12383), .B(n12385), .Z(N12861) );
  XNOR U14758 ( .A(n12381), .B(n12384), .Z(n12385) );
  AND U14759 ( .A(n12386), .B(n12387), .Z(n12384) );
  NANDN U14760 ( .A(n12388), .B(n12389), .Z(n12387) );
  NANDN U14761 ( .A(n12390), .B(n12391), .Z(n12389) );
  NANDN U14762 ( .A(n12391), .B(n12390), .Z(n12386) );
  NAND U14763 ( .A(n12392), .B(n12393), .Z(n12381) );
  NANDN U14764 ( .A(n12394), .B(n12395), .Z(n12393) );
  OR U14765 ( .A(n12396), .B(n12397), .Z(n12395) );
  NAND U14766 ( .A(n12397), .B(n12396), .Z(n12392) );
  AND U14767 ( .A(n12398), .B(n12399), .Z(n12383) );
  NANDN U14768 ( .A(n12400), .B(n12401), .Z(n12399) );
  NANDN U14769 ( .A(n12402), .B(n12403), .Z(n12401) );
  NANDN U14770 ( .A(n12403), .B(n12402), .Z(n12398) );
  XOR U14771 ( .A(n12397), .B(n12404), .Z(N12860) );
  XOR U14772 ( .A(n12394), .B(n12396), .Z(n12404) );
  XNOR U14773 ( .A(n12390), .B(n12405), .Z(n12396) );
  XNOR U14774 ( .A(n12388), .B(n12391), .Z(n12405) );
  NAND U14775 ( .A(n12406), .B(n12407), .Z(n12391) );
  NAND U14776 ( .A(n12408), .B(n12409), .Z(n12407) );
  OR U14777 ( .A(n12410), .B(n12411), .Z(n12408) );
  NANDN U14778 ( .A(n12412), .B(n12410), .Z(n12406) );
  IV U14779 ( .A(n12411), .Z(n12412) );
  NAND U14780 ( .A(n12413), .B(n12414), .Z(n12388) );
  NAND U14781 ( .A(n12415), .B(n12416), .Z(n12414) );
  NANDN U14782 ( .A(n12417), .B(n12418), .Z(n12415) );
  NANDN U14783 ( .A(n12418), .B(n12417), .Z(n12413) );
  AND U14784 ( .A(n12419), .B(n12420), .Z(n12390) );
  NAND U14785 ( .A(n12421), .B(n12422), .Z(n12420) );
  OR U14786 ( .A(n12423), .B(n12424), .Z(n12421) );
  NANDN U14787 ( .A(n12425), .B(n12423), .Z(n12419) );
  NAND U14788 ( .A(n12426), .B(n12427), .Z(n12394) );
  NANDN U14789 ( .A(n12428), .B(n12429), .Z(n12427) );
  OR U14790 ( .A(n12430), .B(n12431), .Z(n12429) );
  NANDN U14791 ( .A(n12432), .B(n12430), .Z(n12426) );
  IV U14792 ( .A(n12431), .Z(n12432) );
  XNOR U14793 ( .A(n12402), .B(n12433), .Z(n12397) );
  XNOR U14794 ( .A(n12400), .B(n12403), .Z(n12433) );
  NAND U14795 ( .A(n12434), .B(n12435), .Z(n12403) );
  NAND U14796 ( .A(n12436), .B(n12437), .Z(n12435) );
  OR U14797 ( .A(n12438), .B(n12439), .Z(n12436) );
  NANDN U14798 ( .A(n12440), .B(n12438), .Z(n12434) );
  IV U14799 ( .A(n12439), .Z(n12440) );
  NAND U14800 ( .A(n12441), .B(n12442), .Z(n12400) );
  NAND U14801 ( .A(n12443), .B(n12444), .Z(n12442) );
  NANDN U14802 ( .A(n12445), .B(n12446), .Z(n12443) );
  NANDN U14803 ( .A(n12446), .B(n12445), .Z(n12441) );
  AND U14804 ( .A(n12447), .B(n12448), .Z(n12402) );
  NAND U14805 ( .A(n12449), .B(n12450), .Z(n12448) );
  OR U14806 ( .A(n12451), .B(n12452), .Z(n12449) );
  NANDN U14807 ( .A(n12453), .B(n12451), .Z(n12447) );
  XNOR U14808 ( .A(n12428), .B(n12454), .Z(N12859) );
  XOR U14809 ( .A(n12430), .B(n12431), .Z(n12454) );
  XNOR U14810 ( .A(n12444), .B(n12455), .Z(n12431) );
  XOR U14811 ( .A(n12445), .B(n12446), .Z(n12455) );
  XOR U14812 ( .A(n12451), .B(n12456), .Z(n12446) );
  XOR U14813 ( .A(n12450), .B(n12453), .Z(n12456) );
  IV U14814 ( .A(n12452), .Z(n12453) );
  NAND U14815 ( .A(n12457), .B(n12458), .Z(n12452) );
  OR U14816 ( .A(n12459), .B(n12460), .Z(n12458) );
  OR U14817 ( .A(n12461), .B(n12462), .Z(n12457) );
  NAND U14818 ( .A(n12463), .B(n12464), .Z(n12450) );
  OR U14819 ( .A(n12465), .B(n12466), .Z(n12464) );
  OR U14820 ( .A(n12467), .B(n12468), .Z(n12463) );
  NOR U14821 ( .A(n12469), .B(n12470), .Z(n12451) );
  ANDN U14822 ( .B(n12471), .A(n12472), .Z(n12445) );
  XNOR U14823 ( .A(n12438), .B(n12473), .Z(n12444) );
  XNOR U14824 ( .A(n12437), .B(n12439), .Z(n12473) );
  NAND U14825 ( .A(n12474), .B(n12475), .Z(n12439) );
  OR U14826 ( .A(n12476), .B(n12477), .Z(n12475) );
  OR U14827 ( .A(n12478), .B(n12479), .Z(n12474) );
  NAND U14828 ( .A(n12480), .B(n12481), .Z(n12437) );
  OR U14829 ( .A(n12482), .B(n12483), .Z(n12481) );
  OR U14830 ( .A(n12484), .B(n12485), .Z(n12480) );
  ANDN U14831 ( .B(n12486), .A(n12487), .Z(n12438) );
  IV U14832 ( .A(n12488), .Z(n12486) );
  ANDN U14833 ( .B(n12489), .A(n12490), .Z(n12430) );
  XOR U14834 ( .A(n12416), .B(n12491), .Z(n12428) );
  XOR U14835 ( .A(n12417), .B(n12418), .Z(n12491) );
  XOR U14836 ( .A(n12423), .B(n12492), .Z(n12418) );
  XOR U14837 ( .A(n12422), .B(n12425), .Z(n12492) );
  IV U14838 ( .A(n12424), .Z(n12425) );
  NAND U14839 ( .A(n12493), .B(n12494), .Z(n12424) );
  OR U14840 ( .A(n12495), .B(n12496), .Z(n12494) );
  OR U14841 ( .A(n12497), .B(n12498), .Z(n12493) );
  NAND U14842 ( .A(n12499), .B(n12500), .Z(n12422) );
  OR U14843 ( .A(n12501), .B(n12502), .Z(n12500) );
  OR U14844 ( .A(n12503), .B(n12504), .Z(n12499) );
  NOR U14845 ( .A(n12505), .B(n12506), .Z(n12423) );
  ANDN U14846 ( .B(n12507), .A(n12508), .Z(n12417) );
  IV U14847 ( .A(n12509), .Z(n12507) );
  XNOR U14848 ( .A(n12410), .B(n12510), .Z(n12416) );
  XNOR U14849 ( .A(n12409), .B(n12411), .Z(n12510) );
  NAND U14850 ( .A(n12511), .B(n12512), .Z(n12411) );
  OR U14851 ( .A(n12513), .B(n12514), .Z(n12512) );
  OR U14852 ( .A(n12515), .B(n12516), .Z(n12511) );
  NAND U14853 ( .A(n12517), .B(n12518), .Z(n12409) );
  OR U14854 ( .A(n12519), .B(n12520), .Z(n12518) );
  OR U14855 ( .A(n12521), .B(n12522), .Z(n12517) );
  ANDN U14856 ( .B(n12523), .A(n12524), .Z(n12410) );
  IV U14857 ( .A(n12525), .Z(n12523) );
  XNOR U14858 ( .A(n12490), .B(n12489), .Z(N12858) );
  XOR U14859 ( .A(n12509), .B(n12508), .Z(n12489) );
  XNOR U14860 ( .A(n12524), .B(n12525), .Z(n12508) );
  XNOR U14861 ( .A(n12519), .B(n12520), .Z(n12525) );
  XNOR U14862 ( .A(n12521), .B(n12522), .Z(n12520) );
  XNOR U14863 ( .A(y[181]), .B(x[181]), .Z(n12522) );
  XNOR U14864 ( .A(y[182]), .B(x[182]), .Z(n12521) );
  XNOR U14865 ( .A(y[180]), .B(x[180]), .Z(n12519) );
  XNOR U14866 ( .A(n12513), .B(n12514), .Z(n12524) );
  XNOR U14867 ( .A(y[177]), .B(x[177]), .Z(n12514) );
  XNOR U14868 ( .A(n12515), .B(n12516), .Z(n12513) );
  XNOR U14869 ( .A(y[178]), .B(x[178]), .Z(n12516) );
  XNOR U14870 ( .A(y[179]), .B(x[179]), .Z(n12515) );
  XNOR U14871 ( .A(n12506), .B(n12505), .Z(n12509) );
  XNOR U14872 ( .A(n12501), .B(n12502), .Z(n12505) );
  XNOR U14873 ( .A(y[174]), .B(x[174]), .Z(n12502) );
  XNOR U14874 ( .A(n12503), .B(n12504), .Z(n12501) );
  XNOR U14875 ( .A(y[175]), .B(x[175]), .Z(n12504) );
  XNOR U14876 ( .A(y[176]), .B(x[176]), .Z(n12503) );
  XNOR U14877 ( .A(n12495), .B(n12496), .Z(n12506) );
  XNOR U14878 ( .A(y[171]), .B(x[171]), .Z(n12496) );
  XNOR U14879 ( .A(n12497), .B(n12498), .Z(n12495) );
  XNOR U14880 ( .A(y[172]), .B(x[172]), .Z(n12498) );
  XNOR U14881 ( .A(y[173]), .B(x[173]), .Z(n12497) );
  XOR U14882 ( .A(n12471), .B(n12472), .Z(n12490) );
  XNOR U14883 ( .A(n12487), .B(n12488), .Z(n12472) );
  XNOR U14884 ( .A(n12482), .B(n12483), .Z(n12488) );
  XNOR U14885 ( .A(n12484), .B(n12485), .Z(n12483) );
  XNOR U14886 ( .A(y[169]), .B(x[169]), .Z(n12485) );
  XNOR U14887 ( .A(y[170]), .B(x[170]), .Z(n12484) );
  XNOR U14888 ( .A(y[168]), .B(x[168]), .Z(n12482) );
  XNOR U14889 ( .A(n12476), .B(n12477), .Z(n12487) );
  XNOR U14890 ( .A(y[165]), .B(x[165]), .Z(n12477) );
  XNOR U14891 ( .A(n12478), .B(n12479), .Z(n12476) );
  XNOR U14892 ( .A(y[166]), .B(x[166]), .Z(n12479) );
  XNOR U14893 ( .A(y[167]), .B(x[167]), .Z(n12478) );
  XOR U14894 ( .A(n12470), .B(n12469), .Z(n12471) );
  XNOR U14895 ( .A(n12465), .B(n12466), .Z(n12469) );
  XNOR U14896 ( .A(y[162]), .B(x[162]), .Z(n12466) );
  XNOR U14897 ( .A(n12467), .B(n12468), .Z(n12465) );
  XNOR U14898 ( .A(y[163]), .B(x[163]), .Z(n12468) );
  XNOR U14899 ( .A(y[164]), .B(x[164]), .Z(n12467) );
  XNOR U14900 ( .A(n12459), .B(n12460), .Z(n12470) );
  XNOR U14901 ( .A(y[159]), .B(x[159]), .Z(n12460) );
  XNOR U14902 ( .A(n12461), .B(n12462), .Z(n12459) );
  XNOR U14903 ( .A(y[160]), .B(x[160]), .Z(n12462) );
  XNOR U14904 ( .A(y[161]), .B(x[161]), .Z(n12461) );
  NAND U14905 ( .A(n12526), .B(n12527), .Z(N12851) );
  NANDN U14906 ( .A(n12528), .B(n12529), .Z(n12527) );
  OR U14907 ( .A(n12530), .B(n12531), .Z(n12529) );
  NAND U14908 ( .A(n12530), .B(n12531), .Z(n12526) );
  XOR U14909 ( .A(n12530), .B(n12532), .Z(N12850) );
  XNOR U14910 ( .A(n12528), .B(n12531), .Z(n12532) );
  AND U14911 ( .A(n12533), .B(n12534), .Z(n12531) );
  NANDN U14912 ( .A(n12535), .B(n12536), .Z(n12534) );
  NANDN U14913 ( .A(n12537), .B(n12538), .Z(n12536) );
  NANDN U14914 ( .A(n12538), .B(n12537), .Z(n12533) );
  NAND U14915 ( .A(n12539), .B(n12540), .Z(n12528) );
  NANDN U14916 ( .A(n12541), .B(n12542), .Z(n12540) );
  OR U14917 ( .A(n12543), .B(n12544), .Z(n12542) );
  NAND U14918 ( .A(n12544), .B(n12543), .Z(n12539) );
  AND U14919 ( .A(n12545), .B(n12546), .Z(n12530) );
  NANDN U14920 ( .A(n12547), .B(n12548), .Z(n12546) );
  NANDN U14921 ( .A(n12549), .B(n12550), .Z(n12548) );
  NANDN U14922 ( .A(n12550), .B(n12549), .Z(n12545) );
  XOR U14923 ( .A(n12544), .B(n12551), .Z(N12849) );
  XOR U14924 ( .A(n12541), .B(n12543), .Z(n12551) );
  XNOR U14925 ( .A(n12537), .B(n12552), .Z(n12543) );
  XNOR U14926 ( .A(n12535), .B(n12538), .Z(n12552) );
  NAND U14927 ( .A(n12553), .B(n12554), .Z(n12538) );
  NAND U14928 ( .A(n12555), .B(n12556), .Z(n12554) );
  OR U14929 ( .A(n12557), .B(n12558), .Z(n12555) );
  NANDN U14930 ( .A(n12559), .B(n12557), .Z(n12553) );
  IV U14931 ( .A(n12558), .Z(n12559) );
  NAND U14932 ( .A(n12560), .B(n12561), .Z(n12535) );
  NAND U14933 ( .A(n12562), .B(n12563), .Z(n12561) );
  NANDN U14934 ( .A(n12564), .B(n12565), .Z(n12562) );
  NANDN U14935 ( .A(n12565), .B(n12564), .Z(n12560) );
  AND U14936 ( .A(n12566), .B(n12567), .Z(n12537) );
  NAND U14937 ( .A(n12568), .B(n12569), .Z(n12567) );
  OR U14938 ( .A(n12570), .B(n12571), .Z(n12568) );
  NANDN U14939 ( .A(n12572), .B(n12570), .Z(n12566) );
  NAND U14940 ( .A(n12573), .B(n12574), .Z(n12541) );
  NANDN U14941 ( .A(n12575), .B(n12576), .Z(n12574) );
  OR U14942 ( .A(n12577), .B(n12578), .Z(n12576) );
  NANDN U14943 ( .A(n12579), .B(n12577), .Z(n12573) );
  IV U14944 ( .A(n12578), .Z(n12579) );
  XNOR U14945 ( .A(n12549), .B(n12580), .Z(n12544) );
  XNOR U14946 ( .A(n12547), .B(n12550), .Z(n12580) );
  NAND U14947 ( .A(n12581), .B(n12582), .Z(n12550) );
  NAND U14948 ( .A(n12583), .B(n12584), .Z(n12582) );
  OR U14949 ( .A(n12585), .B(n12586), .Z(n12583) );
  NANDN U14950 ( .A(n12587), .B(n12585), .Z(n12581) );
  IV U14951 ( .A(n12586), .Z(n12587) );
  NAND U14952 ( .A(n12588), .B(n12589), .Z(n12547) );
  NAND U14953 ( .A(n12590), .B(n12591), .Z(n12589) );
  NANDN U14954 ( .A(n12592), .B(n12593), .Z(n12590) );
  NANDN U14955 ( .A(n12593), .B(n12592), .Z(n12588) );
  AND U14956 ( .A(n12594), .B(n12595), .Z(n12549) );
  NAND U14957 ( .A(n12596), .B(n12597), .Z(n12595) );
  OR U14958 ( .A(n12598), .B(n12599), .Z(n12596) );
  NANDN U14959 ( .A(n12600), .B(n12598), .Z(n12594) );
  XNOR U14960 ( .A(n12575), .B(n12601), .Z(N12848) );
  XOR U14961 ( .A(n12577), .B(n12578), .Z(n12601) );
  XNOR U14962 ( .A(n12591), .B(n12602), .Z(n12578) );
  XOR U14963 ( .A(n12592), .B(n12593), .Z(n12602) );
  XOR U14964 ( .A(n12598), .B(n12603), .Z(n12593) );
  XOR U14965 ( .A(n12597), .B(n12600), .Z(n12603) );
  IV U14966 ( .A(n12599), .Z(n12600) );
  NAND U14967 ( .A(n12604), .B(n12605), .Z(n12599) );
  OR U14968 ( .A(n12606), .B(n12607), .Z(n12605) );
  OR U14969 ( .A(n12608), .B(n12609), .Z(n12604) );
  NAND U14970 ( .A(n12610), .B(n12611), .Z(n12597) );
  OR U14971 ( .A(n12612), .B(n12613), .Z(n12611) );
  OR U14972 ( .A(n12614), .B(n12615), .Z(n12610) );
  NOR U14973 ( .A(n12616), .B(n12617), .Z(n12598) );
  ANDN U14974 ( .B(n12618), .A(n12619), .Z(n12592) );
  XNOR U14975 ( .A(n12585), .B(n12620), .Z(n12591) );
  XNOR U14976 ( .A(n12584), .B(n12586), .Z(n12620) );
  NAND U14977 ( .A(n12621), .B(n12622), .Z(n12586) );
  OR U14978 ( .A(n12623), .B(n12624), .Z(n12622) );
  OR U14979 ( .A(n12625), .B(n12626), .Z(n12621) );
  NAND U14980 ( .A(n12627), .B(n12628), .Z(n12584) );
  OR U14981 ( .A(n12629), .B(n12630), .Z(n12628) );
  OR U14982 ( .A(n12631), .B(n12632), .Z(n12627) );
  ANDN U14983 ( .B(n12633), .A(n12634), .Z(n12585) );
  IV U14984 ( .A(n12635), .Z(n12633) );
  ANDN U14985 ( .B(n12636), .A(n12637), .Z(n12577) );
  XOR U14986 ( .A(n12563), .B(n12638), .Z(n12575) );
  XOR U14987 ( .A(n12564), .B(n12565), .Z(n12638) );
  XOR U14988 ( .A(n12570), .B(n12639), .Z(n12565) );
  XOR U14989 ( .A(n12569), .B(n12572), .Z(n12639) );
  IV U14990 ( .A(n12571), .Z(n12572) );
  NAND U14991 ( .A(n12640), .B(n12641), .Z(n12571) );
  OR U14992 ( .A(n12642), .B(n12643), .Z(n12641) );
  OR U14993 ( .A(n12644), .B(n12645), .Z(n12640) );
  NAND U14994 ( .A(n12646), .B(n12647), .Z(n12569) );
  OR U14995 ( .A(n12648), .B(n12649), .Z(n12647) );
  OR U14996 ( .A(n12650), .B(n12651), .Z(n12646) );
  NOR U14997 ( .A(n12652), .B(n12653), .Z(n12570) );
  ANDN U14998 ( .B(n12654), .A(n12655), .Z(n12564) );
  IV U14999 ( .A(n12656), .Z(n12654) );
  XNOR U15000 ( .A(n12557), .B(n12657), .Z(n12563) );
  XNOR U15001 ( .A(n12556), .B(n12558), .Z(n12657) );
  NAND U15002 ( .A(n12658), .B(n12659), .Z(n12558) );
  OR U15003 ( .A(n12660), .B(n12661), .Z(n12659) );
  OR U15004 ( .A(n12662), .B(n12663), .Z(n12658) );
  NAND U15005 ( .A(n12664), .B(n12665), .Z(n12556) );
  OR U15006 ( .A(n12666), .B(n12667), .Z(n12665) );
  OR U15007 ( .A(n12668), .B(n12669), .Z(n12664) );
  ANDN U15008 ( .B(n12670), .A(n12671), .Z(n12557) );
  IV U15009 ( .A(n12672), .Z(n12670) );
  XNOR U15010 ( .A(n12637), .B(n12636), .Z(N12847) );
  XOR U15011 ( .A(n12656), .B(n12655), .Z(n12636) );
  XNOR U15012 ( .A(n12671), .B(n12672), .Z(n12655) );
  XNOR U15013 ( .A(n12666), .B(n12667), .Z(n12672) );
  XNOR U15014 ( .A(n12668), .B(n12669), .Z(n12667) );
  XNOR U15015 ( .A(y[157]), .B(x[157]), .Z(n12669) );
  XNOR U15016 ( .A(y[158]), .B(x[158]), .Z(n12668) );
  XNOR U15017 ( .A(y[156]), .B(x[156]), .Z(n12666) );
  XNOR U15018 ( .A(n12660), .B(n12661), .Z(n12671) );
  XNOR U15019 ( .A(y[153]), .B(x[153]), .Z(n12661) );
  XNOR U15020 ( .A(n12662), .B(n12663), .Z(n12660) );
  XNOR U15021 ( .A(y[154]), .B(x[154]), .Z(n12663) );
  XNOR U15022 ( .A(y[155]), .B(x[155]), .Z(n12662) );
  XNOR U15023 ( .A(n12653), .B(n12652), .Z(n12656) );
  XNOR U15024 ( .A(n12648), .B(n12649), .Z(n12652) );
  XNOR U15025 ( .A(y[150]), .B(x[150]), .Z(n12649) );
  XNOR U15026 ( .A(n12650), .B(n12651), .Z(n12648) );
  XNOR U15027 ( .A(y[151]), .B(x[151]), .Z(n12651) );
  XNOR U15028 ( .A(y[152]), .B(x[152]), .Z(n12650) );
  XNOR U15029 ( .A(n12642), .B(n12643), .Z(n12653) );
  XNOR U15030 ( .A(y[147]), .B(x[147]), .Z(n12643) );
  XNOR U15031 ( .A(n12644), .B(n12645), .Z(n12642) );
  XNOR U15032 ( .A(y[148]), .B(x[148]), .Z(n12645) );
  XNOR U15033 ( .A(y[149]), .B(x[149]), .Z(n12644) );
  XOR U15034 ( .A(n12618), .B(n12619), .Z(n12637) );
  XNOR U15035 ( .A(n12634), .B(n12635), .Z(n12619) );
  XNOR U15036 ( .A(n12629), .B(n12630), .Z(n12635) );
  XNOR U15037 ( .A(n12631), .B(n12632), .Z(n12630) );
  XNOR U15038 ( .A(y[145]), .B(x[145]), .Z(n12632) );
  XNOR U15039 ( .A(y[146]), .B(x[146]), .Z(n12631) );
  XNOR U15040 ( .A(y[144]), .B(x[144]), .Z(n12629) );
  XNOR U15041 ( .A(n12623), .B(n12624), .Z(n12634) );
  XNOR U15042 ( .A(y[141]), .B(x[141]), .Z(n12624) );
  XNOR U15043 ( .A(n12625), .B(n12626), .Z(n12623) );
  XNOR U15044 ( .A(y[142]), .B(x[142]), .Z(n12626) );
  XNOR U15045 ( .A(y[143]), .B(x[143]), .Z(n12625) );
  XOR U15046 ( .A(n12617), .B(n12616), .Z(n12618) );
  XNOR U15047 ( .A(n12612), .B(n12613), .Z(n12616) );
  XNOR U15048 ( .A(y[138]), .B(x[138]), .Z(n12613) );
  XNOR U15049 ( .A(n12614), .B(n12615), .Z(n12612) );
  XNOR U15050 ( .A(y[139]), .B(x[139]), .Z(n12615) );
  XNOR U15051 ( .A(y[140]), .B(x[140]), .Z(n12614) );
  XNOR U15052 ( .A(n12606), .B(n12607), .Z(n12617) );
  XNOR U15053 ( .A(y[135]), .B(x[135]), .Z(n12607) );
  XNOR U15054 ( .A(n12608), .B(n12609), .Z(n12606) );
  XNOR U15055 ( .A(y[136]), .B(x[136]), .Z(n12609) );
  XNOR U15056 ( .A(y[137]), .B(x[137]), .Z(n12608) );
  NAND U15057 ( .A(n12673), .B(n12674), .Z(N12840) );
  NANDN U15058 ( .A(n12675), .B(n12676), .Z(n12674) );
  OR U15059 ( .A(n12677), .B(n12678), .Z(n12676) );
  NAND U15060 ( .A(n12677), .B(n12678), .Z(n12673) );
  XOR U15061 ( .A(n12677), .B(n12679), .Z(N12839) );
  XNOR U15062 ( .A(n12675), .B(n12678), .Z(n12679) );
  AND U15063 ( .A(n12680), .B(n12681), .Z(n12678) );
  NANDN U15064 ( .A(n12682), .B(n12683), .Z(n12681) );
  NANDN U15065 ( .A(n12684), .B(n12685), .Z(n12683) );
  NANDN U15066 ( .A(n12685), .B(n12684), .Z(n12680) );
  NAND U15067 ( .A(n12686), .B(n12687), .Z(n12675) );
  NANDN U15068 ( .A(n12688), .B(n12689), .Z(n12687) );
  OR U15069 ( .A(n12690), .B(n12691), .Z(n12689) );
  NAND U15070 ( .A(n12691), .B(n12690), .Z(n12686) );
  AND U15071 ( .A(n12692), .B(n12693), .Z(n12677) );
  NANDN U15072 ( .A(n12694), .B(n12695), .Z(n12693) );
  NANDN U15073 ( .A(n12696), .B(n12697), .Z(n12695) );
  NANDN U15074 ( .A(n12697), .B(n12696), .Z(n12692) );
  XOR U15075 ( .A(n12691), .B(n12698), .Z(N12838) );
  XOR U15076 ( .A(n12688), .B(n12690), .Z(n12698) );
  XNOR U15077 ( .A(n12684), .B(n12699), .Z(n12690) );
  XNOR U15078 ( .A(n12682), .B(n12685), .Z(n12699) );
  NAND U15079 ( .A(n12700), .B(n12701), .Z(n12685) );
  NAND U15080 ( .A(n12702), .B(n12703), .Z(n12701) );
  OR U15081 ( .A(n12704), .B(n12705), .Z(n12702) );
  NANDN U15082 ( .A(n12706), .B(n12704), .Z(n12700) );
  IV U15083 ( .A(n12705), .Z(n12706) );
  NAND U15084 ( .A(n12707), .B(n12708), .Z(n12682) );
  NAND U15085 ( .A(n12709), .B(n12710), .Z(n12708) );
  NANDN U15086 ( .A(n12711), .B(n12712), .Z(n12709) );
  NANDN U15087 ( .A(n12712), .B(n12711), .Z(n12707) );
  AND U15088 ( .A(n12713), .B(n12714), .Z(n12684) );
  NAND U15089 ( .A(n12715), .B(n12716), .Z(n12714) );
  OR U15090 ( .A(n12717), .B(n12718), .Z(n12715) );
  NANDN U15091 ( .A(n12719), .B(n12717), .Z(n12713) );
  NAND U15092 ( .A(n12720), .B(n12721), .Z(n12688) );
  NANDN U15093 ( .A(n12722), .B(n12723), .Z(n12721) );
  OR U15094 ( .A(n12724), .B(n12725), .Z(n12723) );
  NANDN U15095 ( .A(n12726), .B(n12724), .Z(n12720) );
  IV U15096 ( .A(n12725), .Z(n12726) );
  XNOR U15097 ( .A(n12696), .B(n12727), .Z(n12691) );
  XNOR U15098 ( .A(n12694), .B(n12697), .Z(n12727) );
  NAND U15099 ( .A(n12728), .B(n12729), .Z(n12697) );
  NAND U15100 ( .A(n12730), .B(n12731), .Z(n12729) );
  OR U15101 ( .A(n12732), .B(n12733), .Z(n12730) );
  NANDN U15102 ( .A(n12734), .B(n12732), .Z(n12728) );
  IV U15103 ( .A(n12733), .Z(n12734) );
  NAND U15104 ( .A(n12735), .B(n12736), .Z(n12694) );
  NAND U15105 ( .A(n12737), .B(n12738), .Z(n12736) );
  NANDN U15106 ( .A(n12739), .B(n12740), .Z(n12737) );
  NANDN U15107 ( .A(n12740), .B(n12739), .Z(n12735) );
  AND U15108 ( .A(n12741), .B(n12742), .Z(n12696) );
  NAND U15109 ( .A(n12743), .B(n12744), .Z(n12742) );
  OR U15110 ( .A(n12745), .B(n12746), .Z(n12743) );
  NANDN U15111 ( .A(n12747), .B(n12745), .Z(n12741) );
  XNOR U15112 ( .A(n12722), .B(n12748), .Z(N12837) );
  XOR U15113 ( .A(n12724), .B(n12725), .Z(n12748) );
  XNOR U15114 ( .A(n12738), .B(n12749), .Z(n12725) );
  XOR U15115 ( .A(n12739), .B(n12740), .Z(n12749) );
  XOR U15116 ( .A(n12745), .B(n12750), .Z(n12740) );
  XOR U15117 ( .A(n12744), .B(n12747), .Z(n12750) );
  IV U15118 ( .A(n12746), .Z(n12747) );
  NAND U15119 ( .A(n12751), .B(n12752), .Z(n12746) );
  OR U15120 ( .A(n12753), .B(n12754), .Z(n12752) );
  OR U15121 ( .A(n12755), .B(n12756), .Z(n12751) );
  NAND U15122 ( .A(n12757), .B(n12758), .Z(n12744) );
  OR U15123 ( .A(n12759), .B(n12760), .Z(n12758) );
  OR U15124 ( .A(n12761), .B(n12762), .Z(n12757) );
  NOR U15125 ( .A(n12763), .B(n12764), .Z(n12745) );
  ANDN U15126 ( .B(n12765), .A(n12766), .Z(n12739) );
  XNOR U15127 ( .A(n12732), .B(n12767), .Z(n12738) );
  XNOR U15128 ( .A(n12731), .B(n12733), .Z(n12767) );
  NAND U15129 ( .A(n12768), .B(n12769), .Z(n12733) );
  OR U15130 ( .A(n12770), .B(n12771), .Z(n12769) );
  OR U15131 ( .A(n12772), .B(n12773), .Z(n12768) );
  NAND U15132 ( .A(n12774), .B(n12775), .Z(n12731) );
  OR U15133 ( .A(n12776), .B(n12777), .Z(n12775) );
  OR U15134 ( .A(n12778), .B(n12779), .Z(n12774) );
  ANDN U15135 ( .B(n12780), .A(n12781), .Z(n12732) );
  IV U15136 ( .A(n12782), .Z(n12780) );
  ANDN U15137 ( .B(n12783), .A(n12784), .Z(n12724) );
  XOR U15138 ( .A(n12710), .B(n12785), .Z(n12722) );
  XOR U15139 ( .A(n12711), .B(n12712), .Z(n12785) );
  XOR U15140 ( .A(n12717), .B(n12786), .Z(n12712) );
  XOR U15141 ( .A(n12716), .B(n12719), .Z(n12786) );
  IV U15142 ( .A(n12718), .Z(n12719) );
  NAND U15143 ( .A(n12787), .B(n12788), .Z(n12718) );
  OR U15144 ( .A(n12789), .B(n12790), .Z(n12788) );
  OR U15145 ( .A(n12791), .B(n12792), .Z(n12787) );
  NAND U15146 ( .A(n12793), .B(n12794), .Z(n12716) );
  OR U15147 ( .A(n12795), .B(n12796), .Z(n12794) );
  OR U15148 ( .A(n12797), .B(n12798), .Z(n12793) );
  NOR U15149 ( .A(n12799), .B(n12800), .Z(n12717) );
  ANDN U15150 ( .B(n12801), .A(n12802), .Z(n12711) );
  IV U15151 ( .A(n12803), .Z(n12801) );
  XNOR U15152 ( .A(n12704), .B(n12804), .Z(n12710) );
  XNOR U15153 ( .A(n12703), .B(n12705), .Z(n12804) );
  NAND U15154 ( .A(n12805), .B(n12806), .Z(n12705) );
  OR U15155 ( .A(n12807), .B(n12808), .Z(n12806) );
  OR U15156 ( .A(n12809), .B(n12810), .Z(n12805) );
  NAND U15157 ( .A(n12811), .B(n12812), .Z(n12703) );
  OR U15158 ( .A(n12813), .B(n12814), .Z(n12812) );
  OR U15159 ( .A(n12815), .B(n12816), .Z(n12811) );
  ANDN U15160 ( .B(n12817), .A(n12818), .Z(n12704) );
  IV U15161 ( .A(n12819), .Z(n12817) );
  XNOR U15162 ( .A(n12784), .B(n12783), .Z(N12836) );
  XOR U15163 ( .A(n12803), .B(n12802), .Z(n12783) );
  XNOR U15164 ( .A(n12818), .B(n12819), .Z(n12802) );
  XNOR U15165 ( .A(n12813), .B(n12814), .Z(n12819) );
  XNOR U15166 ( .A(n12815), .B(n12816), .Z(n12814) );
  XNOR U15167 ( .A(y[133]), .B(x[133]), .Z(n12816) );
  XNOR U15168 ( .A(y[134]), .B(x[134]), .Z(n12815) );
  XNOR U15169 ( .A(y[132]), .B(x[132]), .Z(n12813) );
  XNOR U15170 ( .A(n12807), .B(n12808), .Z(n12818) );
  XNOR U15171 ( .A(y[129]), .B(x[129]), .Z(n12808) );
  XNOR U15172 ( .A(n12809), .B(n12810), .Z(n12807) );
  XNOR U15173 ( .A(y[130]), .B(x[130]), .Z(n12810) );
  XNOR U15174 ( .A(y[131]), .B(x[131]), .Z(n12809) );
  XNOR U15175 ( .A(n12800), .B(n12799), .Z(n12803) );
  XNOR U15176 ( .A(n12795), .B(n12796), .Z(n12799) );
  XNOR U15177 ( .A(y[126]), .B(x[126]), .Z(n12796) );
  XNOR U15178 ( .A(n12797), .B(n12798), .Z(n12795) );
  XNOR U15179 ( .A(y[127]), .B(x[127]), .Z(n12798) );
  XNOR U15180 ( .A(y[128]), .B(x[128]), .Z(n12797) );
  XNOR U15181 ( .A(n12789), .B(n12790), .Z(n12800) );
  XNOR U15182 ( .A(y[123]), .B(x[123]), .Z(n12790) );
  XNOR U15183 ( .A(n12791), .B(n12792), .Z(n12789) );
  XNOR U15184 ( .A(y[124]), .B(x[124]), .Z(n12792) );
  XNOR U15185 ( .A(y[125]), .B(x[125]), .Z(n12791) );
  XOR U15186 ( .A(n12765), .B(n12766), .Z(n12784) );
  XNOR U15187 ( .A(n12781), .B(n12782), .Z(n12766) );
  XNOR U15188 ( .A(n12776), .B(n12777), .Z(n12782) );
  XNOR U15189 ( .A(n12778), .B(n12779), .Z(n12777) );
  XNOR U15190 ( .A(y[121]), .B(x[121]), .Z(n12779) );
  XNOR U15191 ( .A(y[122]), .B(x[122]), .Z(n12778) );
  XNOR U15192 ( .A(y[120]), .B(x[120]), .Z(n12776) );
  XNOR U15193 ( .A(n12770), .B(n12771), .Z(n12781) );
  XNOR U15194 ( .A(y[117]), .B(x[117]), .Z(n12771) );
  XNOR U15195 ( .A(n12772), .B(n12773), .Z(n12770) );
  XNOR U15196 ( .A(y[118]), .B(x[118]), .Z(n12773) );
  XNOR U15197 ( .A(y[119]), .B(x[119]), .Z(n12772) );
  XOR U15198 ( .A(n12764), .B(n12763), .Z(n12765) );
  XNOR U15199 ( .A(n12759), .B(n12760), .Z(n12763) );
  XNOR U15200 ( .A(y[114]), .B(x[114]), .Z(n12760) );
  XNOR U15201 ( .A(n12761), .B(n12762), .Z(n12759) );
  XNOR U15202 ( .A(y[115]), .B(x[115]), .Z(n12762) );
  XNOR U15203 ( .A(y[116]), .B(x[116]), .Z(n12761) );
  XNOR U15204 ( .A(n12753), .B(n12754), .Z(n12764) );
  XNOR U15205 ( .A(y[111]), .B(x[111]), .Z(n12754) );
  XNOR U15206 ( .A(n12755), .B(n12756), .Z(n12753) );
  XNOR U15207 ( .A(y[112]), .B(x[112]), .Z(n12756) );
  XNOR U15208 ( .A(y[113]), .B(x[113]), .Z(n12755) );
  NAND U15209 ( .A(n12820), .B(n12821), .Z(N12829) );
  NANDN U15210 ( .A(n12822), .B(n12823), .Z(n12821) );
  OR U15211 ( .A(n12824), .B(n12825), .Z(n12823) );
  NAND U15212 ( .A(n12824), .B(n12825), .Z(n12820) );
  XOR U15213 ( .A(n12824), .B(n12826), .Z(N12828) );
  XNOR U15214 ( .A(n12822), .B(n12825), .Z(n12826) );
  AND U15215 ( .A(n12827), .B(n12828), .Z(n12825) );
  NANDN U15216 ( .A(n12829), .B(n12830), .Z(n12828) );
  NANDN U15217 ( .A(n12831), .B(n12832), .Z(n12830) );
  NANDN U15218 ( .A(n12832), .B(n12831), .Z(n12827) );
  NAND U15219 ( .A(n12833), .B(n12834), .Z(n12822) );
  NANDN U15220 ( .A(n12835), .B(n12836), .Z(n12834) );
  OR U15221 ( .A(n12837), .B(n12838), .Z(n12836) );
  NAND U15222 ( .A(n12838), .B(n12837), .Z(n12833) );
  AND U15223 ( .A(n12839), .B(n12840), .Z(n12824) );
  NANDN U15224 ( .A(n12841), .B(n12842), .Z(n12840) );
  NANDN U15225 ( .A(n12843), .B(n12844), .Z(n12842) );
  NANDN U15226 ( .A(n12844), .B(n12843), .Z(n12839) );
  XOR U15227 ( .A(n12838), .B(n12845), .Z(N12827) );
  XOR U15228 ( .A(n12835), .B(n12837), .Z(n12845) );
  XNOR U15229 ( .A(n12831), .B(n12846), .Z(n12837) );
  XNOR U15230 ( .A(n12829), .B(n12832), .Z(n12846) );
  NAND U15231 ( .A(n12847), .B(n12848), .Z(n12832) );
  NAND U15232 ( .A(n12849), .B(n12850), .Z(n12848) );
  OR U15233 ( .A(n12851), .B(n12852), .Z(n12849) );
  NANDN U15234 ( .A(n12853), .B(n12851), .Z(n12847) );
  IV U15235 ( .A(n12852), .Z(n12853) );
  NAND U15236 ( .A(n12854), .B(n12855), .Z(n12829) );
  NAND U15237 ( .A(n12856), .B(n12857), .Z(n12855) );
  NANDN U15238 ( .A(n12858), .B(n12859), .Z(n12856) );
  NANDN U15239 ( .A(n12859), .B(n12858), .Z(n12854) );
  AND U15240 ( .A(n12860), .B(n12861), .Z(n12831) );
  NAND U15241 ( .A(n12862), .B(n12863), .Z(n12861) );
  OR U15242 ( .A(n12864), .B(n12865), .Z(n12862) );
  NANDN U15243 ( .A(n12866), .B(n12864), .Z(n12860) );
  NAND U15244 ( .A(n12867), .B(n12868), .Z(n12835) );
  NANDN U15245 ( .A(n12869), .B(n12870), .Z(n12868) );
  OR U15246 ( .A(n12871), .B(n12872), .Z(n12870) );
  NANDN U15247 ( .A(n12873), .B(n12871), .Z(n12867) );
  IV U15248 ( .A(n12872), .Z(n12873) );
  XNOR U15249 ( .A(n12843), .B(n12874), .Z(n12838) );
  XNOR U15250 ( .A(n12841), .B(n12844), .Z(n12874) );
  NAND U15251 ( .A(n12875), .B(n12876), .Z(n12844) );
  NAND U15252 ( .A(n12877), .B(n12878), .Z(n12876) );
  OR U15253 ( .A(n12879), .B(n12880), .Z(n12877) );
  NANDN U15254 ( .A(n12881), .B(n12879), .Z(n12875) );
  IV U15255 ( .A(n12880), .Z(n12881) );
  NAND U15256 ( .A(n12882), .B(n12883), .Z(n12841) );
  NAND U15257 ( .A(n12884), .B(n12885), .Z(n12883) );
  NANDN U15258 ( .A(n12886), .B(n12887), .Z(n12884) );
  NANDN U15259 ( .A(n12887), .B(n12886), .Z(n12882) );
  AND U15260 ( .A(n12888), .B(n12889), .Z(n12843) );
  NAND U15261 ( .A(n12890), .B(n12891), .Z(n12889) );
  OR U15262 ( .A(n12892), .B(n12893), .Z(n12890) );
  NANDN U15263 ( .A(n12894), .B(n12892), .Z(n12888) );
  XNOR U15264 ( .A(n12869), .B(n12895), .Z(N12826) );
  XOR U15265 ( .A(n12871), .B(n12872), .Z(n12895) );
  XNOR U15266 ( .A(n12885), .B(n12896), .Z(n12872) );
  XOR U15267 ( .A(n12886), .B(n12887), .Z(n12896) );
  XOR U15268 ( .A(n12892), .B(n12897), .Z(n12887) );
  XOR U15269 ( .A(n12891), .B(n12894), .Z(n12897) );
  IV U15270 ( .A(n12893), .Z(n12894) );
  NAND U15271 ( .A(n12898), .B(n12899), .Z(n12893) );
  OR U15272 ( .A(n12900), .B(n12901), .Z(n12899) );
  OR U15273 ( .A(n12902), .B(n12903), .Z(n12898) );
  NAND U15274 ( .A(n12904), .B(n12905), .Z(n12891) );
  OR U15275 ( .A(n12906), .B(n12907), .Z(n12905) );
  OR U15276 ( .A(n12908), .B(n12909), .Z(n12904) );
  NOR U15277 ( .A(n12910), .B(n12911), .Z(n12892) );
  ANDN U15278 ( .B(n12912), .A(n12913), .Z(n12886) );
  XNOR U15279 ( .A(n12879), .B(n12914), .Z(n12885) );
  XNOR U15280 ( .A(n12878), .B(n12880), .Z(n12914) );
  NAND U15281 ( .A(n12915), .B(n12916), .Z(n12880) );
  OR U15282 ( .A(n12917), .B(n12918), .Z(n12916) );
  OR U15283 ( .A(n12919), .B(n12920), .Z(n12915) );
  NAND U15284 ( .A(n12921), .B(n12922), .Z(n12878) );
  OR U15285 ( .A(n12923), .B(n12924), .Z(n12922) );
  OR U15286 ( .A(n12925), .B(n12926), .Z(n12921) );
  ANDN U15287 ( .B(n12927), .A(n12928), .Z(n12879) );
  IV U15288 ( .A(n12929), .Z(n12927) );
  ANDN U15289 ( .B(n12930), .A(n12931), .Z(n12871) );
  XOR U15290 ( .A(n12857), .B(n12932), .Z(n12869) );
  XOR U15291 ( .A(n12858), .B(n12859), .Z(n12932) );
  XOR U15292 ( .A(n12864), .B(n12933), .Z(n12859) );
  XOR U15293 ( .A(n12863), .B(n12866), .Z(n12933) );
  IV U15294 ( .A(n12865), .Z(n12866) );
  NAND U15295 ( .A(n12934), .B(n12935), .Z(n12865) );
  OR U15296 ( .A(n12936), .B(n12937), .Z(n12935) );
  OR U15297 ( .A(n12938), .B(n12939), .Z(n12934) );
  NAND U15298 ( .A(n12940), .B(n12941), .Z(n12863) );
  OR U15299 ( .A(n12942), .B(n12943), .Z(n12941) );
  OR U15300 ( .A(n12944), .B(n12945), .Z(n12940) );
  NOR U15301 ( .A(n12946), .B(n12947), .Z(n12864) );
  ANDN U15302 ( .B(n12948), .A(n12949), .Z(n12858) );
  IV U15303 ( .A(n12950), .Z(n12948) );
  XNOR U15304 ( .A(n12851), .B(n12951), .Z(n12857) );
  XNOR U15305 ( .A(n12850), .B(n12852), .Z(n12951) );
  NAND U15306 ( .A(n12952), .B(n12953), .Z(n12852) );
  OR U15307 ( .A(n12954), .B(n12955), .Z(n12953) );
  OR U15308 ( .A(n12956), .B(n12957), .Z(n12952) );
  NAND U15309 ( .A(n12958), .B(n12959), .Z(n12850) );
  OR U15310 ( .A(n12960), .B(n12961), .Z(n12959) );
  OR U15311 ( .A(n12962), .B(n12963), .Z(n12958) );
  ANDN U15312 ( .B(n12964), .A(n12965), .Z(n12851) );
  IV U15313 ( .A(n12966), .Z(n12964) );
  XNOR U15314 ( .A(n12931), .B(n12930), .Z(N12825) );
  XOR U15315 ( .A(n12950), .B(n12949), .Z(n12930) );
  XNOR U15316 ( .A(n12965), .B(n12966), .Z(n12949) );
  XNOR U15317 ( .A(n12960), .B(n12961), .Z(n12966) );
  XNOR U15318 ( .A(n12962), .B(n12963), .Z(n12961) );
  XNOR U15319 ( .A(y[109]), .B(x[109]), .Z(n12963) );
  XNOR U15320 ( .A(y[110]), .B(x[110]), .Z(n12962) );
  XNOR U15321 ( .A(y[108]), .B(x[108]), .Z(n12960) );
  XNOR U15322 ( .A(n12954), .B(n12955), .Z(n12965) );
  XNOR U15323 ( .A(y[105]), .B(x[105]), .Z(n12955) );
  XNOR U15324 ( .A(n12956), .B(n12957), .Z(n12954) );
  XNOR U15325 ( .A(y[106]), .B(x[106]), .Z(n12957) );
  XNOR U15326 ( .A(y[107]), .B(x[107]), .Z(n12956) );
  XNOR U15327 ( .A(n12947), .B(n12946), .Z(n12950) );
  XNOR U15328 ( .A(n12942), .B(n12943), .Z(n12946) );
  XNOR U15329 ( .A(y[102]), .B(x[102]), .Z(n12943) );
  XNOR U15330 ( .A(n12944), .B(n12945), .Z(n12942) );
  XNOR U15331 ( .A(y[103]), .B(x[103]), .Z(n12945) );
  XNOR U15332 ( .A(y[104]), .B(x[104]), .Z(n12944) );
  XNOR U15333 ( .A(n12936), .B(n12937), .Z(n12947) );
  XNOR U15334 ( .A(y[99]), .B(x[99]), .Z(n12937) );
  XNOR U15335 ( .A(n12938), .B(n12939), .Z(n12936) );
  XNOR U15336 ( .A(y[100]), .B(x[100]), .Z(n12939) );
  XNOR U15337 ( .A(y[101]), .B(x[101]), .Z(n12938) );
  XOR U15338 ( .A(n12912), .B(n12913), .Z(n12931) );
  XNOR U15339 ( .A(n12928), .B(n12929), .Z(n12913) );
  XNOR U15340 ( .A(n12923), .B(n12924), .Z(n12929) );
  XNOR U15341 ( .A(n12925), .B(n12926), .Z(n12924) );
  XNOR U15342 ( .A(y[97]), .B(x[97]), .Z(n12926) );
  XNOR U15343 ( .A(y[98]), .B(x[98]), .Z(n12925) );
  XNOR U15344 ( .A(y[96]), .B(x[96]), .Z(n12923) );
  XNOR U15345 ( .A(n12917), .B(n12918), .Z(n12928) );
  XNOR U15346 ( .A(y[93]), .B(x[93]), .Z(n12918) );
  XNOR U15347 ( .A(n12919), .B(n12920), .Z(n12917) );
  XNOR U15348 ( .A(y[94]), .B(x[94]), .Z(n12920) );
  XNOR U15349 ( .A(y[95]), .B(x[95]), .Z(n12919) );
  XOR U15350 ( .A(n12911), .B(n12910), .Z(n12912) );
  XNOR U15351 ( .A(n12906), .B(n12907), .Z(n12910) );
  XNOR U15352 ( .A(y[90]), .B(x[90]), .Z(n12907) );
  XNOR U15353 ( .A(n12908), .B(n12909), .Z(n12906) );
  XNOR U15354 ( .A(y[91]), .B(x[91]), .Z(n12909) );
  XNOR U15355 ( .A(y[92]), .B(x[92]), .Z(n12908) );
  XNOR U15356 ( .A(n12900), .B(n12901), .Z(n12911) );
  XNOR U15357 ( .A(y[87]), .B(x[87]), .Z(n12901) );
  XNOR U15358 ( .A(n12902), .B(n12903), .Z(n12900) );
  XNOR U15359 ( .A(y[88]), .B(x[88]), .Z(n12903) );
  XNOR U15360 ( .A(y[89]), .B(x[89]), .Z(n12902) );
  NAND U15361 ( .A(n12967), .B(n12968), .Z(N12818) );
  NANDN U15362 ( .A(n12969), .B(n12970), .Z(n12968) );
  OR U15363 ( .A(n12971), .B(n12972), .Z(n12970) );
  NAND U15364 ( .A(n12971), .B(n12972), .Z(n12967) );
  XOR U15365 ( .A(n12971), .B(n12973), .Z(N12817) );
  XNOR U15366 ( .A(n12969), .B(n12972), .Z(n12973) );
  AND U15367 ( .A(n12974), .B(n12975), .Z(n12972) );
  NANDN U15368 ( .A(n12976), .B(n12977), .Z(n12975) );
  NANDN U15369 ( .A(n12978), .B(n12979), .Z(n12977) );
  NANDN U15370 ( .A(n12979), .B(n12978), .Z(n12974) );
  NAND U15371 ( .A(n12980), .B(n12981), .Z(n12969) );
  NANDN U15372 ( .A(n12982), .B(n12983), .Z(n12981) );
  OR U15373 ( .A(n12984), .B(n12985), .Z(n12983) );
  NAND U15374 ( .A(n12985), .B(n12984), .Z(n12980) );
  AND U15375 ( .A(n12986), .B(n12987), .Z(n12971) );
  NANDN U15376 ( .A(n12988), .B(n12989), .Z(n12987) );
  NANDN U15377 ( .A(n12990), .B(n12991), .Z(n12989) );
  NANDN U15378 ( .A(n12991), .B(n12990), .Z(n12986) );
  XOR U15379 ( .A(n12985), .B(n12992), .Z(N12816) );
  XOR U15380 ( .A(n12982), .B(n12984), .Z(n12992) );
  XNOR U15381 ( .A(n12978), .B(n12993), .Z(n12984) );
  XNOR U15382 ( .A(n12976), .B(n12979), .Z(n12993) );
  NAND U15383 ( .A(n12994), .B(n12995), .Z(n12979) );
  NAND U15384 ( .A(n12996), .B(n12997), .Z(n12995) );
  OR U15385 ( .A(n12998), .B(n12999), .Z(n12996) );
  NANDN U15386 ( .A(n13000), .B(n12998), .Z(n12994) );
  IV U15387 ( .A(n12999), .Z(n13000) );
  NAND U15388 ( .A(n13001), .B(n13002), .Z(n12976) );
  NAND U15389 ( .A(n13003), .B(n13004), .Z(n13002) );
  NANDN U15390 ( .A(n13005), .B(n13006), .Z(n13003) );
  NANDN U15391 ( .A(n13006), .B(n13005), .Z(n13001) );
  AND U15392 ( .A(n13007), .B(n13008), .Z(n12978) );
  NAND U15393 ( .A(n13009), .B(n13010), .Z(n13008) );
  OR U15394 ( .A(n13011), .B(n13012), .Z(n13009) );
  NANDN U15395 ( .A(n13013), .B(n13011), .Z(n13007) );
  NAND U15396 ( .A(n13014), .B(n13015), .Z(n12982) );
  NANDN U15397 ( .A(n13016), .B(n13017), .Z(n13015) );
  OR U15398 ( .A(n13018), .B(n13019), .Z(n13017) );
  NANDN U15399 ( .A(n13020), .B(n13018), .Z(n13014) );
  IV U15400 ( .A(n13019), .Z(n13020) );
  XNOR U15401 ( .A(n12990), .B(n13021), .Z(n12985) );
  XNOR U15402 ( .A(n12988), .B(n12991), .Z(n13021) );
  NAND U15403 ( .A(n13022), .B(n13023), .Z(n12991) );
  NAND U15404 ( .A(n13024), .B(n13025), .Z(n13023) );
  OR U15405 ( .A(n13026), .B(n13027), .Z(n13024) );
  NANDN U15406 ( .A(n13028), .B(n13026), .Z(n13022) );
  IV U15407 ( .A(n13027), .Z(n13028) );
  NAND U15408 ( .A(n13029), .B(n13030), .Z(n12988) );
  NAND U15409 ( .A(n13031), .B(n13032), .Z(n13030) );
  NANDN U15410 ( .A(n13033), .B(n13034), .Z(n13031) );
  NANDN U15411 ( .A(n13034), .B(n13033), .Z(n13029) );
  AND U15412 ( .A(n13035), .B(n13036), .Z(n12990) );
  NAND U15413 ( .A(n13037), .B(n13038), .Z(n13036) );
  OR U15414 ( .A(n13039), .B(n13040), .Z(n13037) );
  NANDN U15415 ( .A(n13041), .B(n13039), .Z(n13035) );
  XNOR U15416 ( .A(n13016), .B(n13042), .Z(N12815) );
  XOR U15417 ( .A(n13018), .B(n13019), .Z(n13042) );
  XNOR U15418 ( .A(n13032), .B(n13043), .Z(n13019) );
  XOR U15419 ( .A(n13033), .B(n13034), .Z(n13043) );
  XOR U15420 ( .A(n13039), .B(n13044), .Z(n13034) );
  XOR U15421 ( .A(n13038), .B(n13041), .Z(n13044) );
  IV U15422 ( .A(n13040), .Z(n13041) );
  NAND U15423 ( .A(n13045), .B(n13046), .Z(n13040) );
  OR U15424 ( .A(n13047), .B(n13048), .Z(n13046) );
  OR U15425 ( .A(n13049), .B(n13050), .Z(n13045) );
  NAND U15426 ( .A(n13051), .B(n13052), .Z(n13038) );
  OR U15427 ( .A(n13053), .B(n13054), .Z(n13052) );
  OR U15428 ( .A(n13055), .B(n13056), .Z(n13051) );
  NOR U15429 ( .A(n13057), .B(n13058), .Z(n13039) );
  ANDN U15430 ( .B(n13059), .A(n13060), .Z(n13033) );
  XNOR U15431 ( .A(n13026), .B(n13061), .Z(n13032) );
  XNOR U15432 ( .A(n13025), .B(n13027), .Z(n13061) );
  NAND U15433 ( .A(n13062), .B(n13063), .Z(n13027) );
  OR U15434 ( .A(n13064), .B(n13065), .Z(n13063) );
  OR U15435 ( .A(n13066), .B(n13067), .Z(n13062) );
  NAND U15436 ( .A(n13068), .B(n13069), .Z(n13025) );
  OR U15437 ( .A(n13070), .B(n13071), .Z(n13069) );
  OR U15438 ( .A(n13072), .B(n13073), .Z(n13068) );
  ANDN U15439 ( .B(n13074), .A(n13075), .Z(n13026) );
  IV U15440 ( .A(n13076), .Z(n13074) );
  ANDN U15441 ( .B(n13077), .A(n13078), .Z(n13018) );
  XOR U15442 ( .A(n13004), .B(n13079), .Z(n13016) );
  XOR U15443 ( .A(n13005), .B(n13006), .Z(n13079) );
  XOR U15444 ( .A(n13011), .B(n13080), .Z(n13006) );
  XOR U15445 ( .A(n13010), .B(n13013), .Z(n13080) );
  IV U15446 ( .A(n13012), .Z(n13013) );
  NAND U15447 ( .A(n13081), .B(n13082), .Z(n13012) );
  OR U15448 ( .A(n13083), .B(n13084), .Z(n13082) );
  OR U15449 ( .A(n13085), .B(n13086), .Z(n13081) );
  NAND U15450 ( .A(n13087), .B(n13088), .Z(n13010) );
  OR U15451 ( .A(n13089), .B(n13090), .Z(n13088) );
  OR U15452 ( .A(n13091), .B(n13092), .Z(n13087) );
  NOR U15453 ( .A(n13093), .B(n13094), .Z(n13011) );
  ANDN U15454 ( .B(n13095), .A(n13096), .Z(n13005) );
  IV U15455 ( .A(n13097), .Z(n13095) );
  XNOR U15456 ( .A(n12998), .B(n13098), .Z(n13004) );
  XNOR U15457 ( .A(n12997), .B(n12999), .Z(n13098) );
  NAND U15458 ( .A(n13099), .B(n13100), .Z(n12999) );
  OR U15459 ( .A(n13101), .B(n13102), .Z(n13100) );
  OR U15460 ( .A(n13103), .B(n13104), .Z(n13099) );
  NAND U15461 ( .A(n13105), .B(n13106), .Z(n12997) );
  OR U15462 ( .A(n13107), .B(n13108), .Z(n13106) );
  OR U15463 ( .A(n13109), .B(n13110), .Z(n13105) );
  ANDN U15464 ( .B(n13111), .A(n13112), .Z(n12998) );
  IV U15465 ( .A(n13113), .Z(n13111) );
  XNOR U15466 ( .A(n13078), .B(n13077), .Z(N12814) );
  XOR U15467 ( .A(n13097), .B(n13096), .Z(n13077) );
  XNOR U15468 ( .A(n13112), .B(n13113), .Z(n13096) );
  XNOR U15469 ( .A(n13107), .B(n13108), .Z(n13113) );
  XNOR U15470 ( .A(n13109), .B(n13110), .Z(n13108) );
  XNOR U15471 ( .A(y[85]), .B(x[85]), .Z(n13110) );
  XNOR U15472 ( .A(y[86]), .B(x[86]), .Z(n13109) );
  XNOR U15473 ( .A(y[84]), .B(x[84]), .Z(n13107) );
  XNOR U15474 ( .A(n13101), .B(n13102), .Z(n13112) );
  XNOR U15475 ( .A(y[81]), .B(x[81]), .Z(n13102) );
  XNOR U15476 ( .A(n13103), .B(n13104), .Z(n13101) );
  XNOR U15477 ( .A(y[82]), .B(x[82]), .Z(n13104) );
  XNOR U15478 ( .A(y[83]), .B(x[83]), .Z(n13103) );
  XNOR U15479 ( .A(n13094), .B(n13093), .Z(n13097) );
  XNOR U15480 ( .A(n13089), .B(n13090), .Z(n13093) );
  XNOR U15481 ( .A(y[78]), .B(x[78]), .Z(n13090) );
  XNOR U15482 ( .A(n13091), .B(n13092), .Z(n13089) );
  XNOR U15483 ( .A(y[79]), .B(x[79]), .Z(n13092) );
  XNOR U15484 ( .A(y[80]), .B(x[80]), .Z(n13091) );
  XNOR U15485 ( .A(n13083), .B(n13084), .Z(n13094) );
  XNOR U15486 ( .A(y[75]), .B(x[75]), .Z(n13084) );
  XNOR U15487 ( .A(n13085), .B(n13086), .Z(n13083) );
  XNOR U15488 ( .A(y[76]), .B(x[76]), .Z(n13086) );
  XNOR U15489 ( .A(y[77]), .B(x[77]), .Z(n13085) );
  XOR U15490 ( .A(n13059), .B(n13060), .Z(n13078) );
  XNOR U15491 ( .A(n13075), .B(n13076), .Z(n13060) );
  XNOR U15492 ( .A(n13070), .B(n13071), .Z(n13076) );
  XNOR U15493 ( .A(n13072), .B(n13073), .Z(n13071) );
  XNOR U15494 ( .A(y[73]), .B(x[73]), .Z(n13073) );
  XNOR U15495 ( .A(y[74]), .B(x[74]), .Z(n13072) );
  XNOR U15496 ( .A(y[72]), .B(x[72]), .Z(n13070) );
  XNOR U15497 ( .A(n13064), .B(n13065), .Z(n13075) );
  XNOR U15498 ( .A(y[69]), .B(x[69]), .Z(n13065) );
  XNOR U15499 ( .A(n13066), .B(n13067), .Z(n13064) );
  XNOR U15500 ( .A(y[70]), .B(x[70]), .Z(n13067) );
  XNOR U15501 ( .A(y[71]), .B(x[71]), .Z(n13066) );
  XOR U15502 ( .A(n13058), .B(n13057), .Z(n13059) );
  XNOR U15503 ( .A(n13053), .B(n13054), .Z(n13057) );
  XNOR U15504 ( .A(y[66]), .B(x[66]), .Z(n13054) );
  XNOR U15505 ( .A(n13055), .B(n13056), .Z(n13053) );
  XNOR U15506 ( .A(y[67]), .B(x[67]), .Z(n13056) );
  XNOR U15507 ( .A(y[68]), .B(x[68]), .Z(n13055) );
  XNOR U15508 ( .A(n13047), .B(n13048), .Z(n13058) );
  XNOR U15509 ( .A(y[63]), .B(x[63]), .Z(n13048) );
  XNOR U15510 ( .A(n13049), .B(n13050), .Z(n13047) );
  XNOR U15511 ( .A(y[64]), .B(x[64]), .Z(n13050) );
  XNOR U15512 ( .A(y[65]), .B(x[65]), .Z(n13049) );
  NAND U15513 ( .A(n13114), .B(n13115), .Z(N12807) );
  NANDN U15514 ( .A(n13116), .B(n13117), .Z(n13115) );
  OR U15515 ( .A(n13118), .B(n13119), .Z(n13117) );
  NAND U15516 ( .A(n13118), .B(n13119), .Z(n13114) );
  XOR U15517 ( .A(n13118), .B(n13120), .Z(N12806) );
  XNOR U15518 ( .A(n13116), .B(n13119), .Z(n13120) );
  AND U15519 ( .A(n13121), .B(n13122), .Z(n13119) );
  NANDN U15520 ( .A(n13123), .B(n13124), .Z(n13122) );
  NANDN U15521 ( .A(n13125), .B(n13126), .Z(n13124) );
  NANDN U15522 ( .A(n13126), .B(n13125), .Z(n13121) );
  NAND U15523 ( .A(n13127), .B(n13128), .Z(n13116) );
  NANDN U15524 ( .A(n13129), .B(n13130), .Z(n13128) );
  OR U15525 ( .A(n13131), .B(n13132), .Z(n13130) );
  NAND U15526 ( .A(n13132), .B(n13131), .Z(n13127) );
  AND U15527 ( .A(n13133), .B(n13134), .Z(n13118) );
  NANDN U15528 ( .A(n13135), .B(n13136), .Z(n13134) );
  NANDN U15529 ( .A(n13137), .B(n13138), .Z(n13136) );
  NANDN U15530 ( .A(n13138), .B(n13137), .Z(n13133) );
  XOR U15531 ( .A(n13132), .B(n13139), .Z(N12805) );
  XOR U15532 ( .A(n13129), .B(n13131), .Z(n13139) );
  XNOR U15533 ( .A(n13125), .B(n13140), .Z(n13131) );
  XNOR U15534 ( .A(n13123), .B(n13126), .Z(n13140) );
  NAND U15535 ( .A(n13141), .B(n13142), .Z(n13126) );
  NAND U15536 ( .A(n13143), .B(n13144), .Z(n13142) );
  OR U15537 ( .A(n13145), .B(n13146), .Z(n13143) );
  NANDN U15538 ( .A(n13147), .B(n13145), .Z(n13141) );
  IV U15539 ( .A(n13146), .Z(n13147) );
  NAND U15540 ( .A(n13148), .B(n13149), .Z(n13123) );
  NAND U15541 ( .A(n13150), .B(n13151), .Z(n13149) );
  NANDN U15542 ( .A(n13152), .B(n13153), .Z(n13150) );
  NANDN U15543 ( .A(n13153), .B(n13152), .Z(n13148) );
  AND U15544 ( .A(n13154), .B(n13155), .Z(n13125) );
  NAND U15545 ( .A(n13156), .B(n13157), .Z(n13155) );
  OR U15546 ( .A(n13158), .B(n13159), .Z(n13156) );
  NANDN U15547 ( .A(n13160), .B(n13158), .Z(n13154) );
  NAND U15548 ( .A(n13161), .B(n13162), .Z(n13129) );
  NANDN U15549 ( .A(n13163), .B(n13164), .Z(n13162) );
  OR U15550 ( .A(n13165), .B(n13166), .Z(n13164) );
  NANDN U15551 ( .A(n13167), .B(n13165), .Z(n13161) );
  IV U15552 ( .A(n13166), .Z(n13167) );
  XNOR U15553 ( .A(n13137), .B(n13168), .Z(n13132) );
  XNOR U15554 ( .A(n13135), .B(n13138), .Z(n13168) );
  NAND U15555 ( .A(n13169), .B(n13170), .Z(n13138) );
  NAND U15556 ( .A(n13171), .B(n13172), .Z(n13170) );
  OR U15557 ( .A(n13173), .B(n13174), .Z(n13171) );
  NANDN U15558 ( .A(n13175), .B(n13173), .Z(n13169) );
  IV U15559 ( .A(n13174), .Z(n13175) );
  NAND U15560 ( .A(n13176), .B(n13177), .Z(n13135) );
  NAND U15561 ( .A(n13178), .B(n13179), .Z(n13177) );
  NANDN U15562 ( .A(n13180), .B(n13181), .Z(n13178) );
  NANDN U15563 ( .A(n13181), .B(n13180), .Z(n13176) );
  AND U15564 ( .A(n13182), .B(n13183), .Z(n13137) );
  NAND U15565 ( .A(n13184), .B(n13185), .Z(n13183) );
  OR U15566 ( .A(n13186), .B(n13187), .Z(n13184) );
  NANDN U15567 ( .A(n13188), .B(n13186), .Z(n13182) );
  XNOR U15568 ( .A(n13163), .B(n13189), .Z(N12804) );
  XOR U15569 ( .A(n13165), .B(n13166), .Z(n13189) );
  XNOR U15570 ( .A(n13179), .B(n13190), .Z(n13166) );
  XOR U15571 ( .A(n13180), .B(n13181), .Z(n13190) );
  XOR U15572 ( .A(n13186), .B(n13191), .Z(n13181) );
  XOR U15573 ( .A(n13185), .B(n13188), .Z(n13191) );
  IV U15574 ( .A(n13187), .Z(n13188) );
  NAND U15575 ( .A(n13192), .B(n13193), .Z(n13187) );
  OR U15576 ( .A(n13194), .B(n13195), .Z(n13193) );
  OR U15577 ( .A(n13196), .B(n13197), .Z(n13192) );
  NAND U15578 ( .A(n13198), .B(n13199), .Z(n13185) );
  OR U15579 ( .A(n13200), .B(n13201), .Z(n13199) );
  OR U15580 ( .A(n13202), .B(n13203), .Z(n13198) );
  NOR U15581 ( .A(n13204), .B(n13205), .Z(n13186) );
  ANDN U15582 ( .B(n13206), .A(n13207), .Z(n13180) );
  XNOR U15583 ( .A(n13173), .B(n13208), .Z(n13179) );
  XNOR U15584 ( .A(n13172), .B(n13174), .Z(n13208) );
  NAND U15585 ( .A(n13209), .B(n13210), .Z(n13174) );
  OR U15586 ( .A(n13211), .B(n13212), .Z(n13210) );
  OR U15587 ( .A(n13213), .B(n13214), .Z(n13209) );
  NAND U15588 ( .A(n13215), .B(n13216), .Z(n13172) );
  OR U15589 ( .A(n13217), .B(n13218), .Z(n13216) );
  OR U15590 ( .A(n13219), .B(n13220), .Z(n13215) );
  ANDN U15591 ( .B(n13221), .A(n13222), .Z(n13173) );
  IV U15592 ( .A(n13223), .Z(n13221) );
  ANDN U15593 ( .B(n13224), .A(n13225), .Z(n13165) );
  XOR U15594 ( .A(n13151), .B(n13226), .Z(n13163) );
  XOR U15595 ( .A(n13152), .B(n13153), .Z(n13226) );
  XOR U15596 ( .A(n13158), .B(n13227), .Z(n13153) );
  XOR U15597 ( .A(n13157), .B(n13160), .Z(n13227) );
  IV U15598 ( .A(n13159), .Z(n13160) );
  NAND U15599 ( .A(n13228), .B(n13229), .Z(n13159) );
  OR U15600 ( .A(n13230), .B(n13231), .Z(n13229) );
  OR U15601 ( .A(n13232), .B(n13233), .Z(n13228) );
  NAND U15602 ( .A(n13234), .B(n13235), .Z(n13157) );
  OR U15603 ( .A(n13236), .B(n13237), .Z(n13235) );
  OR U15604 ( .A(n13238), .B(n13239), .Z(n13234) );
  NOR U15605 ( .A(n13240), .B(n13241), .Z(n13158) );
  ANDN U15606 ( .B(n13242), .A(n13243), .Z(n13152) );
  IV U15607 ( .A(n13244), .Z(n13242) );
  XNOR U15608 ( .A(n13145), .B(n13245), .Z(n13151) );
  XNOR U15609 ( .A(n13144), .B(n13146), .Z(n13245) );
  NAND U15610 ( .A(n13246), .B(n13247), .Z(n13146) );
  OR U15611 ( .A(n13248), .B(n13249), .Z(n13247) );
  OR U15612 ( .A(n13250), .B(n13251), .Z(n13246) );
  NAND U15613 ( .A(n13252), .B(n13253), .Z(n13144) );
  OR U15614 ( .A(n13254), .B(n13255), .Z(n13253) );
  OR U15615 ( .A(n13256), .B(n13257), .Z(n13252) );
  ANDN U15616 ( .B(n13258), .A(n13259), .Z(n13145) );
  IV U15617 ( .A(n13260), .Z(n13258) );
  XNOR U15618 ( .A(n13225), .B(n13224), .Z(N12803) );
  XOR U15619 ( .A(n13244), .B(n13243), .Z(n13224) );
  XNOR U15620 ( .A(n13259), .B(n13260), .Z(n13243) );
  XNOR U15621 ( .A(n13254), .B(n13255), .Z(n13260) );
  XNOR U15622 ( .A(n13256), .B(n13257), .Z(n13255) );
  XNOR U15623 ( .A(y[61]), .B(x[61]), .Z(n13257) );
  XNOR U15624 ( .A(y[62]), .B(x[62]), .Z(n13256) );
  XNOR U15625 ( .A(y[60]), .B(x[60]), .Z(n13254) );
  XNOR U15626 ( .A(n13248), .B(n13249), .Z(n13259) );
  XNOR U15627 ( .A(y[57]), .B(x[57]), .Z(n13249) );
  XNOR U15628 ( .A(n13250), .B(n13251), .Z(n13248) );
  XNOR U15629 ( .A(y[58]), .B(x[58]), .Z(n13251) );
  XNOR U15630 ( .A(y[59]), .B(x[59]), .Z(n13250) );
  XNOR U15631 ( .A(n13241), .B(n13240), .Z(n13244) );
  XNOR U15632 ( .A(n13236), .B(n13237), .Z(n13240) );
  XNOR U15633 ( .A(y[54]), .B(x[54]), .Z(n13237) );
  XNOR U15634 ( .A(n13238), .B(n13239), .Z(n13236) );
  XNOR U15635 ( .A(y[55]), .B(x[55]), .Z(n13239) );
  XNOR U15636 ( .A(y[56]), .B(x[56]), .Z(n13238) );
  XNOR U15637 ( .A(n13230), .B(n13231), .Z(n13241) );
  XNOR U15638 ( .A(y[51]), .B(x[51]), .Z(n13231) );
  XNOR U15639 ( .A(n13232), .B(n13233), .Z(n13230) );
  XNOR U15640 ( .A(y[52]), .B(x[52]), .Z(n13233) );
  XNOR U15641 ( .A(y[53]), .B(x[53]), .Z(n13232) );
  XOR U15642 ( .A(n13206), .B(n13207), .Z(n13225) );
  XNOR U15643 ( .A(n13222), .B(n13223), .Z(n13207) );
  XNOR U15644 ( .A(n13217), .B(n13218), .Z(n13223) );
  XNOR U15645 ( .A(n13219), .B(n13220), .Z(n13218) );
  XNOR U15646 ( .A(y[49]), .B(x[49]), .Z(n13220) );
  XNOR U15647 ( .A(y[50]), .B(x[50]), .Z(n13219) );
  XNOR U15648 ( .A(y[48]), .B(x[48]), .Z(n13217) );
  XNOR U15649 ( .A(n13211), .B(n13212), .Z(n13222) );
  XNOR U15650 ( .A(y[45]), .B(x[45]), .Z(n13212) );
  XNOR U15651 ( .A(n13213), .B(n13214), .Z(n13211) );
  XNOR U15652 ( .A(y[46]), .B(x[46]), .Z(n13214) );
  XNOR U15653 ( .A(y[47]), .B(x[47]), .Z(n13213) );
  XOR U15654 ( .A(n13205), .B(n13204), .Z(n13206) );
  XNOR U15655 ( .A(n13200), .B(n13201), .Z(n13204) );
  XNOR U15656 ( .A(y[42]), .B(x[42]), .Z(n13201) );
  XNOR U15657 ( .A(n13202), .B(n13203), .Z(n13200) );
  XNOR U15658 ( .A(y[43]), .B(x[43]), .Z(n13203) );
  XNOR U15659 ( .A(y[44]), .B(x[44]), .Z(n13202) );
  XNOR U15660 ( .A(n13194), .B(n13195), .Z(n13205) );
  XNOR U15661 ( .A(y[39]), .B(x[39]), .Z(n13195) );
  XNOR U15662 ( .A(n13196), .B(n13197), .Z(n13194) );
  XNOR U15663 ( .A(y[40]), .B(x[40]), .Z(n13197) );
  XNOR U15664 ( .A(y[41]), .B(x[41]), .Z(n13196) );
  NAND U15665 ( .A(n13261), .B(n13262), .Z(N12796) );
  NANDN U15666 ( .A(n13263), .B(n13264), .Z(n13262) );
  OR U15667 ( .A(n13265), .B(n13266), .Z(n13264) );
  NAND U15668 ( .A(n13265), .B(n13266), .Z(n13261) );
  XOR U15669 ( .A(n13265), .B(n13267), .Z(N12795) );
  XNOR U15670 ( .A(n13263), .B(n13266), .Z(n13267) );
  AND U15671 ( .A(n13268), .B(n13269), .Z(n13266) );
  NANDN U15672 ( .A(n13270), .B(n13271), .Z(n13269) );
  NANDN U15673 ( .A(n13272), .B(n13273), .Z(n13271) );
  NANDN U15674 ( .A(n13273), .B(n13272), .Z(n13268) );
  NAND U15675 ( .A(n13274), .B(n13275), .Z(n13263) );
  NANDN U15676 ( .A(n13276), .B(n13277), .Z(n13275) );
  OR U15677 ( .A(n13278), .B(n13279), .Z(n13277) );
  NAND U15678 ( .A(n13279), .B(n13278), .Z(n13274) );
  AND U15679 ( .A(n13280), .B(n13281), .Z(n13265) );
  NANDN U15680 ( .A(n13282), .B(n13283), .Z(n13281) );
  NANDN U15681 ( .A(n13284), .B(n13285), .Z(n13283) );
  NANDN U15682 ( .A(n13285), .B(n13284), .Z(n13280) );
  XOR U15683 ( .A(n13279), .B(n13286), .Z(N12794) );
  XOR U15684 ( .A(n13276), .B(n13278), .Z(n13286) );
  XNOR U15685 ( .A(n13272), .B(n13287), .Z(n13278) );
  XNOR U15686 ( .A(n13270), .B(n13273), .Z(n13287) );
  NAND U15687 ( .A(n13288), .B(n13289), .Z(n13273) );
  NAND U15688 ( .A(n13290), .B(n13291), .Z(n13289) );
  OR U15689 ( .A(n13292), .B(n13293), .Z(n13290) );
  NANDN U15690 ( .A(n13294), .B(n13292), .Z(n13288) );
  IV U15691 ( .A(n13293), .Z(n13294) );
  NAND U15692 ( .A(n13295), .B(n13296), .Z(n13270) );
  NAND U15693 ( .A(n13297), .B(n13298), .Z(n13296) );
  NANDN U15694 ( .A(n13299), .B(n13300), .Z(n13297) );
  NANDN U15695 ( .A(n13300), .B(n13299), .Z(n13295) );
  AND U15696 ( .A(n13301), .B(n13302), .Z(n13272) );
  NAND U15697 ( .A(n13303), .B(n13304), .Z(n13302) );
  OR U15698 ( .A(n13305), .B(n13306), .Z(n13303) );
  NANDN U15699 ( .A(n13307), .B(n13305), .Z(n13301) );
  NAND U15700 ( .A(n13308), .B(n13309), .Z(n13276) );
  NANDN U15701 ( .A(n13310), .B(n13311), .Z(n13309) );
  OR U15702 ( .A(n13312), .B(n13313), .Z(n13311) );
  NANDN U15703 ( .A(n13314), .B(n13312), .Z(n13308) );
  IV U15704 ( .A(n13313), .Z(n13314) );
  XNOR U15705 ( .A(n13284), .B(n13315), .Z(n13279) );
  XNOR U15706 ( .A(n13282), .B(n13285), .Z(n13315) );
  NAND U15707 ( .A(n13316), .B(n13317), .Z(n13285) );
  NAND U15708 ( .A(n13318), .B(n13319), .Z(n13317) );
  OR U15709 ( .A(n13320), .B(n13321), .Z(n13318) );
  NANDN U15710 ( .A(n13322), .B(n13320), .Z(n13316) );
  IV U15711 ( .A(n13321), .Z(n13322) );
  NAND U15712 ( .A(n13323), .B(n13324), .Z(n13282) );
  NAND U15713 ( .A(n13325), .B(n13326), .Z(n13324) );
  NANDN U15714 ( .A(n13327), .B(n13328), .Z(n13325) );
  NANDN U15715 ( .A(n13328), .B(n13327), .Z(n13323) );
  AND U15716 ( .A(n13329), .B(n13330), .Z(n13284) );
  NAND U15717 ( .A(n13331), .B(n13332), .Z(n13330) );
  OR U15718 ( .A(n13333), .B(n13334), .Z(n13331) );
  NANDN U15719 ( .A(n13335), .B(n13333), .Z(n13329) );
  XNOR U15720 ( .A(n13310), .B(n13336), .Z(N12793) );
  XOR U15721 ( .A(n13312), .B(n13313), .Z(n13336) );
  XNOR U15722 ( .A(n13326), .B(n13337), .Z(n13313) );
  XOR U15723 ( .A(n13327), .B(n13328), .Z(n13337) );
  XOR U15724 ( .A(n13333), .B(n13338), .Z(n13328) );
  XOR U15725 ( .A(n13332), .B(n13335), .Z(n13338) );
  IV U15726 ( .A(n13334), .Z(n13335) );
  NAND U15727 ( .A(n13339), .B(n13340), .Z(n13334) );
  OR U15728 ( .A(n13341), .B(n13342), .Z(n13340) );
  OR U15729 ( .A(n13343), .B(n13344), .Z(n13339) );
  NAND U15730 ( .A(n13345), .B(n13346), .Z(n13332) );
  OR U15731 ( .A(n13347), .B(n13348), .Z(n13346) );
  OR U15732 ( .A(n13349), .B(n13350), .Z(n13345) );
  NOR U15733 ( .A(n13351), .B(n13352), .Z(n13333) );
  ANDN U15734 ( .B(n13353), .A(n13354), .Z(n13327) );
  XNOR U15735 ( .A(n13320), .B(n13355), .Z(n13326) );
  XNOR U15736 ( .A(n13319), .B(n13321), .Z(n13355) );
  NAND U15737 ( .A(n13356), .B(n13357), .Z(n13321) );
  OR U15738 ( .A(n13358), .B(n13359), .Z(n13357) );
  OR U15739 ( .A(n13360), .B(n13361), .Z(n13356) );
  NAND U15740 ( .A(n13362), .B(n13363), .Z(n13319) );
  OR U15741 ( .A(n13364), .B(n13365), .Z(n13363) );
  OR U15742 ( .A(n13366), .B(n13367), .Z(n13362) );
  ANDN U15743 ( .B(n13368), .A(n13369), .Z(n13320) );
  IV U15744 ( .A(n13370), .Z(n13368) );
  ANDN U15745 ( .B(n13371), .A(n13372), .Z(n13312) );
  XOR U15746 ( .A(n13298), .B(n13373), .Z(n13310) );
  XOR U15747 ( .A(n13299), .B(n13300), .Z(n13373) );
  XOR U15748 ( .A(n13305), .B(n13374), .Z(n13300) );
  XOR U15749 ( .A(n13304), .B(n13307), .Z(n13374) );
  IV U15750 ( .A(n13306), .Z(n13307) );
  NAND U15751 ( .A(n13375), .B(n13376), .Z(n13306) );
  OR U15752 ( .A(n13377), .B(n13378), .Z(n13376) );
  OR U15753 ( .A(n13379), .B(n13380), .Z(n13375) );
  NAND U15754 ( .A(n13381), .B(n13382), .Z(n13304) );
  OR U15755 ( .A(n13383), .B(n13384), .Z(n13382) );
  OR U15756 ( .A(n13385), .B(n13386), .Z(n13381) );
  NOR U15757 ( .A(n13387), .B(n13388), .Z(n13305) );
  ANDN U15758 ( .B(n13389), .A(n13390), .Z(n13299) );
  IV U15759 ( .A(n13391), .Z(n13389) );
  XNOR U15760 ( .A(n13292), .B(n13392), .Z(n13298) );
  XNOR U15761 ( .A(n13291), .B(n13293), .Z(n13392) );
  NAND U15762 ( .A(n13393), .B(n13394), .Z(n13293) );
  OR U15763 ( .A(n13395), .B(n13396), .Z(n13394) );
  OR U15764 ( .A(n13397), .B(n13398), .Z(n13393) );
  NAND U15765 ( .A(n13399), .B(n13400), .Z(n13291) );
  OR U15766 ( .A(n13401), .B(n13402), .Z(n13400) );
  OR U15767 ( .A(n13403), .B(n13404), .Z(n13399) );
  ANDN U15768 ( .B(n13405), .A(n13406), .Z(n13292) );
  IV U15769 ( .A(n13407), .Z(n13405) );
  XNOR U15770 ( .A(n13372), .B(n13371), .Z(N12792) );
  XOR U15771 ( .A(n13391), .B(n13390), .Z(n13371) );
  XNOR U15772 ( .A(n13406), .B(n13407), .Z(n13390) );
  XNOR U15773 ( .A(n13401), .B(n13402), .Z(n13407) );
  XNOR U15774 ( .A(n13403), .B(n13404), .Z(n13402) );
  XNOR U15775 ( .A(y[37]), .B(x[37]), .Z(n13404) );
  XNOR U15776 ( .A(y[38]), .B(x[38]), .Z(n13403) );
  XNOR U15777 ( .A(y[36]), .B(x[36]), .Z(n13401) );
  XNOR U15778 ( .A(n13395), .B(n13396), .Z(n13406) );
  XNOR U15779 ( .A(y[33]), .B(x[33]), .Z(n13396) );
  XNOR U15780 ( .A(n13397), .B(n13398), .Z(n13395) );
  XNOR U15781 ( .A(y[34]), .B(x[34]), .Z(n13398) );
  XNOR U15782 ( .A(y[35]), .B(x[35]), .Z(n13397) );
  XNOR U15783 ( .A(n13388), .B(n13387), .Z(n13391) );
  XNOR U15784 ( .A(n13383), .B(n13384), .Z(n13387) );
  XNOR U15785 ( .A(y[30]), .B(x[30]), .Z(n13384) );
  XNOR U15786 ( .A(n13385), .B(n13386), .Z(n13383) );
  XNOR U15787 ( .A(y[31]), .B(x[31]), .Z(n13386) );
  XNOR U15788 ( .A(y[32]), .B(x[32]), .Z(n13385) );
  XNOR U15789 ( .A(n13377), .B(n13378), .Z(n13388) );
  XNOR U15790 ( .A(y[27]), .B(x[27]), .Z(n13378) );
  XNOR U15791 ( .A(n13379), .B(n13380), .Z(n13377) );
  XNOR U15792 ( .A(y[28]), .B(x[28]), .Z(n13380) );
  XNOR U15793 ( .A(y[29]), .B(x[29]), .Z(n13379) );
  XOR U15794 ( .A(n13353), .B(n13354), .Z(n13372) );
  XNOR U15795 ( .A(n13369), .B(n13370), .Z(n13354) );
  XNOR U15796 ( .A(n13364), .B(n13365), .Z(n13370) );
  XNOR U15797 ( .A(n13366), .B(n13367), .Z(n13365) );
  XNOR U15798 ( .A(y[25]), .B(x[25]), .Z(n13367) );
  XNOR U15799 ( .A(y[26]), .B(x[26]), .Z(n13366) );
  XNOR U15800 ( .A(y[24]), .B(x[24]), .Z(n13364) );
  XNOR U15801 ( .A(n13358), .B(n13359), .Z(n13369) );
  XNOR U15802 ( .A(y[21]), .B(x[21]), .Z(n13359) );
  XNOR U15803 ( .A(n13360), .B(n13361), .Z(n13358) );
  XNOR U15804 ( .A(y[22]), .B(x[22]), .Z(n13361) );
  XNOR U15805 ( .A(y[23]), .B(x[23]), .Z(n13360) );
  XOR U15806 ( .A(n13352), .B(n13351), .Z(n13353) );
  XNOR U15807 ( .A(n13347), .B(n13348), .Z(n13351) );
  XNOR U15808 ( .A(y[18]), .B(x[18]), .Z(n13348) );
  XNOR U15809 ( .A(n13349), .B(n13350), .Z(n13347) );
  XNOR U15810 ( .A(y[19]), .B(x[19]), .Z(n13350) );
  XNOR U15811 ( .A(y[20]), .B(x[20]), .Z(n13349) );
  XNOR U15812 ( .A(n13341), .B(n13342), .Z(n13352) );
  XNOR U15813 ( .A(y[15]), .B(x[15]), .Z(n13342) );
  XNOR U15814 ( .A(n13343), .B(n13344), .Z(n13341) );
  XNOR U15815 ( .A(y[16]), .B(x[16]), .Z(n13344) );
  XNOR U15816 ( .A(y[17]), .B(x[17]), .Z(n13343) );
  NAND U15817 ( .A(n13408), .B(n13409), .Z(N12785) );
  OR U15818 ( .A(n13410), .B(n13411), .Z(n13409) );
  OR U15819 ( .A(n13411), .B(n13412), .Z(n13408) );
  XNOR U15820 ( .A(n13412), .B(n13413), .Z(N12784) );
  XOR U15821 ( .A(n13410), .B(n13411), .Z(n13413) );
  NAND U15822 ( .A(n13414), .B(n13415), .Z(n13411) );
  NANDN U15823 ( .A(n13416), .B(n13417), .Z(n13415) );
  NANDN U15824 ( .A(n13418), .B(n13419), .Z(n13417) );
  NANDN U15825 ( .A(n13419), .B(n13418), .Z(n13414) );
  NAND U15826 ( .A(n13420), .B(n13421), .Z(n13410) );
  NANDN U15827 ( .A(n13422), .B(n13423), .Z(n13421) );
  OR U15828 ( .A(n13424), .B(n13425), .Z(n13423) );
  NANDN U15829 ( .A(n13426), .B(n13424), .Z(n13420) );
  IV U15830 ( .A(n13425), .Z(n13426) );
  NANDN U15831 ( .A(n13427), .B(n13428), .Z(n13412) );
  XOR U15832 ( .A(n13425), .B(n13429), .Z(N12783) );
  XOR U15833 ( .A(n13422), .B(n13424), .Z(n13429) );
  XNOR U15834 ( .A(n13418), .B(n13430), .Z(n13424) );
  XNOR U15835 ( .A(n13416), .B(n13419), .Z(n13430) );
  NAND U15836 ( .A(n13431), .B(n13432), .Z(n13419) );
  NAND U15837 ( .A(n13433), .B(n13434), .Z(n13432) );
  OR U15838 ( .A(n13435), .B(n13436), .Z(n13433) );
  NANDN U15839 ( .A(n13437), .B(n13435), .Z(n13431) );
  IV U15840 ( .A(n13436), .Z(n13437) );
  NAND U15841 ( .A(n13438), .B(n13439), .Z(n13416) );
  NAND U15842 ( .A(n13440), .B(n13441), .Z(n13439) );
  NANDN U15843 ( .A(n13442), .B(n13443), .Z(n13440) );
  NANDN U15844 ( .A(n13443), .B(n13442), .Z(n13438) );
  AND U15845 ( .A(n13444), .B(n13445), .Z(n13418) );
  NAND U15846 ( .A(n13446), .B(n13447), .Z(n13445) );
  NANDN U15847 ( .A(n13448), .B(n13449), .Z(n13444) );
  NAND U15848 ( .A(n13450), .B(n13451), .Z(n13422) );
  NANDN U15849 ( .A(n13452), .B(n13453), .Z(n13451) );
  OR U15850 ( .A(n13454), .B(n13455), .Z(n13453) );
  NAND U15851 ( .A(n13455), .B(n13454), .Z(n13450) );
  XOR U15852 ( .A(n13428), .B(n13427), .Z(n13425) );
  NANDN U15853 ( .A(n13456), .B(n13457), .Z(n13427) );
  NAND U15854 ( .A(n13458), .B(n13459), .Z(n13428) );
  NAND U15855 ( .A(n13460), .B(n13461), .Z(n13459) );
  NAND U15856 ( .A(n13462), .B(n13463), .Z(n13460) );
  OR U15857 ( .A(n13462), .B(n13463), .Z(n13458) );
  XNOR U15858 ( .A(n13452), .B(n13464), .Z(N12782) );
  XOR U15859 ( .A(n13454), .B(n13455), .Z(n13464) );
  XOR U15860 ( .A(n13461), .B(n13465), .Z(n13455) );
  XOR U15861 ( .A(n13463), .B(n13462), .Z(n13465) );
  NANDN U15862 ( .A(n13466), .B(n13467), .Z(n13462) );
  AND U15863 ( .A(n13468), .B(n13469), .Z(n13463) );
  OR U15864 ( .A(n13470), .B(n13471), .Z(n13469) );
  OR U15865 ( .A(n13472), .B(n13473), .Z(n13468) );
  XNOR U15866 ( .A(n13457), .B(n13456), .Z(n13461) );
  AND U15867 ( .A(n13474), .B(n13475), .Z(n13456) );
  OR U15868 ( .A(n13476), .B(n13477), .Z(n13475) );
  OR U15869 ( .A(n13478), .B(n13479), .Z(n13474) );
  NAND U15870 ( .A(n13480), .B(n13481), .Z(n13457) );
  OR U15871 ( .A(n13482), .B(n13483), .Z(n13480) );
  IV U15872 ( .A(n13484), .Z(n13483) );
  ANDN U15873 ( .B(n13485), .A(n13486), .Z(n13454) );
  XOR U15874 ( .A(n13441), .B(n13487), .Z(n13452) );
  XOR U15875 ( .A(n13442), .B(n13443), .Z(n13487) );
  XNOR U15876 ( .A(n13446), .B(n13447), .Z(n13443) );
  XNOR U15877 ( .A(n13449), .B(n13448), .Z(n13447) );
  AND U15878 ( .A(n13488), .B(n13489), .Z(n13448) );
  NANDN U15879 ( .A(n13490), .B(n13491), .Z(n13489) );
  OR U15880 ( .A(n13492), .B(n13493), .Z(n13488) );
  IV U15881 ( .A(n13494), .Z(n13493) );
  NAND U15882 ( .A(n13495), .B(n13496), .Z(n13449) );
  NANDN U15883 ( .A(n13497), .B(n13498), .Z(n13496) );
  OR U15884 ( .A(n13499), .B(n13500), .Z(n13495) );
  IV U15885 ( .A(n13501), .Z(n13500) );
  ANDN U15886 ( .B(n13502), .A(n13503), .Z(n13446) );
  NOR U15887 ( .A(n13504), .B(n13505), .Z(n13442) );
  XNOR U15888 ( .A(n13435), .B(n13506), .Z(n13441) );
  XNOR U15889 ( .A(n13434), .B(n13436), .Z(n13506) );
  NAND U15890 ( .A(n13507), .B(n13508), .Z(n13436) );
  OR U15891 ( .A(n13509), .B(n13510), .Z(n13508) );
  OR U15892 ( .A(n13511), .B(n13512), .Z(n13507) );
  NAND U15893 ( .A(n13513), .B(n13514), .Z(n13434) );
  OR U15894 ( .A(n13515), .B(n13516), .Z(n13514) );
  OR U15895 ( .A(n13517), .B(n13518), .Z(n13513) );
  ANDN U15896 ( .B(n13519), .A(n13520), .Z(n13435) );
  IV U15897 ( .A(n13521), .Z(n13519) );
  XNOR U15898 ( .A(n13486), .B(n13485), .Z(N12781) );
  XOR U15899 ( .A(n13505), .B(n13504), .Z(n13485) );
  XNOR U15900 ( .A(n13520), .B(n13521), .Z(n13504) );
  XNOR U15901 ( .A(n13515), .B(n13516), .Z(n13521) );
  XNOR U15902 ( .A(n13517), .B(n13518), .Z(n13516) );
  XNOR U15903 ( .A(y[13]), .B(x[13]), .Z(n13518) );
  XNOR U15904 ( .A(y[14]), .B(x[14]), .Z(n13517) );
  XNOR U15905 ( .A(y[12]), .B(x[12]), .Z(n13515) );
  XNOR U15906 ( .A(n13509), .B(n13510), .Z(n13520) );
  XNOR U15907 ( .A(y[9]), .B(x[9]), .Z(n13510) );
  XNOR U15908 ( .A(n13511), .B(n13512), .Z(n13509) );
  XNOR U15909 ( .A(y[10]), .B(x[10]), .Z(n13512) );
  XNOR U15910 ( .A(y[11]), .B(x[11]), .Z(n13511) );
  XOR U15911 ( .A(n13502), .B(n13503), .Z(n13505) );
  XOR U15912 ( .A(n13490), .B(n13491), .Z(n13503) );
  XNOR U15913 ( .A(n13492), .B(n13494), .Z(n13491) );
  XOR U15914 ( .A(y[4]), .B(x[4]), .Z(n13494) );
  XNOR U15915 ( .A(y[5]), .B(x[5]), .Z(n13492) );
  XNOR U15916 ( .A(y[3]), .B(x[3]), .Z(n13490) );
  XNOR U15917 ( .A(n13497), .B(n13498), .Z(n13502) );
  XNOR U15918 ( .A(n13499), .B(n13501), .Z(n13498) );
  XOR U15919 ( .A(y[7]), .B(x[7]), .Z(n13501) );
  XNOR U15920 ( .A(y[8]), .B(x[8]), .Z(n13499) );
  XNOR U15921 ( .A(y[6]), .B(x[6]), .Z(n13497) );
  XOR U15922 ( .A(n13466), .B(n13467), .Z(n13486) );
  XNOR U15923 ( .A(n13482), .B(n13484), .Z(n13467) );
  XOR U15924 ( .A(y[1998]), .B(x[1998]), .Z(n13484) );
  NAND U15925 ( .A(n13522), .B(n13481), .Z(n13482) );
  OR U15926 ( .A(n13523), .B(n13524), .Z(n13481) );
  NAND U15927 ( .A(n13524), .B(n13523), .Z(n13522) );
  XNOR U15928 ( .A(y[1999]), .B(x[1999]), .Z(n13523) );
  XOR U15929 ( .A(n13525), .B(n13476), .Z(n13524) );
  XNOR U15930 ( .A(y[0]), .B(x[0]), .Z(n13476) );
  IV U15931 ( .A(n13477), .Z(n13525) );
  XNOR U15932 ( .A(n13479), .B(n13478), .Z(n13477) );
  XNOR U15933 ( .A(y[1]), .B(x[1]), .Z(n13478) );
  XNOR U15934 ( .A(y[2]), .B(x[2]), .Z(n13479) );
  XNOR U15935 ( .A(n13470), .B(n13471), .Z(n13466) );
  XNOR U15936 ( .A(y[1995]), .B(x[1995]), .Z(n13471) );
  XNOR U15937 ( .A(n13472), .B(n13473), .Z(n13470) );
  XNOR U15938 ( .A(y[1996]), .B(x[1996]), .Z(n13473) );
  XNOR U15939 ( .A(y[1997]), .B(x[1997]), .Z(n13472) );
  NAND U15940 ( .A(n13526), .B(n13527), .Z(N12773) );
  NAND U15941 ( .A(n13528), .B(n13529), .Z(n13527) );
  OR U15942 ( .A(n13530), .B(n13531), .Z(n13528) );
  NANDN U15943 ( .A(n13532), .B(n13530), .Z(n13526) );
  XNOR U15944 ( .A(n13530), .B(n13533), .Z(N12772) );
  XOR U15945 ( .A(n13529), .B(n13532), .Z(n13533) );
  IV U15946 ( .A(n13531), .Z(n13532) );
  NAND U15947 ( .A(n13534), .B(n13535), .Z(n13531) );
  NAND U15948 ( .A(n13536), .B(n13537), .Z(n13535) );
  OR U15949 ( .A(n13538), .B(n13539), .Z(n13536) );
  NANDN U15950 ( .A(n13540), .B(n13538), .Z(n13534) );
  IV U15951 ( .A(n13539), .Z(n13540) );
  NAND U15952 ( .A(n13541), .B(n13542), .Z(n13529) );
  NAND U15953 ( .A(n13543), .B(n13544), .Z(n13542) );
  OR U15954 ( .A(n13545), .B(n13546), .Z(n13543) );
  NAND U15955 ( .A(n13546), .B(n13545), .Z(n13541) );
  NAND U15956 ( .A(n13547), .B(n13548), .Z(n13530) );
  NAND U15957 ( .A(n13549), .B(n13550), .Z(n13548) );
  OR U15958 ( .A(n13551), .B(n13552), .Z(n13549) );
  NANDN U15959 ( .A(n13553), .B(n13551), .Z(n13547) );
  XOR U15960 ( .A(n13544), .B(n13554), .Z(N12771) );
  XOR U15961 ( .A(n13545), .B(n13546), .Z(n13554) );
  XNOR U15962 ( .A(n13551), .B(n13555), .Z(n13546) );
  XOR U15963 ( .A(n13550), .B(n13553), .Z(n13555) );
  IV U15964 ( .A(n13552), .Z(n13553) );
  NAND U15965 ( .A(n13556), .B(n13557), .Z(n13552) );
  OR U15966 ( .A(n13558), .B(n13559), .Z(n13557) );
  OR U15967 ( .A(n13560), .B(n13561), .Z(n13556) );
  NAND U15968 ( .A(n13562), .B(n13563), .Z(n13550) );
  OR U15969 ( .A(n13564), .B(n13565), .Z(n13563) );
  OR U15970 ( .A(n13566), .B(n13567), .Z(n13562) );
  NOR U15971 ( .A(n13568), .B(n13569), .Z(n13551) );
  ANDN U15972 ( .B(n13570), .A(n13571), .Z(n13545) );
  XNOR U15973 ( .A(n13538), .B(n13572), .Z(n13544) );
  XNOR U15974 ( .A(n13537), .B(n13539), .Z(n13572) );
  NAND U15975 ( .A(n13573), .B(n13574), .Z(n13539) );
  OR U15976 ( .A(n13575), .B(n13576), .Z(n13574) );
  IV U15977 ( .A(n13577), .Z(n13576) );
  OR U15978 ( .A(n13578), .B(n13579), .Z(n13573) );
  NAND U15979 ( .A(n13580), .B(n13581), .Z(n13537) );
  OR U15980 ( .A(n13582), .B(n13583), .Z(n13581) );
  OR U15981 ( .A(n13584), .B(n13585), .Z(n13580) );
  AND U15982 ( .A(n13586), .B(n13587), .Z(n13538) );
  IV U15983 ( .A(n13588), .Z(n13587) );
  XNOR U15984 ( .A(n13571), .B(n13570), .Z(N12770) );
  XNOR U15985 ( .A(n13588), .B(n13586), .Z(n13570) );
  XOR U15986 ( .A(n13582), .B(n13583), .Z(n13586) );
  XNOR U15987 ( .A(n13584), .B(n13585), .Z(n13583) );
  XNOR U15988 ( .A(y[1993]), .B(x[1993]), .Z(n13585) );
  XNOR U15989 ( .A(y[1994]), .B(x[1994]), .Z(n13584) );
  XNOR U15990 ( .A(y[1992]), .B(x[1992]), .Z(n13582) );
  XOR U15991 ( .A(n13575), .B(n13577), .Z(n13588) );
  XOR U15992 ( .A(n13578), .B(n13579), .Z(n13577) );
  XNOR U15993 ( .A(y[1990]), .B(x[1990]), .Z(n13579) );
  XNOR U15994 ( .A(y[1991]), .B(x[1991]), .Z(n13578) );
  XNOR U15995 ( .A(y[1989]), .B(x[1989]), .Z(n13575) );
  XNOR U15996 ( .A(n13569), .B(n13568), .Z(n13571) );
  XNOR U15997 ( .A(n13564), .B(n13565), .Z(n13568) );
  XNOR U15998 ( .A(y[1986]), .B(x[1986]), .Z(n13565) );
  XNOR U15999 ( .A(n13566), .B(n13567), .Z(n13564) );
  XNOR U16000 ( .A(y[1987]), .B(x[1987]), .Z(n13567) );
  XNOR U16001 ( .A(y[1988]), .B(x[1988]), .Z(n13566) );
  XNOR U16002 ( .A(n13558), .B(n13559), .Z(n13569) );
  XNOR U16003 ( .A(y[1983]), .B(x[1983]), .Z(n13559) );
  XNOR U16004 ( .A(n13560), .B(n13561), .Z(n13558) );
  XNOR U16005 ( .A(y[1984]), .B(x[1984]), .Z(n13561) );
  XNOR U16006 ( .A(y[1985]), .B(x[1985]), .Z(n13560) );
endmodule

