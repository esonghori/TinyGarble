
module sum_N16384_CC64 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U5 ( .B(n4), .A(n5), .Z(n2) );
  XOR U6 ( .A(b[255]), .B(n3), .Z(n4) );
  XNOR U7 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U8 ( .A(b[99]), .B(n7), .Z(c[99]) );
  XNOR U9 ( .A(b[98]), .B(n8), .Z(c[98]) );
  XNOR U10 ( .A(b[97]), .B(n9), .Z(c[97]) );
  XNOR U11 ( .A(b[96]), .B(n10), .Z(c[96]) );
  XNOR U12 ( .A(b[95]), .B(n11), .Z(c[95]) );
  XNOR U13 ( .A(b[94]), .B(n12), .Z(c[94]) );
  XNOR U14 ( .A(b[93]), .B(n13), .Z(c[93]) );
  XNOR U15 ( .A(b[92]), .B(n14), .Z(c[92]) );
  XNOR U16 ( .A(b[91]), .B(n15), .Z(c[91]) );
  XNOR U17 ( .A(b[90]), .B(n16), .Z(c[90]) );
  XNOR U18 ( .A(b[8]), .B(n17), .Z(c[8]) );
  XNOR U19 ( .A(b[89]), .B(n18), .Z(c[89]) );
  XNOR U20 ( .A(b[88]), .B(n19), .Z(c[88]) );
  XNOR U21 ( .A(b[87]), .B(n20), .Z(c[87]) );
  XNOR U22 ( .A(b[86]), .B(n21), .Z(c[86]) );
  XNOR U23 ( .A(b[85]), .B(n22), .Z(c[85]) );
  XNOR U24 ( .A(b[84]), .B(n23), .Z(c[84]) );
  XNOR U25 ( .A(b[83]), .B(n24), .Z(c[83]) );
  XNOR U26 ( .A(b[82]), .B(n25), .Z(c[82]) );
  XNOR U27 ( .A(b[81]), .B(n26), .Z(c[81]) );
  XNOR U28 ( .A(b[80]), .B(n27), .Z(c[80]) );
  XNOR U29 ( .A(b[7]), .B(n28), .Z(c[7]) );
  XNOR U30 ( .A(b[79]), .B(n29), .Z(c[79]) );
  XNOR U31 ( .A(b[78]), .B(n30), .Z(c[78]) );
  XNOR U32 ( .A(b[77]), .B(n31), .Z(c[77]) );
  XNOR U33 ( .A(b[76]), .B(n32), .Z(c[76]) );
  XNOR U34 ( .A(b[75]), .B(n33), .Z(c[75]) );
  XNOR U35 ( .A(b[74]), .B(n34), .Z(c[74]) );
  XNOR U36 ( .A(b[73]), .B(n35), .Z(c[73]) );
  XNOR U37 ( .A(b[72]), .B(n36), .Z(c[72]) );
  XNOR U38 ( .A(b[71]), .B(n37), .Z(c[71]) );
  XNOR U39 ( .A(b[70]), .B(n38), .Z(c[70]) );
  XNOR U40 ( .A(b[6]), .B(n39), .Z(c[6]) );
  XNOR U41 ( .A(b[69]), .B(n40), .Z(c[69]) );
  XNOR U42 ( .A(b[68]), .B(n41), .Z(c[68]) );
  XNOR U43 ( .A(b[67]), .B(n42), .Z(c[67]) );
  XNOR U44 ( .A(b[66]), .B(n43), .Z(c[66]) );
  XNOR U45 ( .A(b[65]), .B(n44), .Z(c[65]) );
  XNOR U46 ( .A(b[64]), .B(n45), .Z(c[64]) );
  XNOR U47 ( .A(b[63]), .B(n46), .Z(c[63]) );
  XNOR U48 ( .A(b[62]), .B(n47), .Z(c[62]) );
  XNOR U49 ( .A(b[61]), .B(n48), .Z(c[61]) );
  XNOR U50 ( .A(b[60]), .B(n49), .Z(c[60]) );
  XNOR U51 ( .A(b[5]), .B(n50), .Z(c[5]) );
  XNOR U52 ( .A(b[59]), .B(n51), .Z(c[59]) );
  XNOR U53 ( .A(b[58]), .B(n52), .Z(c[58]) );
  XNOR U54 ( .A(b[57]), .B(n53), .Z(c[57]) );
  XNOR U55 ( .A(b[56]), .B(n54), .Z(c[56]) );
  XNOR U56 ( .A(b[55]), .B(n55), .Z(c[55]) );
  XNOR U57 ( .A(b[54]), .B(n56), .Z(c[54]) );
  XNOR U58 ( .A(b[53]), .B(n57), .Z(c[53]) );
  XNOR U59 ( .A(b[52]), .B(n58), .Z(c[52]) );
  XNOR U60 ( .A(b[51]), .B(n59), .Z(c[51]) );
  XNOR U61 ( .A(b[50]), .B(n60), .Z(c[50]) );
  XNOR U62 ( .A(b[4]), .B(n61), .Z(c[4]) );
  XNOR U63 ( .A(b[49]), .B(n62), .Z(c[49]) );
  XNOR U64 ( .A(b[48]), .B(n63), .Z(c[48]) );
  XNOR U65 ( .A(b[47]), .B(n64), .Z(c[47]) );
  XNOR U66 ( .A(b[46]), .B(n65), .Z(c[46]) );
  XNOR U67 ( .A(b[45]), .B(n66), .Z(c[45]) );
  XNOR U68 ( .A(b[44]), .B(n67), .Z(c[44]) );
  XNOR U69 ( .A(b[43]), .B(n68), .Z(c[43]) );
  XNOR U70 ( .A(b[42]), .B(n69), .Z(c[42]) );
  XNOR U71 ( .A(b[41]), .B(n70), .Z(c[41]) );
  XNOR U72 ( .A(b[40]), .B(n71), .Z(c[40]) );
  XNOR U73 ( .A(b[3]), .B(n72), .Z(c[3]) );
  XNOR U74 ( .A(b[39]), .B(n73), .Z(c[39]) );
  XNOR U75 ( .A(b[38]), .B(n74), .Z(c[38]) );
  XNOR U76 ( .A(b[37]), .B(n75), .Z(c[37]) );
  XNOR U77 ( .A(b[36]), .B(n76), .Z(c[36]) );
  XNOR U78 ( .A(b[35]), .B(n77), .Z(c[35]) );
  XNOR U79 ( .A(b[34]), .B(n78), .Z(c[34]) );
  XNOR U80 ( .A(b[33]), .B(n79), .Z(c[33]) );
  XNOR U81 ( .A(b[32]), .B(n80), .Z(c[32]) );
  XNOR U82 ( .A(b[31]), .B(n81), .Z(c[31]) );
  XNOR U83 ( .A(b[30]), .B(n82), .Z(c[30]) );
  XNOR U84 ( .A(b[2]), .B(n83), .Z(c[2]) );
  XNOR U85 ( .A(b[29]), .B(n84), .Z(c[29]) );
  XNOR U86 ( .A(b[28]), .B(n85), .Z(c[28]) );
  XNOR U87 ( .A(b[27]), .B(n86), .Z(c[27]) );
  XNOR U88 ( .A(b[26]), .B(n87), .Z(c[26]) );
  XNOR U89 ( .A(b[25]), .B(n88), .Z(c[25]) );
  XNOR U90 ( .A(b[255]), .B(n5), .Z(c[255]) );
  XNOR U91 ( .A(a[255]), .B(n3), .Z(n5) );
  XNOR U92 ( .A(n89), .B(n90), .Z(n3) );
  ANDN U93 ( .B(n91), .A(n92), .Z(n89) );
  XNOR U94 ( .A(b[254]), .B(n90), .Z(n91) );
  XNOR U95 ( .A(b[254]), .B(n92), .Z(c[254]) );
  XNOR U96 ( .A(a[254]), .B(n93), .Z(n92) );
  IV U97 ( .A(n90), .Z(n93) );
  XOR U98 ( .A(n94), .B(n95), .Z(n90) );
  ANDN U99 ( .B(n96), .A(n97), .Z(n94) );
  XNOR U100 ( .A(b[253]), .B(n95), .Z(n96) );
  XNOR U101 ( .A(b[253]), .B(n97), .Z(c[253]) );
  XNOR U102 ( .A(a[253]), .B(n98), .Z(n97) );
  IV U103 ( .A(n95), .Z(n98) );
  XOR U104 ( .A(n99), .B(n100), .Z(n95) );
  ANDN U105 ( .B(n101), .A(n102), .Z(n99) );
  XNOR U106 ( .A(b[252]), .B(n100), .Z(n101) );
  XNOR U107 ( .A(b[252]), .B(n102), .Z(c[252]) );
  XNOR U108 ( .A(a[252]), .B(n103), .Z(n102) );
  IV U109 ( .A(n100), .Z(n103) );
  XOR U110 ( .A(n104), .B(n105), .Z(n100) );
  ANDN U111 ( .B(n106), .A(n107), .Z(n104) );
  XNOR U112 ( .A(b[251]), .B(n105), .Z(n106) );
  XNOR U113 ( .A(b[251]), .B(n107), .Z(c[251]) );
  XNOR U114 ( .A(a[251]), .B(n108), .Z(n107) );
  IV U115 ( .A(n105), .Z(n108) );
  XOR U116 ( .A(n109), .B(n110), .Z(n105) );
  ANDN U117 ( .B(n111), .A(n112), .Z(n109) );
  XNOR U118 ( .A(b[250]), .B(n110), .Z(n111) );
  XNOR U119 ( .A(b[250]), .B(n112), .Z(c[250]) );
  XNOR U120 ( .A(a[250]), .B(n113), .Z(n112) );
  IV U121 ( .A(n110), .Z(n113) );
  XOR U122 ( .A(n114), .B(n115), .Z(n110) );
  ANDN U123 ( .B(n116), .A(n117), .Z(n114) );
  XNOR U124 ( .A(b[249]), .B(n115), .Z(n116) );
  XNOR U125 ( .A(b[24]), .B(n118), .Z(c[24]) );
  XNOR U126 ( .A(b[249]), .B(n117), .Z(c[249]) );
  XNOR U127 ( .A(a[249]), .B(n119), .Z(n117) );
  IV U128 ( .A(n115), .Z(n119) );
  XOR U129 ( .A(n120), .B(n121), .Z(n115) );
  ANDN U130 ( .B(n122), .A(n123), .Z(n120) );
  XNOR U131 ( .A(b[248]), .B(n121), .Z(n122) );
  XNOR U132 ( .A(b[248]), .B(n123), .Z(c[248]) );
  XNOR U133 ( .A(a[248]), .B(n124), .Z(n123) );
  IV U134 ( .A(n121), .Z(n124) );
  XOR U135 ( .A(n125), .B(n126), .Z(n121) );
  ANDN U136 ( .B(n127), .A(n128), .Z(n125) );
  XNOR U137 ( .A(b[247]), .B(n126), .Z(n127) );
  XNOR U138 ( .A(b[247]), .B(n128), .Z(c[247]) );
  XNOR U139 ( .A(a[247]), .B(n129), .Z(n128) );
  IV U140 ( .A(n126), .Z(n129) );
  XOR U141 ( .A(n130), .B(n131), .Z(n126) );
  ANDN U142 ( .B(n132), .A(n133), .Z(n130) );
  XNOR U143 ( .A(b[246]), .B(n131), .Z(n132) );
  XNOR U144 ( .A(b[246]), .B(n133), .Z(c[246]) );
  XNOR U145 ( .A(a[246]), .B(n134), .Z(n133) );
  IV U146 ( .A(n131), .Z(n134) );
  XOR U147 ( .A(n135), .B(n136), .Z(n131) );
  ANDN U148 ( .B(n137), .A(n138), .Z(n135) );
  XNOR U149 ( .A(b[245]), .B(n136), .Z(n137) );
  XNOR U150 ( .A(b[245]), .B(n138), .Z(c[245]) );
  XNOR U151 ( .A(a[245]), .B(n139), .Z(n138) );
  IV U152 ( .A(n136), .Z(n139) );
  XOR U153 ( .A(n140), .B(n141), .Z(n136) );
  ANDN U154 ( .B(n142), .A(n143), .Z(n140) );
  XNOR U155 ( .A(b[244]), .B(n141), .Z(n142) );
  XNOR U156 ( .A(b[244]), .B(n143), .Z(c[244]) );
  XNOR U157 ( .A(a[244]), .B(n144), .Z(n143) );
  IV U158 ( .A(n141), .Z(n144) );
  XOR U159 ( .A(n145), .B(n146), .Z(n141) );
  ANDN U160 ( .B(n147), .A(n148), .Z(n145) );
  XNOR U161 ( .A(b[243]), .B(n146), .Z(n147) );
  XNOR U162 ( .A(b[243]), .B(n148), .Z(c[243]) );
  XNOR U163 ( .A(a[243]), .B(n149), .Z(n148) );
  IV U164 ( .A(n146), .Z(n149) );
  XOR U165 ( .A(n150), .B(n151), .Z(n146) );
  ANDN U166 ( .B(n152), .A(n153), .Z(n150) );
  XNOR U167 ( .A(b[242]), .B(n151), .Z(n152) );
  XNOR U168 ( .A(b[242]), .B(n153), .Z(c[242]) );
  XNOR U169 ( .A(a[242]), .B(n154), .Z(n153) );
  IV U170 ( .A(n151), .Z(n154) );
  XOR U171 ( .A(n155), .B(n156), .Z(n151) );
  ANDN U172 ( .B(n157), .A(n158), .Z(n155) );
  XNOR U173 ( .A(b[241]), .B(n156), .Z(n157) );
  XNOR U174 ( .A(b[241]), .B(n158), .Z(c[241]) );
  XNOR U175 ( .A(a[241]), .B(n159), .Z(n158) );
  IV U176 ( .A(n156), .Z(n159) );
  XOR U177 ( .A(n160), .B(n161), .Z(n156) );
  ANDN U178 ( .B(n162), .A(n163), .Z(n160) );
  XNOR U179 ( .A(b[240]), .B(n161), .Z(n162) );
  XNOR U180 ( .A(b[240]), .B(n163), .Z(c[240]) );
  XNOR U181 ( .A(a[240]), .B(n164), .Z(n163) );
  IV U182 ( .A(n161), .Z(n164) );
  XOR U183 ( .A(n165), .B(n166), .Z(n161) );
  ANDN U184 ( .B(n167), .A(n168), .Z(n165) );
  XNOR U185 ( .A(b[239]), .B(n166), .Z(n167) );
  XNOR U186 ( .A(b[23]), .B(n169), .Z(c[23]) );
  XNOR U187 ( .A(b[239]), .B(n168), .Z(c[239]) );
  XNOR U188 ( .A(a[239]), .B(n170), .Z(n168) );
  IV U189 ( .A(n166), .Z(n170) );
  XOR U190 ( .A(n171), .B(n172), .Z(n166) );
  ANDN U191 ( .B(n173), .A(n174), .Z(n171) );
  XNOR U192 ( .A(b[238]), .B(n172), .Z(n173) );
  XNOR U193 ( .A(b[238]), .B(n174), .Z(c[238]) );
  XNOR U194 ( .A(a[238]), .B(n175), .Z(n174) );
  IV U195 ( .A(n172), .Z(n175) );
  XOR U196 ( .A(n176), .B(n177), .Z(n172) );
  ANDN U197 ( .B(n178), .A(n179), .Z(n176) );
  XNOR U198 ( .A(b[237]), .B(n177), .Z(n178) );
  XNOR U199 ( .A(b[237]), .B(n179), .Z(c[237]) );
  XNOR U200 ( .A(a[237]), .B(n180), .Z(n179) );
  IV U201 ( .A(n177), .Z(n180) );
  XOR U202 ( .A(n181), .B(n182), .Z(n177) );
  ANDN U203 ( .B(n183), .A(n184), .Z(n181) );
  XNOR U204 ( .A(b[236]), .B(n182), .Z(n183) );
  XNOR U205 ( .A(b[236]), .B(n184), .Z(c[236]) );
  XNOR U206 ( .A(a[236]), .B(n185), .Z(n184) );
  IV U207 ( .A(n182), .Z(n185) );
  XOR U208 ( .A(n186), .B(n187), .Z(n182) );
  ANDN U209 ( .B(n188), .A(n189), .Z(n186) );
  XNOR U210 ( .A(b[235]), .B(n187), .Z(n188) );
  XNOR U211 ( .A(b[235]), .B(n189), .Z(c[235]) );
  XNOR U212 ( .A(a[235]), .B(n190), .Z(n189) );
  IV U213 ( .A(n187), .Z(n190) );
  XOR U214 ( .A(n191), .B(n192), .Z(n187) );
  ANDN U215 ( .B(n193), .A(n194), .Z(n191) );
  XNOR U216 ( .A(b[234]), .B(n192), .Z(n193) );
  XNOR U217 ( .A(b[234]), .B(n194), .Z(c[234]) );
  XNOR U218 ( .A(a[234]), .B(n195), .Z(n194) );
  IV U219 ( .A(n192), .Z(n195) );
  XOR U220 ( .A(n196), .B(n197), .Z(n192) );
  ANDN U221 ( .B(n198), .A(n199), .Z(n196) );
  XNOR U222 ( .A(b[233]), .B(n197), .Z(n198) );
  XNOR U223 ( .A(b[233]), .B(n199), .Z(c[233]) );
  XNOR U224 ( .A(a[233]), .B(n200), .Z(n199) );
  IV U225 ( .A(n197), .Z(n200) );
  XOR U226 ( .A(n201), .B(n202), .Z(n197) );
  ANDN U227 ( .B(n203), .A(n204), .Z(n201) );
  XNOR U228 ( .A(b[232]), .B(n202), .Z(n203) );
  XNOR U229 ( .A(b[232]), .B(n204), .Z(c[232]) );
  XNOR U230 ( .A(a[232]), .B(n205), .Z(n204) );
  IV U231 ( .A(n202), .Z(n205) );
  XOR U232 ( .A(n206), .B(n207), .Z(n202) );
  ANDN U233 ( .B(n208), .A(n209), .Z(n206) );
  XNOR U234 ( .A(b[231]), .B(n207), .Z(n208) );
  XNOR U235 ( .A(b[231]), .B(n209), .Z(c[231]) );
  XNOR U236 ( .A(a[231]), .B(n210), .Z(n209) );
  IV U237 ( .A(n207), .Z(n210) );
  XOR U238 ( .A(n211), .B(n212), .Z(n207) );
  ANDN U239 ( .B(n213), .A(n214), .Z(n211) );
  XNOR U240 ( .A(b[230]), .B(n212), .Z(n213) );
  XNOR U241 ( .A(b[230]), .B(n214), .Z(c[230]) );
  XNOR U242 ( .A(a[230]), .B(n215), .Z(n214) );
  IV U243 ( .A(n212), .Z(n215) );
  XOR U244 ( .A(n216), .B(n217), .Z(n212) );
  ANDN U245 ( .B(n218), .A(n219), .Z(n216) );
  XNOR U246 ( .A(b[229]), .B(n217), .Z(n218) );
  XNOR U247 ( .A(b[22]), .B(n220), .Z(c[22]) );
  XNOR U248 ( .A(b[229]), .B(n219), .Z(c[229]) );
  XNOR U249 ( .A(a[229]), .B(n221), .Z(n219) );
  IV U250 ( .A(n217), .Z(n221) );
  XOR U251 ( .A(n222), .B(n223), .Z(n217) );
  ANDN U252 ( .B(n224), .A(n225), .Z(n222) );
  XNOR U253 ( .A(b[228]), .B(n223), .Z(n224) );
  XNOR U254 ( .A(b[228]), .B(n225), .Z(c[228]) );
  XNOR U255 ( .A(a[228]), .B(n226), .Z(n225) );
  IV U256 ( .A(n223), .Z(n226) );
  XOR U257 ( .A(n227), .B(n228), .Z(n223) );
  ANDN U258 ( .B(n229), .A(n230), .Z(n227) );
  XNOR U259 ( .A(b[227]), .B(n228), .Z(n229) );
  XNOR U260 ( .A(b[227]), .B(n230), .Z(c[227]) );
  XNOR U261 ( .A(a[227]), .B(n231), .Z(n230) );
  IV U262 ( .A(n228), .Z(n231) );
  XOR U263 ( .A(n232), .B(n233), .Z(n228) );
  ANDN U264 ( .B(n234), .A(n235), .Z(n232) );
  XNOR U265 ( .A(b[226]), .B(n233), .Z(n234) );
  XNOR U266 ( .A(b[226]), .B(n235), .Z(c[226]) );
  XNOR U267 ( .A(a[226]), .B(n236), .Z(n235) );
  IV U268 ( .A(n233), .Z(n236) );
  XOR U269 ( .A(n237), .B(n238), .Z(n233) );
  ANDN U270 ( .B(n239), .A(n240), .Z(n237) );
  XNOR U271 ( .A(b[225]), .B(n238), .Z(n239) );
  XNOR U272 ( .A(b[225]), .B(n240), .Z(c[225]) );
  XNOR U273 ( .A(a[225]), .B(n241), .Z(n240) );
  IV U274 ( .A(n238), .Z(n241) );
  XOR U275 ( .A(n242), .B(n243), .Z(n238) );
  ANDN U276 ( .B(n244), .A(n245), .Z(n242) );
  XNOR U277 ( .A(b[224]), .B(n243), .Z(n244) );
  XNOR U278 ( .A(b[224]), .B(n245), .Z(c[224]) );
  XNOR U279 ( .A(a[224]), .B(n246), .Z(n245) );
  IV U280 ( .A(n243), .Z(n246) );
  XOR U281 ( .A(n247), .B(n248), .Z(n243) );
  ANDN U282 ( .B(n249), .A(n250), .Z(n247) );
  XNOR U283 ( .A(b[223]), .B(n248), .Z(n249) );
  XNOR U284 ( .A(b[223]), .B(n250), .Z(c[223]) );
  XNOR U285 ( .A(a[223]), .B(n251), .Z(n250) );
  IV U286 ( .A(n248), .Z(n251) );
  XOR U287 ( .A(n252), .B(n253), .Z(n248) );
  ANDN U288 ( .B(n254), .A(n255), .Z(n252) );
  XNOR U289 ( .A(b[222]), .B(n253), .Z(n254) );
  XNOR U290 ( .A(b[222]), .B(n255), .Z(c[222]) );
  XNOR U291 ( .A(a[222]), .B(n256), .Z(n255) );
  IV U292 ( .A(n253), .Z(n256) );
  XOR U293 ( .A(n257), .B(n258), .Z(n253) );
  ANDN U294 ( .B(n259), .A(n260), .Z(n257) );
  XNOR U295 ( .A(b[221]), .B(n258), .Z(n259) );
  XNOR U296 ( .A(b[221]), .B(n260), .Z(c[221]) );
  XNOR U297 ( .A(a[221]), .B(n261), .Z(n260) );
  IV U298 ( .A(n258), .Z(n261) );
  XOR U299 ( .A(n262), .B(n263), .Z(n258) );
  ANDN U300 ( .B(n264), .A(n265), .Z(n262) );
  XNOR U301 ( .A(b[220]), .B(n263), .Z(n264) );
  XNOR U302 ( .A(b[220]), .B(n265), .Z(c[220]) );
  XNOR U303 ( .A(a[220]), .B(n266), .Z(n265) );
  IV U304 ( .A(n263), .Z(n266) );
  XOR U305 ( .A(n267), .B(n268), .Z(n263) );
  ANDN U306 ( .B(n269), .A(n270), .Z(n267) );
  XNOR U307 ( .A(b[219]), .B(n268), .Z(n269) );
  XNOR U308 ( .A(b[21]), .B(n271), .Z(c[21]) );
  XNOR U309 ( .A(b[219]), .B(n270), .Z(c[219]) );
  XNOR U310 ( .A(a[219]), .B(n272), .Z(n270) );
  IV U311 ( .A(n268), .Z(n272) );
  XOR U312 ( .A(n273), .B(n274), .Z(n268) );
  ANDN U313 ( .B(n275), .A(n276), .Z(n273) );
  XNOR U314 ( .A(b[218]), .B(n274), .Z(n275) );
  XNOR U315 ( .A(b[218]), .B(n276), .Z(c[218]) );
  XNOR U316 ( .A(a[218]), .B(n277), .Z(n276) );
  IV U317 ( .A(n274), .Z(n277) );
  XOR U318 ( .A(n278), .B(n279), .Z(n274) );
  ANDN U319 ( .B(n280), .A(n281), .Z(n278) );
  XNOR U320 ( .A(b[217]), .B(n279), .Z(n280) );
  XNOR U321 ( .A(b[217]), .B(n281), .Z(c[217]) );
  XNOR U322 ( .A(a[217]), .B(n282), .Z(n281) );
  IV U323 ( .A(n279), .Z(n282) );
  XOR U324 ( .A(n283), .B(n284), .Z(n279) );
  ANDN U325 ( .B(n285), .A(n286), .Z(n283) );
  XNOR U326 ( .A(b[216]), .B(n284), .Z(n285) );
  XNOR U327 ( .A(b[216]), .B(n286), .Z(c[216]) );
  XNOR U328 ( .A(a[216]), .B(n287), .Z(n286) );
  IV U329 ( .A(n284), .Z(n287) );
  XOR U330 ( .A(n288), .B(n289), .Z(n284) );
  ANDN U331 ( .B(n290), .A(n291), .Z(n288) );
  XNOR U332 ( .A(b[215]), .B(n289), .Z(n290) );
  XNOR U333 ( .A(b[215]), .B(n291), .Z(c[215]) );
  XNOR U334 ( .A(a[215]), .B(n292), .Z(n291) );
  IV U335 ( .A(n289), .Z(n292) );
  XOR U336 ( .A(n293), .B(n294), .Z(n289) );
  ANDN U337 ( .B(n295), .A(n296), .Z(n293) );
  XNOR U338 ( .A(b[214]), .B(n294), .Z(n295) );
  XNOR U339 ( .A(b[214]), .B(n296), .Z(c[214]) );
  XNOR U340 ( .A(a[214]), .B(n297), .Z(n296) );
  IV U341 ( .A(n294), .Z(n297) );
  XOR U342 ( .A(n298), .B(n299), .Z(n294) );
  ANDN U343 ( .B(n300), .A(n301), .Z(n298) );
  XNOR U344 ( .A(b[213]), .B(n299), .Z(n300) );
  XNOR U345 ( .A(b[213]), .B(n301), .Z(c[213]) );
  XNOR U346 ( .A(a[213]), .B(n302), .Z(n301) );
  IV U347 ( .A(n299), .Z(n302) );
  XOR U348 ( .A(n303), .B(n304), .Z(n299) );
  ANDN U349 ( .B(n305), .A(n306), .Z(n303) );
  XNOR U350 ( .A(b[212]), .B(n304), .Z(n305) );
  XNOR U351 ( .A(b[212]), .B(n306), .Z(c[212]) );
  XNOR U352 ( .A(a[212]), .B(n307), .Z(n306) );
  IV U353 ( .A(n304), .Z(n307) );
  XOR U354 ( .A(n308), .B(n309), .Z(n304) );
  ANDN U355 ( .B(n310), .A(n311), .Z(n308) );
  XNOR U356 ( .A(b[211]), .B(n309), .Z(n310) );
  XNOR U357 ( .A(b[211]), .B(n311), .Z(c[211]) );
  XNOR U358 ( .A(a[211]), .B(n312), .Z(n311) );
  IV U359 ( .A(n309), .Z(n312) );
  XOR U360 ( .A(n313), .B(n314), .Z(n309) );
  ANDN U361 ( .B(n315), .A(n316), .Z(n313) );
  XNOR U362 ( .A(b[210]), .B(n314), .Z(n315) );
  XNOR U363 ( .A(b[210]), .B(n316), .Z(c[210]) );
  XNOR U364 ( .A(a[210]), .B(n317), .Z(n316) );
  IV U365 ( .A(n314), .Z(n317) );
  XOR U366 ( .A(n318), .B(n319), .Z(n314) );
  ANDN U367 ( .B(n320), .A(n321), .Z(n318) );
  XNOR U368 ( .A(b[209]), .B(n319), .Z(n320) );
  XNOR U369 ( .A(b[20]), .B(n322), .Z(c[20]) );
  XNOR U370 ( .A(b[209]), .B(n321), .Z(c[209]) );
  XNOR U371 ( .A(a[209]), .B(n323), .Z(n321) );
  IV U372 ( .A(n319), .Z(n323) );
  XOR U373 ( .A(n324), .B(n325), .Z(n319) );
  ANDN U374 ( .B(n326), .A(n327), .Z(n324) );
  XNOR U375 ( .A(b[208]), .B(n325), .Z(n326) );
  XNOR U376 ( .A(b[208]), .B(n327), .Z(c[208]) );
  XNOR U377 ( .A(a[208]), .B(n328), .Z(n327) );
  IV U378 ( .A(n325), .Z(n328) );
  XOR U379 ( .A(n329), .B(n330), .Z(n325) );
  ANDN U380 ( .B(n331), .A(n332), .Z(n329) );
  XNOR U381 ( .A(b[207]), .B(n330), .Z(n331) );
  XNOR U382 ( .A(b[207]), .B(n332), .Z(c[207]) );
  XNOR U383 ( .A(a[207]), .B(n333), .Z(n332) );
  IV U384 ( .A(n330), .Z(n333) );
  XOR U385 ( .A(n334), .B(n335), .Z(n330) );
  ANDN U386 ( .B(n336), .A(n337), .Z(n334) );
  XNOR U387 ( .A(b[206]), .B(n335), .Z(n336) );
  XNOR U388 ( .A(b[206]), .B(n337), .Z(c[206]) );
  XNOR U389 ( .A(a[206]), .B(n338), .Z(n337) );
  IV U390 ( .A(n335), .Z(n338) );
  XOR U391 ( .A(n339), .B(n340), .Z(n335) );
  ANDN U392 ( .B(n341), .A(n342), .Z(n339) );
  XNOR U393 ( .A(b[205]), .B(n340), .Z(n341) );
  XNOR U394 ( .A(b[205]), .B(n342), .Z(c[205]) );
  XNOR U395 ( .A(a[205]), .B(n343), .Z(n342) );
  IV U396 ( .A(n340), .Z(n343) );
  XOR U397 ( .A(n344), .B(n345), .Z(n340) );
  ANDN U398 ( .B(n346), .A(n347), .Z(n344) );
  XNOR U399 ( .A(b[204]), .B(n345), .Z(n346) );
  XNOR U400 ( .A(b[204]), .B(n347), .Z(c[204]) );
  XNOR U401 ( .A(a[204]), .B(n348), .Z(n347) );
  IV U402 ( .A(n345), .Z(n348) );
  XOR U403 ( .A(n349), .B(n350), .Z(n345) );
  ANDN U404 ( .B(n351), .A(n352), .Z(n349) );
  XNOR U405 ( .A(b[203]), .B(n350), .Z(n351) );
  XNOR U406 ( .A(b[203]), .B(n352), .Z(c[203]) );
  XNOR U407 ( .A(a[203]), .B(n353), .Z(n352) );
  IV U408 ( .A(n350), .Z(n353) );
  XOR U409 ( .A(n354), .B(n355), .Z(n350) );
  ANDN U410 ( .B(n356), .A(n357), .Z(n354) );
  XNOR U411 ( .A(b[202]), .B(n355), .Z(n356) );
  XNOR U412 ( .A(b[202]), .B(n357), .Z(c[202]) );
  XNOR U413 ( .A(a[202]), .B(n358), .Z(n357) );
  IV U414 ( .A(n355), .Z(n358) );
  XOR U415 ( .A(n359), .B(n360), .Z(n355) );
  ANDN U416 ( .B(n361), .A(n362), .Z(n359) );
  XNOR U417 ( .A(b[201]), .B(n360), .Z(n361) );
  XNOR U418 ( .A(b[201]), .B(n362), .Z(c[201]) );
  XNOR U419 ( .A(a[201]), .B(n363), .Z(n362) );
  IV U420 ( .A(n360), .Z(n363) );
  XOR U421 ( .A(n364), .B(n365), .Z(n360) );
  ANDN U422 ( .B(n366), .A(n367), .Z(n364) );
  XNOR U423 ( .A(b[200]), .B(n365), .Z(n366) );
  XNOR U424 ( .A(b[200]), .B(n367), .Z(c[200]) );
  XNOR U425 ( .A(a[200]), .B(n368), .Z(n367) );
  IV U426 ( .A(n365), .Z(n368) );
  XOR U427 ( .A(n369), .B(n370), .Z(n365) );
  ANDN U428 ( .B(n371), .A(n372), .Z(n369) );
  XNOR U429 ( .A(b[199]), .B(n370), .Z(n371) );
  XNOR U430 ( .A(b[1]), .B(n373), .Z(c[1]) );
  XNOR U431 ( .A(b[19]), .B(n374), .Z(c[19]) );
  XNOR U432 ( .A(b[199]), .B(n372), .Z(c[199]) );
  XNOR U433 ( .A(a[199]), .B(n375), .Z(n372) );
  IV U434 ( .A(n370), .Z(n375) );
  XOR U435 ( .A(n376), .B(n377), .Z(n370) );
  ANDN U436 ( .B(n378), .A(n379), .Z(n376) );
  XNOR U437 ( .A(b[198]), .B(n377), .Z(n378) );
  XNOR U438 ( .A(b[198]), .B(n379), .Z(c[198]) );
  XNOR U439 ( .A(a[198]), .B(n380), .Z(n379) );
  IV U440 ( .A(n377), .Z(n380) );
  XOR U441 ( .A(n381), .B(n382), .Z(n377) );
  ANDN U442 ( .B(n383), .A(n384), .Z(n381) );
  XNOR U443 ( .A(b[197]), .B(n382), .Z(n383) );
  XNOR U444 ( .A(b[197]), .B(n384), .Z(c[197]) );
  XNOR U445 ( .A(a[197]), .B(n385), .Z(n384) );
  IV U446 ( .A(n382), .Z(n385) );
  XOR U447 ( .A(n386), .B(n387), .Z(n382) );
  ANDN U448 ( .B(n388), .A(n389), .Z(n386) );
  XNOR U449 ( .A(b[196]), .B(n387), .Z(n388) );
  XNOR U450 ( .A(b[196]), .B(n389), .Z(c[196]) );
  XNOR U451 ( .A(a[196]), .B(n390), .Z(n389) );
  IV U452 ( .A(n387), .Z(n390) );
  XOR U453 ( .A(n391), .B(n392), .Z(n387) );
  ANDN U454 ( .B(n393), .A(n394), .Z(n391) );
  XNOR U455 ( .A(b[195]), .B(n392), .Z(n393) );
  XNOR U456 ( .A(b[195]), .B(n394), .Z(c[195]) );
  XNOR U457 ( .A(a[195]), .B(n395), .Z(n394) );
  IV U458 ( .A(n392), .Z(n395) );
  XOR U459 ( .A(n396), .B(n397), .Z(n392) );
  ANDN U460 ( .B(n398), .A(n399), .Z(n396) );
  XNOR U461 ( .A(b[194]), .B(n397), .Z(n398) );
  XNOR U462 ( .A(b[194]), .B(n399), .Z(c[194]) );
  XNOR U463 ( .A(a[194]), .B(n400), .Z(n399) );
  IV U464 ( .A(n397), .Z(n400) );
  XOR U465 ( .A(n401), .B(n402), .Z(n397) );
  ANDN U466 ( .B(n403), .A(n404), .Z(n401) );
  XNOR U467 ( .A(b[193]), .B(n402), .Z(n403) );
  XNOR U468 ( .A(b[193]), .B(n404), .Z(c[193]) );
  XNOR U469 ( .A(a[193]), .B(n405), .Z(n404) );
  IV U470 ( .A(n402), .Z(n405) );
  XOR U471 ( .A(n406), .B(n407), .Z(n402) );
  ANDN U472 ( .B(n408), .A(n409), .Z(n406) );
  XNOR U473 ( .A(b[192]), .B(n407), .Z(n408) );
  XNOR U474 ( .A(b[192]), .B(n409), .Z(c[192]) );
  XNOR U475 ( .A(a[192]), .B(n410), .Z(n409) );
  IV U476 ( .A(n407), .Z(n410) );
  XOR U477 ( .A(n411), .B(n412), .Z(n407) );
  ANDN U478 ( .B(n413), .A(n414), .Z(n411) );
  XNOR U479 ( .A(b[191]), .B(n412), .Z(n413) );
  XNOR U480 ( .A(b[191]), .B(n414), .Z(c[191]) );
  XNOR U481 ( .A(a[191]), .B(n415), .Z(n414) );
  IV U482 ( .A(n412), .Z(n415) );
  XOR U483 ( .A(n416), .B(n417), .Z(n412) );
  ANDN U484 ( .B(n418), .A(n419), .Z(n416) );
  XNOR U485 ( .A(b[190]), .B(n417), .Z(n418) );
  XNOR U486 ( .A(b[190]), .B(n419), .Z(c[190]) );
  XNOR U487 ( .A(a[190]), .B(n420), .Z(n419) );
  IV U488 ( .A(n417), .Z(n420) );
  XOR U489 ( .A(n421), .B(n422), .Z(n417) );
  ANDN U490 ( .B(n423), .A(n424), .Z(n421) );
  XNOR U491 ( .A(b[189]), .B(n422), .Z(n423) );
  XNOR U492 ( .A(b[18]), .B(n425), .Z(c[18]) );
  XNOR U493 ( .A(b[189]), .B(n424), .Z(c[189]) );
  XNOR U494 ( .A(a[189]), .B(n426), .Z(n424) );
  IV U495 ( .A(n422), .Z(n426) );
  XOR U496 ( .A(n427), .B(n428), .Z(n422) );
  ANDN U497 ( .B(n429), .A(n430), .Z(n427) );
  XNOR U498 ( .A(b[188]), .B(n428), .Z(n429) );
  XNOR U499 ( .A(b[188]), .B(n430), .Z(c[188]) );
  XNOR U500 ( .A(a[188]), .B(n431), .Z(n430) );
  IV U501 ( .A(n428), .Z(n431) );
  XOR U502 ( .A(n432), .B(n433), .Z(n428) );
  ANDN U503 ( .B(n434), .A(n435), .Z(n432) );
  XNOR U504 ( .A(b[187]), .B(n433), .Z(n434) );
  XNOR U505 ( .A(b[187]), .B(n435), .Z(c[187]) );
  XNOR U506 ( .A(a[187]), .B(n436), .Z(n435) );
  IV U507 ( .A(n433), .Z(n436) );
  XOR U508 ( .A(n437), .B(n438), .Z(n433) );
  ANDN U509 ( .B(n439), .A(n440), .Z(n437) );
  XNOR U510 ( .A(b[186]), .B(n438), .Z(n439) );
  XNOR U511 ( .A(b[186]), .B(n440), .Z(c[186]) );
  XNOR U512 ( .A(a[186]), .B(n441), .Z(n440) );
  IV U513 ( .A(n438), .Z(n441) );
  XOR U514 ( .A(n442), .B(n443), .Z(n438) );
  ANDN U515 ( .B(n444), .A(n445), .Z(n442) );
  XNOR U516 ( .A(b[185]), .B(n443), .Z(n444) );
  XNOR U517 ( .A(b[185]), .B(n445), .Z(c[185]) );
  XNOR U518 ( .A(a[185]), .B(n446), .Z(n445) );
  IV U519 ( .A(n443), .Z(n446) );
  XOR U520 ( .A(n447), .B(n448), .Z(n443) );
  ANDN U521 ( .B(n449), .A(n450), .Z(n447) );
  XNOR U522 ( .A(b[184]), .B(n448), .Z(n449) );
  XNOR U523 ( .A(b[184]), .B(n450), .Z(c[184]) );
  XNOR U524 ( .A(a[184]), .B(n451), .Z(n450) );
  IV U525 ( .A(n448), .Z(n451) );
  XOR U526 ( .A(n452), .B(n453), .Z(n448) );
  ANDN U527 ( .B(n454), .A(n455), .Z(n452) );
  XNOR U528 ( .A(b[183]), .B(n453), .Z(n454) );
  XNOR U529 ( .A(b[183]), .B(n455), .Z(c[183]) );
  XNOR U530 ( .A(a[183]), .B(n456), .Z(n455) );
  IV U531 ( .A(n453), .Z(n456) );
  XOR U532 ( .A(n457), .B(n458), .Z(n453) );
  ANDN U533 ( .B(n459), .A(n460), .Z(n457) );
  XNOR U534 ( .A(b[182]), .B(n458), .Z(n459) );
  XNOR U535 ( .A(b[182]), .B(n460), .Z(c[182]) );
  XNOR U536 ( .A(a[182]), .B(n461), .Z(n460) );
  IV U537 ( .A(n458), .Z(n461) );
  XOR U538 ( .A(n462), .B(n463), .Z(n458) );
  ANDN U539 ( .B(n464), .A(n465), .Z(n462) );
  XNOR U540 ( .A(b[181]), .B(n463), .Z(n464) );
  XNOR U541 ( .A(b[181]), .B(n465), .Z(c[181]) );
  XNOR U542 ( .A(a[181]), .B(n466), .Z(n465) );
  IV U543 ( .A(n463), .Z(n466) );
  XOR U544 ( .A(n467), .B(n468), .Z(n463) );
  ANDN U545 ( .B(n469), .A(n470), .Z(n467) );
  XNOR U546 ( .A(b[180]), .B(n468), .Z(n469) );
  XNOR U547 ( .A(b[180]), .B(n470), .Z(c[180]) );
  XNOR U548 ( .A(a[180]), .B(n471), .Z(n470) );
  IV U549 ( .A(n468), .Z(n471) );
  XOR U550 ( .A(n472), .B(n473), .Z(n468) );
  ANDN U551 ( .B(n474), .A(n475), .Z(n472) );
  XNOR U552 ( .A(b[179]), .B(n473), .Z(n474) );
  XNOR U553 ( .A(b[17]), .B(n476), .Z(c[17]) );
  XNOR U554 ( .A(b[179]), .B(n475), .Z(c[179]) );
  XNOR U555 ( .A(a[179]), .B(n477), .Z(n475) );
  IV U556 ( .A(n473), .Z(n477) );
  XOR U557 ( .A(n478), .B(n479), .Z(n473) );
  ANDN U558 ( .B(n480), .A(n481), .Z(n478) );
  XNOR U559 ( .A(b[178]), .B(n479), .Z(n480) );
  XNOR U560 ( .A(b[178]), .B(n481), .Z(c[178]) );
  XNOR U561 ( .A(a[178]), .B(n482), .Z(n481) );
  IV U562 ( .A(n479), .Z(n482) );
  XOR U563 ( .A(n483), .B(n484), .Z(n479) );
  ANDN U564 ( .B(n485), .A(n486), .Z(n483) );
  XNOR U565 ( .A(b[177]), .B(n484), .Z(n485) );
  XNOR U566 ( .A(b[177]), .B(n486), .Z(c[177]) );
  XNOR U567 ( .A(a[177]), .B(n487), .Z(n486) );
  IV U568 ( .A(n484), .Z(n487) );
  XOR U569 ( .A(n488), .B(n489), .Z(n484) );
  ANDN U570 ( .B(n490), .A(n491), .Z(n488) );
  XNOR U571 ( .A(b[176]), .B(n489), .Z(n490) );
  XNOR U572 ( .A(b[176]), .B(n491), .Z(c[176]) );
  XNOR U573 ( .A(a[176]), .B(n492), .Z(n491) );
  IV U574 ( .A(n489), .Z(n492) );
  XOR U575 ( .A(n493), .B(n494), .Z(n489) );
  ANDN U576 ( .B(n495), .A(n496), .Z(n493) );
  XNOR U577 ( .A(b[175]), .B(n494), .Z(n495) );
  XNOR U578 ( .A(b[175]), .B(n496), .Z(c[175]) );
  XNOR U579 ( .A(a[175]), .B(n497), .Z(n496) );
  IV U580 ( .A(n494), .Z(n497) );
  XOR U581 ( .A(n498), .B(n499), .Z(n494) );
  ANDN U582 ( .B(n500), .A(n501), .Z(n498) );
  XNOR U583 ( .A(b[174]), .B(n499), .Z(n500) );
  XNOR U584 ( .A(b[174]), .B(n501), .Z(c[174]) );
  XNOR U585 ( .A(a[174]), .B(n502), .Z(n501) );
  IV U586 ( .A(n499), .Z(n502) );
  XOR U587 ( .A(n503), .B(n504), .Z(n499) );
  ANDN U588 ( .B(n505), .A(n506), .Z(n503) );
  XNOR U589 ( .A(b[173]), .B(n504), .Z(n505) );
  XNOR U590 ( .A(b[173]), .B(n506), .Z(c[173]) );
  XNOR U591 ( .A(a[173]), .B(n507), .Z(n506) );
  IV U592 ( .A(n504), .Z(n507) );
  XOR U593 ( .A(n508), .B(n509), .Z(n504) );
  ANDN U594 ( .B(n510), .A(n511), .Z(n508) );
  XNOR U595 ( .A(b[172]), .B(n509), .Z(n510) );
  XNOR U596 ( .A(b[172]), .B(n511), .Z(c[172]) );
  XNOR U597 ( .A(a[172]), .B(n512), .Z(n511) );
  IV U598 ( .A(n509), .Z(n512) );
  XOR U599 ( .A(n513), .B(n514), .Z(n509) );
  ANDN U600 ( .B(n515), .A(n516), .Z(n513) );
  XNOR U601 ( .A(b[171]), .B(n514), .Z(n515) );
  XNOR U602 ( .A(b[171]), .B(n516), .Z(c[171]) );
  XNOR U603 ( .A(a[171]), .B(n517), .Z(n516) );
  IV U604 ( .A(n514), .Z(n517) );
  XOR U605 ( .A(n518), .B(n519), .Z(n514) );
  ANDN U606 ( .B(n520), .A(n521), .Z(n518) );
  XNOR U607 ( .A(b[170]), .B(n519), .Z(n520) );
  XNOR U608 ( .A(b[170]), .B(n521), .Z(c[170]) );
  XNOR U609 ( .A(a[170]), .B(n522), .Z(n521) );
  IV U610 ( .A(n519), .Z(n522) );
  XOR U611 ( .A(n523), .B(n524), .Z(n519) );
  ANDN U612 ( .B(n525), .A(n526), .Z(n523) );
  XNOR U613 ( .A(b[169]), .B(n524), .Z(n525) );
  XNOR U614 ( .A(b[16]), .B(n527), .Z(c[16]) );
  XNOR U615 ( .A(b[169]), .B(n526), .Z(c[169]) );
  XNOR U616 ( .A(a[169]), .B(n528), .Z(n526) );
  IV U617 ( .A(n524), .Z(n528) );
  XOR U618 ( .A(n529), .B(n530), .Z(n524) );
  ANDN U619 ( .B(n531), .A(n532), .Z(n529) );
  XNOR U620 ( .A(b[168]), .B(n530), .Z(n531) );
  XNOR U621 ( .A(b[168]), .B(n532), .Z(c[168]) );
  XNOR U622 ( .A(a[168]), .B(n533), .Z(n532) );
  IV U623 ( .A(n530), .Z(n533) );
  XOR U624 ( .A(n534), .B(n535), .Z(n530) );
  ANDN U625 ( .B(n536), .A(n537), .Z(n534) );
  XNOR U626 ( .A(b[167]), .B(n535), .Z(n536) );
  XNOR U627 ( .A(b[167]), .B(n537), .Z(c[167]) );
  XNOR U628 ( .A(a[167]), .B(n538), .Z(n537) );
  IV U629 ( .A(n535), .Z(n538) );
  XOR U630 ( .A(n539), .B(n540), .Z(n535) );
  ANDN U631 ( .B(n541), .A(n542), .Z(n539) );
  XNOR U632 ( .A(b[166]), .B(n540), .Z(n541) );
  XNOR U633 ( .A(b[166]), .B(n542), .Z(c[166]) );
  XNOR U634 ( .A(a[166]), .B(n543), .Z(n542) );
  IV U635 ( .A(n540), .Z(n543) );
  XOR U636 ( .A(n544), .B(n545), .Z(n540) );
  ANDN U637 ( .B(n546), .A(n547), .Z(n544) );
  XNOR U638 ( .A(b[165]), .B(n545), .Z(n546) );
  XNOR U639 ( .A(b[165]), .B(n547), .Z(c[165]) );
  XNOR U640 ( .A(a[165]), .B(n548), .Z(n547) );
  IV U641 ( .A(n545), .Z(n548) );
  XOR U642 ( .A(n549), .B(n550), .Z(n545) );
  ANDN U643 ( .B(n551), .A(n552), .Z(n549) );
  XNOR U644 ( .A(b[164]), .B(n550), .Z(n551) );
  XNOR U645 ( .A(b[164]), .B(n552), .Z(c[164]) );
  XNOR U646 ( .A(a[164]), .B(n553), .Z(n552) );
  IV U647 ( .A(n550), .Z(n553) );
  XOR U648 ( .A(n554), .B(n555), .Z(n550) );
  ANDN U649 ( .B(n556), .A(n557), .Z(n554) );
  XNOR U650 ( .A(b[163]), .B(n555), .Z(n556) );
  XNOR U651 ( .A(b[163]), .B(n557), .Z(c[163]) );
  XNOR U652 ( .A(a[163]), .B(n558), .Z(n557) );
  IV U653 ( .A(n555), .Z(n558) );
  XOR U654 ( .A(n559), .B(n560), .Z(n555) );
  ANDN U655 ( .B(n561), .A(n562), .Z(n559) );
  XNOR U656 ( .A(b[162]), .B(n560), .Z(n561) );
  XNOR U657 ( .A(b[162]), .B(n562), .Z(c[162]) );
  XNOR U658 ( .A(a[162]), .B(n563), .Z(n562) );
  IV U659 ( .A(n560), .Z(n563) );
  XOR U660 ( .A(n564), .B(n565), .Z(n560) );
  ANDN U661 ( .B(n566), .A(n567), .Z(n564) );
  XNOR U662 ( .A(b[161]), .B(n565), .Z(n566) );
  XNOR U663 ( .A(b[161]), .B(n567), .Z(c[161]) );
  XNOR U664 ( .A(a[161]), .B(n568), .Z(n567) );
  IV U665 ( .A(n565), .Z(n568) );
  XOR U666 ( .A(n569), .B(n570), .Z(n565) );
  ANDN U667 ( .B(n571), .A(n572), .Z(n569) );
  XNOR U668 ( .A(b[160]), .B(n570), .Z(n571) );
  XNOR U669 ( .A(b[160]), .B(n572), .Z(c[160]) );
  XNOR U670 ( .A(a[160]), .B(n573), .Z(n572) );
  IV U671 ( .A(n570), .Z(n573) );
  XOR U672 ( .A(n574), .B(n575), .Z(n570) );
  ANDN U673 ( .B(n576), .A(n577), .Z(n574) );
  XNOR U674 ( .A(b[159]), .B(n575), .Z(n576) );
  XNOR U675 ( .A(b[15]), .B(n578), .Z(c[15]) );
  XNOR U676 ( .A(b[159]), .B(n577), .Z(c[159]) );
  XNOR U677 ( .A(a[159]), .B(n579), .Z(n577) );
  IV U678 ( .A(n575), .Z(n579) );
  XOR U679 ( .A(n580), .B(n581), .Z(n575) );
  ANDN U680 ( .B(n582), .A(n583), .Z(n580) );
  XNOR U681 ( .A(b[158]), .B(n581), .Z(n582) );
  XNOR U682 ( .A(b[158]), .B(n583), .Z(c[158]) );
  XNOR U683 ( .A(a[158]), .B(n584), .Z(n583) );
  IV U684 ( .A(n581), .Z(n584) );
  XOR U685 ( .A(n585), .B(n586), .Z(n581) );
  ANDN U686 ( .B(n587), .A(n588), .Z(n585) );
  XNOR U687 ( .A(b[157]), .B(n586), .Z(n587) );
  XNOR U688 ( .A(b[157]), .B(n588), .Z(c[157]) );
  XNOR U689 ( .A(a[157]), .B(n589), .Z(n588) );
  IV U690 ( .A(n586), .Z(n589) );
  XOR U691 ( .A(n590), .B(n591), .Z(n586) );
  ANDN U692 ( .B(n592), .A(n593), .Z(n590) );
  XNOR U693 ( .A(b[156]), .B(n591), .Z(n592) );
  XNOR U694 ( .A(b[156]), .B(n593), .Z(c[156]) );
  XNOR U695 ( .A(a[156]), .B(n594), .Z(n593) );
  IV U696 ( .A(n591), .Z(n594) );
  XOR U697 ( .A(n595), .B(n596), .Z(n591) );
  ANDN U698 ( .B(n597), .A(n598), .Z(n595) );
  XNOR U699 ( .A(b[155]), .B(n596), .Z(n597) );
  XNOR U700 ( .A(b[155]), .B(n598), .Z(c[155]) );
  XNOR U701 ( .A(a[155]), .B(n599), .Z(n598) );
  IV U702 ( .A(n596), .Z(n599) );
  XOR U703 ( .A(n600), .B(n601), .Z(n596) );
  ANDN U704 ( .B(n602), .A(n603), .Z(n600) );
  XNOR U705 ( .A(b[154]), .B(n601), .Z(n602) );
  XNOR U706 ( .A(b[154]), .B(n603), .Z(c[154]) );
  XNOR U707 ( .A(a[154]), .B(n604), .Z(n603) );
  IV U708 ( .A(n601), .Z(n604) );
  XOR U709 ( .A(n605), .B(n606), .Z(n601) );
  ANDN U710 ( .B(n607), .A(n608), .Z(n605) );
  XNOR U711 ( .A(b[153]), .B(n606), .Z(n607) );
  XNOR U712 ( .A(b[153]), .B(n608), .Z(c[153]) );
  XNOR U713 ( .A(a[153]), .B(n609), .Z(n608) );
  IV U714 ( .A(n606), .Z(n609) );
  XOR U715 ( .A(n610), .B(n611), .Z(n606) );
  ANDN U716 ( .B(n612), .A(n613), .Z(n610) );
  XNOR U717 ( .A(b[152]), .B(n611), .Z(n612) );
  XNOR U718 ( .A(b[152]), .B(n613), .Z(c[152]) );
  XNOR U719 ( .A(a[152]), .B(n614), .Z(n613) );
  IV U720 ( .A(n611), .Z(n614) );
  XOR U721 ( .A(n615), .B(n616), .Z(n611) );
  ANDN U722 ( .B(n617), .A(n618), .Z(n615) );
  XNOR U723 ( .A(b[151]), .B(n616), .Z(n617) );
  XNOR U724 ( .A(b[151]), .B(n618), .Z(c[151]) );
  XNOR U725 ( .A(a[151]), .B(n619), .Z(n618) );
  IV U726 ( .A(n616), .Z(n619) );
  XOR U727 ( .A(n620), .B(n621), .Z(n616) );
  ANDN U728 ( .B(n622), .A(n623), .Z(n620) );
  XNOR U729 ( .A(b[150]), .B(n621), .Z(n622) );
  XNOR U730 ( .A(b[150]), .B(n623), .Z(c[150]) );
  XNOR U731 ( .A(a[150]), .B(n624), .Z(n623) );
  IV U732 ( .A(n621), .Z(n624) );
  XOR U733 ( .A(n625), .B(n626), .Z(n621) );
  ANDN U734 ( .B(n627), .A(n628), .Z(n625) );
  XNOR U735 ( .A(b[149]), .B(n626), .Z(n627) );
  XNOR U736 ( .A(b[14]), .B(n629), .Z(c[14]) );
  XNOR U737 ( .A(b[149]), .B(n628), .Z(c[149]) );
  XNOR U738 ( .A(a[149]), .B(n630), .Z(n628) );
  IV U739 ( .A(n626), .Z(n630) );
  XOR U740 ( .A(n631), .B(n632), .Z(n626) );
  ANDN U741 ( .B(n633), .A(n634), .Z(n631) );
  XNOR U742 ( .A(b[148]), .B(n632), .Z(n633) );
  XNOR U743 ( .A(b[148]), .B(n634), .Z(c[148]) );
  XNOR U744 ( .A(a[148]), .B(n635), .Z(n634) );
  IV U745 ( .A(n632), .Z(n635) );
  XOR U746 ( .A(n636), .B(n637), .Z(n632) );
  ANDN U747 ( .B(n638), .A(n639), .Z(n636) );
  XNOR U748 ( .A(b[147]), .B(n637), .Z(n638) );
  XNOR U749 ( .A(b[147]), .B(n639), .Z(c[147]) );
  XNOR U750 ( .A(a[147]), .B(n640), .Z(n639) );
  IV U751 ( .A(n637), .Z(n640) );
  XOR U752 ( .A(n641), .B(n642), .Z(n637) );
  ANDN U753 ( .B(n643), .A(n644), .Z(n641) );
  XNOR U754 ( .A(b[146]), .B(n642), .Z(n643) );
  XNOR U755 ( .A(b[146]), .B(n644), .Z(c[146]) );
  XNOR U756 ( .A(a[146]), .B(n645), .Z(n644) );
  IV U757 ( .A(n642), .Z(n645) );
  XOR U758 ( .A(n646), .B(n647), .Z(n642) );
  ANDN U759 ( .B(n648), .A(n649), .Z(n646) );
  XNOR U760 ( .A(b[145]), .B(n647), .Z(n648) );
  XNOR U761 ( .A(b[145]), .B(n649), .Z(c[145]) );
  XNOR U762 ( .A(a[145]), .B(n650), .Z(n649) );
  IV U763 ( .A(n647), .Z(n650) );
  XOR U764 ( .A(n651), .B(n652), .Z(n647) );
  ANDN U765 ( .B(n653), .A(n654), .Z(n651) );
  XNOR U766 ( .A(b[144]), .B(n652), .Z(n653) );
  XNOR U767 ( .A(b[144]), .B(n654), .Z(c[144]) );
  XNOR U768 ( .A(a[144]), .B(n655), .Z(n654) );
  IV U769 ( .A(n652), .Z(n655) );
  XOR U770 ( .A(n656), .B(n657), .Z(n652) );
  ANDN U771 ( .B(n658), .A(n659), .Z(n656) );
  XNOR U772 ( .A(b[143]), .B(n657), .Z(n658) );
  XNOR U773 ( .A(b[143]), .B(n659), .Z(c[143]) );
  XNOR U774 ( .A(a[143]), .B(n660), .Z(n659) );
  IV U775 ( .A(n657), .Z(n660) );
  XOR U776 ( .A(n661), .B(n662), .Z(n657) );
  ANDN U777 ( .B(n663), .A(n664), .Z(n661) );
  XNOR U778 ( .A(b[142]), .B(n662), .Z(n663) );
  XNOR U779 ( .A(b[142]), .B(n664), .Z(c[142]) );
  XNOR U780 ( .A(a[142]), .B(n665), .Z(n664) );
  IV U781 ( .A(n662), .Z(n665) );
  XOR U782 ( .A(n666), .B(n667), .Z(n662) );
  ANDN U783 ( .B(n668), .A(n669), .Z(n666) );
  XNOR U784 ( .A(b[141]), .B(n667), .Z(n668) );
  XNOR U785 ( .A(b[141]), .B(n669), .Z(c[141]) );
  XNOR U786 ( .A(a[141]), .B(n670), .Z(n669) );
  IV U787 ( .A(n667), .Z(n670) );
  XOR U788 ( .A(n671), .B(n672), .Z(n667) );
  ANDN U789 ( .B(n673), .A(n674), .Z(n671) );
  XNOR U790 ( .A(b[140]), .B(n672), .Z(n673) );
  XNOR U791 ( .A(b[140]), .B(n674), .Z(c[140]) );
  XNOR U792 ( .A(a[140]), .B(n675), .Z(n674) );
  IV U793 ( .A(n672), .Z(n675) );
  XOR U794 ( .A(n676), .B(n677), .Z(n672) );
  ANDN U795 ( .B(n678), .A(n679), .Z(n676) );
  XNOR U796 ( .A(b[139]), .B(n677), .Z(n678) );
  XNOR U797 ( .A(b[13]), .B(n680), .Z(c[13]) );
  XNOR U798 ( .A(b[139]), .B(n679), .Z(c[139]) );
  XNOR U799 ( .A(a[139]), .B(n681), .Z(n679) );
  IV U800 ( .A(n677), .Z(n681) );
  XOR U801 ( .A(n682), .B(n683), .Z(n677) );
  ANDN U802 ( .B(n684), .A(n685), .Z(n682) );
  XNOR U803 ( .A(b[138]), .B(n683), .Z(n684) );
  XNOR U804 ( .A(b[138]), .B(n685), .Z(c[138]) );
  XNOR U805 ( .A(a[138]), .B(n686), .Z(n685) );
  IV U806 ( .A(n683), .Z(n686) );
  XOR U807 ( .A(n687), .B(n688), .Z(n683) );
  ANDN U808 ( .B(n689), .A(n690), .Z(n687) );
  XNOR U809 ( .A(b[137]), .B(n688), .Z(n689) );
  XNOR U810 ( .A(b[137]), .B(n690), .Z(c[137]) );
  XNOR U811 ( .A(a[137]), .B(n691), .Z(n690) );
  IV U812 ( .A(n688), .Z(n691) );
  XOR U813 ( .A(n692), .B(n693), .Z(n688) );
  ANDN U814 ( .B(n694), .A(n695), .Z(n692) );
  XNOR U815 ( .A(b[136]), .B(n693), .Z(n694) );
  XNOR U816 ( .A(b[136]), .B(n695), .Z(c[136]) );
  XNOR U817 ( .A(a[136]), .B(n696), .Z(n695) );
  IV U818 ( .A(n693), .Z(n696) );
  XOR U819 ( .A(n697), .B(n698), .Z(n693) );
  ANDN U820 ( .B(n699), .A(n700), .Z(n697) );
  XNOR U821 ( .A(b[135]), .B(n698), .Z(n699) );
  XNOR U822 ( .A(b[135]), .B(n700), .Z(c[135]) );
  XNOR U823 ( .A(a[135]), .B(n701), .Z(n700) );
  IV U824 ( .A(n698), .Z(n701) );
  XOR U825 ( .A(n702), .B(n703), .Z(n698) );
  ANDN U826 ( .B(n704), .A(n705), .Z(n702) );
  XNOR U827 ( .A(b[134]), .B(n703), .Z(n704) );
  XNOR U828 ( .A(b[134]), .B(n705), .Z(c[134]) );
  XNOR U829 ( .A(a[134]), .B(n706), .Z(n705) );
  IV U830 ( .A(n703), .Z(n706) );
  XOR U831 ( .A(n707), .B(n708), .Z(n703) );
  ANDN U832 ( .B(n709), .A(n710), .Z(n707) );
  XNOR U833 ( .A(b[133]), .B(n708), .Z(n709) );
  XNOR U834 ( .A(b[133]), .B(n710), .Z(c[133]) );
  XNOR U835 ( .A(a[133]), .B(n711), .Z(n710) );
  IV U836 ( .A(n708), .Z(n711) );
  XOR U837 ( .A(n712), .B(n713), .Z(n708) );
  ANDN U838 ( .B(n714), .A(n715), .Z(n712) );
  XNOR U839 ( .A(b[132]), .B(n713), .Z(n714) );
  XNOR U840 ( .A(b[132]), .B(n715), .Z(c[132]) );
  XNOR U841 ( .A(a[132]), .B(n716), .Z(n715) );
  IV U842 ( .A(n713), .Z(n716) );
  XOR U843 ( .A(n717), .B(n718), .Z(n713) );
  ANDN U844 ( .B(n719), .A(n720), .Z(n717) );
  XNOR U845 ( .A(b[131]), .B(n718), .Z(n719) );
  XNOR U846 ( .A(b[131]), .B(n720), .Z(c[131]) );
  XNOR U847 ( .A(a[131]), .B(n721), .Z(n720) );
  IV U848 ( .A(n718), .Z(n721) );
  XOR U849 ( .A(n722), .B(n723), .Z(n718) );
  ANDN U850 ( .B(n724), .A(n725), .Z(n722) );
  XNOR U851 ( .A(b[130]), .B(n723), .Z(n724) );
  XNOR U852 ( .A(b[130]), .B(n725), .Z(c[130]) );
  XNOR U853 ( .A(a[130]), .B(n726), .Z(n725) );
  IV U854 ( .A(n723), .Z(n726) );
  XOR U855 ( .A(n727), .B(n728), .Z(n723) );
  ANDN U856 ( .B(n729), .A(n730), .Z(n727) );
  XNOR U857 ( .A(b[129]), .B(n728), .Z(n729) );
  XNOR U858 ( .A(b[12]), .B(n731), .Z(c[12]) );
  XNOR U859 ( .A(b[129]), .B(n730), .Z(c[129]) );
  XNOR U860 ( .A(a[129]), .B(n732), .Z(n730) );
  IV U861 ( .A(n728), .Z(n732) );
  XOR U862 ( .A(n733), .B(n734), .Z(n728) );
  ANDN U863 ( .B(n735), .A(n736), .Z(n733) );
  XNOR U864 ( .A(b[128]), .B(n734), .Z(n735) );
  XNOR U865 ( .A(b[128]), .B(n736), .Z(c[128]) );
  XNOR U866 ( .A(a[128]), .B(n737), .Z(n736) );
  IV U867 ( .A(n734), .Z(n737) );
  XOR U868 ( .A(n738), .B(n739), .Z(n734) );
  ANDN U869 ( .B(n740), .A(n741), .Z(n738) );
  XNOR U870 ( .A(b[127]), .B(n739), .Z(n740) );
  XNOR U871 ( .A(b[127]), .B(n741), .Z(c[127]) );
  XNOR U872 ( .A(a[127]), .B(n742), .Z(n741) );
  IV U873 ( .A(n739), .Z(n742) );
  XOR U874 ( .A(n743), .B(n744), .Z(n739) );
  ANDN U875 ( .B(n745), .A(n746), .Z(n743) );
  XNOR U876 ( .A(b[126]), .B(n744), .Z(n745) );
  XNOR U877 ( .A(b[126]), .B(n746), .Z(c[126]) );
  XNOR U878 ( .A(a[126]), .B(n747), .Z(n746) );
  IV U879 ( .A(n744), .Z(n747) );
  XOR U880 ( .A(n748), .B(n749), .Z(n744) );
  ANDN U881 ( .B(n750), .A(n751), .Z(n748) );
  XNOR U882 ( .A(b[125]), .B(n749), .Z(n750) );
  XNOR U883 ( .A(b[125]), .B(n751), .Z(c[125]) );
  XNOR U884 ( .A(a[125]), .B(n752), .Z(n751) );
  IV U885 ( .A(n749), .Z(n752) );
  XOR U886 ( .A(n753), .B(n754), .Z(n749) );
  ANDN U887 ( .B(n755), .A(n756), .Z(n753) );
  XNOR U888 ( .A(b[124]), .B(n754), .Z(n755) );
  XNOR U889 ( .A(b[124]), .B(n756), .Z(c[124]) );
  XNOR U890 ( .A(a[124]), .B(n757), .Z(n756) );
  IV U891 ( .A(n754), .Z(n757) );
  XOR U892 ( .A(n758), .B(n759), .Z(n754) );
  ANDN U893 ( .B(n760), .A(n761), .Z(n758) );
  XNOR U894 ( .A(b[123]), .B(n759), .Z(n760) );
  XNOR U895 ( .A(b[123]), .B(n761), .Z(c[123]) );
  XNOR U896 ( .A(a[123]), .B(n762), .Z(n761) );
  IV U897 ( .A(n759), .Z(n762) );
  XOR U898 ( .A(n763), .B(n764), .Z(n759) );
  ANDN U899 ( .B(n765), .A(n766), .Z(n763) );
  XNOR U900 ( .A(b[122]), .B(n764), .Z(n765) );
  XNOR U901 ( .A(b[122]), .B(n766), .Z(c[122]) );
  XNOR U902 ( .A(a[122]), .B(n767), .Z(n766) );
  IV U903 ( .A(n764), .Z(n767) );
  XOR U904 ( .A(n768), .B(n769), .Z(n764) );
  ANDN U905 ( .B(n770), .A(n771), .Z(n768) );
  XNOR U906 ( .A(b[121]), .B(n769), .Z(n770) );
  XNOR U907 ( .A(b[121]), .B(n771), .Z(c[121]) );
  XNOR U908 ( .A(a[121]), .B(n772), .Z(n771) );
  IV U909 ( .A(n769), .Z(n772) );
  XOR U910 ( .A(n773), .B(n774), .Z(n769) );
  ANDN U911 ( .B(n775), .A(n776), .Z(n773) );
  XNOR U912 ( .A(b[120]), .B(n774), .Z(n775) );
  XNOR U913 ( .A(b[120]), .B(n776), .Z(c[120]) );
  XNOR U914 ( .A(a[120]), .B(n777), .Z(n776) );
  IV U915 ( .A(n774), .Z(n777) );
  XOR U916 ( .A(n778), .B(n779), .Z(n774) );
  ANDN U917 ( .B(n780), .A(n781), .Z(n778) );
  XNOR U918 ( .A(b[119]), .B(n779), .Z(n780) );
  XNOR U919 ( .A(b[11]), .B(n782), .Z(c[11]) );
  XNOR U920 ( .A(b[119]), .B(n781), .Z(c[119]) );
  XNOR U921 ( .A(a[119]), .B(n783), .Z(n781) );
  IV U922 ( .A(n779), .Z(n783) );
  XOR U923 ( .A(n784), .B(n785), .Z(n779) );
  ANDN U924 ( .B(n786), .A(n787), .Z(n784) );
  XNOR U925 ( .A(b[118]), .B(n785), .Z(n786) );
  XNOR U926 ( .A(b[118]), .B(n787), .Z(c[118]) );
  XNOR U927 ( .A(a[118]), .B(n788), .Z(n787) );
  IV U928 ( .A(n785), .Z(n788) );
  XOR U929 ( .A(n789), .B(n790), .Z(n785) );
  ANDN U930 ( .B(n791), .A(n792), .Z(n789) );
  XNOR U931 ( .A(b[117]), .B(n790), .Z(n791) );
  XNOR U932 ( .A(b[117]), .B(n792), .Z(c[117]) );
  XNOR U933 ( .A(a[117]), .B(n793), .Z(n792) );
  IV U934 ( .A(n790), .Z(n793) );
  XOR U935 ( .A(n794), .B(n795), .Z(n790) );
  ANDN U936 ( .B(n796), .A(n797), .Z(n794) );
  XNOR U937 ( .A(b[116]), .B(n795), .Z(n796) );
  XNOR U938 ( .A(b[116]), .B(n797), .Z(c[116]) );
  XNOR U939 ( .A(a[116]), .B(n798), .Z(n797) );
  IV U940 ( .A(n795), .Z(n798) );
  XOR U941 ( .A(n799), .B(n800), .Z(n795) );
  ANDN U942 ( .B(n801), .A(n802), .Z(n799) );
  XNOR U943 ( .A(b[115]), .B(n800), .Z(n801) );
  XNOR U944 ( .A(b[115]), .B(n802), .Z(c[115]) );
  XNOR U945 ( .A(a[115]), .B(n803), .Z(n802) );
  IV U946 ( .A(n800), .Z(n803) );
  XOR U947 ( .A(n804), .B(n805), .Z(n800) );
  ANDN U948 ( .B(n806), .A(n807), .Z(n804) );
  XNOR U949 ( .A(b[114]), .B(n805), .Z(n806) );
  XNOR U950 ( .A(b[114]), .B(n807), .Z(c[114]) );
  XNOR U951 ( .A(a[114]), .B(n808), .Z(n807) );
  IV U952 ( .A(n805), .Z(n808) );
  XOR U953 ( .A(n809), .B(n810), .Z(n805) );
  ANDN U954 ( .B(n811), .A(n812), .Z(n809) );
  XNOR U955 ( .A(b[113]), .B(n810), .Z(n811) );
  XNOR U956 ( .A(b[113]), .B(n812), .Z(c[113]) );
  XNOR U957 ( .A(a[113]), .B(n813), .Z(n812) );
  IV U958 ( .A(n810), .Z(n813) );
  XOR U959 ( .A(n814), .B(n815), .Z(n810) );
  ANDN U960 ( .B(n816), .A(n817), .Z(n814) );
  XNOR U961 ( .A(b[112]), .B(n815), .Z(n816) );
  XNOR U962 ( .A(b[112]), .B(n817), .Z(c[112]) );
  XNOR U963 ( .A(a[112]), .B(n818), .Z(n817) );
  IV U964 ( .A(n815), .Z(n818) );
  XOR U965 ( .A(n819), .B(n820), .Z(n815) );
  ANDN U966 ( .B(n821), .A(n822), .Z(n819) );
  XNOR U967 ( .A(b[111]), .B(n820), .Z(n821) );
  XNOR U968 ( .A(b[111]), .B(n822), .Z(c[111]) );
  XNOR U969 ( .A(a[111]), .B(n823), .Z(n822) );
  IV U970 ( .A(n820), .Z(n823) );
  XOR U971 ( .A(n824), .B(n825), .Z(n820) );
  ANDN U972 ( .B(n826), .A(n827), .Z(n824) );
  XNOR U973 ( .A(b[110]), .B(n825), .Z(n826) );
  XNOR U974 ( .A(b[110]), .B(n827), .Z(c[110]) );
  XNOR U975 ( .A(a[110]), .B(n828), .Z(n827) );
  IV U976 ( .A(n825), .Z(n828) );
  XOR U977 ( .A(n829), .B(n830), .Z(n825) );
  ANDN U978 ( .B(n831), .A(n832), .Z(n829) );
  XNOR U979 ( .A(b[109]), .B(n830), .Z(n831) );
  XNOR U980 ( .A(b[10]), .B(n833), .Z(c[10]) );
  XNOR U981 ( .A(b[109]), .B(n832), .Z(c[109]) );
  XNOR U982 ( .A(a[109]), .B(n834), .Z(n832) );
  IV U983 ( .A(n830), .Z(n834) );
  XOR U984 ( .A(n835), .B(n836), .Z(n830) );
  ANDN U985 ( .B(n837), .A(n838), .Z(n835) );
  XNOR U986 ( .A(b[108]), .B(n836), .Z(n837) );
  XNOR U987 ( .A(b[108]), .B(n838), .Z(c[108]) );
  XNOR U988 ( .A(a[108]), .B(n839), .Z(n838) );
  IV U989 ( .A(n836), .Z(n839) );
  XOR U990 ( .A(n840), .B(n841), .Z(n836) );
  ANDN U991 ( .B(n842), .A(n843), .Z(n840) );
  XNOR U992 ( .A(b[107]), .B(n841), .Z(n842) );
  XNOR U993 ( .A(b[107]), .B(n843), .Z(c[107]) );
  XNOR U994 ( .A(a[107]), .B(n844), .Z(n843) );
  IV U995 ( .A(n841), .Z(n844) );
  XOR U996 ( .A(n845), .B(n846), .Z(n841) );
  ANDN U997 ( .B(n847), .A(n848), .Z(n845) );
  XNOR U998 ( .A(b[106]), .B(n846), .Z(n847) );
  XNOR U999 ( .A(b[106]), .B(n848), .Z(c[106]) );
  XNOR U1000 ( .A(a[106]), .B(n849), .Z(n848) );
  IV U1001 ( .A(n846), .Z(n849) );
  XOR U1002 ( .A(n850), .B(n851), .Z(n846) );
  ANDN U1003 ( .B(n852), .A(n853), .Z(n850) );
  XNOR U1004 ( .A(b[105]), .B(n851), .Z(n852) );
  XNOR U1005 ( .A(b[105]), .B(n853), .Z(c[105]) );
  XNOR U1006 ( .A(a[105]), .B(n854), .Z(n853) );
  IV U1007 ( .A(n851), .Z(n854) );
  XOR U1008 ( .A(n855), .B(n856), .Z(n851) );
  ANDN U1009 ( .B(n857), .A(n858), .Z(n855) );
  XNOR U1010 ( .A(b[104]), .B(n856), .Z(n857) );
  XNOR U1011 ( .A(b[104]), .B(n858), .Z(c[104]) );
  XNOR U1012 ( .A(a[104]), .B(n859), .Z(n858) );
  IV U1013 ( .A(n856), .Z(n859) );
  XOR U1014 ( .A(n860), .B(n861), .Z(n856) );
  ANDN U1015 ( .B(n862), .A(n863), .Z(n860) );
  XNOR U1016 ( .A(b[103]), .B(n861), .Z(n862) );
  XNOR U1017 ( .A(b[103]), .B(n863), .Z(c[103]) );
  XNOR U1018 ( .A(a[103]), .B(n864), .Z(n863) );
  IV U1019 ( .A(n861), .Z(n864) );
  XOR U1020 ( .A(n865), .B(n866), .Z(n861) );
  ANDN U1021 ( .B(n867), .A(n868), .Z(n865) );
  XNOR U1022 ( .A(b[102]), .B(n866), .Z(n867) );
  XNOR U1023 ( .A(b[102]), .B(n868), .Z(c[102]) );
  XNOR U1024 ( .A(a[102]), .B(n869), .Z(n868) );
  IV U1025 ( .A(n866), .Z(n869) );
  XOR U1026 ( .A(n870), .B(n871), .Z(n866) );
  ANDN U1027 ( .B(n872), .A(n873), .Z(n870) );
  XNOR U1028 ( .A(b[101]), .B(n871), .Z(n872) );
  XNOR U1029 ( .A(b[101]), .B(n873), .Z(c[101]) );
  XNOR U1030 ( .A(a[101]), .B(n874), .Z(n873) );
  IV U1031 ( .A(n871), .Z(n874) );
  XOR U1032 ( .A(n875), .B(n876), .Z(n871) );
  ANDN U1033 ( .B(n877), .A(n878), .Z(n875) );
  XNOR U1034 ( .A(b[100]), .B(n876), .Z(n877) );
  XNOR U1035 ( .A(b[100]), .B(n878), .Z(c[100]) );
  XNOR U1036 ( .A(a[100]), .B(n879), .Z(n878) );
  IV U1037 ( .A(n876), .Z(n879) );
  XOR U1038 ( .A(n880), .B(n881), .Z(n876) );
  ANDN U1039 ( .B(n882), .A(n7), .Z(n880) );
  XNOR U1040 ( .A(a[99]), .B(n883), .Z(n7) );
  IV U1041 ( .A(n881), .Z(n883) );
  XNOR U1042 ( .A(b[99]), .B(n881), .Z(n882) );
  XOR U1043 ( .A(n884), .B(n885), .Z(n881) );
  ANDN U1044 ( .B(n886), .A(n8), .Z(n884) );
  XNOR U1045 ( .A(a[98]), .B(n887), .Z(n8) );
  IV U1046 ( .A(n885), .Z(n887) );
  XNOR U1047 ( .A(b[98]), .B(n885), .Z(n886) );
  XOR U1048 ( .A(n888), .B(n889), .Z(n885) );
  ANDN U1049 ( .B(n890), .A(n9), .Z(n888) );
  XNOR U1050 ( .A(a[97]), .B(n891), .Z(n9) );
  IV U1051 ( .A(n889), .Z(n891) );
  XNOR U1052 ( .A(b[97]), .B(n889), .Z(n890) );
  XOR U1053 ( .A(n892), .B(n893), .Z(n889) );
  ANDN U1054 ( .B(n894), .A(n10), .Z(n892) );
  XNOR U1055 ( .A(a[96]), .B(n895), .Z(n10) );
  IV U1056 ( .A(n893), .Z(n895) );
  XNOR U1057 ( .A(b[96]), .B(n893), .Z(n894) );
  XOR U1058 ( .A(n896), .B(n897), .Z(n893) );
  ANDN U1059 ( .B(n898), .A(n11), .Z(n896) );
  XNOR U1060 ( .A(a[95]), .B(n899), .Z(n11) );
  IV U1061 ( .A(n897), .Z(n899) );
  XNOR U1062 ( .A(b[95]), .B(n897), .Z(n898) );
  XOR U1063 ( .A(n900), .B(n901), .Z(n897) );
  ANDN U1064 ( .B(n902), .A(n12), .Z(n900) );
  XNOR U1065 ( .A(a[94]), .B(n903), .Z(n12) );
  IV U1066 ( .A(n901), .Z(n903) );
  XNOR U1067 ( .A(b[94]), .B(n901), .Z(n902) );
  XOR U1068 ( .A(n904), .B(n905), .Z(n901) );
  ANDN U1069 ( .B(n906), .A(n13), .Z(n904) );
  XNOR U1070 ( .A(a[93]), .B(n907), .Z(n13) );
  IV U1071 ( .A(n905), .Z(n907) );
  XNOR U1072 ( .A(b[93]), .B(n905), .Z(n906) );
  XOR U1073 ( .A(n908), .B(n909), .Z(n905) );
  ANDN U1074 ( .B(n910), .A(n14), .Z(n908) );
  XNOR U1075 ( .A(a[92]), .B(n911), .Z(n14) );
  IV U1076 ( .A(n909), .Z(n911) );
  XNOR U1077 ( .A(b[92]), .B(n909), .Z(n910) );
  XOR U1078 ( .A(n912), .B(n913), .Z(n909) );
  ANDN U1079 ( .B(n914), .A(n15), .Z(n912) );
  XNOR U1080 ( .A(a[91]), .B(n915), .Z(n15) );
  IV U1081 ( .A(n913), .Z(n915) );
  XNOR U1082 ( .A(b[91]), .B(n913), .Z(n914) );
  XOR U1083 ( .A(n916), .B(n917), .Z(n913) );
  ANDN U1084 ( .B(n918), .A(n16), .Z(n916) );
  XNOR U1085 ( .A(a[90]), .B(n919), .Z(n16) );
  IV U1086 ( .A(n917), .Z(n919) );
  XNOR U1087 ( .A(b[90]), .B(n917), .Z(n918) );
  XOR U1088 ( .A(n920), .B(n921), .Z(n917) );
  ANDN U1089 ( .B(n922), .A(n18), .Z(n920) );
  XNOR U1090 ( .A(a[89]), .B(n923), .Z(n18) );
  IV U1091 ( .A(n921), .Z(n923) );
  XNOR U1092 ( .A(b[89]), .B(n921), .Z(n922) );
  XOR U1093 ( .A(n924), .B(n925), .Z(n921) );
  ANDN U1094 ( .B(n926), .A(n19), .Z(n924) );
  XNOR U1095 ( .A(a[88]), .B(n927), .Z(n19) );
  IV U1096 ( .A(n925), .Z(n927) );
  XNOR U1097 ( .A(b[88]), .B(n925), .Z(n926) );
  XOR U1098 ( .A(n928), .B(n929), .Z(n925) );
  ANDN U1099 ( .B(n930), .A(n20), .Z(n928) );
  XNOR U1100 ( .A(a[87]), .B(n931), .Z(n20) );
  IV U1101 ( .A(n929), .Z(n931) );
  XNOR U1102 ( .A(b[87]), .B(n929), .Z(n930) );
  XOR U1103 ( .A(n932), .B(n933), .Z(n929) );
  ANDN U1104 ( .B(n934), .A(n21), .Z(n932) );
  XNOR U1105 ( .A(a[86]), .B(n935), .Z(n21) );
  IV U1106 ( .A(n933), .Z(n935) );
  XNOR U1107 ( .A(b[86]), .B(n933), .Z(n934) );
  XOR U1108 ( .A(n936), .B(n937), .Z(n933) );
  ANDN U1109 ( .B(n938), .A(n22), .Z(n936) );
  XNOR U1110 ( .A(a[85]), .B(n939), .Z(n22) );
  IV U1111 ( .A(n937), .Z(n939) );
  XNOR U1112 ( .A(b[85]), .B(n937), .Z(n938) );
  XOR U1113 ( .A(n940), .B(n941), .Z(n937) );
  ANDN U1114 ( .B(n942), .A(n23), .Z(n940) );
  XNOR U1115 ( .A(a[84]), .B(n943), .Z(n23) );
  IV U1116 ( .A(n941), .Z(n943) );
  XNOR U1117 ( .A(b[84]), .B(n941), .Z(n942) );
  XOR U1118 ( .A(n944), .B(n945), .Z(n941) );
  ANDN U1119 ( .B(n946), .A(n24), .Z(n944) );
  XNOR U1120 ( .A(a[83]), .B(n947), .Z(n24) );
  IV U1121 ( .A(n945), .Z(n947) );
  XNOR U1122 ( .A(b[83]), .B(n945), .Z(n946) );
  XOR U1123 ( .A(n948), .B(n949), .Z(n945) );
  ANDN U1124 ( .B(n950), .A(n25), .Z(n948) );
  XNOR U1125 ( .A(a[82]), .B(n951), .Z(n25) );
  IV U1126 ( .A(n949), .Z(n951) );
  XNOR U1127 ( .A(b[82]), .B(n949), .Z(n950) );
  XOR U1128 ( .A(n952), .B(n953), .Z(n949) );
  ANDN U1129 ( .B(n954), .A(n26), .Z(n952) );
  XNOR U1130 ( .A(a[81]), .B(n955), .Z(n26) );
  IV U1131 ( .A(n953), .Z(n955) );
  XNOR U1132 ( .A(b[81]), .B(n953), .Z(n954) );
  XOR U1133 ( .A(n956), .B(n957), .Z(n953) );
  ANDN U1134 ( .B(n958), .A(n27), .Z(n956) );
  XNOR U1135 ( .A(a[80]), .B(n959), .Z(n27) );
  IV U1136 ( .A(n957), .Z(n959) );
  XNOR U1137 ( .A(b[80]), .B(n957), .Z(n958) );
  XOR U1138 ( .A(n960), .B(n961), .Z(n957) );
  ANDN U1139 ( .B(n962), .A(n29), .Z(n960) );
  XNOR U1140 ( .A(a[79]), .B(n963), .Z(n29) );
  IV U1141 ( .A(n961), .Z(n963) );
  XNOR U1142 ( .A(b[79]), .B(n961), .Z(n962) );
  XOR U1143 ( .A(n964), .B(n965), .Z(n961) );
  ANDN U1144 ( .B(n966), .A(n30), .Z(n964) );
  XNOR U1145 ( .A(a[78]), .B(n967), .Z(n30) );
  IV U1146 ( .A(n965), .Z(n967) );
  XNOR U1147 ( .A(b[78]), .B(n965), .Z(n966) );
  XOR U1148 ( .A(n968), .B(n969), .Z(n965) );
  ANDN U1149 ( .B(n970), .A(n31), .Z(n968) );
  XNOR U1150 ( .A(a[77]), .B(n971), .Z(n31) );
  IV U1151 ( .A(n969), .Z(n971) );
  XNOR U1152 ( .A(b[77]), .B(n969), .Z(n970) );
  XOR U1153 ( .A(n972), .B(n973), .Z(n969) );
  ANDN U1154 ( .B(n974), .A(n32), .Z(n972) );
  XNOR U1155 ( .A(a[76]), .B(n975), .Z(n32) );
  IV U1156 ( .A(n973), .Z(n975) );
  XNOR U1157 ( .A(b[76]), .B(n973), .Z(n974) );
  XOR U1158 ( .A(n976), .B(n977), .Z(n973) );
  ANDN U1159 ( .B(n978), .A(n33), .Z(n976) );
  XNOR U1160 ( .A(a[75]), .B(n979), .Z(n33) );
  IV U1161 ( .A(n977), .Z(n979) );
  XNOR U1162 ( .A(b[75]), .B(n977), .Z(n978) );
  XOR U1163 ( .A(n980), .B(n981), .Z(n977) );
  ANDN U1164 ( .B(n982), .A(n34), .Z(n980) );
  XNOR U1165 ( .A(a[74]), .B(n983), .Z(n34) );
  IV U1166 ( .A(n981), .Z(n983) );
  XNOR U1167 ( .A(b[74]), .B(n981), .Z(n982) );
  XOR U1168 ( .A(n984), .B(n985), .Z(n981) );
  ANDN U1169 ( .B(n986), .A(n35), .Z(n984) );
  XNOR U1170 ( .A(a[73]), .B(n987), .Z(n35) );
  IV U1171 ( .A(n985), .Z(n987) );
  XNOR U1172 ( .A(b[73]), .B(n985), .Z(n986) );
  XOR U1173 ( .A(n988), .B(n989), .Z(n985) );
  ANDN U1174 ( .B(n990), .A(n36), .Z(n988) );
  XNOR U1175 ( .A(a[72]), .B(n991), .Z(n36) );
  IV U1176 ( .A(n989), .Z(n991) );
  XNOR U1177 ( .A(b[72]), .B(n989), .Z(n990) );
  XOR U1178 ( .A(n992), .B(n993), .Z(n989) );
  ANDN U1179 ( .B(n994), .A(n37), .Z(n992) );
  XNOR U1180 ( .A(a[71]), .B(n995), .Z(n37) );
  IV U1181 ( .A(n993), .Z(n995) );
  XNOR U1182 ( .A(b[71]), .B(n993), .Z(n994) );
  XOR U1183 ( .A(n996), .B(n997), .Z(n993) );
  ANDN U1184 ( .B(n998), .A(n38), .Z(n996) );
  XNOR U1185 ( .A(a[70]), .B(n999), .Z(n38) );
  IV U1186 ( .A(n997), .Z(n999) );
  XNOR U1187 ( .A(b[70]), .B(n997), .Z(n998) );
  XOR U1188 ( .A(n1000), .B(n1001), .Z(n997) );
  ANDN U1189 ( .B(n1002), .A(n40), .Z(n1000) );
  XNOR U1190 ( .A(a[69]), .B(n1003), .Z(n40) );
  IV U1191 ( .A(n1001), .Z(n1003) );
  XNOR U1192 ( .A(b[69]), .B(n1001), .Z(n1002) );
  XOR U1193 ( .A(n1004), .B(n1005), .Z(n1001) );
  ANDN U1194 ( .B(n1006), .A(n41), .Z(n1004) );
  XNOR U1195 ( .A(a[68]), .B(n1007), .Z(n41) );
  IV U1196 ( .A(n1005), .Z(n1007) );
  XNOR U1197 ( .A(b[68]), .B(n1005), .Z(n1006) );
  XOR U1198 ( .A(n1008), .B(n1009), .Z(n1005) );
  ANDN U1199 ( .B(n1010), .A(n42), .Z(n1008) );
  XNOR U1200 ( .A(a[67]), .B(n1011), .Z(n42) );
  IV U1201 ( .A(n1009), .Z(n1011) );
  XNOR U1202 ( .A(b[67]), .B(n1009), .Z(n1010) );
  XOR U1203 ( .A(n1012), .B(n1013), .Z(n1009) );
  ANDN U1204 ( .B(n1014), .A(n43), .Z(n1012) );
  XNOR U1205 ( .A(a[66]), .B(n1015), .Z(n43) );
  IV U1206 ( .A(n1013), .Z(n1015) );
  XNOR U1207 ( .A(b[66]), .B(n1013), .Z(n1014) );
  XOR U1208 ( .A(n1016), .B(n1017), .Z(n1013) );
  ANDN U1209 ( .B(n1018), .A(n44), .Z(n1016) );
  XNOR U1210 ( .A(a[65]), .B(n1019), .Z(n44) );
  IV U1211 ( .A(n1017), .Z(n1019) );
  XNOR U1212 ( .A(b[65]), .B(n1017), .Z(n1018) );
  XOR U1213 ( .A(n1020), .B(n1021), .Z(n1017) );
  ANDN U1214 ( .B(n1022), .A(n45), .Z(n1020) );
  XNOR U1215 ( .A(a[64]), .B(n1023), .Z(n45) );
  IV U1216 ( .A(n1021), .Z(n1023) );
  XNOR U1217 ( .A(b[64]), .B(n1021), .Z(n1022) );
  XOR U1218 ( .A(n1024), .B(n1025), .Z(n1021) );
  ANDN U1219 ( .B(n1026), .A(n46), .Z(n1024) );
  XNOR U1220 ( .A(a[63]), .B(n1027), .Z(n46) );
  IV U1221 ( .A(n1025), .Z(n1027) );
  XNOR U1222 ( .A(b[63]), .B(n1025), .Z(n1026) );
  XOR U1223 ( .A(n1028), .B(n1029), .Z(n1025) );
  ANDN U1224 ( .B(n1030), .A(n47), .Z(n1028) );
  XNOR U1225 ( .A(a[62]), .B(n1031), .Z(n47) );
  IV U1226 ( .A(n1029), .Z(n1031) );
  XNOR U1227 ( .A(b[62]), .B(n1029), .Z(n1030) );
  XOR U1228 ( .A(n1032), .B(n1033), .Z(n1029) );
  ANDN U1229 ( .B(n1034), .A(n48), .Z(n1032) );
  XNOR U1230 ( .A(a[61]), .B(n1035), .Z(n48) );
  IV U1231 ( .A(n1033), .Z(n1035) );
  XNOR U1232 ( .A(b[61]), .B(n1033), .Z(n1034) );
  XOR U1233 ( .A(n1036), .B(n1037), .Z(n1033) );
  ANDN U1234 ( .B(n1038), .A(n49), .Z(n1036) );
  XNOR U1235 ( .A(a[60]), .B(n1039), .Z(n49) );
  IV U1236 ( .A(n1037), .Z(n1039) );
  XNOR U1237 ( .A(b[60]), .B(n1037), .Z(n1038) );
  XOR U1238 ( .A(n1040), .B(n1041), .Z(n1037) );
  ANDN U1239 ( .B(n1042), .A(n51), .Z(n1040) );
  XNOR U1240 ( .A(a[59]), .B(n1043), .Z(n51) );
  IV U1241 ( .A(n1041), .Z(n1043) );
  XNOR U1242 ( .A(b[59]), .B(n1041), .Z(n1042) );
  XOR U1243 ( .A(n1044), .B(n1045), .Z(n1041) );
  ANDN U1244 ( .B(n1046), .A(n52), .Z(n1044) );
  XNOR U1245 ( .A(a[58]), .B(n1047), .Z(n52) );
  IV U1246 ( .A(n1045), .Z(n1047) );
  XNOR U1247 ( .A(b[58]), .B(n1045), .Z(n1046) );
  XOR U1248 ( .A(n1048), .B(n1049), .Z(n1045) );
  ANDN U1249 ( .B(n1050), .A(n53), .Z(n1048) );
  XNOR U1250 ( .A(a[57]), .B(n1051), .Z(n53) );
  IV U1251 ( .A(n1049), .Z(n1051) );
  XNOR U1252 ( .A(b[57]), .B(n1049), .Z(n1050) );
  XOR U1253 ( .A(n1052), .B(n1053), .Z(n1049) );
  ANDN U1254 ( .B(n1054), .A(n54), .Z(n1052) );
  XNOR U1255 ( .A(a[56]), .B(n1055), .Z(n54) );
  IV U1256 ( .A(n1053), .Z(n1055) );
  XNOR U1257 ( .A(b[56]), .B(n1053), .Z(n1054) );
  XOR U1258 ( .A(n1056), .B(n1057), .Z(n1053) );
  ANDN U1259 ( .B(n1058), .A(n55), .Z(n1056) );
  XNOR U1260 ( .A(a[55]), .B(n1059), .Z(n55) );
  IV U1261 ( .A(n1057), .Z(n1059) );
  XNOR U1262 ( .A(b[55]), .B(n1057), .Z(n1058) );
  XOR U1263 ( .A(n1060), .B(n1061), .Z(n1057) );
  ANDN U1264 ( .B(n1062), .A(n56), .Z(n1060) );
  XNOR U1265 ( .A(a[54]), .B(n1063), .Z(n56) );
  IV U1266 ( .A(n1061), .Z(n1063) );
  XNOR U1267 ( .A(b[54]), .B(n1061), .Z(n1062) );
  XOR U1268 ( .A(n1064), .B(n1065), .Z(n1061) );
  ANDN U1269 ( .B(n1066), .A(n57), .Z(n1064) );
  XNOR U1270 ( .A(a[53]), .B(n1067), .Z(n57) );
  IV U1271 ( .A(n1065), .Z(n1067) );
  XNOR U1272 ( .A(b[53]), .B(n1065), .Z(n1066) );
  XOR U1273 ( .A(n1068), .B(n1069), .Z(n1065) );
  ANDN U1274 ( .B(n1070), .A(n58), .Z(n1068) );
  XNOR U1275 ( .A(a[52]), .B(n1071), .Z(n58) );
  IV U1276 ( .A(n1069), .Z(n1071) );
  XNOR U1277 ( .A(b[52]), .B(n1069), .Z(n1070) );
  XOR U1278 ( .A(n1072), .B(n1073), .Z(n1069) );
  ANDN U1279 ( .B(n1074), .A(n59), .Z(n1072) );
  XNOR U1280 ( .A(a[51]), .B(n1075), .Z(n59) );
  IV U1281 ( .A(n1073), .Z(n1075) );
  XNOR U1282 ( .A(b[51]), .B(n1073), .Z(n1074) );
  XOR U1283 ( .A(n1076), .B(n1077), .Z(n1073) );
  ANDN U1284 ( .B(n1078), .A(n60), .Z(n1076) );
  XNOR U1285 ( .A(a[50]), .B(n1079), .Z(n60) );
  IV U1286 ( .A(n1077), .Z(n1079) );
  XNOR U1287 ( .A(b[50]), .B(n1077), .Z(n1078) );
  XOR U1288 ( .A(n1080), .B(n1081), .Z(n1077) );
  ANDN U1289 ( .B(n1082), .A(n62), .Z(n1080) );
  XNOR U1290 ( .A(a[49]), .B(n1083), .Z(n62) );
  IV U1291 ( .A(n1081), .Z(n1083) );
  XNOR U1292 ( .A(b[49]), .B(n1081), .Z(n1082) );
  XOR U1293 ( .A(n1084), .B(n1085), .Z(n1081) );
  ANDN U1294 ( .B(n1086), .A(n63), .Z(n1084) );
  XNOR U1295 ( .A(a[48]), .B(n1087), .Z(n63) );
  IV U1296 ( .A(n1085), .Z(n1087) );
  XNOR U1297 ( .A(b[48]), .B(n1085), .Z(n1086) );
  XOR U1298 ( .A(n1088), .B(n1089), .Z(n1085) );
  ANDN U1299 ( .B(n1090), .A(n64), .Z(n1088) );
  XNOR U1300 ( .A(a[47]), .B(n1091), .Z(n64) );
  IV U1301 ( .A(n1089), .Z(n1091) );
  XNOR U1302 ( .A(b[47]), .B(n1089), .Z(n1090) );
  XOR U1303 ( .A(n1092), .B(n1093), .Z(n1089) );
  ANDN U1304 ( .B(n1094), .A(n65), .Z(n1092) );
  XNOR U1305 ( .A(a[46]), .B(n1095), .Z(n65) );
  IV U1306 ( .A(n1093), .Z(n1095) );
  XNOR U1307 ( .A(b[46]), .B(n1093), .Z(n1094) );
  XOR U1308 ( .A(n1096), .B(n1097), .Z(n1093) );
  ANDN U1309 ( .B(n1098), .A(n66), .Z(n1096) );
  XNOR U1310 ( .A(a[45]), .B(n1099), .Z(n66) );
  IV U1311 ( .A(n1097), .Z(n1099) );
  XNOR U1312 ( .A(b[45]), .B(n1097), .Z(n1098) );
  XOR U1313 ( .A(n1100), .B(n1101), .Z(n1097) );
  ANDN U1314 ( .B(n1102), .A(n67), .Z(n1100) );
  XNOR U1315 ( .A(a[44]), .B(n1103), .Z(n67) );
  IV U1316 ( .A(n1101), .Z(n1103) );
  XNOR U1317 ( .A(b[44]), .B(n1101), .Z(n1102) );
  XOR U1318 ( .A(n1104), .B(n1105), .Z(n1101) );
  ANDN U1319 ( .B(n1106), .A(n68), .Z(n1104) );
  XNOR U1320 ( .A(a[43]), .B(n1107), .Z(n68) );
  IV U1321 ( .A(n1105), .Z(n1107) );
  XNOR U1322 ( .A(b[43]), .B(n1105), .Z(n1106) );
  XOR U1323 ( .A(n1108), .B(n1109), .Z(n1105) );
  ANDN U1324 ( .B(n1110), .A(n69), .Z(n1108) );
  XNOR U1325 ( .A(a[42]), .B(n1111), .Z(n69) );
  IV U1326 ( .A(n1109), .Z(n1111) );
  XNOR U1327 ( .A(b[42]), .B(n1109), .Z(n1110) );
  XOR U1328 ( .A(n1112), .B(n1113), .Z(n1109) );
  ANDN U1329 ( .B(n1114), .A(n70), .Z(n1112) );
  XNOR U1330 ( .A(a[41]), .B(n1115), .Z(n70) );
  IV U1331 ( .A(n1113), .Z(n1115) );
  XNOR U1332 ( .A(b[41]), .B(n1113), .Z(n1114) );
  XOR U1333 ( .A(n1116), .B(n1117), .Z(n1113) );
  ANDN U1334 ( .B(n1118), .A(n71), .Z(n1116) );
  XNOR U1335 ( .A(a[40]), .B(n1119), .Z(n71) );
  IV U1336 ( .A(n1117), .Z(n1119) );
  XNOR U1337 ( .A(b[40]), .B(n1117), .Z(n1118) );
  XOR U1338 ( .A(n1120), .B(n1121), .Z(n1117) );
  ANDN U1339 ( .B(n1122), .A(n73), .Z(n1120) );
  XNOR U1340 ( .A(a[39]), .B(n1123), .Z(n73) );
  IV U1341 ( .A(n1121), .Z(n1123) );
  XNOR U1342 ( .A(b[39]), .B(n1121), .Z(n1122) );
  XOR U1343 ( .A(n1124), .B(n1125), .Z(n1121) );
  ANDN U1344 ( .B(n1126), .A(n74), .Z(n1124) );
  XNOR U1345 ( .A(a[38]), .B(n1127), .Z(n74) );
  IV U1346 ( .A(n1125), .Z(n1127) );
  XNOR U1347 ( .A(b[38]), .B(n1125), .Z(n1126) );
  XOR U1348 ( .A(n1128), .B(n1129), .Z(n1125) );
  ANDN U1349 ( .B(n1130), .A(n75), .Z(n1128) );
  XNOR U1350 ( .A(a[37]), .B(n1131), .Z(n75) );
  IV U1351 ( .A(n1129), .Z(n1131) );
  XNOR U1352 ( .A(b[37]), .B(n1129), .Z(n1130) );
  XOR U1353 ( .A(n1132), .B(n1133), .Z(n1129) );
  ANDN U1354 ( .B(n1134), .A(n76), .Z(n1132) );
  XNOR U1355 ( .A(a[36]), .B(n1135), .Z(n76) );
  IV U1356 ( .A(n1133), .Z(n1135) );
  XNOR U1357 ( .A(b[36]), .B(n1133), .Z(n1134) );
  XOR U1358 ( .A(n1136), .B(n1137), .Z(n1133) );
  ANDN U1359 ( .B(n1138), .A(n77), .Z(n1136) );
  XNOR U1360 ( .A(a[35]), .B(n1139), .Z(n77) );
  IV U1361 ( .A(n1137), .Z(n1139) );
  XNOR U1362 ( .A(b[35]), .B(n1137), .Z(n1138) );
  XOR U1363 ( .A(n1140), .B(n1141), .Z(n1137) );
  ANDN U1364 ( .B(n1142), .A(n78), .Z(n1140) );
  XNOR U1365 ( .A(a[34]), .B(n1143), .Z(n78) );
  IV U1366 ( .A(n1141), .Z(n1143) );
  XNOR U1367 ( .A(b[34]), .B(n1141), .Z(n1142) );
  XOR U1368 ( .A(n1144), .B(n1145), .Z(n1141) );
  ANDN U1369 ( .B(n1146), .A(n79), .Z(n1144) );
  XNOR U1370 ( .A(a[33]), .B(n1147), .Z(n79) );
  IV U1371 ( .A(n1145), .Z(n1147) );
  XNOR U1372 ( .A(b[33]), .B(n1145), .Z(n1146) );
  XOR U1373 ( .A(n1148), .B(n1149), .Z(n1145) );
  ANDN U1374 ( .B(n1150), .A(n80), .Z(n1148) );
  XNOR U1375 ( .A(a[32]), .B(n1151), .Z(n80) );
  IV U1376 ( .A(n1149), .Z(n1151) );
  XNOR U1377 ( .A(b[32]), .B(n1149), .Z(n1150) );
  XOR U1378 ( .A(n1152), .B(n1153), .Z(n1149) );
  ANDN U1379 ( .B(n1154), .A(n81), .Z(n1152) );
  XNOR U1380 ( .A(a[31]), .B(n1155), .Z(n81) );
  IV U1381 ( .A(n1153), .Z(n1155) );
  XNOR U1382 ( .A(b[31]), .B(n1153), .Z(n1154) );
  XOR U1383 ( .A(n1156), .B(n1157), .Z(n1153) );
  ANDN U1384 ( .B(n1158), .A(n82), .Z(n1156) );
  XNOR U1385 ( .A(a[30]), .B(n1159), .Z(n82) );
  IV U1386 ( .A(n1157), .Z(n1159) );
  XNOR U1387 ( .A(b[30]), .B(n1157), .Z(n1158) );
  XOR U1388 ( .A(n1160), .B(n1161), .Z(n1157) );
  ANDN U1389 ( .B(n1162), .A(n84), .Z(n1160) );
  XNOR U1390 ( .A(a[29]), .B(n1163), .Z(n84) );
  IV U1391 ( .A(n1161), .Z(n1163) );
  XNOR U1392 ( .A(b[29]), .B(n1161), .Z(n1162) );
  XOR U1393 ( .A(n1164), .B(n1165), .Z(n1161) );
  ANDN U1394 ( .B(n1166), .A(n85), .Z(n1164) );
  XNOR U1395 ( .A(a[28]), .B(n1167), .Z(n85) );
  IV U1396 ( .A(n1165), .Z(n1167) );
  XNOR U1397 ( .A(b[28]), .B(n1165), .Z(n1166) );
  XOR U1398 ( .A(n1168), .B(n1169), .Z(n1165) );
  ANDN U1399 ( .B(n1170), .A(n86), .Z(n1168) );
  XNOR U1400 ( .A(a[27]), .B(n1171), .Z(n86) );
  IV U1401 ( .A(n1169), .Z(n1171) );
  XNOR U1402 ( .A(b[27]), .B(n1169), .Z(n1170) );
  XOR U1403 ( .A(n1172), .B(n1173), .Z(n1169) );
  ANDN U1404 ( .B(n1174), .A(n87), .Z(n1172) );
  XNOR U1405 ( .A(a[26]), .B(n1175), .Z(n87) );
  IV U1406 ( .A(n1173), .Z(n1175) );
  XNOR U1407 ( .A(b[26]), .B(n1173), .Z(n1174) );
  XOR U1408 ( .A(n1176), .B(n1177), .Z(n1173) );
  ANDN U1409 ( .B(n1178), .A(n88), .Z(n1176) );
  XNOR U1410 ( .A(a[25]), .B(n1179), .Z(n88) );
  IV U1411 ( .A(n1177), .Z(n1179) );
  XNOR U1412 ( .A(b[25]), .B(n1177), .Z(n1178) );
  XOR U1413 ( .A(n1180), .B(n1181), .Z(n1177) );
  ANDN U1414 ( .B(n1182), .A(n118), .Z(n1180) );
  XNOR U1415 ( .A(a[24]), .B(n1183), .Z(n118) );
  IV U1416 ( .A(n1181), .Z(n1183) );
  XNOR U1417 ( .A(b[24]), .B(n1181), .Z(n1182) );
  XOR U1418 ( .A(n1184), .B(n1185), .Z(n1181) );
  ANDN U1419 ( .B(n1186), .A(n169), .Z(n1184) );
  XNOR U1420 ( .A(a[23]), .B(n1187), .Z(n169) );
  IV U1421 ( .A(n1185), .Z(n1187) );
  XNOR U1422 ( .A(b[23]), .B(n1185), .Z(n1186) );
  XOR U1423 ( .A(n1188), .B(n1189), .Z(n1185) );
  ANDN U1424 ( .B(n1190), .A(n220), .Z(n1188) );
  XNOR U1425 ( .A(a[22]), .B(n1191), .Z(n220) );
  IV U1426 ( .A(n1189), .Z(n1191) );
  XNOR U1427 ( .A(b[22]), .B(n1189), .Z(n1190) );
  XOR U1428 ( .A(n1192), .B(n1193), .Z(n1189) );
  ANDN U1429 ( .B(n1194), .A(n271), .Z(n1192) );
  XNOR U1430 ( .A(a[21]), .B(n1195), .Z(n271) );
  IV U1431 ( .A(n1193), .Z(n1195) );
  XNOR U1432 ( .A(b[21]), .B(n1193), .Z(n1194) );
  XOR U1433 ( .A(n1196), .B(n1197), .Z(n1193) );
  ANDN U1434 ( .B(n1198), .A(n322), .Z(n1196) );
  XNOR U1435 ( .A(a[20]), .B(n1199), .Z(n322) );
  IV U1436 ( .A(n1197), .Z(n1199) );
  XNOR U1437 ( .A(b[20]), .B(n1197), .Z(n1198) );
  XOR U1438 ( .A(n1200), .B(n1201), .Z(n1197) );
  ANDN U1439 ( .B(n1202), .A(n374), .Z(n1200) );
  XNOR U1440 ( .A(a[19]), .B(n1203), .Z(n374) );
  IV U1441 ( .A(n1201), .Z(n1203) );
  XNOR U1442 ( .A(b[19]), .B(n1201), .Z(n1202) );
  XOR U1443 ( .A(n1204), .B(n1205), .Z(n1201) );
  ANDN U1444 ( .B(n1206), .A(n425), .Z(n1204) );
  XNOR U1445 ( .A(a[18]), .B(n1207), .Z(n425) );
  IV U1446 ( .A(n1205), .Z(n1207) );
  XNOR U1447 ( .A(b[18]), .B(n1205), .Z(n1206) );
  XOR U1448 ( .A(n1208), .B(n1209), .Z(n1205) );
  ANDN U1449 ( .B(n1210), .A(n476), .Z(n1208) );
  XNOR U1450 ( .A(a[17]), .B(n1211), .Z(n476) );
  IV U1451 ( .A(n1209), .Z(n1211) );
  XNOR U1452 ( .A(b[17]), .B(n1209), .Z(n1210) );
  XOR U1453 ( .A(n1212), .B(n1213), .Z(n1209) );
  ANDN U1454 ( .B(n1214), .A(n527), .Z(n1212) );
  XNOR U1455 ( .A(a[16]), .B(n1215), .Z(n527) );
  IV U1456 ( .A(n1213), .Z(n1215) );
  XNOR U1457 ( .A(b[16]), .B(n1213), .Z(n1214) );
  XOR U1458 ( .A(n1216), .B(n1217), .Z(n1213) );
  ANDN U1459 ( .B(n1218), .A(n578), .Z(n1216) );
  XNOR U1460 ( .A(a[15]), .B(n1219), .Z(n578) );
  IV U1461 ( .A(n1217), .Z(n1219) );
  XNOR U1462 ( .A(b[15]), .B(n1217), .Z(n1218) );
  XOR U1463 ( .A(n1220), .B(n1221), .Z(n1217) );
  ANDN U1464 ( .B(n1222), .A(n629), .Z(n1220) );
  XNOR U1465 ( .A(a[14]), .B(n1223), .Z(n629) );
  IV U1466 ( .A(n1221), .Z(n1223) );
  XNOR U1467 ( .A(b[14]), .B(n1221), .Z(n1222) );
  XOR U1468 ( .A(n1224), .B(n1225), .Z(n1221) );
  ANDN U1469 ( .B(n1226), .A(n680), .Z(n1224) );
  XNOR U1470 ( .A(a[13]), .B(n1227), .Z(n680) );
  IV U1471 ( .A(n1225), .Z(n1227) );
  XNOR U1472 ( .A(b[13]), .B(n1225), .Z(n1226) );
  XOR U1473 ( .A(n1228), .B(n1229), .Z(n1225) );
  ANDN U1474 ( .B(n1230), .A(n731), .Z(n1228) );
  XNOR U1475 ( .A(a[12]), .B(n1231), .Z(n731) );
  IV U1476 ( .A(n1229), .Z(n1231) );
  XNOR U1477 ( .A(b[12]), .B(n1229), .Z(n1230) );
  XOR U1478 ( .A(n1232), .B(n1233), .Z(n1229) );
  ANDN U1479 ( .B(n1234), .A(n782), .Z(n1232) );
  XNOR U1480 ( .A(a[11]), .B(n1235), .Z(n782) );
  IV U1481 ( .A(n1233), .Z(n1235) );
  XNOR U1482 ( .A(b[11]), .B(n1233), .Z(n1234) );
  XOR U1483 ( .A(n1236), .B(n1237), .Z(n1233) );
  ANDN U1484 ( .B(n1238), .A(n833), .Z(n1236) );
  XNOR U1485 ( .A(a[10]), .B(n1239), .Z(n833) );
  IV U1486 ( .A(n1237), .Z(n1239) );
  XNOR U1487 ( .A(b[10]), .B(n1237), .Z(n1238) );
  XOR U1488 ( .A(n1240), .B(n1241), .Z(n1237) );
  ANDN U1489 ( .B(n1242), .A(n6), .Z(n1240) );
  XNOR U1490 ( .A(a[9]), .B(n1243), .Z(n6) );
  IV U1491 ( .A(n1241), .Z(n1243) );
  XNOR U1492 ( .A(b[9]), .B(n1241), .Z(n1242) );
  XOR U1493 ( .A(n1244), .B(n1245), .Z(n1241) );
  ANDN U1494 ( .B(n1246), .A(n17), .Z(n1244) );
  XNOR U1495 ( .A(a[8]), .B(n1247), .Z(n17) );
  IV U1496 ( .A(n1245), .Z(n1247) );
  XNOR U1497 ( .A(b[8]), .B(n1245), .Z(n1246) );
  XOR U1498 ( .A(n1248), .B(n1249), .Z(n1245) );
  ANDN U1499 ( .B(n1250), .A(n28), .Z(n1248) );
  XNOR U1500 ( .A(a[7]), .B(n1251), .Z(n28) );
  IV U1501 ( .A(n1249), .Z(n1251) );
  XNOR U1502 ( .A(b[7]), .B(n1249), .Z(n1250) );
  XOR U1503 ( .A(n1252), .B(n1253), .Z(n1249) );
  ANDN U1504 ( .B(n1254), .A(n39), .Z(n1252) );
  XNOR U1505 ( .A(a[6]), .B(n1255), .Z(n39) );
  IV U1506 ( .A(n1253), .Z(n1255) );
  XNOR U1507 ( .A(b[6]), .B(n1253), .Z(n1254) );
  XOR U1508 ( .A(n1256), .B(n1257), .Z(n1253) );
  ANDN U1509 ( .B(n1258), .A(n50), .Z(n1256) );
  XNOR U1510 ( .A(a[5]), .B(n1259), .Z(n50) );
  IV U1511 ( .A(n1257), .Z(n1259) );
  XNOR U1512 ( .A(b[5]), .B(n1257), .Z(n1258) );
  XOR U1513 ( .A(n1260), .B(n1261), .Z(n1257) );
  ANDN U1514 ( .B(n1262), .A(n61), .Z(n1260) );
  XNOR U1515 ( .A(a[4]), .B(n1263), .Z(n61) );
  IV U1516 ( .A(n1261), .Z(n1263) );
  XNOR U1517 ( .A(b[4]), .B(n1261), .Z(n1262) );
  XOR U1518 ( .A(n1264), .B(n1265), .Z(n1261) );
  ANDN U1519 ( .B(n1266), .A(n72), .Z(n1264) );
  XNOR U1520 ( .A(a[3]), .B(n1267), .Z(n72) );
  IV U1521 ( .A(n1265), .Z(n1267) );
  XNOR U1522 ( .A(b[3]), .B(n1265), .Z(n1266) );
  XOR U1523 ( .A(n1268), .B(n1269), .Z(n1265) );
  ANDN U1524 ( .B(n1270), .A(n83), .Z(n1268) );
  XNOR U1525 ( .A(a[2]), .B(n1271), .Z(n83) );
  IV U1526 ( .A(n1269), .Z(n1271) );
  XNOR U1527 ( .A(b[2]), .B(n1269), .Z(n1270) );
  XOR U1528 ( .A(n1272), .B(n1273), .Z(n1269) );
  ANDN U1529 ( .B(n1274), .A(n373), .Z(n1272) );
  XNOR U1530 ( .A(a[1]), .B(n1275), .Z(n373) );
  IV U1531 ( .A(n1273), .Z(n1275) );
  XNOR U1532 ( .A(b[1]), .B(n1273), .Z(n1274) );
  XOR U1533 ( .A(carry_on), .B(n1276), .Z(n1273) );
  NANDN U1534 ( .A(n1277), .B(n1278), .Z(n1276) );
  XOR U1535 ( .A(carry_on), .B(b[0]), .Z(n1278) );
  XNOR U1536 ( .A(b[0]), .B(n1277), .Z(c[0]) );
  XNOR U1537 ( .A(a[0]), .B(carry_on), .Z(n1277) );
endmodule

