
module sum_N128_CC4 ( clk, rst, a, b, c );
  input [31:0] a;
  input [31:0] b;
  output [31:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[0]), .B(b[0]), .Z(n1) );
  XOR U4 ( .A(n1), .B(carry_on), .Z(c[0]) );
  XOR U5 ( .A(a[1]), .B(b[1]), .Z(n4) );
  NAND U6 ( .A(b[0]), .B(a[0]), .Z(n3) );
  NAND U7 ( .A(carry_on), .B(n1), .Z(n2) );
  AND U8 ( .A(n3), .B(n2), .Z(n5) );
  XNOR U9 ( .A(n4), .B(n5), .Z(c[1]) );
  XOR U10 ( .A(a[2]), .B(b[2]), .Z(n8) );
  NAND U11 ( .A(b[1]), .B(a[1]), .Z(n7) );
  NANDN U12 ( .A(n5), .B(n4), .Z(n6) );
  AND U13 ( .A(n7), .B(n6), .Z(n9) );
  XNOR U14 ( .A(n8), .B(n9), .Z(c[2]) );
  XOR U15 ( .A(a[3]), .B(b[3]), .Z(n12) );
  NAND U16 ( .A(b[2]), .B(a[2]), .Z(n11) );
  NANDN U17 ( .A(n9), .B(n8), .Z(n10) );
  AND U18 ( .A(n11), .B(n10), .Z(n13) );
  XNOR U19 ( .A(n12), .B(n13), .Z(c[3]) );
  XOR U20 ( .A(a[4]), .B(b[4]), .Z(n16) );
  NAND U21 ( .A(b[3]), .B(a[3]), .Z(n15) );
  NANDN U22 ( .A(n13), .B(n12), .Z(n14) );
  AND U23 ( .A(n15), .B(n14), .Z(n17) );
  XNOR U24 ( .A(n16), .B(n17), .Z(c[4]) );
  XOR U25 ( .A(a[5]), .B(b[5]), .Z(n20) );
  NAND U26 ( .A(b[4]), .B(a[4]), .Z(n19) );
  NANDN U27 ( .A(n17), .B(n16), .Z(n18) );
  AND U28 ( .A(n19), .B(n18), .Z(n21) );
  XNOR U29 ( .A(n20), .B(n21), .Z(c[5]) );
  XOR U30 ( .A(a[6]), .B(b[6]), .Z(n24) );
  NAND U31 ( .A(b[5]), .B(a[5]), .Z(n23) );
  NANDN U32 ( .A(n21), .B(n20), .Z(n22) );
  AND U33 ( .A(n23), .B(n22), .Z(n25) );
  XNOR U34 ( .A(n24), .B(n25), .Z(c[6]) );
  XOR U35 ( .A(a[7]), .B(b[7]), .Z(n28) );
  NAND U36 ( .A(b[6]), .B(a[6]), .Z(n27) );
  NANDN U37 ( .A(n25), .B(n24), .Z(n26) );
  AND U38 ( .A(n27), .B(n26), .Z(n29) );
  XNOR U39 ( .A(n28), .B(n29), .Z(c[7]) );
  XOR U40 ( .A(a[8]), .B(b[8]), .Z(n32) );
  NAND U41 ( .A(b[7]), .B(a[7]), .Z(n31) );
  NANDN U42 ( .A(n29), .B(n28), .Z(n30) );
  AND U43 ( .A(n31), .B(n30), .Z(n33) );
  XNOR U44 ( .A(n32), .B(n33), .Z(c[8]) );
  XOR U45 ( .A(a[9]), .B(b[9]), .Z(n36) );
  NAND U46 ( .A(b[8]), .B(a[8]), .Z(n35) );
  NANDN U47 ( .A(n33), .B(n32), .Z(n34) );
  AND U48 ( .A(n35), .B(n34), .Z(n37) );
  XNOR U49 ( .A(n36), .B(n37), .Z(c[9]) );
  XOR U50 ( .A(a[10]), .B(b[10]), .Z(n40) );
  NAND U51 ( .A(b[9]), .B(a[9]), .Z(n39) );
  NANDN U52 ( .A(n37), .B(n36), .Z(n38) );
  AND U53 ( .A(n39), .B(n38), .Z(n41) );
  XNOR U54 ( .A(n40), .B(n41), .Z(c[10]) );
  XOR U55 ( .A(a[11]), .B(b[11]), .Z(n44) );
  NAND U56 ( .A(b[10]), .B(a[10]), .Z(n43) );
  NANDN U57 ( .A(n41), .B(n40), .Z(n42) );
  AND U58 ( .A(n43), .B(n42), .Z(n45) );
  XNOR U59 ( .A(n44), .B(n45), .Z(c[11]) );
  XOR U60 ( .A(a[12]), .B(b[12]), .Z(n48) );
  NAND U61 ( .A(b[11]), .B(a[11]), .Z(n47) );
  NANDN U62 ( .A(n45), .B(n44), .Z(n46) );
  AND U63 ( .A(n47), .B(n46), .Z(n49) );
  XNOR U64 ( .A(n48), .B(n49), .Z(c[12]) );
  XOR U65 ( .A(a[13]), .B(b[13]), .Z(n52) );
  NAND U66 ( .A(b[12]), .B(a[12]), .Z(n51) );
  NANDN U67 ( .A(n49), .B(n48), .Z(n50) );
  AND U68 ( .A(n51), .B(n50), .Z(n53) );
  XNOR U69 ( .A(n52), .B(n53), .Z(c[13]) );
  XOR U70 ( .A(a[14]), .B(b[14]), .Z(n56) );
  NAND U71 ( .A(b[13]), .B(a[13]), .Z(n55) );
  NANDN U72 ( .A(n53), .B(n52), .Z(n54) );
  AND U73 ( .A(n55), .B(n54), .Z(n57) );
  XNOR U74 ( .A(n56), .B(n57), .Z(c[14]) );
  XOR U75 ( .A(a[15]), .B(b[15]), .Z(n60) );
  NAND U76 ( .A(b[14]), .B(a[14]), .Z(n59) );
  NANDN U77 ( .A(n57), .B(n56), .Z(n58) );
  AND U78 ( .A(n59), .B(n58), .Z(n61) );
  XNOR U79 ( .A(n60), .B(n61), .Z(c[15]) );
  XOR U80 ( .A(a[16]), .B(b[16]), .Z(n64) );
  NAND U81 ( .A(b[15]), .B(a[15]), .Z(n63) );
  NANDN U82 ( .A(n61), .B(n60), .Z(n62) );
  AND U83 ( .A(n63), .B(n62), .Z(n65) );
  XNOR U84 ( .A(n64), .B(n65), .Z(c[16]) );
  XOR U85 ( .A(a[17]), .B(b[17]), .Z(n68) );
  NAND U86 ( .A(b[16]), .B(a[16]), .Z(n67) );
  NANDN U87 ( .A(n65), .B(n64), .Z(n66) );
  AND U88 ( .A(n67), .B(n66), .Z(n69) );
  XNOR U89 ( .A(n68), .B(n69), .Z(c[17]) );
  XOR U90 ( .A(a[18]), .B(b[18]), .Z(n72) );
  NAND U91 ( .A(b[17]), .B(a[17]), .Z(n71) );
  NANDN U92 ( .A(n69), .B(n68), .Z(n70) );
  AND U93 ( .A(n71), .B(n70), .Z(n73) );
  XNOR U94 ( .A(n72), .B(n73), .Z(c[18]) );
  XOR U95 ( .A(a[19]), .B(b[19]), .Z(n76) );
  NAND U96 ( .A(b[18]), .B(a[18]), .Z(n75) );
  NANDN U97 ( .A(n73), .B(n72), .Z(n74) );
  AND U98 ( .A(n75), .B(n74), .Z(n77) );
  XNOR U99 ( .A(n76), .B(n77), .Z(c[19]) );
  XOR U100 ( .A(a[20]), .B(b[20]), .Z(n80) );
  NAND U101 ( .A(b[19]), .B(a[19]), .Z(n79) );
  NANDN U102 ( .A(n77), .B(n76), .Z(n78) );
  AND U103 ( .A(n79), .B(n78), .Z(n81) );
  XNOR U104 ( .A(n80), .B(n81), .Z(c[20]) );
  XOR U105 ( .A(a[21]), .B(b[21]), .Z(n84) );
  NAND U106 ( .A(b[20]), .B(a[20]), .Z(n83) );
  NANDN U107 ( .A(n81), .B(n80), .Z(n82) );
  AND U108 ( .A(n83), .B(n82), .Z(n85) );
  XNOR U109 ( .A(n84), .B(n85), .Z(c[21]) );
  XOR U110 ( .A(a[22]), .B(b[22]), .Z(n88) );
  NAND U111 ( .A(b[21]), .B(a[21]), .Z(n87) );
  NANDN U112 ( .A(n85), .B(n84), .Z(n86) );
  AND U113 ( .A(n87), .B(n86), .Z(n89) );
  XNOR U114 ( .A(n88), .B(n89), .Z(c[22]) );
  XOR U115 ( .A(a[23]), .B(b[23]), .Z(n92) );
  NAND U116 ( .A(b[22]), .B(a[22]), .Z(n91) );
  NANDN U117 ( .A(n89), .B(n88), .Z(n90) );
  AND U118 ( .A(n91), .B(n90), .Z(n93) );
  XNOR U119 ( .A(n92), .B(n93), .Z(c[23]) );
  XOR U120 ( .A(a[24]), .B(b[24]), .Z(n96) );
  NAND U121 ( .A(b[23]), .B(a[23]), .Z(n95) );
  NANDN U122 ( .A(n93), .B(n92), .Z(n94) );
  AND U123 ( .A(n95), .B(n94), .Z(n97) );
  XNOR U124 ( .A(n96), .B(n97), .Z(c[24]) );
  XOR U125 ( .A(a[25]), .B(b[25]), .Z(n100) );
  NAND U126 ( .A(b[24]), .B(a[24]), .Z(n99) );
  NANDN U127 ( .A(n97), .B(n96), .Z(n98) );
  AND U128 ( .A(n99), .B(n98), .Z(n101) );
  XNOR U129 ( .A(n100), .B(n101), .Z(c[25]) );
  XOR U130 ( .A(a[26]), .B(b[26]), .Z(n104) );
  NAND U131 ( .A(b[25]), .B(a[25]), .Z(n103) );
  NANDN U132 ( .A(n101), .B(n100), .Z(n102) );
  AND U133 ( .A(n103), .B(n102), .Z(n105) );
  XNOR U134 ( .A(n104), .B(n105), .Z(c[26]) );
  XOR U135 ( .A(a[27]), .B(b[27]), .Z(n108) );
  NAND U136 ( .A(b[26]), .B(a[26]), .Z(n107) );
  NANDN U137 ( .A(n105), .B(n104), .Z(n106) );
  AND U138 ( .A(n107), .B(n106), .Z(n109) );
  XNOR U139 ( .A(n108), .B(n109), .Z(c[27]) );
  XOR U140 ( .A(a[28]), .B(b[28]), .Z(n112) );
  NAND U141 ( .A(b[27]), .B(a[27]), .Z(n111) );
  NANDN U142 ( .A(n109), .B(n108), .Z(n110) );
  AND U143 ( .A(n111), .B(n110), .Z(n113) );
  XNOR U144 ( .A(n112), .B(n113), .Z(c[28]) );
  XOR U145 ( .A(a[29]), .B(b[29]), .Z(n116) );
  NAND U146 ( .A(b[28]), .B(a[28]), .Z(n115) );
  NANDN U147 ( .A(n113), .B(n112), .Z(n114) );
  AND U148 ( .A(n115), .B(n114), .Z(n117) );
  XNOR U149 ( .A(n116), .B(n117), .Z(c[29]) );
  XOR U150 ( .A(a[30]), .B(b[30]), .Z(n120) );
  NAND U151 ( .A(b[29]), .B(a[29]), .Z(n119) );
  NANDN U152 ( .A(n117), .B(n116), .Z(n118) );
  AND U153 ( .A(n119), .B(n118), .Z(n121) );
  XNOR U154 ( .A(n120), .B(n121), .Z(c[30]) );
  NAND U155 ( .A(b[30]), .B(a[30]), .Z(n123) );
  NANDN U156 ( .A(n121), .B(n120), .Z(n122) );
  NAND U157 ( .A(n123), .B(n122), .Z(n124) );
  XOR U158 ( .A(a[31]), .B(b[31]), .Z(n125) );
  XOR U159 ( .A(n124), .B(n125), .Z(c[31]) );
  NAND U160 ( .A(b[31]), .B(a[31]), .Z(n127) );
  NAND U161 ( .A(n125), .B(n124), .Z(n126) );
  NAND U162 ( .A(n127), .B(n126), .Z(carry_on_d) );
endmodule

