
module matrixMultSeq ( clk, rst, x, y, o );
  input [31:0] x;
  input [31:0] y;
  output [31:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945;

  DFF \o_reg[31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \o_reg[30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \o_reg[29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \o_reg[28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \o_reg[27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \o_reg[26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \o_reg[25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \o_reg[24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \o_reg[23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \o_reg[22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \o_reg[21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \o_reg[20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \o_reg[19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \o_reg[18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \o_reg[17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \o_reg[16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \o_reg[15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \o_reg[14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \o_reg[13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \o_reg[12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \o_reg[11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \o_reg[10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \o_reg[9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \o_reg[8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \o_reg[7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \o_reg[6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \o_reg[5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \o_reg[4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \o_reg[3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \o_reg[2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \o_reg[1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \o_reg[0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  IV U3 ( .A(y[0]), .Z(n3637) );
  IV U4 ( .A(x[0]), .Z(n3680) );
  NOR U5 ( .A(n3637), .B(n3680), .Z(n1) );
  IV U6 ( .A(n1), .Z(n78) );
  IV U7 ( .A(o[0]), .Z(n3) );
  XOR U8 ( .A(n78), .B(n3), .Z(N33) );
  IV U9 ( .A(x[1]), .Z(n3625) );
  NOR U10 ( .A(n3637), .B(n3625), .Z(n5) );
  IV U11 ( .A(y[1]), .Z(n3773) );
  NOR U12 ( .A(n3773), .B(n3680), .Z(n2) );
  IV U13 ( .A(n2), .Z(n11) );
  XOR U14 ( .A(n11), .B(o[1]), .Z(n6) );
  XOR U15 ( .A(n5), .B(n6), .Z(n8) );
  NOR U16 ( .A(n78), .B(n3), .Z(n4) );
  IV U17 ( .A(n4), .Z(n7) );
  XOR U18 ( .A(n8), .B(n7), .Z(N34) );
  IV U19 ( .A(n5), .Z(n40) );
  NOR U20 ( .A(n40), .B(n6), .Z(n10) );
  NOR U21 ( .A(n8), .B(n7), .Z(n9) );
  NOR U22 ( .A(n10), .B(n9), .Z(n18) );
  IV U23 ( .A(o[1]), .Z(n12) );
  NOR U24 ( .A(n12), .B(n11), .Z(n14) );
  IV U25 ( .A(x[2]), .Z(n3619) );
  NOR U26 ( .A(n3637), .B(n3619), .Z(n24) );
  NOR U27 ( .A(n3773), .B(n3625), .Z(n21) );
  IV U28 ( .A(y[2]), .Z(n3647) );
  NOR U29 ( .A(n3680), .B(n3647), .Z(n13) );
  IV U30 ( .A(n13), .Z(n31) );
  XOR U31 ( .A(n31), .B(o[2]), .Z(n22) );
  XOR U32 ( .A(n21), .B(n22), .Z(n26) );
  XOR U33 ( .A(n24), .B(n26), .Z(n16) );
  XOR U34 ( .A(n14), .B(n16), .Z(n17) );
  XOR U35 ( .A(n18), .B(n17), .Z(N35) );
  IV U36 ( .A(n14), .Z(n15) );
  NOR U37 ( .A(n16), .B(n15), .Z(n20) );
  NOR U38 ( .A(n18), .B(n17), .Z(n19) );
  NOR U39 ( .A(n20), .B(n19), .Z(n37) );
  IV U40 ( .A(n21), .Z(n23) );
  NOR U41 ( .A(n23), .B(n22), .Z(n28) );
  IV U42 ( .A(n24), .Z(n25) );
  NOR U43 ( .A(n26), .B(n25), .Z(n27) );
  NOR U44 ( .A(n28), .B(n27), .Z(n35) );
  IV U45 ( .A(x[3]), .Z(n3635) );
  NOR U46 ( .A(n3635), .B(n3637), .Z(n108) );
  NOR U47 ( .A(n3647), .B(n3625), .Z(n29) );
  XOR U48 ( .A(n108), .B(n29), .Z(n41) );
  IV U49 ( .A(o[2]), .Z(n30) );
  NOR U50 ( .A(n31), .B(n30), .Z(n48) );
  IV U51 ( .A(y[3]), .Z(n3787) );
  NOR U52 ( .A(n3680), .B(n3787), .Z(n46) );
  NOR U53 ( .A(n3773), .B(n3619), .Z(n32) );
  IV U54 ( .A(n32), .Z(n55) );
  XOR U55 ( .A(n55), .B(o[3]), .Z(n47) );
  XOR U56 ( .A(n46), .B(n47), .Z(n50) );
  XOR U57 ( .A(n48), .B(n50), .Z(n42) );
  XOR U58 ( .A(n41), .B(n42), .Z(n34) );
  XOR U59 ( .A(n35), .B(n34), .Z(n33) );
  IV U60 ( .A(n33), .Z(n36) );
  XOR U61 ( .A(n37), .B(n36), .Z(N36) );
  NOR U62 ( .A(n35), .B(n34), .Z(n39) );
  NOR U63 ( .A(n37), .B(n36), .Z(n38) );
  NOR U64 ( .A(n39), .B(n38), .Z(n61) );
  NOR U65 ( .A(n3635), .B(n3647), .Z(n83) );
  IV U66 ( .A(n83), .Z(n333) );
  NOR U67 ( .A(n333), .B(n40), .Z(n45) );
  IV U68 ( .A(n41), .Z(n43) );
  NOR U69 ( .A(n43), .B(n42), .Z(n44) );
  NOR U70 ( .A(n45), .B(n44), .Z(n59) );
  IV U71 ( .A(n59), .Z(n57) );
  IV U72 ( .A(n46), .Z(n211) );
  NOR U73 ( .A(n211), .B(n47), .Z(n52) );
  IV U74 ( .A(n48), .Z(n49) );
  NOR U75 ( .A(n50), .B(n49), .Z(n51) );
  NOR U76 ( .A(n52), .B(n51), .Z(n68) );
  IV U77 ( .A(x[4]), .Z(n3650) );
  NOR U78 ( .A(n3650), .B(n3637), .Z(n156) );
  IV U79 ( .A(y[4]), .Z(n3628) );
  NOR U80 ( .A(n3628), .B(n3680), .Z(n144) );
  XOR U81 ( .A(n156), .B(n144), .Z(n53) );
  IV U82 ( .A(n53), .Z(n80) );
  NOR U83 ( .A(n3625), .B(n3787), .Z(n79) );
  XOR U84 ( .A(n80), .B(n79), .Z(n64) );
  IV U85 ( .A(o[3]), .Z(n54) );
  NOR U86 ( .A(n55), .B(n54), .Z(n73) );
  NOR U87 ( .A(n3647), .B(n3619), .Z(n71) );
  NOR U88 ( .A(n3773), .B(n3635), .Z(n56) );
  IV U89 ( .A(n56), .Z(n85) );
  XOR U90 ( .A(n85), .B(o[4]), .Z(n72) );
  XOR U91 ( .A(n71), .B(n72), .Z(n75) );
  XOR U92 ( .A(n73), .B(n75), .Z(n65) );
  XOR U93 ( .A(n64), .B(n65), .Z(n66) );
  XOR U94 ( .A(n68), .B(n66), .Z(n58) );
  XOR U95 ( .A(n57), .B(n58), .Z(n60) );
  XOR U96 ( .A(n61), .B(n60), .Z(N37) );
  NOR U97 ( .A(n59), .B(n58), .Z(n63) );
  NOR U98 ( .A(n61), .B(n60), .Z(n62) );
  NOR U99 ( .A(n63), .B(n62), .Z(n92) );
  NOR U100 ( .A(n65), .B(n64), .Z(n70) );
  IV U101 ( .A(n66), .Z(n67) );
  NOR U102 ( .A(n68), .B(n67), .Z(n69) );
  NOR U103 ( .A(n70), .B(n69), .Z(n90) );
  IV U104 ( .A(n71), .Z(n416) );
  NOR U105 ( .A(n416), .B(n72), .Z(n77) );
  IV U106 ( .A(n73), .Z(n74) );
  NOR U107 ( .A(n75), .B(n74), .Z(n76) );
  NOR U108 ( .A(n77), .B(n76), .Z(n127) );
  NOR U109 ( .A(n3628), .B(n3650), .Z(n223) );
  IV U110 ( .A(n223), .Z(n915) );
  NOR U111 ( .A(n915), .B(n78), .Z(n82) );
  IV U112 ( .A(n79), .Z(n389) );
  NOR U113 ( .A(n389), .B(n80), .Z(n81) );
  NOR U114 ( .A(n82), .B(n81), .Z(n124) );
  IV U115 ( .A(y[5]), .Z(n3746) );
  NOR U116 ( .A(n3680), .B(n3746), .Z(n103) );
  IV U117 ( .A(n103), .Z(n252) );
  IV U118 ( .A(x[5]), .Z(n3740) );
  NOR U119 ( .A(n3740), .B(n3637), .Z(n264) );
  XOR U120 ( .A(n264), .B(n83), .Z(n110) );
  NOR U121 ( .A(n3625), .B(n3628), .Z(n111) );
  XOR U122 ( .A(n110), .B(n111), .Z(n102) );
  XOR U123 ( .A(n252), .B(n102), .Z(n104) );
  NOR U124 ( .A(n3787), .B(n3619), .Z(n95) );
  NOR U125 ( .A(n3773), .B(n3650), .Z(n84) );
  IV U126 ( .A(n84), .Z(n120) );
  XOR U127 ( .A(n120), .B(o[5]), .Z(n96) );
  XOR U128 ( .A(n95), .B(n96), .Z(n99) );
  IV U129 ( .A(o[4]), .Z(n86) );
  NOR U130 ( .A(n86), .B(n85), .Z(n87) );
  IV U131 ( .A(n87), .Z(n98) );
  XOR U132 ( .A(n99), .B(n98), .Z(n105) );
  XOR U133 ( .A(n104), .B(n105), .Z(n123) );
  XOR U134 ( .A(n124), .B(n123), .Z(n125) );
  XOR U135 ( .A(n127), .B(n125), .Z(n89) );
  XOR U136 ( .A(n90), .B(n89), .Z(n88) );
  IV U137 ( .A(n88), .Z(n91) );
  XOR U138 ( .A(n92), .B(n91), .Z(N38) );
  NOR U139 ( .A(n90), .B(n89), .Z(n94) );
  NOR U140 ( .A(n92), .B(n91), .Z(n93) );
  NOR U141 ( .A(n94), .B(n93), .Z(n172) );
  IV U142 ( .A(n95), .Z(n97) );
  NOR U143 ( .A(n97), .B(n96), .Z(n101) );
  NOR U144 ( .A(n99), .B(n98), .Z(n100) );
  NOR U145 ( .A(n101), .B(n100), .Z(n132) );
  NOR U146 ( .A(n103), .B(n102), .Z(n107) );
  NOR U147 ( .A(n105), .B(n104), .Z(n106) );
  NOR U148 ( .A(n107), .B(n106), .Z(n130) );
  XOR U149 ( .A(n132), .B(n130), .Z(n134) );
  NOR U150 ( .A(n3647), .B(n3740), .Z(n168) );
  IV U151 ( .A(n168), .Z(n198) );
  IV U152 ( .A(n108), .Z(n109) );
  NOR U153 ( .A(n198), .B(n109), .Z(n115) );
  IV U154 ( .A(n110), .Z(n113) );
  IV U155 ( .A(n111), .Z(n112) );
  NOR U156 ( .A(n113), .B(n112), .Z(n114) );
  NOR U157 ( .A(n115), .B(n114), .Z(n141) );
  IV U158 ( .A(x[6]), .Z(n3748) );
  NOR U159 ( .A(n3748), .B(n3637), .Z(n430) );
  NOR U160 ( .A(n3647), .B(n3650), .Z(n116) );
  XOR U161 ( .A(n430), .B(n116), .Z(n159) );
  NOR U162 ( .A(n3619), .B(n3628), .Z(n118) );
  IV U163 ( .A(y[6]), .Z(n3633) );
  NOR U164 ( .A(n3680), .B(n3633), .Z(n117) );
  XOR U165 ( .A(n118), .B(n117), .Z(n119) );
  IV U166 ( .A(n119), .Z(n146) );
  NOR U167 ( .A(n3625), .B(n3746), .Z(n145) );
  XOR U168 ( .A(n146), .B(n145), .Z(n160) );
  XOR U169 ( .A(n159), .B(n160), .Z(n138) );
  IV U170 ( .A(o[5]), .Z(n121) );
  NOR U171 ( .A(n121), .B(n120), .Z(n151) );
  NOR U172 ( .A(n3787), .B(n3635), .Z(n149) );
  NOR U173 ( .A(n3773), .B(n3740), .Z(n122) );
  IV U174 ( .A(n122), .Z(n164) );
  XOR U175 ( .A(n164), .B(o[6]), .Z(n150) );
  XOR U176 ( .A(n149), .B(n150), .Z(n153) );
  XOR U177 ( .A(n151), .B(n153), .Z(n137) );
  XOR U178 ( .A(n138), .B(n137), .Z(n139) );
  XOR U179 ( .A(n141), .B(n139), .Z(n133) );
  XOR U180 ( .A(n134), .B(n133), .Z(n171) );
  NOR U181 ( .A(n124), .B(n123), .Z(n129) );
  IV U182 ( .A(n125), .Z(n126) );
  NOR U183 ( .A(n127), .B(n126), .Z(n128) );
  NOR U184 ( .A(n129), .B(n128), .Z(n169) );
  XOR U185 ( .A(n171), .B(n169), .Z(n174) );
  XOR U186 ( .A(n172), .B(n174), .Z(N39) );
  IV U187 ( .A(n130), .Z(n131) );
  NOR U188 ( .A(n132), .B(n131), .Z(n136) );
  NOR U189 ( .A(n134), .B(n133), .Z(n135) );
  NOR U190 ( .A(n136), .B(n135), .Z(n180) );
  NOR U191 ( .A(n138), .B(n137), .Z(n143) );
  IV U192 ( .A(n139), .Z(n140) );
  NOR U193 ( .A(n141), .B(n140), .Z(n142) );
  NOR U194 ( .A(n143), .B(n142), .Z(n229) );
  NOR U195 ( .A(n3619), .B(n3633), .Z(n218) );
  IV U196 ( .A(n218), .Z(n1155) );
  IV U197 ( .A(n144), .Z(n355) );
  NOR U198 ( .A(n1155), .B(n355), .Z(n148) );
  IV U199 ( .A(n145), .Z(n192) );
  NOR U200 ( .A(n192), .B(n146), .Z(n147) );
  NOR U201 ( .A(n148), .B(n147), .Z(n227) );
  IV U202 ( .A(n149), .Z(n944) );
  NOR U203 ( .A(n944), .B(n150), .Z(n155) );
  IV U204 ( .A(n151), .Z(n152) );
  NOR U205 ( .A(n153), .B(n152), .Z(n154) );
  NOR U206 ( .A(n155), .B(n154), .Z(n189) );
  NOR U207 ( .A(n3748), .B(n3647), .Z(n217) );
  IV U208 ( .A(n217), .Z(n158) );
  IV U209 ( .A(n156), .Z(n157) );
  NOR U210 ( .A(n158), .B(n157), .Z(n163) );
  IV U211 ( .A(n159), .Z(n161) );
  NOR U212 ( .A(n161), .B(n160), .Z(n162) );
  NOR U213 ( .A(n163), .B(n162), .Z(n187) );
  IV U214 ( .A(o[6]), .Z(n165) );
  NOR U215 ( .A(n165), .B(n164), .Z(n206) );
  NOR U216 ( .A(n3628), .B(n3635), .Z(n204) );
  NOR U217 ( .A(n3773), .B(n3748), .Z(n166) );
  IV U218 ( .A(n166), .Z(n220) );
  XOR U219 ( .A(n220), .B(o[7]), .Z(n205) );
  XOR U220 ( .A(n204), .B(n205), .Z(n208) );
  XOR U221 ( .A(n206), .B(n208), .Z(n200) );
  NOR U222 ( .A(n3619), .B(n3746), .Z(n903) );
  NOR U223 ( .A(n3625), .B(n3633), .Z(n712) );
  XOR U224 ( .A(n903), .B(n712), .Z(n193) );
  IV U225 ( .A(y[7]), .Z(n3687) );
  NOR U226 ( .A(n3687), .B(n3680), .Z(n949) );
  NOR U227 ( .A(n3650), .B(n3787), .Z(n605) );
  XOR U228 ( .A(n949), .B(n605), .Z(n167) );
  IV U229 ( .A(n167), .Z(n213) );
  IV U230 ( .A(x[7]), .Z(n3682) );
  NOR U231 ( .A(n3682), .B(n3637), .Z(n212) );
  XOR U232 ( .A(n213), .B(n212), .Z(n195) );
  XOR U233 ( .A(n193), .B(n195), .Z(n199) );
  XOR U234 ( .A(n168), .B(n199), .Z(n201) );
  XOR U235 ( .A(n200), .B(n201), .Z(n185) );
  XOR U236 ( .A(n187), .B(n185), .Z(n188) );
  XOR U237 ( .A(n189), .B(n188), .Z(n225) );
  XOR U238 ( .A(n227), .B(n225), .Z(n228) );
  XOR U239 ( .A(n229), .B(n228), .Z(n178) );
  XOR U240 ( .A(n180), .B(n178), .Z(n182) );
  IV U241 ( .A(n169), .Z(n170) );
  NOR U242 ( .A(n171), .B(n170), .Z(n176) );
  IV U243 ( .A(n172), .Z(n173) );
  NOR U244 ( .A(n174), .B(n173), .Z(n175) );
  NOR U245 ( .A(n176), .B(n175), .Z(n177) );
  IV U246 ( .A(n177), .Z(n181) );
  XOR U247 ( .A(n182), .B(n181), .Z(N40) );
  IV U248 ( .A(n178), .Z(n179) );
  NOR U249 ( .A(n180), .B(n179), .Z(n184) );
  NOR U250 ( .A(n182), .B(n181), .Z(n183) );
  NOR U251 ( .A(n184), .B(n183), .Z(n291) );
  IV U252 ( .A(n185), .Z(n186) );
  NOR U253 ( .A(n187), .B(n186), .Z(n191) );
  NOR U254 ( .A(n189), .B(n188), .Z(n190) );
  NOR U255 ( .A(n191), .B(n190), .Z(n235) );
  NOR U256 ( .A(n1155), .B(n192), .Z(n197) );
  IV U257 ( .A(n193), .Z(n194) );
  NOR U258 ( .A(n195), .B(n194), .Z(n196) );
  NOR U259 ( .A(n197), .B(n196), .Z(n233) );
  NOR U260 ( .A(n199), .B(n198), .Z(n203) );
  NOR U261 ( .A(n201), .B(n200), .Z(n202) );
  NOR U262 ( .A(n203), .B(n202), .Z(n242) );
  IV U263 ( .A(n204), .Z(n1072) );
  NOR U264 ( .A(n1072), .B(n205), .Z(n210) );
  IV U265 ( .A(n206), .Z(n207) );
  NOR U266 ( .A(n208), .B(n207), .Z(n209) );
  NOR U267 ( .A(n210), .B(n209), .Z(n239) );
  NOR U268 ( .A(n3650), .B(n3687), .Z(n424) );
  IV U269 ( .A(n424), .Z(n1640) );
  NOR U270 ( .A(n1640), .B(n211), .Z(n215) );
  IV U271 ( .A(n212), .Z(n820) );
  NOR U272 ( .A(n820), .B(n213), .Z(n214) );
  NOR U273 ( .A(n215), .B(n214), .Z(n249) );
  IV U274 ( .A(x[8]), .Z(n3749) );
  NOR U275 ( .A(n3637), .B(n3749), .Z(n216) );
  NOR U276 ( .A(n3787), .B(n3740), .Z(n769) );
  XOR U277 ( .A(n216), .B(n769), .Z(n266) );
  XOR U278 ( .A(n218), .B(n217), .Z(n272) );
  NOR U279 ( .A(n3625), .B(n3687), .Z(n219) );
  IV U280 ( .A(n219), .Z(n254) );
  IV U281 ( .A(y[8]), .Z(n3462) );
  NOR U282 ( .A(n3462), .B(n3680), .Z(n697) );
  NOR U283 ( .A(n3635), .B(n3746), .Z(n1489) );
  XOR U284 ( .A(n697), .B(n1489), .Z(n253) );
  XOR U285 ( .A(n254), .B(n253), .Z(n274) );
  XOR U286 ( .A(n272), .B(n274), .Z(n268) );
  XOR U287 ( .A(n266), .B(n268), .Z(n246) );
  IV U288 ( .A(o[7]), .Z(n221) );
  NOR U289 ( .A(n221), .B(n220), .Z(n259) );
  NOR U290 ( .A(n3682), .B(n3773), .Z(n222) );
  IV U291 ( .A(n222), .Z(n284) );
  XOR U292 ( .A(n284), .B(o[8]), .Z(n258) );
  XOR U293 ( .A(n223), .B(n258), .Z(n261) );
  XOR U294 ( .A(n259), .B(n261), .Z(n245) );
  XOR U295 ( .A(n246), .B(n245), .Z(n247) );
  XOR U296 ( .A(n249), .B(n247), .Z(n238) );
  XOR U297 ( .A(n239), .B(n238), .Z(n240) );
  XOR U298 ( .A(n242), .B(n240), .Z(n232) );
  XOR U299 ( .A(n233), .B(n232), .Z(n224) );
  IV U300 ( .A(n224), .Z(n234) );
  XOR U301 ( .A(n235), .B(n234), .Z(n290) );
  IV U302 ( .A(n225), .Z(n226) );
  NOR U303 ( .A(n227), .B(n226), .Z(n231) );
  NOR U304 ( .A(n229), .B(n228), .Z(n230) );
  NOR U305 ( .A(n231), .B(n230), .Z(n288) );
  XOR U306 ( .A(n290), .B(n288), .Z(n293) );
  XOR U307 ( .A(n291), .B(n293), .Z(N41) );
  NOR U308 ( .A(n233), .B(n232), .Z(n237) );
  NOR U309 ( .A(n235), .B(n234), .Z(n236) );
  NOR U310 ( .A(n237), .B(n236), .Z(n298) );
  NOR U311 ( .A(n239), .B(n238), .Z(n244) );
  IV U312 ( .A(n240), .Z(n241) );
  NOR U313 ( .A(n242), .B(n241), .Z(n243) );
  NOR U314 ( .A(n244), .B(n243), .Z(n307) );
  NOR U315 ( .A(n246), .B(n245), .Z(n251) );
  IV U316 ( .A(n247), .Z(n248) );
  NOR U317 ( .A(n249), .B(n248), .Z(n250) );
  NOR U318 ( .A(n251), .B(n250), .Z(n304) );
  NOR U319 ( .A(n3462), .B(n3635), .Z(n425) );
  IV U320 ( .A(n425), .Z(n1848) );
  NOR U321 ( .A(n1848), .B(n252), .Z(n257) );
  IV U322 ( .A(n253), .Z(n255) );
  NOR U323 ( .A(n255), .B(n254), .Z(n256) );
  NOR U324 ( .A(n257), .B(n256), .Z(n311) );
  NOR U325 ( .A(n915), .B(n258), .Z(n263) );
  IV U326 ( .A(n259), .Z(n260) );
  NOR U327 ( .A(n261), .B(n260), .Z(n262) );
  NOR U328 ( .A(n263), .B(n262), .Z(n310) );
  XOR U329 ( .A(n311), .B(n310), .Z(n312) );
  NOR U330 ( .A(n3787), .B(n3749), .Z(n435) );
  IV U331 ( .A(n435), .Z(n1621) );
  IV U332 ( .A(n264), .Z(n265) );
  NOR U333 ( .A(n1621), .B(n265), .Z(n270) );
  IV U334 ( .A(n266), .Z(n267) );
  NOR U335 ( .A(n268), .B(n267), .Z(n269) );
  NOR U336 ( .A(n270), .B(n269), .Z(n365) );
  NOR U337 ( .A(n3633), .B(n3748), .Z(n517) );
  IV U338 ( .A(n517), .Z(n271) );
  NOR U339 ( .A(n271), .B(n416), .Z(n276) );
  IV U340 ( .A(n272), .Z(n273) );
  NOR U341 ( .A(n274), .B(n273), .Z(n275) );
  NOR U342 ( .A(n276), .B(n275), .Z(n362) );
  NOR U343 ( .A(n3647), .B(n3682), .Z(n278) );
  NOR U344 ( .A(n3633), .B(n3635), .Z(n277) );
  XOR U345 ( .A(n278), .B(n277), .Z(n335) );
  IV U346 ( .A(x[9]), .Z(n3765) );
  NOR U347 ( .A(n3765), .B(n3637), .Z(n279) );
  IV U348 ( .A(n279), .Z(n357) );
  IV U349 ( .A(y[9]), .Z(n3646) );
  NOR U350 ( .A(n3680), .B(n3646), .Z(n1633) );
  NOR U351 ( .A(n3628), .B(n3740), .Z(n280) );
  XOR U352 ( .A(n1633), .B(n280), .Z(n356) );
  XOR U353 ( .A(n357), .B(n356), .Z(n336) );
  XOR U354 ( .A(n335), .B(n336), .Z(n328) );
  NOR U355 ( .A(n3687), .B(n3619), .Z(n281) );
  IV U356 ( .A(n281), .Z(n343) );
  NOR U357 ( .A(n3462), .B(n3625), .Z(n283) );
  NOR U358 ( .A(n3748), .B(n3787), .Z(n282) );
  XOR U359 ( .A(n283), .B(n282), .Z(n341) );
  XOR U360 ( .A(n343), .B(n341), .Z(n325) );
  IV U361 ( .A(o[8]), .Z(n285) );
  NOR U362 ( .A(n285), .B(n284), .Z(n320) );
  NOR U363 ( .A(n3746), .B(n3650), .Z(n317) );
  NOR U364 ( .A(n3749), .B(n3773), .Z(n286) );
  IV U365 ( .A(n286), .Z(n346) );
  XOR U366 ( .A(n346), .B(o[9]), .Z(n319) );
  XOR U367 ( .A(n317), .B(n319), .Z(n322) );
  XOR U368 ( .A(n320), .B(n322), .Z(n326) );
  XOR U369 ( .A(n325), .B(n326), .Z(n327) );
  XOR U370 ( .A(n328), .B(n327), .Z(n361) );
  XOR U371 ( .A(n362), .B(n361), .Z(n363) );
  XOR U372 ( .A(n365), .B(n363), .Z(n313) );
  XOR U373 ( .A(n312), .B(n313), .Z(n303) );
  XOR U374 ( .A(n304), .B(n303), .Z(n305) );
  XOR U375 ( .A(n307), .B(n305), .Z(n297) );
  XOR U376 ( .A(n298), .B(n297), .Z(n287) );
  IV U377 ( .A(n287), .Z(n300) );
  IV U378 ( .A(n288), .Z(n289) );
  NOR U379 ( .A(n290), .B(n289), .Z(n295) );
  IV U380 ( .A(n291), .Z(n292) );
  NOR U381 ( .A(n293), .B(n292), .Z(n294) );
  NOR U382 ( .A(n295), .B(n294), .Z(n296) );
  IV U383 ( .A(n296), .Z(n299) );
  XOR U384 ( .A(n300), .B(n299), .Z(N42) );
  NOR U385 ( .A(n298), .B(n297), .Z(n302) );
  NOR U386 ( .A(n300), .B(n299), .Z(n301) );
  NOR U387 ( .A(n302), .B(n301), .Z(n444) );
  NOR U388 ( .A(n304), .B(n303), .Z(n309) );
  IV U389 ( .A(n305), .Z(n306) );
  NOR U390 ( .A(n307), .B(n306), .Z(n308) );
  NOR U391 ( .A(n309), .B(n308), .Z(n441) );
  NOR U392 ( .A(n311), .B(n310), .Z(n316) );
  IV U393 ( .A(n312), .Z(n314) );
  NOR U394 ( .A(n314), .B(n313), .Z(n315) );
  NOR U395 ( .A(n316), .B(n315), .Z(n371) );
  IV U396 ( .A(n317), .Z(n318) );
  NOR U397 ( .A(n319), .B(n318), .Z(n324) );
  IV U398 ( .A(n320), .Z(n321) );
  NOR U399 ( .A(n322), .B(n321), .Z(n323) );
  NOR U400 ( .A(n324), .B(n323), .Z(n377) );
  NOR U401 ( .A(n326), .B(n325), .Z(n331) );
  IV U402 ( .A(n327), .Z(n329) );
  NOR U403 ( .A(n329), .B(n328), .Z(n330) );
  NOR U404 ( .A(n331), .B(n330), .Z(n376) );
  XOR U405 ( .A(n377), .B(n376), .Z(n332) );
  IV U406 ( .A(n332), .Z(n378) );
  NOR U407 ( .A(n3682), .B(n3633), .Z(n617) );
  IV U408 ( .A(n617), .Z(n334) );
  NOR U409 ( .A(n334), .B(n333), .Z(n339) );
  IV U410 ( .A(n335), .Z(n337) );
  NOR U411 ( .A(n337), .B(n336), .Z(n338) );
  NOR U412 ( .A(n339), .B(n338), .Z(n340) );
  IV U413 ( .A(n340), .Z(n386) );
  NOR U414 ( .A(n3748), .B(n3462), .Z(n731) );
  IV U415 ( .A(n731), .Z(n806) );
  NOR U416 ( .A(n806), .B(n389), .Z(n345) );
  IV U417 ( .A(n341), .Z(n342) );
  NOR U418 ( .A(n343), .B(n342), .Z(n344) );
  NOR U419 ( .A(n345), .B(n344), .Z(n399) );
  IV U420 ( .A(o[9]), .Z(n347) );
  NOR U421 ( .A(n347), .B(n346), .Z(n405) );
  NOR U422 ( .A(n3746), .B(n3740), .Z(n402) );
  NOR U423 ( .A(n3765), .B(n3773), .Z(n348) );
  IV U424 ( .A(n348), .Z(n429) );
  XOR U425 ( .A(n429), .B(o[10]), .Z(n403) );
  XOR U426 ( .A(n402), .B(n403), .Z(n407) );
  XOR U427 ( .A(n405), .B(n407), .Z(n397) );
  NOR U428 ( .A(n3635), .B(n3687), .Z(n410) );
  NOR U429 ( .A(n3633), .B(n3650), .Z(n349) );
  IV U430 ( .A(n349), .Z(n419) );
  NOR U431 ( .A(n3647), .B(n3749), .Z(n587) );
  NOR U432 ( .A(n3462), .B(n3619), .Z(n350) );
  XOR U433 ( .A(n587), .B(n350), .Z(n418) );
  XOR U434 ( .A(n419), .B(n418), .Z(n411) );
  XOR U435 ( .A(n410), .B(n411), .Z(n412) );
  NOR U436 ( .A(n3625), .B(n3646), .Z(n351) );
  NOR U437 ( .A(n3787), .B(n3682), .Z(n478) );
  XOR U438 ( .A(n351), .B(n478), .Z(n390) );
  IV U439 ( .A(x[10]), .Z(n3779) );
  NOR U440 ( .A(n3637), .B(n3779), .Z(n353) );
  NOR U441 ( .A(n3748), .B(n3628), .Z(n352) );
  XOR U442 ( .A(n353), .B(n352), .Z(n354) );
  IV U443 ( .A(n354), .Z(n432) );
  IV U444 ( .A(y[10]), .Z(n3622) );
  NOR U445 ( .A(n3680), .B(n3622), .Z(n431) );
  XOR U446 ( .A(n432), .B(n431), .Z(n392) );
  XOR U447 ( .A(n390), .B(n392), .Z(n413) );
  XOR U448 ( .A(n412), .B(n413), .Z(n395) );
  XOR U449 ( .A(n397), .B(n395), .Z(n398) );
  XOR U450 ( .A(n399), .B(n398), .Z(n384) );
  NOR U451 ( .A(n3646), .B(n3740), .Z(n719) );
  IV U452 ( .A(n719), .Z(n1459) );
  NOR U453 ( .A(n1459), .B(n355), .Z(n360) );
  IV U454 ( .A(n356), .Z(n358) );
  NOR U455 ( .A(n358), .B(n357), .Z(n359) );
  NOR U456 ( .A(n360), .B(n359), .Z(n382) );
  XOR U457 ( .A(n384), .B(n382), .Z(n385) );
  XOR U458 ( .A(n386), .B(n385), .Z(n379) );
  XOR U459 ( .A(n378), .B(n379), .Z(n370) );
  NOR U460 ( .A(n362), .B(n361), .Z(n367) );
  IV U461 ( .A(n363), .Z(n364) );
  NOR U462 ( .A(n365), .B(n364), .Z(n366) );
  NOR U463 ( .A(n367), .B(n366), .Z(n368) );
  XOR U464 ( .A(n370), .B(n368), .Z(n373) );
  XOR U465 ( .A(n371), .B(n373), .Z(n443) );
  XOR U466 ( .A(n441), .B(n443), .Z(n446) );
  XOR U467 ( .A(n444), .B(n446), .Z(N43) );
  IV U468 ( .A(n368), .Z(n369) );
  NOR U469 ( .A(n370), .B(n369), .Z(n375) );
  IV U470 ( .A(n371), .Z(n372) );
  NOR U471 ( .A(n373), .B(n372), .Z(n374) );
  NOR U472 ( .A(n375), .B(n374), .Z(n450) );
  NOR U473 ( .A(n377), .B(n376), .Z(n381) );
  NOR U474 ( .A(n379), .B(n378), .Z(n380) );
  NOR U475 ( .A(n381), .B(n380), .Z(n461) );
  IV U476 ( .A(n461), .Z(n440) );
  IV U477 ( .A(n382), .Z(n383) );
  NOR U478 ( .A(n384), .B(n383), .Z(n388) );
  NOR U479 ( .A(n386), .B(n385), .Z(n387) );
  NOR U480 ( .A(n388), .B(n387), .Z(n457) );
  NOR U481 ( .A(n3682), .B(n3646), .Z(n927) );
  IV U482 ( .A(n927), .Z(n1015) );
  NOR U483 ( .A(n1015), .B(n389), .Z(n394) );
  IV U484 ( .A(n390), .Z(n391) );
  NOR U485 ( .A(n392), .B(n391), .Z(n393) );
  NOR U486 ( .A(n394), .B(n393), .Z(n465) );
  IV U487 ( .A(n395), .Z(n396) );
  NOR U488 ( .A(n397), .B(n396), .Z(n401) );
  NOR U489 ( .A(n399), .B(n398), .Z(n400) );
  NOR U490 ( .A(n401), .B(n400), .Z(n464) );
  XOR U491 ( .A(n465), .B(n464), .Z(n466) );
  IV U492 ( .A(n402), .Z(n404) );
  NOR U493 ( .A(n404), .B(n403), .Z(n409) );
  IV U494 ( .A(n405), .Z(n406) );
  NOR U495 ( .A(n407), .B(n406), .Z(n408) );
  NOR U496 ( .A(n409), .B(n408), .Z(n472) );
  IV U497 ( .A(n410), .Z(n506) );
  NOR U498 ( .A(n506), .B(n411), .Z(n415) );
  NOR U499 ( .A(n413), .B(n412), .Z(n414) );
  NOR U500 ( .A(n415), .B(n414), .Z(n471) );
  XOR U501 ( .A(n472), .B(n471), .Z(n473) );
  NOR U502 ( .A(n3749), .B(n3462), .Z(n963) );
  IV U503 ( .A(n963), .Z(n417) );
  NOR U504 ( .A(n417), .B(n416), .Z(n422) );
  IV U505 ( .A(n418), .Z(n420) );
  NOR U506 ( .A(n420), .B(n419), .Z(n421) );
  NOR U507 ( .A(n422), .B(n421), .Z(n537) );
  IV U508 ( .A(y[11]), .Z(n3781) );
  NOR U509 ( .A(n3680), .B(n3781), .Z(n423) );
  NOR U510 ( .A(n3625), .B(n3622), .Z(n790) );
  XOR U511 ( .A(n423), .B(n790), .Z(n487) );
  XOR U512 ( .A(n425), .B(n424), .Z(n508) );
  NOR U513 ( .A(n3646), .B(n3619), .Z(n426) );
  IV U514 ( .A(n426), .Z(n1829) );
  XOR U515 ( .A(n508), .B(n1829), .Z(n488) );
  XOR U516 ( .A(n487), .B(n488), .Z(n534) );
  NOR U517 ( .A(n3633), .B(n3740), .Z(n498) );
  NOR U518 ( .A(n3779), .B(n3773), .Z(n427) );
  IV U519 ( .A(n427), .Z(n524) );
  XOR U520 ( .A(n524), .B(o[11]), .Z(n499) );
  XOR U521 ( .A(n498), .B(n499), .Z(n502) );
  IV U522 ( .A(o[10]), .Z(n428) );
  NOR U523 ( .A(n429), .B(n428), .Z(n500) );
  XOR U524 ( .A(n502), .B(n500), .Z(n533) );
  XOR U525 ( .A(n534), .B(n533), .Z(n535) );
  XOR U526 ( .A(n537), .B(n535), .Z(n529) );
  NOR U527 ( .A(n3779), .B(n3628), .Z(n722) );
  IV U528 ( .A(n722), .Z(n772) );
  IV U529 ( .A(n430), .Z(n493) );
  NOR U530 ( .A(n772), .B(n493), .Z(n434) );
  IV U531 ( .A(n431), .Z(n486) );
  NOR U532 ( .A(n486), .B(n432), .Z(n433) );
  NOR U533 ( .A(n434), .B(n433), .Z(n526) );
  NOR U534 ( .A(n3628), .B(n3682), .Z(n436) );
  XOR U535 ( .A(n436), .B(n435), .Z(n481) );
  IV U536 ( .A(x[11]), .Z(n3062) );
  NOR U537 ( .A(n3637), .B(n3062), .Z(n438) );
  NOR U538 ( .A(n3746), .B(n3748), .Z(n437) );
  XOR U539 ( .A(n438), .B(n437), .Z(n439) );
  IV U540 ( .A(n439), .Z(n495) );
  NOR U541 ( .A(n3765), .B(n3647), .Z(n494) );
  XOR U542 ( .A(n495), .B(n494), .Z(n482) );
  XOR U543 ( .A(n481), .B(n482), .Z(n525) );
  XOR U544 ( .A(n526), .B(n525), .Z(n527) );
  XOR U545 ( .A(n529), .B(n527), .Z(n474) );
  XOR U546 ( .A(n473), .B(n474), .Z(n467) );
  XOR U547 ( .A(n466), .B(n467), .Z(n459) );
  XOR U548 ( .A(n457), .B(n459), .Z(n460) );
  XOR U549 ( .A(n440), .B(n460), .Z(n452) );
  XOR U550 ( .A(n450), .B(n452), .Z(n454) );
  IV U551 ( .A(n441), .Z(n442) );
  NOR U552 ( .A(n443), .B(n442), .Z(n448) );
  IV U553 ( .A(n444), .Z(n445) );
  NOR U554 ( .A(n446), .B(n445), .Z(n447) );
  NOR U555 ( .A(n448), .B(n447), .Z(n449) );
  IV U556 ( .A(n449), .Z(n453) );
  XOR U557 ( .A(n454), .B(n453), .Z(N44) );
  IV U558 ( .A(n450), .Z(n451) );
  NOR U559 ( .A(n452), .B(n451), .Z(n456) );
  NOR U560 ( .A(n454), .B(n453), .Z(n455) );
  NOR U561 ( .A(n456), .B(n455), .Z(n630) );
  IV U562 ( .A(n457), .Z(n458) );
  NOR U563 ( .A(n459), .B(n458), .Z(n463) );
  NOR U564 ( .A(n461), .B(n460), .Z(n462) );
  NOR U565 ( .A(n463), .B(n462), .Z(n627) );
  NOR U566 ( .A(n465), .B(n464), .Z(n470) );
  IV U567 ( .A(n466), .Z(n468) );
  NOR U568 ( .A(n468), .B(n467), .Z(n469) );
  NOR U569 ( .A(n470), .B(n469), .Z(n544) );
  NOR U570 ( .A(n472), .B(n471), .Z(n477) );
  IV U571 ( .A(n473), .Z(n475) );
  NOR U572 ( .A(n475), .B(n474), .Z(n476) );
  NOR U573 ( .A(n477), .B(n476), .Z(n541) );
  NOR U574 ( .A(n3749), .B(n3628), .Z(n512) );
  IV U575 ( .A(n512), .Z(n480) );
  IV U576 ( .A(n478), .Z(n479) );
  NOR U577 ( .A(n480), .B(n479), .Z(n485) );
  IV U578 ( .A(n481), .Z(n483) );
  NOR U579 ( .A(n483), .B(n482), .Z(n484) );
  NOR U580 ( .A(n485), .B(n484), .Z(n558) );
  IV U581 ( .A(n558), .Z(n492) );
  NOR U582 ( .A(n3781), .B(n3625), .Z(n521) );
  IV U583 ( .A(n521), .Z(n1511) );
  NOR U584 ( .A(n1511), .B(n486), .Z(n491) );
  IV U585 ( .A(n487), .Z(n489) );
  NOR U586 ( .A(n489), .B(n488), .Z(n490) );
  NOR U587 ( .A(n491), .B(n490), .Z(n557) );
  XOR U588 ( .A(n492), .B(n557), .Z(n560) );
  NOR U589 ( .A(n3062), .B(n3746), .Z(n923) );
  IV U590 ( .A(n923), .Z(n1038) );
  NOR U591 ( .A(n1038), .B(n493), .Z(n497) );
  IV U592 ( .A(n494), .Z(n1056) );
  NOR U593 ( .A(n1056), .B(n495), .Z(n496) );
  NOR U594 ( .A(n497), .B(n496), .Z(n565) );
  IV U595 ( .A(n498), .Z(n1861) );
  NOR U596 ( .A(n1861), .B(n499), .Z(n504) );
  IV U597 ( .A(n500), .Z(n501) );
  NOR U598 ( .A(n502), .B(n501), .Z(n503) );
  NOR U599 ( .A(n504), .B(n503), .Z(n564) );
  XOR U600 ( .A(n565), .B(n564), .Z(n505) );
  IV U601 ( .A(n505), .Z(n568) );
  NOR U602 ( .A(n3462), .B(n3650), .Z(n518) );
  IV U603 ( .A(n518), .Z(n507) );
  NOR U604 ( .A(n507), .B(n506), .Z(n511) );
  IV U605 ( .A(n508), .Z(n509) );
  NOR U606 ( .A(n1829), .B(n509), .Z(n510) );
  NOR U607 ( .A(n511), .B(n510), .Z(n575) );
  NOR U608 ( .A(n3647), .B(n3779), .Z(n513) );
  XOR U609 ( .A(n513), .B(n512), .Z(n588) );
  IV U610 ( .A(y[12]), .Z(n3688) );
  NOR U611 ( .A(n3688), .B(n3680), .Z(n514) );
  IV U612 ( .A(n514), .Z(n620) );
  NOR U613 ( .A(n3746), .B(n3682), .Z(n515) );
  IV U614 ( .A(x[12]), .Z(n3548) );
  NOR U615 ( .A(n3637), .B(n3548), .Z(n1358) );
  XOR U616 ( .A(n515), .B(n1358), .Z(n619) );
  XOR U617 ( .A(n620), .B(n619), .Z(n590) );
  XOR U618 ( .A(n588), .B(n590), .Z(n596) );
  NOR U619 ( .A(n3646), .B(n3635), .Z(n593) );
  NOR U620 ( .A(n3622), .B(n3619), .Z(n516) );
  XOR U621 ( .A(n517), .B(n516), .Z(n600) );
  NOR U622 ( .A(n3787), .B(n3765), .Z(n519) );
  XOR U623 ( .A(n519), .B(n518), .Z(n520) );
  IV U624 ( .A(n520), .Z(n607) );
  XOR U625 ( .A(n607), .B(n521), .Z(n602) );
  XOR U626 ( .A(n600), .B(n602), .Z(n594) );
  XOR U627 ( .A(n593), .B(n594), .Z(n595) );
  XOR U628 ( .A(n596), .B(n595), .Z(n571) );
  NOR U629 ( .A(n3740), .B(n3687), .Z(n579) );
  NOR U630 ( .A(n3062), .B(n3773), .Z(n522) );
  IV U631 ( .A(n522), .Z(n624) );
  XOR U632 ( .A(n624), .B(o[12]), .Z(n580) );
  XOR U633 ( .A(n579), .B(n580), .Z(n584) );
  IV U634 ( .A(o[11]), .Z(n523) );
  NOR U635 ( .A(n524), .B(n523), .Z(n582) );
  XOR U636 ( .A(n584), .B(n582), .Z(n572) );
  XOR U637 ( .A(n571), .B(n572), .Z(n574) );
  XOR U638 ( .A(n575), .B(n574), .Z(n566) );
  XOR U639 ( .A(n568), .B(n566), .Z(n559) );
  XOR U640 ( .A(n560), .B(n559), .Z(n553) );
  NOR U641 ( .A(n526), .B(n525), .Z(n531) );
  IV U642 ( .A(n527), .Z(n528) );
  NOR U643 ( .A(n529), .B(n528), .Z(n530) );
  NOR U644 ( .A(n531), .B(n530), .Z(n532) );
  IV U645 ( .A(n532), .Z(n551) );
  NOR U646 ( .A(n534), .B(n533), .Z(n539) );
  IV U647 ( .A(n535), .Z(n536) );
  NOR U648 ( .A(n537), .B(n536), .Z(n538) );
  NOR U649 ( .A(n539), .B(n538), .Z(n549) );
  XOR U650 ( .A(n551), .B(n549), .Z(n552) );
  XOR U651 ( .A(n553), .B(n552), .Z(n540) );
  IV U652 ( .A(n540), .Z(n543) );
  XOR U653 ( .A(n541), .B(n543), .Z(n546) );
  XOR U654 ( .A(n544), .B(n546), .Z(n629) );
  XOR U655 ( .A(n627), .B(n629), .Z(n632) );
  XOR U656 ( .A(n630), .B(n632), .Z(N45) );
  IV U657 ( .A(n541), .Z(n542) );
  NOR U658 ( .A(n543), .B(n542), .Z(n548) );
  IV U659 ( .A(n544), .Z(n545) );
  NOR U660 ( .A(n546), .B(n545), .Z(n547) );
  NOR U661 ( .A(n548), .B(n547), .Z(n636) );
  IV U662 ( .A(n549), .Z(n550) );
  NOR U663 ( .A(n551), .B(n550), .Z(n555) );
  NOR U664 ( .A(n553), .B(n552), .Z(n554) );
  NOR U665 ( .A(n555), .B(n554), .Z(n556) );
  IV U666 ( .A(n556), .Z(n647) );
  NOR U667 ( .A(n558), .B(n557), .Z(n562) );
  NOR U668 ( .A(n560), .B(n559), .Z(n561) );
  NOR U669 ( .A(n562), .B(n561), .Z(n563) );
  IV U670 ( .A(n563), .Z(n654) );
  NOR U671 ( .A(n565), .B(n564), .Z(n570) );
  IV U672 ( .A(n566), .Z(n567) );
  NOR U673 ( .A(n568), .B(n567), .Z(n569) );
  NOR U674 ( .A(n570), .B(n569), .Z(n650) );
  IV U675 ( .A(n571), .Z(n573) );
  NOR U676 ( .A(n573), .B(n572), .Z(n577) );
  NOR U677 ( .A(n575), .B(n574), .Z(n576) );
  NOR U678 ( .A(n577), .B(n576), .Z(n578) );
  IV U679 ( .A(n578), .Z(n651) );
  XOR U680 ( .A(n650), .B(n651), .Z(n653) );
  XOR U681 ( .A(n654), .B(n653), .Z(n644) );
  IV U682 ( .A(n579), .Z(n581) );
  NOR U683 ( .A(n581), .B(n580), .Z(n586) );
  IV U684 ( .A(n582), .Z(n583) );
  NOR U685 ( .A(n584), .B(n583), .Z(n585) );
  NOR U686 ( .A(n586), .B(n585), .Z(n658) );
  IV U687 ( .A(n587), .Z(n733) );
  NOR U688 ( .A(n772), .B(n733), .Z(n592) );
  IV U689 ( .A(n588), .Z(n589) );
  NOR U690 ( .A(n590), .B(n589), .Z(n591) );
  NOR U691 ( .A(n592), .B(n591), .Z(n657) );
  XOR U692 ( .A(n658), .B(n657), .Z(n659) );
  IV U693 ( .A(n593), .Z(n1333) );
  NOR U694 ( .A(n1333), .B(n594), .Z(n598) );
  NOR U695 ( .A(n596), .B(n595), .Z(n597) );
  NOR U696 ( .A(n598), .B(n597), .Z(n668) );
  NOR U697 ( .A(n3748), .B(n3622), .Z(n920) );
  IV U698 ( .A(n920), .Z(n599) );
  NOR U699 ( .A(n1155), .B(n599), .Z(n604) );
  IV U700 ( .A(n600), .Z(n601) );
  NOR U701 ( .A(n602), .B(n601), .Z(n603) );
  NOR U702 ( .A(n604), .B(n603), .Z(n665) );
  NOR U703 ( .A(n3765), .B(n3462), .Z(n1070) );
  IV U704 ( .A(n1070), .Z(n606) );
  IV U705 ( .A(n605), .Z(n1037) );
  NOR U706 ( .A(n606), .B(n1037), .Z(n609) );
  NOR U707 ( .A(n1511), .B(n607), .Z(n608) );
  NOR U708 ( .A(n609), .B(n608), .Z(n682) );
  NOR U709 ( .A(n3647), .B(n3062), .Z(n611) );
  NOR U710 ( .A(n3746), .B(n3749), .Z(n610) );
  XOR U711 ( .A(n611), .B(n610), .Z(n734) );
  IV U712 ( .A(y[13]), .Z(n3763) );
  NOR U713 ( .A(n3763), .B(n3680), .Z(n613) );
  NOR U714 ( .A(n3462), .B(n3740), .Z(n612) );
  XOR U715 ( .A(n613), .B(n612), .Z(n614) );
  IV U716 ( .A(n614), .Z(n700) );
  IV U717 ( .A(x[13]), .Z(n3546) );
  NOR U718 ( .A(n3546), .B(n3637), .Z(n699) );
  XOR U719 ( .A(n700), .B(n699), .Z(n735) );
  XOR U720 ( .A(n734), .B(n735), .Z(n679) );
  NOR U721 ( .A(n3650), .B(n3646), .Z(n615) );
  NOR U722 ( .A(n3787), .B(n3779), .Z(n1297) );
  XOR U723 ( .A(n615), .B(n1297), .Z(n692) );
  NOR U724 ( .A(n3622), .B(n3635), .Z(n1606) );
  NOR U725 ( .A(n3628), .B(n3765), .Z(n1822) );
  XOR U726 ( .A(n1606), .B(n1822), .Z(n686) );
  NOR U727 ( .A(n3688), .B(n3625), .Z(n616) );
  XOR U728 ( .A(n617), .B(n616), .Z(n618) );
  IV U729 ( .A(n618), .Z(n715) );
  NOR U730 ( .A(n3781), .B(n3619), .Z(n714) );
  XOR U731 ( .A(n715), .B(n714), .Z(n688) );
  XOR U732 ( .A(n686), .B(n688), .Z(n694) );
  XOR U733 ( .A(n692), .B(n694), .Z(n678) );
  XOR U734 ( .A(n679), .B(n678), .Z(n680) );
  XOR U735 ( .A(n682), .B(n680), .Z(n675) );
  NOR U736 ( .A(n3746), .B(n3548), .Z(n1069) );
  IV U737 ( .A(n1069), .Z(n784) );
  NOR U738 ( .A(n784), .B(n820), .Z(n623) );
  IV U739 ( .A(n619), .Z(n621) );
  NOR U740 ( .A(n621), .B(n620), .Z(n622) );
  NOR U741 ( .A(n623), .B(n622), .Z(n672) );
  IV U742 ( .A(o[12]), .Z(n625) );
  NOR U743 ( .A(n625), .B(n624), .Z(n706) );
  NOR U744 ( .A(n3748), .B(n3687), .Z(n703) );
  NOR U745 ( .A(n3773), .B(n3548), .Z(n626) );
  IV U746 ( .A(n626), .Z(n728) );
  XOR U747 ( .A(n728), .B(o[13]), .Z(n705) );
  XOR U748 ( .A(n703), .B(n705), .Z(n708) );
  XOR U749 ( .A(n706), .B(n708), .Z(n671) );
  XOR U750 ( .A(n672), .B(n671), .Z(n673) );
  XOR U751 ( .A(n675), .B(n673), .Z(n664) );
  XOR U752 ( .A(n665), .B(n664), .Z(n666) );
  XOR U753 ( .A(n668), .B(n666), .Z(n661) );
  XOR U754 ( .A(n659), .B(n661), .Z(n643) );
  XOR U755 ( .A(n644), .B(n643), .Z(n645) );
  XOR U756 ( .A(n647), .B(n645), .Z(n638) );
  XOR U757 ( .A(n636), .B(n638), .Z(n640) );
  IV U758 ( .A(n627), .Z(n628) );
  NOR U759 ( .A(n629), .B(n628), .Z(n634) );
  IV U760 ( .A(n630), .Z(n631) );
  NOR U761 ( .A(n632), .B(n631), .Z(n633) );
  NOR U762 ( .A(n634), .B(n633), .Z(n635) );
  IV U763 ( .A(n635), .Z(n639) );
  XOR U764 ( .A(n640), .B(n639), .Z(N46) );
  IV U765 ( .A(n636), .Z(n637) );
  NOR U766 ( .A(n638), .B(n637), .Z(n642) );
  NOR U767 ( .A(n640), .B(n639), .Z(n641) );
  NOR U768 ( .A(n642), .B(n641), .Z(n846) );
  NOR U769 ( .A(n644), .B(n643), .Z(n649) );
  IV U770 ( .A(n645), .Z(n646) );
  NOR U771 ( .A(n647), .B(n646), .Z(n648) );
  NOR U772 ( .A(n649), .B(n648), .Z(n843) );
  IV U773 ( .A(n650), .Z(n652) );
  NOR U774 ( .A(n652), .B(n651), .Z(n656) );
  NOR U775 ( .A(n654), .B(n653), .Z(n655) );
  NOR U776 ( .A(n656), .B(n655), .Z(n744) );
  IV U777 ( .A(n744), .Z(n739) );
  NOR U778 ( .A(n658), .B(n657), .Z(n663) );
  IV U779 ( .A(n659), .Z(n660) );
  NOR U780 ( .A(n661), .B(n660), .Z(n662) );
  NOR U781 ( .A(n663), .B(n662), .Z(n740) );
  NOR U782 ( .A(n665), .B(n664), .Z(n670) );
  IV U783 ( .A(n666), .Z(n667) );
  NOR U784 ( .A(n668), .B(n667), .Z(n669) );
  NOR U785 ( .A(n670), .B(n669), .Z(n750) );
  NOR U786 ( .A(n672), .B(n671), .Z(n677) );
  IV U787 ( .A(n673), .Z(n674) );
  NOR U788 ( .A(n675), .B(n674), .Z(n676) );
  NOR U789 ( .A(n677), .B(n676), .Z(n747) );
  NOR U790 ( .A(n679), .B(n678), .Z(n684) );
  IV U791 ( .A(n680), .Z(n681) );
  NOR U792 ( .A(n682), .B(n681), .Z(n683) );
  NOR U793 ( .A(n684), .B(n683), .Z(n685) );
  IV U794 ( .A(n685), .Z(n757) );
  NOR U795 ( .A(n3765), .B(n3622), .Z(n1391) );
  IV U796 ( .A(n1391), .Z(n1503) );
  NOR U797 ( .A(n1503), .B(n1072), .Z(n690) );
  IV U798 ( .A(n686), .Z(n687) );
  NOR U799 ( .A(n688), .B(n687), .Z(n689) );
  NOR U800 ( .A(n690), .B(n689), .Z(n755) );
  XOR U801 ( .A(n757), .B(n755), .Z(n760) );
  NOR U802 ( .A(n3646), .B(n3779), .Z(n691) );
  IV U803 ( .A(n691), .Z(n1386) );
  NOR U804 ( .A(n1386), .B(n1037), .Z(n696) );
  IV U805 ( .A(n692), .Z(n693) );
  NOR U806 ( .A(n694), .B(n693), .Z(n695) );
  NOR U807 ( .A(n696), .B(n695), .Z(n833) );
  IV U808 ( .A(n697), .Z(n1476) );
  NOR U809 ( .A(n3763), .B(n3740), .Z(n1169) );
  IV U810 ( .A(n1169), .Z(n698) );
  NOR U811 ( .A(n1476), .B(n698), .Z(n702) );
  IV U812 ( .A(n699), .Z(n1162) );
  NOR U813 ( .A(n1162), .B(n700), .Z(n701) );
  NOR U814 ( .A(n702), .B(n701), .Z(n831) );
  IV U815 ( .A(n831), .Z(n711) );
  IV U816 ( .A(n703), .Z(n704) );
  NOR U817 ( .A(n705), .B(n704), .Z(n710) );
  IV U818 ( .A(n706), .Z(n707) );
  NOR U819 ( .A(n708), .B(n707), .Z(n709) );
  NOR U820 ( .A(n710), .B(n709), .Z(n830) );
  XOR U821 ( .A(n711), .B(n830), .Z(n832) );
  XOR U822 ( .A(n833), .B(n832), .Z(n840) );
  NOR U823 ( .A(n3682), .B(n3688), .Z(n1344) );
  IV U824 ( .A(n1344), .Z(n713) );
  IV U825 ( .A(n712), .Z(n1022) );
  NOR U826 ( .A(n713), .B(n1022), .Z(n717) );
  IV U827 ( .A(n714), .Z(n813) );
  NOR U828 ( .A(n813), .B(n715), .Z(n716) );
  NOR U829 ( .A(n717), .B(n716), .Z(n766) );
  NOR U830 ( .A(n3763), .B(n3625), .Z(n1613) );
  NOR U831 ( .A(n3650), .B(n3622), .Z(n718) );
  XOR U832 ( .A(n1613), .B(n718), .Z(n792) );
  NOR U833 ( .A(n3787), .B(n3062), .Z(n720) );
  XOR U834 ( .A(n720), .B(n719), .Z(n721) );
  IV U835 ( .A(n721), .Z(n773) );
  XOR U836 ( .A(n773), .B(n722), .Z(n794) );
  XOR U837 ( .A(n792), .B(n794), .Z(n764) );
  NOR U838 ( .A(n3746), .B(n3765), .Z(n1147) );
  NOR U839 ( .A(n3548), .B(n3647), .Z(n1451) );
  XOR U840 ( .A(n1147), .B(n1451), .Z(n785) );
  IV U841 ( .A(y[14]), .Z(n3467) );
  NOR U842 ( .A(n3680), .B(n3467), .Z(n723) );
  IV U843 ( .A(n723), .Z(n822) );
  NOR U844 ( .A(n3687), .B(n3682), .Z(n724) );
  IV U845 ( .A(x[14]), .Z(n3776) );
  NOR U846 ( .A(n3776), .B(n3637), .Z(n1807) );
  XOR U847 ( .A(n724), .B(n1807), .Z(n821) );
  XOR U848 ( .A(n822), .B(n821), .Z(n787) );
  XOR U849 ( .A(n785), .B(n787), .Z(n802) );
  NOR U850 ( .A(n3749), .B(n3633), .Z(n725) );
  IV U851 ( .A(n725), .Z(n816) );
  NOR U852 ( .A(n3619), .B(n3688), .Z(n727) );
  NOR U853 ( .A(n3635), .B(n3781), .Z(n726) );
  XOR U854 ( .A(n727), .B(n726), .Z(n815) );
  XOR U855 ( .A(n816), .B(n815), .Z(n799) );
  IV U856 ( .A(o[13]), .Z(n729) );
  NOR U857 ( .A(n729), .B(n728), .Z(n807) );
  NOR U858 ( .A(n3773), .B(n3546), .Z(n730) );
  IV U859 ( .A(n730), .Z(n827) );
  XOR U860 ( .A(n827), .B(o[14]), .Z(n805) );
  XOR U861 ( .A(n731), .B(n805), .Z(n809) );
  XOR U862 ( .A(n807), .B(n809), .Z(n798) );
  XOR U863 ( .A(n799), .B(n798), .Z(n800) );
  XOR U864 ( .A(n802), .B(n800), .Z(n763) );
  XOR U865 ( .A(n764), .B(n763), .Z(n732) );
  IV U866 ( .A(n732), .Z(n765) );
  XOR U867 ( .A(n766), .B(n765), .Z(n838) );
  NOR U868 ( .A(n1038), .B(n733), .Z(n738) );
  IV U869 ( .A(n734), .Z(n736) );
  NOR U870 ( .A(n736), .B(n735), .Z(n737) );
  NOR U871 ( .A(n738), .B(n737), .Z(n836) );
  XOR U872 ( .A(n838), .B(n836), .Z(n839) );
  XOR U873 ( .A(n840), .B(n839), .Z(n758) );
  XOR U874 ( .A(n760), .B(n758), .Z(n749) );
  XOR U875 ( .A(n747), .B(n749), .Z(n752) );
  XOR U876 ( .A(n750), .B(n752), .Z(n741) );
  XOR U877 ( .A(n740), .B(n741), .Z(n743) );
  XOR U878 ( .A(n739), .B(n743), .Z(n845) );
  XOR U879 ( .A(n843), .B(n845), .Z(n848) );
  XOR U880 ( .A(n846), .B(n848), .Z(N47) );
  IV U881 ( .A(n740), .Z(n742) );
  NOR U882 ( .A(n742), .B(n741), .Z(n746) );
  NOR U883 ( .A(n744), .B(n743), .Z(n745) );
  NOR U884 ( .A(n746), .B(n745), .Z(n852) );
  IV U885 ( .A(n747), .Z(n748) );
  NOR U886 ( .A(n749), .B(n748), .Z(n754) );
  IV U887 ( .A(n750), .Z(n751) );
  NOR U888 ( .A(n752), .B(n751), .Z(n753) );
  NOR U889 ( .A(n754), .B(n753), .Z(n862) );
  IV U890 ( .A(n755), .Z(n756) );
  NOR U891 ( .A(n757), .B(n756), .Z(n762) );
  IV U892 ( .A(n758), .Z(n759) );
  NOR U893 ( .A(n760), .B(n759), .Z(n761) );
  NOR U894 ( .A(n762), .B(n761), .Z(n859) );
  NOR U895 ( .A(n764), .B(n763), .Z(n768) );
  NOR U896 ( .A(n766), .B(n765), .Z(n767) );
  NOR U897 ( .A(n768), .B(n767), .Z(n878) );
  NOR U898 ( .A(n3062), .B(n3646), .Z(n1465) );
  IV U899 ( .A(n1465), .Z(n771) );
  IV U900 ( .A(n769), .Z(n770) );
  NOR U901 ( .A(n771), .B(n770), .Z(n775) );
  NOR U902 ( .A(n773), .B(n772), .Z(n774) );
  NOR U903 ( .A(n775), .B(n774), .Z(n970) );
  NOR U904 ( .A(n3746), .B(n3779), .Z(n776) );
  NOR U905 ( .A(n3763), .B(n3619), .Z(n2056) );
  XOR U906 ( .A(n776), .B(n2056), .Z(n904) );
  NOR U907 ( .A(n3467), .B(n3625), .Z(n777) );
  IV U908 ( .A(n777), .Z(n952) );
  NOR U909 ( .A(n3687), .B(n3749), .Z(n779) );
  IV U910 ( .A(y[15]), .Z(n3741) );
  NOR U911 ( .A(n3680), .B(n3741), .Z(n778) );
  XOR U912 ( .A(n779), .B(n778), .Z(n951) );
  XOR U913 ( .A(n952), .B(n951), .Z(n906) );
  XOR U914 ( .A(n904), .B(n906), .Z(n968) );
  NOR U915 ( .A(n3647), .B(n3546), .Z(n2041) );
  NOR U916 ( .A(n3765), .B(n3633), .Z(n2198) );
  XOR U917 ( .A(n2041), .B(n2198), .Z(n909) );
  NOR U918 ( .A(n3688), .B(n3635), .Z(n812) );
  NOR U919 ( .A(n3548), .B(n3787), .Z(n780) );
  XOR U920 ( .A(n812), .B(n780), .Z(n781) );
  IV U921 ( .A(n781), .Z(n946) );
  IV U922 ( .A(x[15]), .Z(n3465) );
  NOR U923 ( .A(n3465), .B(n3637), .Z(n945) );
  XOR U924 ( .A(n946), .B(n945), .Z(n911) );
  XOR U925 ( .A(n909), .B(n911), .Z(n941) );
  NOR U926 ( .A(n3646), .B(n3748), .Z(n937) );
  NOR U927 ( .A(n3628), .B(n3062), .Z(n782) );
  NOR U928 ( .A(n3781), .B(n3650), .Z(n1310) );
  XOR U929 ( .A(n782), .B(n1310), .Z(n783) );
  IV U930 ( .A(n783), .Z(n917) );
  NOR U931 ( .A(n3740), .B(n3622), .Z(n916) );
  XOR U932 ( .A(n917), .B(n916), .Z(n939) );
  XOR U933 ( .A(n937), .B(n939), .Z(n940) );
  XOR U934 ( .A(n941), .B(n940), .Z(n966) );
  XOR U935 ( .A(n968), .B(n966), .Z(n969) );
  XOR U936 ( .A(n970), .B(n969), .Z(n898) );
  NOR U937 ( .A(n784), .B(n1056), .Z(n789) );
  IV U938 ( .A(n785), .Z(n786) );
  NOR U939 ( .A(n787), .B(n786), .Z(n788) );
  NOR U940 ( .A(n789), .B(n788), .Z(n896) );
  XOR U941 ( .A(n898), .B(n896), .Z(n900) );
  NOR U942 ( .A(n3763), .B(n3650), .Z(n1071) );
  IV U943 ( .A(n1071), .Z(n1203) );
  IV U944 ( .A(n790), .Z(n791) );
  NOR U945 ( .A(n1203), .B(n791), .Z(n796) );
  IV U946 ( .A(n792), .Z(n793) );
  NOR U947 ( .A(n794), .B(n793), .Z(n795) );
  NOR U948 ( .A(n796), .B(n795), .Z(n797) );
  IV U949 ( .A(n797), .Z(n899) );
  XOR U950 ( .A(n900), .B(n899), .Z(n876) );
  NOR U951 ( .A(n799), .B(n798), .Z(n804) );
  IV U952 ( .A(n800), .Z(n801) );
  NOR U953 ( .A(n802), .B(n801), .Z(n803) );
  NOR U954 ( .A(n804), .B(n803), .Z(n885) );
  NOR U955 ( .A(n806), .B(n805), .Z(n811) );
  IV U956 ( .A(n807), .Z(n808) );
  NOR U957 ( .A(n809), .B(n808), .Z(n810) );
  NOR U958 ( .A(n811), .B(n810), .Z(n882) );
  IV U959 ( .A(n812), .Z(n814) );
  NOR U960 ( .A(n814), .B(n813), .Z(n819) );
  IV U961 ( .A(n815), .Z(n817) );
  NOR U962 ( .A(n817), .B(n816), .Z(n818) );
  NOR U963 ( .A(n819), .B(n818), .Z(n893) );
  NOR U964 ( .A(n3776), .B(n3687), .Z(n1626) );
  IV U965 ( .A(n1626), .Z(n1057) );
  NOR U966 ( .A(n1057), .B(n820), .Z(n825) );
  IV U967 ( .A(n821), .Z(n823) );
  NOR U968 ( .A(n823), .B(n822), .Z(n824) );
  NOR U969 ( .A(n825), .B(n824), .Z(n890) );
  IV U970 ( .A(o[14]), .Z(n826) );
  NOR U971 ( .A(n827), .B(n826), .Z(n932) );
  NOR U972 ( .A(n3682), .B(n3462), .Z(n929) );
  NOR U973 ( .A(n3773), .B(n3776), .Z(n828) );
  IV U974 ( .A(n828), .Z(n924) );
  XOR U975 ( .A(n924), .B(o[15]), .Z(n931) );
  XOR U976 ( .A(n929), .B(n931), .Z(n934) );
  XOR U977 ( .A(n932), .B(n934), .Z(n889) );
  XOR U978 ( .A(n890), .B(n889), .Z(n891) );
  XOR U979 ( .A(n893), .B(n891), .Z(n881) );
  XOR U980 ( .A(n882), .B(n881), .Z(n883) );
  XOR U981 ( .A(n885), .B(n883), .Z(n875) );
  XOR U982 ( .A(n876), .B(n875), .Z(n829) );
  IV U983 ( .A(n829), .Z(n877) );
  XOR U984 ( .A(n878), .B(n877), .Z(n870) );
  NOR U985 ( .A(n831), .B(n830), .Z(n835) );
  NOR U986 ( .A(n833), .B(n832), .Z(n834) );
  NOR U987 ( .A(n835), .B(n834), .Z(n869) );
  IV U988 ( .A(n836), .Z(n837) );
  NOR U989 ( .A(n838), .B(n837), .Z(n842) );
  NOR U990 ( .A(n840), .B(n839), .Z(n841) );
  NOR U991 ( .A(n842), .B(n841), .Z(n867) );
  XOR U992 ( .A(n869), .B(n867), .Z(n871) );
  XOR U993 ( .A(n870), .B(n871), .Z(n861) );
  XOR U994 ( .A(n859), .B(n861), .Z(n863) );
  XOR U995 ( .A(n862), .B(n863), .Z(n854) );
  XOR U996 ( .A(n852), .B(n854), .Z(n856) );
  IV U997 ( .A(n843), .Z(n844) );
  NOR U998 ( .A(n845), .B(n844), .Z(n850) );
  IV U999 ( .A(n846), .Z(n847) );
  NOR U1000 ( .A(n848), .B(n847), .Z(n849) );
  NOR U1001 ( .A(n850), .B(n849), .Z(n851) );
  IV U1002 ( .A(n851), .Z(n855) );
  XOR U1003 ( .A(n856), .B(n855), .Z(N48) );
  IV U1004 ( .A(n852), .Z(n853) );
  NOR U1005 ( .A(n854), .B(n853), .Z(n858) );
  NOR U1006 ( .A(n856), .B(n855), .Z(n857) );
  NOR U1007 ( .A(n858), .B(n857), .Z(n1098) );
  IV U1008 ( .A(n859), .Z(n860) );
  NOR U1009 ( .A(n861), .B(n860), .Z(n866) );
  IV U1010 ( .A(n862), .Z(n864) );
  NOR U1011 ( .A(n864), .B(n863), .Z(n865) );
  NOR U1012 ( .A(n866), .B(n865), .Z(n1095) );
  IV U1013 ( .A(n867), .Z(n868) );
  NOR U1014 ( .A(n869), .B(n868), .Z(n874) );
  IV U1015 ( .A(n870), .Z(n872) );
  NOR U1016 ( .A(n872), .B(n871), .Z(n873) );
  NOR U1017 ( .A(n874), .B(n873), .Z(n976) );
  NOR U1018 ( .A(n876), .B(n875), .Z(n880) );
  NOR U1019 ( .A(n878), .B(n877), .Z(n879) );
  NOR U1020 ( .A(n880), .B(n879), .Z(n973) );
  NOR U1021 ( .A(n882), .B(n881), .Z(n887) );
  IV U1022 ( .A(n883), .Z(n884) );
  NOR U1023 ( .A(n885), .B(n884), .Z(n886) );
  NOR U1024 ( .A(n887), .B(n886), .Z(n888) );
  IV U1025 ( .A(n888), .Z(n983) );
  NOR U1026 ( .A(n890), .B(n889), .Z(n895) );
  IV U1027 ( .A(n891), .Z(n892) );
  NOR U1028 ( .A(n893), .B(n892), .Z(n894) );
  NOR U1029 ( .A(n895), .B(n894), .Z(n981) );
  XOR U1030 ( .A(n983), .B(n981), .Z(n986) );
  IV U1031 ( .A(n896), .Z(n897) );
  NOR U1032 ( .A(n898), .B(n897), .Z(n902) );
  NOR U1033 ( .A(n900), .B(n899), .Z(n901) );
  NOR U1034 ( .A(n902), .B(n901), .Z(n993) );
  NOR U1035 ( .A(n3779), .B(n3763), .Z(n2055) );
  IV U1036 ( .A(n2055), .Z(n2240) );
  IV U1037 ( .A(n903), .Z(n1305) );
  NOR U1038 ( .A(n2240), .B(n1305), .Z(n908) );
  IV U1039 ( .A(n904), .Z(n905) );
  NOR U1040 ( .A(n906), .B(n905), .Z(n907) );
  NOR U1041 ( .A(n908), .B(n907), .Z(n997) );
  NOR U1042 ( .A(n3633), .B(n3546), .Z(n1349) );
  IV U1043 ( .A(n1349), .Z(n1500) );
  NOR U1044 ( .A(n1500), .B(n1056), .Z(n913) );
  IV U1045 ( .A(n909), .Z(n910) );
  NOR U1046 ( .A(n911), .B(n910), .Z(n912) );
  NOR U1047 ( .A(n913), .B(n912), .Z(n996) );
  XOR U1048 ( .A(n997), .B(n996), .Z(n914) );
  IV U1049 ( .A(n914), .Z(n998) );
  NOR U1050 ( .A(n3062), .B(n3781), .Z(n1845) );
  IV U1051 ( .A(n1845), .Z(n1989) );
  NOR U1052 ( .A(n1989), .B(n915), .Z(n919) );
  IV U1053 ( .A(n916), .Z(n1086) );
  NOR U1054 ( .A(n1086), .B(n917), .Z(n918) );
  NOR U1055 ( .A(n919), .B(n918), .Z(n1012) );
  NOR U1056 ( .A(n3740), .B(n3781), .Z(n1218) );
  XOR U1057 ( .A(n1218), .B(n920), .Z(n1088) );
  NOR U1058 ( .A(n3650), .B(n3688), .Z(n1482) );
  NOR U1059 ( .A(n3787), .B(n3546), .Z(n921) );
  XOR U1060 ( .A(n1482), .B(n921), .Z(n922) );
  IV U1061 ( .A(n922), .Z(n1039) );
  XOR U1062 ( .A(n1039), .B(n923), .Z(n1089) );
  XOR U1063 ( .A(n1088), .B(n1089), .Z(n1010) );
  IV U1064 ( .A(o[15]), .Z(n925) );
  NOR U1065 ( .A(n925), .B(n924), .Z(n1017) );
  NOR U1066 ( .A(n3465), .B(n3773), .Z(n926) );
  IV U1067 ( .A(n926), .Z(n1033) );
  XOR U1068 ( .A(n1033), .B(o[16]), .Z(n1016) );
  XOR U1069 ( .A(n927), .B(n1016), .Z(n1019) );
  XOR U1070 ( .A(n1017), .B(n1019), .Z(n1009) );
  XOR U1071 ( .A(n1010), .B(n1009), .Z(n928) );
  IV U1072 ( .A(n928), .Z(n1011) );
  XOR U1073 ( .A(n1012), .B(n1011), .Z(n1004) );
  IV U1074 ( .A(n929), .Z(n930) );
  NOR U1075 ( .A(n931), .B(n930), .Z(n936) );
  IV U1076 ( .A(n932), .Z(n933) );
  NOR U1077 ( .A(n934), .B(n933), .Z(n935) );
  NOR U1078 ( .A(n936), .B(n935), .Z(n1002) );
  XOR U1079 ( .A(n1004), .B(n1002), .Z(n1005) );
  IV U1080 ( .A(n937), .Z(n938) );
  NOR U1081 ( .A(n939), .B(n938), .Z(n943) );
  NOR U1082 ( .A(n941), .B(n940), .Z(n942) );
  NOR U1083 ( .A(n943), .B(n942), .Z(n1053) );
  NOR U1084 ( .A(n3688), .B(n3548), .Z(n2222) );
  IV U1085 ( .A(n2222), .Z(n2323) );
  NOR U1086 ( .A(n2323), .B(n944), .Z(n948) );
  IV U1087 ( .A(n945), .Z(n2148) );
  NOR U1088 ( .A(n2148), .B(n946), .Z(n947) );
  NOR U1089 ( .A(n948), .B(n947), .Z(n1051) );
  NOR U1090 ( .A(n3749), .B(n3741), .Z(n2027) );
  IV U1091 ( .A(n2027), .Z(n950) );
  IV U1092 ( .A(n949), .Z(n1352) );
  NOR U1093 ( .A(n950), .B(n1352), .Z(n955) );
  IV U1094 ( .A(n951), .Z(n953) );
  NOR U1095 ( .A(n953), .B(n952), .Z(n954) );
  NOR U1096 ( .A(n955), .B(n954), .Z(n1046) );
  NOR U1097 ( .A(n3548), .B(n3628), .Z(n957) );
  NOR U1098 ( .A(n3763), .B(n3635), .Z(n956) );
  XOR U1099 ( .A(n957), .B(n956), .Z(n1074) );
  NOR U1100 ( .A(n3467), .B(n3619), .Z(n958) );
  IV U1101 ( .A(n958), .Z(n1024) );
  NOR U1102 ( .A(n3779), .B(n3633), .Z(n960) );
  NOR U1103 ( .A(n3741), .B(n3625), .Z(n959) );
  XOR U1104 ( .A(n960), .B(n959), .Z(n1023) );
  XOR U1105 ( .A(n1024), .B(n1023), .Z(n1076) );
  XOR U1106 ( .A(n1074), .B(n1076), .Z(n1043) );
  NOR U1107 ( .A(n3687), .B(n3765), .Z(n961) );
  NOR U1108 ( .A(n3776), .B(n3647), .Z(n1210) );
  XOR U1109 ( .A(n961), .B(n1210), .Z(n1058) );
  IV U1110 ( .A(x[16]), .Z(n3742) );
  NOR U1111 ( .A(n3742), .B(n3637), .Z(n962) );
  IV U1112 ( .A(n962), .Z(n1081) );
  IV U1113 ( .A(y[16]), .Z(n2764) );
  NOR U1114 ( .A(n3680), .B(n2764), .Z(n964) );
  XOR U1115 ( .A(n964), .B(n963), .Z(n1080) );
  XOR U1116 ( .A(n1081), .B(n1080), .Z(n1059) );
  XOR U1117 ( .A(n1058), .B(n1059), .Z(n1042) );
  XOR U1118 ( .A(n1043), .B(n1042), .Z(n1044) );
  XOR U1119 ( .A(n1046), .B(n1044), .Z(n1050) );
  XOR U1120 ( .A(n1051), .B(n1050), .Z(n965) );
  IV U1121 ( .A(n965), .Z(n1052) );
  XOR U1122 ( .A(n1053), .B(n1052), .Z(n1006) );
  XOR U1123 ( .A(n1005), .B(n1006), .Z(n999) );
  XOR U1124 ( .A(n998), .B(n999), .Z(n991) );
  IV U1125 ( .A(n966), .Z(n967) );
  NOR U1126 ( .A(n968), .B(n967), .Z(n972) );
  NOR U1127 ( .A(n970), .B(n969), .Z(n971) );
  NOR U1128 ( .A(n972), .B(n971), .Z(n989) );
  XOR U1129 ( .A(n991), .B(n989), .Z(n992) );
  XOR U1130 ( .A(n993), .B(n992), .Z(n984) );
  XOR U1131 ( .A(n986), .B(n984), .Z(n975) );
  XOR U1132 ( .A(n973), .B(n975), .Z(n978) );
  XOR U1133 ( .A(n976), .B(n978), .Z(n1097) );
  XOR U1134 ( .A(n1095), .B(n1097), .Z(n1100) );
  XOR U1135 ( .A(n1098), .B(n1100), .Z(N49) );
  IV U1136 ( .A(n973), .Z(n974) );
  NOR U1137 ( .A(n975), .B(n974), .Z(n980) );
  IV U1138 ( .A(n976), .Z(n977) );
  NOR U1139 ( .A(n978), .B(n977), .Z(n979) );
  NOR U1140 ( .A(n980), .B(n979), .Z(n1104) );
  IV U1141 ( .A(n981), .Z(n982) );
  NOR U1142 ( .A(n983), .B(n982), .Z(n988) );
  IV U1143 ( .A(n984), .Z(n985) );
  NOR U1144 ( .A(n986), .B(n985), .Z(n987) );
  NOR U1145 ( .A(n988), .B(n987), .Z(n1114) );
  IV U1146 ( .A(n989), .Z(n990) );
  NOR U1147 ( .A(n991), .B(n990), .Z(n995) );
  NOR U1148 ( .A(n993), .B(n992), .Z(n994) );
  NOR U1149 ( .A(n995), .B(n994), .Z(n1111) );
  NOR U1150 ( .A(n997), .B(n996), .Z(n1001) );
  NOR U1151 ( .A(n999), .B(n998), .Z(n1000) );
  NOR U1152 ( .A(n1001), .B(n1000), .Z(n1123) );
  IV U1153 ( .A(n1123), .Z(n1094) );
  IV U1154 ( .A(n1002), .Z(n1003) );
  NOR U1155 ( .A(n1004), .B(n1003), .Z(n1008) );
  NOR U1156 ( .A(n1006), .B(n1005), .Z(n1007) );
  NOR U1157 ( .A(n1008), .B(n1007), .Z(n1119) );
  NOR U1158 ( .A(n1010), .B(n1009), .Z(n1014) );
  NOR U1159 ( .A(n1012), .B(n1011), .Z(n1013) );
  NOR U1160 ( .A(n1014), .B(n1013), .Z(n1233) );
  NOR U1161 ( .A(n1016), .B(n1015), .Z(n1021) );
  IV U1162 ( .A(n1017), .Z(n1018) );
  NOR U1163 ( .A(n1019), .B(n1018), .Z(n1020) );
  NOR U1164 ( .A(n1021), .B(n1020), .Z(n1198) );
  NOR U1165 ( .A(n3779), .B(n3741), .Z(n2436) );
  IV U1166 ( .A(n2436), .Z(n2551) );
  NOR U1167 ( .A(n2551), .B(n1022), .Z(n1027) );
  IV U1168 ( .A(n1023), .Z(n1025) );
  NOR U1169 ( .A(n1025), .B(n1024), .Z(n1026) );
  NOR U1170 ( .A(n1027), .B(n1026), .Z(n1230) );
  NOR U1171 ( .A(n3633), .B(n3062), .Z(n1029) );
  NOR U1172 ( .A(n3741), .B(n3619), .Z(n1028) );
  XOR U1173 ( .A(n1029), .B(n1028), .Z(n1156) );
  NOR U1174 ( .A(n2764), .B(n3625), .Z(n1030) );
  IV U1175 ( .A(n1030), .Z(n1134) );
  IV U1176 ( .A(y[17]), .Z(n3775) );
  NOR U1177 ( .A(n3680), .B(n3775), .Z(n1032) );
  NOR U1178 ( .A(n3779), .B(n3687), .Z(n1031) );
  XOR U1179 ( .A(n1032), .B(n1031), .Z(n1133) );
  XOR U1180 ( .A(n1134), .B(n1133), .Z(n1158) );
  XOR U1181 ( .A(n1156), .B(n1158), .Z(n1228) );
  IV U1182 ( .A(o[16]), .Z(n1034) );
  NOR U1183 ( .A(n1034), .B(n1033), .Z(n1182) );
  NOR U1184 ( .A(n3749), .B(n3646), .Z(n1179) );
  NOR U1185 ( .A(n3773), .B(n3742), .Z(n1035) );
  IV U1186 ( .A(n1035), .Z(n1175) );
  XOR U1187 ( .A(n1175), .B(o[17]), .Z(n1181) );
  XOR U1188 ( .A(n1179), .B(n1181), .Z(n1184) );
  XOR U1189 ( .A(n1182), .B(n1184), .Z(n1227) );
  XOR U1190 ( .A(n1228), .B(n1227), .Z(n1036) );
  IV U1191 ( .A(n1036), .Z(n1229) );
  XOR U1192 ( .A(n1230), .B(n1229), .Z(n1197) );
  NOR U1193 ( .A(n3688), .B(n3546), .Z(n2431) );
  IV U1194 ( .A(n2431), .Z(n2594) );
  NOR U1195 ( .A(n2594), .B(n1037), .Z(n1041) );
  NOR U1196 ( .A(n1039), .B(n1038), .Z(n1040) );
  NOR U1197 ( .A(n1041), .B(n1040), .Z(n1195) );
  XOR U1198 ( .A(n1197), .B(n1195), .Z(n1200) );
  XOR U1199 ( .A(n1198), .B(n1200), .Z(n1235) );
  XOR U1200 ( .A(n1233), .B(n1235), .Z(n1237) );
  NOR U1201 ( .A(n1043), .B(n1042), .Z(n1048) );
  IV U1202 ( .A(n1044), .Z(n1045) );
  NOR U1203 ( .A(n1046), .B(n1045), .Z(n1047) );
  NOR U1204 ( .A(n1048), .B(n1047), .Z(n1049) );
  IV U1205 ( .A(n1049), .Z(n1236) );
  XOR U1206 ( .A(n1237), .B(n1236), .Z(n1245) );
  IV U1207 ( .A(n1245), .Z(n1093) );
  NOR U1208 ( .A(n1051), .B(n1050), .Z(n1055) );
  NOR U1209 ( .A(n1053), .B(n1052), .Z(n1054) );
  NOR U1210 ( .A(n1055), .B(n1054), .Z(n1243) );
  NOR U1211 ( .A(n1057), .B(n1056), .Z(n1062) );
  IV U1212 ( .A(n1058), .Z(n1060) );
  NOR U1213 ( .A(n1060), .B(n1059), .Z(n1061) );
  NOR U1214 ( .A(n1062), .B(n1061), .Z(n1190) );
  NOR U1215 ( .A(n3647), .B(n3465), .Z(n1064) );
  NOR U1216 ( .A(n3787), .B(n3776), .Z(n1063) );
  XOR U1217 ( .A(n1064), .B(n1063), .Z(n1212) );
  NOR U1218 ( .A(n3467), .B(n3635), .Z(n1065) );
  IV U1219 ( .A(n1065), .Z(n1165) );
  IV U1220 ( .A(x[17]), .Z(n3529) );
  NOR U1221 ( .A(n3637), .B(n3529), .Z(n1067) );
  NOR U1222 ( .A(n3546), .B(n3628), .Z(n1066) );
  XOR U1223 ( .A(n1067), .B(n1066), .Z(n1164) );
  XOR U1224 ( .A(n1165), .B(n1164), .Z(n1214) );
  XOR U1225 ( .A(n1212), .B(n1214), .Z(n1206) );
  NOR U1226 ( .A(n3740), .B(n3688), .Z(n1365) );
  NOR U1227 ( .A(n3781), .B(n3748), .Z(n1085) );
  XOR U1228 ( .A(n1365), .B(n1085), .Z(n1221) );
  NOR U1229 ( .A(n3682), .B(n3622), .Z(n1068) );
  IV U1230 ( .A(n1068), .Z(n1151) );
  XOR U1231 ( .A(n1070), .B(n1069), .Z(n1150) );
  XOR U1232 ( .A(n1151), .B(n1150), .Z(n1222) );
  XOR U1233 ( .A(n1221), .B(n1222), .Z(n1204) );
  XOR U1234 ( .A(n1071), .B(n1204), .Z(n1205) );
  XOR U1235 ( .A(n1206), .B(n1205), .Z(n1188) );
  XOR U1236 ( .A(n1190), .B(n1188), .Z(n1192) );
  NOR U1237 ( .A(n3548), .B(n3763), .Z(n2434) );
  IV U1238 ( .A(n2434), .Z(n1073) );
  NOR U1239 ( .A(n1073), .B(n1072), .Z(n1078) );
  IV U1240 ( .A(n1074), .Z(n1075) );
  NOR U1241 ( .A(n1076), .B(n1075), .Z(n1077) );
  NOR U1242 ( .A(n1078), .B(n1077), .Z(n1130) );
  NOR U1243 ( .A(n2764), .B(n3749), .Z(n1079) );
  IV U1244 ( .A(n1079), .Z(n2420) );
  NOR U1245 ( .A(n2420), .B(n1476), .Z(n1084) );
  IV U1246 ( .A(n1080), .Z(n1082) );
  NOR U1247 ( .A(n1082), .B(n1081), .Z(n1083) );
  NOR U1248 ( .A(n1084), .B(n1083), .Z(n1127) );
  IV U1249 ( .A(n1085), .Z(n1087) );
  NOR U1250 ( .A(n1087), .B(n1086), .Z(n1092) );
  IV U1251 ( .A(n1088), .Z(n1090) );
  NOR U1252 ( .A(n1090), .B(n1089), .Z(n1091) );
  NOR U1253 ( .A(n1092), .B(n1091), .Z(n1126) );
  XOR U1254 ( .A(n1127), .B(n1126), .Z(n1128) );
  XOR U1255 ( .A(n1130), .B(n1128), .Z(n1191) );
  XOR U1256 ( .A(n1192), .B(n1191), .Z(n1241) );
  XOR U1257 ( .A(n1243), .B(n1241), .Z(n1244) );
  XOR U1258 ( .A(n1093), .B(n1244), .Z(n1121) );
  XOR U1259 ( .A(n1119), .B(n1121), .Z(n1122) );
  XOR U1260 ( .A(n1094), .B(n1122), .Z(n1113) );
  XOR U1261 ( .A(n1111), .B(n1113), .Z(n1115) );
  XOR U1262 ( .A(n1114), .B(n1115), .Z(n1106) );
  XOR U1263 ( .A(n1104), .B(n1106), .Z(n1108) );
  IV U1264 ( .A(n1095), .Z(n1096) );
  NOR U1265 ( .A(n1097), .B(n1096), .Z(n1102) );
  IV U1266 ( .A(n1098), .Z(n1099) );
  NOR U1267 ( .A(n1100), .B(n1099), .Z(n1101) );
  NOR U1268 ( .A(n1102), .B(n1101), .Z(n1103) );
  IV U1269 ( .A(n1103), .Z(n1107) );
  XOR U1270 ( .A(n1108), .B(n1107), .Z(N50) );
  IV U1271 ( .A(n1104), .Z(n1105) );
  NOR U1272 ( .A(n1106), .B(n1105), .Z(n1110) );
  NOR U1273 ( .A(n1108), .B(n1107), .Z(n1109) );
  NOR U1274 ( .A(n1110), .B(n1109), .Z(n1396) );
  IV U1275 ( .A(n1111), .Z(n1112) );
  NOR U1276 ( .A(n1113), .B(n1112), .Z(n1118) );
  IV U1277 ( .A(n1114), .Z(n1116) );
  NOR U1278 ( .A(n1116), .B(n1115), .Z(n1117) );
  NOR U1279 ( .A(n1118), .B(n1117), .Z(n1393) );
  IV U1280 ( .A(n1119), .Z(n1120) );
  NOR U1281 ( .A(n1121), .B(n1120), .Z(n1125) );
  NOR U1282 ( .A(n1123), .B(n1122), .Z(n1124) );
  NOR U1283 ( .A(n1125), .B(n1124), .Z(n1251) );
  NOR U1284 ( .A(n1127), .B(n1126), .Z(n1132) );
  IV U1285 ( .A(n1128), .Z(n1129) );
  NOR U1286 ( .A(n1130), .B(n1129), .Z(n1131) );
  NOR U1287 ( .A(n1132), .B(n1131), .Z(n1263) );
  NOR U1288 ( .A(n3775), .B(n3779), .Z(n2766) );
  IV U1289 ( .A(n2766), .Z(n3009) );
  NOR U1290 ( .A(n3009), .B(n1352), .Z(n1137) );
  IV U1291 ( .A(n1133), .Z(n1135) );
  NOR U1292 ( .A(n1135), .B(n1134), .Z(n1136) );
  NOR U1293 ( .A(n1137), .B(n1136), .Z(n1323) );
  NOR U1294 ( .A(n3548), .B(n3633), .Z(n1139) );
  IV U1295 ( .A(x[18]), .Z(n3764) );
  NOR U1296 ( .A(n3637), .B(n3764), .Z(n1138) );
  XOR U1297 ( .A(n1139), .B(n1138), .Z(n1359) );
  NOR U1298 ( .A(n3775), .B(n3625), .Z(n1140) );
  IV U1299 ( .A(n1140), .Z(n1354) );
  NOR U1300 ( .A(n3687), .B(n3062), .Z(n1142) );
  IV U1301 ( .A(y[18]), .Z(n3549) );
  NOR U1302 ( .A(n3680), .B(n3549), .Z(n1141) );
  XOR U1303 ( .A(n1142), .B(n1141), .Z(n1353) );
  XOR U1304 ( .A(n1354), .B(n1353), .Z(n1361) );
  XOR U1305 ( .A(n1359), .B(n1361), .Z(n1320) );
  NOR U1306 ( .A(n3787), .B(n3465), .Z(n1209) );
  NOR U1307 ( .A(n3779), .B(n3462), .Z(n1143) );
  XOR U1308 ( .A(n1209), .B(n1143), .Z(n1300) );
  NOR U1309 ( .A(n3619), .B(n2764), .Z(n1145) );
  NOR U1310 ( .A(n3746), .B(n3546), .Z(n1144) );
  XOR U1311 ( .A(n1145), .B(n1144), .Z(n1146) );
  IV U1312 ( .A(n1146), .Z(n1307) );
  NOR U1313 ( .A(n3742), .B(n3647), .Z(n1306) );
  XOR U1314 ( .A(n1307), .B(n1306), .Z(n1301) );
  XOR U1315 ( .A(n1300), .B(n1301), .Z(n1319) );
  XOR U1316 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U1317 ( .A(n1323), .B(n1321), .Z(n1294) );
  NOR U1318 ( .A(n3548), .B(n3462), .Z(n1468) );
  IV U1319 ( .A(n1468), .Z(n1149) );
  IV U1320 ( .A(n1147), .Z(n1148) );
  NOR U1321 ( .A(n1149), .B(n1148), .Z(n1154) );
  IV U1322 ( .A(n1150), .Z(n1152) );
  NOR U1323 ( .A(n1152), .B(n1151), .Z(n1153) );
  NOR U1324 ( .A(n1154), .B(n1153), .Z(n1292) );
  IV U1325 ( .A(n1292), .Z(n1161) );
  NOR U1326 ( .A(n3062), .B(n3741), .Z(n2562) );
  IV U1327 ( .A(n2562), .Z(n2812) );
  NOR U1328 ( .A(n2812), .B(n1155), .Z(n1160) );
  IV U1329 ( .A(n1156), .Z(n1157) );
  NOR U1330 ( .A(n1158), .B(n1157), .Z(n1159) );
  NOR U1331 ( .A(n1160), .B(n1159), .Z(n1291) );
  XOR U1332 ( .A(n1161), .B(n1291), .Z(n1293) );
  XOR U1333 ( .A(n1294), .B(n1293), .Z(n1282) );
  IV U1334 ( .A(n1282), .Z(n1187) );
  NOR U1335 ( .A(n3529), .B(n3628), .Z(n1628) );
  IV U1336 ( .A(n1628), .Z(n1163) );
  NOR U1337 ( .A(n1163), .B(n1162), .Z(n1168) );
  IV U1338 ( .A(n1164), .Z(n1166) );
  NOR U1339 ( .A(n1166), .B(n1165), .Z(n1167) );
  NOR U1340 ( .A(n1168), .B(n1167), .Z(n1329) );
  NOR U1341 ( .A(n3688), .B(n3748), .Z(n1217) );
  XOR U1342 ( .A(n1217), .B(n1169), .Z(n1367) );
  NOR U1343 ( .A(n3650), .B(n3467), .Z(n1171) );
  NOR U1344 ( .A(n3781), .B(n3682), .Z(n1170) );
  XOR U1345 ( .A(n1171), .B(n1170), .Z(n1313) );
  NOR U1346 ( .A(n3628), .B(n3776), .Z(n1172) );
  IV U1347 ( .A(n1172), .Z(n1336) );
  NOR U1348 ( .A(n3765), .B(n3646), .Z(n1174) );
  NOR U1349 ( .A(n3741), .B(n3635), .Z(n1173) );
  XOR U1350 ( .A(n1174), .B(n1173), .Z(n1335) );
  XOR U1351 ( .A(n1336), .B(n1335), .Z(n1315) );
  XOR U1352 ( .A(n1313), .B(n1315), .Z(n1369) );
  XOR U1353 ( .A(n1367), .B(n1369), .Z(n1326) );
  IV U1354 ( .A(o[17]), .Z(n1176) );
  NOR U1355 ( .A(n1176), .B(n1175), .Z(n1375) );
  NOR U1356 ( .A(n3749), .B(n3622), .Z(n1372) );
  NOR U1357 ( .A(n3529), .B(n3773), .Z(n1177) );
  IV U1358 ( .A(n1177), .Z(n1389) );
  XOR U1359 ( .A(n1389), .B(o[18]), .Z(n1374) );
  XOR U1360 ( .A(n1372), .B(n1374), .Z(n1377) );
  XOR U1361 ( .A(n1375), .B(n1377), .Z(n1327) );
  XOR U1362 ( .A(n1326), .B(n1327), .Z(n1178) );
  IV U1363 ( .A(n1178), .Z(n1328) );
  XOR U1364 ( .A(n1329), .B(n1328), .Z(n1280) );
  IV U1365 ( .A(n1179), .Z(n1180) );
  NOR U1366 ( .A(n1181), .B(n1180), .Z(n1186) );
  IV U1367 ( .A(n1182), .Z(n1183) );
  NOR U1368 ( .A(n1184), .B(n1183), .Z(n1185) );
  NOR U1369 ( .A(n1186), .B(n1185), .Z(n1278) );
  XOR U1370 ( .A(n1280), .B(n1278), .Z(n1281) );
  XOR U1371 ( .A(n1187), .B(n1281), .Z(n1265) );
  XOR U1372 ( .A(n1263), .B(n1265), .Z(n1268) );
  IV U1373 ( .A(n1188), .Z(n1189) );
  NOR U1374 ( .A(n1190), .B(n1189), .Z(n1194) );
  NOR U1375 ( .A(n1192), .B(n1191), .Z(n1193) );
  NOR U1376 ( .A(n1194), .B(n1193), .Z(n1266) );
  XOR U1377 ( .A(n1268), .B(n1266), .Z(n1256) );
  IV U1378 ( .A(n1195), .Z(n1196) );
  NOR U1379 ( .A(n1197), .B(n1196), .Z(n1202) );
  IV U1380 ( .A(n1198), .Z(n1199) );
  NOR U1381 ( .A(n1200), .B(n1199), .Z(n1201) );
  NOR U1382 ( .A(n1202), .B(n1201), .Z(n1275) );
  NOR U1383 ( .A(n1204), .B(n1203), .Z(n1208) );
  NOR U1384 ( .A(n1206), .B(n1205), .Z(n1207) );
  NOR U1385 ( .A(n1208), .B(n1207), .Z(n1288) );
  IV U1386 ( .A(n1209), .Z(n1498) );
  IV U1387 ( .A(n1210), .Z(n1211) );
  NOR U1388 ( .A(n1498), .B(n1211), .Z(n1216) );
  IV U1389 ( .A(n1212), .Z(n1213) );
  NOR U1390 ( .A(n1214), .B(n1213), .Z(n1215) );
  NOR U1391 ( .A(n1216), .B(n1215), .Z(n1286) );
  IV U1392 ( .A(n1217), .Z(n1220) );
  IV U1393 ( .A(n1218), .Z(n1219) );
  NOR U1394 ( .A(n1220), .B(n1219), .Z(n1225) );
  IV U1395 ( .A(n1221), .Z(n1223) );
  NOR U1396 ( .A(n1223), .B(n1222), .Z(n1224) );
  NOR U1397 ( .A(n1225), .B(n1224), .Z(n1285) );
  XOR U1398 ( .A(n1286), .B(n1285), .Z(n1226) );
  IV U1399 ( .A(n1226), .Z(n1287) );
  XOR U1400 ( .A(n1288), .B(n1287), .Z(n1273) );
  NOR U1401 ( .A(n1228), .B(n1227), .Z(n1232) );
  NOR U1402 ( .A(n1230), .B(n1229), .Z(n1231) );
  NOR U1403 ( .A(n1232), .B(n1231), .Z(n1271) );
  XOR U1404 ( .A(n1273), .B(n1271), .Z(n1274) );
  XOR U1405 ( .A(n1275), .B(n1274), .Z(n1258) );
  XOR U1406 ( .A(n1256), .B(n1258), .Z(n1260) );
  IV U1407 ( .A(n1233), .Z(n1234) );
  NOR U1408 ( .A(n1235), .B(n1234), .Z(n1239) );
  NOR U1409 ( .A(n1237), .B(n1236), .Z(n1238) );
  NOR U1410 ( .A(n1239), .B(n1238), .Z(n1240) );
  IV U1411 ( .A(n1240), .Z(n1259) );
  XOR U1412 ( .A(n1260), .B(n1259), .Z(n1250) );
  IV U1413 ( .A(n1241), .Z(n1242) );
  NOR U1414 ( .A(n1243), .B(n1242), .Z(n1247) );
  NOR U1415 ( .A(n1245), .B(n1244), .Z(n1246) );
  NOR U1416 ( .A(n1247), .B(n1246), .Z(n1248) );
  XOR U1417 ( .A(n1250), .B(n1248), .Z(n1253) );
  XOR U1418 ( .A(n1251), .B(n1253), .Z(n1395) );
  XOR U1419 ( .A(n1393), .B(n1395), .Z(n1398) );
  XOR U1420 ( .A(n1396), .B(n1398), .Z(N51) );
  IV U1421 ( .A(n1248), .Z(n1249) );
  NOR U1422 ( .A(n1250), .B(n1249), .Z(n1255) );
  IV U1423 ( .A(n1251), .Z(n1252) );
  NOR U1424 ( .A(n1253), .B(n1252), .Z(n1254) );
  NOR U1425 ( .A(n1255), .B(n1254), .Z(n1402) );
  IV U1426 ( .A(n1256), .Z(n1257) );
  NOR U1427 ( .A(n1258), .B(n1257), .Z(n1262) );
  NOR U1428 ( .A(n1260), .B(n1259), .Z(n1261) );
  NOR U1429 ( .A(n1262), .B(n1261), .Z(n1413) );
  IV U1430 ( .A(n1413), .Z(n1392) );
  IV U1431 ( .A(n1263), .Z(n1264) );
  NOR U1432 ( .A(n1265), .B(n1264), .Z(n1270) );
  IV U1433 ( .A(n1266), .Z(n1267) );
  NOR U1434 ( .A(n1268), .B(n1267), .Z(n1269) );
  NOR U1435 ( .A(n1270), .B(n1269), .Z(n1409) );
  IV U1436 ( .A(n1271), .Z(n1272) );
  NOR U1437 ( .A(n1273), .B(n1272), .Z(n1277) );
  NOR U1438 ( .A(n1275), .B(n1274), .Z(n1276) );
  NOR U1439 ( .A(n1277), .B(n1276), .Z(n1419) );
  IV U1440 ( .A(n1278), .Z(n1279) );
  NOR U1441 ( .A(n1280), .B(n1279), .Z(n1284) );
  NOR U1442 ( .A(n1282), .B(n1281), .Z(n1283) );
  NOR U1443 ( .A(n1284), .B(n1283), .Z(n1416) );
  NOR U1444 ( .A(n1286), .B(n1285), .Z(n1290) );
  NOR U1445 ( .A(n1288), .B(n1287), .Z(n1289) );
  NOR U1446 ( .A(n1290), .B(n1289), .Z(n1428) );
  NOR U1447 ( .A(n1292), .B(n1291), .Z(n1296) );
  NOR U1448 ( .A(n1294), .B(n1293), .Z(n1295) );
  NOR U1449 ( .A(n1296), .B(n1295), .Z(n1425) );
  NOR U1450 ( .A(n3465), .B(n3462), .Z(n2024) );
  IV U1451 ( .A(n2024), .Z(n1299) );
  IV U1452 ( .A(n1297), .Z(n1298) );
  NOR U1453 ( .A(n1299), .B(n1298), .Z(n1304) );
  IV U1454 ( .A(n1300), .Z(n1302) );
  NOR U1455 ( .A(n1302), .B(n1301), .Z(n1303) );
  NOR U1456 ( .A(n1304), .B(n1303), .Z(n1539) );
  NOR U1457 ( .A(n2764), .B(n3546), .Z(n3154) );
  IV U1458 ( .A(n3154), .Z(n3470) );
  NOR U1459 ( .A(n3470), .B(n1305), .Z(n1309) );
  IV U1460 ( .A(n1306), .Z(n2214) );
  NOR U1461 ( .A(n2214), .B(n1307), .Z(n1308) );
  NOR U1462 ( .A(n1309), .B(n1308), .Z(n1537) );
  NOR U1463 ( .A(n3682), .B(n3467), .Z(n1645) );
  IV U1464 ( .A(n1645), .Z(n1312) );
  IV U1465 ( .A(n1310), .Z(n1311) );
  NOR U1466 ( .A(n1312), .B(n1311), .Z(n1317) );
  IV U1467 ( .A(n1313), .Z(n1314) );
  NOR U1468 ( .A(n1315), .B(n1314), .Z(n1316) );
  NOR U1469 ( .A(n1317), .B(n1316), .Z(n1536) );
  XOR U1470 ( .A(n1537), .B(n1536), .Z(n1318) );
  IV U1471 ( .A(n1318), .Z(n1538) );
  XOR U1472 ( .A(n1539), .B(n1538), .Z(n1544) );
  NOR U1473 ( .A(n1320), .B(n1319), .Z(n1325) );
  IV U1474 ( .A(n1321), .Z(n1322) );
  NOR U1475 ( .A(n1323), .B(n1322), .Z(n1324) );
  NOR U1476 ( .A(n1325), .B(n1324), .Z(n1542) );
  XOR U1477 ( .A(n1544), .B(n1542), .Z(n1546) );
  NOR U1478 ( .A(n1327), .B(n1326), .Z(n1331) );
  NOR U1479 ( .A(n1329), .B(n1328), .Z(n1330) );
  NOR U1480 ( .A(n1331), .B(n1330), .Z(n1332) );
  IV U1481 ( .A(n1332), .Z(n1545) );
  XOR U1482 ( .A(n1546), .B(n1545), .Z(n1553) );
  NOR U1483 ( .A(n3765), .B(n3741), .Z(n2207) );
  IV U1484 ( .A(n2207), .Z(n1334) );
  NOR U1485 ( .A(n1334), .B(n1333), .Z(n1339) );
  IV U1486 ( .A(n1335), .Z(n1337) );
  NOR U1487 ( .A(n1337), .B(n1336), .Z(n1338) );
  NOR U1488 ( .A(n1339), .B(n1338), .Z(n1448) );
  NOR U1489 ( .A(n3776), .B(n3746), .Z(n1694) );
  NOR U1490 ( .A(n3635), .B(n2764), .Z(n1340) );
  XOR U1491 ( .A(n1694), .B(n1340), .Z(n1491) );
  NOR U1492 ( .A(n3775), .B(n3619), .Z(n1341) );
  IV U1493 ( .A(n1341), .Z(n1514) );
  NOR U1494 ( .A(n3781), .B(n3749), .Z(n1343) );
  NOR U1495 ( .A(n3549), .B(n3625), .Z(n1342) );
  XOR U1496 ( .A(n1343), .B(n1342), .Z(n1512) );
  XOR U1497 ( .A(n1514), .B(n1512), .Z(n1493) );
  XOR U1498 ( .A(n1491), .B(n1493), .Z(n1446) );
  NOR U1499 ( .A(n3650), .B(n3741), .Z(n1345) );
  XOR U1500 ( .A(n1345), .B(n1344), .Z(n1484) );
  NOR U1501 ( .A(n3628), .B(n3465), .Z(n1347) );
  NOR U1502 ( .A(n3787), .B(n3742), .Z(n1346) );
  XOR U1503 ( .A(n1347), .B(n1346), .Z(n1348) );
  IV U1504 ( .A(n1348), .Z(n1499) );
  XOR U1505 ( .A(n1499), .B(n1349), .Z(n1486) );
  XOR U1506 ( .A(n1484), .B(n1486), .Z(n1445) );
  XOR U1507 ( .A(n1446), .B(n1445), .Z(n1350) );
  IV U1508 ( .A(n1350), .Z(n1447) );
  XOR U1509 ( .A(n1448), .B(n1447), .Z(n1531) );
  NOR U1510 ( .A(n3062), .B(n3549), .Z(n1351) );
  IV U1511 ( .A(n1351), .Z(n3483) );
  NOR U1512 ( .A(n3483), .B(n1352), .Z(n1357) );
  IV U1513 ( .A(n1353), .Z(n1355) );
  NOR U1514 ( .A(n1355), .B(n1354), .Z(n1356) );
  NOR U1515 ( .A(n1357), .B(n1356), .Z(n1529) );
  XOR U1516 ( .A(n1531), .B(n1529), .Z(n1533) );
  NOR U1517 ( .A(n3633), .B(n3764), .Z(n2239) );
  IV U1518 ( .A(n2239), .Z(n2309) );
  IV U1519 ( .A(n1358), .Z(n1687) );
  NOR U1520 ( .A(n2309), .B(n1687), .Z(n1363) );
  IV U1521 ( .A(n1359), .Z(n1360) );
  NOR U1522 ( .A(n1361), .B(n1360), .Z(n1362) );
  NOR U1523 ( .A(n1363), .B(n1362), .Z(n1364) );
  IV U1524 ( .A(n1364), .Z(n1532) );
  XOR U1525 ( .A(n1533), .B(n1532), .Z(n1550) );
  NOR U1526 ( .A(n3748), .B(n3763), .Z(n1387) );
  IV U1527 ( .A(n1387), .Z(n1462) );
  IV U1528 ( .A(n1365), .Z(n1366) );
  NOR U1529 ( .A(n1462), .B(n1366), .Z(n1371) );
  IV U1530 ( .A(n1367), .Z(n1368) );
  NOR U1531 ( .A(n1369), .B(n1368), .Z(n1370) );
  NOR U1532 ( .A(n1371), .B(n1370), .Z(n1435) );
  IV U1533 ( .A(n1372), .Z(n1373) );
  NOR U1534 ( .A(n1374), .B(n1373), .Z(n1379) );
  IV U1535 ( .A(n1375), .Z(n1376) );
  NOR U1536 ( .A(n1377), .B(n1376), .Z(n1378) );
  NOR U1537 ( .A(n1379), .B(n1378), .Z(n1432) );
  NOR U1538 ( .A(n3647), .B(n3529), .Z(n1381) );
  NOR U1539 ( .A(n3548), .B(n3687), .Z(n1380) );
  XOR U1540 ( .A(n1381), .B(n1380), .Z(n1454) );
  IV U1541 ( .A(x[19]), .Z(n3689) );
  NOR U1542 ( .A(n3689), .B(n3637), .Z(n1382) );
  IV U1543 ( .A(n1382), .Z(n1478) );
  NOR U1544 ( .A(n3462), .B(n3062), .Z(n1384) );
  IV U1545 ( .A(y[19]), .Z(n3161) );
  NOR U1546 ( .A(n3680), .B(n3161), .Z(n1383) );
  XOR U1547 ( .A(n1384), .B(n1383), .Z(n1477) );
  XOR U1548 ( .A(n1478), .B(n1477), .Z(n1455) );
  XOR U1549 ( .A(n1454), .B(n1455), .Z(n1441) );
  NOR U1550 ( .A(n3467), .B(n3740), .Z(n1385) );
  XOR U1551 ( .A(n1386), .B(n1385), .Z(n1461) );
  XOR U1552 ( .A(n1461), .B(n1387), .Z(n1438) );
  IV U1553 ( .A(o[18]), .Z(n1388) );
  NOR U1554 ( .A(n1389), .B(n1388), .Z(n1505) );
  NOR U1555 ( .A(n3773), .B(n3764), .Z(n1390) );
  IV U1556 ( .A(n1390), .Z(n1525) );
  XOR U1557 ( .A(n1525), .B(o[19]), .Z(n1504) );
  XOR U1558 ( .A(n1391), .B(n1504), .Z(n1507) );
  XOR U1559 ( .A(n1505), .B(n1507), .Z(n1439) );
  XOR U1560 ( .A(n1438), .B(n1439), .Z(n1440) );
  XOR U1561 ( .A(n1441), .B(n1440), .Z(n1431) );
  XOR U1562 ( .A(n1432), .B(n1431), .Z(n1433) );
  XOR U1563 ( .A(n1435), .B(n1433), .Z(n1549) );
  XOR U1564 ( .A(n1550), .B(n1549), .Z(n1551) );
  XOR U1565 ( .A(n1553), .B(n1551), .Z(n1424) );
  XOR U1566 ( .A(n1425), .B(n1424), .Z(n1426) );
  XOR U1567 ( .A(n1428), .B(n1426), .Z(n1418) );
  XOR U1568 ( .A(n1416), .B(n1418), .Z(n1420) );
  XOR U1569 ( .A(n1419), .B(n1420), .Z(n1411) );
  XOR U1570 ( .A(n1409), .B(n1411), .Z(n1412) );
  XOR U1571 ( .A(n1392), .B(n1412), .Z(n1404) );
  XOR U1572 ( .A(n1402), .B(n1404), .Z(n1406) );
  IV U1573 ( .A(n1393), .Z(n1394) );
  NOR U1574 ( .A(n1395), .B(n1394), .Z(n1400) );
  IV U1575 ( .A(n1396), .Z(n1397) );
  NOR U1576 ( .A(n1398), .B(n1397), .Z(n1399) );
  NOR U1577 ( .A(n1400), .B(n1399), .Z(n1401) );
  IV U1578 ( .A(n1401), .Z(n1405) );
  XOR U1579 ( .A(n1406), .B(n1405), .Z(N52) );
  IV U1580 ( .A(n1402), .Z(n1403) );
  NOR U1581 ( .A(n1404), .B(n1403), .Z(n1408) );
  NOR U1582 ( .A(n1406), .B(n1405), .Z(n1407) );
  NOR U1583 ( .A(n1408), .B(n1407), .Z(n1711) );
  IV U1584 ( .A(n1409), .Z(n1410) );
  NOR U1585 ( .A(n1411), .B(n1410), .Z(n1415) );
  NOR U1586 ( .A(n1413), .B(n1412), .Z(n1414) );
  NOR U1587 ( .A(n1415), .B(n1414), .Z(n1708) );
  IV U1588 ( .A(n1416), .Z(n1417) );
  NOR U1589 ( .A(n1418), .B(n1417), .Z(n1423) );
  IV U1590 ( .A(n1419), .Z(n1421) );
  NOR U1591 ( .A(n1421), .B(n1420), .Z(n1422) );
  NOR U1592 ( .A(n1423), .B(n1422), .Z(n1559) );
  NOR U1593 ( .A(n1425), .B(n1424), .Z(n1430) );
  IV U1594 ( .A(n1426), .Z(n1427) );
  NOR U1595 ( .A(n1428), .B(n1427), .Z(n1429) );
  NOR U1596 ( .A(n1430), .B(n1429), .Z(n1556) );
  NOR U1597 ( .A(n1432), .B(n1431), .Z(n1437) );
  IV U1598 ( .A(n1433), .Z(n1434) );
  NOR U1599 ( .A(n1435), .B(n1434), .Z(n1436) );
  NOR U1600 ( .A(n1437), .B(n1436), .Z(n1582) );
  NOR U1601 ( .A(n1439), .B(n1438), .Z(n1444) );
  IV U1602 ( .A(n1440), .Z(n1442) );
  NOR U1603 ( .A(n1442), .B(n1441), .Z(n1443) );
  NOR U1604 ( .A(n1444), .B(n1443), .Z(n1580) );
  IV U1605 ( .A(n1580), .Z(n1528) );
  NOR U1606 ( .A(n1446), .B(n1445), .Z(n1450) );
  NOR U1607 ( .A(n1448), .B(n1447), .Z(n1449) );
  NOR U1608 ( .A(n1450), .B(n1449), .Z(n1591) );
  NOR U1609 ( .A(n3529), .B(n3687), .Z(n2212) );
  IV U1610 ( .A(n2212), .Z(n1453) );
  IV U1611 ( .A(n1451), .Z(n1452) );
  NOR U1612 ( .A(n1453), .B(n1452), .Z(n1458) );
  IV U1613 ( .A(n1454), .Z(n1456) );
  NOR U1614 ( .A(n1456), .B(n1455), .Z(n1457) );
  NOR U1615 ( .A(n1458), .B(n1457), .Z(n1601) );
  NOR U1616 ( .A(n3779), .B(n3467), .Z(n2224) );
  IV U1617 ( .A(n2224), .Z(n1460) );
  NOR U1618 ( .A(n1460), .B(n1459), .Z(n1464) );
  NOR U1619 ( .A(n1462), .B(n1461), .Z(n1463) );
  NOR U1620 ( .A(n1464), .B(n1463), .Z(n1655) );
  IV U1621 ( .A(y[20]), .Z(n3489) );
  NOR U1622 ( .A(n3680), .B(n3489), .Z(n1466) );
  XOR U1623 ( .A(n1466), .B(n1465), .Z(n1635) );
  NOR U1624 ( .A(n3647), .B(n3764), .Z(n1467) );
  IV U1625 ( .A(n1467), .Z(n1689) );
  IV U1626 ( .A(x[20]), .Z(n3782) );
  NOR U1627 ( .A(n3782), .B(n3637), .Z(n1469) );
  XOR U1628 ( .A(n1469), .B(n1468), .Z(n1688) );
  XOR U1629 ( .A(n1689), .B(n1688), .Z(n1637) );
  XOR U1630 ( .A(n1635), .B(n1637), .Z(n1653) );
  NOR U1631 ( .A(n3763), .B(n3682), .Z(n1471) );
  NOR U1632 ( .A(n3625), .B(n3161), .Z(n1470) );
  XOR U1633 ( .A(n1471), .B(n1470), .Z(n1615) );
  NOR U1634 ( .A(n3749), .B(n3688), .Z(n1472) );
  NOR U1635 ( .A(n3529), .B(n3787), .Z(n2315) );
  XOR U1636 ( .A(n1472), .B(n2315), .Z(n1473) );
  IV U1637 ( .A(n1473), .Z(n1622) );
  NOR U1638 ( .A(n3742), .B(n3628), .Z(n1497) );
  XOR U1639 ( .A(n1622), .B(n1497), .Z(n1616) );
  XOR U1640 ( .A(n1615), .B(n1616), .Z(n1652) );
  XOR U1641 ( .A(n1653), .B(n1652), .Z(n1474) );
  IV U1642 ( .A(n1474), .Z(n1654) );
  XOR U1643 ( .A(n1655), .B(n1654), .Z(n1600) );
  NOR U1644 ( .A(n3062), .B(n3161), .Z(n1475) );
  IV U1645 ( .A(n1475), .Z(n3801) );
  NOR U1646 ( .A(n3801), .B(n1476), .Z(n1481) );
  IV U1647 ( .A(n1477), .Z(n1479) );
  NOR U1648 ( .A(n1479), .B(n1478), .Z(n1480) );
  NOR U1649 ( .A(n1481), .B(n1480), .Z(n1598) );
  XOR U1650 ( .A(n1600), .B(n1598), .Z(n1603) );
  XOR U1651 ( .A(n1601), .B(n1603), .Z(n1593) );
  XOR U1652 ( .A(n1591), .B(n1593), .Z(n1594) );
  NOR U1653 ( .A(n3682), .B(n3741), .Z(n1878) );
  IV U1654 ( .A(n1878), .Z(n1801) );
  IV U1655 ( .A(n1482), .Z(n1483) );
  NOR U1656 ( .A(n1801), .B(n1483), .Z(n1488) );
  IV U1657 ( .A(n1484), .Z(n1485) );
  NOR U1658 ( .A(n1486), .B(n1485), .Z(n1487) );
  NOR U1659 ( .A(n1488), .B(n1487), .Z(n1586) );
  IV U1660 ( .A(n1586), .Z(n1496) );
  NOR U1661 ( .A(n2764), .B(n3776), .Z(n3534) );
  IV U1662 ( .A(n3534), .Z(n3821) );
  IV U1663 ( .A(n1489), .Z(n1490) );
  NOR U1664 ( .A(n3821), .B(n1490), .Z(n1495) );
  IV U1665 ( .A(n1491), .Z(n1492) );
  NOR U1666 ( .A(n1493), .B(n1492), .Z(n1494) );
  NOR U1667 ( .A(n1495), .B(n1494), .Z(n1585) );
  XOR U1668 ( .A(n1496), .B(n1585), .Z(n1588) );
  IV U1669 ( .A(n1497), .Z(n2400) );
  NOR U1670 ( .A(n2400), .B(n1498), .Z(n1502) );
  NOR U1671 ( .A(n1500), .B(n1499), .Z(n1501) );
  NOR U1672 ( .A(n1502), .B(n1501), .Z(n1659) );
  NOR U1673 ( .A(n1504), .B(n1503), .Z(n1509) );
  IV U1674 ( .A(n1505), .Z(n1506) );
  NOR U1675 ( .A(n1507), .B(n1506), .Z(n1508) );
  NOR U1676 ( .A(n1509), .B(n1508), .Z(n1658) );
  XOR U1677 ( .A(n1659), .B(n1658), .Z(n1510) );
  IV U1678 ( .A(n1510), .Z(n1662) );
  NOR U1679 ( .A(n3749), .B(n3549), .Z(n2561) );
  IV U1680 ( .A(n2561), .Z(n3022) );
  NOR U1681 ( .A(n3022), .B(n1511), .Z(n1516) );
  IV U1682 ( .A(n1512), .Z(n1513) );
  NOR U1683 ( .A(n1514), .B(n1513), .Z(n1515) );
  NOR U1684 ( .A(n1516), .B(n1515), .Z(n1669) );
  NOR U1685 ( .A(n3622), .B(n3779), .Z(n1518) );
  NOR U1686 ( .A(n3635), .B(n3775), .Z(n1517) );
  XOR U1687 ( .A(n1518), .B(n1517), .Z(n1608) );
  NOR U1688 ( .A(n3549), .B(n3619), .Z(n1519) );
  IV U1689 ( .A(n1519), .Z(n1698) );
  NOR U1690 ( .A(n3746), .B(n3465), .Z(n1521) );
  NOR U1691 ( .A(n3633), .B(n3776), .Z(n1520) );
  XOR U1692 ( .A(n1521), .B(n1520), .Z(n1697) );
  XOR U1693 ( .A(n1698), .B(n1697), .Z(n1610) );
  XOR U1694 ( .A(n1608), .B(n1610), .Z(n1683) );
  NOR U1695 ( .A(n3741), .B(n3740), .Z(n1680) );
  NOR U1696 ( .A(n3650), .B(n2764), .Z(n1523) );
  NOR U1697 ( .A(n3546), .B(n3687), .Z(n1522) );
  XOR U1698 ( .A(n1523), .B(n1522), .Z(n1524) );
  IV U1699 ( .A(n1524), .Z(n1642) );
  NOR U1700 ( .A(n3467), .B(n3748), .Z(n1641) );
  XOR U1701 ( .A(n1642), .B(n1641), .Z(n1681) );
  XOR U1702 ( .A(n1680), .B(n1681), .Z(n1682) );
  XOR U1703 ( .A(n1683), .B(n1682), .Z(n1665) );
  IV U1704 ( .A(o[19]), .Z(n1526) );
  NOR U1705 ( .A(n1526), .B(n1525), .Z(n1675) );
  NOR U1706 ( .A(n3781), .B(n3765), .Z(n1672) );
  NOR U1707 ( .A(n3689), .B(n3773), .Z(n1527) );
  IV U1708 ( .A(n1527), .Z(n1648) );
  XOR U1709 ( .A(n1648), .B(o[20]), .Z(n1673) );
  XOR U1710 ( .A(n1672), .B(n1673), .Z(n1677) );
  XOR U1711 ( .A(n1675), .B(n1677), .Z(n1666) );
  XOR U1712 ( .A(n1665), .B(n1666), .Z(n1668) );
  XOR U1713 ( .A(n1669), .B(n1668), .Z(n1660) );
  XOR U1714 ( .A(n1662), .B(n1660), .Z(n1587) );
  XOR U1715 ( .A(n1588), .B(n1587), .Z(n1595) );
  XOR U1716 ( .A(n1594), .B(n1595), .Z(n1579) );
  XOR U1717 ( .A(n1528), .B(n1579), .Z(n1581) );
  XOR U1718 ( .A(n1582), .B(n1581), .Z(n1576) );
  IV U1719 ( .A(n1529), .Z(n1530) );
  NOR U1720 ( .A(n1531), .B(n1530), .Z(n1535) );
  NOR U1721 ( .A(n1533), .B(n1532), .Z(n1534) );
  NOR U1722 ( .A(n1535), .B(n1534), .Z(n1574) );
  NOR U1723 ( .A(n1537), .B(n1536), .Z(n1541) );
  NOR U1724 ( .A(n1539), .B(n1538), .Z(n1540) );
  NOR U1725 ( .A(n1541), .B(n1540), .Z(n1572) );
  XOR U1726 ( .A(n1574), .B(n1572), .Z(n1575) );
  XOR U1727 ( .A(n1576), .B(n1575), .Z(n1567) );
  IV U1728 ( .A(n1542), .Z(n1543) );
  NOR U1729 ( .A(n1544), .B(n1543), .Z(n1548) );
  NOR U1730 ( .A(n1546), .B(n1545), .Z(n1547) );
  NOR U1731 ( .A(n1548), .B(n1547), .Z(n1566) );
  NOR U1732 ( .A(n1550), .B(n1549), .Z(n1555) );
  IV U1733 ( .A(n1551), .Z(n1552) );
  NOR U1734 ( .A(n1553), .B(n1552), .Z(n1554) );
  NOR U1735 ( .A(n1555), .B(n1554), .Z(n1564) );
  XOR U1736 ( .A(n1566), .B(n1564), .Z(n1568) );
  XOR U1737 ( .A(n1567), .B(n1568), .Z(n1558) );
  XOR U1738 ( .A(n1556), .B(n1558), .Z(n1561) );
  XOR U1739 ( .A(n1559), .B(n1561), .Z(n1710) );
  XOR U1740 ( .A(n1708), .B(n1710), .Z(n1713) );
  XOR U1741 ( .A(n1711), .B(n1713), .Z(N53) );
  IV U1742 ( .A(n1556), .Z(n1557) );
  NOR U1743 ( .A(n1558), .B(n1557), .Z(n1563) );
  IV U1744 ( .A(n1559), .Z(n1560) );
  NOR U1745 ( .A(n1561), .B(n1560), .Z(n1562) );
  NOR U1746 ( .A(n1563), .B(n1562), .Z(n1717) );
  IV U1747 ( .A(n1564), .Z(n1565) );
  NOR U1748 ( .A(n1566), .B(n1565), .Z(n1571) );
  IV U1749 ( .A(n1567), .Z(n1569) );
  NOR U1750 ( .A(n1569), .B(n1568), .Z(n1570) );
  NOR U1751 ( .A(n1571), .B(n1570), .Z(n1727) );
  IV U1752 ( .A(n1572), .Z(n1573) );
  NOR U1753 ( .A(n1574), .B(n1573), .Z(n1578) );
  NOR U1754 ( .A(n1576), .B(n1575), .Z(n1577) );
  NOR U1755 ( .A(n1578), .B(n1577), .Z(n1724) );
  NOR U1756 ( .A(n1580), .B(n1579), .Z(n1584) );
  NOR U1757 ( .A(n1582), .B(n1581), .Z(n1583) );
  NOR U1758 ( .A(n1584), .B(n1583), .Z(n1736) );
  NOR U1759 ( .A(n1586), .B(n1585), .Z(n1590) );
  NOR U1760 ( .A(n1588), .B(n1587), .Z(n1589) );
  NOR U1761 ( .A(n1590), .B(n1589), .Z(n1733) );
  IV U1762 ( .A(n1591), .Z(n1592) );
  NOR U1763 ( .A(n1593), .B(n1592), .Z(n1597) );
  NOR U1764 ( .A(n1595), .B(n1594), .Z(n1596) );
  NOR U1765 ( .A(n1597), .B(n1596), .Z(n1741) );
  IV U1766 ( .A(n1598), .Z(n1599) );
  NOR U1767 ( .A(n1600), .B(n1599), .Z(n1605) );
  IV U1768 ( .A(n1601), .Z(n1602) );
  NOR U1769 ( .A(n1603), .B(n1602), .Z(n1604) );
  NOR U1770 ( .A(n1605), .B(n1604), .Z(n1750) );
  IV U1771 ( .A(n1606), .Z(n1607) );
  NOR U1772 ( .A(n3009), .B(n1607), .Z(n1612) );
  IV U1773 ( .A(n1608), .Z(n1609) );
  NOR U1774 ( .A(n1610), .B(n1609), .Z(n1611) );
  NOR U1775 ( .A(n1612), .B(n1611), .Z(n1761) );
  NOR U1776 ( .A(n3682), .B(n3161), .Z(n2783) );
  IV U1777 ( .A(n2783), .Z(n2785) );
  IV U1778 ( .A(n1613), .Z(n1614) );
  NOR U1779 ( .A(n2785), .B(n1614), .Z(n1619) );
  IV U1780 ( .A(n1615), .Z(n1617) );
  NOR U1781 ( .A(n1617), .B(n1616), .Z(n1618) );
  NOR U1782 ( .A(n1619), .B(n1618), .Z(n1760) );
  XOR U1783 ( .A(n1761), .B(n1760), .Z(n1620) );
  IV U1784 ( .A(n1620), .Z(n1762) );
  NOR U1785 ( .A(n3688), .B(n3529), .Z(n3160) );
  IV U1786 ( .A(n3160), .Z(n3523) );
  NOR U1787 ( .A(n3523), .B(n1621), .Z(n1624) );
  NOR U1788 ( .A(n2400), .B(n1622), .Z(n1623) );
  NOR U1789 ( .A(n1624), .B(n1623), .Z(n1797) );
  NOR U1790 ( .A(n3489), .B(n3625), .Z(n1817) );
  IV U1791 ( .A(y[21]), .Z(n3780) );
  NOR U1792 ( .A(n3680), .B(n3780), .Z(n1625) );
  IV U1793 ( .A(n1625), .Z(n1816) );
  NOR U1794 ( .A(n3062), .B(n3622), .Z(n1814) );
  XOR U1795 ( .A(n1816), .B(n1814), .Z(n1819) );
  XOR U1796 ( .A(n1817), .B(n1819), .Z(n1811) );
  IV U1797 ( .A(x[21]), .Z(n3621) );
  NOR U1798 ( .A(n3621), .B(n3637), .Z(n1627) );
  XOR U1799 ( .A(n1627), .B(n1626), .Z(n1809) );
  XOR U1800 ( .A(n1811), .B(n1809), .Z(n1795) );
  NOR U1801 ( .A(n3765), .B(n3688), .Z(n1629) );
  XOR U1802 ( .A(n1629), .B(n1628), .Z(n1824) );
  NOR U1803 ( .A(n3787), .B(n3764), .Z(n1839) );
  NOR U1804 ( .A(n3775), .B(n3650), .Z(n1630) );
  IV U1805 ( .A(n1630), .Z(n1838) );
  NOR U1806 ( .A(n3742), .B(n3746), .Z(n1836) );
  XOR U1807 ( .A(n1838), .B(n1836), .Z(n1840) );
  XOR U1808 ( .A(n1839), .B(n1840), .Z(n1825) );
  XOR U1809 ( .A(n1824), .B(n1825), .Z(n1794) );
  XOR U1810 ( .A(n1795), .B(n1794), .Z(n1631) );
  IV U1811 ( .A(n1631), .Z(n1796) );
  XOR U1812 ( .A(n1797), .B(n1796), .Z(n1789) );
  NOR U1813 ( .A(n3489), .B(n3062), .Z(n1632) );
  IV U1814 ( .A(n1632), .Z(n3789) );
  IV U1815 ( .A(n1633), .Z(n1634) );
  NOR U1816 ( .A(n3789), .B(n1634), .Z(n1639) );
  IV U1817 ( .A(n1635), .Z(n1636) );
  NOR U1818 ( .A(n1637), .B(n1636), .Z(n1638) );
  NOR U1819 ( .A(n1639), .B(n1638), .Z(n1787) );
  XOR U1820 ( .A(n1789), .B(n1787), .Z(n1790) );
  NOR U1821 ( .A(n3470), .B(n1640), .Z(n1644) );
  IV U1822 ( .A(n1641), .Z(n1800) );
  NOR U1823 ( .A(n1800), .B(n1642), .Z(n1643) );
  NOR U1824 ( .A(n1644), .B(n1643), .Z(n1783) );
  NOR U1825 ( .A(n3741), .B(n3748), .Z(n2004) );
  XOR U1826 ( .A(n1645), .B(n2004), .Z(n1802) );
  NOR U1827 ( .A(n3749), .B(n3763), .Z(n1646) );
  IV U1828 ( .A(n1646), .Z(n1864) );
  NOR U1829 ( .A(n3465), .B(n3633), .Z(n1693) );
  NOR U1830 ( .A(n2764), .B(n3740), .Z(n1647) );
  XOR U1831 ( .A(n1693), .B(n1647), .Z(n1863) );
  XOR U1832 ( .A(n1864), .B(n1863), .Z(n1804) );
  XOR U1833 ( .A(n1802), .B(n1804), .Z(n1781) );
  IV U1834 ( .A(o[20]), .Z(n1649) );
  NOR U1835 ( .A(n1649), .B(n1648), .Z(n1856) );
  NOR U1836 ( .A(n3781), .B(n3779), .Z(n1854) );
  NOR U1837 ( .A(n3773), .B(n3782), .Z(n1650) );
  IV U1838 ( .A(n1650), .Z(n1871) );
  XOR U1839 ( .A(n1871), .B(o[21]), .Z(n1855) );
  XOR U1840 ( .A(n1854), .B(n1855), .Z(n1858) );
  XOR U1841 ( .A(n1856), .B(n1858), .Z(n1780) );
  XOR U1842 ( .A(n1781), .B(n1780), .Z(n1651) );
  IV U1843 ( .A(n1651), .Z(n1782) );
  XOR U1844 ( .A(n1783), .B(n1782), .Z(n1791) );
  XOR U1845 ( .A(n1790), .B(n1791), .Z(n1763) );
  XOR U1846 ( .A(n1762), .B(n1763), .Z(n1748) );
  NOR U1847 ( .A(n1653), .B(n1652), .Z(n1657) );
  NOR U1848 ( .A(n1655), .B(n1654), .Z(n1656) );
  NOR U1849 ( .A(n1657), .B(n1656), .Z(n1746) );
  XOR U1850 ( .A(n1748), .B(n1746), .Z(n1749) );
  XOR U1851 ( .A(n1750), .B(n1749), .Z(n1740) );
  NOR U1852 ( .A(n1659), .B(n1658), .Z(n1664) );
  IV U1853 ( .A(n1660), .Z(n1661) );
  NOR U1854 ( .A(n1662), .B(n1661), .Z(n1663) );
  NOR U1855 ( .A(n1664), .B(n1663), .Z(n1757) );
  IV U1856 ( .A(n1665), .Z(n1667) );
  NOR U1857 ( .A(n1667), .B(n1666), .Z(n1671) );
  NOR U1858 ( .A(n1669), .B(n1668), .Z(n1670) );
  NOR U1859 ( .A(n1671), .B(n1670), .Z(n1754) );
  IV U1860 ( .A(n1672), .Z(n1674) );
  NOR U1861 ( .A(n1674), .B(n1673), .Z(n1679) );
  IV U1862 ( .A(n1675), .Z(n1676) );
  NOR U1863 ( .A(n1677), .B(n1676), .Z(n1678) );
  NOR U1864 ( .A(n1679), .B(n1678), .Z(n1767) );
  IV U1865 ( .A(n1680), .Z(n2423) );
  NOR U1866 ( .A(n2423), .B(n1681), .Z(n1685) );
  NOR U1867 ( .A(n1683), .B(n1682), .Z(n1684) );
  NOR U1868 ( .A(n1685), .B(n1684), .Z(n1766) );
  XOR U1869 ( .A(n1767), .B(n1766), .Z(n1768) );
  NOR U1870 ( .A(n3462), .B(n3782), .Z(n1686) );
  IV U1871 ( .A(n1686), .Z(n3193) );
  NOR U1872 ( .A(n3193), .B(n1687), .Z(n1692) );
  IV U1873 ( .A(n1688), .Z(n1690) );
  NOR U1874 ( .A(n1690), .B(n1689), .Z(n1691) );
  NOR U1875 ( .A(n1692), .B(n1691), .Z(n1777) );
  IV U1876 ( .A(n1693), .Z(n1696) );
  IV U1877 ( .A(n1694), .Z(n1695) );
  NOR U1878 ( .A(n1696), .B(n1695), .Z(n1701) );
  IV U1879 ( .A(n1697), .Z(n1699) );
  NOR U1880 ( .A(n1699), .B(n1698), .Z(n1700) );
  NOR U1881 ( .A(n1701), .B(n1700), .Z(n1774) );
  NOR U1882 ( .A(n3635), .B(n3549), .Z(n1703) );
  NOR U1883 ( .A(n3546), .B(n3462), .Z(n1702) );
  XOR U1884 ( .A(n1703), .B(n1702), .Z(n1849) );
  NOR U1885 ( .A(n3689), .B(n3647), .Z(n1704) );
  IV U1886 ( .A(n1704), .Z(n1832) );
  NOR U1887 ( .A(n3548), .B(n3646), .Z(n1706) );
  NOR U1888 ( .A(n3161), .B(n3619), .Z(n1705) );
  XOR U1889 ( .A(n1706), .B(n1705), .Z(n1831) );
  XOR U1890 ( .A(n1832), .B(n1831), .Z(n1851) );
  XOR U1891 ( .A(n1849), .B(n1851), .Z(n1773) );
  XOR U1892 ( .A(n1774), .B(n1773), .Z(n1775) );
  XOR U1893 ( .A(n1777), .B(n1775), .Z(n1769) );
  XOR U1894 ( .A(n1768), .B(n1769), .Z(n1753) );
  XOR U1895 ( .A(n1754), .B(n1753), .Z(n1755) );
  XOR U1896 ( .A(n1757), .B(n1755), .Z(n1739) );
  XOR U1897 ( .A(n1740), .B(n1739), .Z(n1707) );
  IV U1898 ( .A(n1707), .Z(n1742) );
  XOR U1899 ( .A(n1741), .B(n1742), .Z(n1732) );
  XOR U1900 ( .A(n1733), .B(n1732), .Z(n1734) );
  XOR U1901 ( .A(n1736), .B(n1734), .Z(n1726) );
  XOR U1902 ( .A(n1724), .B(n1726), .Z(n1728) );
  XOR U1903 ( .A(n1727), .B(n1728), .Z(n1719) );
  XOR U1904 ( .A(n1717), .B(n1719), .Z(n1721) );
  IV U1905 ( .A(n1708), .Z(n1709) );
  NOR U1906 ( .A(n1710), .B(n1709), .Z(n1715) );
  IV U1907 ( .A(n1711), .Z(n1712) );
  NOR U1908 ( .A(n1713), .B(n1712), .Z(n1714) );
  NOR U1909 ( .A(n1715), .B(n1714), .Z(n1716) );
  IV U1910 ( .A(n1716), .Z(n1720) );
  XOR U1911 ( .A(n1721), .B(n1720), .Z(N54) );
  IV U1912 ( .A(n1717), .Z(n1718) );
  NOR U1913 ( .A(n1719), .B(n1718), .Z(n1723) );
  NOR U1914 ( .A(n1721), .B(n1720), .Z(n1722) );
  NOR U1915 ( .A(n1723), .B(n1722), .Z(n1885) );
  IV U1916 ( .A(n1724), .Z(n1725) );
  NOR U1917 ( .A(n1726), .B(n1725), .Z(n1731) );
  IV U1918 ( .A(n1727), .Z(n1729) );
  NOR U1919 ( .A(n1729), .B(n1728), .Z(n1730) );
  NOR U1920 ( .A(n1731), .B(n1730), .Z(n1882) );
  NOR U1921 ( .A(n1733), .B(n1732), .Z(n1738) );
  IV U1922 ( .A(n1734), .Z(n1735) );
  NOR U1923 ( .A(n1736), .B(n1735), .Z(n1737) );
  NOR U1924 ( .A(n1738), .B(n1737), .Z(n1893) );
  NOR U1925 ( .A(n1740), .B(n1739), .Z(n1745) );
  IV U1926 ( .A(n1741), .Z(n1743) );
  NOR U1927 ( .A(n1743), .B(n1742), .Z(n1744) );
  NOR U1928 ( .A(n1745), .B(n1744), .Z(n1890) );
  IV U1929 ( .A(n1746), .Z(n1747) );
  NOR U1930 ( .A(n1748), .B(n1747), .Z(n1752) );
  NOR U1931 ( .A(n1750), .B(n1749), .Z(n1751) );
  NOR U1932 ( .A(n1752), .B(n1751), .Z(n1902) );
  IV U1933 ( .A(n1902), .Z(n1881) );
  NOR U1934 ( .A(n1754), .B(n1753), .Z(n1759) );
  IV U1935 ( .A(n1755), .Z(n1756) );
  NOR U1936 ( .A(n1757), .B(n1756), .Z(n1758) );
  NOR U1937 ( .A(n1759), .B(n1758), .Z(n1898) );
  NOR U1938 ( .A(n1761), .B(n1760), .Z(n1765) );
  NOR U1939 ( .A(n1763), .B(n1762), .Z(n1764) );
  NOR U1940 ( .A(n1765), .B(n1764), .Z(n1909) );
  NOR U1941 ( .A(n1767), .B(n1766), .Z(n1772) );
  IV U1942 ( .A(n1768), .Z(n1770) );
  NOR U1943 ( .A(n1770), .B(n1769), .Z(n1771) );
  NOR U1944 ( .A(n1772), .B(n1771), .Z(n1906) );
  NOR U1945 ( .A(n1774), .B(n1773), .Z(n1779) );
  IV U1946 ( .A(n1775), .Z(n1776) );
  NOR U1947 ( .A(n1777), .B(n1776), .Z(n1778) );
  NOR U1948 ( .A(n1779), .B(n1778), .Z(n1914) );
  NOR U1949 ( .A(n1781), .B(n1780), .Z(n1785) );
  NOR U1950 ( .A(n1783), .B(n1782), .Z(n1784) );
  NOR U1951 ( .A(n1785), .B(n1784), .Z(n1786) );
  IV U1952 ( .A(n1786), .Z(n1915) );
  XOR U1953 ( .A(n1914), .B(n1915), .Z(n1919) );
  IV U1954 ( .A(n1787), .Z(n1788) );
  NOR U1955 ( .A(n1789), .B(n1788), .Z(n1793) );
  NOR U1956 ( .A(n1791), .B(n1790), .Z(n1792) );
  NOR U1957 ( .A(n1793), .B(n1792), .Z(n1927) );
  NOR U1958 ( .A(n1795), .B(n1794), .Z(n1799) );
  NOR U1959 ( .A(n1797), .B(n1796), .Z(n1798) );
  NOR U1960 ( .A(n1799), .B(n1798), .Z(n1923) );
  NOR U1961 ( .A(n1801), .B(n1800), .Z(n1806) );
  IV U1962 ( .A(n1802), .Z(n1803) );
  NOR U1963 ( .A(n1804), .B(n1803), .Z(n1805) );
  NOR U1964 ( .A(n1806), .B(n1805), .Z(n1938) );
  NOR U1965 ( .A(n3621), .B(n3687), .Z(n2961) );
  IV U1966 ( .A(n2961), .Z(n3181) );
  IV U1967 ( .A(n1807), .Z(n1808) );
  NOR U1968 ( .A(n3181), .B(n1808), .Z(n1813) );
  IV U1969 ( .A(n1809), .Z(n1810) );
  NOR U1970 ( .A(n1811), .B(n1810), .Z(n1812) );
  NOR U1971 ( .A(n1813), .B(n1812), .Z(n1937) );
  XOR U1972 ( .A(n1938), .B(n1937), .Z(n1939) );
  IV U1973 ( .A(n1814), .Z(n1815) );
  NOR U1974 ( .A(n1816), .B(n1815), .Z(n1821) );
  IV U1975 ( .A(n1817), .Z(n1818) );
  NOR U1976 ( .A(n1819), .B(n1818), .Z(n1820) );
  NOR U1977 ( .A(n1821), .B(n1820), .Z(n1966) );
  IV U1978 ( .A(n1822), .Z(n1823) );
  NOR U1979 ( .A(n3523), .B(n1823), .Z(n1828) );
  IV U1980 ( .A(n1824), .Z(n1826) );
  NOR U1981 ( .A(n1826), .B(n1825), .Z(n1827) );
  NOR U1982 ( .A(n1828), .B(n1827), .Z(n1965) );
  XOR U1983 ( .A(n1966), .B(n1965), .Z(n1967) );
  NOR U1984 ( .A(n3161), .B(n3548), .Z(n3794) );
  IV U1985 ( .A(n3794), .Z(n1830) );
  NOR U1986 ( .A(n1830), .B(n1829), .Z(n1835) );
  IV U1987 ( .A(n1831), .Z(n1833) );
  NOR U1988 ( .A(n1833), .B(n1832), .Z(n1834) );
  NOR U1989 ( .A(n1835), .B(n1834), .Z(n1954) );
  IV U1990 ( .A(n1954), .Z(n1846) );
  IV U1991 ( .A(n1836), .Z(n1837) );
  NOR U1992 ( .A(n1838), .B(n1837), .Z(n1842) );
  IV U1993 ( .A(n1839), .Z(n2229) );
  NOR U1994 ( .A(n2229), .B(n1840), .Z(n1841) );
  NOR U1995 ( .A(n1842), .B(n1841), .Z(n1952) );
  NOR U1996 ( .A(n3625), .B(n3780), .Z(n2033) );
  NOR U1997 ( .A(n3548), .B(n3622), .Z(n1843) );
  IV U1998 ( .A(n1843), .Z(n2034) );
  XOR U1999 ( .A(n2033), .B(n2034), .Z(n2037) );
  IV U2000 ( .A(x[22]), .Z(n3645) );
  NOR U2001 ( .A(n3645), .B(n3637), .Z(n1991) );
  IV U2002 ( .A(y[22]), .Z(n3766) );
  NOR U2003 ( .A(n3680), .B(n3766), .Z(n1844) );
  IV U2004 ( .A(n1844), .Z(n1990) );
  XOR U2005 ( .A(n1990), .B(n1845), .Z(n1993) );
  XOR U2006 ( .A(n1991), .B(n1993), .Z(n2036) );
  XOR U2007 ( .A(n2037), .B(n2036), .Z(n1950) );
  XOR U2008 ( .A(n1952), .B(n1950), .Z(n1953) );
  XOR U2009 ( .A(n1846), .B(n1953), .Z(n1968) );
  XOR U2010 ( .A(n1967), .B(n1968), .Z(n1940) );
  XOR U2011 ( .A(n1939), .B(n1940), .Z(n1946) );
  NOR U2012 ( .A(n3549), .B(n3546), .Z(n1847) );
  IV U2013 ( .A(n1847), .Z(n3790) );
  NOR U2014 ( .A(n3790), .B(n1848), .Z(n1853) );
  IV U2015 ( .A(n1849), .Z(n1850) );
  NOR U2016 ( .A(n1851), .B(n1850), .Z(n1852) );
  NOR U2017 ( .A(n1853), .B(n1852), .Z(n1945) );
  IV U2018 ( .A(n1854), .Z(n2418) );
  NOR U2019 ( .A(n2418), .B(n1855), .Z(n1860) );
  IV U2020 ( .A(n1856), .Z(n1857) );
  NOR U2021 ( .A(n1858), .B(n1857), .Z(n1859) );
  NOR U2022 ( .A(n1860), .B(n1859), .Z(n1934) );
  NOR U2023 ( .A(n3465), .B(n2764), .Z(n3654) );
  IV U2024 ( .A(n3654), .Z(n1862) );
  NOR U2025 ( .A(n1862), .B(n1861), .Z(n1867) );
  IV U2026 ( .A(n1863), .Z(n1865) );
  NOR U2027 ( .A(n1865), .B(n1864), .Z(n1866) );
  NOR U2028 ( .A(n1867), .B(n1866), .Z(n1961) );
  NOR U2029 ( .A(n3619), .B(n3489), .Z(n1868) );
  NOR U2030 ( .A(n3763), .B(n3765), .Z(n2549) );
  XOR U2031 ( .A(n1868), .B(n2549), .Z(n2059) );
  NOR U2032 ( .A(n3689), .B(n3787), .Z(n1869) );
  IV U2033 ( .A(n1869), .Z(n2044) );
  NOR U2034 ( .A(n3546), .B(n3646), .Z(n1870) );
  NOR U2035 ( .A(n3647), .B(n3782), .Z(n2775) );
  XOR U2036 ( .A(n1870), .B(n2775), .Z(n2043) );
  XOR U2037 ( .A(n2044), .B(n2043), .Z(n2061) );
  XOR U2038 ( .A(n2059), .B(n2061), .Z(n1958) );
  IV U2039 ( .A(o[21]), .Z(n1872) );
  NOR U2040 ( .A(n1872), .B(n1871), .Z(n1984) );
  NOR U2041 ( .A(n3688), .B(n3779), .Z(n1981) );
  NOR U2042 ( .A(n3773), .B(n3621), .Z(n1873) );
  IV U2043 ( .A(n1873), .Z(n2052) );
  XOR U2044 ( .A(n2052), .B(o[22]), .Z(n1983) );
  XOR U2045 ( .A(n1981), .B(n1983), .Z(n1986) );
  XOR U2046 ( .A(n1984), .B(n1986), .Z(n1957) );
  XOR U2047 ( .A(n1958), .B(n1957), .Z(n1959) );
  XOR U2048 ( .A(n1961), .B(n1959), .Z(n1931) );
  NOR U2049 ( .A(n3465), .B(n3687), .Z(n2064) );
  NOR U2050 ( .A(n3161), .B(n3635), .Z(n1874) );
  IV U2051 ( .A(n1874), .Z(n2065) );
  XOR U2052 ( .A(n2064), .B(n2065), .Z(n2067) );
  NOR U2053 ( .A(n3529), .B(n3746), .Z(n1875) );
  IV U2054 ( .A(n1875), .Z(n1997) );
  NOR U2055 ( .A(n3742), .B(n3633), .Z(n1877) );
  NOR U2056 ( .A(n3628), .B(n3764), .Z(n1876) );
  XOR U2057 ( .A(n1877), .B(n1876), .Z(n1996) );
  XOR U2058 ( .A(n1997), .B(n1996), .Z(n2068) );
  XOR U2059 ( .A(n2067), .B(n2068), .Z(n1976) );
  NOR U2060 ( .A(n3775), .B(n3740), .Z(n1973) );
  NOR U2061 ( .A(n3748), .B(n2764), .Z(n2141) );
  XOR U2062 ( .A(n2141), .B(n1878), .Z(n2007) );
  NOR U2063 ( .A(n3749), .B(n3467), .Z(n2015) );
  NOR U2064 ( .A(n3776), .B(n3462), .Z(n1879) );
  IV U2065 ( .A(n1879), .Z(n2014) );
  NOR U2066 ( .A(n3549), .B(n3650), .Z(n2012) );
  XOR U2067 ( .A(n2014), .B(n2012), .Z(n2017) );
  XOR U2068 ( .A(n2015), .B(n2017), .Z(n2009) );
  XOR U2069 ( .A(n2007), .B(n2009), .Z(n1975) );
  XOR U2070 ( .A(n1973), .B(n1975), .Z(n1977) );
  XOR U2071 ( .A(n1976), .B(n1977), .Z(n1930) );
  XOR U2072 ( .A(n1931), .B(n1930), .Z(n1932) );
  XOR U2073 ( .A(n1934), .B(n1932), .Z(n1944) );
  XOR U2074 ( .A(n1945), .B(n1944), .Z(n1880) );
  IV U2075 ( .A(n1880), .Z(n1947) );
  XOR U2076 ( .A(n1946), .B(n1947), .Z(n1925) );
  XOR U2077 ( .A(n1923), .B(n1925), .Z(n1926) );
  XOR U2078 ( .A(n1927), .B(n1926), .Z(n1917) );
  XOR U2079 ( .A(n1919), .B(n1917), .Z(n1908) );
  XOR U2080 ( .A(n1906), .B(n1908), .Z(n1911) );
  XOR U2081 ( .A(n1909), .B(n1911), .Z(n1900) );
  XOR U2082 ( .A(n1898), .B(n1900), .Z(n1901) );
  XOR U2083 ( .A(n1881), .B(n1901), .Z(n1892) );
  XOR U2084 ( .A(n1890), .B(n1892), .Z(n1895) );
  XOR U2085 ( .A(n1893), .B(n1895), .Z(n1884) );
  XOR U2086 ( .A(n1882), .B(n1884), .Z(n1887) );
  XOR U2087 ( .A(n1885), .B(n1887), .Z(N55) );
  IV U2088 ( .A(n1882), .Z(n1883) );
  NOR U2089 ( .A(n1884), .B(n1883), .Z(n1889) );
  IV U2090 ( .A(n1885), .Z(n1886) );
  NOR U2091 ( .A(n1887), .B(n1886), .Z(n1888) );
  NOR U2092 ( .A(n1889), .B(n1888), .Z(n2076) );
  IV U2093 ( .A(n1890), .Z(n1891) );
  NOR U2094 ( .A(n1892), .B(n1891), .Z(n1897) );
  IV U2095 ( .A(n1893), .Z(n1894) );
  NOR U2096 ( .A(n1895), .B(n1894), .Z(n1896) );
  NOR U2097 ( .A(n1897), .B(n1896), .Z(n2073) );
  IV U2098 ( .A(n1898), .Z(n1899) );
  NOR U2099 ( .A(n1900), .B(n1899), .Z(n1904) );
  NOR U2100 ( .A(n1902), .B(n1901), .Z(n1903) );
  NOR U2101 ( .A(n1904), .B(n1903), .Z(n1905) );
  IV U2102 ( .A(n1905), .Z(n2083) );
  IV U2103 ( .A(n1906), .Z(n1907) );
  NOR U2104 ( .A(n1908), .B(n1907), .Z(n1913) );
  IV U2105 ( .A(n1909), .Z(n1910) );
  NOR U2106 ( .A(n1911), .B(n1910), .Z(n1912) );
  NOR U2107 ( .A(n1913), .B(n1912), .Z(n2079) );
  IV U2108 ( .A(n1914), .Z(n1916) );
  NOR U2109 ( .A(n1916), .B(n1915), .Z(n1921) );
  IV U2110 ( .A(n1917), .Z(n1918) );
  NOR U2111 ( .A(n1919), .B(n1918), .Z(n1920) );
  NOR U2112 ( .A(n1921), .B(n1920), .Z(n1922) );
  IV U2113 ( .A(n1922), .Z(n2088) );
  IV U2114 ( .A(n1923), .Z(n1924) );
  NOR U2115 ( .A(n1925), .B(n1924), .Z(n1929) );
  NOR U2116 ( .A(n1927), .B(n1926), .Z(n1928) );
  NOR U2117 ( .A(n1929), .B(n1928), .Z(n2086) );
  XOR U2118 ( .A(n2088), .B(n2086), .Z(n2089) );
  IV U2119 ( .A(n2089), .Z(n2071) );
  NOR U2120 ( .A(n1931), .B(n1930), .Z(n1936) );
  IV U2121 ( .A(n1932), .Z(n1933) );
  NOR U2122 ( .A(n1934), .B(n1933), .Z(n1935) );
  NOR U2123 ( .A(n1936), .B(n1935), .Z(n2094) );
  NOR U2124 ( .A(n1938), .B(n1937), .Z(n1943) );
  IV U2125 ( .A(n1939), .Z(n1941) );
  NOR U2126 ( .A(n1941), .B(n1940), .Z(n1942) );
  NOR U2127 ( .A(n1943), .B(n1942), .Z(n2093) );
  XOR U2128 ( .A(n2094), .B(n2093), .Z(n2095) );
  NOR U2129 ( .A(n1945), .B(n1944), .Z(n1949) );
  NOR U2130 ( .A(n1947), .B(n1946), .Z(n1948) );
  NOR U2131 ( .A(n1949), .B(n1948), .Z(n2104) );
  IV U2132 ( .A(n1950), .Z(n1951) );
  NOR U2133 ( .A(n1952), .B(n1951), .Z(n1956) );
  NOR U2134 ( .A(n1954), .B(n1953), .Z(n1955) );
  NOR U2135 ( .A(n1956), .B(n1955), .Z(n2107) );
  NOR U2136 ( .A(n1958), .B(n1957), .Z(n1963) );
  IV U2137 ( .A(n1959), .Z(n1960) );
  NOR U2138 ( .A(n1961), .B(n1960), .Z(n1962) );
  NOR U2139 ( .A(n1963), .B(n1962), .Z(n1964) );
  IV U2140 ( .A(n1964), .Z(n2108) );
  XOR U2141 ( .A(n2107), .B(n2108), .Z(n2111) );
  NOR U2142 ( .A(n1966), .B(n1965), .Z(n1971) );
  IV U2143 ( .A(n1967), .Z(n1969) );
  NOR U2144 ( .A(n1969), .B(n1968), .Z(n1970) );
  NOR U2145 ( .A(n1971), .B(n1970), .Z(n1972) );
  IV U2146 ( .A(n1972), .Z(n2110) );
  XOR U2147 ( .A(n2111), .B(n2110), .Z(n2101) );
  IV U2148 ( .A(n1973), .Z(n1974) );
  NOR U2149 ( .A(n1975), .B(n1974), .Z(n1980) );
  IV U2150 ( .A(n1976), .Z(n1978) );
  NOR U2151 ( .A(n1978), .B(n1977), .Z(n1979) );
  NOR U2152 ( .A(n1980), .B(n1979), .Z(n2125) );
  IV U2153 ( .A(n1981), .Z(n1982) );
  NOR U2154 ( .A(n1983), .B(n1982), .Z(n1988) );
  IV U2155 ( .A(n1984), .Z(n1985) );
  NOR U2156 ( .A(n1986), .B(n1985), .Z(n1987) );
  NOR U2157 ( .A(n1988), .B(n1987), .Z(n2123) );
  NOR U2158 ( .A(n1990), .B(n1989), .Z(n1995) );
  IV U2159 ( .A(n1991), .Z(n1992) );
  NOR U2160 ( .A(n1993), .B(n1992), .Z(n1994) );
  NOR U2161 ( .A(n1995), .B(n1994), .Z(n2195) );
  NOR U2162 ( .A(n2400), .B(n2309), .Z(n2000) );
  IV U2163 ( .A(n1996), .Z(n1998) );
  NOR U2164 ( .A(n1998), .B(n1997), .Z(n1999) );
  NOR U2165 ( .A(n2000), .B(n1999), .Z(n2193) );
  NOR U2166 ( .A(n3780), .B(n3619), .Z(n2155) );
  NOR U2167 ( .A(n3646), .B(n3776), .Z(n2001) );
  IV U2168 ( .A(n2001), .Z(n2156) );
  XOR U2169 ( .A(n2155), .B(n2156), .Z(n2159) );
  NOR U2170 ( .A(n3625), .B(n3766), .Z(n2251) );
  NOR U2171 ( .A(n3781), .B(n3548), .Z(n2002) );
  IV U2172 ( .A(n2002), .Z(n2250) );
  IV U2173 ( .A(y[23]), .Z(n3750) );
  NOR U2174 ( .A(n3680), .B(n3750), .Z(n2248) );
  XOR U2175 ( .A(n2250), .B(n2248), .Z(n2252) );
  XOR U2176 ( .A(n2251), .B(n2252), .Z(n2158) );
  XOR U2177 ( .A(n2159), .B(n2158), .Z(n2191) );
  XOR U2178 ( .A(n2193), .B(n2191), .Z(n2194) );
  XOR U2179 ( .A(n2195), .B(n2194), .Z(n2121) );
  XOR U2180 ( .A(n2123), .B(n2121), .Z(n2124) );
  XOR U2181 ( .A(n2125), .B(n2124), .Z(n2003) );
  IV U2182 ( .A(n2003), .Z(n2180) );
  NOR U2183 ( .A(n3682), .B(n2764), .Z(n2026) );
  IV U2184 ( .A(n2026), .Z(n2006) );
  IV U2185 ( .A(n2004), .Z(n2005) );
  NOR U2186 ( .A(n2006), .B(n2005), .Z(n2011) );
  IV U2187 ( .A(n2007), .Z(n2008) );
  NOR U2188 ( .A(n2009), .B(n2008), .Z(n2010) );
  NOR U2189 ( .A(n2011), .B(n2010), .Z(n2178) );
  IV U2190 ( .A(n2012), .Z(n2013) );
  NOR U2191 ( .A(n2014), .B(n2013), .Z(n2019) );
  IV U2192 ( .A(n2015), .Z(n2016) );
  NOR U2193 ( .A(n2017), .B(n2016), .Z(n2018) );
  NOR U2194 ( .A(n2019), .B(n2018), .Z(n2173) );
  NOR U2195 ( .A(n3687), .B(n3742), .Z(n2021) );
  NOR U2196 ( .A(n3621), .B(n3647), .Z(n2020) );
  XOR U2197 ( .A(n2021), .B(n2020), .Z(n2215) );
  NOR U2198 ( .A(n3489), .B(n3635), .Z(n2022) );
  IV U2199 ( .A(n2022), .Z(n2152) );
  IV U2200 ( .A(x[23]), .Z(n3461) );
  NOR U2201 ( .A(n3461), .B(n3637), .Z(n2023) );
  XOR U2202 ( .A(n2024), .B(n2023), .Z(n2150) );
  XOR U2203 ( .A(n2152), .B(n2150), .Z(n2217) );
  XOR U2204 ( .A(n2215), .B(n2217), .Z(n2171) );
  NOR U2205 ( .A(n3775), .B(n3748), .Z(n2025) );
  XOR U2206 ( .A(n2026), .B(n2025), .Z(n2143) );
  NOR U2207 ( .A(n3740), .B(n3549), .Z(n2028) );
  XOR U2208 ( .A(n2028), .B(n2027), .Z(n2128) );
  NOR U2209 ( .A(n3688), .B(n3062), .Z(n2029) );
  IV U2210 ( .A(n2029), .Z(n2202) );
  NOR U2211 ( .A(n3529), .B(n3633), .Z(n2031) );
  NOR U2212 ( .A(n3765), .B(n3467), .Z(n2030) );
  XOR U2213 ( .A(n2031), .B(n2030), .Z(n2201) );
  XOR U2214 ( .A(n2202), .B(n2201), .Z(n2130) );
  XOR U2215 ( .A(n2128), .B(n2130), .Z(n2145) );
  XOR U2216 ( .A(n2143), .B(n2145), .Z(n2170) );
  XOR U2217 ( .A(n2171), .B(n2170), .Z(n2032) );
  IV U2218 ( .A(n2032), .Z(n2172) );
  XOR U2219 ( .A(n2173), .B(n2172), .Z(n2186) );
  IV U2220 ( .A(n2033), .Z(n2035) );
  NOR U2221 ( .A(n2035), .B(n2034), .Z(n2039) );
  NOR U2222 ( .A(n2037), .B(n2036), .Z(n2038) );
  NOR U2223 ( .A(n2039), .B(n2038), .Z(n2184) );
  XOR U2224 ( .A(n2186), .B(n2184), .Z(n2187) );
  NOR U2225 ( .A(n3646), .B(n3782), .Z(n2040) );
  IV U2226 ( .A(n2040), .Z(n3497) );
  IV U2227 ( .A(n2041), .Z(n2042) );
  NOR U2228 ( .A(n3497), .B(n2042), .Z(n2047) );
  IV U2229 ( .A(n2043), .Z(n2045) );
  NOR U2230 ( .A(n2045), .B(n2044), .Z(n2046) );
  NOR U2231 ( .A(n2047), .B(n2046), .Z(n2166) );
  NOR U2232 ( .A(n3689), .B(n3628), .Z(n2048) );
  IV U2233 ( .A(n2048), .Z(n2231) );
  NOR U2234 ( .A(n3782), .B(n3787), .Z(n2050) );
  NOR U2235 ( .A(n3746), .B(n3764), .Z(n2049) );
  XOR U2236 ( .A(n2050), .B(n2049), .Z(n2230) );
  XOR U2237 ( .A(n2231), .B(n2230), .Z(n2137) );
  NOR U2238 ( .A(n3161), .B(n3650), .Z(n2133) );
  NOR U2239 ( .A(n3546), .B(n3622), .Z(n2051) );
  IV U2240 ( .A(n2051), .Z(n2134) );
  XOR U2241 ( .A(n2133), .B(n2134), .Z(n2136) );
  XOR U2242 ( .A(n2137), .B(n2136), .Z(n2162) );
  IV U2243 ( .A(o[22]), .Z(n2053) );
  NOR U2244 ( .A(n2053), .B(n2052), .Z(n2242) );
  NOR U2245 ( .A(n3645), .B(n3773), .Z(n2054) );
  IV U2246 ( .A(n2054), .Z(n2226) );
  XOR U2247 ( .A(n2226), .B(o[23]), .Z(n2241) );
  XOR U2248 ( .A(n2055), .B(n2241), .Z(n2244) );
  XOR U2249 ( .A(n2242), .B(n2244), .Z(n2163) );
  XOR U2250 ( .A(n2162), .B(n2163), .Z(n2165) );
  XOR U2251 ( .A(n2166), .B(n2165), .Z(n2188) );
  XOR U2252 ( .A(n2187), .B(n2188), .Z(n2118) );
  NOR U2253 ( .A(n3489), .B(n3765), .Z(n3162) );
  IV U2254 ( .A(n3162), .Z(n2058) );
  IV U2255 ( .A(n2056), .Z(n2057) );
  NOR U2256 ( .A(n2058), .B(n2057), .Z(n2063) );
  IV U2257 ( .A(n2059), .Z(n2060) );
  NOR U2258 ( .A(n2061), .B(n2060), .Z(n2062) );
  NOR U2259 ( .A(n2063), .B(n2062), .Z(n2115) );
  IV U2260 ( .A(n2064), .Z(n2066) );
  NOR U2261 ( .A(n2066), .B(n2065), .Z(n2070) );
  NOR U2262 ( .A(n2068), .B(n2067), .Z(n2069) );
  NOR U2263 ( .A(n2070), .B(n2069), .Z(n2114) );
  XOR U2264 ( .A(n2115), .B(n2114), .Z(n2116) );
  XOR U2265 ( .A(n2118), .B(n2116), .Z(n2177) );
  XOR U2266 ( .A(n2178), .B(n2177), .Z(n2179) );
  XOR U2267 ( .A(n2180), .B(n2179), .Z(n2100) );
  XOR U2268 ( .A(n2101), .B(n2100), .Z(n2102) );
  XOR U2269 ( .A(n2104), .B(n2102), .Z(n2096) );
  XOR U2270 ( .A(n2095), .B(n2096), .Z(n2090) );
  XOR U2271 ( .A(n2071), .B(n2090), .Z(n2081) );
  XOR U2272 ( .A(n2079), .B(n2081), .Z(n2082) );
  XOR U2273 ( .A(n2083), .B(n2082), .Z(n2072) );
  XOR U2274 ( .A(n2073), .B(n2072), .Z(n2074) );
  XOR U2275 ( .A(n2076), .B(n2074), .Z(N56) );
  NOR U2276 ( .A(n2073), .B(n2072), .Z(n2078) );
  IV U2277 ( .A(n2074), .Z(n2075) );
  NOR U2278 ( .A(n2076), .B(n2075), .Z(n2077) );
  NOR U2279 ( .A(n2078), .B(n2077), .Z(n2443) );
  IV U2280 ( .A(n2443), .Z(n2257) );
  IV U2281 ( .A(n2079), .Z(n2080) );
  NOR U2282 ( .A(n2081), .B(n2080), .Z(n2085) );
  NOR U2283 ( .A(n2083), .B(n2082), .Z(n2084) );
  NOR U2284 ( .A(n2085), .B(n2084), .Z(n2439) );
  IV U2285 ( .A(n2086), .Z(n2087) );
  NOR U2286 ( .A(n2088), .B(n2087), .Z(n2092) );
  NOR U2287 ( .A(n2090), .B(n2089), .Z(n2091) );
  NOR U2288 ( .A(n2092), .B(n2091), .Z(n2261) );
  NOR U2289 ( .A(n2094), .B(n2093), .Z(n2099) );
  IV U2290 ( .A(n2095), .Z(n2097) );
  NOR U2291 ( .A(n2097), .B(n2096), .Z(n2098) );
  NOR U2292 ( .A(n2099), .B(n2098), .Z(n2258) );
  NOR U2293 ( .A(n2101), .B(n2100), .Z(n2106) );
  IV U2294 ( .A(n2102), .Z(n2103) );
  NOR U2295 ( .A(n2104), .B(n2103), .Z(n2105) );
  NOR U2296 ( .A(n2106), .B(n2105), .Z(n2269) );
  IV U2297 ( .A(n2107), .Z(n2109) );
  NOR U2298 ( .A(n2109), .B(n2108), .Z(n2113) );
  NOR U2299 ( .A(n2111), .B(n2110), .Z(n2112) );
  NOR U2300 ( .A(n2113), .B(n2112), .Z(n2268) );
  NOR U2301 ( .A(n2115), .B(n2114), .Z(n2120) );
  IV U2302 ( .A(n2116), .Z(n2117) );
  NOR U2303 ( .A(n2118), .B(n2117), .Z(n2119) );
  NOR U2304 ( .A(n2120), .B(n2119), .Z(n2284) );
  IV U2305 ( .A(n2121), .Z(n2122) );
  NOR U2306 ( .A(n2123), .B(n2122), .Z(n2127) );
  NOR U2307 ( .A(n2125), .B(n2124), .Z(n2126) );
  NOR U2308 ( .A(n2127), .B(n2126), .Z(n2281) );
  NOR U2309 ( .A(n3022), .B(n2423), .Z(n2132) );
  IV U2310 ( .A(n2128), .Z(n2129) );
  NOR U2311 ( .A(n2130), .B(n2129), .Z(n2131) );
  NOR U2312 ( .A(n2132), .B(n2131), .Z(n2297) );
  IV U2313 ( .A(n2297), .Z(n2140) );
  IV U2314 ( .A(n2133), .Z(n2135) );
  NOR U2315 ( .A(n2135), .B(n2134), .Z(n2139) );
  NOR U2316 ( .A(n2137), .B(n2136), .Z(n2138) );
  NOR U2317 ( .A(n2139), .B(n2138), .Z(n2296) );
  XOR U2318 ( .A(n2140), .B(n2296), .Z(n2299) );
  NOR U2319 ( .A(n3682), .B(n3775), .Z(n2210) );
  IV U2320 ( .A(n2210), .Z(n2334) );
  IV U2321 ( .A(n2141), .Z(n2142) );
  NOR U2322 ( .A(n2334), .B(n2142), .Z(n2147) );
  IV U2323 ( .A(n2143), .Z(n2144) );
  NOR U2324 ( .A(n2145), .B(n2144), .Z(n2146) );
  NOR U2325 ( .A(n2147), .B(n2146), .Z(n2375) );
  NOR U2326 ( .A(n3461), .B(n3462), .Z(n3751) );
  IV U2327 ( .A(n3751), .Z(n2149) );
  NOR U2328 ( .A(n2149), .B(n2148), .Z(n2154) );
  IV U2329 ( .A(n2150), .Z(n2151) );
  NOR U2330 ( .A(n2152), .B(n2151), .Z(n2153) );
  NOR U2331 ( .A(n2154), .B(n2153), .Z(n2372) );
  IV U2332 ( .A(n2155), .Z(n2157) );
  NOR U2333 ( .A(n2157), .B(n2156), .Z(n2161) );
  NOR U2334 ( .A(n2159), .B(n2158), .Z(n2160) );
  NOR U2335 ( .A(n2161), .B(n2160), .Z(n2371) );
  XOR U2336 ( .A(n2372), .B(n2371), .Z(n2373) );
  XOR U2337 ( .A(n2375), .B(n2373), .Z(n2298) );
  XOR U2338 ( .A(n2299), .B(n2298), .Z(n2360) );
  IV U2339 ( .A(n2162), .Z(n2164) );
  NOR U2340 ( .A(n2164), .B(n2163), .Z(n2168) );
  NOR U2341 ( .A(n2166), .B(n2165), .Z(n2167) );
  NOR U2342 ( .A(n2168), .B(n2167), .Z(n2169) );
  IV U2343 ( .A(n2169), .Z(n2358) );
  NOR U2344 ( .A(n2171), .B(n2170), .Z(n2175) );
  NOR U2345 ( .A(n2173), .B(n2172), .Z(n2174) );
  NOR U2346 ( .A(n2175), .B(n2174), .Z(n2356) );
  XOR U2347 ( .A(n2358), .B(n2356), .Z(n2359) );
  XOR U2348 ( .A(n2360), .B(n2359), .Z(n2176) );
  IV U2349 ( .A(n2176), .Z(n2283) );
  XOR U2350 ( .A(n2281), .B(n2283), .Z(n2286) );
  XOR U2351 ( .A(n2284), .B(n2286), .Z(n2277) );
  NOR U2352 ( .A(n2178), .B(n2177), .Z(n2183) );
  IV U2353 ( .A(n2179), .Z(n2181) );
  NOR U2354 ( .A(n2181), .B(n2180), .Z(n2182) );
  NOR U2355 ( .A(n2183), .B(n2182), .Z(n2274) );
  IV U2356 ( .A(n2184), .Z(n2185) );
  NOR U2357 ( .A(n2186), .B(n2185), .Z(n2190) );
  NOR U2358 ( .A(n2188), .B(n2187), .Z(n2189) );
  NOR U2359 ( .A(n2190), .B(n2189), .Z(n2293) );
  IV U2360 ( .A(n2293), .Z(n2256) );
  IV U2361 ( .A(n2191), .Z(n2192) );
  NOR U2362 ( .A(n2193), .B(n2192), .Z(n2197) );
  NOR U2363 ( .A(n2195), .B(n2194), .Z(n2196) );
  NOR U2364 ( .A(n2197), .B(n2196), .Z(n2289) );
  NOR U2365 ( .A(n3529), .B(n3467), .Z(n3642) );
  IV U2366 ( .A(n3642), .Z(n2200) );
  IV U2367 ( .A(n2198), .Z(n2199) );
  NOR U2368 ( .A(n2200), .B(n2199), .Z(n2205) );
  IV U2369 ( .A(n2201), .Z(n2203) );
  NOR U2370 ( .A(n2203), .B(n2202), .Z(n2204) );
  NOR U2371 ( .A(n2205), .B(n2204), .Z(n2352) );
  NOR U2372 ( .A(n3549), .B(n3748), .Z(n2424) );
  NOR U2373 ( .A(n3740), .B(n3161), .Z(n2206) );
  IV U2374 ( .A(n2206), .Z(n2208) );
  XOR U2375 ( .A(n2208), .B(n2207), .Z(n2426) );
  XOR U2376 ( .A(n2424), .B(n2426), .Z(n2335) );
  NOR U2377 ( .A(n3689), .B(n3746), .Z(n2209) );
  IV U2378 ( .A(n2209), .Z(n2333) );
  XOR U2379 ( .A(n2333), .B(n2210), .Z(n2336) );
  XOR U2380 ( .A(n2335), .B(n2336), .Z(n2348) );
  NOR U2381 ( .A(n3621), .B(n3787), .Z(n2211) );
  XOR U2382 ( .A(n2212), .B(n2211), .Z(n2317) );
  NOR U2383 ( .A(n3645), .B(n3647), .Z(n2409) );
  NOR U2384 ( .A(n3766), .B(n3619), .Z(n2213) );
  IV U2385 ( .A(n2213), .Z(n2408) );
  NOR U2386 ( .A(n3465), .B(n3646), .Z(n2406) );
  XOR U2387 ( .A(n2408), .B(n2406), .Z(n2411) );
  XOR U2388 ( .A(n2409), .B(n2411), .Z(n2319) );
  XOR U2389 ( .A(n2317), .B(n2319), .Z(n2350) );
  XOR U2390 ( .A(n2348), .B(n2350), .Z(n2351) );
  XOR U2391 ( .A(n2352), .B(n2351), .Z(n2365) );
  NOR U2392 ( .A(n3181), .B(n2214), .Z(n2219) );
  IV U2393 ( .A(n2215), .Z(n2216) );
  NOR U2394 ( .A(n2217), .B(n2216), .Z(n2218) );
  NOR U2395 ( .A(n2219), .B(n2218), .Z(n2363) );
  XOR U2396 ( .A(n2365), .B(n2363), .Z(n2368) );
  NOR U2397 ( .A(n3776), .B(n3622), .Z(n2393) );
  IV U2398 ( .A(x[24]), .Z(n3686) );
  NOR U2399 ( .A(n3637), .B(n3686), .Z(n2220) );
  IV U2400 ( .A(n2220), .Z(n2394) );
  XOR U2401 ( .A(n2393), .B(n2394), .Z(n2397) );
  NOR U2402 ( .A(n3625), .B(n3750), .Z(n2325) );
  IV U2403 ( .A(y[24]), .Z(n3683) );
  NOR U2404 ( .A(n3680), .B(n3683), .Z(n2221) );
  IV U2405 ( .A(n2221), .Z(n2324) );
  XOR U2406 ( .A(n2324), .B(n2222), .Z(n2327) );
  XOR U2407 ( .A(n2325), .B(n2327), .Z(n2396) );
  XOR U2408 ( .A(n2397), .B(n2396), .Z(n2342) );
  NOR U2409 ( .A(n3546), .B(n3781), .Z(n2223) );
  IV U2410 ( .A(n2223), .Z(n2225) );
  XOR U2411 ( .A(n2225), .B(n2224), .Z(n2419) );
  XOR U2412 ( .A(n2419), .B(n2420), .Z(n2339) );
  IV U2413 ( .A(o[23]), .Z(n2227) );
  NOR U2414 ( .A(n2227), .B(n2226), .Z(n2388) );
  NOR U2415 ( .A(n3062), .B(n3763), .Z(n2385) );
  NOR U2416 ( .A(n3773), .B(n3461), .Z(n2228) );
  IV U2417 ( .A(n2228), .Z(n2415) );
  XOR U2418 ( .A(n2415), .B(o[24]), .Z(n2386) );
  XOR U2419 ( .A(n2385), .B(n2386), .Z(n2390) );
  XOR U2420 ( .A(n2388), .B(n2390), .Z(n2341) );
  XOR U2421 ( .A(n2339), .B(n2341), .Z(n2343) );
  XOR U2422 ( .A(n2342), .B(n2343), .Z(n2382) );
  NOR U2423 ( .A(n3746), .B(n3782), .Z(n2437) );
  IV U2424 ( .A(n2437), .Z(n2601) );
  NOR U2425 ( .A(n2601), .B(n2229), .Z(n2234) );
  IV U2426 ( .A(n2230), .Z(n2232) );
  NOR U2427 ( .A(n2232), .B(n2231), .Z(n2233) );
  NOR U2428 ( .A(n2234), .B(n2233), .Z(n2380) );
  NOR U2429 ( .A(n3780), .B(n3635), .Z(n2401) );
  NOR U2430 ( .A(n3462), .B(n3742), .Z(n2235) );
  IV U2431 ( .A(n2235), .Z(n2237) );
  NOR U2432 ( .A(n3628), .B(n3782), .Z(n2236) );
  XOR U2433 ( .A(n2237), .B(n2236), .Z(n2403) );
  XOR U2434 ( .A(n2401), .B(n2403), .Z(n2312) );
  NOR U2435 ( .A(n3489), .B(n3650), .Z(n2238) );
  IV U2436 ( .A(n2238), .Z(n2310) );
  XOR U2437 ( .A(n2310), .B(n2239), .Z(n2311) );
  XOR U2438 ( .A(n2312), .B(n2311), .Z(n2378) );
  XOR U2439 ( .A(n2380), .B(n2378), .Z(n2381) );
  XOR U2440 ( .A(n2382), .B(n2381), .Z(n2306) );
  NOR U2441 ( .A(n2241), .B(n2240), .Z(n2246) );
  IV U2442 ( .A(n2242), .Z(n2243) );
  NOR U2443 ( .A(n2244), .B(n2243), .Z(n2245) );
  NOR U2444 ( .A(n2246), .B(n2245), .Z(n2247) );
  IV U2445 ( .A(n2247), .Z(n2304) );
  IV U2446 ( .A(n2248), .Z(n2249) );
  NOR U2447 ( .A(n2250), .B(n2249), .Z(n2255) );
  IV U2448 ( .A(n2251), .Z(n2253) );
  NOR U2449 ( .A(n2253), .B(n2252), .Z(n2254) );
  NOR U2450 ( .A(n2255), .B(n2254), .Z(n2302) );
  XOR U2451 ( .A(n2304), .B(n2302), .Z(n2305) );
  XOR U2452 ( .A(n2306), .B(n2305), .Z(n2366) );
  XOR U2453 ( .A(n2368), .B(n2366), .Z(n2290) );
  XOR U2454 ( .A(n2289), .B(n2290), .Z(n2292) );
  XOR U2455 ( .A(n2256), .B(n2292), .Z(n2276) );
  XOR U2456 ( .A(n2274), .B(n2276), .Z(n2278) );
  XOR U2457 ( .A(n2277), .B(n2278), .Z(n2266) );
  XOR U2458 ( .A(n2268), .B(n2266), .Z(n2271) );
  XOR U2459 ( .A(n2269), .B(n2271), .Z(n2260) );
  XOR U2460 ( .A(n2258), .B(n2260), .Z(n2263) );
  XOR U2461 ( .A(n2261), .B(n2263), .Z(n2441) );
  XOR U2462 ( .A(n2439), .B(n2441), .Z(n2442) );
  XOR U2463 ( .A(n2257), .B(n2442), .Z(N57) );
  IV U2464 ( .A(n2258), .Z(n2259) );
  NOR U2465 ( .A(n2260), .B(n2259), .Z(n2265) );
  IV U2466 ( .A(n2261), .Z(n2262) );
  NOR U2467 ( .A(n2263), .B(n2262), .Z(n2264) );
  NOR U2468 ( .A(n2265), .B(n2264), .Z(n2447) );
  IV U2469 ( .A(n2266), .Z(n2267) );
  NOR U2470 ( .A(n2268), .B(n2267), .Z(n2273) );
  IV U2471 ( .A(n2269), .Z(n2270) );
  NOR U2472 ( .A(n2271), .B(n2270), .Z(n2272) );
  NOR U2473 ( .A(n2273), .B(n2272), .Z(n2457) );
  IV U2474 ( .A(n2274), .Z(n2275) );
  NOR U2475 ( .A(n2276), .B(n2275), .Z(n2280) );
  NOR U2476 ( .A(n2278), .B(n2277), .Z(n2279) );
  NOR U2477 ( .A(n2280), .B(n2279), .Z(n2454) );
  IV U2478 ( .A(n2281), .Z(n2282) );
  NOR U2479 ( .A(n2283), .B(n2282), .Z(n2288) );
  IV U2480 ( .A(n2284), .Z(n2285) );
  NOR U2481 ( .A(n2286), .B(n2285), .Z(n2287) );
  NOR U2482 ( .A(n2288), .B(n2287), .Z(n2464) );
  IV U2483 ( .A(n2289), .Z(n2291) );
  NOR U2484 ( .A(n2291), .B(n2290), .Z(n2295) );
  NOR U2485 ( .A(n2293), .B(n2292), .Z(n2294) );
  NOR U2486 ( .A(n2295), .B(n2294), .Z(n2473) );
  NOR U2487 ( .A(n2297), .B(n2296), .Z(n2301) );
  NOR U2488 ( .A(n2299), .B(n2298), .Z(n2300) );
  NOR U2489 ( .A(n2301), .B(n2300), .Z(n2469) );
  IV U2490 ( .A(n2302), .Z(n2303) );
  NOR U2491 ( .A(n2304), .B(n2303), .Z(n2308) );
  NOR U2492 ( .A(n2306), .B(n2305), .Z(n2307) );
  NOR U2493 ( .A(n2308), .B(n2307), .Z(n2634) );
  IV U2494 ( .A(n2634), .Z(n2355) );
  NOR U2495 ( .A(n2310), .B(n2309), .Z(n2314) );
  NOR U2496 ( .A(n2312), .B(n2311), .Z(n2313) );
  NOR U2497 ( .A(n2314), .B(n2313), .Z(n2485) );
  IV U2498 ( .A(n2315), .Z(n2316) );
  NOR U2499 ( .A(n3181), .B(n2316), .Z(n2321) );
  IV U2500 ( .A(n2317), .Z(n2318) );
  NOR U2501 ( .A(n2319), .B(n2318), .Z(n2320) );
  NOR U2502 ( .A(n2321), .B(n2320), .Z(n2484) );
  XOR U2503 ( .A(n2485), .B(n2484), .Z(n2322) );
  IV U2504 ( .A(n2322), .Z(n2486) );
  NOR U2505 ( .A(n2324), .B(n2323), .Z(n2329) );
  IV U2506 ( .A(n2325), .Z(n2326) );
  NOR U2507 ( .A(n2327), .B(n2326), .Z(n2328) );
  NOR U2508 ( .A(n2329), .B(n2328), .Z(n2517) );
  IV U2509 ( .A(x[25]), .Z(n3634) );
  NOR U2510 ( .A(n3637), .B(n3634), .Z(n2572) );
  NOR U2511 ( .A(n3781), .B(n3776), .Z(n2330) );
  IV U2512 ( .A(n2330), .Z(n2573) );
  XOR U2513 ( .A(n2572), .B(n2573), .Z(n2576) );
  NOR U2514 ( .A(n3625), .B(n3683), .Z(n2538) );
  IV U2515 ( .A(y[25]), .Z(n3747) );
  NOR U2516 ( .A(n3680), .B(n3747), .Z(n2331) );
  IV U2517 ( .A(n2331), .Z(n2537) );
  NOR U2518 ( .A(n3465), .B(n3622), .Z(n2535) );
  XOR U2519 ( .A(n2537), .B(n2535), .Z(n2540) );
  XOR U2520 ( .A(n2538), .B(n2540), .Z(n2575) );
  XOR U2521 ( .A(n2576), .B(n2575), .Z(n2513) );
  NOR U2522 ( .A(n3161), .B(n3748), .Z(n2610) );
  NOR U2523 ( .A(n3628), .B(n3621), .Z(n2609) );
  XOR U2524 ( .A(n2610), .B(n2609), .Z(n2612) );
  NOR U2525 ( .A(n3489), .B(n3740), .Z(n2583) );
  NOR U2526 ( .A(n3780), .B(n3650), .Z(n2332) );
  IV U2527 ( .A(n2332), .Z(n2582) );
  NOR U2528 ( .A(n3633), .B(n3689), .Z(n2580) );
  XOR U2529 ( .A(n2582), .B(n2580), .Z(n2585) );
  XOR U2530 ( .A(n2583), .B(n2585), .Z(n2613) );
  XOR U2531 ( .A(n2612), .B(n2613), .Z(n2514) );
  XOR U2532 ( .A(n2513), .B(n2514), .Z(n2516) );
  XOR U2533 ( .A(n2517), .B(n2516), .Z(n2492) );
  NOR U2534 ( .A(n2334), .B(n2333), .Z(n2338) );
  NOR U2535 ( .A(n2336), .B(n2335), .Z(n2337) );
  NOR U2536 ( .A(n2338), .B(n2337), .Z(n2490) );
  XOR U2537 ( .A(n2492), .B(n2490), .Z(n2494) );
  IV U2538 ( .A(n2339), .Z(n2340) );
  NOR U2539 ( .A(n2341), .B(n2340), .Z(n2346) );
  IV U2540 ( .A(n2342), .Z(n2344) );
  NOR U2541 ( .A(n2344), .B(n2343), .Z(n2345) );
  NOR U2542 ( .A(n2346), .B(n2345), .Z(n2347) );
  IV U2543 ( .A(n2347), .Z(n2493) );
  XOR U2544 ( .A(n2494), .B(n2493), .Z(n2487) );
  XOR U2545 ( .A(n2486), .B(n2487), .Z(n2632) );
  IV U2546 ( .A(n2348), .Z(n2349) );
  NOR U2547 ( .A(n2350), .B(n2349), .Z(n2354) );
  NOR U2548 ( .A(n2352), .B(n2351), .Z(n2353) );
  NOR U2549 ( .A(n2354), .B(n2353), .Z(n2630) );
  XOR U2550 ( .A(n2632), .B(n2630), .Z(n2633) );
  XOR U2551 ( .A(n2355), .B(n2633), .Z(n2470) );
  XOR U2552 ( .A(n2469), .B(n2470), .Z(n2472) );
  XOR U2553 ( .A(n2473), .B(n2472), .Z(n2463) );
  IV U2554 ( .A(n2463), .Z(n2438) );
  IV U2555 ( .A(n2356), .Z(n2357) );
  NOR U2556 ( .A(n2358), .B(n2357), .Z(n2362) );
  NOR U2557 ( .A(n2360), .B(n2359), .Z(n2361) );
  NOR U2558 ( .A(n2362), .B(n2361), .Z(n2479) );
  IV U2559 ( .A(n2363), .Z(n2364) );
  NOR U2560 ( .A(n2365), .B(n2364), .Z(n2370) );
  IV U2561 ( .A(n2366), .Z(n2367) );
  NOR U2562 ( .A(n2368), .B(n2367), .Z(n2369) );
  NOR U2563 ( .A(n2370), .B(n2369), .Z(n2476) );
  NOR U2564 ( .A(n2372), .B(n2371), .Z(n2377) );
  IV U2565 ( .A(n2373), .Z(n2374) );
  NOR U2566 ( .A(n2375), .B(n2374), .Z(n2376) );
  NOR U2567 ( .A(n2377), .B(n2376), .Z(n2641) );
  IV U2568 ( .A(n2378), .Z(n2379) );
  NOR U2569 ( .A(n2380), .B(n2379), .Z(n2384) );
  NOR U2570 ( .A(n2382), .B(n2381), .Z(n2383) );
  NOR U2571 ( .A(n2384), .B(n2383), .Z(n2638) );
  IV U2572 ( .A(n2385), .Z(n2387) );
  NOR U2573 ( .A(n2387), .B(n2386), .Z(n2392) );
  IV U2574 ( .A(n2388), .Z(n2389) );
  NOR U2575 ( .A(n2390), .B(n2389), .Z(n2391) );
  NOR U2576 ( .A(n2392), .B(n2391), .Z(n2646) );
  IV U2577 ( .A(n2393), .Z(n2395) );
  NOR U2578 ( .A(n2395), .B(n2394), .Z(n2399) );
  NOR U2579 ( .A(n2397), .B(n2396), .Z(n2398) );
  NOR U2580 ( .A(n2399), .B(n2398), .Z(n2645) );
  XOR U2581 ( .A(n2646), .B(n2645), .Z(n2647) );
  NOR U2582 ( .A(n3193), .B(n2400), .Z(n2405) );
  IV U2583 ( .A(n2401), .Z(n2402) );
  NOR U2584 ( .A(n2403), .B(n2402), .Z(n2404) );
  NOR U2585 ( .A(n2405), .B(n2404), .Z(n2627) );
  IV U2586 ( .A(n2406), .Z(n2407) );
  NOR U2587 ( .A(n2408), .B(n2407), .Z(n2413) );
  IV U2588 ( .A(n2409), .Z(n2410) );
  NOR U2589 ( .A(n2411), .B(n2410), .Z(n2412) );
  NOR U2590 ( .A(n2413), .B(n2412), .Z(n2625) );
  IV U2591 ( .A(o[24]), .Z(n2414) );
  NOR U2592 ( .A(n2415), .B(n2414), .Z(n2567) );
  NOR U2593 ( .A(n3062), .B(n3467), .Z(n2564) );
  NOR U2594 ( .A(n3773), .B(n3686), .Z(n2416) );
  IV U2595 ( .A(n2416), .Z(n2555) );
  XOR U2596 ( .A(n2555), .B(o[25]), .Z(n2565) );
  XOR U2597 ( .A(n2564), .B(n2565), .Z(n2569) );
  XOR U2598 ( .A(n2567), .B(n2569), .Z(n2624) );
  XOR U2599 ( .A(n2625), .B(n2624), .Z(n2417) );
  IV U2600 ( .A(n2417), .Z(n2626) );
  XOR U2601 ( .A(n2627), .B(n2626), .Z(n2500) );
  NOR U2602 ( .A(n3546), .B(n3467), .Z(n2730) );
  IV U2603 ( .A(n2730), .Z(n3037) );
  NOR U2604 ( .A(n3037), .B(n2418), .Z(n2422) );
  NOR U2605 ( .A(n2420), .B(n2419), .Z(n2421) );
  NOR U2606 ( .A(n2422), .B(n2421), .Z(n2499) );
  NOR U2607 ( .A(n3765), .B(n3161), .Z(n3060) );
  IV U2608 ( .A(n3060), .Z(n3490) );
  NOR U2609 ( .A(n3490), .B(n2423), .Z(n2428) );
  IV U2610 ( .A(n2424), .Z(n2425) );
  NOR U2611 ( .A(n2426), .B(n2425), .Z(n2427) );
  NOR U2612 ( .A(n2428), .B(n2427), .Z(n2509) );
  NOR U2613 ( .A(n3766), .B(n3635), .Z(n2429) );
  IV U2614 ( .A(n2429), .Z(n2522) );
  NOR U2615 ( .A(n3529), .B(n3462), .Z(n2520) );
  XOR U2616 ( .A(n2522), .B(n2520), .Z(n2524) );
  NOR U2617 ( .A(n3461), .B(n3647), .Z(n2596) );
  NOR U2618 ( .A(n3750), .B(n3619), .Z(n2430) );
  IV U2619 ( .A(n2430), .Z(n2595) );
  XOR U2620 ( .A(n2595), .B(n2431), .Z(n2597) );
  XOR U2621 ( .A(n2596), .B(n2597), .Z(n2523) );
  XOR U2622 ( .A(n2524), .B(n2523), .Z(n2505) );
  NOR U2623 ( .A(n3646), .B(n3742), .Z(n2617) );
  NOR U2624 ( .A(n3749), .B(n3775), .Z(n2432) );
  IV U2625 ( .A(n2432), .Z(n2618) );
  XOR U2626 ( .A(n2617), .B(n2618), .Z(n2621) );
  NOR U2627 ( .A(n3645), .B(n3787), .Z(n2530) );
  NOR U2628 ( .A(n3687), .B(n3764), .Z(n2433) );
  IV U2629 ( .A(n2433), .Z(n2529) );
  NOR U2630 ( .A(n3682), .B(n3549), .Z(n2527) );
  XOR U2631 ( .A(n2529), .B(n2527), .Z(n2532) );
  XOR U2632 ( .A(n2530), .B(n2532), .Z(n2620) );
  XOR U2633 ( .A(n2621), .B(n2620), .Z(n2603) );
  NOR U2634 ( .A(n3765), .B(n2764), .Z(n2741) );
  XOR U2635 ( .A(n2741), .B(n2434), .Z(n2435) );
  IV U2636 ( .A(n2435), .Z(n2552) );
  XOR U2637 ( .A(n2552), .B(n2436), .Z(n2602) );
  XOR U2638 ( .A(n2437), .B(n2602), .Z(n2604) );
  XOR U2639 ( .A(n2603), .B(n2604), .Z(n2506) );
  XOR U2640 ( .A(n2505), .B(n2506), .Z(n2508) );
  XOR U2641 ( .A(n2509), .B(n2508), .Z(n2497) );
  XOR U2642 ( .A(n2499), .B(n2497), .Z(n2501) );
  XOR U2643 ( .A(n2500), .B(n2501), .Z(n2648) );
  XOR U2644 ( .A(n2647), .B(n2648), .Z(n2637) );
  XOR U2645 ( .A(n2638), .B(n2637), .Z(n2639) );
  XOR U2646 ( .A(n2641), .B(n2639), .Z(n2478) );
  XOR U2647 ( .A(n2476), .B(n2478), .Z(n2480) );
  XOR U2648 ( .A(n2479), .B(n2480), .Z(n2462) );
  XOR U2649 ( .A(n2438), .B(n2462), .Z(n2465) );
  XOR U2650 ( .A(n2464), .B(n2465), .Z(n2456) );
  XOR U2651 ( .A(n2454), .B(n2456), .Z(n2458) );
  XOR U2652 ( .A(n2457), .B(n2458), .Z(n2449) );
  XOR U2653 ( .A(n2447), .B(n2449), .Z(n2451) );
  IV U2654 ( .A(n2439), .Z(n2440) );
  NOR U2655 ( .A(n2441), .B(n2440), .Z(n2445) );
  NOR U2656 ( .A(n2443), .B(n2442), .Z(n2444) );
  NOR U2657 ( .A(n2445), .B(n2444), .Z(n2446) );
  IV U2658 ( .A(n2446), .Z(n2450) );
  XOR U2659 ( .A(n2451), .B(n2450), .Z(N58) );
  IV U2660 ( .A(n2447), .Z(n2448) );
  NOR U2661 ( .A(n2449), .B(n2448), .Z(n2453) );
  NOR U2662 ( .A(n2451), .B(n2450), .Z(n2452) );
  NOR U2663 ( .A(n2453), .B(n2452), .Z(n2856) );
  IV U2664 ( .A(n2454), .Z(n2455) );
  NOR U2665 ( .A(n2456), .B(n2455), .Z(n2461) );
  IV U2666 ( .A(n2457), .Z(n2459) );
  NOR U2667 ( .A(n2459), .B(n2458), .Z(n2460) );
  NOR U2668 ( .A(n2461), .B(n2460), .Z(n2853) );
  NOR U2669 ( .A(n2463), .B(n2462), .Z(n2468) );
  IV U2670 ( .A(n2464), .Z(n2466) );
  NOR U2671 ( .A(n2466), .B(n2465), .Z(n2467) );
  NOR U2672 ( .A(n2468), .B(n2467), .Z(n2655) );
  IV U2673 ( .A(n2469), .Z(n2471) );
  NOR U2674 ( .A(n2471), .B(n2470), .Z(n2475) );
  NOR U2675 ( .A(n2473), .B(n2472), .Z(n2474) );
  NOR U2676 ( .A(n2475), .B(n2474), .Z(n2654) );
  IV U2677 ( .A(n2654), .Z(n2652) );
  IV U2678 ( .A(n2476), .Z(n2477) );
  NOR U2679 ( .A(n2478), .B(n2477), .Z(n2483) );
  IV U2680 ( .A(n2479), .Z(n2481) );
  NOR U2681 ( .A(n2481), .B(n2480), .Z(n2482) );
  NOR U2682 ( .A(n2483), .B(n2482), .Z(n2663) );
  NOR U2683 ( .A(n2485), .B(n2484), .Z(n2489) );
  NOR U2684 ( .A(n2487), .B(n2486), .Z(n2488) );
  NOR U2685 ( .A(n2489), .B(n2488), .Z(n2678) );
  IV U2686 ( .A(n2490), .Z(n2491) );
  NOR U2687 ( .A(n2492), .B(n2491), .Z(n2496) );
  NOR U2688 ( .A(n2494), .B(n2493), .Z(n2495) );
  NOR U2689 ( .A(n2496), .B(n2495), .Z(n2677) );
  IV U2690 ( .A(n2497), .Z(n2498) );
  NOR U2691 ( .A(n2499), .B(n2498), .Z(n2504) );
  IV U2692 ( .A(n2500), .Z(n2502) );
  NOR U2693 ( .A(n2502), .B(n2501), .Z(n2503) );
  NOR U2694 ( .A(n2504), .B(n2503), .Z(n2691) );
  IV U2695 ( .A(n2505), .Z(n2507) );
  NOR U2696 ( .A(n2507), .B(n2506), .Z(n2511) );
  NOR U2697 ( .A(n2509), .B(n2508), .Z(n2510) );
  NOR U2698 ( .A(n2511), .B(n2510), .Z(n2512) );
  IV U2699 ( .A(n2512), .Z(n2692) );
  XOR U2700 ( .A(n2691), .B(n2692), .Z(n2695) );
  IV U2701 ( .A(n2513), .Z(n2515) );
  NOR U2702 ( .A(n2515), .B(n2514), .Z(n2519) );
  NOR U2703 ( .A(n2517), .B(n2516), .Z(n2518) );
  NOR U2704 ( .A(n2519), .B(n2518), .Z(n2686) );
  IV U2705 ( .A(n2520), .Z(n2521) );
  NOR U2706 ( .A(n2522), .B(n2521), .Z(n2526) );
  NOR U2707 ( .A(n2524), .B(n2523), .Z(n2525) );
  NOR U2708 ( .A(n2526), .B(n2525), .Z(n2699) );
  IV U2709 ( .A(n2527), .Z(n2528) );
  NOR U2710 ( .A(n2529), .B(n2528), .Z(n2534) );
  IV U2711 ( .A(n2530), .Z(n2531) );
  NOR U2712 ( .A(n2532), .B(n2531), .Z(n2533) );
  NOR U2713 ( .A(n2534), .B(n2533), .Z(n2845) );
  IV U2714 ( .A(n2535), .Z(n2536) );
  NOR U2715 ( .A(n2537), .B(n2536), .Z(n2542) );
  IV U2716 ( .A(n2538), .Z(n2539) );
  NOR U2717 ( .A(n2540), .B(n2539), .Z(n2541) );
  NOR U2718 ( .A(n2542), .B(n2541), .Z(n2738) );
  NOR U2719 ( .A(n3646), .B(n3529), .Z(n2704) );
  NOR U2720 ( .A(n3787), .B(n3461), .Z(n2543) );
  IV U2721 ( .A(n2543), .Z(n2705) );
  XOR U2722 ( .A(n2704), .B(n2705), .Z(n2708) );
  NOR U2723 ( .A(n3645), .B(n3628), .Z(n2544) );
  IV U2724 ( .A(n2544), .Z(n2707) );
  XOR U2725 ( .A(n2708), .B(n2707), .Z(n2787) );
  NOR U2726 ( .A(n3546), .B(n3763), .Z(n2782) );
  IV U2727 ( .A(n2782), .Z(n2784) );
  XOR U2728 ( .A(n2785), .B(n2784), .Z(n2545) );
  XOR U2729 ( .A(n2787), .B(n2545), .Z(n2734) );
  NOR U2730 ( .A(n3689), .B(n3687), .Z(n2804) );
  NOR U2731 ( .A(n3766), .B(n3650), .Z(n2546) );
  IV U2732 ( .A(n2546), .Z(n2805) );
  XOR U2733 ( .A(n2804), .B(n2805), .Z(n2808) );
  NOR U2734 ( .A(n3635), .B(n3750), .Z(n2751) );
  NOR U2735 ( .A(n3688), .B(n3776), .Z(n2547) );
  IV U2736 ( .A(n2547), .Z(n2750) );
  NOR U2737 ( .A(n3683), .B(n3619), .Z(n2748) );
  XOR U2738 ( .A(n2750), .B(n2748), .Z(n2753) );
  XOR U2739 ( .A(n2751), .B(n2753), .Z(n2807) );
  XOR U2740 ( .A(n2808), .B(n2807), .Z(n2548) );
  IV U2741 ( .A(n2548), .Z(n2735) );
  XOR U2742 ( .A(n2734), .B(n2735), .Z(n2737) );
  XOR U2743 ( .A(n2738), .B(n2737), .Z(n2847) );
  XOR U2744 ( .A(n2845), .B(n2847), .Z(n2848) );
  NOR U2745 ( .A(n2764), .B(n3548), .Z(n3045) );
  IV U2746 ( .A(n3045), .Z(n3187) );
  IV U2747 ( .A(n2549), .Z(n2550) );
  NOR U2748 ( .A(n3187), .B(n2550), .Z(n2554) );
  NOR U2749 ( .A(n2552), .B(n2551), .Z(n2553) );
  NOR U2750 ( .A(n2554), .B(n2553), .Z(n2800) );
  IV U2751 ( .A(o[25]), .Z(n2556) );
  NOR U2752 ( .A(n2556), .B(n2555), .Z(n2714) );
  NOR U2753 ( .A(n3467), .B(n3548), .Z(n2711) );
  NOR U2754 ( .A(n3773), .B(n3634), .Z(n2557) );
  IV U2755 ( .A(n2557), .Z(n2731) );
  XOR U2756 ( .A(n2731), .B(o[26]), .Z(n2713) );
  XOR U2757 ( .A(n2711), .B(n2713), .Z(n2716) );
  XOR U2758 ( .A(n2714), .B(n2716), .Z(n2797) );
  NOR U2759 ( .A(n3779), .B(n2764), .Z(n2559) );
  NOR U2760 ( .A(n3775), .B(n3765), .Z(n2558) );
  XOR U2761 ( .A(n2559), .B(n2558), .Z(n2743) );
  NOR U2762 ( .A(n3462), .B(n3764), .Z(n2560) );
  IV U2763 ( .A(n2560), .Z(n2811) );
  XOR U2764 ( .A(n2811), .B(n2561), .Z(n2813) );
  XOR U2765 ( .A(n2562), .B(n2813), .Z(n2745) );
  XOR U2766 ( .A(n2743), .B(n2745), .Z(n2798) );
  XOR U2767 ( .A(n2797), .B(n2798), .Z(n2563) );
  IV U2768 ( .A(n2563), .Z(n2799) );
  XOR U2769 ( .A(n2800), .B(n2799), .Z(n2849) );
  XOR U2770 ( .A(n2848), .B(n2849), .Z(n2828) );
  IV U2771 ( .A(n2564), .Z(n2566) );
  NOR U2772 ( .A(n2566), .B(n2565), .Z(n2571) );
  IV U2773 ( .A(n2567), .Z(n2568) );
  NOR U2774 ( .A(n2569), .B(n2568), .Z(n2570) );
  NOR U2775 ( .A(n2571), .B(n2570), .Z(n2825) );
  IV U2776 ( .A(n2572), .Z(n2574) );
  NOR U2777 ( .A(n2574), .B(n2573), .Z(n2578) );
  NOR U2778 ( .A(n2576), .B(n2575), .Z(n2577) );
  NOR U2779 ( .A(n2578), .B(n2577), .Z(n2824) );
  XOR U2780 ( .A(n2825), .B(n2824), .Z(n2826) );
  XOR U2781 ( .A(n2828), .B(n2826), .Z(n2698) );
  XOR U2782 ( .A(n2699), .B(n2698), .Z(n2579) );
  IV U2783 ( .A(n2579), .Z(n2701) );
  IV U2784 ( .A(n2580), .Z(n2581) );
  NOR U2785 ( .A(n2582), .B(n2581), .Z(n2587) );
  IV U2786 ( .A(n2583), .Z(n2584) );
  NOR U2787 ( .A(n2585), .B(n2584), .Z(n2586) );
  NOR U2788 ( .A(n2587), .B(n2586), .Z(n2794) );
  NOR U2789 ( .A(n3746), .B(n3621), .Z(n2768) );
  NOR U2790 ( .A(n3489), .B(n3748), .Z(n2588) );
  IV U2791 ( .A(n2588), .Z(n2769) );
  XOR U2792 ( .A(n2768), .B(n2769), .Z(n2771) );
  NOR U2793 ( .A(n3780), .B(n3740), .Z(n2589) );
  IV U2794 ( .A(n2589), .Z(n2778) );
  NOR U2795 ( .A(n3782), .B(n3633), .Z(n2591) );
  NOR U2796 ( .A(n3647), .B(n3686), .Z(n2590) );
  XOR U2797 ( .A(n2591), .B(n2590), .Z(n2777) );
  XOR U2798 ( .A(n2778), .B(n2777), .Z(n2772) );
  XOR U2799 ( .A(n2771), .B(n2772), .Z(n2790) );
  IV U2800 ( .A(y[26]), .Z(n3739) );
  NOR U2801 ( .A(n3680), .B(n3739), .Z(n2723) );
  IV U2802 ( .A(x[26]), .Z(n3745) );
  NOR U2803 ( .A(n3745), .B(n3637), .Z(n2592) );
  IV U2804 ( .A(n2592), .Z(n2722) );
  NOR U2805 ( .A(n3465), .B(n3781), .Z(n2720) );
  XOR U2806 ( .A(n2722), .B(n2720), .Z(n2725) );
  XOR U2807 ( .A(n2723), .B(n2725), .Z(n2820) );
  NOR U2808 ( .A(n3625), .B(n3747), .Z(n2819) );
  IV U2809 ( .A(n2819), .Z(n2817) );
  NOR U2810 ( .A(n3742), .B(n3622), .Z(n2818) );
  IV U2811 ( .A(n2818), .Z(n2816) );
  XOR U2812 ( .A(n2817), .B(n2816), .Z(n2593) );
  XOR U2813 ( .A(n2820), .B(n2593), .Z(n2792) );
  XOR U2814 ( .A(n2790), .B(n2792), .Z(n2793) );
  XOR U2815 ( .A(n2794), .B(n2793), .Z(n2833) );
  NOR U2816 ( .A(n2595), .B(n2594), .Z(n2600) );
  IV U2817 ( .A(n2596), .Z(n2598) );
  NOR U2818 ( .A(n2598), .B(n2597), .Z(n2599) );
  NOR U2819 ( .A(n2600), .B(n2599), .Z(n2831) );
  XOR U2820 ( .A(n2833), .B(n2831), .Z(n2835) );
  NOR U2821 ( .A(n2602), .B(n2601), .Z(n2607) );
  IV U2822 ( .A(n2603), .Z(n2605) );
  NOR U2823 ( .A(n2605), .B(n2604), .Z(n2606) );
  NOR U2824 ( .A(n2607), .B(n2606), .Z(n2608) );
  IV U2825 ( .A(n2608), .Z(n2834) );
  XOR U2826 ( .A(n2835), .B(n2834), .Z(n2842) );
  IV U2827 ( .A(n2609), .Z(n3016) );
  IV U2828 ( .A(n2610), .Z(n2611) );
  NOR U2829 ( .A(n3016), .B(n2611), .Z(n2616) );
  IV U2830 ( .A(n2612), .Z(n2614) );
  NOR U2831 ( .A(n2614), .B(n2613), .Z(n2615) );
  NOR U2832 ( .A(n2616), .B(n2615), .Z(n2839) );
  IV U2833 ( .A(n2617), .Z(n2619) );
  NOR U2834 ( .A(n2619), .B(n2618), .Z(n2623) );
  NOR U2835 ( .A(n2621), .B(n2620), .Z(n2622) );
  NOR U2836 ( .A(n2623), .B(n2622), .Z(n2838) );
  XOR U2837 ( .A(n2839), .B(n2838), .Z(n2840) );
  XOR U2838 ( .A(n2842), .B(n2840), .Z(n2700) );
  XOR U2839 ( .A(n2701), .B(n2700), .Z(n2685) );
  NOR U2840 ( .A(n2625), .B(n2624), .Z(n2629) );
  NOR U2841 ( .A(n2627), .B(n2626), .Z(n2628) );
  NOR U2842 ( .A(n2629), .B(n2628), .Z(n2683) );
  XOR U2843 ( .A(n2685), .B(n2683), .Z(n2688) );
  XOR U2844 ( .A(n2686), .B(n2688), .Z(n2694) );
  XOR U2845 ( .A(n2695), .B(n2694), .Z(n2675) );
  XOR U2846 ( .A(n2677), .B(n2675), .Z(n2680) );
  XOR U2847 ( .A(n2678), .B(n2680), .Z(n2661) );
  IV U2848 ( .A(n2630), .Z(n2631) );
  NOR U2849 ( .A(n2632), .B(n2631), .Z(n2636) );
  NOR U2850 ( .A(n2634), .B(n2633), .Z(n2635) );
  NOR U2851 ( .A(n2636), .B(n2635), .Z(n2672) );
  NOR U2852 ( .A(n2638), .B(n2637), .Z(n2643) );
  IV U2853 ( .A(n2639), .Z(n2640) );
  NOR U2854 ( .A(n2641), .B(n2640), .Z(n2642) );
  NOR U2855 ( .A(n2643), .B(n2642), .Z(n2644) );
  IV U2856 ( .A(n2644), .Z(n2670) );
  NOR U2857 ( .A(n2646), .B(n2645), .Z(n2651) );
  IV U2858 ( .A(n2647), .Z(n2649) );
  NOR U2859 ( .A(n2649), .B(n2648), .Z(n2650) );
  NOR U2860 ( .A(n2651), .B(n2650), .Z(n2668) );
  XOR U2861 ( .A(n2670), .B(n2668), .Z(n2671) );
  XOR U2862 ( .A(n2672), .B(n2671), .Z(n2660) );
  XOR U2863 ( .A(n2661), .B(n2660), .Z(n2665) );
  XOR U2864 ( .A(n2663), .B(n2665), .Z(n2653) );
  XOR U2865 ( .A(n2652), .B(n2653), .Z(n2657) );
  XOR U2866 ( .A(n2655), .B(n2657), .Z(n2855) );
  XOR U2867 ( .A(n2853), .B(n2855), .Z(n2858) );
  XOR U2868 ( .A(n2856), .B(n2858), .Z(N59) );
  NOR U2869 ( .A(n2654), .B(n2653), .Z(n2659) );
  IV U2870 ( .A(n2655), .Z(n2656) );
  NOR U2871 ( .A(n2657), .B(n2656), .Z(n2658) );
  NOR U2872 ( .A(n2659), .B(n2658), .Z(n2862) );
  IV U2873 ( .A(n2660), .Z(n2662) );
  NOR U2874 ( .A(n2662), .B(n2661), .Z(n2667) );
  IV U2875 ( .A(n2663), .Z(n2664) );
  NOR U2876 ( .A(n2665), .B(n2664), .Z(n2666) );
  NOR U2877 ( .A(n2667), .B(n2666), .Z(n2872) );
  IV U2878 ( .A(n2668), .Z(n2669) );
  NOR U2879 ( .A(n2670), .B(n2669), .Z(n2674) );
  NOR U2880 ( .A(n2672), .B(n2671), .Z(n2673) );
  NOR U2881 ( .A(n2674), .B(n2673), .Z(n2869) );
  IV U2882 ( .A(n2675), .Z(n2676) );
  NOR U2883 ( .A(n2677), .B(n2676), .Z(n2682) );
  IV U2884 ( .A(n2678), .Z(n2679) );
  NOR U2885 ( .A(n2680), .B(n2679), .Z(n2681) );
  NOR U2886 ( .A(n2682), .B(n2681), .Z(n2880) );
  IV U2887 ( .A(n2683), .Z(n2684) );
  NOR U2888 ( .A(n2685), .B(n2684), .Z(n2690) );
  IV U2889 ( .A(n2686), .Z(n2687) );
  NOR U2890 ( .A(n2688), .B(n2687), .Z(n2689) );
  NOR U2891 ( .A(n2690), .B(n2689), .Z(n2877) );
  IV U2892 ( .A(n2691), .Z(n2693) );
  NOR U2893 ( .A(n2693), .B(n2692), .Z(n2697) );
  NOR U2894 ( .A(n2695), .B(n2694), .Z(n2696) );
  NOR U2895 ( .A(n2697), .B(n2696), .Z(n2887) );
  NOR U2896 ( .A(n2699), .B(n2698), .Z(n2703) );
  NOR U2897 ( .A(n2701), .B(n2700), .Z(n2702) );
  NOR U2898 ( .A(n2703), .B(n2702), .Z(n2886) );
  IV U2899 ( .A(n2704), .Z(n2706) );
  NOR U2900 ( .A(n2706), .B(n2705), .Z(n2710) );
  NOR U2901 ( .A(n2708), .B(n2707), .Z(n2709) );
  NOR U2902 ( .A(n2710), .B(n2709), .Z(n2989) );
  IV U2903 ( .A(n2711), .Z(n2712) );
  NOR U2904 ( .A(n2713), .B(n2712), .Z(n2718) );
  IV U2905 ( .A(n2714), .Z(n2715) );
  NOR U2906 ( .A(n2716), .B(n2715), .Z(n2717) );
  NOR U2907 ( .A(n2718), .B(n2717), .Z(n2988) );
  XOR U2908 ( .A(n2989), .B(n2988), .Z(n2719) );
  IV U2909 ( .A(n2719), .Z(n2991) );
  IV U2910 ( .A(n2720), .Z(n2721) );
  NOR U2911 ( .A(n2722), .B(n2721), .Z(n2727) );
  IV U2912 ( .A(n2723), .Z(n2724) );
  NOR U2913 ( .A(n2725), .B(n2724), .Z(n2726) );
  NOR U2914 ( .A(n2727), .B(n2726), .Z(n3006) );
  NOR U2915 ( .A(n3646), .B(n3764), .Z(n2943) );
  NOR U2916 ( .A(n3747), .B(n3619), .Z(n2728) );
  IV U2917 ( .A(n2728), .Z(n2944) );
  XOR U2918 ( .A(n2943), .B(n2944), .Z(n2947) );
  NOR U2919 ( .A(n3787), .B(n3686), .Z(n3038) );
  NOR U2920 ( .A(n3625), .B(n3739), .Z(n2729) );
  IV U2921 ( .A(n2729), .Z(n3036) );
  XOR U2922 ( .A(n3036), .B(n2730), .Z(n3040) );
  XOR U2923 ( .A(n3038), .B(n3040), .Z(n2946) );
  XOR U2924 ( .A(n2947), .B(n2946), .Z(n3002) );
  IV U2925 ( .A(o[26]), .Z(n2732) );
  NOR U2926 ( .A(n2732), .B(n2731), .Z(n2981) );
  NOR U2927 ( .A(n3741), .B(n3548), .Z(n2978) );
  NOR U2928 ( .A(n3773), .B(n3745), .Z(n2733) );
  IV U2929 ( .A(n2733), .Z(n3058) );
  XOR U2930 ( .A(n3058), .B(o[27]), .Z(n2979) );
  XOR U2931 ( .A(n2978), .B(n2979), .Z(n2983) );
  XOR U2932 ( .A(n2981), .B(n2983), .Z(n3003) );
  XOR U2933 ( .A(n3002), .B(n3003), .Z(n3005) );
  XOR U2934 ( .A(n3006), .B(n3005), .Z(n2990) );
  XOR U2935 ( .A(n2991), .B(n2990), .Z(n2904) );
  IV U2936 ( .A(n2904), .Z(n2767) );
  IV U2937 ( .A(n2734), .Z(n2736) );
  NOR U2938 ( .A(n2736), .B(n2735), .Z(n2740) );
  NOR U2939 ( .A(n2738), .B(n2737), .Z(n2739) );
  NOR U2940 ( .A(n2740), .B(n2739), .Z(n2902) );
  IV U2941 ( .A(n2741), .Z(n2742) );
  NOR U2942 ( .A(n3009), .B(n2742), .Z(n2747) );
  IV U2943 ( .A(n2743), .Z(n2744) );
  NOR U2944 ( .A(n2745), .B(n2744), .Z(n2746) );
  NOR U2945 ( .A(n2747), .B(n2746), .Z(n2933) );
  IV U2946 ( .A(n2748), .Z(n2749) );
  NOR U2947 ( .A(n2750), .B(n2749), .Z(n2755) );
  IV U2948 ( .A(n2751), .Z(n2752) );
  NOR U2949 ( .A(n2753), .B(n2752), .Z(n2754) );
  NOR U2950 ( .A(n2755), .B(n2754), .Z(n2931) );
  NOR U2951 ( .A(n3628), .B(n3461), .Z(n2757) );
  NOR U2952 ( .A(n3621), .B(n3633), .Z(n2756) );
  XOR U2953 ( .A(n2757), .B(n2756), .Z(n3017) );
  NOR U2954 ( .A(n3650), .B(n3750), .Z(n2953) );
  NOR U2955 ( .A(n3689), .B(n3462), .Z(n2758) );
  IV U2956 ( .A(n2758), .Z(n2952) );
  NOR U2957 ( .A(n3635), .B(n3683), .Z(n2950) );
  XOR U2958 ( .A(n2952), .B(n2950), .Z(n2955) );
  XOR U2959 ( .A(n2953), .B(n2955), .Z(n3019) );
  XOR U2960 ( .A(n3017), .B(n3019), .Z(n2938) );
  NOR U2961 ( .A(n3529), .B(n3622), .Z(n2963) );
  NOR U2962 ( .A(n3647), .B(n3634), .Z(n2759) );
  IV U2963 ( .A(n2759), .Z(n2964) );
  XOR U2964 ( .A(n2963), .B(n2964), .Z(n2966) );
  IV U2965 ( .A(y[27]), .Z(n3649) );
  NOR U2966 ( .A(n3680), .B(n3649), .Z(n3069) );
  NOR U2967 ( .A(n3781), .B(n3742), .Z(n2760) );
  IV U2968 ( .A(n2760), .Z(n3068) );
  IV U2969 ( .A(x[27]), .Z(n3627) );
  NOR U2970 ( .A(n3627), .B(n3637), .Z(n3066) );
  XOR U2971 ( .A(n3068), .B(n3066), .Z(n3071) );
  XOR U2972 ( .A(n3069), .B(n3071), .Z(n2967) );
  XOR U2973 ( .A(n2966), .B(n2967), .Z(n2936) );
  XOR U2974 ( .A(n2938), .B(n2936), .Z(n2939) );
  NOR U2975 ( .A(n3766), .B(n3740), .Z(n2970) );
  NOR U2976 ( .A(n3687), .B(n3782), .Z(n2761) );
  IV U2977 ( .A(n2761), .Z(n2971) );
  XOR U2978 ( .A(n2970), .B(n2971), .Z(n2975) );
  NOR U2979 ( .A(n3748), .B(n3780), .Z(n2973) );
  XOR U2980 ( .A(n2975), .B(n2973), .Z(n3032) );
  NOR U2981 ( .A(n3645), .B(n3746), .Z(n3028) );
  NOR U2982 ( .A(n3763), .B(n3776), .Z(n2762) );
  IV U2983 ( .A(n2762), .Z(n3029) );
  XOR U2984 ( .A(n3028), .B(n3029), .Z(n3031) );
  XOR U2985 ( .A(n3032), .B(n3031), .Z(n3011) );
  NOR U2986 ( .A(n3549), .B(n3765), .Z(n3208) );
  NOR U2987 ( .A(n3161), .B(n3749), .Z(n2763) );
  XOR U2988 ( .A(n3208), .B(n2763), .Z(n3023) );
  NOR U2989 ( .A(n3062), .B(n2764), .Z(n3052) );
  NOR U2990 ( .A(n3682), .B(n3489), .Z(n2765) );
  IV U2991 ( .A(n2765), .Z(n3051) );
  NOR U2992 ( .A(n3465), .B(n3688), .Z(n3049) );
  XOR U2993 ( .A(n3051), .B(n3049), .Z(n3054) );
  XOR U2994 ( .A(n3052), .B(n3054), .Z(n3025) );
  XOR U2995 ( .A(n3023), .B(n3025), .Z(n3010) );
  XOR U2996 ( .A(n2766), .B(n3010), .Z(n3012) );
  XOR U2997 ( .A(n3011), .B(n3012), .Z(n2940) );
  XOR U2998 ( .A(n2939), .B(n2940), .Z(n2929) );
  XOR U2999 ( .A(n2931), .B(n2929), .Z(n2932) );
  XOR U3000 ( .A(n2933), .B(n2932), .Z(n2900) );
  XOR U3001 ( .A(n2902), .B(n2900), .Z(n2903) );
  XOR U3002 ( .A(n2767), .B(n2903), .Z(n2910) );
  IV U3003 ( .A(n2768), .Z(n2770) );
  NOR U3004 ( .A(n2770), .B(n2769), .Z(n2774) );
  NOR U3005 ( .A(n2772), .B(n2771), .Z(n2773) );
  NOR U3006 ( .A(n2774), .B(n2773), .Z(n2999) );
  NOR U3007 ( .A(n3633), .B(n3686), .Z(n3544) );
  IV U3008 ( .A(n3544), .Z(n3670) );
  IV U3009 ( .A(n2775), .Z(n2776) );
  NOR U3010 ( .A(n3670), .B(n2776), .Z(n2781) );
  IV U3011 ( .A(n2777), .Z(n2779) );
  NOR U3012 ( .A(n2779), .B(n2778), .Z(n2780) );
  NOR U3013 ( .A(n2781), .B(n2780), .Z(n2997) );
  NOR U3014 ( .A(n2783), .B(n2782), .Z(n2789) );
  NOR U3015 ( .A(n2785), .B(n2784), .Z(n2786) );
  NOR U3016 ( .A(n2787), .B(n2786), .Z(n2788) );
  NOR U3017 ( .A(n2789), .B(n2788), .Z(n2995) );
  XOR U3018 ( .A(n2997), .B(n2995), .Z(n2998) );
  XOR U3019 ( .A(n2999), .B(n2998), .Z(n2917) );
  IV U3020 ( .A(n2790), .Z(n2791) );
  NOR U3021 ( .A(n2792), .B(n2791), .Z(n2796) );
  NOR U3022 ( .A(n2794), .B(n2793), .Z(n2795) );
  NOR U3023 ( .A(n2796), .B(n2795), .Z(n2915) );
  XOR U3024 ( .A(n2917), .B(n2915), .Z(n2919) );
  NOR U3025 ( .A(n2798), .B(n2797), .Z(n2802) );
  NOR U3026 ( .A(n2800), .B(n2799), .Z(n2801) );
  NOR U3027 ( .A(n2802), .B(n2801), .Z(n2803) );
  IV U3028 ( .A(n2803), .Z(n2918) );
  XOR U3029 ( .A(n2919), .B(n2918), .Z(n2908) );
  IV U3030 ( .A(n2804), .Z(n2806) );
  NOR U3031 ( .A(n2806), .B(n2805), .Z(n2810) );
  NOR U3032 ( .A(n2808), .B(n2807), .Z(n2809) );
  NOR U3033 ( .A(n2810), .B(n2809), .Z(n2926) );
  NOR U3034 ( .A(n3022), .B(n2811), .Z(n2815) );
  NOR U3035 ( .A(n2813), .B(n2812), .Z(n2814) );
  NOR U3036 ( .A(n2815), .B(n2814), .Z(n2923) );
  NOR U3037 ( .A(n2817), .B(n2816), .Z(n2823) );
  NOR U3038 ( .A(n2819), .B(n2818), .Z(n2821) );
  NOR U3039 ( .A(n2821), .B(n2820), .Z(n2822) );
  NOR U3040 ( .A(n2823), .B(n2822), .Z(n2922) );
  XOR U3041 ( .A(n2923), .B(n2922), .Z(n2924) );
  XOR U3042 ( .A(n2926), .B(n2924), .Z(n2907) );
  XOR U3043 ( .A(n2908), .B(n2907), .Z(n2909) );
  XOR U3044 ( .A(n2910), .B(n2909), .Z(n3078) );
  NOR U3045 ( .A(n2825), .B(n2824), .Z(n2830) );
  IV U3046 ( .A(n2826), .Z(n2827) );
  NOR U3047 ( .A(n2828), .B(n2827), .Z(n2829) );
  NOR U3048 ( .A(n2830), .B(n2829), .Z(n3077) );
  IV U3049 ( .A(n2831), .Z(n2832) );
  NOR U3050 ( .A(n2833), .B(n2832), .Z(n2837) );
  NOR U3051 ( .A(n2835), .B(n2834), .Z(n2836) );
  NOR U3052 ( .A(n2837), .B(n2836), .Z(n3075) );
  XOR U3053 ( .A(n3077), .B(n3075), .Z(n3079) );
  XOR U3054 ( .A(n3078), .B(n3079), .Z(n2895) );
  NOR U3055 ( .A(n2839), .B(n2838), .Z(n2844) );
  IV U3056 ( .A(n2840), .Z(n2841) );
  NOR U3057 ( .A(n2842), .B(n2841), .Z(n2843) );
  NOR U3058 ( .A(n2844), .B(n2843), .Z(n2894) );
  IV U3059 ( .A(n2845), .Z(n2846) );
  NOR U3060 ( .A(n2847), .B(n2846), .Z(n2851) );
  NOR U3061 ( .A(n2849), .B(n2848), .Z(n2850) );
  NOR U3062 ( .A(n2851), .B(n2850), .Z(n2892) );
  XOR U3063 ( .A(n2894), .B(n2892), .Z(n2896) );
  XOR U3064 ( .A(n2895), .B(n2896), .Z(n2885) );
  XOR U3065 ( .A(n2886), .B(n2885), .Z(n2852) );
  IV U3066 ( .A(n2852), .Z(n2889) );
  XOR U3067 ( .A(n2887), .B(n2889), .Z(n2878) );
  XOR U3068 ( .A(n2877), .B(n2878), .Z(n2881) );
  XOR U3069 ( .A(n2880), .B(n2881), .Z(n2871) );
  XOR U3070 ( .A(n2869), .B(n2871), .Z(n2873) );
  XOR U3071 ( .A(n2872), .B(n2873), .Z(n2864) );
  XOR U3072 ( .A(n2862), .B(n2864), .Z(n2866) );
  IV U3073 ( .A(n2853), .Z(n2854) );
  NOR U3074 ( .A(n2855), .B(n2854), .Z(n2860) );
  IV U3075 ( .A(n2856), .Z(n2857) );
  NOR U3076 ( .A(n2858), .B(n2857), .Z(n2859) );
  NOR U3077 ( .A(n2860), .B(n2859), .Z(n2861) );
  IV U3078 ( .A(n2861), .Z(n2865) );
  XOR U3079 ( .A(n2866), .B(n2865), .Z(N60) );
  IV U3080 ( .A(n2862), .Z(n2863) );
  NOR U3081 ( .A(n2864), .B(n2863), .Z(n2868) );
  NOR U3082 ( .A(n2866), .B(n2865), .Z(n2867) );
  NOR U3083 ( .A(n2868), .B(n2867), .Z(n3307) );
  IV U3084 ( .A(n2869), .Z(n2870) );
  NOR U3085 ( .A(n2871), .B(n2870), .Z(n2876) );
  IV U3086 ( .A(n2872), .Z(n2874) );
  NOR U3087 ( .A(n2874), .B(n2873), .Z(n2875) );
  NOR U3088 ( .A(n2876), .B(n2875), .Z(n3304) );
  IV U3089 ( .A(n2877), .Z(n2879) );
  NOR U3090 ( .A(n2879), .B(n2878), .Z(n2884) );
  IV U3091 ( .A(n2880), .Z(n2882) );
  NOR U3092 ( .A(n2882), .B(n2881), .Z(n2883) );
  NOR U3093 ( .A(n2884), .B(n2883), .Z(n3085) );
  NOR U3094 ( .A(n2886), .B(n2885), .Z(n2891) );
  IV U3095 ( .A(n2887), .Z(n2888) );
  NOR U3096 ( .A(n2889), .B(n2888), .Z(n2890) );
  NOR U3097 ( .A(n2891), .B(n2890), .Z(n3082) );
  IV U3098 ( .A(n2892), .Z(n2893) );
  NOR U3099 ( .A(n2894), .B(n2893), .Z(n2899) );
  IV U3100 ( .A(n2895), .Z(n2897) );
  NOR U3101 ( .A(n2897), .B(n2896), .Z(n2898) );
  NOR U3102 ( .A(n2899), .B(n2898), .Z(n3093) );
  IV U3103 ( .A(n2900), .Z(n2901) );
  NOR U3104 ( .A(n2902), .B(n2901), .Z(n2906) );
  NOR U3105 ( .A(n2904), .B(n2903), .Z(n2905) );
  NOR U3106 ( .A(n2906), .B(n2905), .Z(n3099) );
  NOR U3107 ( .A(n2908), .B(n2907), .Z(n2913) );
  IV U3108 ( .A(n2909), .Z(n2911) );
  NOR U3109 ( .A(n2911), .B(n2910), .Z(n2912) );
  NOR U3110 ( .A(n2913), .B(n2912), .Z(n3098) );
  XOR U3111 ( .A(n3099), .B(n3098), .Z(n2914) );
  IV U3112 ( .A(n2914), .Z(n3100) );
  IV U3113 ( .A(n2915), .Z(n2916) );
  NOR U3114 ( .A(n2917), .B(n2916), .Z(n2921) );
  NOR U3115 ( .A(n2919), .B(n2918), .Z(n2920) );
  NOR U3116 ( .A(n2921), .B(n2920), .Z(n3108) );
  NOR U3117 ( .A(n2923), .B(n2922), .Z(n2928) );
  IV U3118 ( .A(n2924), .Z(n2925) );
  NOR U3119 ( .A(n2926), .B(n2925), .Z(n2927) );
  NOR U3120 ( .A(n2928), .B(n2927), .Z(n3104) );
  IV U3121 ( .A(n2929), .Z(n2930) );
  NOR U3122 ( .A(n2931), .B(n2930), .Z(n2935) );
  NOR U3123 ( .A(n2933), .B(n2932), .Z(n2934) );
  NOR U3124 ( .A(n2935), .B(n2934), .Z(n3114) );
  IV U3125 ( .A(n2936), .Z(n2937) );
  NOR U3126 ( .A(n2938), .B(n2937), .Z(n2942) );
  NOR U3127 ( .A(n2940), .B(n2939), .Z(n2941) );
  NOR U3128 ( .A(n2942), .B(n2941), .Z(n3112) );
  IV U3129 ( .A(n3112), .Z(n2987) );
  IV U3130 ( .A(n2943), .Z(n2945) );
  NOR U3131 ( .A(n2945), .B(n2944), .Z(n2949) );
  NOR U3132 ( .A(n2947), .B(n2946), .Z(n2948) );
  NOR U3133 ( .A(n2949), .B(n2948), .Z(n3237) );
  IV U3134 ( .A(n2950), .Z(n2951) );
  NOR U3135 ( .A(n2952), .B(n2951), .Z(n2957) );
  IV U3136 ( .A(n2953), .Z(n2954) );
  NOR U3137 ( .A(n2955), .B(n2954), .Z(n2956) );
  NOR U3138 ( .A(n2957), .B(n2956), .Z(n3277) );
  NOR U3139 ( .A(n3688), .B(n3742), .Z(n3171) );
  IV U3140 ( .A(y[28]), .Z(n3636) );
  NOR U3141 ( .A(n3680), .B(n3636), .Z(n2958) );
  IV U3142 ( .A(n2958), .Z(n3172) );
  XOR U3143 ( .A(n3171), .B(n3172), .Z(n3176) );
  NOR U3144 ( .A(n3649), .B(n3625), .Z(n3174) );
  XOR U3145 ( .A(n3176), .B(n3174), .Z(n3269) );
  NOR U3146 ( .A(n3739), .B(n3619), .Z(n3265) );
  NOR U3147 ( .A(n3622), .B(n3764), .Z(n2959) );
  IV U3148 ( .A(n2959), .Z(n3266) );
  XOR U3149 ( .A(n3265), .B(n3266), .Z(n3268) );
  XOR U3150 ( .A(n3269), .B(n3268), .Z(n3273) );
  NOR U3151 ( .A(n3750), .B(n3740), .Z(n2960) );
  IV U3152 ( .A(n2960), .Z(n3180) );
  XOR U3153 ( .A(n2961), .B(n3180), .Z(n3183) );
  NOR U3154 ( .A(n3787), .B(n3634), .Z(n3192) );
  XOR U3155 ( .A(n3192), .B(n3193), .Z(n3197) );
  NOR U3156 ( .A(n3683), .B(n3650), .Z(n3195) );
  XOR U3157 ( .A(n3197), .B(n3195), .Z(n3182) );
  XOR U3158 ( .A(n3183), .B(n3182), .Z(n2962) );
  IV U3159 ( .A(n2962), .Z(n3274) );
  XOR U3160 ( .A(n3273), .B(n3274), .Z(n3276) );
  XOR U3161 ( .A(n3277), .B(n3276), .Z(n3239) );
  XOR U3162 ( .A(n3237), .B(n3239), .Z(n3240) );
  IV U3163 ( .A(n2963), .Z(n2965) );
  NOR U3164 ( .A(n2965), .B(n2964), .Z(n2969) );
  NOR U3165 ( .A(n2967), .B(n2966), .Z(n2968) );
  NOR U3166 ( .A(n2969), .B(n2968), .Z(n3284) );
  IV U3167 ( .A(n2970), .Z(n2972) );
  NOR U3168 ( .A(n2972), .B(n2971), .Z(n2977) );
  IV U3169 ( .A(n2973), .Z(n2974) );
  NOR U3170 ( .A(n2975), .B(n2974), .Z(n2976) );
  NOR U3171 ( .A(n2977), .B(n2976), .Z(n3282) );
  IV U3172 ( .A(n2978), .Z(n2980) );
  NOR U3173 ( .A(n2980), .B(n2979), .Z(n2985) );
  IV U3174 ( .A(n2981), .Z(n2982) );
  NOR U3175 ( .A(n2983), .B(n2982), .Z(n2984) );
  NOR U3176 ( .A(n2985), .B(n2984), .Z(n3281) );
  XOR U3177 ( .A(n3282), .B(n3281), .Z(n2986) );
  IV U3178 ( .A(n2986), .Z(n3283) );
  XOR U3179 ( .A(n3284), .B(n3283), .Z(n3241) );
  XOR U3180 ( .A(n3240), .B(n3241), .Z(n3111) );
  XOR U3181 ( .A(n2987), .B(n3111), .Z(n3113) );
  XOR U3182 ( .A(n3114), .B(n3113), .Z(n3121) );
  NOR U3183 ( .A(n2989), .B(n2988), .Z(n2994) );
  IV U3184 ( .A(n2990), .Z(n2992) );
  NOR U3185 ( .A(n2992), .B(n2991), .Z(n2993) );
  NOR U3186 ( .A(n2994), .B(n2993), .Z(n3117) );
  IV U3187 ( .A(n2995), .Z(n2996) );
  NOR U3188 ( .A(n2997), .B(n2996), .Z(n3001) );
  NOR U3189 ( .A(n2999), .B(n2998), .Z(n3000) );
  NOR U3190 ( .A(n3001), .B(n3000), .Z(n3127) );
  IV U3191 ( .A(n3002), .Z(n3004) );
  NOR U3192 ( .A(n3004), .B(n3003), .Z(n3008) );
  NOR U3193 ( .A(n3006), .B(n3005), .Z(n3007) );
  NOR U3194 ( .A(n3008), .B(n3007), .Z(n3124) );
  NOR U3195 ( .A(n3010), .B(n3009), .Z(n3015) );
  IV U3196 ( .A(n3011), .Z(n3013) );
  NOR U3197 ( .A(n3013), .B(n3012), .Z(n3014) );
  NOR U3198 ( .A(n3015), .B(n3014), .Z(n3299) );
  NOR U3199 ( .A(n3633), .B(n3461), .Z(n3232) );
  IV U3200 ( .A(n3232), .Z(n3484) );
  NOR U3201 ( .A(n3016), .B(n3484), .Z(n3021) );
  IV U3202 ( .A(n3017), .Z(n3018) );
  NOR U3203 ( .A(n3019), .B(n3018), .Z(n3020) );
  NOR U3204 ( .A(n3021), .B(n3020), .Z(n3296) );
  NOR U3205 ( .A(n3490), .B(n3022), .Z(n3027) );
  IV U3206 ( .A(n3023), .Z(n3024) );
  NOR U3207 ( .A(n3025), .B(n3024), .Z(n3026) );
  NOR U3208 ( .A(n3027), .B(n3026), .Z(n3295) );
  XOR U3209 ( .A(n3296), .B(n3295), .Z(n3297) );
  XOR U3210 ( .A(n3299), .B(n3297), .Z(n3135) );
  IV U3211 ( .A(n3028), .Z(n3030) );
  NOR U3212 ( .A(n3030), .B(n3029), .Z(n3034) );
  NOR U3213 ( .A(n3032), .B(n3031), .Z(n3033) );
  NOR U3214 ( .A(n3034), .B(n3033), .Z(n3035) );
  IV U3215 ( .A(n3035), .Z(n3134) );
  NOR U3216 ( .A(n3037), .B(n3036), .Z(n3042) );
  IV U3217 ( .A(n3038), .Z(n3039) );
  NOR U3218 ( .A(n3040), .B(n3039), .Z(n3041) );
  NOR U3219 ( .A(n3042), .B(n3041), .Z(n3144) );
  NOR U3220 ( .A(n3461), .B(n3746), .Z(n3216) );
  NOR U3221 ( .A(n3766), .B(n3748), .Z(n3043) );
  IV U3222 ( .A(n3043), .Z(n3454) );
  XOR U3223 ( .A(n3216), .B(n3454), .Z(n3220) );
  NOR U3224 ( .A(n3686), .B(n3628), .Z(n3218) );
  XOR U3225 ( .A(n3220), .B(n3218), .Z(n3189) );
  NOR U3226 ( .A(n3682), .B(n3780), .Z(n3044) );
  IV U3227 ( .A(n3044), .Z(n3186) );
  XOR U3228 ( .A(n3045), .B(n3186), .Z(n3188) );
  XOR U3229 ( .A(n3189), .B(n3188), .Z(n3140) );
  IV U3230 ( .A(x[28]), .Z(n3788) );
  NOR U3231 ( .A(n3637), .B(n3788), .Z(n3257) );
  NOR U3232 ( .A(n3465), .B(n3763), .Z(n3046) );
  IV U3233 ( .A(n3046), .Z(n3258) );
  XOR U3234 ( .A(n3257), .B(n3258), .Z(n3262) );
  NOR U3235 ( .A(n3745), .B(n3647), .Z(n3260) );
  XOR U3236 ( .A(n3262), .B(n3260), .Z(n3254) );
  NOR U3237 ( .A(n3747), .B(n3635), .Z(n3250) );
  NOR U3238 ( .A(n3467), .B(n3776), .Z(n3047) );
  IV U3239 ( .A(n3047), .Z(n3251) );
  XOR U3240 ( .A(n3250), .B(n3251), .Z(n3253) );
  XOR U3241 ( .A(n3254), .B(n3253), .Z(n3048) );
  IV U3242 ( .A(n3048), .Z(n3141) );
  XOR U3243 ( .A(n3140), .B(n3141), .Z(n3143) );
  XOR U3244 ( .A(n3144), .B(n3143), .Z(n3292) );
  IV U3245 ( .A(n3049), .Z(n3050) );
  NOR U3246 ( .A(n3051), .B(n3050), .Z(n3056) );
  IV U3247 ( .A(n3052), .Z(n3053) );
  NOR U3248 ( .A(n3054), .B(n3053), .Z(n3055) );
  NOR U3249 ( .A(n3056), .B(n3055), .Z(n3247) );
  NOR U3250 ( .A(n3773), .B(n3627), .Z(n3149) );
  IV U3251 ( .A(o[28]), .Z(n3150) );
  XOR U3252 ( .A(n3149), .B(n3150), .Z(n3165) );
  NOR U3253 ( .A(n3741), .B(n3546), .Z(n3163) );
  XOR U3254 ( .A(n3165), .B(n3163), .Z(n3168) );
  IV U3255 ( .A(o[27]), .Z(n3057) );
  NOR U3256 ( .A(n3058), .B(n3057), .Z(n3166) );
  XOR U3257 ( .A(n3168), .B(n3166), .Z(n3244) );
  NOR U3258 ( .A(n3549), .B(n3779), .Z(n3059) );
  IV U3259 ( .A(n3059), .Z(n3061) );
  XOR U3260 ( .A(n3061), .B(n3060), .Z(n3212) );
  NOR U3261 ( .A(n3781), .B(n3529), .Z(n3200) );
  NOR U3262 ( .A(n3062), .B(n3775), .Z(n3063) );
  IV U3263 ( .A(n3063), .Z(n3201) );
  XOR U3264 ( .A(n3200), .B(n3201), .Z(n3203) );
  NOR U3265 ( .A(n3689), .B(n3646), .Z(n3226) );
  NOR U3266 ( .A(n3489), .B(n3749), .Z(n3064) );
  IV U3267 ( .A(n3064), .Z(n3225) );
  NOR U3268 ( .A(n3645), .B(n3633), .Z(n3223) );
  XOR U3269 ( .A(n3225), .B(n3223), .Z(n3228) );
  XOR U3270 ( .A(n3226), .B(n3228), .Z(n3204) );
  XOR U3271 ( .A(n3203), .B(n3204), .Z(n3211) );
  XOR U3272 ( .A(n3212), .B(n3211), .Z(n3245) );
  XOR U3273 ( .A(n3244), .B(n3245), .Z(n3065) );
  IV U3274 ( .A(n3065), .Z(n3246) );
  XOR U3275 ( .A(n3247), .B(n3246), .Z(n3290) );
  IV U3276 ( .A(n3066), .Z(n3067) );
  NOR U3277 ( .A(n3068), .B(n3067), .Z(n3073) );
  IV U3278 ( .A(n3069), .Z(n3070) );
  NOR U3279 ( .A(n3071), .B(n3070), .Z(n3072) );
  NOR U3280 ( .A(n3073), .B(n3072), .Z(n3288) );
  XOR U3281 ( .A(n3290), .B(n3288), .Z(n3291) );
  XOR U3282 ( .A(n3292), .B(n3291), .Z(n3132) );
  XOR U3283 ( .A(n3134), .B(n3132), .Z(n3136) );
  XOR U3284 ( .A(n3135), .B(n3136), .Z(n3126) );
  XOR U3285 ( .A(n3124), .B(n3126), .Z(n3129) );
  XOR U3286 ( .A(n3127), .B(n3129), .Z(n3119) );
  XOR U3287 ( .A(n3117), .B(n3119), .Z(n3120) );
  XOR U3288 ( .A(n3121), .B(n3120), .Z(n3074) );
  IV U3289 ( .A(n3074), .Z(n3106) );
  XOR U3290 ( .A(n3104), .B(n3106), .Z(n3107) );
  XOR U3291 ( .A(n3108), .B(n3107), .Z(n3101) );
  XOR U3292 ( .A(n3100), .B(n3101), .Z(n3092) );
  IV U3293 ( .A(n3075), .Z(n3076) );
  NOR U3294 ( .A(n3077), .B(n3076), .Z(n3081) );
  NOR U3295 ( .A(n3079), .B(n3078), .Z(n3080) );
  NOR U3296 ( .A(n3081), .B(n3080), .Z(n3090) );
  XOR U3297 ( .A(n3092), .B(n3090), .Z(n3095) );
  XOR U3298 ( .A(n3093), .B(n3095), .Z(n3084) );
  XOR U3299 ( .A(n3082), .B(n3084), .Z(n3087) );
  XOR U3300 ( .A(n3085), .B(n3087), .Z(n3306) );
  XOR U3301 ( .A(n3304), .B(n3306), .Z(n3309) );
  XOR U3302 ( .A(n3307), .B(n3309), .Z(N61) );
  IV U3303 ( .A(n3082), .Z(n3083) );
  NOR U3304 ( .A(n3084), .B(n3083), .Z(n3089) );
  IV U3305 ( .A(n3085), .Z(n3086) );
  NOR U3306 ( .A(n3087), .B(n3086), .Z(n3088) );
  NOR U3307 ( .A(n3089), .B(n3088), .Z(n3313) );
  IV U3308 ( .A(n3090), .Z(n3091) );
  NOR U3309 ( .A(n3092), .B(n3091), .Z(n3097) );
  IV U3310 ( .A(n3093), .Z(n3094) );
  NOR U3311 ( .A(n3095), .B(n3094), .Z(n3096) );
  NOR U3312 ( .A(n3097), .B(n3096), .Z(n3322) );
  NOR U3313 ( .A(n3099), .B(n3098), .Z(n3103) );
  NOR U3314 ( .A(n3101), .B(n3100), .Z(n3102) );
  NOR U3315 ( .A(n3103), .B(n3102), .Z(n3321) );
  IV U3316 ( .A(n3321), .Z(n3303) );
  IV U3317 ( .A(n3104), .Z(n3105) );
  NOR U3318 ( .A(n3106), .B(n3105), .Z(n3110) );
  NOR U3319 ( .A(n3108), .B(n3107), .Z(n3109) );
  NOR U3320 ( .A(n3110), .B(n3109), .Z(n3329) );
  NOR U3321 ( .A(n3112), .B(n3111), .Z(n3116) );
  NOR U3322 ( .A(n3114), .B(n3113), .Z(n3115) );
  NOR U3323 ( .A(n3116), .B(n3115), .Z(n3328) );
  IV U3324 ( .A(n3328), .Z(n3302) );
  IV U3325 ( .A(n3117), .Z(n3118) );
  NOR U3326 ( .A(n3119), .B(n3118), .Z(n3123) );
  NOR U3327 ( .A(n3121), .B(n3120), .Z(n3122) );
  NOR U3328 ( .A(n3123), .B(n3122), .Z(n3337) );
  IV U3329 ( .A(n3124), .Z(n3125) );
  NOR U3330 ( .A(n3126), .B(n3125), .Z(n3131) );
  IV U3331 ( .A(n3127), .Z(n3128) );
  NOR U3332 ( .A(n3129), .B(n3128), .Z(n3130) );
  NOR U3333 ( .A(n3131), .B(n3130), .Z(n3334) );
  IV U3334 ( .A(n3132), .Z(n3133) );
  NOR U3335 ( .A(n3134), .B(n3133), .Z(n3139) );
  IV U3336 ( .A(n3135), .Z(n3137) );
  NOR U3337 ( .A(n3137), .B(n3136), .Z(n3138) );
  NOR U3338 ( .A(n3139), .B(n3138), .Z(n3360) );
  IV U3339 ( .A(n3140), .Z(n3142) );
  NOR U3340 ( .A(n3142), .B(n3141), .Z(n3146) );
  NOR U3341 ( .A(n3144), .B(n3143), .Z(n3145) );
  NOR U3342 ( .A(n3146), .B(n3145), .Z(n3410) );
  IV U3343 ( .A(x[29]), .Z(n3648) );
  NOR U3344 ( .A(n3637), .B(n3648), .Z(n3512) );
  NOR U3345 ( .A(n3465), .B(n3467), .Z(n3147) );
  IV U3346 ( .A(n3147), .Z(n3513) );
  XOR U3347 ( .A(n3512), .B(n3513), .Z(n3517) );
  IV U3348 ( .A(y[29]), .Z(n3620) );
  NOR U3349 ( .A(n3680), .B(n3620), .Z(n3515) );
  XOR U3350 ( .A(n3517), .B(n3515), .Z(n3508) );
  NOR U3351 ( .A(n3627), .B(n3647), .Z(n3504) );
  NOR U3352 ( .A(n3781), .B(n3764), .Z(n3148) );
  IV U3353 ( .A(n3148), .Z(n3505) );
  XOR U3354 ( .A(n3504), .B(n3505), .Z(n3507) );
  XOR U3355 ( .A(n3508), .B(n3507), .Z(n3478) );
  IV U3356 ( .A(n3149), .Z(n3151) );
  NOR U3357 ( .A(n3151), .B(n3150), .Z(n3152) );
  IV U3358 ( .A(n3152), .Z(n3472) );
  NOR U3359 ( .A(n3773), .B(n3788), .Z(n3153) );
  IV U3360 ( .A(n3153), .Z(n3532) );
  XOR U3361 ( .A(o[29]), .B(n3532), .Z(n3469) );
  XOR U3362 ( .A(n3154), .B(n3469), .Z(n3471) );
  XOR U3363 ( .A(n3472), .B(n3471), .Z(n3475) );
  NOR U3364 ( .A(n3750), .B(n3748), .Z(n3156) );
  NOR U3365 ( .A(n3766), .B(n3682), .Z(n3155) );
  XOR U3366 ( .A(n3156), .B(n3155), .Z(n3455) );
  NOR U3367 ( .A(n3749), .B(n3780), .Z(n3157) );
  IV U3368 ( .A(n3157), .Z(n3456) );
  XOR U3369 ( .A(n3455), .B(n3456), .Z(n3476) );
  XOR U3370 ( .A(n3475), .B(n3476), .Z(n3479) );
  XOR U3371 ( .A(n3478), .B(n3479), .Z(n3397) );
  NOR U3372 ( .A(n3628), .B(n3634), .Z(n3437) );
  NOR U3373 ( .A(n3645), .B(n3687), .Z(n3158) );
  IV U3374 ( .A(n3158), .Z(n3438) );
  XOR U3375 ( .A(n3437), .B(n3438), .Z(n3441) );
  NOR U3376 ( .A(n3739), .B(n3635), .Z(n3496) );
  XOR U3377 ( .A(n3496), .B(n3497), .Z(n3501) );
  NOR U3378 ( .A(n3747), .B(n3650), .Z(n3499) );
  XOR U3379 ( .A(n3501), .B(n3499), .Z(n3440) );
  XOR U3380 ( .A(n3441), .B(n3440), .Z(n3393) );
  NOR U3381 ( .A(n3689), .B(n3622), .Z(n3520) );
  NOR U3382 ( .A(n3775), .B(n3548), .Z(n3159) );
  IV U3383 ( .A(n3159), .Z(n3521) );
  XOR U3384 ( .A(n3520), .B(n3521), .Z(n3524) );
  XOR U3385 ( .A(n3524), .B(n3160), .Z(n3493) );
  NOR U3386 ( .A(n3161), .B(n3779), .Z(n3207) );
  XOR U3387 ( .A(n3207), .B(n3162), .Z(n3491) );
  XOR U3388 ( .A(n3493), .B(n3491), .Z(n3394) );
  XOR U3389 ( .A(n3393), .B(n3394), .Z(n3396) );
  XOR U3390 ( .A(n3397), .B(n3396), .Z(n3374) );
  IV U3391 ( .A(n3163), .Z(n3164) );
  NOR U3392 ( .A(n3165), .B(n3164), .Z(n3170) );
  IV U3393 ( .A(n3166), .Z(n3167) );
  NOR U3394 ( .A(n3168), .B(n3167), .Z(n3169) );
  NOR U3395 ( .A(n3170), .B(n3169), .Z(n3373) );
  IV U3396 ( .A(n3171), .Z(n3173) );
  NOR U3397 ( .A(n3173), .B(n3172), .Z(n3178) );
  IV U3398 ( .A(n3174), .Z(n3175) );
  NOR U3399 ( .A(n3176), .B(n3175), .Z(n3177) );
  NOR U3400 ( .A(n3178), .B(n3177), .Z(n3372) );
  XOR U3401 ( .A(n3373), .B(n3372), .Z(n3179) );
  IV U3402 ( .A(n3179), .Z(n3375) );
  XOR U3403 ( .A(n3374), .B(n3375), .Z(n3409) );
  XOR U3404 ( .A(n3410), .B(n3409), .Z(n3411) );
  NOR U3405 ( .A(n3181), .B(n3180), .Z(n3185) );
  NOR U3406 ( .A(n3183), .B(n3182), .Z(n3184) );
  NOR U3407 ( .A(n3185), .B(n3184), .Z(n3366) );
  NOR U3408 ( .A(n3187), .B(n3186), .Z(n3191) );
  NOR U3409 ( .A(n3189), .B(n3188), .Z(n3190) );
  NOR U3410 ( .A(n3191), .B(n3190), .Z(n3427) );
  IV U3411 ( .A(n3192), .Z(n3194) );
  NOR U3412 ( .A(n3194), .B(n3193), .Z(n3199) );
  IV U3413 ( .A(n3195), .Z(n3196) );
  NOR U3414 ( .A(n3197), .B(n3196), .Z(n3198) );
  NOR U3415 ( .A(n3199), .B(n3198), .Z(n3424) );
  IV U3416 ( .A(n3200), .Z(n3202) );
  NOR U3417 ( .A(n3202), .B(n3201), .Z(n3206) );
  NOR U3418 ( .A(n3204), .B(n3203), .Z(n3205) );
  NOR U3419 ( .A(n3206), .B(n3205), .Z(n3423) );
  XOR U3420 ( .A(n3424), .B(n3423), .Z(n3425) );
  XOR U3421 ( .A(n3427), .B(n3425), .Z(n3365) );
  XOR U3422 ( .A(n3366), .B(n3365), .Z(n3367) );
  IV U3423 ( .A(n3207), .Z(n3210) );
  IV U3424 ( .A(n3208), .Z(n3209) );
  NOR U3425 ( .A(n3210), .B(n3209), .Z(n3215) );
  IV U3426 ( .A(n3211), .Z(n3213) );
  NOR U3427 ( .A(n3213), .B(n3212), .Z(n3214) );
  NOR U3428 ( .A(n3215), .B(n3214), .Z(n3383) );
  IV U3429 ( .A(n3216), .Z(n3217) );
  NOR U3430 ( .A(n3217), .B(n3454), .Z(n3222) );
  IV U3431 ( .A(n3218), .Z(n3219) );
  NOR U3432 ( .A(n3220), .B(n3219), .Z(n3221) );
  NOR U3433 ( .A(n3222), .B(n3221), .Z(n3381) );
  IV U3434 ( .A(n3223), .Z(n3224) );
  NOR U3435 ( .A(n3225), .B(n3224), .Z(n3230) );
  IV U3436 ( .A(n3226), .Z(n3227) );
  NOR U3437 ( .A(n3228), .B(n3227), .Z(n3229) );
  NOR U3438 ( .A(n3230), .B(n3229), .Z(n3390) );
  NOR U3439 ( .A(n3683), .B(n3740), .Z(n3445) );
  NOR U3440 ( .A(n3621), .B(n3462), .Z(n3231) );
  IV U3441 ( .A(n3231), .Z(n3446) );
  XOR U3442 ( .A(n3445), .B(n3446), .Z(n3450) );
  NOR U3443 ( .A(n3686), .B(n3746), .Z(n3448) );
  XOR U3444 ( .A(n3450), .B(n3448), .Z(n3486) );
  XOR U3445 ( .A(n3232), .B(n3483), .Z(n3485) );
  XOR U3446 ( .A(n3486), .B(n3485), .Z(n3386) );
  NOR U3447 ( .A(n3625), .B(n3636), .Z(n3535) );
  NOR U3448 ( .A(n3741), .B(n3776), .Z(n3233) );
  IV U3449 ( .A(n3233), .Z(n3536) );
  XOR U3450 ( .A(n3535), .B(n3536), .Z(n3540) );
  NOR U3451 ( .A(n3745), .B(n3787), .Z(n3538) );
  XOR U3452 ( .A(n3540), .B(n3538), .Z(n3434) );
  NOR U3453 ( .A(n3649), .B(n3619), .Z(n3430) );
  NOR U3454 ( .A(n3742), .B(n3763), .Z(n3234) );
  IV U3455 ( .A(n3234), .Z(n3431) );
  XOR U3456 ( .A(n3430), .B(n3431), .Z(n3433) );
  XOR U3457 ( .A(n3434), .B(n3433), .Z(n3235) );
  IV U3458 ( .A(n3235), .Z(n3387) );
  XOR U3459 ( .A(n3386), .B(n3387), .Z(n3389) );
  XOR U3460 ( .A(n3390), .B(n3389), .Z(n3379) );
  XOR U3461 ( .A(n3381), .B(n3379), .Z(n3382) );
  XOR U3462 ( .A(n3383), .B(n3382), .Z(n3236) );
  IV U3463 ( .A(n3236), .Z(n3368) );
  XOR U3464 ( .A(n3367), .B(n3368), .Z(n3412) );
  XOR U3465 ( .A(n3411), .B(n3412), .Z(n3359) );
  IV U3466 ( .A(n3237), .Z(n3238) );
  NOR U3467 ( .A(n3239), .B(n3238), .Z(n3243) );
  NOR U3468 ( .A(n3241), .B(n3240), .Z(n3242) );
  NOR U3469 ( .A(n3243), .B(n3242), .Z(n3357) );
  XOR U3470 ( .A(n3359), .B(n3357), .Z(n3361) );
  XOR U3471 ( .A(n3360), .B(n3361), .Z(n3345) );
  NOR U3472 ( .A(n3245), .B(n3244), .Z(n3249) );
  NOR U3473 ( .A(n3247), .B(n3246), .Z(n3248) );
  NOR U3474 ( .A(n3249), .B(n3248), .Z(n3401) );
  IV U3475 ( .A(n3250), .Z(n3252) );
  NOR U3476 ( .A(n3252), .B(n3251), .Z(n3256) );
  NOR U3477 ( .A(n3254), .B(n3253), .Z(n3255) );
  NOR U3478 ( .A(n3256), .B(n3255), .Z(n3419) );
  IV U3479 ( .A(n3257), .Z(n3259) );
  NOR U3480 ( .A(n3259), .B(n3258), .Z(n3264) );
  IV U3481 ( .A(n3260), .Z(n3261) );
  NOR U3482 ( .A(n3262), .B(n3261), .Z(n3263) );
  NOR U3483 ( .A(n3264), .B(n3263), .Z(n3417) );
  IV U3484 ( .A(n3265), .Z(n3267) );
  NOR U3485 ( .A(n3267), .B(n3266), .Z(n3271) );
  NOR U3486 ( .A(n3269), .B(n3268), .Z(n3270) );
  NOR U3487 ( .A(n3271), .B(n3270), .Z(n3416) );
  XOR U3488 ( .A(n3417), .B(n3416), .Z(n3272) );
  IV U3489 ( .A(n3272), .Z(n3418) );
  XOR U3490 ( .A(n3419), .B(n3418), .Z(n3403) );
  XOR U3491 ( .A(n3401), .B(n3403), .Z(n3405) );
  IV U3492 ( .A(n3273), .Z(n3275) );
  NOR U3493 ( .A(n3275), .B(n3274), .Z(n3279) );
  NOR U3494 ( .A(n3277), .B(n3276), .Z(n3278) );
  NOR U3495 ( .A(n3279), .B(n3278), .Z(n3280) );
  IV U3496 ( .A(n3280), .Z(n3404) );
  XOR U3497 ( .A(n3405), .B(n3404), .Z(n3343) );
  NOR U3498 ( .A(n3282), .B(n3281), .Z(n3286) );
  NOR U3499 ( .A(n3284), .B(n3283), .Z(n3285) );
  NOR U3500 ( .A(n3286), .B(n3285), .Z(n3287) );
  IV U3501 ( .A(n3287), .Z(n3353) );
  IV U3502 ( .A(n3288), .Z(n3289) );
  NOR U3503 ( .A(n3290), .B(n3289), .Z(n3294) );
  NOR U3504 ( .A(n3292), .B(n3291), .Z(n3293) );
  NOR U3505 ( .A(n3294), .B(n3293), .Z(n3352) );
  NOR U3506 ( .A(n3296), .B(n3295), .Z(n3301) );
  IV U3507 ( .A(n3297), .Z(n3298) );
  NOR U3508 ( .A(n3299), .B(n3298), .Z(n3300) );
  NOR U3509 ( .A(n3301), .B(n3300), .Z(n3350) );
  XOR U3510 ( .A(n3352), .B(n3350), .Z(n3354) );
  XOR U3511 ( .A(n3353), .B(n3354), .Z(n3342) );
  XOR U3512 ( .A(n3343), .B(n3342), .Z(n3344) );
  XOR U3513 ( .A(n3345), .B(n3344), .Z(n3335) );
  XOR U3514 ( .A(n3334), .B(n3335), .Z(n3339) );
  XOR U3515 ( .A(n3337), .B(n3339), .Z(n3327) );
  XOR U3516 ( .A(n3302), .B(n3327), .Z(n3331) );
  XOR U3517 ( .A(n3329), .B(n3331), .Z(n3320) );
  XOR U3518 ( .A(n3303), .B(n3320), .Z(n3324) );
  XOR U3519 ( .A(n3322), .B(n3324), .Z(n3315) );
  XOR U3520 ( .A(n3313), .B(n3315), .Z(n3317) );
  IV U3521 ( .A(n3304), .Z(n3305) );
  NOR U3522 ( .A(n3306), .B(n3305), .Z(n3311) );
  IV U3523 ( .A(n3307), .Z(n3308) );
  NOR U3524 ( .A(n3309), .B(n3308), .Z(n3310) );
  NOR U3525 ( .A(n3311), .B(n3310), .Z(n3312) );
  IV U3526 ( .A(n3312), .Z(n3316) );
  XOR U3527 ( .A(n3317), .B(n3316), .Z(N62) );
  IV U3528 ( .A(n3313), .Z(n3314) );
  NOR U3529 ( .A(n3315), .B(n3314), .Z(n3319) );
  NOR U3530 ( .A(n3317), .B(n3316), .Z(n3318) );
  NOR U3531 ( .A(n3319), .B(n3318), .Z(n3555) );
  NOR U3532 ( .A(n3321), .B(n3320), .Z(n3326) );
  IV U3533 ( .A(n3322), .Z(n3323) );
  NOR U3534 ( .A(n3324), .B(n3323), .Z(n3325) );
  NOR U3535 ( .A(n3326), .B(n3325), .Z(n3552) );
  NOR U3536 ( .A(n3328), .B(n3327), .Z(n3333) );
  IV U3537 ( .A(n3329), .Z(n3330) );
  NOR U3538 ( .A(n3331), .B(n3330), .Z(n3332) );
  NOR U3539 ( .A(n3333), .B(n3332), .Z(n3930) );
  IV U3540 ( .A(n3334), .Z(n3336) );
  NOR U3541 ( .A(n3336), .B(n3335), .Z(n3341) );
  IV U3542 ( .A(n3337), .Z(n3338) );
  NOR U3543 ( .A(n3339), .B(n3338), .Z(n3340) );
  NOR U3544 ( .A(n3341), .B(n3340), .Z(n3927) );
  NOR U3545 ( .A(n3343), .B(n3342), .Z(n3348) );
  IV U3546 ( .A(n3344), .Z(n3346) );
  NOR U3547 ( .A(n3346), .B(n3345), .Z(n3347) );
  NOR U3548 ( .A(n3348), .B(n3347), .Z(n3349) );
  IV U3549 ( .A(n3349), .Z(n3938) );
  IV U3550 ( .A(n3350), .Z(n3351) );
  NOR U3551 ( .A(n3352), .B(n3351), .Z(n3356) );
  NOR U3552 ( .A(n3354), .B(n3353), .Z(n3355) );
  NOR U3553 ( .A(n3356), .B(n3355), .Z(n3936) );
  IV U3554 ( .A(n3357), .Z(n3358) );
  NOR U3555 ( .A(n3359), .B(n3358), .Z(n3364) );
  IV U3556 ( .A(n3360), .Z(n3362) );
  NOR U3557 ( .A(n3362), .B(n3361), .Z(n3363) );
  NOR U3558 ( .A(n3364), .B(n3363), .Z(n3916) );
  NOR U3559 ( .A(n3366), .B(n3365), .Z(n3371) );
  IV U3560 ( .A(n3367), .Z(n3369) );
  NOR U3561 ( .A(n3369), .B(n3368), .Z(n3370) );
  NOR U3562 ( .A(n3371), .B(n3370), .Z(n3895) );
  NOR U3563 ( .A(n3373), .B(n3372), .Z(n3378) );
  IV U3564 ( .A(n3374), .Z(n3376) );
  NOR U3565 ( .A(n3376), .B(n3375), .Z(n3377) );
  NOR U3566 ( .A(n3378), .B(n3377), .Z(n3892) );
  IV U3567 ( .A(n3379), .Z(n3380) );
  NOR U3568 ( .A(n3381), .B(n3380), .Z(n3385) );
  NOR U3569 ( .A(n3383), .B(n3382), .Z(n3384) );
  NOR U3570 ( .A(n3385), .B(n3384), .Z(n3587) );
  IV U3571 ( .A(n3386), .Z(n3388) );
  NOR U3572 ( .A(n3388), .B(n3387), .Z(n3392) );
  NOR U3573 ( .A(n3390), .B(n3389), .Z(n3391) );
  NOR U3574 ( .A(n3392), .B(n3391), .Z(n3584) );
  IV U3575 ( .A(n3393), .Z(n3395) );
  NOR U3576 ( .A(n3395), .B(n3394), .Z(n3399) );
  NOR U3577 ( .A(n3397), .B(n3396), .Z(n3398) );
  NOR U3578 ( .A(n3399), .B(n3398), .Z(n3583) );
  XOR U3579 ( .A(n3584), .B(n3583), .Z(n3585) );
  XOR U3580 ( .A(n3587), .B(n3585), .Z(n3891) );
  XOR U3581 ( .A(n3892), .B(n3891), .Z(n3893) );
  XOR U3582 ( .A(n3895), .B(n3893), .Z(n3915) );
  XOR U3583 ( .A(n3916), .B(n3915), .Z(n3400) );
  IV U3584 ( .A(n3400), .Z(n3918) );
  IV U3585 ( .A(n3401), .Z(n3402) );
  NOR U3586 ( .A(n3403), .B(n3402), .Z(n3407) );
  NOR U3587 ( .A(n3405), .B(n3404), .Z(n3406) );
  NOR U3588 ( .A(n3407), .B(n3406), .Z(n3408) );
  IV U3589 ( .A(n3408), .Z(n3912) );
  NOR U3590 ( .A(n3410), .B(n3409), .Z(n3415) );
  IV U3591 ( .A(n3411), .Z(n3413) );
  NOR U3592 ( .A(n3413), .B(n3412), .Z(n3414) );
  NOR U3593 ( .A(n3415), .B(n3414), .Z(n3909) );
  NOR U3594 ( .A(n3417), .B(n3416), .Z(n3421) );
  NOR U3595 ( .A(n3419), .B(n3418), .Z(n3420) );
  NOR U3596 ( .A(n3421), .B(n3420), .Z(n3422) );
  IV U3597 ( .A(n3422), .Z(n3563) );
  NOR U3598 ( .A(n3424), .B(n3423), .Z(n3429) );
  IV U3599 ( .A(n3425), .Z(n3426) );
  NOR U3600 ( .A(n3427), .B(n3426), .Z(n3428) );
  NOR U3601 ( .A(n3429), .B(n3428), .Z(n3560) );
  IV U3602 ( .A(n3430), .Z(n3432) );
  NOR U3603 ( .A(n3432), .B(n3431), .Z(n3436) );
  NOR U3604 ( .A(n3434), .B(n3433), .Z(n3435) );
  NOR U3605 ( .A(n3436), .B(n3435), .Z(n3576) );
  IV U3606 ( .A(n3437), .Z(n3439) );
  NOR U3607 ( .A(n3439), .B(n3438), .Z(n3443) );
  NOR U3608 ( .A(n3441), .B(n3440), .Z(n3442) );
  NOR U3609 ( .A(n3443), .B(n3442), .Z(n3575) );
  XOR U3610 ( .A(n3576), .B(n3575), .Z(n3444) );
  IV U3611 ( .A(n3444), .Z(n3577) );
  IV U3612 ( .A(n3445), .Z(n3447) );
  NOR U3613 ( .A(n3447), .B(n3446), .Z(n3452) );
  IV U3614 ( .A(n3448), .Z(n3449) );
  NOR U3615 ( .A(n3450), .B(n3449), .Z(n3451) );
  NOR U3616 ( .A(n3452), .B(n3451), .Z(n3453) );
  IV U3617 ( .A(n3453), .Z(n3875) );
  NOR U3618 ( .A(n3682), .B(n3750), .Z(n3531) );
  IV U3619 ( .A(n3531), .Z(n3802) );
  NOR U3620 ( .A(n3454), .B(n3802), .Z(n3459) );
  IV U3621 ( .A(n3455), .Z(n3457) );
  NOR U3622 ( .A(n3457), .B(n3456), .Z(n3458) );
  NOR U3623 ( .A(n3459), .B(n3458), .Z(n3601) );
  NOR U3624 ( .A(n3649), .B(n3635), .Z(n3731) );
  NOR U3625 ( .A(n3782), .B(n3622), .Z(n3460) );
  IV U3626 ( .A(n3460), .Z(n3732) );
  XOR U3627 ( .A(n3731), .B(n3732), .Z(n3736) );
  NOR U3628 ( .A(n3461), .B(n3687), .Z(n3734) );
  XOR U3629 ( .A(n3736), .B(n3734), .Z(n3608) );
  NOR U3630 ( .A(n3739), .B(n3650), .Z(n3604) );
  NOR U3631 ( .A(n3645), .B(n3462), .Z(n3463) );
  IV U3632 ( .A(n3463), .Z(n3605) );
  XOR U3633 ( .A(n3604), .B(n3605), .Z(n3607) );
  XOR U3634 ( .A(n3608), .B(n3607), .Z(n3464) );
  IV U3635 ( .A(n3464), .Z(n3599) );
  NOR U3636 ( .A(n3627), .B(n3787), .Z(n3703) );
  NOR U3637 ( .A(n3465), .B(n3741), .Z(n3466) );
  IV U3638 ( .A(n3466), .Z(n3704) );
  XOR U3639 ( .A(n3703), .B(n3704), .Z(n3706) );
  NOR U3640 ( .A(n3788), .B(n3647), .Z(n3614) );
  NOR U3641 ( .A(n3742), .B(n3467), .Z(n3468) );
  IV U3642 ( .A(n3468), .Z(n3613) );
  IV U3643 ( .A(x[30]), .Z(n3774) );
  NOR U3644 ( .A(n3637), .B(n3774), .Z(n3611) );
  XOR U3645 ( .A(n3613), .B(n3611), .Z(n3616) );
  XOR U3646 ( .A(n3614), .B(n3616), .Z(n3707) );
  XOR U3647 ( .A(n3706), .B(n3707), .Z(n3597) );
  XOR U3648 ( .A(n3599), .B(n3597), .Z(n3600) );
  XOR U3649 ( .A(n3601), .B(n3600), .Z(n3873) );
  NOR U3650 ( .A(n3470), .B(n3469), .Z(n3474) );
  NOR U3651 ( .A(n3472), .B(n3471), .Z(n3473) );
  NOR U3652 ( .A(n3474), .B(n3473), .Z(n3871) );
  XOR U3653 ( .A(n3873), .B(n3871), .Z(n3874) );
  XOR U3654 ( .A(n3875), .B(n3874), .Z(n3578) );
  XOR U3655 ( .A(n3577), .B(n3578), .Z(n3888) );
  IV U3656 ( .A(n3475), .Z(n3477) );
  NOR U3657 ( .A(n3477), .B(n3476), .Z(n3482) );
  IV U3658 ( .A(n3478), .Z(n3480) );
  NOR U3659 ( .A(n3480), .B(n3479), .Z(n3481) );
  NOR U3660 ( .A(n3482), .B(n3481), .Z(n3868) );
  NOR U3661 ( .A(n3484), .B(n3483), .Z(n3488) );
  NOR U3662 ( .A(n3486), .B(n3485), .Z(n3487) );
  NOR U3663 ( .A(n3488), .B(n3487), .Z(n3866) );
  NOR U3664 ( .A(n3489), .B(n3779), .Z(n3528) );
  IV U3665 ( .A(n3528), .Z(n3809) );
  NOR U3666 ( .A(n3490), .B(n3809), .Z(n3495) );
  IV U3667 ( .A(n3491), .Z(n3492) );
  NOR U3668 ( .A(n3493), .B(n3492), .Z(n3494) );
  NOR U3669 ( .A(n3495), .B(n3494), .Z(n3594) );
  IV U3670 ( .A(n3496), .Z(n3498) );
  NOR U3671 ( .A(n3498), .B(n3497), .Z(n3503) );
  IV U3672 ( .A(n3499), .Z(n3500) );
  NOR U3673 ( .A(n3501), .B(n3500), .Z(n3502) );
  NOR U3674 ( .A(n3503), .B(n3502), .Z(n3591) );
  IV U3675 ( .A(n3504), .Z(n3506) );
  NOR U3676 ( .A(n3506), .B(n3505), .Z(n3510) );
  NOR U3677 ( .A(n3508), .B(n3507), .Z(n3509) );
  NOR U3678 ( .A(n3510), .B(n3509), .Z(n3590) );
  XOR U3679 ( .A(n3591), .B(n3590), .Z(n3592) );
  XOR U3680 ( .A(n3594), .B(n3592), .Z(n3865) );
  XOR U3681 ( .A(n3866), .B(n3865), .Z(n3511) );
  IV U3682 ( .A(n3511), .Z(n3867) );
  XOR U3683 ( .A(n3868), .B(n3867), .Z(n3885) );
  IV U3684 ( .A(n3512), .Z(n3514) );
  NOR U3685 ( .A(n3514), .B(n3513), .Z(n3519) );
  IV U3686 ( .A(n3515), .Z(n3516) );
  NOR U3687 ( .A(n3517), .B(n3516), .Z(n3518) );
  NOR U3688 ( .A(n3519), .B(n3518), .Z(n3568) );
  IV U3689 ( .A(n3520), .Z(n3522) );
  NOR U3690 ( .A(n3522), .B(n3521), .Z(n3526) );
  NOR U3691 ( .A(n3524), .B(n3523), .Z(n3525) );
  NOR U3692 ( .A(n3526), .B(n3525), .Z(n3849) );
  NOR U3693 ( .A(n3747), .B(n3740), .Z(n3527) );
  IV U3694 ( .A(n3527), .Z(n3808) );
  XOR U3695 ( .A(n3528), .B(n3808), .Z(n3812) );
  NOR U3696 ( .A(n3646), .B(n3621), .Z(n3810) );
  XOR U3697 ( .A(n3812), .B(n3810), .Z(n3832) );
  NOR U3698 ( .A(n3748), .B(n3683), .Z(n3828) );
  NOR U3699 ( .A(n3529), .B(n3763), .Z(n3530) );
  IV U3700 ( .A(n3530), .Z(n3829) );
  XOR U3701 ( .A(n3828), .B(n3829), .Z(n3831) );
  XOR U3702 ( .A(n3832), .B(n3831), .Z(n3719) );
  XOR U3703 ( .A(n3531), .B(n3801), .Z(n3805) );
  NOR U3704 ( .A(n3765), .B(n3780), .Z(n3803) );
  XOR U3705 ( .A(n3805), .B(n3803), .Z(n3718) );
  NOR U3706 ( .A(n3749), .B(n3766), .Z(n3716) );
  XOR U3707 ( .A(n3718), .B(n3716), .Z(n3720) );
  XOR U3708 ( .A(n3719), .B(n3720), .Z(n3846) );
  IV U3709 ( .A(o[29]), .Z(n3533) );
  NOR U3710 ( .A(n3533), .B(n3532), .Z(n3823) );
  NOR U3711 ( .A(n3773), .B(n3648), .Z(n3760) );
  IV U3712 ( .A(o[30]), .Z(n3761) );
  XOR U3713 ( .A(n3760), .B(n3761), .Z(n3822) );
  XOR U3714 ( .A(n3822), .B(n3534), .Z(n3824) );
  XOR U3715 ( .A(n3823), .B(n3824), .Z(n3845) );
  XOR U3716 ( .A(n3846), .B(n3845), .Z(n3847) );
  XOR U3717 ( .A(n3849), .B(n3847), .Z(n3567) );
  XOR U3718 ( .A(n3568), .B(n3567), .Z(n3570) );
  IV U3719 ( .A(n3535), .Z(n3537) );
  NOR U3720 ( .A(n3537), .B(n3536), .Z(n3542) );
  IV U3721 ( .A(n3538), .Z(n3539) );
  NOR U3722 ( .A(n3540), .B(n3539), .Z(n3541) );
  NOR U3723 ( .A(n3542), .B(n3541), .Z(n3856) );
  NOR U3724 ( .A(n3689), .B(n3781), .Z(n3543) );
  IV U3725 ( .A(n3543), .Z(n3669) );
  XOR U3726 ( .A(n3544), .B(n3669), .Z(n3673) );
  NOR U3727 ( .A(n3625), .B(n3620), .Z(n3671) );
  XOR U3728 ( .A(n3673), .B(n3671), .Z(n3728) );
  NOR U3729 ( .A(n3636), .B(n3619), .Z(n3724) );
  NOR U3730 ( .A(n3688), .B(n3764), .Z(n3545) );
  IV U3731 ( .A(n3545), .Z(n3725) );
  XOR U3732 ( .A(n3724), .B(n3725), .Z(n3727) );
  XOR U3733 ( .A(n3728), .B(n3727), .Z(n3852) );
  IV U3734 ( .A(y[30]), .Z(n3626) );
  NOR U3735 ( .A(n3680), .B(n3626), .Z(n3661) );
  NOR U3736 ( .A(n3775), .B(n3546), .Z(n3547) );
  IV U3737 ( .A(n3547), .Z(n3662) );
  XOR U3738 ( .A(n3661), .B(n3662), .Z(n3666) );
  NOR U3739 ( .A(n3745), .B(n3628), .Z(n3664) );
  XOR U3740 ( .A(n3666), .B(n3664), .Z(n3700) );
  NOR U3741 ( .A(n3746), .B(n3634), .Z(n3696) );
  NOR U3742 ( .A(n3549), .B(n3548), .Z(n3550) );
  IV U3743 ( .A(n3550), .Z(n3697) );
  XOR U3744 ( .A(n3696), .B(n3697), .Z(n3699) );
  XOR U3745 ( .A(n3700), .B(n3699), .Z(n3551) );
  IV U3746 ( .A(n3551), .Z(n3853) );
  XOR U3747 ( .A(n3852), .B(n3853), .Z(n3855) );
  XOR U3748 ( .A(n3856), .B(n3855), .Z(n3569) );
  XOR U3749 ( .A(n3570), .B(n3569), .Z(n3884) );
  XOR U3750 ( .A(n3885), .B(n3884), .Z(n3886) );
  XOR U3751 ( .A(n3888), .B(n3886), .Z(n3561) );
  XOR U3752 ( .A(n3560), .B(n3561), .Z(n3564) );
  XOR U3753 ( .A(n3563), .B(n3564), .Z(n3908) );
  XOR U3754 ( .A(n3909), .B(n3908), .Z(n3910) );
  XOR U3755 ( .A(n3912), .B(n3910), .Z(n3917) );
  XOR U3756 ( .A(n3918), .B(n3917), .Z(n3935) );
  XOR U3757 ( .A(n3936), .B(n3935), .Z(n3937) );
  XOR U3758 ( .A(n3938), .B(n3937), .Z(n3929) );
  XOR U3759 ( .A(n3927), .B(n3929), .Z(n3932) );
  XOR U3760 ( .A(n3930), .B(n3932), .Z(n3554) );
  XOR U3761 ( .A(n3552), .B(n3554), .Z(n3557) );
  XOR U3762 ( .A(n3555), .B(n3557), .Z(N63) );
  IV U3763 ( .A(n3552), .Z(n3553) );
  NOR U3764 ( .A(n3554), .B(n3553), .Z(n3559) );
  IV U3765 ( .A(n3555), .Z(n3556) );
  NOR U3766 ( .A(n3557), .B(n3556), .Z(n3558) );
  NOR U3767 ( .A(n3559), .B(n3558), .Z(n3926) );
  IV U3768 ( .A(n3560), .Z(n3562) );
  NOR U3769 ( .A(n3562), .B(n3561), .Z(n3566) );
  NOR U3770 ( .A(n3564), .B(n3563), .Z(n3565) );
  NOR U3771 ( .A(n3566), .B(n3565), .Z(n3907) );
  NOR U3772 ( .A(n3568), .B(n3567), .Z(n3574) );
  IV U3773 ( .A(n3569), .Z(n3572) );
  IV U3774 ( .A(n3570), .Z(n3571) );
  NOR U3775 ( .A(n3572), .B(n3571), .Z(n3573) );
  NOR U3776 ( .A(n3574), .B(n3573), .Z(n3582) );
  NOR U3777 ( .A(n3576), .B(n3575), .Z(n3580) );
  NOR U3778 ( .A(n3578), .B(n3577), .Z(n3579) );
  NOR U3779 ( .A(n3580), .B(n3579), .Z(n3581) );
  XOR U3780 ( .A(n3582), .B(n3581), .Z(n3905) );
  NOR U3781 ( .A(n3584), .B(n3583), .Z(n3589) );
  IV U3782 ( .A(n3585), .Z(n3586) );
  NOR U3783 ( .A(n3587), .B(n3586), .Z(n3588) );
  NOR U3784 ( .A(n3589), .B(n3588), .Z(n3903) );
  NOR U3785 ( .A(n3591), .B(n3590), .Z(n3596) );
  IV U3786 ( .A(n3592), .Z(n3593) );
  NOR U3787 ( .A(n3594), .B(n3593), .Z(n3595) );
  NOR U3788 ( .A(n3596), .B(n3595), .Z(n3883) );
  IV U3789 ( .A(n3597), .Z(n3598) );
  NOR U3790 ( .A(n3599), .B(n3598), .Z(n3603) );
  NOR U3791 ( .A(n3601), .B(n3600), .Z(n3602) );
  NOR U3792 ( .A(n3603), .B(n3602), .Z(n3864) );
  IV U3793 ( .A(n3604), .Z(n3606) );
  NOR U3794 ( .A(n3606), .B(n3605), .Z(n3610) );
  NOR U3795 ( .A(n3608), .B(n3607), .Z(n3609) );
  NOR U3796 ( .A(n3610), .B(n3609), .Z(n3844) );
  IV U3797 ( .A(n3611), .Z(n3612) );
  NOR U3798 ( .A(n3613), .B(n3612), .Z(n3618) );
  IV U3799 ( .A(n3614), .Z(n3615) );
  NOR U3800 ( .A(n3616), .B(n3615), .Z(n3617) );
  NOR U3801 ( .A(n3618), .B(n3617), .Z(n3715) );
  NOR U3802 ( .A(n3620), .B(n3619), .Z(n3624) );
  NOR U3803 ( .A(n3622), .B(n3621), .Z(n3623) );
  XOR U3804 ( .A(n3624), .B(n3623), .Z(n3632) );
  NOR U3805 ( .A(n3626), .B(n3625), .Z(n3630) );
  NOR U3806 ( .A(n3628), .B(n3627), .Z(n3629) );
  XOR U3807 ( .A(n3630), .B(n3629), .Z(n3631) );
  XOR U3808 ( .A(n3632), .B(n3631), .Z(n3660) );
  NOR U3809 ( .A(n3634), .B(n3633), .Z(n3644) );
  NOR U3810 ( .A(n3636), .B(n3635), .Z(n3640) );
  IV U3811 ( .A(x[31]), .Z(n3638) );
  NOR U3812 ( .A(n3638), .B(n3637), .Z(n3639) );
  XOR U3813 ( .A(n3640), .B(n3639), .Z(n3641) );
  XOR U3814 ( .A(n3642), .B(n3641), .Z(n3643) );
  XOR U3815 ( .A(n3644), .B(n3643), .Z(n3658) );
  NOR U3816 ( .A(n3646), .B(n3645), .Z(n3656) );
  NOR U3817 ( .A(n3648), .B(n3647), .Z(n3652) );
  NOR U3818 ( .A(n3650), .B(n3649), .Z(n3651) );
  XOR U3819 ( .A(n3652), .B(n3651), .Z(n3653) );
  XOR U3820 ( .A(n3654), .B(n3653), .Z(n3655) );
  XOR U3821 ( .A(n3656), .B(n3655), .Z(n3657) );
  XOR U3822 ( .A(n3658), .B(n3657), .Z(n3659) );
  XOR U3823 ( .A(n3660), .B(n3659), .Z(n3679) );
  IV U3824 ( .A(n3661), .Z(n3663) );
  NOR U3825 ( .A(n3663), .B(n3662), .Z(n3668) );
  IV U3826 ( .A(n3664), .Z(n3665) );
  NOR U3827 ( .A(n3666), .B(n3665), .Z(n3667) );
  NOR U3828 ( .A(n3668), .B(n3667), .Z(n3677) );
  NOR U3829 ( .A(n3670), .B(n3669), .Z(n3675) );
  IV U3830 ( .A(n3671), .Z(n3672) );
  NOR U3831 ( .A(n3673), .B(n3672), .Z(n3674) );
  NOR U3832 ( .A(n3675), .B(n3674), .Z(n3676) );
  XOR U3833 ( .A(n3677), .B(n3676), .Z(n3678) );
  XOR U3834 ( .A(n3679), .B(n3678), .Z(n3695) );
  IV U3835 ( .A(y[31]), .Z(n3681) );
  NOR U3836 ( .A(n3681), .B(n3680), .Z(n3685) );
  NOR U3837 ( .A(n3683), .B(n3682), .Z(n3684) );
  XOR U3838 ( .A(n3685), .B(n3684), .Z(n3693) );
  NOR U3839 ( .A(n3687), .B(n3686), .Z(n3691) );
  NOR U3840 ( .A(n3689), .B(n3688), .Z(n3690) );
  XOR U3841 ( .A(n3691), .B(n3690), .Z(n3692) );
  XOR U3842 ( .A(n3693), .B(n3692), .Z(n3694) );
  XOR U3843 ( .A(n3695), .B(n3694), .Z(n3713) );
  IV U3844 ( .A(n3696), .Z(n3698) );
  NOR U3845 ( .A(n3698), .B(n3697), .Z(n3702) );
  NOR U3846 ( .A(n3700), .B(n3699), .Z(n3701) );
  NOR U3847 ( .A(n3702), .B(n3701), .Z(n3711) );
  IV U3848 ( .A(n3703), .Z(n3705) );
  NOR U3849 ( .A(n3705), .B(n3704), .Z(n3709) );
  NOR U3850 ( .A(n3707), .B(n3706), .Z(n3708) );
  NOR U3851 ( .A(n3709), .B(n3708), .Z(n3710) );
  XOR U3852 ( .A(n3711), .B(n3710), .Z(n3712) );
  XOR U3853 ( .A(n3713), .B(n3712), .Z(n3714) );
  XOR U3854 ( .A(n3715), .B(n3714), .Z(n3842) );
  IV U3855 ( .A(n3716), .Z(n3717) );
  NOR U3856 ( .A(n3718), .B(n3717), .Z(n3723) );
  IV U3857 ( .A(n3719), .Z(n3721) );
  NOR U3858 ( .A(n3721), .B(n3720), .Z(n3722) );
  NOR U3859 ( .A(n3723), .B(n3722), .Z(n3840) );
  IV U3860 ( .A(n3724), .Z(n3726) );
  NOR U3861 ( .A(n3726), .B(n3725), .Z(n3730) );
  NOR U3862 ( .A(n3728), .B(n3727), .Z(n3729) );
  NOR U3863 ( .A(n3730), .B(n3729), .Z(n3820) );
  IV U3864 ( .A(n3731), .Z(n3733) );
  NOR U3865 ( .A(n3733), .B(n3732), .Z(n3738) );
  IV U3866 ( .A(n3734), .Z(n3735) );
  NOR U3867 ( .A(n3736), .B(n3735), .Z(n3737) );
  NOR U3868 ( .A(n3738), .B(n3737), .Z(n3800) );
  NOR U3869 ( .A(n3740), .B(n3739), .Z(n3744) );
  NOR U3870 ( .A(n3742), .B(n3741), .Z(n3743) );
  XOR U3871 ( .A(n3744), .B(n3743), .Z(n3759) );
  NOR U3872 ( .A(n3746), .B(n3745), .Z(n3757) );
  NOR U3873 ( .A(n3748), .B(n3747), .Z(n3755) );
  NOR U3874 ( .A(n3750), .B(n3749), .Z(n3753) );
  XOR U3875 ( .A(n3751), .B(o[31]), .Z(n3752) );
  XOR U3876 ( .A(n3753), .B(n3752), .Z(n3754) );
  XOR U3877 ( .A(n3755), .B(n3754), .Z(n3756) );
  XOR U3878 ( .A(n3757), .B(n3756), .Z(n3758) );
  XOR U3879 ( .A(n3759), .B(n3758), .Z(n3772) );
  IV U3880 ( .A(n3760), .Z(n3762) );
  NOR U3881 ( .A(n3762), .B(n3761), .Z(n3770) );
  NOR U3882 ( .A(n3764), .B(n3763), .Z(n3768) );
  NOR U3883 ( .A(n3766), .B(n3765), .Z(n3767) );
  XOR U3884 ( .A(n3768), .B(n3767), .Z(n3769) );
  XOR U3885 ( .A(n3770), .B(n3769), .Z(n3771) );
  XOR U3886 ( .A(n3772), .B(n3771), .Z(n3798) );
  NOR U3887 ( .A(n3774), .B(n3773), .Z(n3778) );
  NOR U3888 ( .A(n3776), .B(n3775), .Z(n3777) );
  XOR U3889 ( .A(n3778), .B(n3777), .Z(n3786) );
  NOR U3890 ( .A(n3780), .B(n3779), .Z(n3784) );
  NOR U3891 ( .A(n3782), .B(n3781), .Z(n3783) );
  XOR U3892 ( .A(n3784), .B(n3783), .Z(n3785) );
  XOR U3893 ( .A(n3786), .B(n3785), .Z(n3796) );
  NOR U3894 ( .A(n3788), .B(n3787), .Z(n3792) );
  XOR U3895 ( .A(n3790), .B(n3789), .Z(n3791) );
  XOR U3896 ( .A(n3792), .B(n3791), .Z(n3793) );
  XOR U3897 ( .A(n3794), .B(n3793), .Z(n3795) );
  XOR U3898 ( .A(n3796), .B(n3795), .Z(n3797) );
  XOR U3899 ( .A(n3798), .B(n3797), .Z(n3799) );
  XOR U3900 ( .A(n3800), .B(n3799), .Z(n3818) );
  NOR U3901 ( .A(n3802), .B(n3801), .Z(n3807) );
  IV U3902 ( .A(n3803), .Z(n3804) );
  NOR U3903 ( .A(n3805), .B(n3804), .Z(n3806) );
  NOR U3904 ( .A(n3807), .B(n3806), .Z(n3816) );
  NOR U3905 ( .A(n3809), .B(n3808), .Z(n3814) );
  IV U3906 ( .A(n3810), .Z(n3811) );
  NOR U3907 ( .A(n3812), .B(n3811), .Z(n3813) );
  NOR U3908 ( .A(n3814), .B(n3813), .Z(n3815) );
  XOR U3909 ( .A(n3816), .B(n3815), .Z(n3817) );
  XOR U3910 ( .A(n3818), .B(n3817), .Z(n3819) );
  XOR U3911 ( .A(n3820), .B(n3819), .Z(n3838) );
  NOR U3912 ( .A(n3822), .B(n3821), .Z(n3827) );
  IV U3913 ( .A(n3823), .Z(n3825) );
  NOR U3914 ( .A(n3825), .B(n3824), .Z(n3826) );
  NOR U3915 ( .A(n3827), .B(n3826), .Z(n3836) );
  IV U3916 ( .A(n3828), .Z(n3830) );
  NOR U3917 ( .A(n3830), .B(n3829), .Z(n3834) );
  NOR U3918 ( .A(n3832), .B(n3831), .Z(n3833) );
  NOR U3919 ( .A(n3834), .B(n3833), .Z(n3835) );
  XOR U3920 ( .A(n3836), .B(n3835), .Z(n3837) );
  XOR U3921 ( .A(n3838), .B(n3837), .Z(n3839) );
  XOR U3922 ( .A(n3840), .B(n3839), .Z(n3841) );
  XOR U3923 ( .A(n3842), .B(n3841), .Z(n3843) );
  XOR U3924 ( .A(n3844), .B(n3843), .Z(n3862) );
  NOR U3925 ( .A(n3846), .B(n3845), .Z(n3851) );
  IV U3926 ( .A(n3847), .Z(n3848) );
  NOR U3927 ( .A(n3849), .B(n3848), .Z(n3850) );
  NOR U3928 ( .A(n3851), .B(n3850), .Z(n3860) );
  IV U3929 ( .A(n3852), .Z(n3854) );
  NOR U3930 ( .A(n3854), .B(n3853), .Z(n3858) );
  NOR U3931 ( .A(n3856), .B(n3855), .Z(n3857) );
  NOR U3932 ( .A(n3858), .B(n3857), .Z(n3859) );
  XOR U3933 ( .A(n3860), .B(n3859), .Z(n3861) );
  XOR U3934 ( .A(n3862), .B(n3861), .Z(n3863) );
  XOR U3935 ( .A(n3864), .B(n3863), .Z(n3881) );
  NOR U3936 ( .A(n3866), .B(n3865), .Z(n3870) );
  NOR U3937 ( .A(n3868), .B(n3867), .Z(n3869) );
  NOR U3938 ( .A(n3870), .B(n3869), .Z(n3879) );
  IV U3939 ( .A(n3871), .Z(n3872) );
  NOR U3940 ( .A(n3873), .B(n3872), .Z(n3877) );
  NOR U3941 ( .A(n3875), .B(n3874), .Z(n3876) );
  NOR U3942 ( .A(n3877), .B(n3876), .Z(n3878) );
  XOR U3943 ( .A(n3879), .B(n3878), .Z(n3880) );
  XOR U3944 ( .A(n3881), .B(n3880), .Z(n3882) );
  XOR U3945 ( .A(n3883), .B(n3882), .Z(n3901) );
  NOR U3946 ( .A(n3885), .B(n3884), .Z(n3890) );
  IV U3947 ( .A(n3886), .Z(n3887) );
  NOR U3948 ( .A(n3888), .B(n3887), .Z(n3889) );
  NOR U3949 ( .A(n3890), .B(n3889), .Z(n3899) );
  NOR U3950 ( .A(n3892), .B(n3891), .Z(n3897) );
  IV U3951 ( .A(n3893), .Z(n3894) );
  NOR U3952 ( .A(n3895), .B(n3894), .Z(n3896) );
  NOR U3953 ( .A(n3897), .B(n3896), .Z(n3898) );
  XOR U3954 ( .A(n3899), .B(n3898), .Z(n3900) );
  XOR U3955 ( .A(n3901), .B(n3900), .Z(n3902) );
  XOR U3956 ( .A(n3903), .B(n3902), .Z(n3904) );
  XOR U3957 ( .A(n3905), .B(n3904), .Z(n3906) );
  XOR U3958 ( .A(n3907), .B(n3906), .Z(n3924) );
  NOR U3959 ( .A(n3909), .B(n3908), .Z(n3914) );
  IV U3960 ( .A(n3910), .Z(n3911) );
  NOR U3961 ( .A(n3912), .B(n3911), .Z(n3913) );
  NOR U3962 ( .A(n3914), .B(n3913), .Z(n3922) );
  NOR U3963 ( .A(n3916), .B(n3915), .Z(n3920) );
  NOR U3964 ( .A(n3918), .B(n3917), .Z(n3919) );
  NOR U3965 ( .A(n3920), .B(n3919), .Z(n3921) );
  XOR U3966 ( .A(n3922), .B(n3921), .Z(n3923) );
  XOR U3967 ( .A(n3924), .B(n3923), .Z(n3925) );
  XOR U3968 ( .A(n3926), .B(n3925), .Z(n3945) );
  IV U3969 ( .A(n3927), .Z(n3928) );
  NOR U3970 ( .A(n3929), .B(n3928), .Z(n3934) );
  IV U3971 ( .A(n3930), .Z(n3931) );
  NOR U3972 ( .A(n3932), .B(n3931), .Z(n3933) );
  NOR U3973 ( .A(n3934), .B(n3933), .Z(n3943) );
  NOR U3974 ( .A(n3936), .B(n3935), .Z(n3941) );
  IV U3975 ( .A(n3937), .Z(n3939) );
  NOR U3976 ( .A(n3939), .B(n3938), .Z(n3940) );
  NOR U3977 ( .A(n3941), .B(n3940), .Z(n3942) );
  XOR U3978 ( .A(n3943), .B(n3942), .Z(n3944) );
  XOR U3979 ( .A(n3945), .B(n3944), .Z(N64) );
endmodule

