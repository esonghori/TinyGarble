
module mult_N64_CC8 ( clk, rst, a, b, c );
  input [63:0] a;
  input [7:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720;
  wire   [127:0] sreg;

  DFF \sreg_reg[119]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[61]) );
  DFF \sreg_reg[60]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[60]) );
  DFF \sreg_reg[59]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[59]) );
  DFF \sreg_reg[58]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[58]) );
  DFF \sreg_reg[57]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[57]) );
  DFF \sreg_reg[56]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[56]) );
  DFF \sreg_reg[55]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U11 ( .A(n553), .B(n551), .Z(n1) );
  XOR U12 ( .A(n551), .B(n553), .Z(n2) );
  NANDN U13 ( .A(n552), .B(n2), .Z(n3) );
  NAND U14 ( .A(n1), .B(n3), .Z(n603) );
  NAND U15 ( .A(n794), .B(n795), .Z(n4) );
  NANDN U16 ( .A(n793), .B(n792), .Z(n5) );
  NAND U17 ( .A(n4), .B(n5), .Z(n802) );
  NAND U18 ( .A(n1241), .B(n1242), .Z(n6) );
  NANDN U19 ( .A(n1240), .B(n1239), .Z(n7) );
  NAND U20 ( .A(n6), .B(n7), .Z(n1249) );
  NAND U21 ( .A(n620), .B(n621), .Z(n8) );
  NANDN U22 ( .A(n619), .B(n618), .Z(n9) );
  NAND U23 ( .A(n8), .B(n9), .Z(n680) );
  NAND U24 ( .A(n844), .B(n845), .Z(n10) );
  NANDN U25 ( .A(n843), .B(n842), .Z(n11) );
  NAND U26 ( .A(n10), .B(n11), .Z(n904) );
  NAND U27 ( .A(n1068), .B(n1069), .Z(n12) );
  NANDN U28 ( .A(n1067), .B(n1066), .Z(n13) );
  NAND U29 ( .A(n12), .B(n13), .Z(n1128) );
  NAND U30 ( .A(n1291), .B(n1292), .Z(n14) );
  NANDN U31 ( .A(n1290), .B(n1289), .Z(n15) );
  NAND U32 ( .A(n14), .B(n15), .Z(n1351) );
  NAND U33 ( .A(n1402), .B(n1403), .Z(n16) );
  NANDN U34 ( .A(n1401), .B(n1400), .Z(n17) );
  NAND U35 ( .A(n16), .B(n17), .Z(n1462) );
  NAND U36 ( .A(n1513), .B(n1514), .Z(n18) );
  NANDN U37 ( .A(n1512), .B(n1511), .Z(n19) );
  NAND U38 ( .A(n18), .B(n19), .Z(n1573) );
  NAND U39 ( .A(n1624), .B(n1625), .Z(n20) );
  NANDN U40 ( .A(n1623), .B(n1622), .Z(n21) );
  NAND U41 ( .A(n20), .B(n21), .Z(n1684) );
  NAND U42 ( .A(n1735), .B(n1736), .Z(n22) );
  NANDN U43 ( .A(n1734), .B(n1733), .Z(n23) );
  NAND U44 ( .A(n22), .B(n23), .Z(n1795) );
  NAND U45 ( .A(n1846), .B(n1847), .Z(n24) );
  NANDN U46 ( .A(n1845), .B(n1844), .Z(n25) );
  NAND U47 ( .A(n24), .B(n25), .Z(n1906) );
  NAND U48 ( .A(n1957), .B(n1958), .Z(n26) );
  NANDN U49 ( .A(n1956), .B(n1955), .Z(n27) );
  NAND U50 ( .A(n26), .B(n27), .Z(n2017) );
  NAND U51 ( .A(n2068), .B(n2069), .Z(n28) );
  NANDN U52 ( .A(n2067), .B(n2066), .Z(n29) );
  NAND U53 ( .A(n28), .B(n29), .Z(n2128) );
  NAND U54 ( .A(n2179), .B(n2180), .Z(n30) );
  NANDN U55 ( .A(n2178), .B(n2177), .Z(n31) );
  NAND U56 ( .A(n30), .B(n31), .Z(n2239) );
  NAND U57 ( .A(n2290), .B(n2291), .Z(n32) );
  NANDN U58 ( .A(n2289), .B(n2288), .Z(n33) );
  NAND U59 ( .A(n32), .B(n33), .Z(n2350) );
  NOR U60 ( .A(b[4]), .B(n248), .Z(n34) );
  NANDN U61 ( .A(n247), .B(n2658), .Z(n35) );
  NAND U62 ( .A(n34), .B(n35), .Z(n36) );
  NANDN U63 ( .A(a[0]), .B(n2628), .Z(n37) );
  NAND U64 ( .A(n36), .B(n37), .Z(n332) );
  NAND U65 ( .A(n2402), .B(n2403), .Z(n38) );
  NANDN U66 ( .A(n2401), .B(n2400), .Z(n39) );
  NAND U67 ( .A(n38), .B(n39), .Z(n2464) );
  XOR U68 ( .A(n300), .B(n299), .Z(n40) );
  NANDN U69 ( .A(n298), .B(n40), .Z(n41) );
  NAND U70 ( .A(n300), .B(n299), .Z(n42) );
  AND U71 ( .A(n41), .B(n42), .Z(n330) );
  NAND U72 ( .A(n616), .B(n617), .Z(n43) );
  NANDN U73 ( .A(n615), .B(n614), .Z(n44) );
  NAND U74 ( .A(n43), .B(n44), .Z(n654) );
  NAND U75 ( .A(n728), .B(n729), .Z(n45) );
  NANDN U76 ( .A(n727), .B(n726), .Z(n46) );
  NAND U77 ( .A(n45), .B(n46), .Z(n768) );
  NAND U78 ( .A(n840), .B(n841), .Z(n47) );
  NANDN U79 ( .A(n839), .B(n838), .Z(n48) );
  NAND U80 ( .A(n47), .B(n48), .Z(n878) );
  NAND U81 ( .A(n951), .B(n952), .Z(n49) );
  NANDN U82 ( .A(n950), .B(n949), .Z(n50) );
  NAND U83 ( .A(n49), .B(n50), .Z(n991) );
  NAND U84 ( .A(n1064), .B(n1065), .Z(n51) );
  NANDN U85 ( .A(n1063), .B(n1062), .Z(n52) );
  NAND U86 ( .A(n51), .B(n52), .Z(n1102) );
  NAND U87 ( .A(n1176), .B(n1177), .Z(n53) );
  NANDN U88 ( .A(n1175), .B(n1174), .Z(n54) );
  NAND U89 ( .A(n53), .B(n54), .Z(n1216) );
  NAND U90 ( .A(n1287), .B(n1288), .Z(n55) );
  NANDN U91 ( .A(n1286), .B(n1285), .Z(n56) );
  NAND U92 ( .A(n55), .B(n56), .Z(n1325) );
  NAND U93 ( .A(n1398), .B(n1399), .Z(n57) );
  NANDN U94 ( .A(n1397), .B(n1396), .Z(n58) );
  NAND U95 ( .A(n57), .B(n58), .Z(n1436) );
  NAND U96 ( .A(n1509), .B(n1510), .Z(n59) );
  NANDN U97 ( .A(n1508), .B(n1507), .Z(n60) );
  NAND U98 ( .A(n59), .B(n60), .Z(n1547) );
  NAND U99 ( .A(n1620), .B(n1621), .Z(n61) );
  NANDN U100 ( .A(n1619), .B(n1618), .Z(n62) );
  NAND U101 ( .A(n61), .B(n62), .Z(n1658) );
  NAND U102 ( .A(n1731), .B(n1732), .Z(n63) );
  NANDN U103 ( .A(n1730), .B(n1729), .Z(n64) );
  NAND U104 ( .A(n63), .B(n64), .Z(n1769) );
  NAND U105 ( .A(n1842), .B(n1843), .Z(n65) );
  NANDN U106 ( .A(n1841), .B(n1840), .Z(n66) );
  NAND U107 ( .A(n65), .B(n66), .Z(n1880) );
  NAND U108 ( .A(n1953), .B(n1954), .Z(n67) );
  NANDN U109 ( .A(n1952), .B(n1951), .Z(n68) );
  NAND U110 ( .A(n67), .B(n68), .Z(n1991) );
  NAND U111 ( .A(n2064), .B(n2065), .Z(n69) );
  NANDN U112 ( .A(n2063), .B(n2062), .Z(n70) );
  NAND U113 ( .A(n69), .B(n70), .Z(n2102) );
  NAND U114 ( .A(n2175), .B(n2176), .Z(n71) );
  NANDN U115 ( .A(n2174), .B(n2173), .Z(n72) );
  NAND U116 ( .A(n71), .B(n72), .Z(n2213) );
  NAND U117 ( .A(n2286), .B(n2287), .Z(n73) );
  NANDN U118 ( .A(n2285), .B(n2284), .Z(n74) );
  NAND U119 ( .A(n73), .B(n74), .Z(n2324) );
  NAND U120 ( .A(n2398), .B(n2399), .Z(n75) );
  NANDN U121 ( .A(n2397), .B(n2396), .Z(n76) );
  NAND U122 ( .A(n75), .B(n76), .Z(n2437) );
  NAND U123 ( .A(n549), .B(n550), .Z(n77) );
  NANDN U124 ( .A(n548), .B(n547), .Z(n78) );
  NAND U125 ( .A(n77), .B(n78), .Z(n606) );
  NAND U126 ( .A(n657), .B(n658), .Z(n79) );
  NANDN U127 ( .A(n656), .B(n655), .Z(n80) );
  NAND U128 ( .A(n79), .B(n80), .Z(n718) );
  NAND U129 ( .A(n771), .B(n772), .Z(n81) );
  NANDN U130 ( .A(n770), .B(n769), .Z(n82) );
  NAND U131 ( .A(n81), .B(n82), .Z(n830) );
  NAND U132 ( .A(n881), .B(n882), .Z(n83) );
  NANDN U133 ( .A(n880), .B(n879), .Z(n84) );
  NAND U134 ( .A(n83), .B(n84), .Z(n941) );
  NAND U135 ( .A(n994), .B(n995), .Z(n85) );
  NANDN U136 ( .A(n993), .B(n992), .Z(n86) );
  NAND U137 ( .A(n85), .B(n86), .Z(n1054) );
  NAND U138 ( .A(n1105), .B(n1106), .Z(n87) );
  NANDN U139 ( .A(n1104), .B(n1103), .Z(n88) );
  NAND U140 ( .A(n87), .B(n88), .Z(n1166) );
  NAND U141 ( .A(n1219), .B(n1220), .Z(n89) );
  NANDN U142 ( .A(n1218), .B(n1217), .Z(n90) );
  NAND U143 ( .A(n89), .B(n90), .Z(n1277) );
  NAND U144 ( .A(n1328), .B(n1329), .Z(n91) );
  NANDN U145 ( .A(n1327), .B(n1326), .Z(n92) );
  NAND U146 ( .A(n91), .B(n92), .Z(n1388) );
  NAND U147 ( .A(n1439), .B(n1440), .Z(n93) );
  NANDN U148 ( .A(n1438), .B(n1437), .Z(n94) );
  NAND U149 ( .A(n93), .B(n94), .Z(n1499) );
  NAND U150 ( .A(n1550), .B(n1551), .Z(n95) );
  NANDN U151 ( .A(n1549), .B(n1548), .Z(n96) );
  NAND U152 ( .A(n95), .B(n96), .Z(n1610) );
  NAND U153 ( .A(n1661), .B(n1662), .Z(n97) );
  NANDN U154 ( .A(n1660), .B(n1659), .Z(n98) );
  NAND U155 ( .A(n97), .B(n98), .Z(n1721) );
  NAND U156 ( .A(n1772), .B(n1773), .Z(n99) );
  NANDN U157 ( .A(n1771), .B(n1770), .Z(n100) );
  NAND U158 ( .A(n99), .B(n100), .Z(n1832) );
  NAND U159 ( .A(n1883), .B(n1884), .Z(n101) );
  NANDN U160 ( .A(n1882), .B(n1881), .Z(n102) );
  NAND U161 ( .A(n101), .B(n102), .Z(n1943) );
  NAND U162 ( .A(n1994), .B(n1995), .Z(n103) );
  NANDN U163 ( .A(n1993), .B(n1992), .Z(n104) );
  NAND U164 ( .A(n103), .B(n104), .Z(n2054) );
  NAND U165 ( .A(n2105), .B(n2106), .Z(n105) );
  NANDN U166 ( .A(n2104), .B(n2103), .Z(n106) );
  NAND U167 ( .A(n105), .B(n106), .Z(n2165) );
  NAND U168 ( .A(n2216), .B(n2217), .Z(n107) );
  NANDN U169 ( .A(n2215), .B(n2214), .Z(n108) );
  NAND U170 ( .A(n107), .B(n108), .Z(n2276) );
  NAND U171 ( .A(n2327), .B(n2328), .Z(n109) );
  NANDN U172 ( .A(n2326), .B(n2325), .Z(n110) );
  NAND U173 ( .A(n109), .B(n110), .Z(n2388) );
  NAND U174 ( .A(n355), .B(n356), .Z(n111) );
  NANDN U175 ( .A(n354), .B(n353), .Z(n112) );
  NAND U176 ( .A(n111), .B(n112), .Z(n397) );
  NAND U177 ( .A(n2440), .B(n2441), .Z(n113) );
  NANDN U178 ( .A(n2439), .B(n2438), .Z(n114) );
  NAND U179 ( .A(n113), .B(n114), .Z(n2479) );
  NANDN U180 ( .A(n335), .B(n334), .Z(n115) );
  NANDN U181 ( .A(n333), .B(n332), .Z(n116) );
  NAND U182 ( .A(n115), .B(n116), .Z(n347) );
  NAND U183 ( .A(n545), .B(n546), .Z(n117) );
  NANDN U184 ( .A(n544), .B(n543), .Z(n118) );
  NAND U185 ( .A(n117), .B(n118), .Z(n580) );
  NAND U186 ( .A(n653), .B(n654), .Z(n119) );
  NANDN U187 ( .A(n652), .B(n651), .Z(n120) );
  NAND U188 ( .A(n119), .B(n120), .Z(n691) );
  NAND U189 ( .A(n767), .B(n768), .Z(n121) );
  NANDN U190 ( .A(n766), .B(n765), .Z(n122) );
  NAND U191 ( .A(n121), .B(n122), .Z(n804) );
  NAND U192 ( .A(n877), .B(n878), .Z(n123) );
  NANDN U193 ( .A(n876), .B(n875), .Z(n124) );
  NAND U194 ( .A(n123), .B(n124), .Z(n915) );
  NAND U195 ( .A(n990), .B(n991), .Z(n125) );
  NANDN U196 ( .A(n989), .B(n988), .Z(n126) );
  NAND U197 ( .A(n125), .B(n126), .Z(n1028) );
  NAND U198 ( .A(n1101), .B(n1102), .Z(n127) );
  NANDN U199 ( .A(n1100), .B(n1099), .Z(n128) );
  NAND U200 ( .A(n127), .B(n128), .Z(n1139) );
  NAND U201 ( .A(n1215), .B(n1216), .Z(n129) );
  NANDN U202 ( .A(n1214), .B(n1213), .Z(n130) );
  NAND U203 ( .A(n129), .B(n130), .Z(n1251) );
  NAND U204 ( .A(n1324), .B(n1325), .Z(n131) );
  NANDN U205 ( .A(n1323), .B(n1322), .Z(n132) );
  NAND U206 ( .A(n131), .B(n132), .Z(n1362) );
  NAND U207 ( .A(n1435), .B(n1436), .Z(n133) );
  NANDN U208 ( .A(n1434), .B(n1433), .Z(n134) );
  NAND U209 ( .A(n133), .B(n134), .Z(n1473) );
  NAND U210 ( .A(n1546), .B(n1547), .Z(n135) );
  NANDN U211 ( .A(n1545), .B(n1544), .Z(n136) );
  NAND U212 ( .A(n135), .B(n136), .Z(n1584) );
  NAND U213 ( .A(n1657), .B(n1658), .Z(n137) );
  NANDN U214 ( .A(n1656), .B(n1655), .Z(n138) );
  NAND U215 ( .A(n137), .B(n138), .Z(n1695) );
  NAND U216 ( .A(n1768), .B(n1769), .Z(n139) );
  NANDN U217 ( .A(n1767), .B(n1766), .Z(n140) );
  NAND U218 ( .A(n139), .B(n140), .Z(n1806) );
  NAND U219 ( .A(n1879), .B(n1880), .Z(n141) );
  NANDN U220 ( .A(n1878), .B(n1877), .Z(n142) );
  NAND U221 ( .A(n141), .B(n142), .Z(n1917) );
  NAND U222 ( .A(n1990), .B(n1991), .Z(n143) );
  NANDN U223 ( .A(n1989), .B(n1988), .Z(n144) );
  NAND U224 ( .A(n143), .B(n144), .Z(n2028) );
  NAND U225 ( .A(n2101), .B(n2102), .Z(n145) );
  NANDN U226 ( .A(n2100), .B(n2099), .Z(n146) );
  NAND U227 ( .A(n145), .B(n146), .Z(n2139) );
  NAND U228 ( .A(n2212), .B(n2213), .Z(n147) );
  NANDN U229 ( .A(n2211), .B(n2210), .Z(n148) );
  NAND U230 ( .A(n147), .B(n148), .Z(n2250) );
  NAND U231 ( .A(n2323), .B(n2324), .Z(n149) );
  NANDN U232 ( .A(n2322), .B(n2321), .Z(n150) );
  NAND U233 ( .A(n149), .B(n150), .Z(n2361) );
  NAND U234 ( .A(n2436), .B(n2437), .Z(n151) );
  NANDN U235 ( .A(n2435), .B(n2434), .Z(n152) );
  NAND U236 ( .A(n151), .B(n152), .Z(n2475) );
  NAND U237 ( .A(n287), .B(n286), .Z(n153) );
  XOR U238 ( .A(n286), .B(n287), .Z(n154) );
  NANDN U239 ( .A(n288), .B(n154), .Z(n155) );
  NAND U240 ( .A(n153), .B(n155), .Z(n300) );
  XNOR U241 ( .A(n2691), .B(n2692), .Z(n2687) );
  NANDN U242 ( .A(n248), .B(a[0]), .Z(n156) );
  ANDN U243 ( .B(n156), .A(n2695), .Z(n157) );
  XNOR U244 ( .A(a[0]), .B(n248), .Z(n158) );
  NAND U245 ( .A(n158), .B(b[6]), .Z(n159) );
  NAND U246 ( .A(n157), .B(n159), .Z(n400) );
  NAND U247 ( .A(n470), .B(n471), .Z(n160) );
  NANDN U248 ( .A(n469), .B(n468), .Z(n161) );
  NAND U249 ( .A(n160), .B(n161), .Z(n535) );
  NAND U250 ( .A(n583), .B(n584), .Z(n162) );
  NANDN U251 ( .A(n582), .B(n581), .Z(n163) );
  NAND U252 ( .A(n162), .B(n163), .Z(n643) );
  NAND U253 ( .A(n694), .B(n695), .Z(n164) );
  NANDN U254 ( .A(n693), .B(n692), .Z(n165) );
  NAND U255 ( .A(n164), .B(n165), .Z(n757) );
  NAND U256 ( .A(n807), .B(n808), .Z(n166) );
  NANDN U257 ( .A(n806), .B(n805), .Z(n167) );
  NAND U258 ( .A(n166), .B(n167), .Z(n867) );
  NAND U259 ( .A(n918), .B(n919), .Z(n168) );
  NANDN U260 ( .A(n917), .B(n916), .Z(n169) );
  NAND U261 ( .A(n168), .B(n169), .Z(n980) );
  NAND U262 ( .A(n1031), .B(n1032), .Z(n170) );
  NANDN U263 ( .A(n1030), .B(n1029), .Z(n171) );
  NAND U264 ( .A(n170), .B(n171), .Z(n1091) );
  NAND U265 ( .A(n1142), .B(n1143), .Z(n172) );
  NANDN U266 ( .A(n1141), .B(n1140), .Z(n173) );
  NAND U267 ( .A(n172), .B(n173), .Z(n1205) );
  NAND U268 ( .A(n1254), .B(n1255), .Z(n174) );
  NANDN U269 ( .A(n1253), .B(n1252), .Z(n175) );
  NAND U270 ( .A(n174), .B(n175), .Z(n1314) );
  NAND U271 ( .A(n1365), .B(n1366), .Z(n176) );
  NANDN U272 ( .A(n1364), .B(n1363), .Z(n177) );
  NAND U273 ( .A(n176), .B(n177), .Z(n1425) );
  NAND U274 ( .A(n1476), .B(n1477), .Z(n178) );
  NANDN U275 ( .A(n1475), .B(n1474), .Z(n179) );
  NAND U276 ( .A(n178), .B(n179), .Z(n1536) );
  NAND U277 ( .A(n1587), .B(n1588), .Z(n180) );
  NANDN U278 ( .A(n1586), .B(n1585), .Z(n181) );
  NAND U279 ( .A(n180), .B(n181), .Z(n1647) );
  NAND U280 ( .A(n1698), .B(n1699), .Z(n182) );
  NANDN U281 ( .A(n1697), .B(n1696), .Z(n183) );
  NAND U282 ( .A(n182), .B(n183), .Z(n1758) );
  NAND U283 ( .A(n1809), .B(n1810), .Z(n184) );
  NANDN U284 ( .A(n1808), .B(n1807), .Z(n185) );
  NAND U285 ( .A(n184), .B(n185), .Z(n1869) );
  NAND U286 ( .A(n1920), .B(n1921), .Z(n186) );
  NANDN U287 ( .A(n1919), .B(n1918), .Z(n187) );
  NAND U288 ( .A(n186), .B(n187), .Z(n1980) );
  NAND U289 ( .A(n2031), .B(n2032), .Z(n188) );
  NANDN U290 ( .A(n2030), .B(n2029), .Z(n189) );
  NAND U291 ( .A(n188), .B(n189), .Z(n2091) );
  NAND U292 ( .A(n2142), .B(n2143), .Z(n190) );
  NANDN U293 ( .A(n2141), .B(n2140), .Z(n191) );
  NAND U294 ( .A(n190), .B(n191), .Z(n2202) );
  NAND U295 ( .A(n2253), .B(n2254), .Z(n192) );
  NANDN U296 ( .A(n2252), .B(n2251), .Z(n193) );
  NAND U297 ( .A(n192), .B(n193), .Z(n2313) );
  NAND U298 ( .A(n2364), .B(n2365), .Z(n194) );
  NANDN U299 ( .A(n2363), .B(n2362), .Z(n195) );
  NAND U300 ( .A(n194), .B(n195), .Z(n2426) );
  NOR U301 ( .A(n336), .B(n337), .Z(n375) );
  NAND U302 ( .A(n2484), .B(n2485), .Z(n196) );
  NANDN U303 ( .A(n2483), .B(n2482), .Z(n197) );
  NAND U304 ( .A(n196), .B(n197), .Z(n2541) );
  XNOR U305 ( .A(n2524), .B(n2525), .Z(n2517) );
  ANDN U306 ( .B(n417), .A(n247), .Z(n198) );
  AND U307 ( .A(n2561), .B(n198), .Z(n199) );
  ANDN U308 ( .B(n2602), .A(n247), .Z(n200) );
  NAND U309 ( .A(n200), .B(n2537), .Z(n201) );
  NANDN U310 ( .A(n199), .B(n201), .Z(n286) );
  NAND U311 ( .A(n579), .B(n580), .Z(n202) );
  NANDN U312 ( .A(n578), .B(n577), .Z(n203) );
  NAND U313 ( .A(n202), .B(n203), .Z(n617) );
  NAND U314 ( .A(n690), .B(n691), .Z(n204) );
  NANDN U315 ( .A(n689), .B(n688), .Z(n205) );
  NAND U316 ( .A(n204), .B(n205), .Z(n729) );
  NAND U317 ( .A(n803), .B(n804), .Z(n206) );
  NANDN U318 ( .A(n802), .B(n801), .Z(n207) );
  NAND U319 ( .A(n206), .B(n207), .Z(n841) );
  NAND U320 ( .A(n914), .B(n915), .Z(n208) );
  NANDN U321 ( .A(n913), .B(n912), .Z(n209) );
  NAND U322 ( .A(n208), .B(n209), .Z(n952) );
  NAND U323 ( .A(n1027), .B(n1028), .Z(n210) );
  NANDN U324 ( .A(n1026), .B(n1025), .Z(n211) );
  NAND U325 ( .A(n210), .B(n211), .Z(n1065) );
  NAND U326 ( .A(n1138), .B(n1139), .Z(n212) );
  NANDN U327 ( .A(n1137), .B(n1136), .Z(n213) );
  NAND U328 ( .A(n212), .B(n213), .Z(n1177) );
  NAND U329 ( .A(n1250), .B(n1251), .Z(n214) );
  NANDN U330 ( .A(n1249), .B(n1248), .Z(n215) );
  NAND U331 ( .A(n214), .B(n215), .Z(n1288) );
  NAND U332 ( .A(n1361), .B(n1362), .Z(n216) );
  NANDN U333 ( .A(n1360), .B(n1359), .Z(n217) );
  NAND U334 ( .A(n216), .B(n217), .Z(n1399) );
  NAND U335 ( .A(n1472), .B(n1473), .Z(n218) );
  NANDN U336 ( .A(n1471), .B(n1470), .Z(n219) );
  NAND U337 ( .A(n218), .B(n219), .Z(n1510) );
  NAND U338 ( .A(n1583), .B(n1584), .Z(n220) );
  NANDN U339 ( .A(n1582), .B(n1581), .Z(n221) );
  NAND U340 ( .A(n220), .B(n221), .Z(n1621) );
  NAND U341 ( .A(n1694), .B(n1695), .Z(n222) );
  NANDN U342 ( .A(n1693), .B(n1692), .Z(n223) );
  NAND U343 ( .A(n222), .B(n223), .Z(n1732) );
  NAND U344 ( .A(n1805), .B(n1806), .Z(n224) );
  NANDN U345 ( .A(n1804), .B(n1803), .Z(n225) );
  NAND U346 ( .A(n224), .B(n225), .Z(n1843) );
  NAND U347 ( .A(n1916), .B(n1917), .Z(n226) );
  NANDN U348 ( .A(n1915), .B(n1914), .Z(n227) );
  NAND U349 ( .A(n226), .B(n227), .Z(n1954) );
  NAND U350 ( .A(n2027), .B(n2028), .Z(n228) );
  NANDN U351 ( .A(n2026), .B(n2025), .Z(n229) );
  NAND U352 ( .A(n228), .B(n229), .Z(n2065) );
  NAND U353 ( .A(n2138), .B(n2139), .Z(n230) );
  NANDN U354 ( .A(n2137), .B(n2136), .Z(n231) );
  NAND U355 ( .A(n230), .B(n231), .Z(n2176) );
  NAND U356 ( .A(n2249), .B(n2250), .Z(n232) );
  NANDN U357 ( .A(n2248), .B(n2247), .Z(n233) );
  NAND U358 ( .A(n232), .B(n233), .Z(n2287) );
  NAND U359 ( .A(n2360), .B(n2361), .Z(n234) );
  NANDN U360 ( .A(n2359), .B(n2358), .Z(n235) );
  NAND U361 ( .A(n234), .B(n235), .Z(n2399) );
  NAND U362 ( .A(n330), .B(n331), .Z(n236) );
  NANDN U363 ( .A(n329), .B(n328), .Z(n237) );
  NAND U364 ( .A(n236), .B(n237), .Z(n350) );
  NAND U365 ( .A(n2474), .B(n2475), .Z(n238) );
  NANDN U366 ( .A(n2473), .B(n2472), .Z(n239) );
  NAND U367 ( .A(n238), .B(n239), .Z(n2513) );
  NAND U368 ( .A(n2584), .B(n2582), .Z(n240) );
  XOR U369 ( .A(n2582), .B(n2584), .Z(n241) );
  NANDN U370 ( .A(n2583), .B(n241), .Z(n242) );
  NAND U371 ( .A(n240), .B(n242), .Z(n2615) );
  XOR U372 ( .A(n2688), .B(n2687), .Z(n243) );
  NANDN U373 ( .A(n2686), .B(n243), .Z(n244) );
  NAND U374 ( .A(n2688), .B(n2687), .Z(n245) );
  AND U375 ( .A(n244), .B(n245), .Z(n2702) );
  IV U376 ( .A(b[0]), .Z(n246) );
  IV U377 ( .A(b[3]), .Z(n247) );
  IV U378 ( .A(b[5]), .Z(n248) );
  NANDN U379 ( .A(n246), .B(a[0]), .Z(n250) );
  XNOR U380 ( .A(n250), .B(sreg[56]), .Z(c[56]) );
  ANDN U381 ( .B(a[1]), .A(n246), .Z(n254) );
  IV U382 ( .A(b[1]), .Z(n2537) );
  NANDN U383 ( .A(n2537), .B(a[0]), .Z(n249) );
  XNOR U384 ( .A(n254), .B(n249), .Z(n256) );
  XNOR U385 ( .A(sreg[57]), .B(n256), .Z(n258) );
  NANDN U386 ( .A(n250), .B(sreg[56]), .Z(n257) );
  XOR U387 ( .A(n258), .B(n257), .Z(c[57]) );
  NANDN U388 ( .A(n246), .B(a[2]), .Z(n251) );
  XOR U389 ( .A(n2537), .B(n251), .Z(n253) );
  NANDN U390 ( .A(b[0]), .B(a[1]), .Z(n252) );
  AND U391 ( .A(n253), .B(n252), .Z(n261) );
  IV U392 ( .A(a[0]), .Z(n417) );
  IV U393 ( .A(b[2]), .Z(n2602) );
  XOR U394 ( .A(n2602), .B(n2537), .Z(n2561) );
  NANDN U395 ( .A(n417), .B(n2561), .Z(n262) );
  XOR U396 ( .A(n261), .B(n262), .Z(n264) );
  ANDN U397 ( .B(n417), .A(n254), .Z(n255) );
  NANDN U398 ( .A(n2537), .B(n255), .Z(n263) );
  XOR U399 ( .A(n264), .B(n263), .Z(n277) );
  NAND U400 ( .A(sreg[57]), .B(n256), .Z(n260) );
  OR U401 ( .A(n258), .B(n257), .Z(n259) );
  NAND U402 ( .A(n260), .B(n259), .Z(n276) );
  XNOR U403 ( .A(n276), .B(sreg[58]), .Z(n278) );
  XNOR U404 ( .A(n277), .B(n278), .Z(c[58]) );
  NANDN U405 ( .A(n262), .B(n261), .Z(n266) );
  OR U406 ( .A(n264), .B(n263), .Z(n265) );
  AND U407 ( .A(n266), .B(n265), .Z(n288) );
  XNOR U408 ( .A(n247), .B(a[0]), .Z(n269) );
  XOR U409 ( .A(n247), .B(n2602), .Z(n268) );
  XNOR U410 ( .A(n247), .B(b[1]), .Z(n267) );
  AND U411 ( .A(n268), .B(n267), .Z(n2563) );
  NAND U412 ( .A(n269), .B(n2563), .Z(n271) );
  XNOR U413 ( .A(n247), .B(a[1]), .Z(n294) );
  NAND U414 ( .A(n294), .B(n2561), .Z(n270) );
  NAND U415 ( .A(n271), .B(n270), .Z(n290) );
  NANDN U416 ( .A(n246), .B(a[3]), .Z(n272) );
  XOR U417 ( .A(n2537), .B(n272), .Z(n274) );
  NANDN U418 ( .A(b[0]), .B(a[2]), .Z(n273) );
  NAND U419 ( .A(n274), .B(n273), .Z(n289) );
  XNOR U420 ( .A(n290), .B(n289), .Z(n287) );
  XOR U421 ( .A(n286), .B(n287), .Z(n275) );
  XNOR U422 ( .A(n288), .B(n275), .Z(n281) );
  XOR U423 ( .A(sreg[59]), .B(n281), .Z(n282) );
  NAND U424 ( .A(n276), .B(sreg[58]), .Z(n280) );
  NANDN U425 ( .A(n278), .B(n277), .Z(n279) );
  NAND U426 ( .A(n280), .B(n279), .Z(n283) );
  XOR U427 ( .A(n282), .B(n283), .Z(c[59]) );
  OR U428 ( .A(n281), .B(sreg[59]), .Z(n285) );
  NANDN U429 ( .A(n283), .B(n282), .Z(n284) );
  AND U430 ( .A(n285), .B(n284), .Z(n318) );
  XNOR U431 ( .A(sreg[60]), .B(n318), .Z(n320) );
  ANDN U432 ( .B(n290), .A(n289), .Z(n299) );
  NANDN U433 ( .A(n246), .B(a[4]), .Z(n291) );
  XOR U434 ( .A(n2537), .B(n291), .Z(n293) );
  IV U435 ( .A(a[3]), .Z(n358) );
  NANDN U436 ( .A(n358), .B(n246), .Z(n292) );
  AND U437 ( .A(n293), .B(n292), .Z(n312) );
  XNOR U438 ( .A(b[3]), .B(a[2]), .Z(n301) );
  NANDN U439 ( .A(n301), .B(n2561), .Z(n296) );
  NAND U440 ( .A(n294), .B(n2563), .Z(n295) );
  AND U441 ( .A(n296), .B(n295), .Z(n313) );
  XOR U442 ( .A(n312), .B(n313), .Z(n315) );
  XNOR U443 ( .A(b[4]), .B(b[3]), .Z(n2608) );
  NANDN U444 ( .A(n2608), .B(a[0]), .Z(n314) );
  XNOR U445 ( .A(n315), .B(n314), .Z(n298) );
  XNOR U446 ( .A(n299), .B(n298), .Z(n297) );
  XNOR U447 ( .A(n300), .B(n297), .Z(n319) );
  XOR U448 ( .A(n320), .B(n319), .Z(c[60]) );
  XOR U449 ( .A(b[3]), .B(n358), .Z(n338) );
  NANDN U450 ( .A(n338), .B(n2561), .Z(n303) );
  NANDN U451 ( .A(n301), .B(n2563), .Z(n302) );
  AND U452 ( .A(n303), .B(n302), .Z(n333) );
  IV U453 ( .A(b[4]), .Z(n2658) );
  ANDN U454 ( .B(b[5]), .A(n2608), .Z(n2628) );
  XNOR U455 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U456 ( .A(n248), .B(a[0]), .Z(n306) );
  XNOR U457 ( .A(n248), .B(b[4]), .Z(n305) );
  XNOR U458 ( .A(n248), .B(b[3]), .Z(n304) );
  AND U459 ( .A(n305), .B(n304), .Z(n2625) );
  NAND U460 ( .A(n306), .B(n2625), .Z(n308) );
  XNOR U461 ( .A(n248), .B(a[1]), .Z(n344) );
  ANDN U462 ( .B(n344), .A(n2608), .Z(n307) );
  ANDN U463 ( .B(n308), .A(n307), .Z(n337) );
  NANDN U464 ( .A(n246), .B(a[5]), .Z(n309) );
  XOR U465 ( .A(n2537), .B(n309), .Z(n311) );
  NANDN U466 ( .A(b[0]), .B(a[4]), .Z(n310) );
  NAND U467 ( .A(n311), .B(n310), .Z(n336) );
  XNOR U468 ( .A(n337), .B(n336), .Z(n335) );
  XOR U469 ( .A(n334), .B(n335), .Z(n328) );
  NANDN U470 ( .A(n313), .B(n312), .Z(n317) );
  OR U471 ( .A(n315), .B(n314), .Z(n316) );
  NAND U472 ( .A(n317), .B(n316), .Z(n329) );
  XNOR U473 ( .A(n328), .B(n329), .Z(n331) );
  XOR U474 ( .A(n330), .B(n331), .Z(n323) );
  XOR U475 ( .A(n323), .B(sreg[61]), .Z(n325) );
  NAND U476 ( .A(n318), .B(sreg[60]), .Z(n322) );
  OR U477 ( .A(n320), .B(n319), .Z(n321) );
  AND U478 ( .A(n322), .B(n321), .Z(n324) );
  XOR U479 ( .A(n325), .B(n324), .Z(c[61]) );
  NANDN U480 ( .A(n323), .B(sreg[61]), .Z(n327) );
  OR U481 ( .A(n325), .B(n324), .Z(n326) );
  NAND U482 ( .A(n327), .B(n326), .Z(n378) );
  XNOR U483 ( .A(n378), .B(sreg[62]), .Z(n380) );
  XNOR U484 ( .A(n247), .B(a[4]), .Z(n369) );
  NAND U485 ( .A(n369), .B(n2561), .Z(n340) );
  NANDN U486 ( .A(n338), .B(n2563), .Z(n339) );
  NAND U487 ( .A(n340), .B(n339), .Z(n356) );
  NANDN U488 ( .A(n246), .B(a[6]), .Z(n341) );
  XOR U489 ( .A(n2537), .B(n341), .Z(n343) );
  NANDN U490 ( .A(b[0]), .B(a[5]), .Z(n342) );
  AND U491 ( .A(n343), .B(n342), .Z(n353) );
  XNOR U492 ( .A(n248), .B(b[6]), .Z(n2665) );
  NANDN U493 ( .A(n417), .B(n2665), .Z(n354) );
  XNOR U494 ( .A(n353), .B(n354), .Z(n355) );
  XNOR U495 ( .A(n356), .B(n355), .Z(n372) );
  XNOR U496 ( .A(b[5]), .B(a[2]), .Z(n357) );
  OR U497 ( .A(n357), .B(n2608), .Z(n346) );
  NAND U498 ( .A(n2625), .B(n344), .Z(n345) );
  NAND U499 ( .A(n346), .B(n345), .Z(n373) );
  XNOR U500 ( .A(n372), .B(n373), .Z(n374) );
  XOR U501 ( .A(n375), .B(n374), .Z(n348) );
  XOR U502 ( .A(n347), .B(n348), .Z(n349) );
  XOR U503 ( .A(n350), .B(n349), .Z(n379) );
  XOR U504 ( .A(n380), .B(n379), .Z(c[62]) );
  OR U505 ( .A(n348), .B(n347), .Z(n352) );
  NAND U506 ( .A(n350), .B(n349), .Z(n351) );
  NAND U507 ( .A(n352), .B(n351), .Z(n391) );
  NANDN U508 ( .A(n357), .B(n2625), .Z(n360) );
  XOR U509 ( .A(n248), .B(n358), .Z(n418) );
  NANDN U510 ( .A(n2608), .B(n418), .Z(n359) );
  NAND U511 ( .A(n360), .B(n359), .Z(n407) );
  IV U512 ( .A(b[7]), .Z(n2695) );
  XNOR U513 ( .A(n2695), .B(a[0]), .Z(n363) );
  XNOR U514 ( .A(n2695), .B(b[5]), .Z(n362) );
  XNOR U515 ( .A(n2695), .B(b[6]), .Z(n361) );
  AND U516 ( .A(n362), .B(n361), .Z(n2666) );
  NAND U517 ( .A(n363), .B(n2666), .Z(n365) );
  XNOR U518 ( .A(n2695), .B(a[1]), .Z(n408) );
  NAND U519 ( .A(n408), .B(n2665), .Z(n364) );
  NAND U520 ( .A(n365), .B(n364), .Z(n406) );
  XNOR U521 ( .A(n407), .B(n406), .Z(n403) );
  NANDN U522 ( .A(n246), .B(a[7]), .Z(n366) );
  XOR U523 ( .A(n2537), .B(n366), .Z(n368) );
  NANDN U524 ( .A(b[0]), .B(a[6]), .Z(n367) );
  AND U525 ( .A(n368), .B(n367), .Z(n401) );
  XNOR U526 ( .A(n400), .B(n401), .Z(n402) );
  XOR U527 ( .A(n403), .B(n402), .Z(n394) );
  XOR U528 ( .A(n247), .B(a[5]), .Z(n411) );
  NANDN U529 ( .A(n411), .B(n2561), .Z(n371) );
  NAND U530 ( .A(n2563), .B(n369), .Z(n370) );
  AND U531 ( .A(n371), .B(n370), .Z(n395) );
  XNOR U532 ( .A(n394), .B(n395), .Z(n396) );
  XNOR U533 ( .A(n397), .B(n396), .Z(n388) );
  NANDN U534 ( .A(n373), .B(n372), .Z(n377) );
  NANDN U535 ( .A(n375), .B(n374), .Z(n376) );
  NAND U536 ( .A(n377), .B(n376), .Z(n389) );
  XNOR U537 ( .A(n388), .B(n389), .Z(n390) );
  XNOR U538 ( .A(n391), .B(n390), .Z(n383) );
  XNOR U539 ( .A(sreg[63]), .B(n383), .Z(n385) );
  NAND U540 ( .A(n378), .B(sreg[62]), .Z(n382) );
  OR U541 ( .A(n380), .B(n379), .Z(n381) );
  AND U542 ( .A(n382), .B(n381), .Z(n384) );
  XOR U543 ( .A(n385), .B(n384), .Z(c[63]) );
  NAND U544 ( .A(sreg[63]), .B(n383), .Z(n387) );
  OR U545 ( .A(n385), .B(n384), .Z(n386) );
  NAND U546 ( .A(n387), .B(n386), .Z(n457) );
  XNOR U547 ( .A(n457), .B(sreg[64]), .Z(n459) );
  NANDN U548 ( .A(n389), .B(n388), .Z(n393) );
  NANDN U549 ( .A(n391), .B(n390), .Z(n392) );
  NAND U550 ( .A(n393), .B(n392), .Z(n454) );
  NAND U551 ( .A(n395), .B(n394), .Z(n399) );
  OR U552 ( .A(n397), .B(n396), .Z(n398) );
  NAND U553 ( .A(n399), .B(n398), .Z(n452) );
  NANDN U554 ( .A(n401), .B(n400), .Z(n405) );
  NAND U555 ( .A(n403), .B(n402), .Z(n404) );
  NAND U556 ( .A(n405), .B(n404), .Z(n445) );
  NAND U557 ( .A(n407), .B(n406), .Z(n442) );
  NAND U558 ( .A(n408), .B(n2666), .Z(n410) );
  XNOR U559 ( .A(n2695), .B(a[2]), .Z(n421) );
  NAND U560 ( .A(n421), .B(n2665), .Z(n409) );
  NAND U561 ( .A(n410), .B(n409), .Z(n440) );
  XNOR U562 ( .A(b[3]), .B(a[6]), .Z(n424) );
  NANDN U563 ( .A(n424), .B(n2561), .Z(n413) );
  NANDN U564 ( .A(n411), .B(n2563), .Z(n412) );
  AND U565 ( .A(n413), .B(n412), .Z(n439) );
  XNOR U566 ( .A(n440), .B(n439), .Z(n441) );
  XNOR U567 ( .A(n442), .B(n441), .Z(n446) );
  XNOR U568 ( .A(n445), .B(n446), .Z(n447) );
  NANDN U569 ( .A(n246), .B(a[8]), .Z(n414) );
  XOR U570 ( .A(n2537), .B(n414), .Z(n416) );
  NANDN U571 ( .A(b[0]), .B(a[7]), .Z(n415) );
  AND U572 ( .A(n416), .B(n415), .Z(n436) );
  ANDN U573 ( .B(b[7]), .A(n417), .Z(n433) );
  XNOR U574 ( .A(b[5]), .B(a[4]), .Z(n430) );
  OR U575 ( .A(n430), .B(n2608), .Z(n420) );
  NAND U576 ( .A(n2625), .B(n418), .Z(n419) );
  NAND U577 ( .A(n420), .B(n419), .Z(n434) );
  XOR U578 ( .A(n433), .B(n434), .Z(n435) );
  XOR U579 ( .A(n436), .B(n435), .Z(n448) );
  XNOR U580 ( .A(n447), .B(n448), .Z(n451) );
  XNOR U581 ( .A(n452), .B(n451), .Z(n453) );
  XOR U582 ( .A(n454), .B(n453), .Z(n458) );
  XOR U583 ( .A(n459), .B(n458), .Z(c[64]) );
  NAND U584 ( .A(n421), .B(n2666), .Z(n423) );
  XNOR U585 ( .A(n2695), .B(a[3]), .Z(n484) );
  NAND U586 ( .A(n484), .B(n2665), .Z(n422) );
  NAND U587 ( .A(n423), .B(n422), .Z(n468) );
  XNOR U588 ( .A(b[3]), .B(a[7]), .Z(n487) );
  NANDN U589 ( .A(n487), .B(n2561), .Z(n426) );
  NANDN U590 ( .A(n424), .B(n2563), .Z(n425) );
  AND U591 ( .A(n426), .B(n425), .Z(n469) );
  XNOR U592 ( .A(n468), .B(n469), .Z(n470) );
  NANDN U593 ( .A(n246), .B(a[9]), .Z(n427) );
  XOR U594 ( .A(n2537), .B(n427), .Z(n429) );
  IV U595 ( .A(a[8]), .Z(n702) );
  NANDN U596 ( .A(n702), .B(n246), .Z(n428) );
  AND U597 ( .A(n429), .B(n428), .Z(n474) );
  NANDN U598 ( .A(n430), .B(n2625), .Z(n432) );
  XNOR U599 ( .A(b[5]), .B(a[5]), .Z(n481) );
  OR U600 ( .A(n481), .B(n2608), .Z(n431) );
  NAND U601 ( .A(n432), .B(n431), .Z(n472) );
  NANDN U602 ( .A(n2695), .B(a[1]), .Z(n473) );
  XNOR U603 ( .A(n472), .B(n473), .Z(n475) );
  XOR U604 ( .A(n474), .B(n475), .Z(n471) );
  XOR U605 ( .A(n470), .B(n471), .Z(n490) );
  OR U606 ( .A(n434), .B(n433), .Z(n438) );
  NANDN U607 ( .A(n436), .B(n435), .Z(n437) );
  AND U608 ( .A(n438), .B(n437), .Z(n491) );
  XNOR U609 ( .A(n490), .B(n491), .Z(n493) );
  NANDN U610 ( .A(n440), .B(n439), .Z(n444) );
  NAND U611 ( .A(n442), .B(n441), .Z(n443) );
  AND U612 ( .A(n444), .B(n443), .Z(n492) );
  XNOR U613 ( .A(n493), .B(n492), .Z(n462) );
  NANDN U614 ( .A(n446), .B(n445), .Z(n450) );
  NANDN U615 ( .A(n448), .B(n447), .Z(n449) );
  AND U616 ( .A(n450), .B(n449), .Z(n463) );
  XNOR U617 ( .A(n462), .B(n463), .Z(n465) );
  NAND U618 ( .A(n452), .B(n451), .Z(n456) );
  OR U619 ( .A(n454), .B(n453), .Z(n455) );
  AND U620 ( .A(n456), .B(n455), .Z(n464) );
  XNOR U621 ( .A(n465), .B(n464), .Z(n496) );
  XNOR U622 ( .A(sreg[65]), .B(n496), .Z(n498) );
  NAND U623 ( .A(n457), .B(sreg[64]), .Z(n461) );
  OR U624 ( .A(n459), .B(n458), .Z(n460) );
  AND U625 ( .A(n461), .B(n460), .Z(n497) );
  XOR U626 ( .A(n498), .B(n497), .Z(c[65]) );
  NAND U627 ( .A(n463), .B(n462), .Z(n467) );
  NANDN U628 ( .A(n465), .B(n464), .Z(n466) );
  NAND U629 ( .A(n467), .B(n466), .Z(n503) );
  NANDN U630 ( .A(n473), .B(n472), .Z(n477) );
  NAND U631 ( .A(n475), .B(n474), .Z(n476) );
  NAND U632 ( .A(n477), .B(n476), .Z(n533) );
  NANDN U633 ( .A(n246), .B(a[10]), .Z(n478) );
  XOR U634 ( .A(n2537), .B(n478), .Z(n480) );
  NANDN U635 ( .A(b[0]), .B(a[9]), .Z(n479) );
  AND U636 ( .A(n480), .B(n479), .Z(n515) );
  NANDN U637 ( .A(n481), .B(n2625), .Z(n483) );
  XNOR U638 ( .A(n248), .B(a[6]), .Z(n522) );
  NANDN U639 ( .A(n2608), .B(n522), .Z(n482) );
  NAND U640 ( .A(n483), .B(n482), .Z(n513) );
  NANDN U641 ( .A(n2695), .B(a[2]), .Z(n514) );
  XNOR U642 ( .A(n513), .B(n514), .Z(n516) );
  XOR U643 ( .A(n515), .B(n516), .Z(n509) );
  NAND U644 ( .A(n484), .B(n2666), .Z(n486) );
  XNOR U645 ( .A(n2695), .B(a[4]), .Z(n526) );
  NAND U646 ( .A(n526), .B(n2665), .Z(n485) );
  NAND U647 ( .A(n486), .B(n485), .Z(n507) );
  XOR U648 ( .A(b[3]), .B(n702), .Z(n529) );
  NANDN U649 ( .A(n529), .B(n2561), .Z(n489) );
  NANDN U650 ( .A(n487), .B(n2563), .Z(n488) );
  AND U651 ( .A(n489), .B(n488), .Z(n508) );
  XOR U652 ( .A(n507), .B(n508), .Z(n510) );
  XNOR U653 ( .A(n509), .B(n510), .Z(n532) );
  XOR U654 ( .A(n533), .B(n532), .Z(n534) );
  XNOR U655 ( .A(n535), .B(n534), .Z(n501) );
  NAND U656 ( .A(n491), .B(n490), .Z(n495) );
  NANDN U657 ( .A(n493), .B(n492), .Z(n494) );
  NAND U658 ( .A(n495), .B(n494), .Z(n502) );
  XOR U659 ( .A(n501), .B(n502), .Z(n504) );
  XNOR U660 ( .A(n503), .B(n504), .Z(n538) );
  XNOR U661 ( .A(n538), .B(sreg[66]), .Z(n540) );
  NAND U662 ( .A(sreg[65]), .B(n496), .Z(n500) );
  OR U663 ( .A(n498), .B(n497), .Z(n499) );
  AND U664 ( .A(n500), .B(n499), .Z(n539) );
  XOR U665 ( .A(n540), .B(n539), .Z(c[66]) );
  NANDN U666 ( .A(n502), .B(n501), .Z(n506) );
  OR U667 ( .A(n504), .B(n503), .Z(n505) );
  NAND U668 ( .A(n506), .B(n505), .Z(n546) );
  NANDN U669 ( .A(n508), .B(n507), .Z(n512) );
  NANDN U670 ( .A(n510), .B(n509), .Z(n511) );
  NAND U671 ( .A(n512), .B(n511), .Z(n569) );
  NANDN U672 ( .A(n514), .B(n513), .Z(n518) );
  NAND U673 ( .A(n516), .B(n515), .Z(n517) );
  NAND U674 ( .A(n518), .B(n517), .Z(n567) );
  NANDN U675 ( .A(n246), .B(a[11]), .Z(n519) );
  XOR U676 ( .A(n2537), .B(n519), .Z(n521) );
  NANDN U677 ( .A(b[0]), .B(a[10]), .Z(n520) );
  AND U678 ( .A(n521), .B(n520), .Z(n553) );
  XNOR U679 ( .A(b[5]), .B(a[7]), .Z(n563) );
  OR U680 ( .A(n563), .B(n2608), .Z(n524) );
  NAND U681 ( .A(n2625), .B(n522), .Z(n523) );
  AND U682 ( .A(n524), .B(n523), .Z(n552) );
  AND U683 ( .A(a[3]), .B(b[7]), .Z(n551) );
  XNOR U684 ( .A(n552), .B(n551), .Z(n525) );
  XOR U685 ( .A(n553), .B(n525), .Z(n550) );
  NAND U686 ( .A(n526), .B(n2666), .Z(n528) );
  XNOR U687 ( .A(n2695), .B(a[5]), .Z(n554) );
  NAND U688 ( .A(n554), .B(n2665), .Z(n527) );
  NAND U689 ( .A(n528), .B(n527), .Z(n547) );
  XNOR U690 ( .A(b[3]), .B(a[9]), .Z(n557) );
  NANDN U691 ( .A(n557), .B(n2561), .Z(n531) );
  NANDN U692 ( .A(n529), .B(n2563), .Z(n530) );
  AND U693 ( .A(n531), .B(n530), .Z(n548) );
  XNOR U694 ( .A(n547), .B(n548), .Z(n549) );
  XOR U695 ( .A(n550), .B(n549), .Z(n566) );
  XOR U696 ( .A(n567), .B(n566), .Z(n568) );
  XNOR U697 ( .A(n569), .B(n568), .Z(n543) );
  NAND U698 ( .A(n533), .B(n532), .Z(n537) );
  NAND U699 ( .A(n535), .B(n534), .Z(n536) );
  NAND U700 ( .A(n537), .B(n536), .Z(n544) );
  XNOR U701 ( .A(n543), .B(n544), .Z(n545) );
  XNOR U702 ( .A(n546), .B(n545), .Z(n572) );
  XNOR U703 ( .A(n572), .B(sreg[67]), .Z(n574) );
  NAND U704 ( .A(n538), .B(sreg[66]), .Z(n542) );
  OR U705 ( .A(n540), .B(n539), .Z(n541) );
  AND U706 ( .A(n542), .B(n541), .Z(n573) );
  XOR U707 ( .A(n574), .B(n573), .Z(c[67]) );
  NAND U708 ( .A(n554), .B(n2666), .Z(n556) );
  XNOR U709 ( .A(n2695), .B(a[6]), .Z(n591) );
  NAND U710 ( .A(n591), .B(n2665), .Z(n555) );
  NAND U711 ( .A(n556), .B(n555), .Z(n581) );
  XNOR U712 ( .A(b[3]), .B(a[10]), .Z(n594) );
  NANDN U713 ( .A(n594), .B(n2561), .Z(n559) );
  NANDN U714 ( .A(n557), .B(n2563), .Z(n558) );
  AND U715 ( .A(n559), .B(n558), .Z(n582) );
  XNOR U716 ( .A(n581), .B(n582), .Z(n583) );
  NANDN U717 ( .A(n246), .B(a[12]), .Z(n560) );
  XOR U718 ( .A(n2537), .B(n560), .Z(n562) );
  NANDN U719 ( .A(b[0]), .B(a[11]), .Z(n561) );
  AND U720 ( .A(n562), .B(n561), .Z(n587) );
  NANDN U721 ( .A(n563), .B(n2625), .Z(n565) );
  XOR U722 ( .A(b[5]), .B(n702), .Z(n600) );
  OR U723 ( .A(n600), .B(n2608), .Z(n564) );
  NAND U724 ( .A(n565), .B(n564), .Z(n585) );
  NANDN U725 ( .A(n2695), .B(a[4]), .Z(n586) );
  XNOR U726 ( .A(n585), .B(n586), .Z(n588) );
  XOR U727 ( .A(n587), .B(n588), .Z(n584) );
  XOR U728 ( .A(n583), .B(n584), .Z(n604) );
  XOR U729 ( .A(n603), .B(n604), .Z(n605) );
  XNOR U730 ( .A(n606), .B(n605), .Z(n577) );
  NAND U731 ( .A(n567), .B(n566), .Z(n571) );
  NAND U732 ( .A(n569), .B(n568), .Z(n570) );
  NAND U733 ( .A(n571), .B(n570), .Z(n578) );
  XNOR U734 ( .A(n577), .B(n578), .Z(n579) );
  XNOR U735 ( .A(n580), .B(n579), .Z(n609) );
  XNOR U736 ( .A(n609), .B(sreg[68]), .Z(n611) );
  NAND U737 ( .A(n572), .B(sreg[67]), .Z(n576) );
  OR U738 ( .A(n574), .B(n573), .Z(n575) );
  AND U739 ( .A(n576), .B(n575), .Z(n610) );
  XOR U740 ( .A(n611), .B(n610), .Z(c[68]) );
  NANDN U741 ( .A(n586), .B(n585), .Z(n590) );
  NAND U742 ( .A(n588), .B(n587), .Z(n589) );
  NAND U743 ( .A(n590), .B(n589), .Z(n641) );
  NAND U744 ( .A(n591), .B(n2666), .Z(n593) );
  XNOR U745 ( .A(n2695), .B(a[7]), .Z(n628) );
  NAND U746 ( .A(n628), .B(n2665), .Z(n592) );
  NAND U747 ( .A(n593), .B(n592), .Z(n618) );
  XNOR U748 ( .A(b[3]), .B(a[11]), .Z(n631) );
  NANDN U749 ( .A(n631), .B(n2561), .Z(n596) );
  NANDN U750 ( .A(n594), .B(n2563), .Z(n595) );
  AND U751 ( .A(n596), .B(n595), .Z(n619) );
  XNOR U752 ( .A(n618), .B(n619), .Z(n620) );
  NANDN U753 ( .A(n246), .B(a[13]), .Z(n597) );
  XOR U754 ( .A(n2537), .B(n597), .Z(n599) );
  NANDN U755 ( .A(b[0]), .B(a[12]), .Z(n598) );
  AND U756 ( .A(n599), .B(n598), .Z(n624) );
  NANDN U757 ( .A(n600), .B(n2625), .Z(n602) );
  XNOR U758 ( .A(b[5]), .B(a[9]), .Z(n637) );
  OR U759 ( .A(n637), .B(n2608), .Z(n601) );
  NAND U760 ( .A(n602), .B(n601), .Z(n622) );
  NANDN U761 ( .A(n2695), .B(a[5]), .Z(n623) );
  XNOR U762 ( .A(n622), .B(n623), .Z(n625) );
  XOR U763 ( .A(n624), .B(n625), .Z(n621) );
  XOR U764 ( .A(n620), .B(n621), .Z(n640) );
  XOR U765 ( .A(n641), .B(n640), .Z(n642) );
  XNOR U766 ( .A(n643), .B(n642), .Z(n614) );
  NAND U767 ( .A(n604), .B(n603), .Z(n608) );
  NAND U768 ( .A(n606), .B(n605), .Z(n607) );
  NAND U769 ( .A(n608), .B(n607), .Z(n615) );
  XNOR U770 ( .A(n614), .B(n615), .Z(n616) );
  XNOR U771 ( .A(n617), .B(n616), .Z(n646) );
  XNOR U772 ( .A(n646), .B(sreg[69]), .Z(n648) );
  NAND U773 ( .A(n609), .B(sreg[68]), .Z(n613) );
  OR U774 ( .A(n611), .B(n610), .Z(n612) );
  AND U775 ( .A(n613), .B(n612), .Z(n647) );
  XOR U776 ( .A(n648), .B(n647), .Z(c[69]) );
  NANDN U777 ( .A(n623), .B(n622), .Z(n627) );
  NAND U778 ( .A(n625), .B(n624), .Z(n626) );
  NAND U779 ( .A(n627), .B(n626), .Z(n678) );
  NAND U780 ( .A(n628), .B(n2666), .Z(n630) );
  XNOR U781 ( .A(n2695), .B(a[8]), .Z(n665) );
  NAND U782 ( .A(n665), .B(n2665), .Z(n629) );
  NAND U783 ( .A(n630), .B(n629), .Z(n655) );
  XNOR U784 ( .A(b[3]), .B(a[12]), .Z(n668) );
  NANDN U785 ( .A(n668), .B(n2561), .Z(n633) );
  NANDN U786 ( .A(n631), .B(n2563), .Z(n632) );
  AND U787 ( .A(n633), .B(n632), .Z(n656) );
  XNOR U788 ( .A(n655), .B(n656), .Z(n657) );
  NANDN U789 ( .A(n246), .B(a[14]), .Z(n634) );
  XOR U790 ( .A(n2537), .B(n634), .Z(n636) );
  NANDN U791 ( .A(b[0]), .B(a[13]), .Z(n635) );
  AND U792 ( .A(n636), .B(n635), .Z(n661) );
  NANDN U793 ( .A(n637), .B(n2625), .Z(n639) );
  XNOR U794 ( .A(b[5]), .B(a[10]), .Z(n674) );
  OR U795 ( .A(n674), .B(n2608), .Z(n638) );
  NAND U796 ( .A(n639), .B(n638), .Z(n659) );
  NANDN U797 ( .A(n2695), .B(a[6]), .Z(n660) );
  XNOR U798 ( .A(n659), .B(n660), .Z(n662) );
  XOR U799 ( .A(n661), .B(n662), .Z(n658) );
  XOR U800 ( .A(n657), .B(n658), .Z(n677) );
  XOR U801 ( .A(n678), .B(n677), .Z(n679) );
  XNOR U802 ( .A(n680), .B(n679), .Z(n651) );
  NAND U803 ( .A(n641), .B(n640), .Z(n645) );
  NAND U804 ( .A(n643), .B(n642), .Z(n644) );
  NAND U805 ( .A(n645), .B(n644), .Z(n652) );
  XNOR U806 ( .A(n651), .B(n652), .Z(n653) );
  XNOR U807 ( .A(n654), .B(n653), .Z(n683) );
  XNOR U808 ( .A(n683), .B(sreg[70]), .Z(n685) );
  NAND U809 ( .A(n646), .B(sreg[69]), .Z(n650) );
  OR U810 ( .A(n648), .B(n647), .Z(n649) );
  AND U811 ( .A(n650), .B(n649), .Z(n684) );
  XOR U812 ( .A(n685), .B(n684), .Z(c[70]) );
  NANDN U813 ( .A(n660), .B(n659), .Z(n664) );
  NAND U814 ( .A(n662), .B(n661), .Z(n663) );
  NAND U815 ( .A(n664), .B(n663), .Z(n716) );
  NAND U816 ( .A(n665), .B(n2666), .Z(n667) );
  XNOR U817 ( .A(n2695), .B(a[9]), .Z(n709) );
  NAND U818 ( .A(n709), .B(n2665), .Z(n666) );
  NAND U819 ( .A(n667), .B(n666), .Z(n692) );
  XNOR U820 ( .A(b[3]), .B(a[13]), .Z(n712) );
  NANDN U821 ( .A(n712), .B(n2561), .Z(n670) );
  NANDN U822 ( .A(n668), .B(n2563), .Z(n669) );
  AND U823 ( .A(n670), .B(n669), .Z(n693) );
  XNOR U824 ( .A(n692), .B(n693), .Z(n694) );
  NANDN U825 ( .A(n246), .B(a[15]), .Z(n671) );
  XOR U826 ( .A(n2537), .B(n671), .Z(n673) );
  IV U827 ( .A(a[14]), .Z(n789) );
  NANDN U828 ( .A(n789), .B(n246), .Z(n672) );
  AND U829 ( .A(n673), .B(n672), .Z(n698) );
  NANDN U830 ( .A(n674), .B(n2625), .Z(n676) );
  XNOR U831 ( .A(n248), .B(a[11]), .Z(n703) );
  NANDN U832 ( .A(n2608), .B(n703), .Z(n675) );
  NAND U833 ( .A(n676), .B(n675), .Z(n696) );
  NANDN U834 ( .A(n2695), .B(a[7]), .Z(n697) );
  XNOR U835 ( .A(n696), .B(n697), .Z(n699) );
  XOR U836 ( .A(n698), .B(n699), .Z(n695) );
  XOR U837 ( .A(n694), .B(n695), .Z(n715) );
  XOR U838 ( .A(n716), .B(n715), .Z(n717) );
  XNOR U839 ( .A(n718), .B(n717), .Z(n688) );
  NAND U840 ( .A(n678), .B(n677), .Z(n682) );
  NAND U841 ( .A(n680), .B(n679), .Z(n681) );
  NAND U842 ( .A(n682), .B(n681), .Z(n689) );
  XNOR U843 ( .A(n688), .B(n689), .Z(n690) );
  XNOR U844 ( .A(n691), .B(n690), .Z(n721) );
  XNOR U845 ( .A(n721), .B(sreg[71]), .Z(n723) );
  NAND U846 ( .A(n683), .B(sreg[70]), .Z(n687) );
  OR U847 ( .A(n685), .B(n684), .Z(n686) );
  AND U848 ( .A(n687), .B(n686), .Z(n722) );
  XOR U849 ( .A(n723), .B(n722), .Z(c[71]) );
  NANDN U850 ( .A(n697), .B(n696), .Z(n701) );
  NAND U851 ( .A(n699), .B(n698), .Z(n700) );
  NAND U852 ( .A(n701), .B(n700), .Z(n754) );
  ANDN U853 ( .B(b[7]), .A(n702), .Z(n736) );
  XNOR U854 ( .A(b[5]), .B(a[12]), .Z(n751) );
  OR U855 ( .A(n751), .B(n2608), .Z(n705) );
  NAND U856 ( .A(n2625), .B(n703), .Z(n704) );
  NAND U857 ( .A(n705), .B(n704), .Z(n737) );
  XOR U858 ( .A(n736), .B(n737), .Z(n738) );
  NANDN U859 ( .A(n246), .B(a[16]), .Z(n706) );
  XOR U860 ( .A(n2537), .B(n706), .Z(n708) );
  NANDN U861 ( .A(b[0]), .B(a[15]), .Z(n707) );
  AND U862 ( .A(n708), .B(n707), .Z(n739) );
  XOR U863 ( .A(n738), .B(n739), .Z(n733) );
  NAND U864 ( .A(n709), .B(n2666), .Z(n711) );
  XNOR U865 ( .A(n2695), .B(a[10]), .Z(n742) );
  NAND U866 ( .A(n742), .B(n2665), .Z(n710) );
  NAND U867 ( .A(n711), .B(n710), .Z(n730) );
  XOR U868 ( .A(b[3]), .B(n789), .Z(n745) );
  NANDN U869 ( .A(n745), .B(n2561), .Z(n714) );
  NANDN U870 ( .A(n712), .B(n2563), .Z(n713) );
  AND U871 ( .A(n714), .B(n713), .Z(n731) );
  XNOR U872 ( .A(n730), .B(n731), .Z(n732) );
  XNOR U873 ( .A(n733), .B(n732), .Z(n755) );
  XNOR U874 ( .A(n754), .B(n755), .Z(n756) );
  XNOR U875 ( .A(n757), .B(n756), .Z(n726) );
  NAND U876 ( .A(n716), .B(n715), .Z(n720) );
  NAND U877 ( .A(n718), .B(n717), .Z(n719) );
  NAND U878 ( .A(n720), .B(n719), .Z(n727) );
  XNOR U879 ( .A(n726), .B(n727), .Z(n728) );
  XNOR U880 ( .A(n729), .B(n728), .Z(n760) );
  XNOR U881 ( .A(n760), .B(sreg[72]), .Z(n762) );
  NAND U882 ( .A(n721), .B(sreg[71]), .Z(n725) );
  OR U883 ( .A(n723), .B(n722), .Z(n724) );
  AND U884 ( .A(n725), .B(n724), .Z(n761) );
  XOR U885 ( .A(n762), .B(n761), .Z(c[72]) );
  NANDN U886 ( .A(n731), .B(n730), .Z(n735) );
  NAND U887 ( .A(n733), .B(n732), .Z(n734) );
  NAND U888 ( .A(n735), .B(n734), .Z(n795) );
  OR U889 ( .A(n737), .B(n736), .Z(n741) );
  NANDN U890 ( .A(n739), .B(n738), .Z(n740) );
  NAND U891 ( .A(n741), .B(n740), .Z(n793) );
  NAND U892 ( .A(n742), .B(n2666), .Z(n744) );
  XNOR U893 ( .A(n2695), .B(a[11]), .Z(n779) );
  NAND U894 ( .A(n779), .B(n2665), .Z(n743) );
  NAND U895 ( .A(n744), .B(n743), .Z(n769) );
  XNOR U896 ( .A(b[3]), .B(a[15]), .Z(n782) );
  NANDN U897 ( .A(n782), .B(n2561), .Z(n747) );
  NANDN U898 ( .A(n745), .B(n2563), .Z(n746) );
  AND U899 ( .A(n747), .B(n746), .Z(n770) );
  XNOR U900 ( .A(n769), .B(n770), .Z(n771) );
  NANDN U901 ( .A(n246), .B(a[17]), .Z(n748) );
  XOR U902 ( .A(n2537), .B(n748), .Z(n750) );
  NANDN U903 ( .A(b[0]), .B(a[16]), .Z(n749) );
  AND U904 ( .A(n750), .B(n749), .Z(n775) );
  NANDN U905 ( .A(n751), .B(n2625), .Z(n753) );
  XNOR U906 ( .A(b[5]), .B(a[13]), .Z(n788) );
  OR U907 ( .A(n788), .B(n2608), .Z(n752) );
  NAND U908 ( .A(n753), .B(n752), .Z(n773) );
  NANDN U909 ( .A(n2695), .B(a[9]), .Z(n774) );
  XNOR U910 ( .A(n773), .B(n774), .Z(n776) );
  XOR U911 ( .A(n775), .B(n776), .Z(n772) );
  XOR U912 ( .A(n771), .B(n772), .Z(n792) );
  XNOR U913 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U914 ( .A(n795), .B(n794), .Z(n765) );
  NANDN U915 ( .A(n755), .B(n754), .Z(n759) );
  NAND U916 ( .A(n757), .B(n756), .Z(n758) );
  NAND U917 ( .A(n759), .B(n758), .Z(n766) );
  XNOR U918 ( .A(n765), .B(n766), .Z(n767) );
  XNOR U919 ( .A(n768), .B(n767), .Z(n796) );
  XNOR U920 ( .A(n796), .B(sreg[73]), .Z(n798) );
  NAND U921 ( .A(n760), .B(sreg[72]), .Z(n764) );
  OR U922 ( .A(n762), .B(n761), .Z(n763) );
  AND U923 ( .A(n764), .B(n763), .Z(n797) );
  XOR U924 ( .A(n798), .B(n797), .Z(c[73]) );
  NANDN U925 ( .A(n774), .B(n773), .Z(n778) );
  NAND U926 ( .A(n776), .B(n775), .Z(n777) );
  NAND U927 ( .A(n778), .B(n777), .Z(n828) );
  NAND U928 ( .A(n779), .B(n2666), .Z(n781) );
  XNOR U929 ( .A(n2695), .B(a[12]), .Z(n815) );
  NAND U930 ( .A(n815), .B(n2665), .Z(n780) );
  NAND U931 ( .A(n781), .B(n780), .Z(n805) );
  XNOR U932 ( .A(b[3]), .B(a[16]), .Z(n818) );
  NANDN U933 ( .A(n818), .B(n2561), .Z(n784) );
  NANDN U934 ( .A(n782), .B(n2563), .Z(n783) );
  AND U935 ( .A(n784), .B(n783), .Z(n806) );
  XNOR U936 ( .A(n805), .B(n806), .Z(n807) );
  NANDN U937 ( .A(n246), .B(a[18]), .Z(n785) );
  XOR U938 ( .A(n2537), .B(n785), .Z(n787) );
  NANDN U939 ( .A(b[0]), .B(a[17]), .Z(n786) );
  AND U940 ( .A(n787), .B(n786), .Z(n811) );
  NANDN U941 ( .A(n788), .B(n2625), .Z(n791) );
  XOR U942 ( .A(b[5]), .B(n789), .Z(n824) );
  OR U943 ( .A(n824), .B(n2608), .Z(n790) );
  NAND U944 ( .A(n791), .B(n790), .Z(n809) );
  NANDN U945 ( .A(n2695), .B(a[10]), .Z(n810) );
  XNOR U946 ( .A(n809), .B(n810), .Z(n812) );
  XOR U947 ( .A(n811), .B(n812), .Z(n808) );
  XOR U948 ( .A(n807), .B(n808), .Z(n827) );
  XOR U949 ( .A(n828), .B(n827), .Z(n829) );
  XNOR U950 ( .A(n830), .B(n829), .Z(n801) );
  XNOR U951 ( .A(n801), .B(n802), .Z(n803) );
  XNOR U952 ( .A(n804), .B(n803), .Z(n833) );
  XNOR U953 ( .A(n833), .B(sreg[74]), .Z(n835) );
  NAND U954 ( .A(n796), .B(sreg[73]), .Z(n800) );
  OR U955 ( .A(n798), .B(n797), .Z(n799) );
  AND U956 ( .A(n800), .B(n799), .Z(n834) );
  XOR U957 ( .A(n835), .B(n834), .Z(c[74]) );
  NANDN U958 ( .A(n810), .B(n809), .Z(n814) );
  NAND U959 ( .A(n812), .B(n811), .Z(n813) );
  NAND U960 ( .A(n814), .B(n813), .Z(n865) );
  NAND U961 ( .A(n815), .B(n2666), .Z(n817) );
  XNOR U962 ( .A(n2695), .B(a[13]), .Z(n852) );
  NAND U963 ( .A(n852), .B(n2665), .Z(n816) );
  NAND U964 ( .A(n817), .B(n816), .Z(n842) );
  XNOR U965 ( .A(b[3]), .B(a[17]), .Z(n855) );
  NANDN U966 ( .A(n855), .B(n2561), .Z(n820) );
  NANDN U967 ( .A(n818), .B(n2563), .Z(n819) );
  AND U968 ( .A(n820), .B(n819), .Z(n843) );
  XNOR U969 ( .A(n842), .B(n843), .Z(n844) );
  NANDN U970 ( .A(n246), .B(a[19]), .Z(n821) );
  XOR U971 ( .A(n2537), .B(n821), .Z(n823) );
  NANDN U972 ( .A(b[0]), .B(a[18]), .Z(n822) );
  AND U973 ( .A(n823), .B(n822), .Z(n848) );
  NANDN U974 ( .A(n824), .B(n2625), .Z(n826) );
  XNOR U975 ( .A(b[5]), .B(a[15]), .Z(n861) );
  OR U976 ( .A(n861), .B(n2608), .Z(n825) );
  NAND U977 ( .A(n826), .B(n825), .Z(n846) );
  NANDN U978 ( .A(n2695), .B(a[11]), .Z(n847) );
  XNOR U979 ( .A(n846), .B(n847), .Z(n849) );
  XOR U980 ( .A(n848), .B(n849), .Z(n845) );
  XOR U981 ( .A(n844), .B(n845), .Z(n864) );
  XOR U982 ( .A(n865), .B(n864), .Z(n866) );
  XNOR U983 ( .A(n867), .B(n866), .Z(n838) );
  NAND U984 ( .A(n828), .B(n827), .Z(n832) );
  NAND U985 ( .A(n830), .B(n829), .Z(n831) );
  NAND U986 ( .A(n832), .B(n831), .Z(n839) );
  XNOR U987 ( .A(n838), .B(n839), .Z(n840) );
  XNOR U988 ( .A(n841), .B(n840), .Z(n870) );
  XNOR U989 ( .A(n870), .B(sreg[75]), .Z(n872) );
  NAND U990 ( .A(n833), .B(sreg[74]), .Z(n837) );
  OR U991 ( .A(n835), .B(n834), .Z(n836) );
  AND U992 ( .A(n837), .B(n836), .Z(n871) );
  XOR U993 ( .A(n872), .B(n871), .Z(c[75]) );
  NANDN U994 ( .A(n847), .B(n846), .Z(n851) );
  NAND U995 ( .A(n849), .B(n848), .Z(n850) );
  NAND U996 ( .A(n851), .B(n850), .Z(n902) );
  NAND U997 ( .A(n852), .B(n2666), .Z(n854) );
  XNOR U998 ( .A(n2695), .B(a[14]), .Z(n889) );
  NAND U999 ( .A(n889), .B(n2665), .Z(n853) );
  NAND U1000 ( .A(n854), .B(n853), .Z(n879) );
  XNOR U1001 ( .A(b[3]), .B(a[18]), .Z(n892) );
  NANDN U1002 ( .A(n892), .B(n2561), .Z(n857) );
  NANDN U1003 ( .A(n855), .B(n2563), .Z(n856) );
  AND U1004 ( .A(n857), .B(n856), .Z(n880) );
  XNOR U1005 ( .A(n879), .B(n880), .Z(n881) );
  NANDN U1006 ( .A(n246), .B(a[20]), .Z(n858) );
  XOR U1007 ( .A(n2537), .B(n858), .Z(n860) );
  NANDN U1008 ( .A(b[0]), .B(a[19]), .Z(n859) );
  AND U1009 ( .A(n860), .B(n859), .Z(n885) );
  NANDN U1010 ( .A(n861), .B(n2625), .Z(n863) );
  XNOR U1011 ( .A(b[5]), .B(a[16]), .Z(n898) );
  OR U1012 ( .A(n898), .B(n2608), .Z(n862) );
  NAND U1013 ( .A(n863), .B(n862), .Z(n883) );
  NANDN U1014 ( .A(n2695), .B(a[12]), .Z(n884) );
  XNOR U1015 ( .A(n883), .B(n884), .Z(n886) );
  XOR U1016 ( .A(n885), .B(n886), .Z(n882) );
  XOR U1017 ( .A(n881), .B(n882), .Z(n901) );
  XOR U1018 ( .A(n902), .B(n901), .Z(n903) );
  XNOR U1019 ( .A(n904), .B(n903), .Z(n875) );
  NAND U1020 ( .A(n865), .B(n864), .Z(n869) );
  NAND U1021 ( .A(n867), .B(n866), .Z(n868) );
  NAND U1022 ( .A(n869), .B(n868), .Z(n876) );
  XNOR U1023 ( .A(n875), .B(n876), .Z(n877) );
  XNOR U1024 ( .A(n878), .B(n877), .Z(n907) );
  XNOR U1025 ( .A(n907), .B(sreg[76]), .Z(n909) );
  NAND U1026 ( .A(n870), .B(sreg[75]), .Z(n874) );
  OR U1027 ( .A(n872), .B(n871), .Z(n873) );
  AND U1028 ( .A(n874), .B(n873), .Z(n908) );
  XOR U1029 ( .A(n909), .B(n908), .Z(c[76]) );
  NANDN U1030 ( .A(n884), .B(n883), .Z(n888) );
  NAND U1031 ( .A(n886), .B(n885), .Z(n887) );
  NAND U1032 ( .A(n888), .B(n887), .Z(n939) );
  NAND U1033 ( .A(n889), .B(n2666), .Z(n891) );
  XNOR U1034 ( .A(n2695), .B(a[15]), .Z(n932) );
  NAND U1035 ( .A(n932), .B(n2665), .Z(n890) );
  NAND U1036 ( .A(n891), .B(n890), .Z(n916) );
  XNOR U1037 ( .A(b[3]), .B(a[19]), .Z(n935) );
  NANDN U1038 ( .A(n935), .B(n2561), .Z(n894) );
  NANDN U1039 ( .A(n892), .B(n2563), .Z(n893) );
  AND U1040 ( .A(n894), .B(n893), .Z(n917) );
  XNOR U1041 ( .A(n916), .B(n917), .Z(n918) );
  NANDN U1042 ( .A(n246), .B(a[21]), .Z(n895) );
  XOR U1043 ( .A(n2537), .B(n895), .Z(n897) );
  IV U1044 ( .A(a[20]), .Z(n1150) );
  NANDN U1045 ( .A(n1150), .B(n246), .Z(n896) );
  AND U1046 ( .A(n897), .B(n896), .Z(n922) );
  NANDN U1047 ( .A(n898), .B(n2625), .Z(n900) );
  XNOR U1048 ( .A(n248), .B(a[17]), .Z(n926) );
  NANDN U1049 ( .A(n2608), .B(n926), .Z(n899) );
  NAND U1050 ( .A(n900), .B(n899), .Z(n920) );
  NANDN U1051 ( .A(n2695), .B(a[13]), .Z(n921) );
  XNOR U1052 ( .A(n920), .B(n921), .Z(n923) );
  XOR U1053 ( .A(n922), .B(n923), .Z(n919) );
  XOR U1054 ( .A(n918), .B(n919), .Z(n938) );
  XOR U1055 ( .A(n939), .B(n938), .Z(n940) );
  XNOR U1056 ( .A(n941), .B(n940), .Z(n912) );
  NAND U1057 ( .A(n902), .B(n901), .Z(n906) );
  NAND U1058 ( .A(n904), .B(n903), .Z(n905) );
  NAND U1059 ( .A(n906), .B(n905), .Z(n913) );
  XNOR U1060 ( .A(n912), .B(n913), .Z(n914) );
  XNOR U1061 ( .A(n915), .B(n914), .Z(n944) );
  XNOR U1062 ( .A(n944), .B(sreg[77]), .Z(n946) );
  NAND U1063 ( .A(n907), .B(sreg[76]), .Z(n911) );
  OR U1064 ( .A(n909), .B(n908), .Z(n910) );
  AND U1065 ( .A(n911), .B(n910), .Z(n945) );
  XOR U1066 ( .A(n946), .B(n945), .Z(c[77]) );
  NANDN U1067 ( .A(n921), .B(n920), .Z(n925) );
  NAND U1068 ( .A(n923), .B(n922), .Z(n924) );
  NAND U1069 ( .A(n925), .B(n924), .Z(n977) );
  AND U1070 ( .A(a[14]), .B(b[7]), .Z(n972) );
  XNOR U1071 ( .A(b[5]), .B(a[18]), .Z(n962) );
  OR U1072 ( .A(n962), .B(n2608), .Z(n928) );
  NAND U1073 ( .A(n2625), .B(n926), .Z(n927) );
  NAND U1074 ( .A(n928), .B(n927), .Z(n971) );
  XOR U1075 ( .A(n972), .B(n971), .Z(n973) );
  NANDN U1076 ( .A(n246), .B(a[22]), .Z(n929) );
  XOR U1077 ( .A(n2537), .B(n929), .Z(n931) );
  NANDN U1078 ( .A(b[0]), .B(a[21]), .Z(n930) );
  AND U1079 ( .A(n931), .B(n930), .Z(n974) );
  XOR U1080 ( .A(n973), .B(n974), .Z(n968) );
  NAND U1081 ( .A(n932), .B(n2666), .Z(n934) );
  XNOR U1082 ( .A(n2695), .B(a[16]), .Z(n953) );
  NAND U1083 ( .A(n953), .B(n2665), .Z(n933) );
  NAND U1084 ( .A(n934), .B(n933), .Z(n965) );
  XOR U1085 ( .A(b[3]), .B(n1150), .Z(n956) );
  NANDN U1086 ( .A(n956), .B(n2561), .Z(n937) );
  NANDN U1087 ( .A(n935), .B(n2563), .Z(n936) );
  AND U1088 ( .A(n937), .B(n936), .Z(n966) );
  XNOR U1089 ( .A(n965), .B(n966), .Z(n967) );
  XNOR U1090 ( .A(n968), .B(n967), .Z(n978) );
  XNOR U1091 ( .A(n977), .B(n978), .Z(n979) );
  XNOR U1092 ( .A(n980), .B(n979), .Z(n949) );
  NAND U1093 ( .A(n939), .B(n938), .Z(n943) );
  NAND U1094 ( .A(n941), .B(n940), .Z(n942) );
  NAND U1095 ( .A(n943), .B(n942), .Z(n950) );
  XNOR U1096 ( .A(n949), .B(n950), .Z(n951) );
  XNOR U1097 ( .A(n952), .B(n951), .Z(n983) );
  XNOR U1098 ( .A(n983), .B(sreg[78]), .Z(n985) );
  NAND U1099 ( .A(n944), .B(sreg[77]), .Z(n948) );
  OR U1100 ( .A(n946), .B(n945), .Z(n947) );
  AND U1101 ( .A(n948), .B(n947), .Z(n984) );
  XOR U1102 ( .A(n985), .B(n984), .Z(c[78]) );
  NAND U1103 ( .A(n953), .B(n2666), .Z(n955) );
  XNOR U1104 ( .A(n2695), .B(a[17]), .Z(n1002) );
  NAND U1105 ( .A(n1002), .B(n2665), .Z(n954) );
  NAND U1106 ( .A(n955), .B(n954), .Z(n992) );
  XNOR U1107 ( .A(b[3]), .B(a[21]), .Z(n1005) );
  NANDN U1108 ( .A(n1005), .B(n2561), .Z(n958) );
  NANDN U1109 ( .A(n956), .B(n2563), .Z(n957) );
  AND U1110 ( .A(n958), .B(n957), .Z(n993) );
  XNOR U1111 ( .A(n992), .B(n993), .Z(n994) );
  NANDN U1112 ( .A(n246), .B(a[23]), .Z(n959) );
  XOR U1113 ( .A(n2537), .B(n959), .Z(n961) );
  NANDN U1114 ( .A(b[0]), .B(a[22]), .Z(n960) );
  AND U1115 ( .A(n961), .B(n960), .Z(n998) );
  NANDN U1116 ( .A(n962), .B(n2625), .Z(n964) );
  XNOR U1117 ( .A(b[5]), .B(a[19]), .Z(n1011) );
  OR U1118 ( .A(n1011), .B(n2608), .Z(n963) );
  NAND U1119 ( .A(n964), .B(n963), .Z(n996) );
  NANDN U1120 ( .A(n2695), .B(a[15]), .Z(n997) );
  XNOR U1121 ( .A(n996), .B(n997), .Z(n999) );
  XOR U1122 ( .A(n998), .B(n999), .Z(n995) );
  XOR U1123 ( .A(n994), .B(n995), .Z(n1016) );
  NANDN U1124 ( .A(n966), .B(n965), .Z(n970) );
  NAND U1125 ( .A(n968), .B(n967), .Z(n969) );
  NAND U1126 ( .A(n970), .B(n969), .Z(n1014) );
  OR U1127 ( .A(n972), .B(n971), .Z(n976) );
  NANDN U1128 ( .A(n974), .B(n973), .Z(n975) );
  NAND U1129 ( .A(n976), .B(n975), .Z(n1015) );
  XNOR U1130 ( .A(n1014), .B(n1015), .Z(n1017) );
  XNOR U1131 ( .A(n1016), .B(n1017), .Z(n988) );
  NANDN U1132 ( .A(n978), .B(n977), .Z(n982) );
  NAND U1133 ( .A(n980), .B(n979), .Z(n981) );
  NAND U1134 ( .A(n982), .B(n981), .Z(n989) );
  XNOR U1135 ( .A(n988), .B(n989), .Z(n990) );
  XNOR U1136 ( .A(n991), .B(n990), .Z(n1020) );
  XNOR U1137 ( .A(n1020), .B(sreg[79]), .Z(n1022) );
  NAND U1138 ( .A(n983), .B(sreg[78]), .Z(n987) );
  OR U1139 ( .A(n985), .B(n984), .Z(n986) );
  AND U1140 ( .A(n987), .B(n986), .Z(n1021) );
  XOR U1141 ( .A(n1022), .B(n1021), .Z(c[79]) );
  NANDN U1142 ( .A(n997), .B(n996), .Z(n1001) );
  NAND U1143 ( .A(n999), .B(n998), .Z(n1000) );
  NAND U1144 ( .A(n1001), .B(n1000), .Z(n1052) );
  NAND U1145 ( .A(n1002), .B(n2666), .Z(n1004) );
  XNOR U1146 ( .A(n2695), .B(a[18]), .Z(n1039) );
  NAND U1147 ( .A(n1039), .B(n2665), .Z(n1003) );
  NAND U1148 ( .A(n1004), .B(n1003), .Z(n1029) );
  XNOR U1149 ( .A(b[3]), .B(a[22]), .Z(n1042) );
  NANDN U1150 ( .A(n1042), .B(n2561), .Z(n1007) );
  NANDN U1151 ( .A(n1005), .B(n2563), .Z(n1006) );
  AND U1152 ( .A(n1007), .B(n1006), .Z(n1030) );
  XNOR U1153 ( .A(n1029), .B(n1030), .Z(n1031) );
  NANDN U1154 ( .A(n246), .B(a[24]), .Z(n1008) );
  XOR U1155 ( .A(n2537), .B(n1008), .Z(n1010) );
  NANDN U1156 ( .A(b[0]), .B(a[23]), .Z(n1009) );
  AND U1157 ( .A(n1010), .B(n1009), .Z(n1035) );
  NANDN U1158 ( .A(n1011), .B(n2625), .Z(n1013) );
  XOR U1159 ( .A(b[5]), .B(n1150), .Z(n1048) );
  OR U1160 ( .A(n1048), .B(n2608), .Z(n1012) );
  NAND U1161 ( .A(n1013), .B(n1012), .Z(n1033) );
  NANDN U1162 ( .A(n2695), .B(a[16]), .Z(n1034) );
  XNOR U1163 ( .A(n1033), .B(n1034), .Z(n1036) );
  XOR U1164 ( .A(n1035), .B(n1036), .Z(n1032) );
  XOR U1165 ( .A(n1031), .B(n1032), .Z(n1051) );
  XOR U1166 ( .A(n1052), .B(n1051), .Z(n1053) );
  XNOR U1167 ( .A(n1054), .B(n1053), .Z(n1025) );
  NANDN U1168 ( .A(n1015), .B(n1014), .Z(n1019) );
  NAND U1169 ( .A(n1017), .B(n1016), .Z(n1018) );
  NAND U1170 ( .A(n1019), .B(n1018), .Z(n1026) );
  XNOR U1171 ( .A(n1025), .B(n1026), .Z(n1027) );
  XNOR U1172 ( .A(n1028), .B(n1027), .Z(n1057) );
  XNOR U1173 ( .A(n1057), .B(sreg[80]), .Z(n1059) );
  NAND U1174 ( .A(n1020), .B(sreg[79]), .Z(n1024) );
  OR U1175 ( .A(n1022), .B(n1021), .Z(n1023) );
  AND U1176 ( .A(n1024), .B(n1023), .Z(n1058) );
  XOR U1177 ( .A(n1059), .B(n1058), .Z(c[80]) );
  NANDN U1178 ( .A(n1034), .B(n1033), .Z(n1038) );
  NAND U1179 ( .A(n1036), .B(n1035), .Z(n1037) );
  NAND U1180 ( .A(n1038), .B(n1037), .Z(n1089) );
  NAND U1181 ( .A(n1039), .B(n2666), .Z(n1041) );
  XNOR U1182 ( .A(n2695), .B(a[19]), .Z(n1076) );
  NAND U1183 ( .A(n1076), .B(n2665), .Z(n1040) );
  NAND U1184 ( .A(n1041), .B(n1040), .Z(n1066) );
  XNOR U1185 ( .A(b[3]), .B(a[23]), .Z(n1079) );
  NANDN U1186 ( .A(n1079), .B(n2561), .Z(n1044) );
  NANDN U1187 ( .A(n1042), .B(n2563), .Z(n1043) );
  AND U1188 ( .A(n1044), .B(n1043), .Z(n1067) );
  XNOR U1189 ( .A(n1066), .B(n1067), .Z(n1068) );
  NANDN U1190 ( .A(n246), .B(a[25]), .Z(n1045) );
  XOR U1191 ( .A(n2537), .B(n1045), .Z(n1047) );
  NANDN U1192 ( .A(b[0]), .B(a[24]), .Z(n1046) );
  AND U1193 ( .A(n1047), .B(n1046), .Z(n1072) );
  NANDN U1194 ( .A(n1048), .B(n2625), .Z(n1050) );
  XNOR U1195 ( .A(b[5]), .B(a[21]), .Z(n1085) );
  OR U1196 ( .A(n1085), .B(n2608), .Z(n1049) );
  NAND U1197 ( .A(n1050), .B(n1049), .Z(n1070) );
  NANDN U1198 ( .A(n2695), .B(a[17]), .Z(n1071) );
  XNOR U1199 ( .A(n1070), .B(n1071), .Z(n1073) );
  XOR U1200 ( .A(n1072), .B(n1073), .Z(n1069) );
  XOR U1201 ( .A(n1068), .B(n1069), .Z(n1088) );
  XOR U1202 ( .A(n1089), .B(n1088), .Z(n1090) );
  XNOR U1203 ( .A(n1091), .B(n1090), .Z(n1062) );
  NAND U1204 ( .A(n1052), .B(n1051), .Z(n1056) );
  NAND U1205 ( .A(n1054), .B(n1053), .Z(n1055) );
  NAND U1206 ( .A(n1056), .B(n1055), .Z(n1063) );
  XNOR U1207 ( .A(n1062), .B(n1063), .Z(n1064) );
  XNOR U1208 ( .A(n1065), .B(n1064), .Z(n1094) );
  XNOR U1209 ( .A(n1094), .B(sreg[81]), .Z(n1096) );
  NAND U1210 ( .A(n1057), .B(sreg[80]), .Z(n1061) );
  OR U1211 ( .A(n1059), .B(n1058), .Z(n1060) );
  AND U1212 ( .A(n1061), .B(n1060), .Z(n1095) );
  XOR U1213 ( .A(n1096), .B(n1095), .Z(c[81]) );
  NANDN U1214 ( .A(n1071), .B(n1070), .Z(n1075) );
  NAND U1215 ( .A(n1073), .B(n1072), .Z(n1074) );
  NAND U1216 ( .A(n1075), .B(n1074), .Z(n1126) );
  NAND U1217 ( .A(n1076), .B(n2666), .Z(n1078) );
  XNOR U1218 ( .A(n2695), .B(a[20]), .Z(n1113) );
  NAND U1219 ( .A(n1113), .B(n2665), .Z(n1077) );
  NAND U1220 ( .A(n1078), .B(n1077), .Z(n1103) );
  XNOR U1221 ( .A(b[3]), .B(a[24]), .Z(n1116) );
  NANDN U1222 ( .A(n1116), .B(n2561), .Z(n1081) );
  NANDN U1223 ( .A(n1079), .B(n2563), .Z(n1080) );
  AND U1224 ( .A(n1081), .B(n1080), .Z(n1104) );
  XNOR U1225 ( .A(n1103), .B(n1104), .Z(n1105) );
  NANDN U1226 ( .A(n246), .B(a[26]), .Z(n1082) );
  XOR U1227 ( .A(n2537), .B(n1082), .Z(n1084) );
  NANDN U1228 ( .A(b[0]), .B(a[25]), .Z(n1083) );
  AND U1229 ( .A(n1084), .B(n1083), .Z(n1109) );
  NANDN U1230 ( .A(n1085), .B(n2625), .Z(n1087) );
  XNOR U1231 ( .A(b[5]), .B(a[22]), .Z(n1122) );
  OR U1232 ( .A(n1122), .B(n2608), .Z(n1086) );
  NAND U1233 ( .A(n1087), .B(n1086), .Z(n1107) );
  NANDN U1234 ( .A(n2695), .B(a[18]), .Z(n1108) );
  XNOR U1235 ( .A(n1107), .B(n1108), .Z(n1110) );
  XOR U1236 ( .A(n1109), .B(n1110), .Z(n1106) );
  XOR U1237 ( .A(n1105), .B(n1106), .Z(n1125) );
  XOR U1238 ( .A(n1126), .B(n1125), .Z(n1127) );
  XNOR U1239 ( .A(n1128), .B(n1127), .Z(n1099) );
  NAND U1240 ( .A(n1089), .B(n1088), .Z(n1093) );
  NAND U1241 ( .A(n1091), .B(n1090), .Z(n1092) );
  NAND U1242 ( .A(n1093), .B(n1092), .Z(n1100) );
  XNOR U1243 ( .A(n1099), .B(n1100), .Z(n1101) );
  XNOR U1244 ( .A(n1102), .B(n1101), .Z(n1131) );
  XNOR U1245 ( .A(n1131), .B(sreg[82]), .Z(n1133) );
  NAND U1246 ( .A(n1094), .B(sreg[81]), .Z(n1098) );
  OR U1247 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U1248 ( .A(n1098), .B(n1097), .Z(n1132) );
  XOR U1249 ( .A(n1133), .B(n1132), .Z(c[82]) );
  NANDN U1250 ( .A(n1108), .B(n1107), .Z(n1112) );
  NAND U1251 ( .A(n1110), .B(n1109), .Z(n1111) );
  NAND U1252 ( .A(n1112), .B(n1111), .Z(n1164) );
  NAND U1253 ( .A(n1113), .B(n2666), .Z(n1115) );
  XNOR U1254 ( .A(n2695), .B(a[21]), .Z(n1157) );
  NAND U1255 ( .A(n1157), .B(n2665), .Z(n1114) );
  NAND U1256 ( .A(n1115), .B(n1114), .Z(n1140) );
  XNOR U1257 ( .A(b[3]), .B(a[25]), .Z(n1160) );
  NANDN U1258 ( .A(n1160), .B(n2561), .Z(n1118) );
  NANDN U1259 ( .A(n1116), .B(n2563), .Z(n1117) );
  AND U1260 ( .A(n1118), .B(n1117), .Z(n1141) );
  XNOR U1261 ( .A(n1140), .B(n1141), .Z(n1142) );
  NANDN U1262 ( .A(n246), .B(a[27]), .Z(n1119) );
  XOR U1263 ( .A(n2537), .B(n1119), .Z(n1121) );
  NANDN U1264 ( .A(b[0]), .B(a[26]), .Z(n1120) );
  AND U1265 ( .A(n1121), .B(n1120), .Z(n1146) );
  NANDN U1266 ( .A(n1122), .B(n2625), .Z(n1124) );
  XNOR U1267 ( .A(n248), .B(a[23]), .Z(n1151) );
  NANDN U1268 ( .A(n2608), .B(n1151), .Z(n1123) );
  NAND U1269 ( .A(n1124), .B(n1123), .Z(n1144) );
  NANDN U1270 ( .A(n2695), .B(a[19]), .Z(n1145) );
  XNOR U1271 ( .A(n1144), .B(n1145), .Z(n1147) );
  XOR U1272 ( .A(n1146), .B(n1147), .Z(n1143) );
  XOR U1273 ( .A(n1142), .B(n1143), .Z(n1163) );
  XOR U1274 ( .A(n1164), .B(n1163), .Z(n1165) );
  XNOR U1275 ( .A(n1166), .B(n1165), .Z(n1136) );
  NAND U1276 ( .A(n1126), .B(n1125), .Z(n1130) );
  NAND U1277 ( .A(n1128), .B(n1127), .Z(n1129) );
  NAND U1278 ( .A(n1130), .B(n1129), .Z(n1137) );
  XNOR U1279 ( .A(n1136), .B(n1137), .Z(n1138) );
  XNOR U1280 ( .A(n1139), .B(n1138), .Z(n1169) );
  XNOR U1281 ( .A(n1169), .B(sreg[83]), .Z(n1171) );
  NAND U1282 ( .A(n1131), .B(sreg[82]), .Z(n1135) );
  OR U1283 ( .A(n1133), .B(n1132), .Z(n1134) );
  AND U1284 ( .A(n1135), .B(n1134), .Z(n1170) );
  XOR U1285 ( .A(n1171), .B(n1170), .Z(c[83]) );
  NANDN U1286 ( .A(n1145), .B(n1144), .Z(n1149) );
  NAND U1287 ( .A(n1147), .B(n1146), .Z(n1148) );
  NAND U1288 ( .A(n1149), .B(n1148), .Z(n1202) );
  ANDN U1289 ( .B(b[7]), .A(n1150), .Z(n1184) );
  XNOR U1290 ( .A(b[5]), .B(a[24]), .Z(n1199) );
  OR U1291 ( .A(n1199), .B(n2608), .Z(n1153) );
  NAND U1292 ( .A(n2625), .B(n1151), .Z(n1152) );
  NAND U1293 ( .A(n1153), .B(n1152), .Z(n1185) );
  XOR U1294 ( .A(n1184), .B(n1185), .Z(n1186) );
  NANDN U1295 ( .A(n246), .B(a[28]), .Z(n1154) );
  XOR U1296 ( .A(n2537), .B(n1154), .Z(n1156) );
  NANDN U1297 ( .A(b[0]), .B(a[27]), .Z(n1155) );
  AND U1298 ( .A(n1156), .B(n1155), .Z(n1187) );
  XOR U1299 ( .A(n1186), .B(n1187), .Z(n1181) );
  NAND U1300 ( .A(n1157), .B(n2666), .Z(n1159) );
  XNOR U1301 ( .A(n2695), .B(a[22]), .Z(n1190) );
  NAND U1302 ( .A(n1190), .B(n2665), .Z(n1158) );
  NAND U1303 ( .A(n1159), .B(n1158), .Z(n1178) );
  XNOR U1304 ( .A(b[3]), .B(a[26]), .Z(n1193) );
  NANDN U1305 ( .A(n1193), .B(n2561), .Z(n1162) );
  NANDN U1306 ( .A(n1160), .B(n2563), .Z(n1161) );
  AND U1307 ( .A(n1162), .B(n1161), .Z(n1179) );
  XNOR U1308 ( .A(n1178), .B(n1179), .Z(n1180) );
  XNOR U1309 ( .A(n1181), .B(n1180), .Z(n1203) );
  XNOR U1310 ( .A(n1202), .B(n1203), .Z(n1204) );
  XNOR U1311 ( .A(n1205), .B(n1204), .Z(n1174) );
  NAND U1312 ( .A(n1164), .B(n1163), .Z(n1168) );
  NAND U1313 ( .A(n1166), .B(n1165), .Z(n1167) );
  NAND U1314 ( .A(n1168), .B(n1167), .Z(n1175) );
  XNOR U1315 ( .A(n1174), .B(n1175), .Z(n1176) );
  XNOR U1316 ( .A(n1177), .B(n1176), .Z(n1208) );
  XNOR U1317 ( .A(n1208), .B(sreg[84]), .Z(n1210) );
  NAND U1318 ( .A(n1169), .B(sreg[83]), .Z(n1173) );
  OR U1319 ( .A(n1171), .B(n1170), .Z(n1172) );
  AND U1320 ( .A(n1173), .B(n1172), .Z(n1209) );
  XOR U1321 ( .A(n1210), .B(n1209), .Z(c[84]) );
  NANDN U1322 ( .A(n1179), .B(n1178), .Z(n1183) );
  NAND U1323 ( .A(n1181), .B(n1180), .Z(n1182) );
  NAND U1324 ( .A(n1183), .B(n1182), .Z(n1242) );
  OR U1325 ( .A(n1185), .B(n1184), .Z(n1189) );
  NANDN U1326 ( .A(n1187), .B(n1186), .Z(n1188) );
  NAND U1327 ( .A(n1189), .B(n1188), .Z(n1240) );
  NAND U1328 ( .A(n1190), .B(n2666), .Z(n1192) );
  XNOR U1329 ( .A(n2695), .B(a[23]), .Z(n1227) );
  NAND U1330 ( .A(n1227), .B(n2665), .Z(n1191) );
  NAND U1331 ( .A(n1192), .B(n1191), .Z(n1217) );
  XNOR U1332 ( .A(b[3]), .B(a[27]), .Z(n1230) );
  NANDN U1333 ( .A(n1230), .B(n2561), .Z(n1195) );
  NANDN U1334 ( .A(n1193), .B(n2563), .Z(n1194) );
  AND U1335 ( .A(n1195), .B(n1194), .Z(n1218) );
  XNOR U1336 ( .A(n1217), .B(n1218), .Z(n1219) );
  NANDN U1337 ( .A(n246), .B(a[29]), .Z(n1196) );
  XOR U1338 ( .A(n2537), .B(n1196), .Z(n1198) );
  NANDN U1339 ( .A(b[0]), .B(a[28]), .Z(n1197) );
  AND U1340 ( .A(n1198), .B(n1197), .Z(n1223) );
  NANDN U1341 ( .A(n1199), .B(n2625), .Z(n1201) );
  XNOR U1342 ( .A(b[5]), .B(a[25]), .Z(n1236) );
  OR U1343 ( .A(n1236), .B(n2608), .Z(n1200) );
  NAND U1344 ( .A(n1201), .B(n1200), .Z(n1221) );
  NANDN U1345 ( .A(n2695), .B(a[21]), .Z(n1222) );
  XNOR U1346 ( .A(n1221), .B(n1222), .Z(n1224) );
  XOR U1347 ( .A(n1223), .B(n1224), .Z(n1220) );
  XOR U1348 ( .A(n1219), .B(n1220), .Z(n1239) );
  XNOR U1349 ( .A(n1240), .B(n1239), .Z(n1241) );
  XNOR U1350 ( .A(n1242), .B(n1241), .Z(n1213) );
  NANDN U1351 ( .A(n1203), .B(n1202), .Z(n1207) );
  NAND U1352 ( .A(n1205), .B(n1204), .Z(n1206) );
  NAND U1353 ( .A(n1207), .B(n1206), .Z(n1214) );
  XNOR U1354 ( .A(n1213), .B(n1214), .Z(n1215) );
  XNOR U1355 ( .A(n1216), .B(n1215), .Z(n1243) );
  XNOR U1356 ( .A(n1243), .B(sreg[85]), .Z(n1245) );
  NAND U1357 ( .A(n1208), .B(sreg[84]), .Z(n1212) );
  OR U1358 ( .A(n1210), .B(n1209), .Z(n1211) );
  AND U1359 ( .A(n1212), .B(n1211), .Z(n1244) );
  XOR U1360 ( .A(n1245), .B(n1244), .Z(c[85]) );
  NANDN U1361 ( .A(n1222), .B(n1221), .Z(n1226) );
  NAND U1362 ( .A(n1224), .B(n1223), .Z(n1225) );
  NAND U1363 ( .A(n1226), .B(n1225), .Z(n1275) );
  NAND U1364 ( .A(n1227), .B(n2666), .Z(n1229) );
  XNOR U1365 ( .A(n2695), .B(a[24]), .Z(n1262) );
  NAND U1366 ( .A(n1262), .B(n2665), .Z(n1228) );
  NAND U1367 ( .A(n1229), .B(n1228), .Z(n1252) );
  XNOR U1368 ( .A(b[3]), .B(a[28]), .Z(n1265) );
  NANDN U1369 ( .A(n1265), .B(n2561), .Z(n1232) );
  NANDN U1370 ( .A(n1230), .B(n2563), .Z(n1231) );
  AND U1371 ( .A(n1232), .B(n1231), .Z(n1253) );
  XNOR U1372 ( .A(n1252), .B(n1253), .Z(n1254) );
  NANDN U1373 ( .A(n246), .B(a[30]), .Z(n1233) );
  XOR U1374 ( .A(n2537), .B(n1233), .Z(n1235) );
  NANDN U1375 ( .A(b[0]), .B(a[29]), .Z(n1234) );
  AND U1376 ( .A(n1235), .B(n1234), .Z(n1258) );
  NANDN U1377 ( .A(n1236), .B(n2625), .Z(n1238) );
  XNOR U1378 ( .A(b[5]), .B(a[26]), .Z(n1271) );
  OR U1379 ( .A(n1271), .B(n2608), .Z(n1237) );
  NAND U1380 ( .A(n1238), .B(n1237), .Z(n1256) );
  NANDN U1381 ( .A(n2695), .B(a[22]), .Z(n1257) );
  XNOR U1382 ( .A(n1256), .B(n1257), .Z(n1259) );
  XOR U1383 ( .A(n1258), .B(n1259), .Z(n1255) );
  XOR U1384 ( .A(n1254), .B(n1255), .Z(n1274) );
  XOR U1385 ( .A(n1275), .B(n1274), .Z(n1276) );
  XNOR U1386 ( .A(n1277), .B(n1276), .Z(n1248) );
  XNOR U1387 ( .A(n1248), .B(n1249), .Z(n1250) );
  XNOR U1388 ( .A(n1251), .B(n1250), .Z(n1280) );
  XNOR U1389 ( .A(n1280), .B(sreg[86]), .Z(n1282) );
  NAND U1390 ( .A(n1243), .B(sreg[85]), .Z(n1247) );
  OR U1391 ( .A(n1245), .B(n1244), .Z(n1246) );
  AND U1392 ( .A(n1247), .B(n1246), .Z(n1281) );
  XOR U1393 ( .A(n1282), .B(n1281), .Z(c[86]) );
  NANDN U1394 ( .A(n1257), .B(n1256), .Z(n1261) );
  NAND U1395 ( .A(n1259), .B(n1258), .Z(n1260) );
  NAND U1396 ( .A(n1261), .B(n1260), .Z(n1312) );
  NAND U1397 ( .A(n1262), .B(n2666), .Z(n1264) );
  XNOR U1398 ( .A(n2695), .B(a[25]), .Z(n1299) );
  NAND U1399 ( .A(n1299), .B(n2665), .Z(n1263) );
  NAND U1400 ( .A(n1264), .B(n1263), .Z(n1289) );
  XNOR U1401 ( .A(b[3]), .B(a[29]), .Z(n1302) );
  NANDN U1402 ( .A(n1302), .B(n2561), .Z(n1267) );
  NANDN U1403 ( .A(n1265), .B(n2563), .Z(n1266) );
  AND U1404 ( .A(n1267), .B(n1266), .Z(n1290) );
  XNOR U1405 ( .A(n1289), .B(n1290), .Z(n1291) );
  NANDN U1406 ( .A(n246), .B(a[31]), .Z(n1268) );
  XOR U1407 ( .A(n2537), .B(n1268), .Z(n1270) );
  NANDN U1408 ( .A(b[0]), .B(a[30]), .Z(n1269) );
  AND U1409 ( .A(n1270), .B(n1269), .Z(n1295) );
  NANDN U1410 ( .A(n1271), .B(n2625), .Z(n1273) );
  XNOR U1411 ( .A(b[5]), .B(a[27]), .Z(n1308) );
  OR U1412 ( .A(n1308), .B(n2608), .Z(n1272) );
  NAND U1413 ( .A(n1273), .B(n1272), .Z(n1293) );
  NANDN U1414 ( .A(n2695), .B(a[23]), .Z(n1294) );
  XNOR U1415 ( .A(n1293), .B(n1294), .Z(n1296) );
  XOR U1416 ( .A(n1295), .B(n1296), .Z(n1292) );
  XOR U1417 ( .A(n1291), .B(n1292), .Z(n1311) );
  XOR U1418 ( .A(n1312), .B(n1311), .Z(n1313) );
  XNOR U1419 ( .A(n1314), .B(n1313), .Z(n1285) );
  NAND U1420 ( .A(n1275), .B(n1274), .Z(n1279) );
  NAND U1421 ( .A(n1277), .B(n1276), .Z(n1278) );
  NAND U1422 ( .A(n1279), .B(n1278), .Z(n1286) );
  XNOR U1423 ( .A(n1285), .B(n1286), .Z(n1287) );
  XNOR U1424 ( .A(n1288), .B(n1287), .Z(n1317) );
  XNOR U1425 ( .A(n1317), .B(sreg[87]), .Z(n1319) );
  NAND U1426 ( .A(n1280), .B(sreg[86]), .Z(n1284) );
  OR U1427 ( .A(n1282), .B(n1281), .Z(n1283) );
  AND U1428 ( .A(n1284), .B(n1283), .Z(n1318) );
  XOR U1429 ( .A(n1319), .B(n1318), .Z(c[87]) );
  NANDN U1430 ( .A(n1294), .B(n1293), .Z(n1298) );
  NAND U1431 ( .A(n1296), .B(n1295), .Z(n1297) );
  NAND U1432 ( .A(n1298), .B(n1297), .Z(n1349) );
  NAND U1433 ( .A(n1299), .B(n2666), .Z(n1301) );
  XNOR U1434 ( .A(n2695), .B(a[26]), .Z(n1336) );
  NAND U1435 ( .A(n1336), .B(n2665), .Z(n1300) );
  NAND U1436 ( .A(n1301), .B(n1300), .Z(n1326) );
  XNOR U1437 ( .A(b[3]), .B(a[30]), .Z(n1339) );
  NANDN U1438 ( .A(n1339), .B(n2561), .Z(n1304) );
  NANDN U1439 ( .A(n1302), .B(n2563), .Z(n1303) );
  AND U1440 ( .A(n1304), .B(n1303), .Z(n1327) );
  XNOR U1441 ( .A(n1326), .B(n1327), .Z(n1328) );
  NANDN U1442 ( .A(n246), .B(a[32]), .Z(n1305) );
  XOR U1443 ( .A(n2537), .B(n1305), .Z(n1307) );
  NANDN U1444 ( .A(b[0]), .B(a[31]), .Z(n1306) );
  AND U1445 ( .A(n1307), .B(n1306), .Z(n1332) );
  NANDN U1446 ( .A(n1308), .B(n2625), .Z(n1310) );
  XNOR U1447 ( .A(b[5]), .B(a[28]), .Z(n1345) );
  OR U1448 ( .A(n1345), .B(n2608), .Z(n1309) );
  NAND U1449 ( .A(n1310), .B(n1309), .Z(n1330) );
  NANDN U1450 ( .A(n2695), .B(a[24]), .Z(n1331) );
  XNOR U1451 ( .A(n1330), .B(n1331), .Z(n1333) );
  XOR U1452 ( .A(n1332), .B(n1333), .Z(n1329) );
  XOR U1453 ( .A(n1328), .B(n1329), .Z(n1348) );
  XOR U1454 ( .A(n1349), .B(n1348), .Z(n1350) );
  XNOR U1455 ( .A(n1351), .B(n1350), .Z(n1322) );
  NAND U1456 ( .A(n1312), .B(n1311), .Z(n1316) );
  NAND U1457 ( .A(n1314), .B(n1313), .Z(n1315) );
  NAND U1458 ( .A(n1316), .B(n1315), .Z(n1323) );
  XNOR U1459 ( .A(n1322), .B(n1323), .Z(n1324) );
  XNOR U1460 ( .A(n1325), .B(n1324), .Z(n1354) );
  XNOR U1461 ( .A(n1354), .B(sreg[88]), .Z(n1356) );
  NAND U1462 ( .A(n1317), .B(sreg[87]), .Z(n1321) );
  OR U1463 ( .A(n1319), .B(n1318), .Z(n1320) );
  AND U1464 ( .A(n1321), .B(n1320), .Z(n1355) );
  XOR U1465 ( .A(n1356), .B(n1355), .Z(c[88]) );
  NANDN U1466 ( .A(n1331), .B(n1330), .Z(n1335) );
  NAND U1467 ( .A(n1333), .B(n1332), .Z(n1334) );
  NAND U1468 ( .A(n1335), .B(n1334), .Z(n1386) );
  NAND U1469 ( .A(n1336), .B(n2666), .Z(n1338) );
  XNOR U1470 ( .A(n2695), .B(a[27]), .Z(n1373) );
  NAND U1471 ( .A(n1373), .B(n2665), .Z(n1337) );
  NAND U1472 ( .A(n1338), .B(n1337), .Z(n1363) );
  XNOR U1473 ( .A(b[3]), .B(a[31]), .Z(n1376) );
  NANDN U1474 ( .A(n1376), .B(n2561), .Z(n1341) );
  NANDN U1475 ( .A(n1339), .B(n2563), .Z(n1340) );
  AND U1476 ( .A(n1341), .B(n1340), .Z(n1364) );
  XNOR U1477 ( .A(n1363), .B(n1364), .Z(n1365) );
  NANDN U1478 ( .A(n246), .B(a[33]), .Z(n1342) );
  XOR U1479 ( .A(n2537), .B(n1342), .Z(n1344) );
  NANDN U1480 ( .A(b[0]), .B(a[32]), .Z(n1343) );
  AND U1481 ( .A(n1344), .B(n1343), .Z(n1369) );
  NANDN U1482 ( .A(n1345), .B(n2625), .Z(n1347) );
  XNOR U1483 ( .A(b[5]), .B(a[29]), .Z(n1382) );
  OR U1484 ( .A(n1382), .B(n2608), .Z(n1346) );
  NAND U1485 ( .A(n1347), .B(n1346), .Z(n1367) );
  NANDN U1486 ( .A(n2695), .B(a[25]), .Z(n1368) );
  XNOR U1487 ( .A(n1367), .B(n1368), .Z(n1370) );
  XOR U1488 ( .A(n1369), .B(n1370), .Z(n1366) );
  XOR U1489 ( .A(n1365), .B(n1366), .Z(n1385) );
  XOR U1490 ( .A(n1386), .B(n1385), .Z(n1387) );
  XNOR U1491 ( .A(n1388), .B(n1387), .Z(n1359) );
  NAND U1492 ( .A(n1349), .B(n1348), .Z(n1353) );
  NAND U1493 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U1494 ( .A(n1353), .B(n1352), .Z(n1360) );
  XNOR U1495 ( .A(n1359), .B(n1360), .Z(n1361) );
  XNOR U1496 ( .A(n1362), .B(n1361), .Z(n1391) );
  XNOR U1497 ( .A(n1391), .B(sreg[89]), .Z(n1393) );
  NAND U1498 ( .A(n1354), .B(sreg[88]), .Z(n1358) );
  OR U1499 ( .A(n1356), .B(n1355), .Z(n1357) );
  AND U1500 ( .A(n1358), .B(n1357), .Z(n1392) );
  XOR U1501 ( .A(n1393), .B(n1392), .Z(c[89]) );
  NANDN U1502 ( .A(n1368), .B(n1367), .Z(n1372) );
  NAND U1503 ( .A(n1370), .B(n1369), .Z(n1371) );
  NAND U1504 ( .A(n1372), .B(n1371), .Z(n1423) );
  NAND U1505 ( .A(n1373), .B(n2666), .Z(n1375) );
  XNOR U1506 ( .A(n2695), .B(a[28]), .Z(n1410) );
  NAND U1507 ( .A(n1410), .B(n2665), .Z(n1374) );
  NAND U1508 ( .A(n1375), .B(n1374), .Z(n1400) );
  XNOR U1509 ( .A(b[3]), .B(a[32]), .Z(n1413) );
  NANDN U1510 ( .A(n1413), .B(n2561), .Z(n1378) );
  NANDN U1511 ( .A(n1376), .B(n2563), .Z(n1377) );
  AND U1512 ( .A(n1378), .B(n1377), .Z(n1401) );
  XNOR U1513 ( .A(n1400), .B(n1401), .Z(n1402) );
  NANDN U1514 ( .A(n246), .B(a[34]), .Z(n1379) );
  XOR U1515 ( .A(n2537), .B(n1379), .Z(n1381) );
  NANDN U1516 ( .A(b[0]), .B(a[33]), .Z(n1380) );
  AND U1517 ( .A(n1381), .B(n1380), .Z(n1406) );
  NANDN U1518 ( .A(n1382), .B(n2625), .Z(n1384) );
  XNOR U1519 ( .A(b[5]), .B(a[30]), .Z(n1419) );
  OR U1520 ( .A(n1419), .B(n2608), .Z(n1383) );
  NAND U1521 ( .A(n1384), .B(n1383), .Z(n1404) );
  NANDN U1522 ( .A(n2695), .B(a[26]), .Z(n1405) );
  XNOR U1523 ( .A(n1404), .B(n1405), .Z(n1407) );
  XOR U1524 ( .A(n1406), .B(n1407), .Z(n1403) );
  XOR U1525 ( .A(n1402), .B(n1403), .Z(n1422) );
  XOR U1526 ( .A(n1423), .B(n1422), .Z(n1424) );
  XNOR U1527 ( .A(n1425), .B(n1424), .Z(n1396) );
  NAND U1528 ( .A(n1386), .B(n1385), .Z(n1390) );
  NAND U1529 ( .A(n1388), .B(n1387), .Z(n1389) );
  NAND U1530 ( .A(n1390), .B(n1389), .Z(n1397) );
  XNOR U1531 ( .A(n1396), .B(n1397), .Z(n1398) );
  XNOR U1532 ( .A(n1399), .B(n1398), .Z(n1428) );
  XNOR U1533 ( .A(n1428), .B(sreg[90]), .Z(n1430) );
  NAND U1534 ( .A(n1391), .B(sreg[89]), .Z(n1395) );
  OR U1535 ( .A(n1393), .B(n1392), .Z(n1394) );
  AND U1536 ( .A(n1395), .B(n1394), .Z(n1429) );
  XOR U1537 ( .A(n1430), .B(n1429), .Z(c[90]) );
  NANDN U1538 ( .A(n1405), .B(n1404), .Z(n1409) );
  NAND U1539 ( .A(n1407), .B(n1406), .Z(n1408) );
  NAND U1540 ( .A(n1409), .B(n1408), .Z(n1460) );
  NAND U1541 ( .A(n1410), .B(n2666), .Z(n1412) );
  XNOR U1542 ( .A(n2695), .B(a[29]), .Z(n1447) );
  NAND U1543 ( .A(n1447), .B(n2665), .Z(n1411) );
  NAND U1544 ( .A(n1412), .B(n1411), .Z(n1437) );
  XNOR U1545 ( .A(b[3]), .B(a[33]), .Z(n1450) );
  NANDN U1546 ( .A(n1450), .B(n2561), .Z(n1415) );
  NANDN U1547 ( .A(n1413), .B(n2563), .Z(n1414) );
  AND U1548 ( .A(n1415), .B(n1414), .Z(n1438) );
  XNOR U1549 ( .A(n1437), .B(n1438), .Z(n1439) );
  NANDN U1550 ( .A(n246), .B(a[35]), .Z(n1416) );
  XOR U1551 ( .A(n2537), .B(n1416), .Z(n1418) );
  NANDN U1552 ( .A(b[0]), .B(a[34]), .Z(n1417) );
  AND U1553 ( .A(n1418), .B(n1417), .Z(n1443) );
  NANDN U1554 ( .A(n1419), .B(n2625), .Z(n1421) );
  XNOR U1555 ( .A(b[5]), .B(a[31]), .Z(n1456) );
  OR U1556 ( .A(n1456), .B(n2608), .Z(n1420) );
  NAND U1557 ( .A(n1421), .B(n1420), .Z(n1441) );
  NANDN U1558 ( .A(n2695), .B(a[27]), .Z(n1442) );
  XNOR U1559 ( .A(n1441), .B(n1442), .Z(n1444) );
  XOR U1560 ( .A(n1443), .B(n1444), .Z(n1440) );
  XOR U1561 ( .A(n1439), .B(n1440), .Z(n1459) );
  XOR U1562 ( .A(n1460), .B(n1459), .Z(n1461) );
  XNOR U1563 ( .A(n1462), .B(n1461), .Z(n1433) );
  NAND U1564 ( .A(n1423), .B(n1422), .Z(n1427) );
  NAND U1565 ( .A(n1425), .B(n1424), .Z(n1426) );
  NAND U1566 ( .A(n1427), .B(n1426), .Z(n1434) );
  XNOR U1567 ( .A(n1433), .B(n1434), .Z(n1435) );
  XNOR U1568 ( .A(n1436), .B(n1435), .Z(n1465) );
  XNOR U1569 ( .A(n1465), .B(sreg[91]), .Z(n1467) );
  NAND U1570 ( .A(n1428), .B(sreg[90]), .Z(n1432) );
  OR U1571 ( .A(n1430), .B(n1429), .Z(n1431) );
  AND U1572 ( .A(n1432), .B(n1431), .Z(n1466) );
  XOR U1573 ( .A(n1467), .B(n1466), .Z(c[91]) );
  NANDN U1574 ( .A(n1442), .B(n1441), .Z(n1446) );
  NAND U1575 ( .A(n1444), .B(n1443), .Z(n1445) );
  NAND U1576 ( .A(n1446), .B(n1445), .Z(n1497) );
  NAND U1577 ( .A(n1447), .B(n2666), .Z(n1449) );
  XNOR U1578 ( .A(n2695), .B(a[30]), .Z(n1484) );
  NAND U1579 ( .A(n1484), .B(n2665), .Z(n1448) );
  NAND U1580 ( .A(n1449), .B(n1448), .Z(n1474) );
  XNOR U1581 ( .A(b[3]), .B(a[34]), .Z(n1487) );
  NANDN U1582 ( .A(n1487), .B(n2561), .Z(n1452) );
  NANDN U1583 ( .A(n1450), .B(n2563), .Z(n1451) );
  AND U1584 ( .A(n1452), .B(n1451), .Z(n1475) );
  XNOR U1585 ( .A(n1474), .B(n1475), .Z(n1476) );
  NANDN U1586 ( .A(n246), .B(a[36]), .Z(n1453) );
  XOR U1587 ( .A(n2537), .B(n1453), .Z(n1455) );
  NANDN U1588 ( .A(b[0]), .B(a[35]), .Z(n1454) );
  AND U1589 ( .A(n1455), .B(n1454), .Z(n1480) );
  NANDN U1590 ( .A(n1456), .B(n2625), .Z(n1458) );
  XNOR U1591 ( .A(b[5]), .B(a[32]), .Z(n1493) );
  OR U1592 ( .A(n1493), .B(n2608), .Z(n1457) );
  NAND U1593 ( .A(n1458), .B(n1457), .Z(n1478) );
  NANDN U1594 ( .A(n2695), .B(a[28]), .Z(n1479) );
  XNOR U1595 ( .A(n1478), .B(n1479), .Z(n1481) );
  XOR U1596 ( .A(n1480), .B(n1481), .Z(n1477) );
  XOR U1597 ( .A(n1476), .B(n1477), .Z(n1496) );
  XOR U1598 ( .A(n1497), .B(n1496), .Z(n1498) );
  XNOR U1599 ( .A(n1499), .B(n1498), .Z(n1470) );
  NAND U1600 ( .A(n1460), .B(n1459), .Z(n1464) );
  NAND U1601 ( .A(n1462), .B(n1461), .Z(n1463) );
  NAND U1602 ( .A(n1464), .B(n1463), .Z(n1471) );
  XNOR U1603 ( .A(n1470), .B(n1471), .Z(n1472) );
  XNOR U1604 ( .A(n1473), .B(n1472), .Z(n1502) );
  XNOR U1605 ( .A(n1502), .B(sreg[92]), .Z(n1504) );
  NAND U1606 ( .A(n1465), .B(sreg[91]), .Z(n1469) );
  OR U1607 ( .A(n1467), .B(n1466), .Z(n1468) );
  AND U1608 ( .A(n1469), .B(n1468), .Z(n1503) );
  XOR U1609 ( .A(n1504), .B(n1503), .Z(c[92]) );
  NANDN U1610 ( .A(n1479), .B(n1478), .Z(n1483) );
  NAND U1611 ( .A(n1481), .B(n1480), .Z(n1482) );
  NAND U1612 ( .A(n1483), .B(n1482), .Z(n1534) );
  NAND U1613 ( .A(n1484), .B(n2666), .Z(n1486) );
  XNOR U1614 ( .A(n2695), .B(a[31]), .Z(n1521) );
  NAND U1615 ( .A(n1521), .B(n2665), .Z(n1485) );
  NAND U1616 ( .A(n1486), .B(n1485), .Z(n1511) );
  XNOR U1617 ( .A(b[3]), .B(a[35]), .Z(n1524) );
  NANDN U1618 ( .A(n1524), .B(n2561), .Z(n1489) );
  NANDN U1619 ( .A(n1487), .B(n2563), .Z(n1488) );
  AND U1620 ( .A(n1489), .B(n1488), .Z(n1512) );
  XNOR U1621 ( .A(n1511), .B(n1512), .Z(n1513) );
  NANDN U1622 ( .A(n246), .B(a[37]), .Z(n1490) );
  XOR U1623 ( .A(n2537), .B(n1490), .Z(n1492) );
  NANDN U1624 ( .A(b[0]), .B(a[36]), .Z(n1491) );
  AND U1625 ( .A(n1492), .B(n1491), .Z(n1517) );
  NANDN U1626 ( .A(n1493), .B(n2625), .Z(n1495) );
  XNOR U1627 ( .A(b[5]), .B(a[33]), .Z(n1530) );
  OR U1628 ( .A(n1530), .B(n2608), .Z(n1494) );
  NAND U1629 ( .A(n1495), .B(n1494), .Z(n1515) );
  NANDN U1630 ( .A(n2695), .B(a[29]), .Z(n1516) );
  XNOR U1631 ( .A(n1515), .B(n1516), .Z(n1518) );
  XOR U1632 ( .A(n1517), .B(n1518), .Z(n1514) );
  XOR U1633 ( .A(n1513), .B(n1514), .Z(n1533) );
  XOR U1634 ( .A(n1534), .B(n1533), .Z(n1535) );
  XNOR U1635 ( .A(n1536), .B(n1535), .Z(n1507) );
  NAND U1636 ( .A(n1497), .B(n1496), .Z(n1501) );
  NAND U1637 ( .A(n1499), .B(n1498), .Z(n1500) );
  NAND U1638 ( .A(n1501), .B(n1500), .Z(n1508) );
  XNOR U1639 ( .A(n1507), .B(n1508), .Z(n1509) );
  XNOR U1640 ( .A(n1510), .B(n1509), .Z(n1539) );
  XNOR U1641 ( .A(n1539), .B(sreg[93]), .Z(n1541) );
  NAND U1642 ( .A(n1502), .B(sreg[92]), .Z(n1506) );
  OR U1643 ( .A(n1504), .B(n1503), .Z(n1505) );
  AND U1644 ( .A(n1506), .B(n1505), .Z(n1540) );
  XOR U1645 ( .A(n1541), .B(n1540), .Z(c[93]) );
  NANDN U1646 ( .A(n1516), .B(n1515), .Z(n1520) );
  NAND U1647 ( .A(n1518), .B(n1517), .Z(n1519) );
  NAND U1648 ( .A(n1520), .B(n1519), .Z(n1571) );
  NAND U1649 ( .A(n1521), .B(n2666), .Z(n1523) );
  XNOR U1650 ( .A(n2695), .B(a[32]), .Z(n1558) );
  NAND U1651 ( .A(n1558), .B(n2665), .Z(n1522) );
  NAND U1652 ( .A(n1523), .B(n1522), .Z(n1548) );
  XNOR U1653 ( .A(b[3]), .B(a[36]), .Z(n1561) );
  NANDN U1654 ( .A(n1561), .B(n2561), .Z(n1526) );
  NANDN U1655 ( .A(n1524), .B(n2563), .Z(n1525) );
  AND U1656 ( .A(n1526), .B(n1525), .Z(n1549) );
  XNOR U1657 ( .A(n1548), .B(n1549), .Z(n1550) );
  NANDN U1658 ( .A(n246), .B(a[38]), .Z(n1527) );
  XOR U1659 ( .A(n2537), .B(n1527), .Z(n1529) );
  NANDN U1660 ( .A(b[0]), .B(a[37]), .Z(n1528) );
  AND U1661 ( .A(n1529), .B(n1528), .Z(n1554) );
  NANDN U1662 ( .A(n1530), .B(n2625), .Z(n1532) );
  XNOR U1663 ( .A(b[5]), .B(a[34]), .Z(n1567) );
  OR U1664 ( .A(n1567), .B(n2608), .Z(n1531) );
  NAND U1665 ( .A(n1532), .B(n1531), .Z(n1552) );
  NANDN U1666 ( .A(n2695), .B(a[30]), .Z(n1553) );
  XNOR U1667 ( .A(n1552), .B(n1553), .Z(n1555) );
  XOR U1668 ( .A(n1554), .B(n1555), .Z(n1551) );
  XOR U1669 ( .A(n1550), .B(n1551), .Z(n1570) );
  XOR U1670 ( .A(n1571), .B(n1570), .Z(n1572) );
  XNOR U1671 ( .A(n1573), .B(n1572), .Z(n1544) );
  NAND U1672 ( .A(n1534), .B(n1533), .Z(n1538) );
  NAND U1673 ( .A(n1536), .B(n1535), .Z(n1537) );
  NAND U1674 ( .A(n1538), .B(n1537), .Z(n1545) );
  XNOR U1675 ( .A(n1544), .B(n1545), .Z(n1546) );
  XNOR U1676 ( .A(n1547), .B(n1546), .Z(n1576) );
  XNOR U1677 ( .A(n1576), .B(sreg[94]), .Z(n1578) );
  NAND U1678 ( .A(n1539), .B(sreg[93]), .Z(n1543) );
  OR U1679 ( .A(n1541), .B(n1540), .Z(n1542) );
  AND U1680 ( .A(n1543), .B(n1542), .Z(n1577) );
  XOR U1681 ( .A(n1578), .B(n1577), .Z(c[94]) );
  NANDN U1682 ( .A(n1553), .B(n1552), .Z(n1557) );
  NAND U1683 ( .A(n1555), .B(n1554), .Z(n1556) );
  NAND U1684 ( .A(n1557), .B(n1556), .Z(n1608) );
  NAND U1685 ( .A(n1558), .B(n2666), .Z(n1560) );
  XNOR U1686 ( .A(n2695), .B(a[33]), .Z(n1595) );
  NAND U1687 ( .A(n1595), .B(n2665), .Z(n1559) );
  NAND U1688 ( .A(n1560), .B(n1559), .Z(n1585) );
  XNOR U1689 ( .A(b[3]), .B(a[37]), .Z(n1598) );
  NANDN U1690 ( .A(n1598), .B(n2561), .Z(n1563) );
  NANDN U1691 ( .A(n1561), .B(n2563), .Z(n1562) );
  AND U1692 ( .A(n1563), .B(n1562), .Z(n1586) );
  XNOR U1693 ( .A(n1585), .B(n1586), .Z(n1587) );
  NANDN U1694 ( .A(n246), .B(a[39]), .Z(n1564) );
  XOR U1695 ( .A(n2537), .B(n1564), .Z(n1566) );
  NANDN U1696 ( .A(b[0]), .B(a[38]), .Z(n1565) );
  AND U1697 ( .A(n1566), .B(n1565), .Z(n1591) );
  NANDN U1698 ( .A(n1567), .B(n2625), .Z(n1569) );
  XNOR U1699 ( .A(b[5]), .B(a[35]), .Z(n1604) );
  OR U1700 ( .A(n1604), .B(n2608), .Z(n1568) );
  NAND U1701 ( .A(n1569), .B(n1568), .Z(n1589) );
  NANDN U1702 ( .A(n2695), .B(a[31]), .Z(n1590) );
  XNOR U1703 ( .A(n1589), .B(n1590), .Z(n1592) );
  XOR U1704 ( .A(n1591), .B(n1592), .Z(n1588) );
  XOR U1705 ( .A(n1587), .B(n1588), .Z(n1607) );
  XOR U1706 ( .A(n1608), .B(n1607), .Z(n1609) );
  XNOR U1707 ( .A(n1610), .B(n1609), .Z(n1581) );
  NAND U1708 ( .A(n1571), .B(n1570), .Z(n1575) );
  NAND U1709 ( .A(n1573), .B(n1572), .Z(n1574) );
  NAND U1710 ( .A(n1575), .B(n1574), .Z(n1582) );
  XNOR U1711 ( .A(n1581), .B(n1582), .Z(n1583) );
  XNOR U1712 ( .A(n1584), .B(n1583), .Z(n1613) );
  XNOR U1713 ( .A(n1613), .B(sreg[95]), .Z(n1615) );
  NAND U1714 ( .A(n1576), .B(sreg[94]), .Z(n1580) );
  OR U1715 ( .A(n1578), .B(n1577), .Z(n1579) );
  AND U1716 ( .A(n1580), .B(n1579), .Z(n1614) );
  XOR U1717 ( .A(n1615), .B(n1614), .Z(c[95]) );
  NANDN U1718 ( .A(n1590), .B(n1589), .Z(n1594) );
  NAND U1719 ( .A(n1592), .B(n1591), .Z(n1593) );
  NAND U1720 ( .A(n1594), .B(n1593), .Z(n1645) );
  NAND U1721 ( .A(n1595), .B(n2666), .Z(n1597) );
  XNOR U1722 ( .A(n2695), .B(a[34]), .Z(n1632) );
  NAND U1723 ( .A(n1632), .B(n2665), .Z(n1596) );
  NAND U1724 ( .A(n1597), .B(n1596), .Z(n1622) );
  XNOR U1725 ( .A(b[3]), .B(a[38]), .Z(n1635) );
  NANDN U1726 ( .A(n1635), .B(n2561), .Z(n1600) );
  NANDN U1727 ( .A(n1598), .B(n2563), .Z(n1599) );
  AND U1728 ( .A(n1600), .B(n1599), .Z(n1623) );
  XNOR U1729 ( .A(n1622), .B(n1623), .Z(n1624) );
  NANDN U1730 ( .A(n246), .B(a[40]), .Z(n1601) );
  XOR U1731 ( .A(n2537), .B(n1601), .Z(n1603) );
  NANDN U1732 ( .A(b[0]), .B(a[39]), .Z(n1602) );
  AND U1733 ( .A(n1603), .B(n1602), .Z(n1628) );
  NANDN U1734 ( .A(n1604), .B(n2625), .Z(n1606) );
  XNOR U1735 ( .A(b[5]), .B(a[36]), .Z(n1641) );
  OR U1736 ( .A(n1641), .B(n2608), .Z(n1605) );
  NAND U1737 ( .A(n1606), .B(n1605), .Z(n1626) );
  NANDN U1738 ( .A(n2695), .B(a[32]), .Z(n1627) );
  XNOR U1739 ( .A(n1626), .B(n1627), .Z(n1629) );
  XOR U1740 ( .A(n1628), .B(n1629), .Z(n1625) );
  XOR U1741 ( .A(n1624), .B(n1625), .Z(n1644) );
  XOR U1742 ( .A(n1645), .B(n1644), .Z(n1646) );
  XNOR U1743 ( .A(n1647), .B(n1646), .Z(n1618) );
  NAND U1744 ( .A(n1608), .B(n1607), .Z(n1612) );
  NAND U1745 ( .A(n1610), .B(n1609), .Z(n1611) );
  NAND U1746 ( .A(n1612), .B(n1611), .Z(n1619) );
  XNOR U1747 ( .A(n1618), .B(n1619), .Z(n1620) );
  XNOR U1748 ( .A(n1621), .B(n1620), .Z(n1650) );
  XNOR U1749 ( .A(n1650), .B(sreg[96]), .Z(n1652) );
  NAND U1750 ( .A(n1613), .B(sreg[95]), .Z(n1617) );
  OR U1751 ( .A(n1615), .B(n1614), .Z(n1616) );
  AND U1752 ( .A(n1617), .B(n1616), .Z(n1651) );
  XOR U1753 ( .A(n1652), .B(n1651), .Z(c[96]) );
  NANDN U1754 ( .A(n1627), .B(n1626), .Z(n1631) );
  NAND U1755 ( .A(n1629), .B(n1628), .Z(n1630) );
  NAND U1756 ( .A(n1631), .B(n1630), .Z(n1682) );
  NAND U1757 ( .A(n1632), .B(n2666), .Z(n1634) );
  XNOR U1758 ( .A(n2695), .B(a[35]), .Z(n1669) );
  NAND U1759 ( .A(n1669), .B(n2665), .Z(n1633) );
  NAND U1760 ( .A(n1634), .B(n1633), .Z(n1659) );
  XNOR U1761 ( .A(b[3]), .B(a[39]), .Z(n1672) );
  NANDN U1762 ( .A(n1672), .B(n2561), .Z(n1637) );
  NANDN U1763 ( .A(n1635), .B(n2563), .Z(n1636) );
  AND U1764 ( .A(n1637), .B(n1636), .Z(n1660) );
  XNOR U1765 ( .A(n1659), .B(n1660), .Z(n1661) );
  NANDN U1766 ( .A(n246), .B(a[41]), .Z(n1638) );
  XOR U1767 ( .A(n2537), .B(n1638), .Z(n1640) );
  NANDN U1768 ( .A(b[0]), .B(a[40]), .Z(n1639) );
  AND U1769 ( .A(n1640), .B(n1639), .Z(n1665) );
  NANDN U1770 ( .A(n1641), .B(n2625), .Z(n1643) );
  XNOR U1771 ( .A(b[5]), .B(a[37]), .Z(n1678) );
  OR U1772 ( .A(n1678), .B(n2608), .Z(n1642) );
  NAND U1773 ( .A(n1643), .B(n1642), .Z(n1663) );
  NANDN U1774 ( .A(n2695), .B(a[33]), .Z(n1664) );
  XNOR U1775 ( .A(n1663), .B(n1664), .Z(n1666) );
  XOR U1776 ( .A(n1665), .B(n1666), .Z(n1662) );
  XOR U1777 ( .A(n1661), .B(n1662), .Z(n1681) );
  XOR U1778 ( .A(n1682), .B(n1681), .Z(n1683) );
  XNOR U1779 ( .A(n1684), .B(n1683), .Z(n1655) );
  NAND U1780 ( .A(n1645), .B(n1644), .Z(n1649) );
  NAND U1781 ( .A(n1647), .B(n1646), .Z(n1648) );
  NAND U1782 ( .A(n1649), .B(n1648), .Z(n1656) );
  XNOR U1783 ( .A(n1655), .B(n1656), .Z(n1657) );
  XNOR U1784 ( .A(n1658), .B(n1657), .Z(n1687) );
  XNOR U1785 ( .A(n1687), .B(sreg[97]), .Z(n1689) );
  NAND U1786 ( .A(n1650), .B(sreg[96]), .Z(n1654) );
  OR U1787 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U1788 ( .A(n1654), .B(n1653), .Z(n1688) );
  XOR U1789 ( .A(n1689), .B(n1688), .Z(c[97]) );
  NANDN U1790 ( .A(n1664), .B(n1663), .Z(n1668) );
  NAND U1791 ( .A(n1666), .B(n1665), .Z(n1667) );
  NAND U1792 ( .A(n1668), .B(n1667), .Z(n1719) );
  NAND U1793 ( .A(n1669), .B(n2666), .Z(n1671) );
  XNOR U1794 ( .A(n2695), .B(a[36]), .Z(n1706) );
  NAND U1795 ( .A(n1706), .B(n2665), .Z(n1670) );
  NAND U1796 ( .A(n1671), .B(n1670), .Z(n1696) );
  XNOR U1797 ( .A(b[3]), .B(a[40]), .Z(n1709) );
  NANDN U1798 ( .A(n1709), .B(n2561), .Z(n1674) );
  NANDN U1799 ( .A(n1672), .B(n2563), .Z(n1673) );
  AND U1800 ( .A(n1674), .B(n1673), .Z(n1697) );
  XNOR U1801 ( .A(n1696), .B(n1697), .Z(n1698) );
  NANDN U1802 ( .A(n246), .B(a[42]), .Z(n1675) );
  XOR U1803 ( .A(n2537), .B(n1675), .Z(n1677) );
  NANDN U1804 ( .A(b[0]), .B(a[41]), .Z(n1676) );
  AND U1805 ( .A(n1677), .B(n1676), .Z(n1702) );
  NANDN U1806 ( .A(n1678), .B(n2625), .Z(n1680) );
  XNOR U1807 ( .A(b[5]), .B(a[38]), .Z(n1715) );
  OR U1808 ( .A(n1715), .B(n2608), .Z(n1679) );
  NAND U1809 ( .A(n1680), .B(n1679), .Z(n1700) );
  NANDN U1810 ( .A(n2695), .B(a[34]), .Z(n1701) );
  XNOR U1811 ( .A(n1700), .B(n1701), .Z(n1703) );
  XOR U1812 ( .A(n1702), .B(n1703), .Z(n1699) );
  XOR U1813 ( .A(n1698), .B(n1699), .Z(n1718) );
  XOR U1814 ( .A(n1719), .B(n1718), .Z(n1720) );
  XNOR U1815 ( .A(n1721), .B(n1720), .Z(n1692) );
  NAND U1816 ( .A(n1682), .B(n1681), .Z(n1686) );
  NAND U1817 ( .A(n1684), .B(n1683), .Z(n1685) );
  NAND U1818 ( .A(n1686), .B(n1685), .Z(n1693) );
  XNOR U1819 ( .A(n1692), .B(n1693), .Z(n1694) );
  XNOR U1820 ( .A(n1695), .B(n1694), .Z(n1724) );
  XNOR U1821 ( .A(n1724), .B(sreg[98]), .Z(n1726) );
  NAND U1822 ( .A(n1687), .B(sreg[97]), .Z(n1691) );
  OR U1823 ( .A(n1689), .B(n1688), .Z(n1690) );
  AND U1824 ( .A(n1691), .B(n1690), .Z(n1725) );
  XOR U1825 ( .A(n1726), .B(n1725), .Z(c[98]) );
  NANDN U1826 ( .A(n1701), .B(n1700), .Z(n1705) );
  NAND U1827 ( .A(n1703), .B(n1702), .Z(n1704) );
  NAND U1828 ( .A(n1705), .B(n1704), .Z(n1756) );
  NAND U1829 ( .A(n1706), .B(n2666), .Z(n1708) );
  XNOR U1830 ( .A(n2695), .B(a[37]), .Z(n1743) );
  NAND U1831 ( .A(n1743), .B(n2665), .Z(n1707) );
  NAND U1832 ( .A(n1708), .B(n1707), .Z(n1733) );
  XNOR U1833 ( .A(b[3]), .B(a[41]), .Z(n1746) );
  NANDN U1834 ( .A(n1746), .B(n2561), .Z(n1711) );
  NANDN U1835 ( .A(n1709), .B(n2563), .Z(n1710) );
  AND U1836 ( .A(n1711), .B(n1710), .Z(n1734) );
  XNOR U1837 ( .A(n1733), .B(n1734), .Z(n1735) );
  NANDN U1838 ( .A(n246), .B(a[43]), .Z(n1712) );
  XOR U1839 ( .A(n2537), .B(n1712), .Z(n1714) );
  NANDN U1840 ( .A(b[0]), .B(a[42]), .Z(n1713) );
  AND U1841 ( .A(n1714), .B(n1713), .Z(n1739) );
  NANDN U1842 ( .A(n1715), .B(n2625), .Z(n1717) );
  XNOR U1843 ( .A(b[5]), .B(a[39]), .Z(n1752) );
  OR U1844 ( .A(n1752), .B(n2608), .Z(n1716) );
  NAND U1845 ( .A(n1717), .B(n1716), .Z(n1737) );
  NANDN U1846 ( .A(n2695), .B(a[35]), .Z(n1738) );
  XNOR U1847 ( .A(n1737), .B(n1738), .Z(n1740) );
  XOR U1848 ( .A(n1739), .B(n1740), .Z(n1736) );
  XOR U1849 ( .A(n1735), .B(n1736), .Z(n1755) );
  XOR U1850 ( .A(n1756), .B(n1755), .Z(n1757) );
  XNOR U1851 ( .A(n1758), .B(n1757), .Z(n1729) );
  NAND U1852 ( .A(n1719), .B(n1718), .Z(n1723) );
  NAND U1853 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U1854 ( .A(n1723), .B(n1722), .Z(n1730) );
  XNOR U1855 ( .A(n1729), .B(n1730), .Z(n1731) );
  XNOR U1856 ( .A(n1732), .B(n1731), .Z(n1761) );
  XNOR U1857 ( .A(n1761), .B(sreg[99]), .Z(n1763) );
  NAND U1858 ( .A(n1724), .B(sreg[98]), .Z(n1728) );
  OR U1859 ( .A(n1726), .B(n1725), .Z(n1727) );
  AND U1860 ( .A(n1728), .B(n1727), .Z(n1762) );
  XOR U1861 ( .A(n1763), .B(n1762), .Z(c[99]) );
  NANDN U1862 ( .A(n1738), .B(n1737), .Z(n1742) );
  NAND U1863 ( .A(n1740), .B(n1739), .Z(n1741) );
  NAND U1864 ( .A(n1742), .B(n1741), .Z(n1793) );
  NAND U1865 ( .A(n1743), .B(n2666), .Z(n1745) );
  XNOR U1866 ( .A(n2695), .B(a[38]), .Z(n1780) );
  NAND U1867 ( .A(n1780), .B(n2665), .Z(n1744) );
  NAND U1868 ( .A(n1745), .B(n1744), .Z(n1770) );
  XNOR U1869 ( .A(b[3]), .B(a[42]), .Z(n1783) );
  NANDN U1870 ( .A(n1783), .B(n2561), .Z(n1748) );
  NANDN U1871 ( .A(n1746), .B(n2563), .Z(n1747) );
  AND U1872 ( .A(n1748), .B(n1747), .Z(n1771) );
  XNOR U1873 ( .A(n1770), .B(n1771), .Z(n1772) );
  NANDN U1874 ( .A(n246), .B(a[44]), .Z(n1749) );
  XOR U1875 ( .A(n2537), .B(n1749), .Z(n1751) );
  NANDN U1876 ( .A(b[0]), .B(a[43]), .Z(n1750) );
  AND U1877 ( .A(n1751), .B(n1750), .Z(n1776) );
  NANDN U1878 ( .A(n1752), .B(n2625), .Z(n1754) );
  XNOR U1879 ( .A(b[5]), .B(a[40]), .Z(n1789) );
  OR U1880 ( .A(n1789), .B(n2608), .Z(n1753) );
  NAND U1881 ( .A(n1754), .B(n1753), .Z(n1774) );
  NANDN U1882 ( .A(n2695), .B(a[36]), .Z(n1775) );
  XNOR U1883 ( .A(n1774), .B(n1775), .Z(n1777) );
  XOR U1884 ( .A(n1776), .B(n1777), .Z(n1773) );
  XOR U1885 ( .A(n1772), .B(n1773), .Z(n1792) );
  XOR U1886 ( .A(n1793), .B(n1792), .Z(n1794) );
  XNOR U1887 ( .A(n1795), .B(n1794), .Z(n1766) );
  NAND U1888 ( .A(n1756), .B(n1755), .Z(n1760) );
  NAND U1889 ( .A(n1758), .B(n1757), .Z(n1759) );
  NAND U1890 ( .A(n1760), .B(n1759), .Z(n1767) );
  XNOR U1891 ( .A(n1766), .B(n1767), .Z(n1768) );
  XNOR U1892 ( .A(n1769), .B(n1768), .Z(n1798) );
  XNOR U1893 ( .A(n1798), .B(sreg[100]), .Z(n1800) );
  NAND U1894 ( .A(n1761), .B(sreg[99]), .Z(n1765) );
  OR U1895 ( .A(n1763), .B(n1762), .Z(n1764) );
  AND U1896 ( .A(n1765), .B(n1764), .Z(n1799) );
  XOR U1897 ( .A(n1800), .B(n1799), .Z(c[100]) );
  NANDN U1898 ( .A(n1775), .B(n1774), .Z(n1779) );
  NAND U1899 ( .A(n1777), .B(n1776), .Z(n1778) );
  NAND U1900 ( .A(n1779), .B(n1778), .Z(n1830) );
  NAND U1901 ( .A(n1780), .B(n2666), .Z(n1782) );
  XNOR U1902 ( .A(n2695), .B(a[39]), .Z(n1817) );
  NAND U1903 ( .A(n1817), .B(n2665), .Z(n1781) );
  NAND U1904 ( .A(n1782), .B(n1781), .Z(n1807) );
  XNOR U1905 ( .A(b[3]), .B(a[43]), .Z(n1820) );
  NANDN U1906 ( .A(n1820), .B(n2561), .Z(n1785) );
  NANDN U1907 ( .A(n1783), .B(n2563), .Z(n1784) );
  AND U1908 ( .A(n1785), .B(n1784), .Z(n1808) );
  XNOR U1909 ( .A(n1807), .B(n1808), .Z(n1809) );
  NANDN U1910 ( .A(n246), .B(a[45]), .Z(n1786) );
  XOR U1911 ( .A(n2537), .B(n1786), .Z(n1788) );
  NANDN U1912 ( .A(b[0]), .B(a[44]), .Z(n1787) );
  AND U1913 ( .A(n1788), .B(n1787), .Z(n1813) );
  NANDN U1914 ( .A(n1789), .B(n2625), .Z(n1791) );
  XNOR U1915 ( .A(b[5]), .B(a[41]), .Z(n1826) );
  OR U1916 ( .A(n1826), .B(n2608), .Z(n1790) );
  NAND U1917 ( .A(n1791), .B(n1790), .Z(n1811) );
  NANDN U1918 ( .A(n2695), .B(a[37]), .Z(n1812) );
  XNOR U1919 ( .A(n1811), .B(n1812), .Z(n1814) );
  XOR U1920 ( .A(n1813), .B(n1814), .Z(n1810) );
  XOR U1921 ( .A(n1809), .B(n1810), .Z(n1829) );
  XOR U1922 ( .A(n1830), .B(n1829), .Z(n1831) );
  XNOR U1923 ( .A(n1832), .B(n1831), .Z(n1803) );
  NAND U1924 ( .A(n1793), .B(n1792), .Z(n1797) );
  NAND U1925 ( .A(n1795), .B(n1794), .Z(n1796) );
  NAND U1926 ( .A(n1797), .B(n1796), .Z(n1804) );
  XNOR U1927 ( .A(n1803), .B(n1804), .Z(n1805) );
  XNOR U1928 ( .A(n1806), .B(n1805), .Z(n1835) );
  XNOR U1929 ( .A(n1835), .B(sreg[101]), .Z(n1837) );
  NAND U1930 ( .A(n1798), .B(sreg[100]), .Z(n1802) );
  OR U1931 ( .A(n1800), .B(n1799), .Z(n1801) );
  AND U1932 ( .A(n1802), .B(n1801), .Z(n1836) );
  XOR U1933 ( .A(n1837), .B(n1836), .Z(c[101]) );
  NANDN U1934 ( .A(n1812), .B(n1811), .Z(n1816) );
  NAND U1935 ( .A(n1814), .B(n1813), .Z(n1815) );
  NAND U1936 ( .A(n1816), .B(n1815), .Z(n1867) );
  NAND U1937 ( .A(n1817), .B(n2666), .Z(n1819) );
  XNOR U1938 ( .A(n2695), .B(a[40]), .Z(n1854) );
  NAND U1939 ( .A(n1854), .B(n2665), .Z(n1818) );
  NAND U1940 ( .A(n1819), .B(n1818), .Z(n1844) );
  XNOR U1941 ( .A(b[3]), .B(a[44]), .Z(n1857) );
  NANDN U1942 ( .A(n1857), .B(n2561), .Z(n1822) );
  NANDN U1943 ( .A(n1820), .B(n2563), .Z(n1821) );
  AND U1944 ( .A(n1822), .B(n1821), .Z(n1845) );
  XNOR U1945 ( .A(n1844), .B(n1845), .Z(n1846) );
  NANDN U1946 ( .A(n246), .B(a[46]), .Z(n1823) );
  XOR U1947 ( .A(n2537), .B(n1823), .Z(n1825) );
  NANDN U1948 ( .A(b[0]), .B(a[45]), .Z(n1824) );
  AND U1949 ( .A(n1825), .B(n1824), .Z(n1850) );
  NANDN U1950 ( .A(n1826), .B(n2625), .Z(n1828) );
  XNOR U1951 ( .A(b[5]), .B(a[42]), .Z(n1863) );
  OR U1952 ( .A(n1863), .B(n2608), .Z(n1827) );
  NAND U1953 ( .A(n1828), .B(n1827), .Z(n1848) );
  NANDN U1954 ( .A(n2695), .B(a[38]), .Z(n1849) );
  XNOR U1955 ( .A(n1848), .B(n1849), .Z(n1851) );
  XOR U1956 ( .A(n1850), .B(n1851), .Z(n1847) );
  XOR U1957 ( .A(n1846), .B(n1847), .Z(n1866) );
  XOR U1958 ( .A(n1867), .B(n1866), .Z(n1868) );
  XNOR U1959 ( .A(n1869), .B(n1868), .Z(n1840) );
  NAND U1960 ( .A(n1830), .B(n1829), .Z(n1834) );
  NAND U1961 ( .A(n1832), .B(n1831), .Z(n1833) );
  NAND U1962 ( .A(n1834), .B(n1833), .Z(n1841) );
  XNOR U1963 ( .A(n1840), .B(n1841), .Z(n1842) );
  XNOR U1964 ( .A(n1843), .B(n1842), .Z(n1872) );
  XNOR U1965 ( .A(n1872), .B(sreg[102]), .Z(n1874) );
  NAND U1966 ( .A(n1835), .B(sreg[101]), .Z(n1839) );
  OR U1967 ( .A(n1837), .B(n1836), .Z(n1838) );
  AND U1968 ( .A(n1839), .B(n1838), .Z(n1873) );
  XOR U1969 ( .A(n1874), .B(n1873), .Z(c[102]) );
  NANDN U1970 ( .A(n1849), .B(n1848), .Z(n1853) );
  NAND U1971 ( .A(n1851), .B(n1850), .Z(n1852) );
  NAND U1972 ( .A(n1853), .B(n1852), .Z(n1904) );
  NAND U1973 ( .A(n1854), .B(n2666), .Z(n1856) );
  XNOR U1974 ( .A(n2695), .B(a[41]), .Z(n1891) );
  NAND U1975 ( .A(n1891), .B(n2665), .Z(n1855) );
  NAND U1976 ( .A(n1856), .B(n1855), .Z(n1881) );
  XNOR U1977 ( .A(b[3]), .B(a[45]), .Z(n1894) );
  NANDN U1978 ( .A(n1894), .B(n2561), .Z(n1859) );
  NANDN U1979 ( .A(n1857), .B(n2563), .Z(n1858) );
  AND U1980 ( .A(n1859), .B(n1858), .Z(n1882) );
  XNOR U1981 ( .A(n1881), .B(n1882), .Z(n1883) );
  NANDN U1982 ( .A(n246), .B(a[47]), .Z(n1860) );
  XOR U1983 ( .A(n2537), .B(n1860), .Z(n1862) );
  NANDN U1984 ( .A(b[0]), .B(a[46]), .Z(n1861) );
  AND U1985 ( .A(n1862), .B(n1861), .Z(n1887) );
  NANDN U1986 ( .A(n1863), .B(n2625), .Z(n1865) );
  XNOR U1987 ( .A(b[5]), .B(a[43]), .Z(n1900) );
  OR U1988 ( .A(n1900), .B(n2608), .Z(n1864) );
  NAND U1989 ( .A(n1865), .B(n1864), .Z(n1885) );
  NANDN U1990 ( .A(n2695), .B(a[39]), .Z(n1886) );
  XNOR U1991 ( .A(n1885), .B(n1886), .Z(n1888) );
  XOR U1992 ( .A(n1887), .B(n1888), .Z(n1884) );
  XOR U1993 ( .A(n1883), .B(n1884), .Z(n1903) );
  XOR U1994 ( .A(n1904), .B(n1903), .Z(n1905) );
  XNOR U1995 ( .A(n1906), .B(n1905), .Z(n1877) );
  NAND U1996 ( .A(n1867), .B(n1866), .Z(n1871) );
  NAND U1997 ( .A(n1869), .B(n1868), .Z(n1870) );
  NAND U1998 ( .A(n1871), .B(n1870), .Z(n1878) );
  XNOR U1999 ( .A(n1877), .B(n1878), .Z(n1879) );
  XNOR U2000 ( .A(n1880), .B(n1879), .Z(n1909) );
  XNOR U2001 ( .A(n1909), .B(sreg[103]), .Z(n1911) );
  NAND U2002 ( .A(n1872), .B(sreg[102]), .Z(n1876) );
  OR U2003 ( .A(n1874), .B(n1873), .Z(n1875) );
  AND U2004 ( .A(n1876), .B(n1875), .Z(n1910) );
  XOR U2005 ( .A(n1911), .B(n1910), .Z(c[103]) );
  NANDN U2006 ( .A(n1886), .B(n1885), .Z(n1890) );
  NAND U2007 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U2008 ( .A(n1890), .B(n1889), .Z(n1941) );
  NAND U2009 ( .A(n1891), .B(n2666), .Z(n1893) );
  XNOR U2010 ( .A(n2695), .B(a[42]), .Z(n1928) );
  NAND U2011 ( .A(n1928), .B(n2665), .Z(n1892) );
  NAND U2012 ( .A(n1893), .B(n1892), .Z(n1918) );
  XNOR U2013 ( .A(b[3]), .B(a[46]), .Z(n1931) );
  NANDN U2014 ( .A(n1931), .B(n2561), .Z(n1896) );
  NANDN U2015 ( .A(n1894), .B(n2563), .Z(n1895) );
  AND U2016 ( .A(n1896), .B(n1895), .Z(n1919) );
  XNOR U2017 ( .A(n1918), .B(n1919), .Z(n1920) );
  NANDN U2018 ( .A(n246), .B(a[48]), .Z(n1897) );
  XOR U2019 ( .A(n2537), .B(n1897), .Z(n1899) );
  NANDN U2020 ( .A(b[0]), .B(a[47]), .Z(n1898) );
  AND U2021 ( .A(n1899), .B(n1898), .Z(n1924) );
  NANDN U2022 ( .A(n1900), .B(n2625), .Z(n1902) );
  XNOR U2023 ( .A(b[5]), .B(a[44]), .Z(n1937) );
  OR U2024 ( .A(n1937), .B(n2608), .Z(n1901) );
  NAND U2025 ( .A(n1902), .B(n1901), .Z(n1922) );
  NANDN U2026 ( .A(n2695), .B(a[40]), .Z(n1923) );
  XNOR U2027 ( .A(n1922), .B(n1923), .Z(n1925) );
  XOR U2028 ( .A(n1924), .B(n1925), .Z(n1921) );
  XOR U2029 ( .A(n1920), .B(n1921), .Z(n1940) );
  XOR U2030 ( .A(n1941), .B(n1940), .Z(n1942) );
  XNOR U2031 ( .A(n1943), .B(n1942), .Z(n1914) );
  NAND U2032 ( .A(n1904), .B(n1903), .Z(n1908) );
  NAND U2033 ( .A(n1906), .B(n1905), .Z(n1907) );
  NAND U2034 ( .A(n1908), .B(n1907), .Z(n1915) );
  XNOR U2035 ( .A(n1914), .B(n1915), .Z(n1916) );
  XNOR U2036 ( .A(n1917), .B(n1916), .Z(n1946) );
  XNOR U2037 ( .A(n1946), .B(sreg[104]), .Z(n1948) );
  NAND U2038 ( .A(n1909), .B(sreg[103]), .Z(n1913) );
  OR U2039 ( .A(n1911), .B(n1910), .Z(n1912) );
  AND U2040 ( .A(n1913), .B(n1912), .Z(n1947) );
  XOR U2041 ( .A(n1948), .B(n1947), .Z(c[104]) );
  NANDN U2042 ( .A(n1923), .B(n1922), .Z(n1927) );
  NAND U2043 ( .A(n1925), .B(n1924), .Z(n1926) );
  NAND U2044 ( .A(n1927), .B(n1926), .Z(n1978) );
  NAND U2045 ( .A(n1928), .B(n2666), .Z(n1930) );
  XNOR U2046 ( .A(n2695), .B(a[43]), .Z(n1965) );
  NAND U2047 ( .A(n1965), .B(n2665), .Z(n1929) );
  NAND U2048 ( .A(n1930), .B(n1929), .Z(n1955) );
  XNOR U2049 ( .A(b[3]), .B(a[47]), .Z(n1968) );
  NANDN U2050 ( .A(n1968), .B(n2561), .Z(n1933) );
  NANDN U2051 ( .A(n1931), .B(n2563), .Z(n1932) );
  AND U2052 ( .A(n1933), .B(n1932), .Z(n1956) );
  XNOR U2053 ( .A(n1955), .B(n1956), .Z(n1957) );
  NANDN U2054 ( .A(n246), .B(a[49]), .Z(n1934) );
  XOR U2055 ( .A(n2537), .B(n1934), .Z(n1936) );
  NANDN U2056 ( .A(b[0]), .B(a[48]), .Z(n1935) );
  AND U2057 ( .A(n1936), .B(n1935), .Z(n1961) );
  NANDN U2058 ( .A(n1937), .B(n2625), .Z(n1939) );
  XNOR U2059 ( .A(b[5]), .B(a[45]), .Z(n1974) );
  OR U2060 ( .A(n1974), .B(n2608), .Z(n1938) );
  NAND U2061 ( .A(n1939), .B(n1938), .Z(n1959) );
  NANDN U2062 ( .A(n2695), .B(a[41]), .Z(n1960) );
  XNOR U2063 ( .A(n1959), .B(n1960), .Z(n1962) );
  XOR U2064 ( .A(n1961), .B(n1962), .Z(n1958) );
  XOR U2065 ( .A(n1957), .B(n1958), .Z(n1977) );
  XOR U2066 ( .A(n1978), .B(n1977), .Z(n1979) );
  XNOR U2067 ( .A(n1980), .B(n1979), .Z(n1951) );
  NAND U2068 ( .A(n1941), .B(n1940), .Z(n1945) );
  NAND U2069 ( .A(n1943), .B(n1942), .Z(n1944) );
  NAND U2070 ( .A(n1945), .B(n1944), .Z(n1952) );
  XNOR U2071 ( .A(n1951), .B(n1952), .Z(n1953) );
  XNOR U2072 ( .A(n1954), .B(n1953), .Z(n1983) );
  XNOR U2073 ( .A(n1983), .B(sreg[105]), .Z(n1985) );
  NAND U2074 ( .A(n1946), .B(sreg[104]), .Z(n1950) );
  OR U2075 ( .A(n1948), .B(n1947), .Z(n1949) );
  AND U2076 ( .A(n1950), .B(n1949), .Z(n1984) );
  XOR U2077 ( .A(n1985), .B(n1984), .Z(c[105]) );
  NANDN U2078 ( .A(n1960), .B(n1959), .Z(n1964) );
  NAND U2079 ( .A(n1962), .B(n1961), .Z(n1963) );
  NAND U2080 ( .A(n1964), .B(n1963), .Z(n2015) );
  NAND U2081 ( .A(n1965), .B(n2666), .Z(n1967) );
  XNOR U2082 ( .A(n2695), .B(a[44]), .Z(n2002) );
  NAND U2083 ( .A(n2002), .B(n2665), .Z(n1966) );
  NAND U2084 ( .A(n1967), .B(n1966), .Z(n1992) );
  XNOR U2085 ( .A(b[3]), .B(a[48]), .Z(n2005) );
  NANDN U2086 ( .A(n2005), .B(n2561), .Z(n1970) );
  NANDN U2087 ( .A(n1968), .B(n2563), .Z(n1969) );
  AND U2088 ( .A(n1970), .B(n1969), .Z(n1993) );
  XNOR U2089 ( .A(n1992), .B(n1993), .Z(n1994) );
  NANDN U2090 ( .A(n246), .B(a[50]), .Z(n1971) );
  XOR U2091 ( .A(n2537), .B(n1971), .Z(n1973) );
  NANDN U2092 ( .A(b[0]), .B(a[49]), .Z(n1972) );
  AND U2093 ( .A(n1973), .B(n1972), .Z(n1998) );
  NANDN U2094 ( .A(n1974), .B(n2625), .Z(n1976) );
  XNOR U2095 ( .A(b[5]), .B(a[46]), .Z(n2011) );
  OR U2096 ( .A(n2011), .B(n2608), .Z(n1975) );
  NAND U2097 ( .A(n1976), .B(n1975), .Z(n1996) );
  NANDN U2098 ( .A(n2695), .B(a[42]), .Z(n1997) );
  XNOR U2099 ( .A(n1996), .B(n1997), .Z(n1999) );
  XOR U2100 ( .A(n1998), .B(n1999), .Z(n1995) );
  XOR U2101 ( .A(n1994), .B(n1995), .Z(n2014) );
  XOR U2102 ( .A(n2015), .B(n2014), .Z(n2016) );
  XNOR U2103 ( .A(n2017), .B(n2016), .Z(n1988) );
  NAND U2104 ( .A(n1978), .B(n1977), .Z(n1982) );
  NAND U2105 ( .A(n1980), .B(n1979), .Z(n1981) );
  NAND U2106 ( .A(n1982), .B(n1981), .Z(n1989) );
  XNOR U2107 ( .A(n1988), .B(n1989), .Z(n1990) );
  XNOR U2108 ( .A(n1991), .B(n1990), .Z(n2020) );
  XNOR U2109 ( .A(n2020), .B(sreg[106]), .Z(n2022) );
  NAND U2110 ( .A(n1983), .B(sreg[105]), .Z(n1987) );
  OR U2111 ( .A(n1985), .B(n1984), .Z(n1986) );
  AND U2112 ( .A(n1987), .B(n1986), .Z(n2021) );
  XOR U2113 ( .A(n2022), .B(n2021), .Z(c[106]) );
  NANDN U2114 ( .A(n1997), .B(n1996), .Z(n2001) );
  NAND U2115 ( .A(n1999), .B(n1998), .Z(n2000) );
  NAND U2116 ( .A(n2001), .B(n2000), .Z(n2052) );
  NAND U2117 ( .A(n2002), .B(n2666), .Z(n2004) );
  XNOR U2118 ( .A(n2695), .B(a[45]), .Z(n2039) );
  NAND U2119 ( .A(n2039), .B(n2665), .Z(n2003) );
  NAND U2120 ( .A(n2004), .B(n2003), .Z(n2029) );
  XNOR U2121 ( .A(b[3]), .B(a[49]), .Z(n2042) );
  NANDN U2122 ( .A(n2042), .B(n2561), .Z(n2007) );
  NANDN U2123 ( .A(n2005), .B(n2563), .Z(n2006) );
  AND U2124 ( .A(n2007), .B(n2006), .Z(n2030) );
  XNOR U2125 ( .A(n2029), .B(n2030), .Z(n2031) );
  NANDN U2126 ( .A(n246), .B(a[51]), .Z(n2008) );
  XOR U2127 ( .A(n2537), .B(n2008), .Z(n2010) );
  NANDN U2128 ( .A(b[0]), .B(a[50]), .Z(n2009) );
  AND U2129 ( .A(n2010), .B(n2009), .Z(n2035) );
  NANDN U2130 ( .A(n2011), .B(n2625), .Z(n2013) );
  XNOR U2131 ( .A(b[5]), .B(a[47]), .Z(n2048) );
  OR U2132 ( .A(n2048), .B(n2608), .Z(n2012) );
  NAND U2133 ( .A(n2013), .B(n2012), .Z(n2033) );
  NANDN U2134 ( .A(n2695), .B(a[43]), .Z(n2034) );
  XNOR U2135 ( .A(n2033), .B(n2034), .Z(n2036) );
  XOR U2136 ( .A(n2035), .B(n2036), .Z(n2032) );
  XOR U2137 ( .A(n2031), .B(n2032), .Z(n2051) );
  XOR U2138 ( .A(n2052), .B(n2051), .Z(n2053) );
  XNOR U2139 ( .A(n2054), .B(n2053), .Z(n2025) );
  NAND U2140 ( .A(n2015), .B(n2014), .Z(n2019) );
  NAND U2141 ( .A(n2017), .B(n2016), .Z(n2018) );
  NAND U2142 ( .A(n2019), .B(n2018), .Z(n2026) );
  XNOR U2143 ( .A(n2025), .B(n2026), .Z(n2027) );
  XNOR U2144 ( .A(n2028), .B(n2027), .Z(n2057) );
  XNOR U2145 ( .A(n2057), .B(sreg[107]), .Z(n2059) );
  NAND U2146 ( .A(n2020), .B(sreg[106]), .Z(n2024) );
  OR U2147 ( .A(n2022), .B(n2021), .Z(n2023) );
  AND U2148 ( .A(n2024), .B(n2023), .Z(n2058) );
  XOR U2149 ( .A(n2059), .B(n2058), .Z(c[107]) );
  NANDN U2150 ( .A(n2034), .B(n2033), .Z(n2038) );
  NAND U2151 ( .A(n2036), .B(n2035), .Z(n2037) );
  NAND U2152 ( .A(n2038), .B(n2037), .Z(n2089) );
  NAND U2153 ( .A(n2039), .B(n2666), .Z(n2041) );
  XNOR U2154 ( .A(n2695), .B(a[46]), .Z(n2076) );
  NAND U2155 ( .A(n2076), .B(n2665), .Z(n2040) );
  NAND U2156 ( .A(n2041), .B(n2040), .Z(n2066) );
  XNOR U2157 ( .A(b[3]), .B(a[50]), .Z(n2079) );
  NANDN U2158 ( .A(n2079), .B(n2561), .Z(n2044) );
  NANDN U2159 ( .A(n2042), .B(n2563), .Z(n2043) );
  AND U2160 ( .A(n2044), .B(n2043), .Z(n2067) );
  XNOR U2161 ( .A(n2066), .B(n2067), .Z(n2068) );
  NANDN U2162 ( .A(n246), .B(a[52]), .Z(n2045) );
  XOR U2163 ( .A(n2537), .B(n2045), .Z(n2047) );
  NANDN U2164 ( .A(b[0]), .B(a[51]), .Z(n2046) );
  AND U2165 ( .A(n2047), .B(n2046), .Z(n2072) );
  NANDN U2166 ( .A(n2048), .B(n2625), .Z(n2050) );
  XNOR U2167 ( .A(b[5]), .B(a[48]), .Z(n2085) );
  OR U2168 ( .A(n2085), .B(n2608), .Z(n2049) );
  NAND U2169 ( .A(n2050), .B(n2049), .Z(n2070) );
  NANDN U2170 ( .A(n2695), .B(a[44]), .Z(n2071) );
  XNOR U2171 ( .A(n2070), .B(n2071), .Z(n2073) );
  XOR U2172 ( .A(n2072), .B(n2073), .Z(n2069) );
  XOR U2173 ( .A(n2068), .B(n2069), .Z(n2088) );
  XOR U2174 ( .A(n2089), .B(n2088), .Z(n2090) );
  XNOR U2175 ( .A(n2091), .B(n2090), .Z(n2062) );
  NAND U2176 ( .A(n2052), .B(n2051), .Z(n2056) );
  NAND U2177 ( .A(n2054), .B(n2053), .Z(n2055) );
  NAND U2178 ( .A(n2056), .B(n2055), .Z(n2063) );
  XNOR U2179 ( .A(n2062), .B(n2063), .Z(n2064) );
  XNOR U2180 ( .A(n2065), .B(n2064), .Z(n2094) );
  XNOR U2181 ( .A(n2094), .B(sreg[108]), .Z(n2096) );
  NAND U2182 ( .A(n2057), .B(sreg[107]), .Z(n2061) );
  OR U2183 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U2184 ( .A(n2061), .B(n2060), .Z(n2095) );
  XOR U2185 ( .A(n2096), .B(n2095), .Z(c[108]) );
  NANDN U2186 ( .A(n2071), .B(n2070), .Z(n2075) );
  NAND U2187 ( .A(n2073), .B(n2072), .Z(n2074) );
  NAND U2188 ( .A(n2075), .B(n2074), .Z(n2126) );
  NAND U2189 ( .A(n2076), .B(n2666), .Z(n2078) );
  XNOR U2190 ( .A(n2695), .B(a[47]), .Z(n2113) );
  NAND U2191 ( .A(n2113), .B(n2665), .Z(n2077) );
  NAND U2192 ( .A(n2078), .B(n2077), .Z(n2103) );
  XNOR U2193 ( .A(b[3]), .B(a[51]), .Z(n2116) );
  NANDN U2194 ( .A(n2116), .B(n2561), .Z(n2081) );
  NANDN U2195 ( .A(n2079), .B(n2563), .Z(n2080) );
  AND U2196 ( .A(n2081), .B(n2080), .Z(n2104) );
  XNOR U2197 ( .A(n2103), .B(n2104), .Z(n2105) );
  NANDN U2198 ( .A(n246), .B(a[53]), .Z(n2082) );
  XOR U2199 ( .A(n2537), .B(n2082), .Z(n2084) );
  NANDN U2200 ( .A(b[0]), .B(a[52]), .Z(n2083) );
  AND U2201 ( .A(n2084), .B(n2083), .Z(n2109) );
  NANDN U2202 ( .A(n2085), .B(n2625), .Z(n2087) );
  XNOR U2203 ( .A(b[5]), .B(a[49]), .Z(n2122) );
  OR U2204 ( .A(n2122), .B(n2608), .Z(n2086) );
  NAND U2205 ( .A(n2087), .B(n2086), .Z(n2107) );
  NANDN U2206 ( .A(n2695), .B(a[45]), .Z(n2108) );
  XNOR U2207 ( .A(n2107), .B(n2108), .Z(n2110) );
  XOR U2208 ( .A(n2109), .B(n2110), .Z(n2106) );
  XOR U2209 ( .A(n2105), .B(n2106), .Z(n2125) );
  XOR U2210 ( .A(n2126), .B(n2125), .Z(n2127) );
  XNOR U2211 ( .A(n2128), .B(n2127), .Z(n2099) );
  NAND U2212 ( .A(n2089), .B(n2088), .Z(n2093) );
  NAND U2213 ( .A(n2091), .B(n2090), .Z(n2092) );
  NAND U2214 ( .A(n2093), .B(n2092), .Z(n2100) );
  XNOR U2215 ( .A(n2099), .B(n2100), .Z(n2101) );
  XNOR U2216 ( .A(n2102), .B(n2101), .Z(n2131) );
  XNOR U2217 ( .A(n2131), .B(sreg[109]), .Z(n2133) );
  NAND U2218 ( .A(n2094), .B(sreg[108]), .Z(n2098) );
  OR U2219 ( .A(n2096), .B(n2095), .Z(n2097) );
  AND U2220 ( .A(n2098), .B(n2097), .Z(n2132) );
  XOR U2221 ( .A(n2133), .B(n2132), .Z(c[109]) );
  NANDN U2222 ( .A(n2108), .B(n2107), .Z(n2112) );
  NAND U2223 ( .A(n2110), .B(n2109), .Z(n2111) );
  NAND U2224 ( .A(n2112), .B(n2111), .Z(n2163) );
  NAND U2225 ( .A(n2113), .B(n2666), .Z(n2115) );
  XNOR U2226 ( .A(n2695), .B(a[48]), .Z(n2150) );
  NAND U2227 ( .A(n2150), .B(n2665), .Z(n2114) );
  NAND U2228 ( .A(n2115), .B(n2114), .Z(n2140) );
  XNOR U2229 ( .A(b[3]), .B(a[52]), .Z(n2153) );
  NANDN U2230 ( .A(n2153), .B(n2561), .Z(n2118) );
  NANDN U2231 ( .A(n2116), .B(n2563), .Z(n2117) );
  AND U2232 ( .A(n2118), .B(n2117), .Z(n2141) );
  XNOR U2233 ( .A(n2140), .B(n2141), .Z(n2142) );
  NANDN U2234 ( .A(n246), .B(a[54]), .Z(n2119) );
  XOR U2235 ( .A(n2537), .B(n2119), .Z(n2121) );
  NANDN U2236 ( .A(b[0]), .B(a[53]), .Z(n2120) );
  AND U2237 ( .A(n2121), .B(n2120), .Z(n2146) );
  NANDN U2238 ( .A(n2122), .B(n2625), .Z(n2124) );
  XNOR U2239 ( .A(b[5]), .B(a[50]), .Z(n2159) );
  OR U2240 ( .A(n2159), .B(n2608), .Z(n2123) );
  NAND U2241 ( .A(n2124), .B(n2123), .Z(n2144) );
  NANDN U2242 ( .A(n2695), .B(a[46]), .Z(n2145) );
  XNOR U2243 ( .A(n2144), .B(n2145), .Z(n2147) );
  XOR U2244 ( .A(n2146), .B(n2147), .Z(n2143) );
  XOR U2245 ( .A(n2142), .B(n2143), .Z(n2162) );
  XOR U2246 ( .A(n2163), .B(n2162), .Z(n2164) );
  XNOR U2247 ( .A(n2165), .B(n2164), .Z(n2136) );
  NAND U2248 ( .A(n2126), .B(n2125), .Z(n2130) );
  NAND U2249 ( .A(n2128), .B(n2127), .Z(n2129) );
  NAND U2250 ( .A(n2130), .B(n2129), .Z(n2137) );
  XNOR U2251 ( .A(n2136), .B(n2137), .Z(n2138) );
  XNOR U2252 ( .A(n2139), .B(n2138), .Z(n2168) );
  XNOR U2253 ( .A(n2168), .B(sreg[110]), .Z(n2170) );
  NAND U2254 ( .A(n2131), .B(sreg[109]), .Z(n2135) );
  OR U2255 ( .A(n2133), .B(n2132), .Z(n2134) );
  AND U2256 ( .A(n2135), .B(n2134), .Z(n2169) );
  XOR U2257 ( .A(n2170), .B(n2169), .Z(c[110]) );
  NANDN U2258 ( .A(n2145), .B(n2144), .Z(n2149) );
  NAND U2259 ( .A(n2147), .B(n2146), .Z(n2148) );
  NAND U2260 ( .A(n2149), .B(n2148), .Z(n2200) );
  NAND U2261 ( .A(n2150), .B(n2666), .Z(n2152) );
  XNOR U2262 ( .A(n2695), .B(a[49]), .Z(n2187) );
  NAND U2263 ( .A(n2187), .B(n2665), .Z(n2151) );
  NAND U2264 ( .A(n2152), .B(n2151), .Z(n2177) );
  XNOR U2265 ( .A(b[3]), .B(a[53]), .Z(n2190) );
  NANDN U2266 ( .A(n2190), .B(n2561), .Z(n2155) );
  NANDN U2267 ( .A(n2153), .B(n2563), .Z(n2154) );
  AND U2268 ( .A(n2155), .B(n2154), .Z(n2178) );
  XNOR U2269 ( .A(n2177), .B(n2178), .Z(n2179) );
  NANDN U2270 ( .A(n246), .B(a[55]), .Z(n2156) );
  XOR U2271 ( .A(n2537), .B(n2156), .Z(n2158) );
  NANDN U2272 ( .A(b[0]), .B(a[54]), .Z(n2157) );
  AND U2273 ( .A(n2158), .B(n2157), .Z(n2183) );
  NANDN U2274 ( .A(n2159), .B(n2625), .Z(n2161) );
  XNOR U2275 ( .A(b[5]), .B(a[51]), .Z(n2196) );
  OR U2276 ( .A(n2196), .B(n2608), .Z(n2160) );
  NAND U2277 ( .A(n2161), .B(n2160), .Z(n2181) );
  NANDN U2278 ( .A(n2695), .B(a[47]), .Z(n2182) );
  XNOR U2279 ( .A(n2181), .B(n2182), .Z(n2184) );
  XOR U2280 ( .A(n2183), .B(n2184), .Z(n2180) );
  XOR U2281 ( .A(n2179), .B(n2180), .Z(n2199) );
  XOR U2282 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U2283 ( .A(n2202), .B(n2201), .Z(n2173) );
  NAND U2284 ( .A(n2163), .B(n2162), .Z(n2167) );
  NAND U2285 ( .A(n2165), .B(n2164), .Z(n2166) );
  NAND U2286 ( .A(n2167), .B(n2166), .Z(n2174) );
  XNOR U2287 ( .A(n2173), .B(n2174), .Z(n2175) );
  XNOR U2288 ( .A(n2176), .B(n2175), .Z(n2205) );
  XNOR U2289 ( .A(n2205), .B(sreg[111]), .Z(n2207) );
  NAND U2290 ( .A(n2168), .B(sreg[110]), .Z(n2172) );
  OR U2291 ( .A(n2170), .B(n2169), .Z(n2171) );
  AND U2292 ( .A(n2172), .B(n2171), .Z(n2206) );
  XOR U2293 ( .A(n2207), .B(n2206), .Z(c[111]) );
  NANDN U2294 ( .A(n2182), .B(n2181), .Z(n2186) );
  NAND U2295 ( .A(n2184), .B(n2183), .Z(n2185) );
  NAND U2296 ( .A(n2186), .B(n2185), .Z(n2237) );
  NAND U2297 ( .A(n2187), .B(n2666), .Z(n2189) );
  XNOR U2298 ( .A(n2695), .B(a[50]), .Z(n2224) );
  NAND U2299 ( .A(n2224), .B(n2665), .Z(n2188) );
  NAND U2300 ( .A(n2189), .B(n2188), .Z(n2214) );
  XNOR U2301 ( .A(b[3]), .B(a[54]), .Z(n2227) );
  NANDN U2302 ( .A(n2227), .B(n2561), .Z(n2192) );
  NANDN U2303 ( .A(n2190), .B(n2563), .Z(n2191) );
  AND U2304 ( .A(n2192), .B(n2191), .Z(n2215) );
  XNOR U2305 ( .A(n2214), .B(n2215), .Z(n2216) );
  NANDN U2306 ( .A(n246), .B(a[56]), .Z(n2193) );
  XOR U2307 ( .A(n2537), .B(n2193), .Z(n2195) );
  IV U2308 ( .A(a[55]), .Z(n2448) );
  NANDN U2309 ( .A(n2448), .B(n246), .Z(n2194) );
  AND U2310 ( .A(n2195), .B(n2194), .Z(n2220) );
  NANDN U2311 ( .A(n2196), .B(n2625), .Z(n2198) );
  XNOR U2312 ( .A(b[5]), .B(a[52]), .Z(n2233) );
  OR U2313 ( .A(n2233), .B(n2608), .Z(n2197) );
  NAND U2314 ( .A(n2198), .B(n2197), .Z(n2218) );
  NANDN U2315 ( .A(n2695), .B(a[48]), .Z(n2219) );
  XNOR U2316 ( .A(n2218), .B(n2219), .Z(n2221) );
  XOR U2317 ( .A(n2220), .B(n2221), .Z(n2217) );
  XOR U2318 ( .A(n2216), .B(n2217), .Z(n2236) );
  XOR U2319 ( .A(n2237), .B(n2236), .Z(n2238) );
  XNOR U2320 ( .A(n2239), .B(n2238), .Z(n2210) );
  NAND U2321 ( .A(n2200), .B(n2199), .Z(n2204) );
  NAND U2322 ( .A(n2202), .B(n2201), .Z(n2203) );
  NAND U2323 ( .A(n2204), .B(n2203), .Z(n2211) );
  XNOR U2324 ( .A(n2210), .B(n2211), .Z(n2212) );
  XNOR U2325 ( .A(n2213), .B(n2212), .Z(n2242) );
  XNOR U2326 ( .A(n2242), .B(sreg[112]), .Z(n2244) );
  NAND U2327 ( .A(n2205), .B(sreg[111]), .Z(n2209) );
  OR U2328 ( .A(n2207), .B(n2206), .Z(n2208) );
  AND U2329 ( .A(n2209), .B(n2208), .Z(n2243) );
  XOR U2330 ( .A(n2244), .B(n2243), .Z(c[112]) );
  NANDN U2331 ( .A(n2219), .B(n2218), .Z(n2223) );
  NAND U2332 ( .A(n2221), .B(n2220), .Z(n2222) );
  NAND U2333 ( .A(n2223), .B(n2222), .Z(n2274) );
  NAND U2334 ( .A(n2224), .B(n2666), .Z(n2226) );
  XNOR U2335 ( .A(n2695), .B(a[51]), .Z(n2261) );
  NAND U2336 ( .A(n2261), .B(n2665), .Z(n2225) );
  NAND U2337 ( .A(n2226), .B(n2225), .Z(n2251) );
  XOR U2338 ( .A(b[3]), .B(n2448), .Z(n2264) );
  NANDN U2339 ( .A(n2264), .B(n2561), .Z(n2229) );
  NANDN U2340 ( .A(n2227), .B(n2563), .Z(n2228) );
  AND U2341 ( .A(n2229), .B(n2228), .Z(n2252) );
  XNOR U2342 ( .A(n2251), .B(n2252), .Z(n2253) );
  NANDN U2343 ( .A(n246), .B(a[57]), .Z(n2230) );
  XOR U2344 ( .A(n2537), .B(n2230), .Z(n2232) );
  NANDN U2345 ( .A(b[0]), .B(a[56]), .Z(n2231) );
  AND U2346 ( .A(n2232), .B(n2231), .Z(n2257) );
  NANDN U2347 ( .A(n2233), .B(n2625), .Z(n2235) );
  XNOR U2348 ( .A(b[5]), .B(a[53]), .Z(n2270) );
  OR U2349 ( .A(n2270), .B(n2608), .Z(n2234) );
  NAND U2350 ( .A(n2235), .B(n2234), .Z(n2255) );
  NANDN U2351 ( .A(n2695), .B(a[49]), .Z(n2256) );
  XNOR U2352 ( .A(n2255), .B(n2256), .Z(n2258) );
  XOR U2353 ( .A(n2257), .B(n2258), .Z(n2254) );
  XOR U2354 ( .A(n2253), .B(n2254), .Z(n2273) );
  XOR U2355 ( .A(n2274), .B(n2273), .Z(n2275) );
  XNOR U2356 ( .A(n2276), .B(n2275), .Z(n2247) );
  NAND U2357 ( .A(n2237), .B(n2236), .Z(n2241) );
  NAND U2358 ( .A(n2239), .B(n2238), .Z(n2240) );
  NAND U2359 ( .A(n2241), .B(n2240), .Z(n2248) );
  XNOR U2360 ( .A(n2247), .B(n2248), .Z(n2249) );
  XNOR U2361 ( .A(n2250), .B(n2249), .Z(n2279) );
  XNOR U2362 ( .A(n2279), .B(sreg[113]), .Z(n2281) );
  NAND U2363 ( .A(n2242), .B(sreg[112]), .Z(n2246) );
  OR U2364 ( .A(n2244), .B(n2243), .Z(n2245) );
  AND U2365 ( .A(n2246), .B(n2245), .Z(n2280) );
  XOR U2366 ( .A(n2281), .B(n2280), .Z(c[113]) );
  NANDN U2367 ( .A(n2256), .B(n2255), .Z(n2260) );
  NAND U2368 ( .A(n2258), .B(n2257), .Z(n2259) );
  NAND U2369 ( .A(n2260), .B(n2259), .Z(n2311) );
  NAND U2370 ( .A(n2261), .B(n2666), .Z(n2263) );
  XNOR U2371 ( .A(n2695), .B(a[52]), .Z(n2298) );
  NAND U2372 ( .A(n2298), .B(n2665), .Z(n2262) );
  NAND U2373 ( .A(n2263), .B(n2262), .Z(n2288) );
  XNOR U2374 ( .A(b[3]), .B(a[56]), .Z(n2301) );
  NANDN U2375 ( .A(n2301), .B(n2561), .Z(n2266) );
  NANDN U2376 ( .A(n2264), .B(n2563), .Z(n2265) );
  AND U2377 ( .A(n2266), .B(n2265), .Z(n2289) );
  XNOR U2378 ( .A(n2288), .B(n2289), .Z(n2290) );
  NANDN U2379 ( .A(n246), .B(a[58]), .Z(n2267) );
  XOR U2380 ( .A(n2537), .B(n2267), .Z(n2269) );
  IV U2381 ( .A(a[57]), .Z(n2382) );
  NANDN U2382 ( .A(n2382), .B(n246), .Z(n2268) );
  AND U2383 ( .A(n2269), .B(n2268), .Z(n2294) );
  NANDN U2384 ( .A(n2270), .B(n2625), .Z(n2272) );
  XNOR U2385 ( .A(b[5]), .B(a[54]), .Z(n2307) );
  OR U2386 ( .A(n2307), .B(n2608), .Z(n2271) );
  NAND U2387 ( .A(n2272), .B(n2271), .Z(n2292) );
  NANDN U2388 ( .A(n2695), .B(a[50]), .Z(n2293) );
  XNOR U2389 ( .A(n2292), .B(n2293), .Z(n2295) );
  XOR U2390 ( .A(n2294), .B(n2295), .Z(n2291) );
  XOR U2391 ( .A(n2290), .B(n2291), .Z(n2310) );
  XOR U2392 ( .A(n2311), .B(n2310), .Z(n2312) );
  XNOR U2393 ( .A(n2313), .B(n2312), .Z(n2284) );
  NAND U2394 ( .A(n2274), .B(n2273), .Z(n2278) );
  NAND U2395 ( .A(n2276), .B(n2275), .Z(n2277) );
  NAND U2396 ( .A(n2278), .B(n2277), .Z(n2285) );
  XNOR U2397 ( .A(n2284), .B(n2285), .Z(n2286) );
  XNOR U2398 ( .A(n2287), .B(n2286), .Z(n2316) );
  XNOR U2399 ( .A(n2316), .B(sreg[114]), .Z(n2318) );
  NAND U2400 ( .A(n2279), .B(sreg[113]), .Z(n2283) );
  OR U2401 ( .A(n2281), .B(n2280), .Z(n2282) );
  AND U2402 ( .A(n2283), .B(n2282), .Z(n2317) );
  XOR U2403 ( .A(n2318), .B(n2317), .Z(c[114]) );
  NANDN U2404 ( .A(n2293), .B(n2292), .Z(n2297) );
  NAND U2405 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2406 ( .A(n2297), .B(n2296), .Z(n2348) );
  NAND U2407 ( .A(n2298), .B(n2666), .Z(n2300) );
  XNOR U2408 ( .A(n2695), .B(a[53]), .Z(n2335) );
  NAND U2409 ( .A(n2335), .B(n2665), .Z(n2299) );
  NAND U2410 ( .A(n2300), .B(n2299), .Z(n2325) );
  XOR U2411 ( .A(b[3]), .B(n2382), .Z(n2338) );
  NANDN U2412 ( .A(n2338), .B(n2561), .Z(n2303) );
  NANDN U2413 ( .A(n2301), .B(n2563), .Z(n2302) );
  AND U2414 ( .A(n2303), .B(n2302), .Z(n2326) );
  XNOR U2415 ( .A(n2325), .B(n2326), .Z(n2327) );
  NANDN U2416 ( .A(n246), .B(a[59]), .Z(n2304) );
  XOR U2417 ( .A(n2537), .B(n2304), .Z(n2306) );
  IV U2418 ( .A(a[58]), .Z(n2420) );
  NANDN U2419 ( .A(n2420), .B(n246), .Z(n2305) );
  AND U2420 ( .A(n2306), .B(n2305), .Z(n2331) );
  NANDN U2421 ( .A(n2307), .B(n2625), .Z(n2309) );
  XOR U2422 ( .A(b[5]), .B(n2448), .Z(n2344) );
  OR U2423 ( .A(n2344), .B(n2608), .Z(n2308) );
  NAND U2424 ( .A(n2309), .B(n2308), .Z(n2329) );
  NANDN U2425 ( .A(n2695), .B(a[51]), .Z(n2330) );
  XNOR U2426 ( .A(n2329), .B(n2330), .Z(n2332) );
  XOR U2427 ( .A(n2331), .B(n2332), .Z(n2328) );
  XOR U2428 ( .A(n2327), .B(n2328), .Z(n2347) );
  XOR U2429 ( .A(n2348), .B(n2347), .Z(n2349) );
  XNOR U2430 ( .A(n2350), .B(n2349), .Z(n2321) );
  NAND U2431 ( .A(n2311), .B(n2310), .Z(n2315) );
  NAND U2432 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U2433 ( .A(n2315), .B(n2314), .Z(n2322) );
  XNOR U2434 ( .A(n2321), .B(n2322), .Z(n2323) );
  XNOR U2435 ( .A(n2324), .B(n2323), .Z(n2353) );
  XNOR U2436 ( .A(n2353), .B(sreg[115]), .Z(n2355) );
  NAND U2437 ( .A(n2316), .B(sreg[114]), .Z(n2320) );
  OR U2438 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U2439 ( .A(n2320), .B(n2319), .Z(n2354) );
  XOR U2440 ( .A(n2355), .B(n2354), .Z(c[115]) );
  NANDN U2441 ( .A(n2330), .B(n2329), .Z(n2334) );
  NAND U2442 ( .A(n2332), .B(n2331), .Z(n2333) );
  NAND U2443 ( .A(n2334), .B(n2333), .Z(n2386) );
  NAND U2444 ( .A(n2335), .B(n2666), .Z(n2337) );
  XNOR U2445 ( .A(n2695), .B(a[54]), .Z(n2372) );
  NAND U2446 ( .A(n2372), .B(n2665), .Z(n2336) );
  NAND U2447 ( .A(n2337), .B(n2336), .Z(n2362) );
  XOR U2448 ( .A(b[3]), .B(n2420), .Z(n2375) );
  NANDN U2449 ( .A(n2375), .B(n2561), .Z(n2340) );
  NANDN U2450 ( .A(n2338), .B(n2563), .Z(n2339) );
  AND U2451 ( .A(n2340), .B(n2339), .Z(n2363) );
  XNOR U2452 ( .A(n2362), .B(n2363), .Z(n2364) );
  NANDN U2453 ( .A(n246), .B(a[60]), .Z(n2341) );
  XOR U2454 ( .A(n2537), .B(n2341), .Z(n2343) );
  NANDN U2455 ( .A(b[0]), .B(a[59]), .Z(n2342) );
  AND U2456 ( .A(n2343), .B(n2342), .Z(n2368) );
  NANDN U2457 ( .A(n2344), .B(n2625), .Z(n2346) );
  XNOR U2458 ( .A(b[5]), .B(a[56]), .Z(n2381) );
  OR U2459 ( .A(n2381), .B(n2608), .Z(n2345) );
  NAND U2460 ( .A(n2346), .B(n2345), .Z(n2366) );
  NANDN U2461 ( .A(n2695), .B(a[52]), .Z(n2367) );
  XNOR U2462 ( .A(n2366), .B(n2367), .Z(n2369) );
  XOR U2463 ( .A(n2368), .B(n2369), .Z(n2365) );
  XOR U2464 ( .A(n2364), .B(n2365), .Z(n2385) );
  XOR U2465 ( .A(n2386), .B(n2385), .Z(n2387) );
  XNOR U2466 ( .A(n2388), .B(n2387), .Z(n2358) );
  NAND U2467 ( .A(n2348), .B(n2347), .Z(n2352) );
  NAND U2468 ( .A(n2350), .B(n2349), .Z(n2351) );
  NAND U2469 ( .A(n2352), .B(n2351), .Z(n2359) );
  XNOR U2470 ( .A(n2358), .B(n2359), .Z(n2360) );
  XNOR U2471 ( .A(n2361), .B(n2360), .Z(n2391) );
  XNOR U2472 ( .A(n2391), .B(sreg[116]), .Z(n2393) );
  NAND U2473 ( .A(n2353), .B(sreg[115]), .Z(n2357) );
  OR U2474 ( .A(n2355), .B(n2354), .Z(n2356) );
  AND U2475 ( .A(n2357), .B(n2356), .Z(n2392) );
  XOR U2476 ( .A(n2393), .B(n2392), .Z(c[116]) );
  NANDN U2477 ( .A(n2367), .B(n2366), .Z(n2371) );
  NAND U2478 ( .A(n2369), .B(n2368), .Z(n2370) );
  NAND U2479 ( .A(n2371), .B(n2370), .Z(n2424) );
  NAND U2480 ( .A(n2372), .B(n2666), .Z(n2374) );
  XNOR U2481 ( .A(n2695), .B(a[55]), .Z(n2410) );
  NAND U2482 ( .A(n2410), .B(n2665), .Z(n2373) );
  NAND U2483 ( .A(n2374), .B(n2373), .Z(n2400) );
  XNOR U2484 ( .A(b[3]), .B(a[59]), .Z(n2413) );
  NANDN U2485 ( .A(n2413), .B(n2561), .Z(n2377) );
  NANDN U2486 ( .A(n2375), .B(n2563), .Z(n2376) );
  AND U2487 ( .A(n2377), .B(n2376), .Z(n2401) );
  XNOR U2488 ( .A(n2400), .B(n2401), .Z(n2402) );
  NANDN U2489 ( .A(n246), .B(a[61]), .Z(n2378) );
  XOR U2490 ( .A(n2537), .B(n2378), .Z(n2380) );
  IV U2491 ( .A(a[60]), .Z(n2629) );
  NANDN U2492 ( .A(n2629), .B(n246), .Z(n2379) );
  AND U2493 ( .A(n2380), .B(n2379), .Z(n2406) );
  NANDN U2494 ( .A(n2381), .B(n2625), .Z(n2384) );
  XOR U2495 ( .A(b[5]), .B(n2382), .Z(n2419) );
  OR U2496 ( .A(n2419), .B(n2608), .Z(n2383) );
  NAND U2497 ( .A(n2384), .B(n2383), .Z(n2404) );
  NANDN U2498 ( .A(n2695), .B(a[53]), .Z(n2405) );
  XNOR U2499 ( .A(n2404), .B(n2405), .Z(n2407) );
  XOR U2500 ( .A(n2406), .B(n2407), .Z(n2403) );
  XOR U2501 ( .A(n2402), .B(n2403), .Z(n2423) );
  XOR U2502 ( .A(n2424), .B(n2423), .Z(n2425) );
  XNOR U2503 ( .A(n2426), .B(n2425), .Z(n2396) );
  NAND U2504 ( .A(n2386), .B(n2385), .Z(n2390) );
  NAND U2505 ( .A(n2388), .B(n2387), .Z(n2389) );
  NAND U2506 ( .A(n2390), .B(n2389), .Z(n2397) );
  XNOR U2507 ( .A(n2396), .B(n2397), .Z(n2398) );
  XNOR U2508 ( .A(n2399), .B(n2398), .Z(n2429) );
  XNOR U2509 ( .A(n2429), .B(sreg[117]), .Z(n2431) );
  NAND U2510 ( .A(n2391), .B(sreg[116]), .Z(n2395) );
  OR U2511 ( .A(n2393), .B(n2392), .Z(n2394) );
  AND U2512 ( .A(n2395), .B(n2394), .Z(n2430) );
  XOR U2513 ( .A(n2431), .B(n2430), .Z(c[117]) );
  NANDN U2514 ( .A(n2405), .B(n2404), .Z(n2409) );
  NAND U2515 ( .A(n2407), .B(n2406), .Z(n2408) );
  NAND U2516 ( .A(n2409), .B(n2408), .Z(n2462) );
  NAND U2517 ( .A(n2410), .B(n2666), .Z(n2412) );
  XNOR U2518 ( .A(n2695), .B(a[56]), .Z(n2455) );
  NAND U2519 ( .A(n2455), .B(n2665), .Z(n2411) );
  NAND U2520 ( .A(n2412), .B(n2411), .Z(n2438) );
  XOR U2521 ( .A(b[3]), .B(n2629), .Z(n2458) );
  NANDN U2522 ( .A(n2458), .B(n2561), .Z(n2415) );
  NANDN U2523 ( .A(n2413), .B(n2563), .Z(n2414) );
  AND U2524 ( .A(n2415), .B(n2414), .Z(n2439) );
  XNOR U2525 ( .A(n2438), .B(n2439), .Z(n2440) );
  IV U2526 ( .A(a[62]), .Z(n2631) );
  NANDN U2527 ( .A(n2631), .B(b[0]), .Z(n2416) );
  XOR U2528 ( .A(n2537), .B(n2416), .Z(n2418) );
  NANDN U2529 ( .A(b[0]), .B(a[61]), .Z(n2417) );
  AND U2530 ( .A(n2418), .B(n2417), .Z(n2444) );
  NANDN U2531 ( .A(n2419), .B(n2625), .Z(n2422) );
  XOR U2532 ( .A(n248), .B(n2420), .Z(n2452) );
  NANDN U2533 ( .A(n2608), .B(n2452), .Z(n2421) );
  NAND U2534 ( .A(n2422), .B(n2421), .Z(n2442) );
  NANDN U2535 ( .A(n2695), .B(a[54]), .Z(n2443) );
  XNOR U2536 ( .A(n2442), .B(n2443), .Z(n2445) );
  XOR U2537 ( .A(n2444), .B(n2445), .Z(n2441) );
  XOR U2538 ( .A(n2440), .B(n2441), .Z(n2461) );
  XOR U2539 ( .A(n2462), .B(n2461), .Z(n2463) );
  XNOR U2540 ( .A(n2464), .B(n2463), .Z(n2434) );
  NAND U2541 ( .A(n2424), .B(n2423), .Z(n2428) );
  NAND U2542 ( .A(n2426), .B(n2425), .Z(n2427) );
  NAND U2543 ( .A(n2428), .B(n2427), .Z(n2435) );
  XNOR U2544 ( .A(n2434), .B(n2435), .Z(n2436) );
  XNOR U2545 ( .A(n2437), .B(n2436), .Z(n2467) );
  XNOR U2546 ( .A(n2467), .B(sreg[118]), .Z(n2469) );
  NAND U2547 ( .A(n2429), .B(sreg[117]), .Z(n2433) );
  OR U2548 ( .A(n2431), .B(n2430), .Z(n2432) );
  AND U2549 ( .A(n2433), .B(n2432), .Z(n2468) );
  XOR U2550 ( .A(n2469), .B(n2468), .Z(c[118]) );
  NANDN U2551 ( .A(n2443), .B(n2442), .Z(n2447) );
  NAND U2552 ( .A(n2445), .B(n2444), .Z(n2446) );
  NAND U2553 ( .A(n2447), .B(n2446), .Z(n2477) );
  ANDN U2554 ( .B(b[7]), .A(n2448), .Z(n2489) );
  NANDN U2555 ( .A(n246), .B(a[63]), .Z(n2449) );
  XOR U2556 ( .A(n2537), .B(n2449), .Z(n2451) );
  NANDN U2557 ( .A(n2631), .B(n246), .Z(n2450) );
  AND U2558 ( .A(n2451), .B(n2450), .Z(n2487) );
  XOR U2559 ( .A(n248), .B(a[59]), .Z(n2500) );
  OR U2560 ( .A(n2500), .B(n2608), .Z(n2454) );
  NAND U2561 ( .A(n2625), .B(n2452), .Z(n2453) );
  AND U2562 ( .A(n2454), .B(n2453), .Z(n2486) );
  XNOR U2563 ( .A(n2487), .B(n2486), .Z(n2488) );
  XOR U2564 ( .A(n2489), .B(n2488), .Z(n2485) );
  NAND U2565 ( .A(n2455), .B(n2666), .Z(n2457) );
  XNOR U2566 ( .A(n2695), .B(a[57]), .Z(n2492) );
  NAND U2567 ( .A(n2492), .B(n2665), .Z(n2456) );
  NAND U2568 ( .A(n2457), .B(n2456), .Z(n2482) );
  XNOR U2569 ( .A(a[61]), .B(b[3]), .Z(n2495) );
  NANDN U2570 ( .A(n2495), .B(n2561), .Z(n2460) );
  NANDN U2571 ( .A(n2458), .B(n2563), .Z(n2459) );
  AND U2572 ( .A(n2460), .B(n2459), .Z(n2483) );
  XNOR U2573 ( .A(n2482), .B(n2483), .Z(n2484) );
  XOR U2574 ( .A(n2485), .B(n2484), .Z(n2476) );
  XOR U2575 ( .A(n2477), .B(n2476), .Z(n2478) );
  XNOR U2576 ( .A(n2479), .B(n2478), .Z(n2472) );
  NAND U2577 ( .A(n2462), .B(n2461), .Z(n2466) );
  NAND U2578 ( .A(n2464), .B(n2463), .Z(n2465) );
  NAND U2579 ( .A(n2466), .B(n2465), .Z(n2473) );
  XNOR U2580 ( .A(n2472), .B(n2473), .Z(n2474) );
  XNOR U2581 ( .A(n2475), .B(n2474), .Z(n2503) );
  XNOR U2582 ( .A(n2503), .B(sreg[119]), .Z(n2505) );
  NAND U2583 ( .A(n2467), .B(sreg[118]), .Z(n2471) );
  OR U2584 ( .A(n2469), .B(n2468), .Z(n2470) );
  AND U2585 ( .A(n2471), .B(n2470), .Z(n2504) );
  XOR U2586 ( .A(n2505), .B(n2504), .Z(c[119]) );
  NAND U2587 ( .A(n2477), .B(n2476), .Z(n2481) );
  NAND U2588 ( .A(n2479), .B(n2478), .Z(n2480) );
  NAND U2589 ( .A(n2481), .B(n2480), .Z(n2510) );
  NANDN U2590 ( .A(n2487), .B(n2486), .Z(n2491) );
  NANDN U2591 ( .A(n2489), .B(n2488), .Z(n2490) );
  NAND U2592 ( .A(n2491), .B(n2490), .Z(n2538) );
  NAND U2593 ( .A(n2492), .B(n2666), .Z(n2494) );
  XNOR U2594 ( .A(n2695), .B(a[58]), .Z(n2528) );
  NAND U2595 ( .A(n2528), .B(n2665), .Z(n2493) );
  NAND U2596 ( .A(n2494), .B(n2493), .Z(n2518) );
  XOR U2597 ( .A(a[62]), .B(n247), .Z(n2534) );
  NANDN U2598 ( .A(n2534), .B(n2561), .Z(n2497) );
  NANDN U2599 ( .A(n2495), .B(n2563), .Z(n2496) );
  NAND U2600 ( .A(n2497), .B(n2496), .Z(n2516) );
  IV U2601 ( .A(a[63]), .Z(n2696) );
  NANDN U2602 ( .A(n2537), .B(n2696), .Z(n2499) );
  NANDN U2603 ( .A(n246), .B(b[1]), .Z(n2498) );
  AND U2604 ( .A(n2499), .B(n2498), .Z(n2522) );
  NANDN U2605 ( .A(n2695), .B(a[56]), .Z(n2523) );
  XNOR U2606 ( .A(n2522), .B(n2523), .Z(n2524) );
  XOR U2607 ( .A(n248), .B(a[60]), .Z(n2531) );
  OR U2608 ( .A(n2531), .B(n2608), .Z(n2502) );
  NANDN U2609 ( .A(n2500), .B(n2625), .Z(n2501) );
  AND U2610 ( .A(n2502), .B(n2501), .Z(n2525) );
  XOR U2611 ( .A(n2516), .B(n2517), .Z(n2519) );
  XNOR U2612 ( .A(n2518), .B(n2519), .Z(n2539) );
  XNOR U2613 ( .A(n2538), .B(n2539), .Z(n2540) );
  XOR U2614 ( .A(n2541), .B(n2540), .Z(n2511) );
  XOR U2615 ( .A(n2510), .B(n2511), .Z(n2512) );
  XOR U2616 ( .A(n2513), .B(n2512), .Z(n2509) );
  NAND U2617 ( .A(n2503), .B(sreg[119]), .Z(n2507) );
  OR U2618 ( .A(n2505), .B(n2504), .Z(n2506) );
  AND U2619 ( .A(n2507), .B(n2506), .Z(n2508) );
  XOR U2620 ( .A(n2509), .B(n2508), .Z(c[120]) );
  OR U2621 ( .A(n2509), .B(n2508), .Z(n2579) );
  OR U2622 ( .A(n2511), .B(n2510), .Z(n2515) );
  NAND U2623 ( .A(n2513), .B(n2512), .Z(n2514) );
  NAND U2624 ( .A(n2515), .B(n2514), .Z(n2547) );
  NANDN U2625 ( .A(n2517), .B(n2516), .Z(n2521) );
  NANDN U2626 ( .A(n2519), .B(n2518), .Z(n2520) );
  NAND U2627 ( .A(n2521), .B(n2520), .Z(n2550) );
  OR U2628 ( .A(n2523), .B(n2522), .Z(n2527) );
  OR U2629 ( .A(n2525), .B(n2524), .Z(n2526) );
  AND U2630 ( .A(n2527), .B(n2526), .Z(n2551) );
  XNOR U2631 ( .A(n2550), .B(n2551), .Z(n2552) );
  NAND U2632 ( .A(n2528), .B(n2666), .Z(n2530) );
  XNOR U2633 ( .A(n2695), .B(a[59]), .Z(n2566) );
  NAND U2634 ( .A(n2566), .B(n2665), .Z(n2529) );
  NAND U2635 ( .A(n2530), .B(n2529), .Z(n2572) );
  AND U2636 ( .A(a[57]), .B(b[7]), .Z(n2636) );
  XOR U2637 ( .A(n2572), .B(n2636), .Z(n2574) );
  XOR U2638 ( .A(a[61]), .B(n248), .Z(n2569) );
  OR U2639 ( .A(n2569), .B(n2608), .Z(n2533) );
  NANDN U2640 ( .A(n2531), .B(n2625), .Z(n2532) );
  NAND U2641 ( .A(n2533), .B(n2532), .Z(n2573) );
  XNOR U2642 ( .A(n2574), .B(n2573), .Z(n2558) );
  XOR U2643 ( .A(n247), .B(n2696), .Z(n2562) );
  NAND U2644 ( .A(n2562), .B(n2561), .Z(n2536) );
  NANDN U2645 ( .A(n2534), .B(n2563), .Z(n2535) );
  AND U2646 ( .A(n2536), .B(n2535), .Z(n2556) );
  XNOR U2647 ( .A(n2537), .B(n2556), .Z(n2557) );
  XNOR U2648 ( .A(n2558), .B(n2557), .Z(n2553) );
  XOR U2649 ( .A(n2552), .B(n2553), .Z(n2544) );
  NANDN U2650 ( .A(n2539), .B(n2538), .Z(n2543) );
  NANDN U2651 ( .A(n2541), .B(n2540), .Z(n2542) );
  AND U2652 ( .A(n2543), .B(n2542), .Z(n2545) );
  XNOR U2653 ( .A(n2544), .B(n2545), .Z(n2546) );
  XOR U2654 ( .A(n2547), .B(n2546), .Z(n2578) );
  XOR U2655 ( .A(n2579), .B(n2578), .Z(c[121]) );
  NANDN U2656 ( .A(n2545), .B(n2544), .Z(n2549) );
  NAND U2657 ( .A(n2547), .B(n2546), .Z(n2548) );
  AND U2658 ( .A(n2549), .B(n2548), .Z(n2584) );
  NANDN U2659 ( .A(n2551), .B(n2550), .Z(n2555) );
  NANDN U2660 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND U2661 ( .A(n2555), .B(n2554), .Z(n2583) );
  OR U2662 ( .A(n2556), .B(b[1]), .Z(n2560) );
  NAND U2663 ( .A(n2558), .B(n2557), .Z(n2559) );
  NAND U2664 ( .A(n2560), .B(n2559), .Z(n2588) );
  NAND U2665 ( .A(a[58]), .B(b[7]), .Z(n2599) );
  NANDN U2666 ( .A(n247), .B(n2561), .Z(n2565) );
  NAND U2667 ( .A(n2563), .B(n2562), .Z(n2564) );
  NAND U2668 ( .A(n2565), .B(n2564), .Z(n2597) );
  XNOR U2669 ( .A(n2597), .B(n2636), .Z(n2598) );
  XNOR U2670 ( .A(n2599), .B(n2598), .Z(n2594) );
  NAND U2671 ( .A(n2566), .B(n2666), .Z(n2568) );
  XNOR U2672 ( .A(n2695), .B(a[60]), .Z(n2604) );
  NAND U2673 ( .A(n2604), .B(n2665), .Z(n2567) );
  NAND U2674 ( .A(n2568), .B(n2567), .Z(n2592) );
  XOR U2675 ( .A(a[62]), .B(n248), .Z(n2607) );
  OR U2676 ( .A(n2607), .B(n2608), .Z(n2571) );
  NANDN U2677 ( .A(n2569), .B(n2625), .Z(n2570) );
  AND U2678 ( .A(n2571), .B(n2570), .Z(n2591) );
  XNOR U2679 ( .A(n2592), .B(n2591), .Z(n2593) );
  XOR U2680 ( .A(n2594), .B(n2593), .Z(n2585) );
  NANDN U2681 ( .A(n2572), .B(n2636), .Z(n2576) );
  OR U2682 ( .A(n2574), .B(n2573), .Z(n2575) );
  NAND U2683 ( .A(n2576), .B(n2575), .Z(n2586) );
  XNOR U2684 ( .A(n2585), .B(n2586), .Z(n2587) );
  XOR U2685 ( .A(n2588), .B(n2587), .Z(n2582) );
  XNOR U2686 ( .A(n2583), .B(n2582), .Z(n2577) );
  XOR U2687 ( .A(n2584), .B(n2577), .Z(n2580) );
  OR U2688 ( .A(n2579), .B(n2578), .Z(n2581) );
  XNOR U2689 ( .A(n2580), .B(n2581), .Z(c[122]) );
  NANDN U2690 ( .A(n2581), .B(n2580), .Z(n2612) );
  NANDN U2691 ( .A(n2586), .B(n2585), .Z(n2590) );
  NAND U2692 ( .A(n2588), .B(n2587), .Z(n2589) );
  NAND U2693 ( .A(n2590), .B(n2589), .Z(n2614) );
  NANDN U2694 ( .A(n2592), .B(n2591), .Z(n2596) );
  NANDN U2695 ( .A(n2594), .B(n2593), .Z(n2595) );
  NAND U2696 ( .A(n2596), .B(n2595), .Z(n2643) );
  NANDN U2697 ( .A(n2597), .B(n2636), .Z(n2601) );
  NAND U2698 ( .A(n2599), .B(n2598), .Z(n2600) );
  NAND U2699 ( .A(n2601), .B(n2600), .Z(n2640) );
  NANDN U2700 ( .A(n2695), .B(a[59]), .Z(n2634) );
  NANDN U2701 ( .A(n2602), .B(b[1]), .Z(n2603) );
  ANDN U2702 ( .B(n2603), .A(n247), .Z(n2635) );
  XOR U2703 ( .A(n2634), .B(n2635), .Z(n2637) );
  XNOR U2704 ( .A(n2636), .B(n2637), .Z(n2621) );
  NAND U2705 ( .A(n2604), .B(n2666), .Z(n2606) );
  XNOR U2706 ( .A(n2695), .B(a[61]), .Z(n2630) );
  NAND U2707 ( .A(n2630), .B(n2665), .Z(n2605) );
  NAND U2708 ( .A(n2606), .B(n2605), .Z(n2619) );
  NANDN U2709 ( .A(n2607), .B(n2625), .Z(n2610) );
  XOR U2710 ( .A(b[5]), .B(n2696), .Z(n2626) );
  OR U2711 ( .A(n2626), .B(n2608), .Z(n2609) );
  AND U2712 ( .A(n2610), .B(n2609), .Z(n2620) );
  XOR U2713 ( .A(n2619), .B(n2620), .Z(n2622) );
  XOR U2714 ( .A(n2621), .B(n2622), .Z(n2641) );
  XNOR U2715 ( .A(n2640), .B(n2641), .Z(n2642) );
  XOR U2716 ( .A(n2643), .B(n2642), .Z(n2613) );
  XOR U2717 ( .A(n2614), .B(n2613), .Z(n2616) );
  XOR U2718 ( .A(n2615), .B(n2616), .Z(n2611) );
  XOR U2719 ( .A(n2612), .B(n2611), .Z(c[123]) );
  OR U2720 ( .A(n2612), .B(n2611), .Z(n2672) );
  NANDN U2721 ( .A(n2614), .B(n2613), .Z(n2618) );
  OR U2722 ( .A(n2616), .B(n2615), .Z(n2617) );
  NAND U2723 ( .A(n2618), .B(n2617), .Z(n2649) );
  NANDN U2724 ( .A(n2620), .B(n2619), .Z(n2624) );
  OR U2725 ( .A(n2622), .B(n2621), .Z(n2623) );
  NAND U2726 ( .A(n2624), .B(n2623), .Z(n2655) );
  NANDN U2727 ( .A(n2626), .B(n2625), .Z(n2627) );
  NANDN U2728 ( .A(n2628), .B(n2627), .Z(n2660) );
  ANDN U2729 ( .B(b[7]), .A(n2629), .Z(n2682) );
  XOR U2730 ( .A(n2660), .B(n2682), .Z(n2662) );
  NAND U2731 ( .A(n2630), .B(n2666), .Z(n2633) );
  XOR U2732 ( .A(b[7]), .B(n2631), .Z(n2667) );
  NANDN U2733 ( .A(n2667), .B(n2665), .Z(n2632) );
  NAND U2734 ( .A(n2633), .B(n2632), .Z(n2661) );
  XNOR U2735 ( .A(n2662), .B(n2661), .Z(n2652) );
  OR U2736 ( .A(n2635), .B(n2634), .Z(n2639) );
  NAND U2737 ( .A(n2637), .B(n2636), .Z(n2638) );
  AND U2738 ( .A(n2639), .B(n2638), .Z(n2653) );
  XNOR U2739 ( .A(n2652), .B(n2653), .Z(n2654) );
  XNOR U2740 ( .A(n2655), .B(n2654), .Z(n2646) );
  NANDN U2741 ( .A(n2641), .B(n2640), .Z(n2645) );
  NAND U2742 ( .A(n2643), .B(n2642), .Z(n2644) );
  AND U2743 ( .A(n2645), .B(n2644), .Z(n2647) );
  XNOR U2744 ( .A(n2646), .B(n2647), .Z(n2648) );
  XOR U2745 ( .A(n2649), .B(n2648), .Z(n2671) );
  XOR U2746 ( .A(n2672), .B(n2671), .Z(c[124]) );
  NANDN U2747 ( .A(n2647), .B(n2646), .Z(n2651) );
  NAND U2748 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U2749 ( .A(n2651), .B(n2650), .Z(n2688) );
  NANDN U2750 ( .A(n2653), .B(n2652), .Z(n2657) );
  NAND U2751 ( .A(n2655), .B(n2654), .Z(n2656) );
  NAND U2752 ( .A(n2657), .B(n2656), .Z(n2686) );
  NANDN U2753 ( .A(n2695), .B(a[61]), .Z(n2681) );
  NANDN U2754 ( .A(n2658), .B(b[3]), .Z(n2659) );
  ANDN U2755 ( .B(n2659), .A(n248), .Z(n2680) );
  XNOR U2756 ( .A(n2681), .B(n2680), .Z(n2683) );
  XOR U2757 ( .A(n2682), .B(n2683), .Z(n2692) );
  NANDN U2758 ( .A(n2660), .B(n2682), .Z(n2664) );
  OR U2759 ( .A(n2662), .B(n2661), .Z(n2663) );
  NAND U2760 ( .A(n2664), .B(n2663), .Z(n2689) );
  XNOR U2761 ( .A(b[7]), .B(a[63]), .Z(n2676) );
  NANDN U2762 ( .A(n2676), .B(n2665), .Z(n2669) );
  NANDN U2763 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U2764 ( .A(n2669), .B(n2668), .Z(n2690) );
  XNOR U2765 ( .A(n2689), .B(n2690), .Z(n2691) );
  XOR U2766 ( .A(n2686), .B(n2687), .Z(n2670) );
  XNOR U2767 ( .A(n2688), .B(n2670), .Z(n2674) );
  OR U2768 ( .A(n2672), .B(n2671), .Z(n2673) );
  XOR U2769 ( .A(n2674), .B(n2673), .Z(c[125]) );
  OR U2770 ( .A(n2674), .B(n2673), .Z(n2708) );
  NANDN U2771 ( .A(n248), .B(b[6]), .Z(n2675) );
  XOR U2772 ( .A(n2695), .B(n2675), .Z(n2679) );
  XOR U2773 ( .A(b[6]), .B(n248), .Z(n2677) );
  NAND U2774 ( .A(n2677), .B(n2676), .Z(n2678) );
  AND U2775 ( .A(n2679), .B(n2678), .Z(n2714) );
  NANDN U2776 ( .A(n2695), .B(a[62]), .Z(n2716) );
  OR U2777 ( .A(n2681), .B(n2680), .Z(n2685) );
  NANDN U2778 ( .A(n2683), .B(n2682), .Z(n2684) );
  AND U2779 ( .A(n2685), .B(n2684), .Z(n2715) );
  XNOR U2780 ( .A(n2716), .B(n2715), .Z(n2713) );
  XNOR U2781 ( .A(n2714), .B(n2713), .Z(n2703) );
  OR U2782 ( .A(n2690), .B(n2689), .Z(n2694) );
  OR U2783 ( .A(n2692), .B(n2691), .Z(n2693) );
  NAND U2784 ( .A(n2694), .B(n2693), .Z(n2701) );
  XOR U2785 ( .A(n2702), .B(n2701), .Z(n2704) );
  XOR U2786 ( .A(n2703), .B(n2704), .Z(n2707) );
  XOR U2787 ( .A(n2708), .B(n2707), .Z(c[126]) );
  NANDN U2788 ( .A(b[5]), .B(n2695), .Z(n2697) );
  ANDN U2789 ( .B(n2697), .A(n2696), .Z(n2700) );
  XNOR U2790 ( .A(n248), .B(b[7]), .Z(n2698) );
  NANDN U2791 ( .A(b[6]), .B(n2698), .Z(n2699) );
  NAND U2792 ( .A(n2700), .B(n2699), .Z(n2712) );
  NOR U2793 ( .A(n2702), .B(n2701), .Z(n2706) );
  AND U2794 ( .A(n2704), .B(n2703), .Z(n2705) );
  OR U2795 ( .A(n2706), .B(n2705), .Z(n2710) );
  OR U2796 ( .A(n2708), .B(n2707), .Z(n2709) );
  NAND U2797 ( .A(n2710), .B(n2709), .Z(n2711) );
  XNOR U2798 ( .A(n2712), .B(n2711), .Z(n2720) );
  OR U2799 ( .A(n2714), .B(n2713), .Z(n2718) );
  OR U2800 ( .A(n2716), .B(n2715), .Z(n2717) );
  NAND U2801 ( .A(n2718), .B(n2717), .Z(n2719) );
  XNOR U2802 ( .A(n2720), .B(n2719), .Z(c[127]) );
endmodule

