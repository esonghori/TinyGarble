
module Bus_Mux ( imm_in, reg_source, a_mux, a_out, reg_target, b_mux, b_out, 
        c_bus, c_memory, c_pc, c_pc_plus4, c_mux, reg_dest_out, branch_func, 
        take_branch );
  input [15:0] imm_in;
  input [31:0] reg_source;
  input [1:0] a_mux;
  output [31:0] a_out;
  input [31:0] reg_target;
  input [1:0] b_mux;
  output [31:0] b_out;
  input [31:0] c_bus;
  input [31:0] c_memory;
  input [31:2] c_pc;
  input [31:2] c_pc_plus4;
  input [2:0] c_mux;
  output [31:0] reg_dest_out;
  input [2:0] branch_func;
  output take_branch;
  wire   n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006;

  NAND U606 ( .A(n507), .B(n508), .Z(take_branch) );
  AND U607 ( .A(n509), .B(n510), .Z(n508) );
  OR U608 ( .A(n511), .B(n512), .Z(n510) );
  MUX U609 ( .IN0(n513), .IN1(n514), .SEL(n515), .F(n509) );
  OR U610 ( .A(n516), .B(branch_func[0]), .Z(n513) );
  AND U611 ( .A(n517), .B(n518), .Z(n507) );
  MUX U612 ( .IN0(n519), .IN1(n514), .SEL(n520), .F(n518) );
  IV U613 ( .A(branch_func[0]), .Z(n520) );
  OR U614 ( .A(n521), .B(c_bus[31]), .Z(n514) );
  OR U615 ( .A(branch_func[1]), .B(n522), .Z(n521) );
  OR U616 ( .A(n515), .B(n511), .Z(n519) );
  OR U617 ( .A(branch_func[1]), .B(branch_func[2]), .Z(n511) );
  MUX U618 ( .IN0(n523), .IN1(n524), .SEL(branch_func[0]), .F(n517) );
  NANDN U619 ( .A(n516), .B(n515), .Z(n524) );
  NAND U620 ( .A(n525), .B(n526), .Z(n515) );
  AND U621 ( .A(n527), .B(n528), .Z(n526) );
  AND U622 ( .A(n529), .B(n530), .Z(n528) );
  AND U623 ( .A(n531), .B(n532), .Z(n530) );
  NOR U624 ( .A(c_bus[9]), .B(c_bus[8]), .Z(n532) );
  NOR U625 ( .A(c_bus[7]), .B(c_bus[6]), .Z(n531) );
  AND U626 ( .A(n533), .B(n534), .Z(n529) );
  NOR U627 ( .A(c_bus[5]), .B(c_bus[4]), .Z(n534) );
  ANDN U628 ( .B(n512), .A(c_bus[3]), .Z(n533) );
  AND U629 ( .A(n535), .B(n536), .Z(n527) );
  AND U630 ( .A(n537), .B(n538), .Z(n536) );
  NOR U631 ( .A(c_bus[30]), .B(c_bus[2]), .Z(n538) );
  NOR U632 ( .A(c_bus[29]), .B(c_bus[28]), .Z(n537) );
  AND U633 ( .A(n539), .B(n540), .Z(n535) );
  NOR U634 ( .A(c_bus[27]), .B(c_bus[26]), .Z(n540) );
  NOR U635 ( .A(c_bus[25]), .B(c_bus[24]), .Z(n539) );
  AND U636 ( .A(n541), .B(n542), .Z(n525) );
  AND U637 ( .A(n543), .B(n544), .Z(n542) );
  AND U638 ( .A(n545), .B(n546), .Z(n544) );
  NOR U639 ( .A(c_bus[23]), .B(c_bus[22]), .Z(n546) );
  NOR U640 ( .A(c_bus[21]), .B(c_bus[20]), .Z(n545) );
  AND U641 ( .A(n547), .B(n548), .Z(n543) );
  NOR U642 ( .A(c_bus[1]), .B(c_bus[19]), .Z(n548) );
  NOR U643 ( .A(c_bus[18]), .B(c_bus[17]), .Z(n547) );
  AND U644 ( .A(n549), .B(n550), .Z(n541) );
  AND U645 ( .A(n551), .B(n552), .Z(n550) );
  NOR U646 ( .A(c_bus[16]), .B(c_bus[15]), .Z(n552) );
  NOR U647 ( .A(c_bus[14]), .B(c_bus[13]), .Z(n551) );
  AND U648 ( .A(n553), .B(n554), .Z(n549) );
  NOR U649 ( .A(c_bus[12]), .B(c_bus[11]), .Z(n554) );
  NOR U650 ( .A(c_bus[10]), .B(c_bus[0]), .Z(n553) );
  NANDN U651 ( .A(branch_func[2]), .B(branch_func[1]), .Z(n516) );
  NANDN U652 ( .A(n522), .B(branch_func[1]), .Z(n523) );
  IV U653 ( .A(branch_func[2]), .Z(n522) );
  NAND U654 ( .A(n555), .B(n556), .Z(reg_dest_out[9]) );
  AND U655 ( .A(n557), .B(n558), .Z(n556) );
  NAND U656 ( .A(n559), .B(c_pc[9]), .Z(n558) );
  AND U657 ( .A(n560), .B(n561), .Z(n557) );
  NAND U658 ( .A(n562), .B(c_bus[9]), .Z(n561) );
  NAND U659 ( .A(n563), .B(c_memory[9]), .Z(n560) );
  AND U660 ( .A(n564), .B(n565), .Z(n555) );
  NAND U661 ( .A(n566), .B(c_pc_plus4[9]), .Z(n565) );
  NAND U662 ( .A(n567), .B(reg_source[9]), .Z(n564) );
  NAND U663 ( .A(n568), .B(n569), .Z(reg_dest_out[8]) );
  AND U664 ( .A(n570), .B(n571), .Z(n569) );
  NAND U665 ( .A(n559), .B(c_pc[8]), .Z(n571) );
  AND U666 ( .A(n572), .B(n573), .Z(n570) );
  NAND U667 ( .A(n562), .B(c_bus[8]), .Z(n573) );
  NAND U668 ( .A(n563), .B(c_memory[8]), .Z(n572) );
  AND U669 ( .A(n574), .B(n575), .Z(n568) );
  NAND U670 ( .A(n566), .B(c_pc_plus4[8]), .Z(n575) );
  NAND U671 ( .A(n567), .B(reg_source[8]), .Z(n574) );
  NAND U672 ( .A(n576), .B(n577), .Z(reg_dest_out[7]) );
  AND U673 ( .A(n578), .B(n579), .Z(n577) );
  NAND U674 ( .A(n559), .B(c_pc[7]), .Z(n579) );
  AND U675 ( .A(n580), .B(n581), .Z(n578) );
  NAND U676 ( .A(n562), .B(c_bus[7]), .Z(n581) );
  NAND U677 ( .A(n563), .B(c_memory[7]), .Z(n580) );
  AND U678 ( .A(n582), .B(n583), .Z(n576) );
  NAND U679 ( .A(n566), .B(c_pc_plus4[7]), .Z(n583) );
  NAND U680 ( .A(n567), .B(reg_source[7]), .Z(n582) );
  NAND U681 ( .A(n584), .B(n585), .Z(reg_dest_out[6]) );
  AND U682 ( .A(n586), .B(n587), .Z(n585) );
  NAND U683 ( .A(n559), .B(c_pc[6]), .Z(n587) );
  AND U684 ( .A(n588), .B(n589), .Z(n586) );
  NAND U685 ( .A(n562), .B(c_bus[6]), .Z(n589) );
  NAND U686 ( .A(n563), .B(c_memory[6]), .Z(n588) );
  AND U687 ( .A(n590), .B(n591), .Z(n584) );
  NAND U688 ( .A(n566), .B(c_pc_plus4[6]), .Z(n591) );
  NAND U689 ( .A(n567), .B(reg_source[6]), .Z(n590) );
  NAND U690 ( .A(n592), .B(n593), .Z(reg_dest_out[5]) );
  AND U691 ( .A(n594), .B(n595), .Z(n593) );
  NAND U692 ( .A(n559), .B(c_pc[5]), .Z(n595) );
  AND U693 ( .A(n596), .B(n597), .Z(n594) );
  NAND U694 ( .A(n562), .B(c_bus[5]), .Z(n597) );
  NAND U695 ( .A(n563), .B(c_memory[5]), .Z(n596) );
  AND U696 ( .A(n598), .B(n599), .Z(n592) );
  NAND U697 ( .A(n566), .B(c_pc_plus4[5]), .Z(n599) );
  NAND U698 ( .A(n567), .B(reg_source[5]), .Z(n598) );
  NAND U699 ( .A(n600), .B(n601), .Z(reg_dest_out[4]) );
  AND U700 ( .A(n602), .B(n603), .Z(n601) );
  NAND U701 ( .A(n559), .B(c_pc[4]), .Z(n603) );
  AND U702 ( .A(n604), .B(n605), .Z(n602) );
  NAND U703 ( .A(n562), .B(c_bus[4]), .Z(n605) );
  NAND U704 ( .A(n563), .B(c_memory[4]), .Z(n604) );
  AND U705 ( .A(n606), .B(n607), .Z(n600) );
  NAND U706 ( .A(n566), .B(c_pc_plus4[4]), .Z(n607) );
  NAND U707 ( .A(n567), .B(reg_source[4]), .Z(n606) );
  NAND U708 ( .A(n608), .B(n609), .Z(reg_dest_out[3]) );
  AND U709 ( .A(n610), .B(n611), .Z(n609) );
  NAND U710 ( .A(n559), .B(c_pc[3]), .Z(n611) );
  AND U711 ( .A(n612), .B(n613), .Z(n610) );
  NAND U712 ( .A(n562), .B(c_bus[3]), .Z(n613) );
  NAND U713 ( .A(n563), .B(c_memory[3]), .Z(n612) );
  AND U714 ( .A(n614), .B(n615), .Z(n608) );
  NAND U715 ( .A(n566), .B(c_pc_plus4[3]), .Z(n615) );
  NAND U716 ( .A(n567), .B(reg_source[3]), .Z(n614) );
  NAND U717 ( .A(n616), .B(n617), .Z(reg_dest_out[31]) );
  AND U718 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U719 ( .A(n512), .B(n562), .Z(n619) );
  IV U720 ( .A(c_bus[31]), .Z(n512) );
  AND U721 ( .A(n620), .B(n621), .Z(n618) );
  NAND U722 ( .A(n563), .B(c_memory[31]), .Z(n621) );
  NAND U723 ( .A(n567), .B(reg_source[31]), .Z(n620) );
  AND U724 ( .A(n622), .B(n623), .Z(n616) );
  NAND U725 ( .A(n559), .B(c_pc[31]), .Z(n623) );
  AND U726 ( .A(n624), .B(n625), .Z(n622) );
  NAND U727 ( .A(n566), .B(c_pc_plus4[31]), .Z(n625) );
  NANDN U728 ( .A(n626), .B(n627), .Z(n624) );
  NAND U729 ( .A(n628), .B(n629), .Z(reg_dest_out[30]) );
  AND U730 ( .A(n630), .B(n631), .Z(n629) );
  NAND U731 ( .A(n562), .B(c_bus[30]), .Z(n631) );
  AND U732 ( .A(n632), .B(n633), .Z(n630) );
  NAND U733 ( .A(n563), .B(c_memory[30]), .Z(n633) );
  NAND U734 ( .A(n567), .B(reg_source[30]), .Z(n632) );
  AND U735 ( .A(n634), .B(n635), .Z(n628) );
  NAND U736 ( .A(n559), .B(c_pc[30]), .Z(n635) );
  AND U737 ( .A(n636), .B(n637), .Z(n634) );
  NAND U738 ( .A(n566), .B(c_pc_plus4[30]), .Z(n637) );
  NAND U739 ( .A(n627), .B(imm_in[14]), .Z(n636) );
  NAND U740 ( .A(n638), .B(n639), .Z(reg_dest_out[2]) );
  AND U741 ( .A(n640), .B(n641), .Z(n639) );
  NAND U742 ( .A(n559), .B(c_pc[2]), .Z(n641) );
  AND U743 ( .A(n642), .B(n643), .Z(n640) );
  NAND U744 ( .A(n562), .B(c_bus[2]), .Z(n643) );
  NAND U745 ( .A(n563), .B(c_memory[2]), .Z(n642) );
  AND U746 ( .A(n644), .B(n645), .Z(n638) );
  NAND U747 ( .A(n566), .B(c_pc_plus4[2]), .Z(n645) );
  NAND U748 ( .A(n567), .B(reg_source[2]), .Z(n644) );
  NAND U749 ( .A(n646), .B(n647), .Z(reg_dest_out[29]) );
  AND U750 ( .A(n648), .B(n649), .Z(n647) );
  NAND U751 ( .A(n562), .B(c_bus[29]), .Z(n649) );
  AND U752 ( .A(n650), .B(n651), .Z(n648) );
  NAND U753 ( .A(n563), .B(c_memory[29]), .Z(n651) );
  NAND U754 ( .A(n567), .B(reg_source[29]), .Z(n650) );
  AND U755 ( .A(n652), .B(n653), .Z(n646) );
  NAND U756 ( .A(n559), .B(c_pc[29]), .Z(n653) );
  AND U757 ( .A(n654), .B(n655), .Z(n652) );
  NAND U758 ( .A(n566), .B(c_pc_plus4[29]), .Z(n655) );
  NAND U759 ( .A(n627), .B(imm_in[13]), .Z(n654) );
  NAND U760 ( .A(n656), .B(n657), .Z(reg_dest_out[28]) );
  AND U761 ( .A(n658), .B(n659), .Z(n657) );
  NAND U762 ( .A(n562), .B(c_bus[28]), .Z(n659) );
  AND U763 ( .A(n660), .B(n661), .Z(n658) );
  NAND U764 ( .A(n563), .B(c_memory[28]), .Z(n661) );
  NAND U765 ( .A(n567), .B(reg_source[28]), .Z(n660) );
  AND U766 ( .A(n662), .B(n663), .Z(n656) );
  NAND U767 ( .A(n559), .B(c_pc[28]), .Z(n663) );
  AND U768 ( .A(n664), .B(n665), .Z(n662) );
  NAND U769 ( .A(n566), .B(c_pc_plus4[28]), .Z(n665) );
  NAND U770 ( .A(n627), .B(imm_in[12]), .Z(n664) );
  NAND U771 ( .A(n666), .B(n667), .Z(reg_dest_out[27]) );
  AND U772 ( .A(n668), .B(n669), .Z(n667) );
  NAND U773 ( .A(n562), .B(c_bus[27]), .Z(n669) );
  AND U774 ( .A(n670), .B(n671), .Z(n668) );
  NAND U775 ( .A(n563), .B(c_memory[27]), .Z(n671) );
  NAND U776 ( .A(n567), .B(reg_source[27]), .Z(n670) );
  AND U777 ( .A(n672), .B(n673), .Z(n666) );
  NAND U778 ( .A(n559), .B(c_pc[27]), .Z(n673) );
  AND U779 ( .A(n674), .B(n675), .Z(n672) );
  NAND U780 ( .A(n566), .B(c_pc_plus4[27]), .Z(n675) );
  NAND U781 ( .A(n627), .B(imm_in[11]), .Z(n674) );
  NAND U782 ( .A(n676), .B(n677), .Z(reg_dest_out[26]) );
  AND U783 ( .A(n678), .B(n679), .Z(n677) );
  NAND U784 ( .A(n562), .B(c_bus[26]), .Z(n679) );
  AND U785 ( .A(n680), .B(n681), .Z(n678) );
  NAND U786 ( .A(n563), .B(c_memory[26]), .Z(n681) );
  NAND U787 ( .A(n567), .B(reg_source[26]), .Z(n680) );
  AND U788 ( .A(n682), .B(n683), .Z(n676) );
  NAND U789 ( .A(n559), .B(c_pc[26]), .Z(n683) );
  AND U790 ( .A(n684), .B(n685), .Z(n682) );
  NAND U791 ( .A(n566), .B(c_pc_plus4[26]), .Z(n685) );
  NAND U792 ( .A(n627), .B(imm_in[10]), .Z(n684) );
  NAND U793 ( .A(n686), .B(n687), .Z(reg_dest_out[25]) );
  AND U794 ( .A(n688), .B(n689), .Z(n687) );
  NAND U795 ( .A(n562), .B(c_bus[25]), .Z(n689) );
  AND U796 ( .A(n690), .B(n691), .Z(n688) );
  NAND U797 ( .A(n563), .B(c_memory[25]), .Z(n691) );
  NAND U798 ( .A(n567), .B(reg_source[25]), .Z(n690) );
  AND U799 ( .A(n692), .B(n693), .Z(n686) );
  NAND U800 ( .A(n559), .B(c_pc[25]), .Z(n693) );
  AND U801 ( .A(n694), .B(n695), .Z(n692) );
  NAND U802 ( .A(n566), .B(c_pc_plus4[25]), .Z(n695) );
  NAND U803 ( .A(n627), .B(imm_in[9]), .Z(n694) );
  NAND U804 ( .A(n696), .B(n697), .Z(reg_dest_out[24]) );
  AND U805 ( .A(n698), .B(n699), .Z(n697) );
  NAND U806 ( .A(n562), .B(c_bus[24]), .Z(n699) );
  AND U807 ( .A(n700), .B(n701), .Z(n698) );
  NAND U808 ( .A(n563), .B(c_memory[24]), .Z(n701) );
  NAND U809 ( .A(n567), .B(reg_source[24]), .Z(n700) );
  AND U810 ( .A(n702), .B(n703), .Z(n696) );
  NAND U811 ( .A(n559), .B(c_pc[24]), .Z(n703) );
  AND U812 ( .A(n704), .B(n705), .Z(n702) );
  NAND U813 ( .A(n566), .B(c_pc_plus4[24]), .Z(n705) );
  NAND U814 ( .A(n627), .B(imm_in[8]), .Z(n704) );
  NAND U815 ( .A(n706), .B(n707), .Z(reg_dest_out[23]) );
  AND U816 ( .A(n708), .B(n709), .Z(n707) );
  NAND U817 ( .A(n562), .B(c_bus[23]), .Z(n709) );
  AND U818 ( .A(n710), .B(n711), .Z(n708) );
  NAND U819 ( .A(n563), .B(c_memory[23]), .Z(n711) );
  NAND U820 ( .A(n567), .B(reg_source[23]), .Z(n710) );
  AND U821 ( .A(n712), .B(n713), .Z(n706) );
  NAND U822 ( .A(n559), .B(c_pc[23]), .Z(n713) );
  AND U823 ( .A(n714), .B(n715), .Z(n712) );
  NAND U824 ( .A(n566), .B(c_pc_plus4[23]), .Z(n715) );
  NAND U825 ( .A(n627), .B(imm_in[7]), .Z(n714) );
  NAND U826 ( .A(n716), .B(n717), .Z(reg_dest_out[22]) );
  AND U827 ( .A(n718), .B(n719), .Z(n717) );
  NAND U828 ( .A(n562), .B(c_bus[22]), .Z(n719) );
  AND U829 ( .A(n720), .B(n721), .Z(n718) );
  NAND U830 ( .A(n563), .B(c_memory[22]), .Z(n721) );
  NAND U831 ( .A(n567), .B(reg_source[22]), .Z(n720) );
  AND U832 ( .A(n722), .B(n723), .Z(n716) );
  NAND U833 ( .A(n559), .B(c_pc[22]), .Z(n723) );
  AND U834 ( .A(n724), .B(n725), .Z(n722) );
  NAND U835 ( .A(n566), .B(c_pc_plus4[22]), .Z(n725) );
  NAND U836 ( .A(n627), .B(imm_in[6]), .Z(n724) );
  NAND U837 ( .A(n726), .B(n727), .Z(reg_dest_out[21]) );
  AND U838 ( .A(n728), .B(n729), .Z(n727) );
  NAND U839 ( .A(n562), .B(c_bus[21]), .Z(n729) );
  AND U840 ( .A(n730), .B(n731), .Z(n728) );
  NAND U841 ( .A(n563), .B(c_memory[21]), .Z(n731) );
  NAND U842 ( .A(n567), .B(reg_source[21]), .Z(n730) );
  AND U843 ( .A(n732), .B(n733), .Z(n726) );
  NAND U844 ( .A(n559), .B(c_pc[21]), .Z(n733) );
  AND U845 ( .A(n734), .B(n735), .Z(n732) );
  NAND U846 ( .A(n566), .B(c_pc_plus4[21]), .Z(n735) );
  NAND U847 ( .A(n627), .B(imm_in[5]), .Z(n734) );
  NAND U848 ( .A(n736), .B(n737), .Z(reg_dest_out[20]) );
  AND U849 ( .A(n738), .B(n739), .Z(n737) );
  NAND U850 ( .A(n562), .B(c_bus[20]), .Z(n739) );
  AND U851 ( .A(n740), .B(n741), .Z(n738) );
  NAND U852 ( .A(n563), .B(c_memory[20]), .Z(n741) );
  NAND U853 ( .A(n567), .B(reg_source[20]), .Z(n740) );
  AND U854 ( .A(n742), .B(n743), .Z(n736) );
  NAND U855 ( .A(n559), .B(c_pc[20]), .Z(n743) );
  AND U856 ( .A(n744), .B(n745), .Z(n742) );
  NAND U857 ( .A(n566), .B(c_pc_plus4[20]), .Z(n745) );
  NAND U858 ( .A(n627), .B(imm_in[4]), .Z(n744) );
  NAND U859 ( .A(n746), .B(n747), .Z(reg_dest_out[1]) );
  NAND U860 ( .A(n562), .B(c_bus[1]), .Z(n747) );
  AND U861 ( .A(n748), .B(n749), .Z(n746) );
  NAND U862 ( .A(n563), .B(c_memory[1]), .Z(n749) );
  NAND U863 ( .A(n567), .B(reg_source[1]), .Z(n748) );
  NAND U864 ( .A(n750), .B(n751), .Z(reg_dest_out[19]) );
  AND U865 ( .A(n752), .B(n753), .Z(n751) );
  NAND U866 ( .A(n562), .B(c_bus[19]), .Z(n753) );
  AND U867 ( .A(n754), .B(n755), .Z(n752) );
  NAND U868 ( .A(n563), .B(c_memory[19]), .Z(n755) );
  NAND U869 ( .A(n567), .B(reg_source[19]), .Z(n754) );
  AND U870 ( .A(n756), .B(n757), .Z(n750) );
  NAND U871 ( .A(n559), .B(c_pc[19]), .Z(n757) );
  AND U872 ( .A(n758), .B(n759), .Z(n756) );
  NAND U873 ( .A(n566), .B(c_pc_plus4[19]), .Z(n759) );
  NAND U874 ( .A(n627), .B(imm_in[3]), .Z(n758) );
  NAND U875 ( .A(n760), .B(n761), .Z(reg_dest_out[18]) );
  AND U876 ( .A(n762), .B(n763), .Z(n761) );
  NAND U877 ( .A(n562), .B(c_bus[18]), .Z(n763) );
  AND U878 ( .A(n764), .B(n765), .Z(n762) );
  NAND U879 ( .A(n563), .B(c_memory[18]), .Z(n765) );
  NAND U880 ( .A(n567), .B(reg_source[18]), .Z(n764) );
  AND U881 ( .A(n766), .B(n767), .Z(n760) );
  NAND U882 ( .A(n559), .B(c_pc[18]), .Z(n767) );
  AND U883 ( .A(n768), .B(n769), .Z(n766) );
  NAND U884 ( .A(n566), .B(c_pc_plus4[18]), .Z(n769) );
  NAND U885 ( .A(n627), .B(imm_in[2]), .Z(n768) );
  NAND U886 ( .A(n770), .B(n771), .Z(reg_dest_out[17]) );
  AND U887 ( .A(n772), .B(n773), .Z(n771) );
  NAND U888 ( .A(n562), .B(c_bus[17]), .Z(n773) );
  AND U889 ( .A(n774), .B(n775), .Z(n772) );
  NAND U890 ( .A(n563), .B(c_memory[17]), .Z(n775) );
  NAND U891 ( .A(n567), .B(reg_source[17]), .Z(n774) );
  AND U892 ( .A(n776), .B(n777), .Z(n770) );
  NAND U893 ( .A(n559), .B(c_pc[17]), .Z(n777) );
  AND U894 ( .A(n778), .B(n779), .Z(n776) );
  NAND U895 ( .A(n566), .B(c_pc_plus4[17]), .Z(n779) );
  NAND U896 ( .A(imm_in[1]), .B(n627), .Z(n778) );
  NAND U897 ( .A(n780), .B(n781), .Z(reg_dest_out[16]) );
  AND U898 ( .A(n782), .B(n783), .Z(n781) );
  NAND U899 ( .A(n562), .B(c_bus[16]), .Z(n783) );
  AND U900 ( .A(n784), .B(n785), .Z(n782) );
  NAND U901 ( .A(n563), .B(c_memory[16]), .Z(n785) );
  NAND U902 ( .A(n567), .B(reg_source[16]), .Z(n784) );
  AND U903 ( .A(n786), .B(n787), .Z(n780) );
  NAND U904 ( .A(n559), .B(c_pc[16]), .Z(n787) );
  AND U905 ( .A(n788), .B(n789), .Z(n786) );
  NAND U906 ( .A(n566), .B(c_pc_plus4[16]), .Z(n789) );
  NAND U907 ( .A(n627), .B(imm_in[0]), .Z(n788) );
  NOR U908 ( .A(n790), .B(n791), .Z(n627) );
  NAND U909 ( .A(n792), .B(n793), .Z(reg_dest_out[15]) );
  AND U910 ( .A(n794), .B(n795), .Z(n793) );
  NAND U911 ( .A(n559), .B(c_pc[15]), .Z(n795) );
  AND U912 ( .A(n796), .B(n797), .Z(n794) );
  NAND U913 ( .A(n562), .B(c_bus[15]), .Z(n797) );
  NAND U914 ( .A(n563), .B(c_memory[15]), .Z(n796) );
  AND U915 ( .A(n798), .B(n799), .Z(n792) );
  NAND U916 ( .A(n566), .B(c_pc_plus4[15]), .Z(n799) );
  NAND U917 ( .A(n567), .B(reg_source[15]), .Z(n798) );
  NAND U918 ( .A(n800), .B(n801), .Z(reg_dest_out[14]) );
  AND U919 ( .A(n802), .B(n803), .Z(n801) );
  NAND U920 ( .A(n559), .B(c_pc[14]), .Z(n803) );
  AND U921 ( .A(n804), .B(n805), .Z(n802) );
  NAND U922 ( .A(n562), .B(c_bus[14]), .Z(n805) );
  NAND U923 ( .A(n563), .B(c_memory[14]), .Z(n804) );
  AND U924 ( .A(n806), .B(n807), .Z(n800) );
  NAND U925 ( .A(n566), .B(c_pc_plus4[14]), .Z(n807) );
  NAND U926 ( .A(n567), .B(reg_source[14]), .Z(n806) );
  NAND U927 ( .A(n808), .B(n809), .Z(reg_dest_out[13]) );
  AND U928 ( .A(n810), .B(n811), .Z(n809) );
  NAND U929 ( .A(n559), .B(c_pc[13]), .Z(n811) );
  AND U930 ( .A(n812), .B(n813), .Z(n810) );
  NAND U931 ( .A(n562), .B(c_bus[13]), .Z(n813) );
  NAND U932 ( .A(n563), .B(c_memory[13]), .Z(n812) );
  AND U933 ( .A(n814), .B(n815), .Z(n808) );
  NAND U934 ( .A(n566), .B(c_pc_plus4[13]), .Z(n815) );
  NAND U935 ( .A(n567), .B(reg_source[13]), .Z(n814) );
  NAND U936 ( .A(n816), .B(n817), .Z(reg_dest_out[12]) );
  AND U937 ( .A(n818), .B(n819), .Z(n817) );
  NAND U938 ( .A(n559), .B(c_pc[12]), .Z(n819) );
  AND U939 ( .A(n820), .B(n821), .Z(n818) );
  NAND U940 ( .A(n562), .B(c_bus[12]), .Z(n821) );
  NAND U941 ( .A(n563), .B(c_memory[12]), .Z(n820) );
  AND U942 ( .A(n822), .B(n823), .Z(n816) );
  NAND U943 ( .A(n566), .B(c_pc_plus4[12]), .Z(n823) );
  NAND U944 ( .A(n567), .B(reg_source[12]), .Z(n822) );
  NAND U945 ( .A(n824), .B(n825), .Z(reg_dest_out[11]) );
  AND U946 ( .A(n826), .B(n827), .Z(n825) );
  NAND U947 ( .A(c_pc[11]), .B(n559), .Z(n827) );
  AND U948 ( .A(n828), .B(n829), .Z(n826) );
  NAND U949 ( .A(n562), .B(c_bus[11]), .Z(n829) );
  NAND U950 ( .A(n563), .B(c_memory[11]), .Z(n828) );
  AND U951 ( .A(n830), .B(n831), .Z(n824) );
  NAND U952 ( .A(c_pc_plus4[11]), .B(n566), .Z(n831) );
  NAND U953 ( .A(n567), .B(reg_source[11]), .Z(n830) );
  NAND U954 ( .A(n832), .B(n833), .Z(reg_dest_out[10]) );
  AND U955 ( .A(n834), .B(n835), .Z(n833) );
  NAND U956 ( .A(n559), .B(c_pc[10]), .Z(n835) );
  NOR U957 ( .A(n790), .B(n836), .Z(n559) );
  AND U958 ( .A(n837), .B(n838), .Z(n834) );
  NAND U959 ( .A(n562), .B(c_bus[10]), .Z(n838) );
  NAND U960 ( .A(c_memory[10]), .B(n563), .Z(n837) );
  AND U961 ( .A(n839), .B(n840), .Z(n832) );
  NAND U962 ( .A(n566), .B(c_pc_plus4[10]), .Z(n840) );
  NOR U963 ( .A(c_mux[0]), .B(n791), .Z(n566) );
  NANDN U964 ( .A(c_mux[1]), .B(c_mux[2]), .Z(n791) );
  NAND U965 ( .A(reg_source[10]), .B(n567), .Z(n839) );
  NAND U966 ( .A(n841), .B(n842), .Z(reg_dest_out[0]) );
  NAND U967 ( .A(n562), .B(c_bus[0]), .Z(n842) );
  ANDN U968 ( .B(n843), .A(n790), .Z(n562) );
  ANDN U969 ( .B(n844), .A(c_mux[2]), .Z(n843) );
  AND U970 ( .A(n845), .B(n846), .Z(n841) );
  NAND U971 ( .A(n563), .B(c_memory[0]), .Z(n846) );
  NOR U972 ( .A(c_mux[0]), .B(n836), .Z(n563) );
  NANDN U973 ( .A(c_mux[2]), .B(c_mux[1]), .Z(n836) );
  NAND U974 ( .A(n567), .B(reg_source[0]), .Z(n845) );
  AND U975 ( .A(n847), .B(c_mux[2]), .Z(n567) );
  ANDN U976 ( .B(n790), .A(n844), .Z(n847) );
  IV U977 ( .A(c_mux[1]), .Z(n844) );
  IV U978 ( .A(c_mux[0]), .Z(n790) );
  NAND U979 ( .A(n848), .B(n849), .Z(b_out[9]) );
  NAND U980 ( .A(n850), .B(reg_target[9]), .Z(n849) );
  AND U981 ( .A(n851), .B(n852), .Z(n848) );
  NAND U982 ( .A(n853), .B(imm_in[9]), .Z(n852) );
  NANDN U983 ( .A(n854), .B(imm_in[7]), .Z(n851) );
  NAND U984 ( .A(n855), .B(n856), .Z(b_out[8]) );
  NAND U985 ( .A(n850), .B(reg_target[8]), .Z(n856) );
  AND U986 ( .A(n857), .B(n858), .Z(n855) );
  NAND U987 ( .A(n853), .B(imm_in[8]), .Z(n858) );
  NANDN U988 ( .A(n854), .B(imm_in[6]), .Z(n857) );
  NAND U989 ( .A(n859), .B(n860), .Z(b_out[7]) );
  NAND U990 ( .A(n850), .B(reg_target[7]), .Z(n860) );
  AND U991 ( .A(n861), .B(n862), .Z(n859) );
  NAND U992 ( .A(n853), .B(imm_in[7]), .Z(n862) );
  NANDN U993 ( .A(n854), .B(imm_in[5]), .Z(n861) );
  NAND U994 ( .A(n863), .B(n864), .Z(b_out[6]) );
  NAND U995 ( .A(n850), .B(reg_target[6]), .Z(n864) );
  AND U996 ( .A(n865), .B(n866), .Z(n863) );
  NAND U997 ( .A(n853), .B(imm_in[6]), .Z(n866) );
  NANDN U998 ( .A(n854), .B(imm_in[4]), .Z(n865) );
  NAND U999 ( .A(n867), .B(n868), .Z(b_out[5]) );
  NAND U1000 ( .A(n850), .B(reg_target[5]), .Z(n868) );
  AND U1001 ( .A(n869), .B(n870), .Z(n867) );
  NAND U1002 ( .A(n853), .B(imm_in[5]), .Z(n870) );
  NANDN U1003 ( .A(n854), .B(imm_in[3]), .Z(n869) );
  NAND U1004 ( .A(n871), .B(n872), .Z(b_out[4]) );
  NAND U1005 ( .A(n850), .B(reg_target[4]), .Z(n872) );
  AND U1006 ( .A(n873), .B(n874), .Z(n871) );
  NAND U1007 ( .A(n853), .B(imm_in[4]), .Z(n874) );
  NANDN U1008 ( .A(n854), .B(imm_in[2]), .Z(n873) );
  NAND U1009 ( .A(n875), .B(n876), .Z(b_out[3]) );
  NAND U1010 ( .A(n850), .B(reg_target[3]), .Z(n876) );
  AND U1011 ( .A(n877), .B(n878), .Z(n875) );
  NAND U1012 ( .A(n853), .B(imm_in[3]), .Z(n878) );
  NANDN U1013 ( .A(n854), .B(imm_in[1]), .Z(n877) );
  NAND U1014 ( .A(n879), .B(n880), .Z(b_out[31]) );
  NAND U1015 ( .A(n850), .B(reg_target[31]), .Z(n879) );
  NAND U1016 ( .A(n881), .B(n880), .Z(b_out[30]) );
  NAND U1017 ( .A(n850), .B(reg_target[30]), .Z(n881) );
  NAND U1018 ( .A(n882), .B(n883), .Z(b_out[2]) );
  NAND U1019 ( .A(n850), .B(reg_target[2]), .Z(n883) );
  AND U1020 ( .A(n884), .B(n885), .Z(n882) );
  NAND U1021 ( .A(n853), .B(imm_in[2]), .Z(n885) );
  NANDN U1022 ( .A(n854), .B(imm_in[0]), .Z(n884) );
  NAND U1023 ( .A(n886), .B(n880), .Z(b_out[29]) );
  NAND U1024 ( .A(n850), .B(reg_target[29]), .Z(n886) );
  NAND U1025 ( .A(n887), .B(n880), .Z(b_out[28]) );
  NAND U1026 ( .A(n850), .B(reg_target[28]), .Z(n887) );
  NAND U1027 ( .A(n888), .B(n880), .Z(b_out[27]) );
  NAND U1028 ( .A(n850), .B(reg_target[27]), .Z(n888) );
  NAND U1029 ( .A(n889), .B(n880), .Z(b_out[26]) );
  NAND U1030 ( .A(n850), .B(reg_target[26]), .Z(n889) );
  NAND U1031 ( .A(n890), .B(n880), .Z(b_out[25]) );
  NAND U1032 ( .A(n850), .B(reg_target[25]), .Z(n890) );
  NAND U1033 ( .A(n891), .B(n880), .Z(b_out[24]) );
  NAND U1034 ( .A(n850), .B(reg_target[24]), .Z(n891) );
  NAND U1035 ( .A(n892), .B(n880), .Z(b_out[23]) );
  NAND U1036 ( .A(n850), .B(reg_target[23]), .Z(n892) );
  NAND U1037 ( .A(n893), .B(n880), .Z(b_out[22]) );
  NAND U1038 ( .A(n850), .B(reg_target[22]), .Z(n893) );
  NAND U1039 ( .A(n894), .B(n880), .Z(b_out[21]) );
  NAND U1040 ( .A(n850), .B(reg_target[21]), .Z(n894) );
  NAND U1041 ( .A(n895), .B(n880), .Z(b_out[20]) );
  NAND U1042 ( .A(n850), .B(reg_target[20]), .Z(n895) );
  NAND U1043 ( .A(n896), .B(n897), .Z(b_out[1]) );
  NAND U1044 ( .A(n853), .B(imm_in[1]), .Z(n897) );
  NAND U1045 ( .A(n850), .B(reg_target[1]), .Z(n896) );
  NAND U1046 ( .A(n898), .B(n880), .Z(b_out[19]) );
  NAND U1047 ( .A(n850), .B(reg_target[19]), .Z(n898) );
  NAND U1048 ( .A(n899), .B(n880), .Z(b_out[18]) );
  NAND U1049 ( .A(n850), .B(reg_target[18]), .Z(n899) );
  NAND U1050 ( .A(n900), .B(n901), .Z(b_out[17]) );
  NANDN U1051 ( .A(n626), .B(b_mux[1]), .Z(n901) );
  NAND U1052 ( .A(n850), .B(reg_target[17]), .Z(n900) );
  NAND U1053 ( .A(n902), .B(n903), .Z(b_out[16]) );
  NAND U1054 ( .A(n850), .B(reg_target[16]), .Z(n903) );
  AND U1055 ( .A(n880), .B(n904), .Z(n902) );
  NANDN U1056 ( .A(n854), .B(imm_in[14]), .Z(n904) );
  NANDN U1057 ( .A(n905), .B(imm_in[15]), .Z(n880) );
  NAND U1058 ( .A(n906), .B(n907), .Z(b_out[15]) );
  NAND U1059 ( .A(n850), .B(reg_target[15]), .Z(n907) );
  AND U1060 ( .A(n908), .B(n909), .Z(n906) );
  NANDN U1061 ( .A(n626), .B(n853), .Z(n909) );
  IV U1062 ( .A(imm_in[15]), .Z(n626) );
  NANDN U1063 ( .A(n854), .B(imm_in[13]), .Z(n908) );
  NAND U1064 ( .A(n910), .B(n911), .Z(b_out[14]) );
  NAND U1065 ( .A(n850), .B(reg_target[14]), .Z(n911) );
  AND U1066 ( .A(n912), .B(n913), .Z(n910) );
  NAND U1067 ( .A(n853), .B(imm_in[14]), .Z(n913) );
  NANDN U1068 ( .A(n854), .B(imm_in[12]), .Z(n912) );
  NAND U1069 ( .A(n914), .B(n915), .Z(b_out[13]) );
  NAND U1070 ( .A(n850), .B(reg_target[13]), .Z(n915) );
  AND U1071 ( .A(n916), .B(n917), .Z(n914) );
  NAND U1072 ( .A(n853), .B(imm_in[13]), .Z(n917) );
  NANDN U1073 ( .A(n854), .B(imm_in[11]), .Z(n916) );
  NAND U1074 ( .A(n918), .B(n919), .Z(b_out[12]) );
  NAND U1075 ( .A(n850), .B(reg_target[12]), .Z(n919) );
  AND U1076 ( .A(n920), .B(n921), .Z(n918) );
  NAND U1077 ( .A(n853), .B(imm_in[12]), .Z(n921) );
  NANDN U1078 ( .A(n854), .B(imm_in[10]), .Z(n920) );
  NAND U1079 ( .A(n922), .B(n923), .Z(b_out[11]) );
  NAND U1080 ( .A(n850), .B(reg_target[11]), .Z(n923) );
  AND U1081 ( .A(n924), .B(n925), .Z(n922) );
  NAND U1082 ( .A(n853), .B(imm_in[11]), .Z(n925) );
  NANDN U1083 ( .A(n854), .B(imm_in[9]), .Z(n924) );
  NAND U1084 ( .A(n926), .B(n927), .Z(b_out[10]) );
  NAND U1085 ( .A(reg_target[10]), .B(n850), .Z(n927) );
  AND U1086 ( .A(n928), .B(n929), .Z(n926) );
  NAND U1087 ( .A(n853), .B(imm_in[10]), .Z(n929) );
  NANDN U1088 ( .A(n854), .B(imm_in[8]), .Z(n928) );
  NAND U1089 ( .A(b_mux[1]), .B(b_mux[0]), .Z(n854) );
  NAND U1090 ( .A(n930), .B(n931), .Z(b_out[0]) );
  NAND U1091 ( .A(n853), .B(imm_in[0]), .Z(n931) );
  NAND U1092 ( .A(n932), .B(n905), .Z(n853) );
  NANDN U1093 ( .A(b_mux[0]), .B(b_mux[1]), .Z(n905) );
  NANDN U1094 ( .A(b_mux[1]), .B(b_mux[0]), .Z(n932) );
  NAND U1095 ( .A(n850), .B(reg_target[0]), .Z(n930) );
  NOR U1096 ( .A(b_mux[1]), .B(b_mux[0]), .Z(n850) );
  NAND U1097 ( .A(n933), .B(n934), .Z(a_out[9]) );
  NAND U1098 ( .A(c_pc[9]), .B(n935), .Z(n934) );
  NAND U1099 ( .A(reg_source[9]), .B(n936), .Z(n933) );
  NAND U1100 ( .A(n937), .B(n938), .Z(a_out[8]) );
  NAND U1101 ( .A(c_pc[8]), .B(n935), .Z(n938) );
  NAND U1102 ( .A(reg_source[8]), .B(n936), .Z(n937) );
  NAND U1103 ( .A(n939), .B(n940), .Z(a_out[7]) );
  NAND U1104 ( .A(c_pc[7]), .B(n935), .Z(n940) );
  NAND U1105 ( .A(reg_source[7]), .B(n936), .Z(n939) );
  NAND U1106 ( .A(n941), .B(n942), .Z(a_out[6]) );
  NAND U1107 ( .A(c_pc[6]), .B(n935), .Z(n942) );
  NAND U1108 ( .A(reg_source[6]), .B(n936), .Z(n941) );
  NAND U1109 ( .A(n943), .B(n944), .Z(a_out[5]) );
  NAND U1110 ( .A(c_pc[5]), .B(n935), .Z(n944) );
  NAND U1111 ( .A(reg_source[5]), .B(n936), .Z(n943) );
  NAND U1112 ( .A(n945), .B(n946), .Z(a_out[4]) );
  NAND U1113 ( .A(reg_source[4]), .B(n936), .Z(n946) );
  AND U1114 ( .A(n947), .B(n948), .Z(n945) );
  NANDN U1115 ( .A(n949), .B(imm_in[10]), .Z(n948) );
  NAND U1116 ( .A(c_pc[4]), .B(n935), .Z(n947) );
  NAND U1117 ( .A(n950), .B(n951), .Z(a_out[3]) );
  NAND U1118 ( .A(reg_source[3]), .B(n936), .Z(n951) );
  AND U1119 ( .A(n952), .B(n953), .Z(n950) );
  NANDN U1120 ( .A(n949), .B(imm_in[9]), .Z(n953) );
  NAND U1121 ( .A(c_pc[3]), .B(n935), .Z(n952) );
  NAND U1122 ( .A(n954), .B(n955), .Z(a_out[31]) );
  NAND U1123 ( .A(c_pc[31]), .B(n935), .Z(n955) );
  NAND U1124 ( .A(reg_source[31]), .B(n936), .Z(n954) );
  NAND U1125 ( .A(n956), .B(n957), .Z(a_out[30]) );
  NAND U1126 ( .A(c_pc[30]), .B(n935), .Z(n957) );
  NAND U1127 ( .A(reg_source[30]), .B(n936), .Z(n956) );
  NAND U1128 ( .A(n958), .B(n959), .Z(a_out[2]) );
  NAND U1129 ( .A(reg_source[2]), .B(n936), .Z(n959) );
  AND U1130 ( .A(n960), .B(n961), .Z(n958) );
  NANDN U1131 ( .A(n949), .B(imm_in[8]), .Z(n961) );
  NAND U1132 ( .A(c_pc[2]), .B(n935), .Z(n960) );
  NAND U1133 ( .A(n962), .B(n963), .Z(a_out[29]) );
  NAND U1134 ( .A(c_pc[29]), .B(n935), .Z(n963) );
  NAND U1135 ( .A(reg_source[29]), .B(n936), .Z(n962) );
  NAND U1136 ( .A(n964), .B(n965), .Z(a_out[28]) );
  NAND U1137 ( .A(c_pc[28]), .B(n935), .Z(n965) );
  NAND U1138 ( .A(reg_source[28]), .B(n936), .Z(n964) );
  NAND U1139 ( .A(n966), .B(n967), .Z(a_out[27]) );
  NAND U1140 ( .A(c_pc[27]), .B(n935), .Z(n967) );
  NAND U1141 ( .A(reg_source[27]), .B(n936), .Z(n966) );
  NAND U1142 ( .A(n968), .B(n969), .Z(a_out[26]) );
  NAND U1143 ( .A(c_pc[26]), .B(n935), .Z(n969) );
  NAND U1144 ( .A(reg_source[26]), .B(n936), .Z(n968) );
  NAND U1145 ( .A(n970), .B(n971), .Z(a_out[25]) );
  NAND U1146 ( .A(c_pc[25]), .B(n935), .Z(n971) );
  NAND U1147 ( .A(reg_source[25]), .B(n936), .Z(n970) );
  NAND U1148 ( .A(n972), .B(n973), .Z(a_out[24]) );
  NAND U1149 ( .A(c_pc[24]), .B(n935), .Z(n973) );
  NAND U1150 ( .A(reg_source[24]), .B(n936), .Z(n972) );
  NAND U1151 ( .A(n974), .B(n975), .Z(a_out[23]) );
  NAND U1152 ( .A(c_pc[23]), .B(n935), .Z(n975) );
  NAND U1153 ( .A(reg_source[23]), .B(n936), .Z(n974) );
  NAND U1154 ( .A(n976), .B(n977), .Z(a_out[22]) );
  NAND U1155 ( .A(c_pc[22]), .B(n935), .Z(n977) );
  NAND U1156 ( .A(reg_source[22]), .B(n936), .Z(n976) );
  NAND U1157 ( .A(n978), .B(n979), .Z(a_out[21]) );
  NAND U1158 ( .A(c_pc[21]), .B(n935), .Z(n979) );
  NAND U1159 ( .A(reg_source[21]), .B(n936), .Z(n978) );
  NAND U1160 ( .A(n980), .B(n981), .Z(a_out[20]) );
  NAND U1161 ( .A(c_pc[20]), .B(n935), .Z(n981) );
  NAND U1162 ( .A(reg_source[20]), .B(n936), .Z(n980) );
  NAND U1163 ( .A(n982), .B(n983), .Z(a_out[1]) );
  NANDN U1164 ( .A(n949), .B(imm_in[7]), .Z(n983) );
  NAND U1165 ( .A(reg_source[1]), .B(n936), .Z(n982) );
  NAND U1166 ( .A(n984), .B(n985), .Z(a_out[19]) );
  NAND U1167 ( .A(c_pc[19]), .B(n935), .Z(n985) );
  NAND U1168 ( .A(reg_source[19]), .B(n936), .Z(n984) );
  NAND U1169 ( .A(n986), .B(n987), .Z(a_out[18]) );
  NAND U1170 ( .A(c_pc[18]), .B(n935), .Z(n987) );
  NAND U1171 ( .A(reg_source[18]), .B(n936), .Z(n986) );
  NAND U1172 ( .A(n988), .B(n989), .Z(a_out[17]) );
  NAND U1173 ( .A(c_pc[17]), .B(n935), .Z(n989) );
  NAND U1174 ( .A(reg_source[17]), .B(n936), .Z(n988) );
  NAND U1175 ( .A(n990), .B(n991), .Z(a_out[16]) );
  NAND U1176 ( .A(c_pc[16]), .B(n935), .Z(n991) );
  NAND U1177 ( .A(reg_source[16]), .B(n936), .Z(n990) );
  NAND U1178 ( .A(n992), .B(n993), .Z(a_out[15]) );
  NAND U1179 ( .A(c_pc[15]), .B(n935), .Z(n993) );
  NAND U1180 ( .A(reg_source[15]), .B(n936), .Z(n992) );
  NAND U1181 ( .A(n994), .B(n995), .Z(a_out[14]) );
  NAND U1182 ( .A(c_pc[14]), .B(n935), .Z(n995) );
  NAND U1183 ( .A(reg_source[14]), .B(n936), .Z(n994) );
  NAND U1184 ( .A(n996), .B(n997), .Z(a_out[13]) );
  NAND U1185 ( .A(c_pc[13]), .B(n935), .Z(n997) );
  NAND U1186 ( .A(reg_source[13]), .B(n936), .Z(n996) );
  NAND U1187 ( .A(n998), .B(n999), .Z(a_out[12]) );
  NAND U1188 ( .A(c_pc[12]), .B(n935), .Z(n999) );
  NAND U1189 ( .A(reg_source[12]), .B(n936), .Z(n998) );
  NAND U1190 ( .A(n1000), .B(n1001), .Z(a_out[11]) );
  NAND U1191 ( .A(n935), .B(c_pc[11]), .Z(n1001) );
  NAND U1192 ( .A(reg_source[11]), .B(n936), .Z(n1000) );
  NAND U1193 ( .A(n1002), .B(n1003), .Z(a_out[10]) );
  NAND U1194 ( .A(n935), .B(c_pc[10]), .Z(n1003) );
  NOR U1195 ( .A(n1004), .B(a_mux[0]), .Z(n935) );
  IV U1196 ( .A(a_mux[1]), .Z(n1004) );
  NAND U1197 ( .A(n936), .B(reg_source[10]), .Z(n1002) );
  NAND U1198 ( .A(n1005), .B(n1006), .Z(a_out[0]) );
  NANDN U1199 ( .A(n949), .B(imm_in[6]), .Z(n1006) );
  NANDN U1200 ( .A(a_mux[1]), .B(a_mux[0]), .Z(n949) );
  NAND U1201 ( .A(n936), .B(reg_source[0]), .Z(n1005) );
  NOR U1202 ( .A(a_mux[1]), .B(a_mux[0]), .Z(n936) );
endmodule

