
module hamming_N160_CC4 ( clk, rst, x, y, o );
  input [39:0] x;
  input [39:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259;
  wire   [7:0] oglobal;

  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U43 ( .A(n93), .B(n92), .Z(n1) );
  NAND U44 ( .A(n90), .B(n91), .Z(n2) );
  NAND U45 ( .A(n1), .B(n2), .Z(n187) );
  NAND U46 ( .A(n223), .B(n224), .Z(n3) );
  XOR U47 ( .A(n223), .B(n224), .Z(n4) );
  NANDN U48 ( .A(n222), .B(n4), .Z(n5) );
  NAND U49 ( .A(n3), .B(n5), .Z(n242) );
  NANDN U50 ( .A(n221), .B(n220), .Z(n6) );
  NANDN U51 ( .A(n219), .B(oglobal[2]), .Z(n7) );
  NAND U52 ( .A(n6), .B(n7), .Z(n243) );
  NAND U53 ( .A(n150), .B(n152), .Z(n8) );
  XOR U54 ( .A(n150), .B(n152), .Z(n9) );
  NAND U55 ( .A(n9), .B(n151), .Z(n10) );
  NAND U56 ( .A(n8), .B(n10), .Z(n199) );
  XOR U57 ( .A(n227), .B(n225), .Z(n11) );
  NANDN U58 ( .A(n226), .B(n11), .Z(n12) );
  NAND U59 ( .A(n227), .B(n225), .Z(n13) );
  AND U60 ( .A(n12), .B(n13), .Z(n241) );
  NAND U61 ( .A(n126), .B(n125), .Z(n14) );
  NAND U62 ( .A(n123), .B(n124), .Z(n15) );
  NAND U63 ( .A(n14), .B(n15), .Z(n208) );
  NAND U64 ( .A(n71), .B(n70), .Z(n16) );
  NAND U65 ( .A(n68), .B(n69), .Z(n17) );
  NAND U66 ( .A(n16), .B(n17), .Z(n206) );
  NAND U67 ( .A(n89), .B(n88), .Z(n18) );
  NAND U68 ( .A(n86), .B(n87), .Z(n19) );
  AND U69 ( .A(n18), .B(n19), .Z(n186) );
  XOR U70 ( .A(n116), .B(n117), .Z(n20) );
  NANDN U71 ( .A(n118), .B(n20), .Z(n21) );
  NAND U72 ( .A(n116), .B(n117), .Z(n22) );
  AND U73 ( .A(n21), .B(n22), .Z(n165) );
  XOR U74 ( .A(n155), .B(n153), .Z(n23) );
  NANDN U75 ( .A(n154), .B(n23), .Z(n24) );
  NAND U76 ( .A(n155), .B(n153), .Z(n25) );
  AND U77 ( .A(n24), .B(n25), .Z(n202) );
  NAND U78 ( .A(n241), .B(n242), .Z(n26) );
  XOR U79 ( .A(n241), .B(n242), .Z(n27) );
  NANDN U80 ( .A(n240), .B(n27), .Z(n28) );
  NAND U81 ( .A(n26), .B(n28), .Z(n247) );
  NAND U82 ( .A(n122), .B(n121), .Z(n29) );
  NAND U83 ( .A(n119), .B(n120), .Z(n30) );
  NAND U84 ( .A(n29), .B(n30), .Z(n209) );
  NAND U85 ( .A(n97), .B(n96), .Z(n31) );
  NAND U86 ( .A(n94), .B(n95), .Z(n32) );
  NAND U87 ( .A(n31), .B(n32), .Z(n189) );
  NAND U88 ( .A(n131), .B(n130), .Z(n33) );
  NAND U89 ( .A(n128), .B(n129), .Z(n34) );
  NAND U90 ( .A(n33), .B(n34), .Z(n183) );
  XOR U91 ( .A(n205), .B(n206), .Z(n35) );
  NANDN U92 ( .A(n207), .B(n35), .Z(n36) );
  NAND U93 ( .A(n205), .B(n206), .Z(n37) );
  AND U94 ( .A(n36), .B(n37), .Z(n221) );
  NAND U95 ( .A(n156), .B(n158), .Z(n38) );
  XOR U96 ( .A(n156), .B(n158), .Z(n39) );
  NAND U97 ( .A(n39), .B(n157), .Z(n40) );
  NAND U98 ( .A(n38), .B(n40), .Z(n200) );
  NAND U99 ( .A(n160), .B(n162), .Z(n41) );
  XOR U100 ( .A(n160), .B(n162), .Z(n42) );
  NAND U101 ( .A(n42), .B(n161), .Z(n43) );
  NAND U102 ( .A(n41), .B(n43), .Z(n180) );
  NAND U103 ( .A(n237), .B(n239), .Z(n44) );
  XOR U104 ( .A(n237), .B(n239), .Z(n45) );
  NAND U105 ( .A(n45), .B(n238), .Z(n46) );
  NAND U106 ( .A(n44), .B(n46), .Z(n245) );
  XOR U107 ( .A(oglobal[1]), .B(n208), .Z(n47) );
  NAND U108 ( .A(n47), .B(n209), .Z(n48) );
  NAND U109 ( .A(oglobal[1]), .B(n208), .Z(n49) );
  AND U110 ( .A(n48), .B(n49), .Z(n219) );
  XOR U111 ( .A(n147), .B(n148), .Z(n50) );
  NANDN U112 ( .A(n149), .B(n50), .Z(n51) );
  NAND U113 ( .A(n147), .B(n148), .Z(n52) );
  AND U114 ( .A(n51), .B(n52), .Z(n171) );
  NAND U115 ( .A(n184), .B(n185), .Z(n53) );
  XOR U116 ( .A(n184), .B(n185), .Z(n54) );
  NANDN U117 ( .A(n183), .B(n54), .Z(n55) );
  NAND U118 ( .A(n53), .B(n55), .Z(n226) );
  NAND U119 ( .A(n177), .B(n178), .Z(n56) );
  XOR U120 ( .A(n177), .B(n178), .Z(n57) );
  NANDN U121 ( .A(n176), .B(n57), .Z(n58) );
  NAND U122 ( .A(n56), .B(n58), .Z(n231) );
  XOR U123 ( .A(n180), .B(n181), .Z(n59) );
  NANDN U124 ( .A(n182), .B(n59), .Z(n60) );
  NAND U125 ( .A(n180), .B(n181), .Z(n61) );
  AND U126 ( .A(n60), .B(n61), .Z(n214) );
  NAND U127 ( .A(n252), .B(n253), .Z(n257) );
  XOR U128 ( .A(x[27]), .B(y[27]), .Z(n126) );
  XOR U129 ( .A(x[39]), .B(y[39]), .Z(n124) );
  XOR U130 ( .A(x[25]), .B(y[25]), .Z(n123) );
  XOR U131 ( .A(n124), .B(n123), .Z(n125) );
  XOR U132 ( .A(n126), .B(n125), .Z(n136) );
  XOR U133 ( .A(x[35]), .B(y[35]), .Z(n133) );
  XOR U134 ( .A(x[33]), .B(y[33]), .Z(n132) );
  XOR U135 ( .A(n133), .B(n132), .Z(n135) );
  XOR U136 ( .A(n136), .B(n135), .Z(n155) );
  XOR U137 ( .A(x[3]), .B(y[3]), .Z(n95) );
  XOR U138 ( .A(x[1]), .B(y[1]), .Z(n94) );
  XOR U139 ( .A(n95), .B(n94), .Z(n97) );
  XOR U140 ( .A(x[5]), .B(y[5]), .Z(n96) );
  XNOR U141 ( .A(n97), .B(n96), .Z(n154) );
  XOR U142 ( .A(x[17]), .B(y[17]), .Z(n143) );
  XOR U143 ( .A(x[13]), .B(y[13]), .Z(n140) );
  XOR U144 ( .A(x[15]), .B(y[15]), .Z(n139) );
  XOR U145 ( .A(n140), .B(n139), .Z(n142) );
  XOR U146 ( .A(n143), .B(n142), .Z(n153) );
  XOR U147 ( .A(n154), .B(n153), .Z(n62) );
  XNOR U148 ( .A(n155), .B(n62), .Z(n162) );
  XOR U149 ( .A(x[24]), .B(y[24]), .Z(n106) );
  XOR U150 ( .A(x[28]), .B(y[28]), .Z(n104) );
  XNOR U151 ( .A(x[26]), .B(y[26]), .Z(n105) );
  XOR U152 ( .A(n104), .B(n105), .Z(n107) );
  XOR U153 ( .A(n106), .B(n107), .Z(n148) );
  XOR U154 ( .A(x[30]), .B(y[30]), .Z(n111) );
  XNOR U155 ( .A(x[32]), .B(y[32]), .Z(n110) );
  XOR U156 ( .A(oglobal[0]), .B(n110), .Z(n112) );
  XNOR U157 ( .A(n111), .B(n112), .Z(n149) );
  XOR U158 ( .A(x[18]), .B(y[18]), .Z(n100) );
  XOR U159 ( .A(x[22]), .B(y[22]), .Z(n98) );
  XNOR U160 ( .A(x[20]), .B(y[20]), .Z(n99) );
  XOR U161 ( .A(n98), .B(n99), .Z(n101) );
  XOR U162 ( .A(n100), .B(n101), .Z(n147) );
  XOR U163 ( .A(n149), .B(n147), .Z(n63) );
  XOR U164 ( .A(n148), .B(n63), .Z(n161) );
  XOR U165 ( .A(x[6]), .B(y[6]), .Z(n71) );
  XOR U166 ( .A(x[8]), .B(y[8]), .Z(n69) );
  XOR U167 ( .A(x[10]), .B(y[10]), .Z(n68) );
  XOR U168 ( .A(n69), .B(n68), .Z(n70) );
  XOR U169 ( .A(n71), .B(n70), .Z(n158) );
  XOR U170 ( .A(x[4]), .B(y[4]), .Z(n91) );
  XOR U171 ( .A(x[2]), .B(y[2]), .Z(n90) );
  XOR U172 ( .A(n91), .B(n90), .Z(n93) );
  XOR U173 ( .A(x[0]), .B(y[0]), .Z(n92) );
  XOR U174 ( .A(n93), .B(n92), .Z(n157) );
  XOR U175 ( .A(x[12]), .B(y[12]), .Z(n75) );
  XOR U176 ( .A(x[14]), .B(y[14]), .Z(n73) );
  XOR U177 ( .A(x[16]), .B(y[16]), .Z(n72) );
  XOR U178 ( .A(n73), .B(n72), .Z(n74) );
  XOR U179 ( .A(n75), .B(n74), .Z(n156) );
  XNOR U180 ( .A(n157), .B(n156), .Z(n64) );
  XOR U181 ( .A(n158), .B(n64), .Z(n117) );
  XOR U182 ( .A(x[23]), .B(y[23]), .Z(n122) );
  XOR U183 ( .A(x[19]), .B(y[19]), .Z(n120) );
  XOR U184 ( .A(x[21]), .B(y[21]), .Z(n119) );
  XOR U185 ( .A(n120), .B(n119), .Z(n121) );
  XOR U186 ( .A(n122), .B(n121), .Z(n152) );
  XOR U187 ( .A(x[9]), .B(y[9]), .Z(n87) );
  XOR U188 ( .A(x[7]), .B(y[7]), .Z(n86) );
  XOR U189 ( .A(n87), .B(n86), .Z(n89) );
  XOR U190 ( .A(x[11]), .B(y[11]), .Z(n88) );
  XOR U191 ( .A(n89), .B(n88), .Z(n151) );
  XOR U192 ( .A(x[31]), .B(y[31]), .Z(n131) );
  XOR U193 ( .A(x[29]), .B(y[29]), .Z(n129) );
  XOR U194 ( .A(x[37]), .B(y[37]), .Z(n128) );
  XOR U195 ( .A(n129), .B(n128), .Z(n130) );
  XOR U196 ( .A(n131), .B(n130), .Z(n150) );
  XNOR U197 ( .A(n151), .B(n150), .Z(n65) );
  XNOR U198 ( .A(n152), .B(n65), .Z(n118) );
  XOR U199 ( .A(x[34]), .B(y[34]), .Z(n81) );
  XOR U200 ( .A(x[38]), .B(y[38]), .Z(n79) );
  XNOR U201 ( .A(x[36]), .B(y[36]), .Z(n80) );
  XOR U202 ( .A(n79), .B(n80), .Z(n82) );
  XOR U203 ( .A(n81), .B(n82), .Z(n116) );
  XOR U204 ( .A(n118), .B(n116), .Z(n66) );
  XOR U205 ( .A(n117), .B(n66), .Z(n160) );
  XNOR U206 ( .A(n161), .B(n160), .Z(n67) );
  XNOR U207 ( .A(n162), .B(n67), .Z(o[0]) );
  NAND U208 ( .A(n73), .B(n72), .Z(n78) );
  IV U209 ( .A(n74), .Z(n76) );
  NANDN U210 ( .A(n76), .B(n75), .Z(n77) );
  AND U211 ( .A(n78), .B(n77), .Z(n207) );
  NANDN U212 ( .A(n80), .B(n79), .Z(n84) );
  NANDN U213 ( .A(n82), .B(n81), .Z(n83) );
  NAND U214 ( .A(n84), .B(n83), .Z(n205) );
  XOR U215 ( .A(n207), .B(n205), .Z(n85) );
  XOR U216 ( .A(n206), .B(n85), .Z(n177) );
  XNOR U217 ( .A(n186), .B(n187), .Z(n188) );
  XNOR U218 ( .A(n188), .B(n189), .Z(n178) );
  NANDN U219 ( .A(n99), .B(n98), .Z(n103) );
  NANDN U220 ( .A(n101), .B(n100), .Z(n102) );
  AND U221 ( .A(n103), .B(n102), .Z(n192) );
  NANDN U222 ( .A(n105), .B(n104), .Z(n109) );
  NANDN U223 ( .A(n107), .B(n106), .Z(n108) );
  NAND U224 ( .A(n109), .B(n108), .Z(n193) );
  XNOR U225 ( .A(n192), .B(n193), .Z(n194) );
  NANDN U226 ( .A(n110), .B(oglobal[0]), .Z(n114) );
  NANDN U227 ( .A(n112), .B(n111), .Z(n113) );
  NAND U228 ( .A(n114), .B(n113), .Z(n195) );
  XOR U229 ( .A(n194), .B(n195), .Z(n176) );
  XOR U230 ( .A(n178), .B(n176), .Z(n115) );
  XNOR U231 ( .A(n177), .B(n115), .Z(n164) );
  XNOR U232 ( .A(n164), .B(n165), .Z(n166) );
  XOR U233 ( .A(n208), .B(oglobal[1]), .Z(n127) );
  XOR U234 ( .A(n209), .B(n127), .Z(n173) );
  IV U235 ( .A(n132), .Z(n134) );
  NANDN U236 ( .A(n134), .B(n133), .Z(n138) );
  NAND U237 ( .A(n136), .B(n135), .Z(n137) );
  AND U238 ( .A(n138), .B(n137), .Z(n185) );
  IV U239 ( .A(n139), .Z(n141) );
  NANDN U240 ( .A(n141), .B(n140), .Z(n145) );
  NAND U241 ( .A(n143), .B(n142), .Z(n144) );
  AND U242 ( .A(n145), .B(n144), .Z(n184) );
  XNOR U243 ( .A(n185), .B(n184), .Z(n146) );
  XOR U244 ( .A(n183), .B(n146), .Z(n170) );
  XNOR U245 ( .A(n170), .B(n171), .Z(n172) );
  XOR U246 ( .A(n173), .B(n172), .Z(n167) );
  XOR U247 ( .A(n166), .B(n167), .Z(n181) );
  XNOR U248 ( .A(n202), .B(n200), .Z(n159) );
  XNOR U249 ( .A(n199), .B(n159), .Z(n182) );
  XNOR U250 ( .A(n182), .B(n180), .Z(n163) );
  XOR U251 ( .A(n181), .B(n163), .Z(o[1]) );
  NANDN U252 ( .A(n165), .B(n164), .Z(n169) );
  NANDN U253 ( .A(n167), .B(n166), .Z(n168) );
  AND U254 ( .A(n169), .B(n168), .Z(n232) );
  NANDN U255 ( .A(n171), .B(n170), .Z(n175) );
  NANDN U256 ( .A(n173), .B(n172), .Z(n174) );
  AND U257 ( .A(n175), .B(n174), .Z(n230) );
  IV U258 ( .A(n230), .Z(n229) );
  XOR U259 ( .A(n229), .B(n231), .Z(n179) );
  XNOR U260 ( .A(n232), .B(n179), .Z(n215) );
  NANDN U261 ( .A(n187), .B(n186), .Z(n191) );
  NANDN U262 ( .A(n189), .B(n188), .Z(n190) );
  AND U263 ( .A(n191), .B(n190), .Z(n227) );
  NANDN U264 ( .A(n193), .B(n192), .Z(n197) );
  NANDN U265 ( .A(n195), .B(n194), .Z(n196) );
  AND U266 ( .A(n197), .B(n196), .Z(n225) );
  XNOR U267 ( .A(n227), .B(n225), .Z(n198) );
  XOR U268 ( .A(n226), .B(n198), .Z(n222) );
  NAND U269 ( .A(n200), .B(n199), .Z(n204) );
  NOR U270 ( .A(n200), .B(n199), .Z(n201) );
  OR U271 ( .A(n202), .B(n201), .Z(n203) );
  AND U272 ( .A(n204), .B(n203), .Z(n224) );
  XNOR U273 ( .A(n219), .B(oglobal[2]), .Z(n220) );
  XOR U274 ( .A(n221), .B(n220), .Z(n223) );
  XOR U275 ( .A(n224), .B(n223), .Z(n210) );
  XOR U276 ( .A(n222), .B(n210), .Z(n213) );
  IV U277 ( .A(n213), .Z(n212) );
  XOR U278 ( .A(n214), .B(n212), .Z(n211) );
  XNOR U279 ( .A(n215), .B(n211), .Z(o[2]) );
  OR U280 ( .A(n214), .B(n212), .Z(n218) );
  ANDN U281 ( .B(n214), .A(n213), .Z(n216) );
  OR U282 ( .A(n216), .B(n215), .Z(n217) );
  AND U283 ( .A(n218), .B(n217), .Z(n237) );
  XOR U284 ( .A(oglobal[3]), .B(n243), .Z(n240) );
  XNOR U285 ( .A(n242), .B(n241), .Z(n228) );
  XOR U286 ( .A(n240), .B(n228), .Z(n239) );
  OR U287 ( .A(n231), .B(n229), .Z(n235) );
  ANDN U288 ( .B(n231), .A(n230), .Z(n233) );
  NANDN U289 ( .A(n233), .B(n232), .Z(n234) );
  AND U290 ( .A(n235), .B(n234), .Z(n238) );
  XOR U291 ( .A(n239), .B(n238), .Z(n236) );
  XNOR U292 ( .A(n237), .B(n236), .Z(o[3]) );
  AND U293 ( .A(oglobal[3]), .B(n243), .Z(n250) );
  XOR U294 ( .A(n250), .B(oglobal[4]), .Z(n246) );
  XNOR U295 ( .A(n247), .B(n246), .Z(n244) );
  XNOR U296 ( .A(n245), .B(n244), .Z(o[4]) );
  NANDN U297 ( .A(n245), .B(n246), .Z(n249) );
  NANDN U298 ( .A(n246), .B(n245), .Z(n248) );
  ANDN U299 ( .B(n248), .A(n247), .Z(n253) );
  ANDN U300 ( .B(n249), .A(n253), .Z(n251) );
  AND U301 ( .A(n250), .B(oglobal[4]), .Z(n252) );
  ANDN U302 ( .B(n251), .A(n252), .Z(n255) );
  NANDN U303 ( .A(n255), .B(n257), .Z(n254) );
  XNOR U304 ( .A(oglobal[5]), .B(n254), .Z(o[5]) );
  NANDN U305 ( .A(n255), .B(oglobal[5]), .Z(n256) );
  AND U306 ( .A(n257), .B(n256), .Z(n258) );
  XNOR U307 ( .A(n258), .B(oglobal[6]), .Z(o[6]) );
  NANDN U308 ( .A(n258), .B(oglobal[6]), .Z(n259) );
  XNOR U309 ( .A(oglobal[7]), .B(n259), .Z(o[7]) );
endmodule

