
module mult_N1024_CC256 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [3:0] b;
  output [2047:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720;
  wire   [2047:0] sreg;

  DFF \sreg_reg[2043]  ( .D(c[2047]), .CLK(clk), .RST(rst), .Q(sreg[2043]) );
  DFF \sreg_reg[2042]  ( .D(c[2046]), .CLK(clk), .RST(rst), .Q(sreg[2042]) );
  DFF \sreg_reg[2041]  ( .D(c[2045]), .CLK(clk), .RST(rst), .Q(sreg[2041]) );
  DFF \sreg_reg[2040]  ( .D(c[2044]), .CLK(clk), .RST(rst), .Q(sreg[2040]) );
  DFF \sreg_reg[2039]  ( .D(c[2043]), .CLK(clk), .RST(rst), .Q(sreg[2039]) );
  DFF \sreg_reg[2038]  ( .D(c[2042]), .CLK(clk), .RST(rst), .Q(sreg[2038]) );
  DFF \sreg_reg[2037]  ( .D(c[2041]), .CLK(clk), .RST(rst), .Q(sreg[2037]) );
  DFF \sreg_reg[2036]  ( .D(c[2040]), .CLK(clk), .RST(rst), .Q(sreg[2036]) );
  DFF \sreg_reg[2035]  ( .D(c[2039]), .CLK(clk), .RST(rst), .Q(sreg[2035]) );
  DFF \sreg_reg[2034]  ( .D(c[2038]), .CLK(clk), .RST(rst), .Q(sreg[2034]) );
  DFF \sreg_reg[2033]  ( .D(c[2037]), .CLK(clk), .RST(rst), .Q(sreg[2033]) );
  DFF \sreg_reg[2032]  ( .D(c[2036]), .CLK(clk), .RST(rst), .Q(sreg[2032]) );
  DFF \sreg_reg[2031]  ( .D(c[2035]), .CLK(clk), .RST(rst), .Q(sreg[2031]) );
  DFF \sreg_reg[2030]  ( .D(c[2034]), .CLK(clk), .RST(rst), .Q(sreg[2030]) );
  DFF \sreg_reg[2029]  ( .D(c[2033]), .CLK(clk), .RST(rst), .Q(sreg[2029]) );
  DFF \sreg_reg[2028]  ( .D(c[2032]), .CLK(clk), .RST(rst), .Q(sreg[2028]) );
  DFF \sreg_reg[2027]  ( .D(c[2031]), .CLK(clk), .RST(rst), .Q(sreg[2027]) );
  DFF \sreg_reg[2026]  ( .D(c[2030]), .CLK(clk), .RST(rst), .Q(sreg[2026]) );
  DFF \sreg_reg[2025]  ( .D(c[2029]), .CLK(clk), .RST(rst), .Q(sreg[2025]) );
  DFF \sreg_reg[2024]  ( .D(c[2028]), .CLK(clk), .RST(rst), .Q(sreg[2024]) );
  DFF \sreg_reg[2023]  ( .D(c[2027]), .CLK(clk), .RST(rst), .Q(sreg[2023]) );
  DFF \sreg_reg[2022]  ( .D(c[2026]), .CLK(clk), .RST(rst), .Q(sreg[2022]) );
  DFF \sreg_reg[2021]  ( .D(c[2025]), .CLK(clk), .RST(rst), .Q(sreg[2021]) );
  DFF \sreg_reg[2020]  ( .D(c[2024]), .CLK(clk), .RST(rst), .Q(sreg[2020]) );
  DFF \sreg_reg[2019]  ( .D(c[2023]), .CLK(clk), .RST(rst), .Q(sreg[2019]) );
  DFF \sreg_reg[2018]  ( .D(c[2022]), .CLK(clk), .RST(rst), .Q(sreg[2018]) );
  DFF \sreg_reg[2017]  ( .D(c[2021]), .CLK(clk), .RST(rst), .Q(sreg[2017]) );
  DFF \sreg_reg[2016]  ( .D(c[2020]), .CLK(clk), .RST(rst), .Q(sreg[2016]) );
  DFF \sreg_reg[2015]  ( .D(c[2019]), .CLK(clk), .RST(rst), .Q(sreg[2015]) );
  DFF \sreg_reg[2014]  ( .D(c[2018]), .CLK(clk), .RST(rst), .Q(sreg[2014]) );
  DFF \sreg_reg[2013]  ( .D(c[2017]), .CLK(clk), .RST(rst), .Q(sreg[2013]) );
  DFF \sreg_reg[2012]  ( .D(c[2016]), .CLK(clk), .RST(rst), .Q(sreg[2012]) );
  DFF \sreg_reg[2011]  ( .D(c[2015]), .CLK(clk), .RST(rst), .Q(sreg[2011]) );
  DFF \sreg_reg[2010]  ( .D(c[2014]), .CLK(clk), .RST(rst), .Q(sreg[2010]) );
  DFF \sreg_reg[2009]  ( .D(c[2013]), .CLK(clk), .RST(rst), .Q(sreg[2009]) );
  DFF \sreg_reg[2008]  ( .D(c[2012]), .CLK(clk), .RST(rst), .Q(sreg[2008]) );
  DFF \sreg_reg[2007]  ( .D(c[2011]), .CLK(clk), .RST(rst), .Q(sreg[2007]) );
  DFF \sreg_reg[2006]  ( .D(c[2010]), .CLK(clk), .RST(rst), .Q(sreg[2006]) );
  DFF \sreg_reg[2005]  ( .D(c[2009]), .CLK(clk), .RST(rst), .Q(sreg[2005]) );
  DFF \sreg_reg[2004]  ( .D(c[2008]), .CLK(clk), .RST(rst), .Q(sreg[2004]) );
  DFF \sreg_reg[2003]  ( .D(c[2007]), .CLK(clk), .RST(rst), .Q(sreg[2003]) );
  DFF \sreg_reg[2002]  ( .D(c[2006]), .CLK(clk), .RST(rst), .Q(sreg[2002]) );
  DFF \sreg_reg[2001]  ( .D(c[2005]), .CLK(clk), .RST(rst), .Q(sreg[2001]) );
  DFF \sreg_reg[2000]  ( .D(c[2004]), .CLK(clk), .RST(rst), .Q(sreg[2000]) );
  DFF \sreg_reg[1999]  ( .D(c[2003]), .CLK(clk), .RST(rst), .Q(sreg[1999]) );
  DFF \sreg_reg[1998]  ( .D(c[2002]), .CLK(clk), .RST(rst), .Q(sreg[1998]) );
  DFF \sreg_reg[1997]  ( .D(c[2001]), .CLK(clk), .RST(rst), .Q(sreg[1997]) );
  DFF \sreg_reg[1996]  ( .D(c[2000]), .CLK(clk), .RST(rst), .Q(sreg[1996]) );
  DFF \sreg_reg[1995]  ( .D(c[1999]), .CLK(clk), .RST(rst), .Q(sreg[1995]) );
  DFF \sreg_reg[1994]  ( .D(c[1998]), .CLK(clk), .RST(rst), .Q(sreg[1994]) );
  DFF \sreg_reg[1993]  ( .D(c[1997]), .CLK(clk), .RST(rst), .Q(sreg[1993]) );
  DFF \sreg_reg[1992]  ( .D(c[1996]), .CLK(clk), .RST(rst), .Q(sreg[1992]) );
  DFF \sreg_reg[1991]  ( .D(c[1995]), .CLK(clk), .RST(rst), .Q(sreg[1991]) );
  DFF \sreg_reg[1990]  ( .D(c[1994]), .CLK(clk), .RST(rst), .Q(sreg[1990]) );
  DFF \sreg_reg[1989]  ( .D(c[1993]), .CLK(clk), .RST(rst), .Q(sreg[1989]) );
  DFF \sreg_reg[1988]  ( .D(c[1992]), .CLK(clk), .RST(rst), .Q(sreg[1988]) );
  DFF \sreg_reg[1987]  ( .D(c[1991]), .CLK(clk), .RST(rst), .Q(sreg[1987]) );
  DFF \sreg_reg[1986]  ( .D(c[1990]), .CLK(clk), .RST(rst), .Q(sreg[1986]) );
  DFF \sreg_reg[1985]  ( .D(c[1989]), .CLK(clk), .RST(rst), .Q(sreg[1985]) );
  DFF \sreg_reg[1984]  ( .D(c[1988]), .CLK(clk), .RST(rst), .Q(sreg[1984]) );
  DFF \sreg_reg[1983]  ( .D(c[1987]), .CLK(clk), .RST(rst), .Q(sreg[1983]) );
  DFF \sreg_reg[1982]  ( .D(c[1986]), .CLK(clk), .RST(rst), .Q(sreg[1982]) );
  DFF \sreg_reg[1981]  ( .D(c[1985]), .CLK(clk), .RST(rst), .Q(sreg[1981]) );
  DFF \sreg_reg[1980]  ( .D(c[1984]), .CLK(clk), .RST(rst), .Q(sreg[1980]) );
  DFF \sreg_reg[1979]  ( .D(c[1983]), .CLK(clk), .RST(rst), .Q(sreg[1979]) );
  DFF \sreg_reg[1978]  ( .D(c[1982]), .CLK(clk), .RST(rst), .Q(sreg[1978]) );
  DFF \sreg_reg[1977]  ( .D(c[1981]), .CLK(clk), .RST(rst), .Q(sreg[1977]) );
  DFF \sreg_reg[1976]  ( .D(c[1980]), .CLK(clk), .RST(rst), .Q(sreg[1976]) );
  DFF \sreg_reg[1975]  ( .D(c[1979]), .CLK(clk), .RST(rst), .Q(sreg[1975]) );
  DFF \sreg_reg[1974]  ( .D(c[1978]), .CLK(clk), .RST(rst), .Q(sreg[1974]) );
  DFF \sreg_reg[1973]  ( .D(c[1977]), .CLK(clk), .RST(rst), .Q(sreg[1973]) );
  DFF \sreg_reg[1972]  ( .D(c[1976]), .CLK(clk), .RST(rst), .Q(sreg[1972]) );
  DFF \sreg_reg[1971]  ( .D(c[1975]), .CLK(clk), .RST(rst), .Q(sreg[1971]) );
  DFF \sreg_reg[1970]  ( .D(c[1974]), .CLK(clk), .RST(rst), .Q(sreg[1970]) );
  DFF \sreg_reg[1969]  ( .D(c[1973]), .CLK(clk), .RST(rst), .Q(sreg[1969]) );
  DFF \sreg_reg[1968]  ( .D(c[1972]), .CLK(clk), .RST(rst), .Q(sreg[1968]) );
  DFF \sreg_reg[1967]  ( .D(c[1971]), .CLK(clk), .RST(rst), .Q(sreg[1967]) );
  DFF \sreg_reg[1966]  ( .D(c[1970]), .CLK(clk), .RST(rst), .Q(sreg[1966]) );
  DFF \sreg_reg[1965]  ( .D(c[1969]), .CLK(clk), .RST(rst), .Q(sreg[1965]) );
  DFF \sreg_reg[1964]  ( .D(c[1968]), .CLK(clk), .RST(rst), .Q(sreg[1964]) );
  DFF \sreg_reg[1963]  ( .D(c[1967]), .CLK(clk), .RST(rst), .Q(sreg[1963]) );
  DFF \sreg_reg[1962]  ( .D(c[1966]), .CLK(clk), .RST(rst), .Q(sreg[1962]) );
  DFF \sreg_reg[1961]  ( .D(c[1965]), .CLK(clk), .RST(rst), .Q(sreg[1961]) );
  DFF \sreg_reg[1960]  ( .D(c[1964]), .CLK(clk), .RST(rst), .Q(sreg[1960]) );
  DFF \sreg_reg[1959]  ( .D(c[1963]), .CLK(clk), .RST(rst), .Q(sreg[1959]) );
  DFF \sreg_reg[1958]  ( .D(c[1962]), .CLK(clk), .RST(rst), .Q(sreg[1958]) );
  DFF \sreg_reg[1957]  ( .D(c[1961]), .CLK(clk), .RST(rst), .Q(sreg[1957]) );
  DFF \sreg_reg[1956]  ( .D(c[1960]), .CLK(clk), .RST(rst), .Q(sreg[1956]) );
  DFF \sreg_reg[1955]  ( .D(c[1959]), .CLK(clk), .RST(rst), .Q(sreg[1955]) );
  DFF \sreg_reg[1954]  ( .D(c[1958]), .CLK(clk), .RST(rst), .Q(sreg[1954]) );
  DFF \sreg_reg[1953]  ( .D(c[1957]), .CLK(clk), .RST(rst), .Q(sreg[1953]) );
  DFF \sreg_reg[1952]  ( .D(c[1956]), .CLK(clk), .RST(rst), .Q(sreg[1952]) );
  DFF \sreg_reg[1951]  ( .D(c[1955]), .CLK(clk), .RST(rst), .Q(sreg[1951]) );
  DFF \sreg_reg[1950]  ( .D(c[1954]), .CLK(clk), .RST(rst), .Q(sreg[1950]) );
  DFF \sreg_reg[1949]  ( .D(c[1953]), .CLK(clk), .RST(rst), .Q(sreg[1949]) );
  DFF \sreg_reg[1948]  ( .D(c[1952]), .CLK(clk), .RST(rst), .Q(sreg[1948]) );
  DFF \sreg_reg[1947]  ( .D(c[1951]), .CLK(clk), .RST(rst), .Q(sreg[1947]) );
  DFF \sreg_reg[1946]  ( .D(c[1950]), .CLK(clk), .RST(rst), .Q(sreg[1946]) );
  DFF \sreg_reg[1945]  ( .D(c[1949]), .CLK(clk), .RST(rst), .Q(sreg[1945]) );
  DFF \sreg_reg[1944]  ( .D(c[1948]), .CLK(clk), .RST(rst), .Q(sreg[1944]) );
  DFF \sreg_reg[1943]  ( .D(c[1947]), .CLK(clk), .RST(rst), .Q(sreg[1943]) );
  DFF \sreg_reg[1942]  ( .D(c[1946]), .CLK(clk), .RST(rst), .Q(sreg[1942]) );
  DFF \sreg_reg[1941]  ( .D(c[1945]), .CLK(clk), .RST(rst), .Q(sreg[1941]) );
  DFF \sreg_reg[1940]  ( .D(c[1944]), .CLK(clk), .RST(rst), .Q(sreg[1940]) );
  DFF \sreg_reg[1939]  ( .D(c[1943]), .CLK(clk), .RST(rst), .Q(sreg[1939]) );
  DFF \sreg_reg[1938]  ( .D(c[1942]), .CLK(clk), .RST(rst), .Q(sreg[1938]) );
  DFF \sreg_reg[1937]  ( .D(c[1941]), .CLK(clk), .RST(rst), .Q(sreg[1937]) );
  DFF \sreg_reg[1936]  ( .D(c[1940]), .CLK(clk), .RST(rst), .Q(sreg[1936]) );
  DFF \sreg_reg[1935]  ( .D(c[1939]), .CLK(clk), .RST(rst), .Q(sreg[1935]) );
  DFF \sreg_reg[1934]  ( .D(c[1938]), .CLK(clk), .RST(rst), .Q(sreg[1934]) );
  DFF \sreg_reg[1933]  ( .D(c[1937]), .CLK(clk), .RST(rst), .Q(sreg[1933]) );
  DFF \sreg_reg[1932]  ( .D(c[1936]), .CLK(clk), .RST(rst), .Q(sreg[1932]) );
  DFF \sreg_reg[1931]  ( .D(c[1935]), .CLK(clk), .RST(rst), .Q(sreg[1931]) );
  DFF \sreg_reg[1930]  ( .D(c[1934]), .CLK(clk), .RST(rst), .Q(sreg[1930]) );
  DFF \sreg_reg[1929]  ( .D(c[1933]), .CLK(clk), .RST(rst), .Q(sreg[1929]) );
  DFF \sreg_reg[1928]  ( .D(c[1932]), .CLK(clk), .RST(rst), .Q(sreg[1928]) );
  DFF \sreg_reg[1927]  ( .D(c[1931]), .CLK(clk), .RST(rst), .Q(sreg[1927]) );
  DFF \sreg_reg[1926]  ( .D(c[1930]), .CLK(clk), .RST(rst), .Q(sreg[1926]) );
  DFF \sreg_reg[1925]  ( .D(c[1929]), .CLK(clk), .RST(rst), .Q(sreg[1925]) );
  DFF \sreg_reg[1924]  ( .D(c[1928]), .CLK(clk), .RST(rst), .Q(sreg[1924]) );
  DFF \sreg_reg[1923]  ( .D(c[1927]), .CLK(clk), .RST(rst), .Q(sreg[1923]) );
  DFF \sreg_reg[1922]  ( .D(c[1926]), .CLK(clk), .RST(rst), .Q(sreg[1922]) );
  DFF \sreg_reg[1921]  ( .D(c[1925]), .CLK(clk), .RST(rst), .Q(sreg[1921]) );
  DFF \sreg_reg[1920]  ( .D(c[1924]), .CLK(clk), .RST(rst), .Q(sreg[1920]) );
  DFF \sreg_reg[1919]  ( .D(c[1923]), .CLK(clk), .RST(rst), .Q(sreg[1919]) );
  DFF \sreg_reg[1918]  ( .D(c[1922]), .CLK(clk), .RST(rst), .Q(sreg[1918]) );
  DFF \sreg_reg[1917]  ( .D(c[1921]), .CLK(clk), .RST(rst), .Q(sreg[1917]) );
  DFF \sreg_reg[1916]  ( .D(c[1920]), .CLK(clk), .RST(rst), .Q(sreg[1916]) );
  DFF \sreg_reg[1915]  ( .D(c[1919]), .CLK(clk), .RST(rst), .Q(sreg[1915]) );
  DFF \sreg_reg[1914]  ( .D(c[1918]), .CLK(clk), .RST(rst), .Q(sreg[1914]) );
  DFF \sreg_reg[1913]  ( .D(c[1917]), .CLK(clk), .RST(rst), .Q(sreg[1913]) );
  DFF \sreg_reg[1912]  ( .D(c[1916]), .CLK(clk), .RST(rst), .Q(sreg[1912]) );
  DFF \sreg_reg[1911]  ( .D(c[1915]), .CLK(clk), .RST(rst), .Q(sreg[1911]) );
  DFF \sreg_reg[1910]  ( .D(c[1914]), .CLK(clk), .RST(rst), .Q(sreg[1910]) );
  DFF \sreg_reg[1909]  ( .D(c[1913]), .CLK(clk), .RST(rst), .Q(sreg[1909]) );
  DFF \sreg_reg[1908]  ( .D(c[1912]), .CLK(clk), .RST(rst), .Q(sreg[1908]) );
  DFF \sreg_reg[1907]  ( .D(c[1911]), .CLK(clk), .RST(rst), .Q(sreg[1907]) );
  DFF \sreg_reg[1906]  ( .D(c[1910]), .CLK(clk), .RST(rst), .Q(sreg[1906]) );
  DFF \sreg_reg[1905]  ( .D(c[1909]), .CLK(clk), .RST(rst), .Q(sreg[1905]) );
  DFF \sreg_reg[1904]  ( .D(c[1908]), .CLK(clk), .RST(rst), .Q(sreg[1904]) );
  DFF \sreg_reg[1903]  ( .D(c[1907]), .CLK(clk), .RST(rst), .Q(sreg[1903]) );
  DFF \sreg_reg[1902]  ( .D(c[1906]), .CLK(clk), .RST(rst), .Q(sreg[1902]) );
  DFF \sreg_reg[1901]  ( .D(c[1905]), .CLK(clk), .RST(rst), .Q(sreg[1901]) );
  DFF \sreg_reg[1900]  ( .D(c[1904]), .CLK(clk), .RST(rst), .Q(sreg[1900]) );
  DFF \sreg_reg[1899]  ( .D(c[1903]), .CLK(clk), .RST(rst), .Q(sreg[1899]) );
  DFF \sreg_reg[1898]  ( .D(c[1902]), .CLK(clk), .RST(rst), .Q(sreg[1898]) );
  DFF \sreg_reg[1897]  ( .D(c[1901]), .CLK(clk), .RST(rst), .Q(sreg[1897]) );
  DFF \sreg_reg[1896]  ( .D(c[1900]), .CLK(clk), .RST(rst), .Q(sreg[1896]) );
  DFF \sreg_reg[1895]  ( .D(c[1899]), .CLK(clk), .RST(rst), .Q(sreg[1895]) );
  DFF \sreg_reg[1894]  ( .D(c[1898]), .CLK(clk), .RST(rst), .Q(sreg[1894]) );
  DFF \sreg_reg[1893]  ( .D(c[1897]), .CLK(clk), .RST(rst), .Q(sreg[1893]) );
  DFF \sreg_reg[1892]  ( .D(c[1896]), .CLK(clk), .RST(rst), .Q(sreg[1892]) );
  DFF \sreg_reg[1891]  ( .D(c[1895]), .CLK(clk), .RST(rst), .Q(sreg[1891]) );
  DFF \sreg_reg[1890]  ( .D(c[1894]), .CLK(clk), .RST(rst), .Q(sreg[1890]) );
  DFF \sreg_reg[1889]  ( .D(c[1893]), .CLK(clk), .RST(rst), .Q(sreg[1889]) );
  DFF \sreg_reg[1888]  ( .D(c[1892]), .CLK(clk), .RST(rst), .Q(sreg[1888]) );
  DFF \sreg_reg[1887]  ( .D(c[1891]), .CLK(clk), .RST(rst), .Q(sreg[1887]) );
  DFF \sreg_reg[1886]  ( .D(c[1890]), .CLK(clk), .RST(rst), .Q(sreg[1886]) );
  DFF \sreg_reg[1885]  ( .D(c[1889]), .CLK(clk), .RST(rst), .Q(sreg[1885]) );
  DFF \sreg_reg[1884]  ( .D(c[1888]), .CLK(clk), .RST(rst), .Q(sreg[1884]) );
  DFF \sreg_reg[1883]  ( .D(c[1887]), .CLK(clk), .RST(rst), .Q(sreg[1883]) );
  DFF \sreg_reg[1882]  ( .D(c[1886]), .CLK(clk), .RST(rst), .Q(sreg[1882]) );
  DFF \sreg_reg[1881]  ( .D(c[1885]), .CLK(clk), .RST(rst), .Q(sreg[1881]) );
  DFF \sreg_reg[1880]  ( .D(c[1884]), .CLK(clk), .RST(rst), .Q(sreg[1880]) );
  DFF \sreg_reg[1879]  ( .D(c[1883]), .CLK(clk), .RST(rst), .Q(sreg[1879]) );
  DFF \sreg_reg[1878]  ( .D(c[1882]), .CLK(clk), .RST(rst), .Q(sreg[1878]) );
  DFF \sreg_reg[1877]  ( .D(c[1881]), .CLK(clk), .RST(rst), .Q(sreg[1877]) );
  DFF \sreg_reg[1876]  ( .D(c[1880]), .CLK(clk), .RST(rst), .Q(sreg[1876]) );
  DFF \sreg_reg[1875]  ( .D(c[1879]), .CLK(clk), .RST(rst), .Q(sreg[1875]) );
  DFF \sreg_reg[1874]  ( .D(c[1878]), .CLK(clk), .RST(rst), .Q(sreg[1874]) );
  DFF \sreg_reg[1873]  ( .D(c[1877]), .CLK(clk), .RST(rst), .Q(sreg[1873]) );
  DFF \sreg_reg[1872]  ( .D(c[1876]), .CLK(clk), .RST(rst), .Q(sreg[1872]) );
  DFF \sreg_reg[1871]  ( .D(c[1875]), .CLK(clk), .RST(rst), .Q(sreg[1871]) );
  DFF \sreg_reg[1870]  ( .D(c[1874]), .CLK(clk), .RST(rst), .Q(sreg[1870]) );
  DFF \sreg_reg[1869]  ( .D(c[1873]), .CLK(clk), .RST(rst), .Q(sreg[1869]) );
  DFF \sreg_reg[1868]  ( .D(c[1872]), .CLK(clk), .RST(rst), .Q(sreg[1868]) );
  DFF \sreg_reg[1867]  ( .D(c[1871]), .CLK(clk), .RST(rst), .Q(sreg[1867]) );
  DFF \sreg_reg[1866]  ( .D(c[1870]), .CLK(clk), .RST(rst), .Q(sreg[1866]) );
  DFF \sreg_reg[1865]  ( .D(c[1869]), .CLK(clk), .RST(rst), .Q(sreg[1865]) );
  DFF \sreg_reg[1864]  ( .D(c[1868]), .CLK(clk), .RST(rst), .Q(sreg[1864]) );
  DFF \sreg_reg[1863]  ( .D(c[1867]), .CLK(clk), .RST(rst), .Q(sreg[1863]) );
  DFF \sreg_reg[1862]  ( .D(c[1866]), .CLK(clk), .RST(rst), .Q(sreg[1862]) );
  DFF \sreg_reg[1861]  ( .D(c[1865]), .CLK(clk), .RST(rst), .Q(sreg[1861]) );
  DFF \sreg_reg[1860]  ( .D(c[1864]), .CLK(clk), .RST(rst), .Q(sreg[1860]) );
  DFF \sreg_reg[1859]  ( .D(c[1863]), .CLK(clk), .RST(rst), .Q(sreg[1859]) );
  DFF \sreg_reg[1858]  ( .D(c[1862]), .CLK(clk), .RST(rst), .Q(sreg[1858]) );
  DFF \sreg_reg[1857]  ( .D(c[1861]), .CLK(clk), .RST(rst), .Q(sreg[1857]) );
  DFF \sreg_reg[1856]  ( .D(c[1860]), .CLK(clk), .RST(rst), .Q(sreg[1856]) );
  DFF \sreg_reg[1855]  ( .D(c[1859]), .CLK(clk), .RST(rst), .Q(sreg[1855]) );
  DFF \sreg_reg[1854]  ( .D(c[1858]), .CLK(clk), .RST(rst), .Q(sreg[1854]) );
  DFF \sreg_reg[1853]  ( .D(c[1857]), .CLK(clk), .RST(rst), .Q(sreg[1853]) );
  DFF \sreg_reg[1852]  ( .D(c[1856]), .CLK(clk), .RST(rst), .Q(sreg[1852]) );
  DFF \sreg_reg[1851]  ( .D(c[1855]), .CLK(clk), .RST(rst), .Q(sreg[1851]) );
  DFF \sreg_reg[1850]  ( .D(c[1854]), .CLK(clk), .RST(rst), .Q(sreg[1850]) );
  DFF \sreg_reg[1849]  ( .D(c[1853]), .CLK(clk), .RST(rst), .Q(sreg[1849]) );
  DFF \sreg_reg[1848]  ( .D(c[1852]), .CLK(clk), .RST(rst), .Q(sreg[1848]) );
  DFF \sreg_reg[1847]  ( .D(c[1851]), .CLK(clk), .RST(rst), .Q(sreg[1847]) );
  DFF \sreg_reg[1846]  ( .D(c[1850]), .CLK(clk), .RST(rst), .Q(sreg[1846]) );
  DFF \sreg_reg[1845]  ( .D(c[1849]), .CLK(clk), .RST(rst), .Q(sreg[1845]) );
  DFF \sreg_reg[1844]  ( .D(c[1848]), .CLK(clk), .RST(rst), .Q(sreg[1844]) );
  DFF \sreg_reg[1843]  ( .D(c[1847]), .CLK(clk), .RST(rst), .Q(sreg[1843]) );
  DFF \sreg_reg[1842]  ( .D(c[1846]), .CLK(clk), .RST(rst), .Q(sreg[1842]) );
  DFF \sreg_reg[1841]  ( .D(c[1845]), .CLK(clk), .RST(rst), .Q(sreg[1841]) );
  DFF \sreg_reg[1840]  ( .D(c[1844]), .CLK(clk), .RST(rst), .Q(sreg[1840]) );
  DFF \sreg_reg[1839]  ( .D(c[1843]), .CLK(clk), .RST(rst), .Q(sreg[1839]) );
  DFF \sreg_reg[1838]  ( .D(c[1842]), .CLK(clk), .RST(rst), .Q(sreg[1838]) );
  DFF \sreg_reg[1837]  ( .D(c[1841]), .CLK(clk), .RST(rst), .Q(sreg[1837]) );
  DFF \sreg_reg[1836]  ( .D(c[1840]), .CLK(clk), .RST(rst), .Q(sreg[1836]) );
  DFF \sreg_reg[1835]  ( .D(c[1839]), .CLK(clk), .RST(rst), .Q(sreg[1835]) );
  DFF \sreg_reg[1834]  ( .D(c[1838]), .CLK(clk), .RST(rst), .Q(sreg[1834]) );
  DFF \sreg_reg[1833]  ( .D(c[1837]), .CLK(clk), .RST(rst), .Q(sreg[1833]) );
  DFF \sreg_reg[1832]  ( .D(c[1836]), .CLK(clk), .RST(rst), .Q(sreg[1832]) );
  DFF \sreg_reg[1831]  ( .D(c[1835]), .CLK(clk), .RST(rst), .Q(sreg[1831]) );
  DFF \sreg_reg[1830]  ( .D(c[1834]), .CLK(clk), .RST(rst), .Q(sreg[1830]) );
  DFF \sreg_reg[1829]  ( .D(c[1833]), .CLK(clk), .RST(rst), .Q(sreg[1829]) );
  DFF \sreg_reg[1828]  ( .D(c[1832]), .CLK(clk), .RST(rst), .Q(sreg[1828]) );
  DFF \sreg_reg[1827]  ( .D(c[1831]), .CLK(clk), .RST(rst), .Q(sreg[1827]) );
  DFF \sreg_reg[1826]  ( .D(c[1830]), .CLK(clk), .RST(rst), .Q(sreg[1826]) );
  DFF \sreg_reg[1825]  ( .D(c[1829]), .CLK(clk), .RST(rst), .Q(sreg[1825]) );
  DFF \sreg_reg[1824]  ( .D(c[1828]), .CLK(clk), .RST(rst), .Q(sreg[1824]) );
  DFF \sreg_reg[1823]  ( .D(c[1827]), .CLK(clk), .RST(rst), .Q(sreg[1823]) );
  DFF \sreg_reg[1822]  ( .D(c[1826]), .CLK(clk), .RST(rst), .Q(sreg[1822]) );
  DFF \sreg_reg[1821]  ( .D(c[1825]), .CLK(clk), .RST(rst), .Q(sreg[1821]) );
  DFF \sreg_reg[1820]  ( .D(c[1824]), .CLK(clk), .RST(rst), .Q(sreg[1820]) );
  DFF \sreg_reg[1819]  ( .D(c[1823]), .CLK(clk), .RST(rst), .Q(sreg[1819]) );
  DFF \sreg_reg[1818]  ( .D(c[1822]), .CLK(clk), .RST(rst), .Q(sreg[1818]) );
  DFF \sreg_reg[1817]  ( .D(c[1821]), .CLK(clk), .RST(rst), .Q(sreg[1817]) );
  DFF \sreg_reg[1816]  ( .D(c[1820]), .CLK(clk), .RST(rst), .Q(sreg[1816]) );
  DFF \sreg_reg[1815]  ( .D(c[1819]), .CLK(clk), .RST(rst), .Q(sreg[1815]) );
  DFF \sreg_reg[1814]  ( .D(c[1818]), .CLK(clk), .RST(rst), .Q(sreg[1814]) );
  DFF \sreg_reg[1813]  ( .D(c[1817]), .CLK(clk), .RST(rst), .Q(sreg[1813]) );
  DFF \sreg_reg[1812]  ( .D(c[1816]), .CLK(clk), .RST(rst), .Q(sreg[1812]) );
  DFF \sreg_reg[1811]  ( .D(c[1815]), .CLK(clk), .RST(rst), .Q(sreg[1811]) );
  DFF \sreg_reg[1810]  ( .D(c[1814]), .CLK(clk), .RST(rst), .Q(sreg[1810]) );
  DFF \sreg_reg[1809]  ( .D(c[1813]), .CLK(clk), .RST(rst), .Q(sreg[1809]) );
  DFF \sreg_reg[1808]  ( .D(c[1812]), .CLK(clk), .RST(rst), .Q(sreg[1808]) );
  DFF \sreg_reg[1807]  ( .D(c[1811]), .CLK(clk), .RST(rst), .Q(sreg[1807]) );
  DFF \sreg_reg[1806]  ( .D(c[1810]), .CLK(clk), .RST(rst), .Q(sreg[1806]) );
  DFF \sreg_reg[1805]  ( .D(c[1809]), .CLK(clk), .RST(rst), .Q(sreg[1805]) );
  DFF \sreg_reg[1804]  ( .D(c[1808]), .CLK(clk), .RST(rst), .Q(sreg[1804]) );
  DFF \sreg_reg[1803]  ( .D(c[1807]), .CLK(clk), .RST(rst), .Q(sreg[1803]) );
  DFF \sreg_reg[1802]  ( .D(c[1806]), .CLK(clk), .RST(rst), .Q(sreg[1802]) );
  DFF \sreg_reg[1801]  ( .D(c[1805]), .CLK(clk), .RST(rst), .Q(sreg[1801]) );
  DFF \sreg_reg[1800]  ( .D(c[1804]), .CLK(clk), .RST(rst), .Q(sreg[1800]) );
  DFF \sreg_reg[1799]  ( .D(c[1803]), .CLK(clk), .RST(rst), .Q(sreg[1799]) );
  DFF \sreg_reg[1798]  ( .D(c[1802]), .CLK(clk), .RST(rst), .Q(sreg[1798]) );
  DFF \sreg_reg[1797]  ( .D(c[1801]), .CLK(clk), .RST(rst), .Q(sreg[1797]) );
  DFF \sreg_reg[1796]  ( .D(c[1800]), .CLK(clk), .RST(rst), .Q(sreg[1796]) );
  DFF \sreg_reg[1795]  ( .D(c[1799]), .CLK(clk), .RST(rst), .Q(sreg[1795]) );
  DFF \sreg_reg[1794]  ( .D(c[1798]), .CLK(clk), .RST(rst), .Q(sreg[1794]) );
  DFF \sreg_reg[1793]  ( .D(c[1797]), .CLK(clk), .RST(rst), .Q(sreg[1793]) );
  DFF \sreg_reg[1792]  ( .D(c[1796]), .CLK(clk), .RST(rst), .Q(sreg[1792]) );
  DFF \sreg_reg[1791]  ( .D(c[1795]), .CLK(clk), .RST(rst), .Q(sreg[1791]) );
  DFF \sreg_reg[1790]  ( .D(c[1794]), .CLK(clk), .RST(rst), .Q(sreg[1790]) );
  DFF \sreg_reg[1789]  ( .D(c[1793]), .CLK(clk), .RST(rst), .Q(sreg[1789]) );
  DFF \sreg_reg[1788]  ( .D(c[1792]), .CLK(clk), .RST(rst), .Q(sreg[1788]) );
  DFF \sreg_reg[1787]  ( .D(c[1791]), .CLK(clk), .RST(rst), .Q(sreg[1787]) );
  DFF \sreg_reg[1786]  ( .D(c[1790]), .CLK(clk), .RST(rst), .Q(sreg[1786]) );
  DFF \sreg_reg[1785]  ( .D(c[1789]), .CLK(clk), .RST(rst), .Q(sreg[1785]) );
  DFF \sreg_reg[1784]  ( .D(c[1788]), .CLK(clk), .RST(rst), .Q(sreg[1784]) );
  DFF \sreg_reg[1783]  ( .D(c[1787]), .CLK(clk), .RST(rst), .Q(sreg[1783]) );
  DFF \sreg_reg[1782]  ( .D(c[1786]), .CLK(clk), .RST(rst), .Q(sreg[1782]) );
  DFF \sreg_reg[1781]  ( .D(c[1785]), .CLK(clk), .RST(rst), .Q(sreg[1781]) );
  DFF \sreg_reg[1780]  ( .D(c[1784]), .CLK(clk), .RST(rst), .Q(sreg[1780]) );
  DFF \sreg_reg[1779]  ( .D(c[1783]), .CLK(clk), .RST(rst), .Q(sreg[1779]) );
  DFF \sreg_reg[1778]  ( .D(c[1782]), .CLK(clk), .RST(rst), .Q(sreg[1778]) );
  DFF \sreg_reg[1777]  ( .D(c[1781]), .CLK(clk), .RST(rst), .Q(sreg[1777]) );
  DFF \sreg_reg[1776]  ( .D(c[1780]), .CLK(clk), .RST(rst), .Q(sreg[1776]) );
  DFF \sreg_reg[1775]  ( .D(c[1779]), .CLK(clk), .RST(rst), .Q(sreg[1775]) );
  DFF \sreg_reg[1774]  ( .D(c[1778]), .CLK(clk), .RST(rst), .Q(sreg[1774]) );
  DFF \sreg_reg[1773]  ( .D(c[1777]), .CLK(clk), .RST(rst), .Q(sreg[1773]) );
  DFF \sreg_reg[1772]  ( .D(c[1776]), .CLK(clk), .RST(rst), .Q(sreg[1772]) );
  DFF \sreg_reg[1771]  ( .D(c[1775]), .CLK(clk), .RST(rst), .Q(sreg[1771]) );
  DFF \sreg_reg[1770]  ( .D(c[1774]), .CLK(clk), .RST(rst), .Q(sreg[1770]) );
  DFF \sreg_reg[1769]  ( .D(c[1773]), .CLK(clk), .RST(rst), .Q(sreg[1769]) );
  DFF \sreg_reg[1768]  ( .D(c[1772]), .CLK(clk), .RST(rst), .Q(sreg[1768]) );
  DFF \sreg_reg[1767]  ( .D(c[1771]), .CLK(clk), .RST(rst), .Q(sreg[1767]) );
  DFF \sreg_reg[1766]  ( .D(c[1770]), .CLK(clk), .RST(rst), .Q(sreg[1766]) );
  DFF \sreg_reg[1765]  ( .D(c[1769]), .CLK(clk), .RST(rst), .Q(sreg[1765]) );
  DFF \sreg_reg[1764]  ( .D(c[1768]), .CLK(clk), .RST(rst), .Q(sreg[1764]) );
  DFF \sreg_reg[1763]  ( .D(c[1767]), .CLK(clk), .RST(rst), .Q(sreg[1763]) );
  DFF \sreg_reg[1762]  ( .D(c[1766]), .CLK(clk), .RST(rst), .Q(sreg[1762]) );
  DFF \sreg_reg[1761]  ( .D(c[1765]), .CLK(clk), .RST(rst), .Q(sreg[1761]) );
  DFF \sreg_reg[1760]  ( .D(c[1764]), .CLK(clk), .RST(rst), .Q(sreg[1760]) );
  DFF \sreg_reg[1759]  ( .D(c[1763]), .CLK(clk), .RST(rst), .Q(sreg[1759]) );
  DFF \sreg_reg[1758]  ( .D(c[1762]), .CLK(clk), .RST(rst), .Q(sreg[1758]) );
  DFF \sreg_reg[1757]  ( .D(c[1761]), .CLK(clk), .RST(rst), .Q(sreg[1757]) );
  DFF \sreg_reg[1756]  ( .D(c[1760]), .CLK(clk), .RST(rst), .Q(sreg[1756]) );
  DFF \sreg_reg[1755]  ( .D(c[1759]), .CLK(clk), .RST(rst), .Q(sreg[1755]) );
  DFF \sreg_reg[1754]  ( .D(c[1758]), .CLK(clk), .RST(rst), .Q(sreg[1754]) );
  DFF \sreg_reg[1753]  ( .D(c[1757]), .CLK(clk), .RST(rst), .Q(sreg[1753]) );
  DFF \sreg_reg[1752]  ( .D(c[1756]), .CLK(clk), .RST(rst), .Q(sreg[1752]) );
  DFF \sreg_reg[1751]  ( .D(c[1755]), .CLK(clk), .RST(rst), .Q(sreg[1751]) );
  DFF \sreg_reg[1750]  ( .D(c[1754]), .CLK(clk), .RST(rst), .Q(sreg[1750]) );
  DFF \sreg_reg[1749]  ( .D(c[1753]), .CLK(clk), .RST(rst), .Q(sreg[1749]) );
  DFF \sreg_reg[1748]  ( .D(c[1752]), .CLK(clk), .RST(rst), .Q(sreg[1748]) );
  DFF \sreg_reg[1747]  ( .D(c[1751]), .CLK(clk), .RST(rst), .Q(sreg[1747]) );
  DFF \sreg_reg[1746]  ( .D(c[1750]), .CLK(clk), .RST(rst), .Q(sreg[1746]) );
  DFF \sreg_reg[1745]  ( .D(c[1749]), .CLK(clk), .RST(rst), .Q(sreg[1745]) );
  DFF \sreg_reg[1744]  ( .D(c[1748]), .CLK(clk), .RST(rst), .Q(sreg[1744]) );
  DFF \sreg_reg[1743]  ( .D(c[1747]), .CLK(clk), .RST(rst), .Q(sreg[1743]) );
  DFF \sreg_reg[1742]  ( .D(c[1746]), .CLK(clk), .RST(rst), .Q(sreg[1742]) );
  DFF \sreg_reg[1741]  ( .D(c[1745]), .CLK(clk), .RST(rst), .Q(sreg[1741]) );
  DFF \sreg_reg[1740]  ( .D(c[1744]), .CLK(clk), .RST(rst), .Q(sreg[1740]) );
  DFF \sreg_reg[1739]  ( .D(c[1743]), .CLK(clk), .RST(rst), .Q(sreg[1739]) );
  DFF \sreg_reg[1738]  ( .D(c[1742]), .CLK(clk), .RST(rst), .Q(sreg[1738]) );
  DFF \sreg_reg[1737]  ( .D(c[1741]), .CLK(clk), .RST(rst), .Q(sreg[1737]) );
  DFF \sreg_reg[1736]  ( .D(c[1740]), .CLK(clk), .RST(rst), .Q(sreg[1736]) );
  DFF \sreg_reg[1735]  ( .D(c[1739]), .CLK(clk), .RST(rst), .Q(sreg[1735]) );
  DFF \sreg_reg[1734]  ( .D(c[1738]), .CLK(clk), .RST(rst), .Q(sreg[1734]) );
  DFF \sreg_reg[1733]  ( .D(c[1737]), .CLK(clk), .RST(rst), .Q(sreg[1733]) );
  DFF \sreg_reg[1732]  ( .D(c[1736]), .CLK(clk), .RST(rst), .Q(sreg[1732]) );
  DFF \sreg_reg[1731]  ( .D(c[1735]), .CLK(clk), .RST(rst), .Q(sreg[1731]) );
  DFF \sreg_reg[1730]  ( .D(c[1734]), .CLK(clk), .RST(rst), .Q(sreg[1730]) );
  DFF \sreg_reg[1729]  ( .D(c[1733]), .CLK(clk), .RST(rst), .Q(sreg[1729]) );
  DFF \sreg_reg[1728]  ( .D(c[1732]), .CLK(clk), .RST(rst), .Q(sreg[1728]) );
  DFF \sreg_reg[1727]  ( .D(c[1731]), .CLK(clk), .RST(rst), .Q(sreg[1727]) );
  DFF \sreg_reg[1726]  ( .D(c[1730]), .CLK(clk), .RST(rst), .Q(sreg[1726]) );
  DFF \sreg_reg[1725]  ( .D(c[1729]), .CLK(clk), .RST(rst), .Q(sreg[1725]) );
  DFF \sreg_reg[1724]  ( .D(c[1728]), .CLK(clk), .RST(rst), .Q(sreg[1724]) );
  DFF \sreg_reg[1723]  ( .D(c[1727]), .CLK(clk), .RST(rst), .Q(sreg[1723]) );
  DFF \sreg_reg[1722]  ( .D(c[1726]), .CLK(clk), .RST(rst), .Q(sreg[1722]) );
  DFF \sreg_reg[1721]  ( .D(c[1725]), .CLK(clk), .RST(rst), .Q(sreg[1721]) );
  DFF \sreg_reg[1720]  ( .D(c[1724]), .CLK(clk), .RST(rst), .Q(sreg[1720]) );
  DFF \sreg_reg[1719]  ( .D(c[1723]), .CLK(clk), .RST(rst), .Q(sreg[1719]) );
  DFF \sreg_reg[1718]  ( .D(c[1722]), .CLK(clk), .RST(rst), .Q(sreg[1718]) );
  DFF \sreg_reg[1717]  ( .D(c[1721]), .CLK(clk), .RST(rst), .Q(sreg[1717]) );
  DFF \sreg_reg[1716]  ( .D(c[1720]), .CLK(clk), .RST(rst), .Q(sreg[1716]) );
  DFF \sreg_reg[1715]  ( .D(c[1719]), .CLK(clk), .RST(rst), .Q(sreg[1715]) );
  DFF \sreg_reg[1714]  ( .D(c[1718]), .CLK(clk), .RST(rst), .Q(sreg[1714]) );
  DFF \sreg_reg[1713]  ( .D(c[1717]), .CLK(clk), .RST(rst), .Q(sreg[1713]) );
  DFF \sreg_reg[1712]  ( .D(c[1716]), .CLK(clk), .RST(rst), .Q(sreg[1712]) );
  DFF \sreg_reg[1711]  ( .D(c[1715]), .CLK(clk), .RST(rst), .Q(sreg[1711]) );
  DFF \sreg_reg[1710]  ( .D(c[1714]), .CLK(clk), .RST(rst), .Q(sreg[1710]) );
  DFF \sreg_reg[1709]  ( .D(c[1713]), .CLK(clk), .RST(rst), .Q(sreg[1709]) );
  DFF \sreg_reg[1708]  ( .D(c[1712]), .CLK(clk), .RST(rst), .Q(sreg[1708]) );
  DFF \sreg_reg[1707]  ( .D(c[1711]), .CLK(clk), .RST(rst), .Q(sreg[1707]) );
  DFF \sreg_reg[1706]  ( .D(c[1710]), .CLK(clk), .RST(rst), .Q(sreg[1706]) );
  DFF \sreg_reg[1705]  ( .D(c[1709]), .CLK(clk), .RST(rst), .Q(sreg[1705]) );
  DFF \sreg_reg[1704]  ( .D(c[1708]), .CLK(clk), .RST(rst), .Q(sreg[1704]) );
  DFF \sreg_reg[1703]  ( .D(c[1707]), .CLK(clk), .RST(rst), .Q(sreg[1703]) );
  DFF \sreg_reg[1702]  ( .D(c[1706]), .CLK(clk), .RST(rst), .Q(sreg[1702]) );
  DFF \sreg_reg[1701]  ( .D(c[1705]), .CLK(clk), .RST(rst), .Q(sreg[1701]) );
  DFF \sreg_reg[1700]  ( .D(c[1704]), .CLK(clk), .RST(rst), .Q(sreg[1700]) );
  DFF \sreg_reg[1699]  ( .D(c[1703]), .CLK(clk), .RST(rst), .Q(sreg[1699]) );
  DFF \sreg_reg[1698]  ( .D(c[1702]), .CLK(clk), .RST(rst), .Q(sreg[1698]) );
  DFF \sreg_reg[1697]  ( .D(c[1701]), .CLK(clk), .RST(rst), .Q(sreg[1697]) );
  DFF \sreg_reg[1696]  ( .D(c[1700]), .CLK(clk), .RST(rst), .Q(sreg[1696]) );
  DFF \sreg_reg[1695]  ( .D(c[1699]), .CLK(clk), .RST(rst), .Q(sreg[1695]) );
  DFF \sreg_reg[1694]  ( .D(c[1698]), .CLK(clk), .RST(rst), .Q(sreg[1694]) );
  DFF \sreg_reg[1693]  ( .D(c[1697]), .CLK(clk), .RST(rst), .Q(sreg[1693]) );
  DFF \sreg_reg[1692]  ( .D(c[1696]), .CLK(clk), .RST(rst), .Q(sreg[1692]) );
  DFF \sreg_reg[1691]  ( .D(c[1695]), .CLK(clk), .RST(rst), .Q(sreg[1691]) );
  DFF \sreg_reg[1690]  ( .D(c[1694]), .CLK(clk), .RST(rst), .Q(sreg[1690]) );
  DFF \sreg_reg[1689]  ( .D(c[1693]), .CLK(clk), .RST(rst), .Q(sreg[1689]) );
  DFF \sreg_reg[1688]  ( .D(c[1692]), .CLK(clk), .RST(rst), .Q(sreg[1688]) );
  DFF \sreg_reg[1687]  ( .D(c[1691]), .CLK(clk), .RST(rst), .Q(sreg[1687]) );
  DFF \sreg_reg[1686]  ( .D(c[1690]), .CLK(clk), .RST(rst), .Q(sreg[1686]) );
  DFF \sreg_reg[1685]  ( .D(c[1689]), .CLK(clk), .RST(rst), .Q(sreg[1685]) );
  DFF \sreg_reg[1684]  ( .D(c[1688]), .CLK(clk), .RST(rst), .Q(sreg[1684]) );
  DFF \sreg_reg[1683]  ( .D(c[1687]), .CLK(clk), .RST(rst), .Q(sreg[1683]) );
  DFF \sreg_reg[1682]  ( .D(c[1686]), .CLK(clk), .RST(rst), .Q(sreg[1682]) );
  DFF \sreg_reg[1681]  ( .D(c[1685]), .CLK(clk), .RST(rst), .Q(sreg[1681]) );
  DFF \sreg_reg[1680]  ( .D(c[1684]), .CLK(clk), .RST(rst), .Q(sreg[1680]) );
  DFF \sreg_reg[1679]  ( .D(c[1683]), .CLK(clk), .RST(rst), .Q(sreg[1679]) );
  DFF \sreg_reg[1678]  ( .D(c[1682]), .CLK(clk), .RST(rst), .Q(sreg[1678]) );
  DFF \sreg_reg[1677]  ( .D(c[1681]), .CLK(clk), .RST(rst), .Q(sreg[1677]) );
  DFF \sreg_reg[1676]  ( .D(c[1680]), .CLK(clk), .RST(rst), .Q(sreg[1676]) );
  DFF \sreg_reg[1675]  ( .D(c[1679]), .CLK(clk), .RST(rst), .Q(sreg[1675]) );
  DFF \sreg_reg[1674]  ( .D(c[1678]), .CLK(clk), .RST(rst), .Q(sreg[1674]) );
  DFF \sreg_reg[1673]  ( .D(c[1677]), .CLK(clk), .RST(rst), .Q(sreg[1673]) );
  DFF \sreg_reg[1672]  ( .D(c[1676]), .CLK(clk), .RST(rst), .Q(sreg[1672]) );
  DFF \sreg_reg[1671]  ( .D(c[1675]), .CLK(clk), .RST(rst), .Q(sreg[1671]) );
  DFF \sreg_reg[1670]  ( .D(c[1674]), .CLK(clk), .RST(rst), .Q(sreg[1670]) );
  DFF \sreg_reg[1669]  ( .D(c[1673]), .CLK(clk), .RST(rst), .Q(sreg[1669]) );
  DFF \sreg_reg[1668]  ( .D(c[1672]), .CLK(clk), .RST(rst), .Q(sreg[1668]) );
  DFF \sreg_reg[1667]  ( .D(c[1671]), .CLK(clk), .RST(rst), .Q(sreg[1667]) );
  DFF \sreg_reg[1666]  ( .D(c[1670]), .CLK(clk), .RST(rst), .Q(sreg[1666]) );
  DFF \sreg_reg[1665]  ( .D(c[1669]), .CLK(clk), .RST(rst), .Q(sreg[1665]) );
  DFF \sreg_reg[1664]  ( .D(c[1668]), .CLK(clk), .RST(rst), .Q(sreg[1664]) );
  DFF \sreg_reg[1663]  ( .D(c[1667]), .CLK(clk), .RST(rst), .Q(sreg[1663]) );
  DFF \sreg_reg[1662]  ( .D(c[1666]), .CLK(clk), .RST(rst), .Q(sreg[1662]) );
  DFF \sreg_reg[1661]  ( .D(c[1665]), .CLK(clk), .RST(rst), .Q(sreg[1661]) );
  DFF \sreg_reg[1660]  ( .D(c[1664]), .CLK(clk), .RST(rst), .Q(sreg[1660]) );
  DFF \sreg_reg[1659]  ( .D(c[1663]), .CLK(clk), .RST(rst), .Q(sreg[1659]) );
  DFF \sreg_reg[1658]  ( .D(c[1662]), .CLK(clk), .RST(rst), .Q(sreg[1658]) );
  DFF \sreg_reg[1657]  ( .D(c[1661]), .CLK(clk), .RST(rst), .Q(sreg[1657]) );
  DFF \sreg_reg[1656]  ( .D(c[1660]), .CLK(clk), .RST(rst), .Q(sreg[1656]) );
  DFF \sreg_reg[1655]  ( .D(c[1659]), .CLK(clk), .RST(rst), .Q(sreg[1655]) );
  DFF \sreg_reg[1654]  ( .D(c[1658]), .CLK(clk), .RST(rst), .Q(sreg[1654]) );
  DFF \sreg_reg[1653]  ( .D(c[1657]), .CLK(clk), .RST(rst), .Q(sreg[1653]) );
  DFF \sreg_reg[1652]  ( .D(c[1656]), .CLK(clk), .RST(rst), .Q(sreg[1652]) );
  DFF \sreg_reg[1651]  ( .D(c[1655]), .CLK(clk), .RST(rst), .Q(sreg[1651]) );
  DFF \sreg_reg[1650]  ( .D(c[1654]), .CLK(clk), .RST(rst), .Q(sreg[1650]) );
  DFF \sreg_reg[1649]  ( .D(c[1653]), .CLK(clk), .RST(rst), .Q(sreg[1649]) );
  DFF \sreg_reg[1648]  ( .D(c[1652]), .CLK(clk), .RST(rst), .Q(sreg[1648]) );
  DFF \sreg_reg[1647]  ( .D(c[1651]), .CLK(clk), .RST(rst), .Q(sreg[1647]) );
  DFF \sreg_reg[1646]  ( .D(c[1650]), .CLK(clk), .RST(rst), .Q(sreg[1646]) );
  DFF \sreg_reg[1645]  ( .D(c[1649]), .CLK(clk), .RST(rst), .Q(sreg[1645]) );
  DFF \sreg_reg[1644]  ( .D(c[1648]), .CLK(clk), .RST(rst), .Q(sreg[1644]) );
  DFF \sreg_reg[1643]  ( .D(c[1647]), .CLK(clk), .RST(rst), .Q(sreg[1643]) );
  DFF \sreg_reg[1642]  ( .D(c[1646]), .CLK(clk), .RST(rst), .Q(sreg[1642]) );
  DFF \sreg_reg[1641]  ( .D(c[1645]), .CLK(clk), .RST(rst), .Q(sreg[1641]) );
  DFF \sreg_reg[1640]  ( .D(c[1644]), .CLK(clk), .RST(rst), .Q(sreg[1640]) );
  DFF \sreg_reg[1639]  ( .D(c[1643]), .CLK(clk), .RST(rst), .Q(sreg[1639]) );
  DFF \sreg_reg[1638]  ( .D(c[1642]), .CLK(clk), .RST(rst), .Q(sreg[1638]) );
  DFF \sreg_reg[1637]  ( .D(c[1641]), .CLK(clk), .RST(rst), .Q(sreg[1637]) );
  DFF \sreg_reg[1636]  ( .D(c[1640]), .CLK(clk), .RST(rst), .Q(sreg[1636]) );
  DFF \sreg_reg[1635]  ( .D(c[1639]), .CLK(clk), .RST(rst), .Q(sreg[1635]) );
  DFF \sreg_reg[1634]  ( .D(c[1638]), .CLK(clk), .RST(rst), .Q(sreg[1634]) );
  DFF \sreg_reg[1633]  ( .D(c[1637]), .CLK(clk), .RST(rst), .Q(sreg[1633]) );
  DFF \sreg_reg[1632]  ( .D(c[1636]), .CLK(clk), .RST(rst), .Q(sreg[1632]) );
  DFF \sreg_reg[1631]  ( .D(c[1635]), .CLK(clk), .RST(rst), .Q(sreg[1631]) );
  DFF \sreg_reg[1630]  ( .D(c[1634]), .CLK(clk), .RST(rst), .Q(sreg[1630]) );
  DFF \sreg_reg[1629]  ( .D(c[1633]), .CLK(clk), .RST(rst), .Q(sreg[1629]) );
  DFF \sreg_reg[1628]  ( .D(c[1632]), .CLK(clk), .RST(rst), .Q(sreg[1628]) );
  DFF \sreg_reg[1627]  ( .D(c[1631]), .CLK(clk), .RST(rst), .Q(sreg[1627]) );
  DFF \sreg_reg[1626]  ( .D(c[1630]), .CLK(clk), .RST(rst), .Q(sreg[1626]) );
  DFF \sreg_reg[1625]  ( .D(c[1629]), .CLK(clk), .RST(rst), .Q(sreg[1625]) );
  DFF \sreg_reg[1624]  ( .D(c[1628]), .CLK(clk), .RST(rst), .Q(sreg[1624]) );
  DFF \sreg_reg[1623]  ( .D(c[1627]), .CLK(clk), .RST(rst), .Q(sreg[1623]) );
  DFF \sreg_reg[1622]  ( .D(c[1626]), .CLK(clk), .RST(rst), .Q(sreg[1622]) );
  DFF \sreg_reg[1621]  ( .D(c[1625]), .CLK(clk), .RST(rst), .Q(sreg[1621]) );
  DFF \sreg_reg[1620]  ( .D(c[1624]), .CLK(clk), .RST(rst), .Q(sreg[1620]) );
  DFF \sreg_reg[1619]  ( .D(c[1623]), .CLK(clk), .RST(rst), .Q(sreg[1619]) );
  DFF \sreg_reg[1618]  ( .D(c[1622]), .CLK(clk), .RST(rst), .Q(sreg[1618]) );
  DFF \sreg_reg[1617]  ( .D(c[1621]), .CLK(clk), .RST(rst), .Q(sreg[1617]) );
  DFF \sreg_reg[1616]  ( .D(c[1620]), .CLK(clk), .RST(rst), .Q(sreg[1616]) );
  DFF \sreg_reg[1615]  ( .D(c[1619]), .CLK(clk), .RST(rst), .Q(sreg[1615]) );
  DFF \sreg_reg[1614]  ( .D(c[1618]), .CLK(clk), .RST(rst), .Q(sreg[1614]) );
  DFF \sreg_reg[1613]  ( .D(c[1617]), .CLK(clk), .RST(rst), .Q(sreg[1613]) );
  DFF \sreg_reg[1612]  ( .D(c[1616]), .CLK(clk), .RST(rst), .Q(sreg[1612]) );
  DFF \sreg_reg[1611]  ( .D(c[1615]), .CLK(clk), .RST(rst), .Q(sreg[1611]) );
  DFF \sreg_reg[1610]  ( .D(c[1614]), .CLK(clk), .RST(rst), .Q(sreg[1610]) );
  DFF \sreg_reg[1609]  ( .D(c[1613]), .CLK(clk), .RST(rst), .Q(sreg[1609]) );
  DFF \sreg_reg[1608]  ( .D(c[1612]), .CLK(clk), .RST(rst), .Q(sreg[1608]) );
  DFF \sreg_reg[1607]  ( .D(c[1611]), .CLK(clk), .RST(rst), .Q(sreg[1607]) );
  DFF \sreg_reg[1606]  ( .D(c[1610]), .CLK(clk), .RST(rst), .Q(sreg[1606]) );
  DFF \sreg_reg[1605]  ( .D(c[1609]), .CLK(clk), .RST(rst), .Q(sreg[1605]) );
  DFF \sreg_reg[1604]  ( .D(c[1608]), .CLK(clk), .RST(rst), .Q(sreg[1604]) );
  DFF \sreg_reg[1603]  ( .D(c[1607]), .CLK(clk), .RST(rst), .Q(sreg[1603]) );
  DFF \sreg_reg[1602]  ( .D(c[1606]), .CLK(clk), .RST(rst), .Q(sreg[1602]) );
  DFF \sreg_reg[1601]  ( .D(c[1605]), .CLK(clk), .RST(rst), .Q(sreg[1601]) );
  DFF \sreg_reg[1600]  ( .D(c[1604]), .CLK(clk), .RST(rst), .Q(sreg[1600]) );
  DFF \sreg_reg[1599]  ( .D(c[1603]), .CLK(clk), .RST(rst), .Q(sreg[1599]) );
  DFF \sreg_reg[1598]  ( .D(c[1602]), .CLK(clk), .RST(rst), .Q(sreg[1598]) );
  DFF \sreg_reg[1597]  ( .D(c[1601]), .CLK(clk), .RST(rst), .Q(sreg[1597]) );
  DFF \sreg_reg[1596]  ( .D(c[1600]), .CLK(clk), .RST(rst), .Q(sreg[1596]) );
  DFF \sreg_reg[1595]  ( .D(c[1599]), .CLK(clk), .RST(rst), .Q(sreg[1595]) );
  DFF \sreg_reg[1594]  ( .D(c[1598]), .CLK(clk), .RST(rst), .Q(sreg[1594]) );
  DFF \sreg_reg[1593]  ( .D(c[1597]), .CLK(clk), .RST(rst), .Q(sreg[1593]) );
  DFF \sreg_reg[1592]  ( .D(c[1596]), .CLK(clk), .RST(rst), .Q(sreg[1592]) );
  DFF \sreg_reg[1591]  ( .D(c[1595]), .CLK(clk), .RST(rst), .Q(sreg[1591]) );
  DFF \sreg_reg[1590]  ( .D(c[1594]), .CLK(clk), .RST(rst), .Q(sreg[1590]) );
  DFF \sreg_reg[1589]  ( .D(c[1593]), .CLK(clk), .RST(rst), .Q(sreg[1589]) );
  DFF \sreg_reg[1588]  ( .D(c[1592]), .CLK(clk), .RST(rst), .Q(sreg[1588]) );
  DFF \sreg_reg[1587]  ( .D(c[1591]), .CLK(clk), .RST(rst), .Q(sreg[1587]) );
  DFF \sreg_reg[1586]  ( .D(c[1590]), .CLK(clk), .RST(rst), .Q(sreg[1586]) );
  DFF \sreg_reg[1585]  ( .D(c[1589]), .CLK(clk), .RST(rst), .Q(sreg[1585]) );
  DFF \sreg_reg[1584]  ( .D(c[1588]), .CLK(clk), .RST(rst), .Q(sreg[1584]) );
  DFF \sreg_reg[1583]  ( .D(c[1587]), .CLK(clk), .RST(rst), .Q(sreg[1583]) );
  DFF \sreg_reg[1582]  ( .D(c[1586]), .CLK(clk), .RST(rst), .Q(sreg[1582]) );
  DFF \sreg_reg[1581]  ( .D(c[1585]), .CLK(clk), .RST(rst), .Q(sreg[1581]) );
  DFF \sreg_reg[1580]  ( .D(c[1584]), .CLK(clk), .RST(rst), .Q(sreg[1580]) );
  DFF \sreg_reg[1579]  ( .D(c[1583]), .CLK(clk), .RST(rst), .Q(sreg[1579]) );
  DFF \sreg_reg[1578]  ( .D(c[1582]), .CLK(clk), .RST(rst), .Q(sreg[1578]) );
  DFF \sreg_reg[1577]  ( .D(c[1581]), .CLK(clk), .RST(rst), .Q(sreg[1577]) );
  DFF \sreg_reg[1576]  ( .D(c[1580]), .CLK(clk), .RST(rst), .Q(sreg[1576]) );
  DFF \sreg_reg[1575]  ( .D(c[1579]), .CLK(clk), .RST(rst), .Q(sreg[1575]) );
  DFF \sreg_reg[1574]  ( .D(c[1578]), .CLK(clk), .RST(rst), .Q(sreg[1574]) );
  DFF \sreg_reg[1573]  ( .D(c[1577]), .CLK(clk), .RST(rst), .Q(sreg[1573]) );
  DFF \sreg_reg[1572]  ( .D(c[1576]), .CLK(clk), .RST(rst), .Q(sreg[1572]) );
  DFF \sreg_reg[1571]  ( .D(c[1575]), .CLK(clk), .RST(rst), .Q(sreg[1571]) );
  DFF \sreg_reg[1570]  ( .D(c[1574]), .CLK(clk), .RST(rst), .Q(sreg[1570]) );
  DFF \sreg_reg[1569]  ( .D(c[1573]), .CLK(clk), .RST(rst), .Q(sreg[1569]) );
  DFF \sreg_reg[1568]  ( .D(c[1572]), .CLK(clk), .RST(rst), .Q(sreg[1568]) );
  DFF \sreg_reg[1567]  ( .D(c[1571]), .CLK(clk), .RST(rst), .Q(sreg[1567]) );
  DFF \sreg_reg[1566]  ( .D(c[1570]), .CLK(clk), .RST(rst), .Q(sreg[1566]) );
  DFF \sreg_reg[1565]  ( .D(c[1569]), .CLK(clk), .RST(rst), .Q(sreg[1565]) );
  DFF \sreg_reg[1564]  ( .D(c[1568]), .CLK(clk), .RST(rst), .Q(sreg[1564]) );
  DFF \sreg_reg[1563]  ( .D(c[1567]), .CLK(clk), .RST(rst), .Q(sreg[1563]) );
  DFF \sreg_reg[1562]  ( .D(c[1566]), .CLK(clk), .RST(rst), .Q(sreg[1562]) );
  DFF \sreg_reg[1561]  ( .D(c[1565]), .CLK(clk), .RST(rst), .Q(sreg[1561]) );
  DFF \sreg_reg[1560]  ( .D(c[1564]), .CLK(clk), .RST(rst), .Q(sreg[1560]) );
  DFF \sreg_reg[1559]  ( .D(c[1563]), .CLK(clk), .RST(rst), .Q(sreg[1559]) );
  DFF \sreg_reg[1558]  ( .D(c[1562]), .CLK(clk), .RST(rst), .Q(sreg[1558]) );
  DFF \sreg_reg[1557]  ( .D(c[1561]), .CLK(clk), .RST(rst), .Q(sreg[1557]) );
  DFF \sreg_reg[1556]  ( .D(c[1560]), .CLK(clk), .RST(rst), .Q(sreg[1556]) );
  DFF \sreg_reg[1555]  ( .D(c[1559]), .CLK(clk), .RST(rst), .Q(sreg[1555]) );
  DFF \sreg_reg[1554]  ( .D(c[1558]), .CLK(clk), .RST(rst), .Q(sreg[1554]) );
  DFF \sreg_reg[1553]  ( .D(c[1557]), .CLK(clk), .RST(rst), .Q(sreg[1553]) );
  DFF \sreg_reg[1552]  ( .D(c[1556]), .CLK(clk), .RST(rst), .Q(sreg[1552]) );
  DFF \sreg_reg[1551]  ( .D(c[1555]), .CLK(clk), .RST(rst), .Q(sreg[1551]) );
  DFF \sreg_reg[1550]  ( .D(c[1554]), .CLK(clk), .RST(rst), .Q(sreg[1550]) );
  DFF \sreg_reg[1549]  ( .D(c[1553]), .CLK(clk), .RST(rst), .Q(sreg[1549]) );
  DFF \sreg_reg[1548]  ( .D(c[1552]), .CLK(clk), .RST(rst), .Q(sreg[1548]) );
  DFF \sreg_reg[1547]  ( .D(c[1551]), .CLK(clk), .RST(rst), .Q(sreg[1547]) );
  DFF \sreg_reg[1546]  ( .D(c[1550]), .CLK(clk), .RST(rst), .Q(sreg[1546]) );
  DFF \sreg_reg[1545]  ( .D(c[1549]), .CLK(clk), .RST(rst), .Q(sreg[1545]) );
  DFF \sreg_reg[1544]  ( .D(c[1548]), .CLK(clk), .RST(rst), .Q(sreg[1544]) );
  DFF \sreg_reg[1543]  ( .D(c[1547]), .CLK(clk), .RST(rst), .Q(sreg[1543]) );
  DFF \sreg_reg[1542]  ( .D(c[1546]), .CLK(clk), .RST(rst), .Q(sreg[1542]) );
  DFF \sreg_reg[1541]  ( .D(c[1545]), .CLK(clk), .RST(rst), .Q(sreg[1541]) );
  DFF \sreg_reg[1540]  ( .D(c[1544]), .CLK(clk), .RST(rst), .Q(sreg[1540]) );
  DFF \sreg_reg[1539]  ( .D(c[1543]), .CLK(clk), .RST(rst), .Q(sreg[1539]) );
  DFF \sreg_reg[1538]  ( .D(c[1542]), .CLK(clk), .RST(rst), .Q(sreg[1538]) );
  DFF \sreg_reg[1537]  ( .D(c[1541]), .CLK(clk), .RST(rst), .Q(sreg[1537]) );
  DFF \sreg_reg[1536]  ( .D(c[1540]), .CLK(clk), .RST(rst), .Q(sreg[1536]) );
  DFF \sreg_reg[1535]  ( .D(c[1539]), .CLK(clk), .RST(rst), .Q(sreg[1535]) );
  DFF \sreg_reg[1534]  ( .D(c[1538]), .CLK(clk), .RST(rst), .Q(sreg[1534]) );
  DFF \sreg_reg[1533]  ( .D(c[1537]), .CLK(clk), .RST(rst), .Q(sreg[1533]) );
  DFF \sreg_reg[1532]  ( .D(c[1536]), .CLK(clk), .RST(rst), .Q(sreg[1532]) );
  DFF \sreg_reg[1531]  ( .D(c[1535]), .CLK(clk), .RST(rst), .Q(sreg[1531]) );
  DFF \sreg_reg[1530]  ( .D(c[1534]), .CLK(clk), .RST(rst), .Q(sreg[1530]) );
  DFF \sreg_reg[1529]  ( .D(c[1533]), .CLK(clk), .RST(rst), .Q(sreg[1529]) );
  DFF \sreg_reg[1528]  ( .D(c[1532]), .CLK(clk), .RST(rst), .Q(sreg[1528]) );
  DFF \sreg_reg[1527]  ( .D(c[1531]), .CLK(clk), .RST(rst), .Q(sreg[1527]) );
  DFF \sreg_reg[1526]  ( .D(c[1530]), .CLK(clk), .RST(rst), .Q(sreg[1526]) );
  DFF \sreg_reg[1525]  ( .D(c[1529]), .CLK(clk), .RST(rst), .Q(sreg[1525]) );
  DFF \sreg_reg[1524]  ( .D(c[1528]), .CLK(clk), .RST(rst), .Q(sreg[1524]) );
  DFF \sreg_reg[1523]  ( .D(c[1527]), .CLK(clk), .RST(rst), .Q(sreg[1523]) );
  DFF \sreg_reg[1522]  ( .D(c[1526]), .CLK(clk), .RST(rst), .Q(sreg[1522]) );
  DFF \sreg_reg[1521]  ( .D(c[1525]), .CLK(clk), .RST(rst), .Q(sreg[1521]) );
  DFF \sreg_reg[1520]  ( .D(c[1524]), .CLK(clk), .RST(rst), .Q(sreg[1520]) );
  DFF \sreg_reg[1519]  ( .D(c[1523]), .CLK(clk), .RST(rst), .Q(sreg[1519]) );
  DFF \sreg_reg[1518]  ( .D(c[1522]), .CLK(clk), .RST(rst), .Q(sreg[1518]) );
  DFF \sreg_reg[1517]  ( .D(c[1521]), .CLK(clk), .RST(rst), .Q(sreg[1517]) );
  DFF \sreg_reg[1516]  ( .D(c[1520]), .CLK(clk), .RST(rst), .Q(sreg[1516]) );
  DFF \sreg_reg[1515]  ( .D(c[1519]), .CLK(clk), .RST(rst), .Q(sreg[1515]) );
  DFF \sreg_reg[1514]  ( .D(c[1518]), .CLK(clk), .RST(rst), .Q(sreg[1514]) );
  DFF \sreg_reg[1513]  ( .D(c[1517]), .CLK(clk), .RST(rst), .Q(sreg[1513]) );
  DFF \sreg_reg[1512]  ( .D(c[1516]), .CLK(clk), .RST(rst), .Q(sreg[1512]) );
  DFF \sreg_reg[1511]  ( .D(c[1515]), .CLK(clk), .RST(rst), .Q(sreg[1511]) );
  DFF \sreg_reg[1510]  ( .D(c[1514]), .CLK(clk), .RST(rst), .Q(sreg[1510]) );
  DFF \sreg_reg[1509]  ( .D(c[1513]), .CLK(clk), .RST(rst), .Q(sreg[1509]) );
  DFF \sreg_reg[1508]  ( .D(c[1512]), .CLK(clk), .RST(rst), .Q(sreg[1508]) );
  DFF \sreg_reg[1507]  ( .D(c[1511]), .CLK(clk), .RST(rst), .Q(sreg[1507]) );
  DFF \sreg_reg[1506]  ( .D(c[1510]), .CLK(clk), .RST(rst), .Q(sreg[1506]) );
  DFF \sreg_reg[1505]  ( .D(c[1509]), .CLK(clk), .RST(rst), .Q(sreg[1505]) );
  DFF \sreg_reg[1504]  ( .D(c[1508]), .CLK(clk), .RST(rst), .Q(sreg[1504]) );
  DFF \sreg_reg[1503]  ( .D(c[1507]), .CLK(clk), .RST(rst), .Q(sreg[1503]) );
  DFF \sreg_reg[1502]  ( .D(c[1506]), .CLK(clk), .RST(rst), .Q(sreg[1502]) );
  DFF \sreg_reg[1501]  ( .D(c[1505]), .CLK(clk), .RST(rst), .Q(sreg[1501]) );
  DFF \sreg_reg[1500]  ( .D(c[1504]), .CLK(clk), .RST(rst), .Q(sreg[1500]) );
  DFF \sreg_reg[1499]  ( .D(c[1503]), .CLK(clk), .RST(rst), .Q(sreg[1499]) );
  DFF \sreg_reg[1498]  ( .D(c[1502]), .CLK(clk), .RST(rst), .Q(sreg[1498]) );
  DFF \sreg_reg[1497]  ( .D(c[1501]), .CLK(clk), .RST(rst), .Q(sreg[1497]) );
  DFF \sreg_reg[1496]  ( .D(c[1500]), .CLK(clk), .RST(rst), .Q(sreg[1496]) );
  DFF \sreg_reg[1495]  ( .D(c[1499]), .CLK(clk), .RST(rst), .Q(sreg[1495]) );
  DFF \sreg_reg[1494]  ( .D(c[1498]), .CLK(clk), .RST(rst), .Q(sreg[1494]) );
  DFF \sreg_reg[1493]  ( .D(c[1497]), .CLK(clk), .RST(rst), .Q(sreg[1493]) );
  DFF \sreg_reg[1492]  ( .D(c[1496]), .CLK(clk), .RST(rst), .Q(sreg[1492]) );
  DFF \sreg_reg[1491]  ( .D(c[1495]), .CLK(clk), .RST(rst), .Q(sreg[1491]) );
  DFF \sreg_reg[1490]  ( .D(c[1494]), .CLK(clk), .RST(rst), .Q(sreg[1490]) );
  DFF \sreg_reg[1489]  ( .D(c[1493]), .CLK(clk), .RST(rst), .Q(sreg[1489]) );
  DFF \sreg_reg[1488]  ( .D(c[1492]), .CLK(clk), .RST(rst), .Q(sreg[1488]) );
  DFF \sreg_reg[1487]  ( .D(c[1491]), .CLK(clk), .RST(rst), .Q(sreg[1487]) );
  DFF \sreg_reg[1486]  ( .D(c[1490]), .CLK(clk), .RST(rst), .Q(sreg[1486]) );
  DFF \sreg_reg[1485]  ( .D(c[1489]), .CLK(clk), .RST(rst), .Q(sreg[1485]) );
  DFF \sreg_reg[1484]  ( .D(c[1488]), .CLK(clk), .RST(rst), .Q(sreg[1484]) );
  DFF \sreg_reg[1483]  ( .D(c[1487]), .CLK(clk), .RST(rst), .Q(sreg[1483]) );
  DFF \sreg_reg[1482]  ( .D(c[1486]), .CLK(clk), .RST(rst), .Q(sreg[1482]) );
  DFF \sreg_reg[1481]  ( .D(c[1485]), .CLK(clk), .RST(rst), .Q(sreg[1481]) );
  DFF \sreg_reg[1480]  ( .D(c[1484]), .CLK(clk), .RST(rst), .Q(sreg[1480]) );
  DFF \sreg_reg[1479]  ( .D(c[1483]), .CLK(clk), .RST(rst), .Q(sreg[1479]) );
  DFF \sreg_reg[1478]  ( .D(c[1482]), .CLK(clk), .RST(rst), .Q(sreg[1478]) );
  DFF \sreg_reg[1477]  ( .D(c[1481]), .CLK(clk), .RST(rst), .Q(sreg[1477]) );
  DFF \sreg_reg[1476]  ( .D(c[1480]), .CLK(clk), .RST(rst), .Q(sreg[1476]) );
  DFF \sreg_reg[1475]  ( .D(c[1479]), .CLK(clk), .RST(rst), .Q(sreg[1475]) );
  DFF \sreg_reg[1474]  ( .D(c[1478]), .CLK(clk), .RST(rst), .Q(sreg[1474]) );
  DFF \sreg_reg[1473]  ( .D(c[1477]), .CLK(clk), .RST(rst), .Q(sreg[1473]) );
  DFF \sreg_reg[1472]  ( .D(c[1476]), .CLK(clk), .RST(rst), .Q(sreg[1472]) );
  DFF \sreg_reg[1471]  ( .D(c[1475]), .CLK(clk), .RST(rst), .Q(sreg[1471]) );
  DFF \sreg_reg[1470]  ( .D(c[1474]), .CLK(clk), .RST(rst), .Q(sreg[1470]) );
  DFF \sreg_reg[1469]  ( .D(c[1473]), .CLK(clk), .RST(rst), .Q(sreg[1469]) );
  DFF \sreg_reg[1468]  ( .D(c[1472]), .CLK(clk), .RST(rst), .Q(sreg[1468]) );
  DFF \sreg_reg[1467]  ( .D(c[1471]), .CLK(clk), .RST(rst), .Q(sreg[1467]) );
  DFF \sreg_reg[1466]  ( .D(c[1470]), .CLK(clk), .RST(rst), .Q(sreg[1466]) );
  DFF \sreg_reg[1465]  ( .D(c[1469]), .CLK(clk), .RST(rst), .Q(sreg[1465]) );
  DFF \sreg_reg[1464]  ( .D(c[1468]), .CLK(clk), .RST(rst), .Q(sreg[1464]) );
  DFF \sreg_reg[1463]  ( .D(c[1467]), .CLK(clk), .RST(rst), .Q(sreg[1463]) );
  DFF \sreg_reg[1462]  ( .D(c[1466]), .CLK(clk), .RST(rst), .Q(sreg[1462]) );
  DFF \sreg_reg[1461]  ( .D(c[1465]), .CLK(clk), .RST(rst), .Q(sreg[1461]) );
  DFF \sreg_reg[1460]  ( .D(c[1464]), .CLK(clk), .RST(rst), .Q(sreg[1460]) );
  DFF \sreg_reg[1459]  ( .D(c[1463]), .CLK(clk), .RST(rst), .Q(sreg[1459]) );
  DFF \sreg_reg[1458]  ( .D(c[1462]), .CLK(clk), .RST(rst), .Q(sreg[1458]) );
  DFF \sreg_reg[1457]  ( .D(c[1461]), .CLK(clk), .RST(rst), .Q(sreg[1457]) );
  DFF \sreg_reg[1456]  ( .D(c[1460]), .CLK(clk), .RST(rst), .Q(sreg[1456]) );
  DFF \sreg_reg[1455]  ( .D(c[1459]), .CLK(clk), .RST(rst), .Q(sreg[1455]) );
  DFF \sreg_reg[1454]  ( .D(c[1458]), .CLK(clk), .RST(rst), .Q(sreg[1454]) );
  DFF \sreg_reg[1453]  ( .D(c[1457]), .CLK(clk), .RST(rst), .Q(sreg[1453]) );
  DFF \sreg_reg[1452]  ( .D(c[1456]), .CLK(clk), .RST(rst), .Q(sreg[1452]) );
  DFF \sreg_reg[1451]  ( .D(c[1455]), .CLK(clk), .RST(rst), .Q(sreg[1451]) );
  DFF \sreg_reg[1450]  ( .D(c[1454]), .CLK(clk), .RST(rst), .Q(sreg[1450]) );
  DFF \sreg_reg[1449]  ( .D(c[1453]), .CLK(clk), .RST(rst), .Q(sreg[1449]) );
  DFF \sreg_reg[1448]  ( .D(c[1452]), .CLK(clk), .RST(rst), .Q(sreg[1448]) );
  DFF \sreg_reg[1447]  ( .D(c[1451]), .CLK(clk), .RST(rst), .Q(sreg[1447]) );
  DFF \sreg_reg[1446]  ( .D(c[1450]), .CLK(clk), .RST(rst), .Q(sreg[1446]) );
  DFF \sreg_reg[1445]  ( .D(c[1449]), .CLK(clk), .RST(rst), .Q(sreg[1445]) );
  DFF \sreg_reg[1444]  ( .D(c[1448]), .CLK(clk), .RST(rst), .Q(sreg[1444]) );
  DFF \sreg_reg[1443]  ( .D(c[1447]), .CLK(clk), .RST(rst), .Q(sreg[1443]) );
  DFF \sreg_reg[1442]  ( .D(c[1446]), .CLK(clk), .RST(rst), .Q(sreg[1442]) );
  DFF \sreg_reg[1441]  ( .D(c[1445]), .CLK(clk), .RST(rst), .Q(sreg[1441]) );
  DFF \sreg_reg[1440]  ( .D(c[1444]), .CLK(clk), .RST(rst), .Q(sreg[1440]) );
  DFF \sreg_reg[1439]  ( .D(c[1443]), .CLK(clk), .RST(rst), .Q(sreg[1439]) );
  DFF \sreg_reg[1438]  ( .D(c[1442]), .CLK(clk), .RST(rst), .Q(sreg[1438]) );
  DFF \sreg_reg[1437]  ( .D(c[1441]), .CLK(clk), .RST(rst), .Q(sreg[1437]) );
  DFF \sreg_reg[1436]  ( .D(c[1440]), .CLK(clk), .RST(rst), .Q(sreg[1436]) );
  DFF \sreg_reg[1435]  ( .D(c[1439]), .CLK(clk), .RST(rst), .Q(sreg[1435]) );
  DFF \sreg_reg[1434]  ( .D(c[1438]), .CLK(clk), .RST(rst), .Q(sreg[1434]) );
  DFF \sreg_reg[1433]  ( .D(c[1437]), .CLK(clk), .RST(rst), .Q(sreg[1433]) );
  DFF \sreg_reg[1432]  ( .D(c[1436]), .CLK(clk), .RST(rst), .Q(sreg[1432]) );
  DFF \sreg_reg[1431]  ( .D(c[1435]), .CLK(clk), .RST(rst), .Q(sreg[1431]) );
  DFF \sreg_reg[1430]  ( .D(c[1434]), .CLK(clk), .RST(rst), .Q(sreg[1430]) );
  DFF \sreg_reg[1429]  ( .D(c[1433]), .CLK(clk), .RST(rst), .Q(sreg[1429]) );
  DFF \sreg_reg[1428]  ( .D(c[1432]), .CLK(clk), .RST(rst), .Q(sreg[1428]) );
  DFF \sreg_reg[1427]  ( .D(c[1431]), .CLK(clk), .RST(rst), .Q(sreg[1427]) );
  DFF \sreg_reg[1426]  ( .D(c[1430]), .CLK(clk), .RST(rst), .Q(sreg[1426]) );
  DFF \sreg_reg[1425]  ( .D(c[1429]), .CLK(clk), .RST(rst), .Q(sreg[1425]) );
  DFF \sreg_reg[1424]  ( .D(c[1428]), .CLK(clk), .RST(rst), .Q(sreg[1424]) );
  DFF \sreg_reg[1423]  ( .D(c[1427]), .CLK(clk), .RST(rst), .Q(sreg[1423]) );
  DFF \sreg_reg[1422]  ( .D(c[1426]), .CLK(clk), .RST(rst), .Q(sreg[1422]) );
  DFF \sreg_reg[1421]  ( .D(c[1425]), .CLK(clk), .RST(rst), .Q(sreg[1421]) );
  DFF \sreg_reg[1420]  ( .D(c[1424]), .CLK(clk), .RST(rst), .Q(sreg[1420]) );
  DFF \sreg_reg[1419]  ( .D(c[1423]), .CLK(clk), .RST(rst), .Q(sreg[1419]) );
  DFF \sreg_reg[1418]  ( .D(c[1422]), .CLK(clk), .RST(rst), .Q(sreg[1418]) );
  DFF \sreg_reg[1417]  ( .D(c[1421]), .CLK(clk), .RST(rst), .Q(sreg[1417]) );
  DFF \sreg_reg[1416]  ( .D(c[1420]), .CLK(clk), .RST(rst), .Q(sreg[1416]) );
  DFF \sreg_reg[1415]  ( .D(c[1419]), .CLK(clk), .RST(rst), .Q(sreg[1415]) );
  DFF \sreg_reg[1414]  ( .D(c[1418]), .CLK(clk), .RST(rst), .Q(sreg[1414]) );
  DFF \sreg_reg[1413]  ( .D(c[1417]), .CLK(clk), .RST(rst), .Q(sreg[1413]) );
  DFF \sreg_reg[1412]  ( .D(c[1416]), .CLK(clk), .RST(rst), .Q(sreg[1412]) );
  DFF \sreg_reg[1411]  ( .D(c[1415]), .CLK(clk), .RST(rst), .Q(sreg[1411]) );
  DFF \sreg_reg[1410]  ( .D(c[1414]), .CLK(clk), .RST(rst), .Q(sreg[1410]) );
  DFF \sreg_reg[1409]  ( .D(c[1413]), .CLK(clk), .RST(rst), .Q(sreg[1409]) );
  DFF \sreg_reg[1408]  ( .D(c[1412]), .CLK(clk), .RST(rst), .Q(sreg[1408]) );
  DFF \sreg_reg[1407]  ( .D(c[1411]), .CLK(clk), .RST(rst), .Q(sreg[1407]) );
  DFF \sreg_reg[1406]  ( .D(c[1410]), .CLK(clk), .RST(rst), .Q(sreg[1406]) );
  DFF \sreg_reg[1405]  ( .D(c[1409]), .CLK(clk), .RST(rst), .Q(sreg[1405]) );
  DFF \sreg_reg[1404]  ( .D(c[1408]), .CLK(clk), .RST(rst), .Q(sreg[1404]) );
  DFF \sreg_reg[1403]  ( .D(c[1407]), .CLK(clk), .RST(rst), .Q(sreg[1403]) );
  DFF \sreg_reg[1402]  ( .D(c[1406]), .CLK(clk), .RST(rst), .Q(sreg[1402]) );
  DFF \sreg_reg[1401]  ( .D(c[1405]), .CLK(clk), .RST(rst), .Q(sreg[1401]) );
  DFF \sreg_reg[1400]  ( .D(c[1404]), .CLK(clk), .RST(rst), .Q(sreg[1400]) );
  DFF \sreg_reg[1399]  ( .D(c[1403]), .CLK(clk), .RST(rst), .Q(sreg[1399]) );
  DFF \sreg_reg[1398]  ( .D(c[1402]), .CLK(clk), .RST(rst), .Q(sreg[1398]) );
  DFF \sreg_reg[1397]  ( .D(c[1401]), .CLK(clk), .RST(rst), .Q(sreg[1397]) );
  DFF \sreg_reg[1396]  ( .D(c[1400]), .CLK(clk), .RST(rst), .Q(sreg[1396]) );
  DFF \sreg_reg[1395]  ( .D(c[1399]), .CLK(clk), .RST(rst), .Q(sreg[1395]) );
  DFF \sreg_reg[1394]  ( .D(c[1398]), .CLK(clk), .RST(rst), .Q(sreg[1394]) );
  DFF \sreg_reg[1393]  ( .D(c[1397]), .CLK(clk), .RST(rst), .Q(sreg[1393]) );
  DFF \sreg_reg[1392]  ( .D(c[1396]), .CLK(clk), .RST(rst), .Q(sreg[1392]) );
  DFF \sreg_reg[1391]  ( .D(c[1395]), .CLK(clk), .RST(rst), .Q(sreg[1391]) );
  DFF \sreg_reg[1390]  ( .D(c[1394]), .CLK(clk), .RST(rst), .Q(sreg[1390]) );
  DFF \sreg_reg[1389]  ( .D(c[1393]), .CLK(clk), .RST(rst), .Q(sreg[1389]) );
  DFF \sreg_reg[1388]  ( .D(c[1392]), .CLK(clk), .RST(rst), .Q(sreg[1388]) );
  DFF \sreg_reg[1387]  ( .D(c[1391]), .CLK(clk), .RST(rst), .Q(sreg[1387]) );
  DFF \sreg_reg[1386]  ( .D(c[1390]), .CLK(clk), .RST(rst), .Q(sreg[1386]) );
  DFF \sreg_reg[1385]  ( .D(c[1389]), .CLK(clk), .RST(rst), .Q(sreg[1385]) );
  DFF \sreg_reg[1384]  ( .D(c[1388]), .CLK(clk), .RST(rst), .Q(sreg[1384]) );
  DFF \sreg_reg[1383]  ( .D(c[1387]), .CLK(clk), .RST(rst), .Q(sreg[1383]) );
  DFF \sreg_reg[1382]  ( .D(c[1386]), .CLK(clk), .RST(rst), .Q(sreg[1382]) );
  DFF \sreg_reg[1381]  ( .D(c[1385]), .CLK(clk), .RST(rst), .Q(sreg[1381]) );
  DFF \sreg_reg[1380]  ( .D(c[1384]), .CLK(clk), .RST(rst), .Q(sreg[1380]) );
  DFF \sreg_reg[1379]  ( .D(c[1383]), .CLK(clk), .RST(rst), .Q(sreg[1379]) );
  DFF \sreg_reg[1378]  ( .D(c[1382]), .CLK(clk), .RST(rst), .Q(sreg[1378]) );
  DFF \sreg_reg[1377]  ( .D(c[1381]), .CLK(clk), .RST(rst), .Q(sreg[1377]) );
  DFF \sreg_reg[1376]  ( .D(c[1380]), .CLK(clk), .RST(rst), .Q(sreg[1376]) );
  DFF \sreg_reg[1375]  ( .D(c[1379]), .CLK(clk), .RST(rst), .Q(sreg[1375]) );
  DFF \sreg_reg[1374]  ( .D(c[1378]), .CLK(clk), .RST(rst), .Q(sreg[1374]) );
  DFF \sreg_reg[1373]  ( .D(c[1377]), .CLK(clk), .RST(rst), .Q(sreg[1373]) );
  DFF \sreg_reg[1372]  ( .D(c[1376]), .CLK(clk), .RST(rst), .Q(sreg[1372]) );
  DFF \sreg_reg[1371]  ( .D(c[1375]), .CLK(clk), .RST(rst), .Q(sreg[1371]) );
  DFF \sreg_reg[1370]  ( .D(c[1374]), .CLK(clk), .RST(rst), .Q(sreg[1370]) );
  DFF \sreg_reg[1369]  ( .D(c[1373]), .CLK(clk), .RST(rst), .Q(sreg[1369]) );
  DFF \sreg_reg[1368]  ( .D(c[1372]), .CLK(clk), .RST(rst), .Q(sreg[1368]) );
  DFF \sreg_reg[1367]  ( .D(c[1371]), .CLK(clk), .RST(rst), .Q(sreg[1367]) );
  DFF \sreg_reg[1366]  ( .D(c[1370]), .CLK(clk), .RST(rst), .Q(sreg[1366]) );
  DFF \sreg_reg[1365]  ( .D(c[1369]), .CLK(clk), .RST(rst), .Q(sreg[1365]) );
  DFF \sreg_reg[1364]  ( .D(c[1368]), .CLK(clk), .RST(rst), .Q(sreg[1364]) );
  DFF \sreg_reg[1363]  ( .D(c[1367]), .CLK(clk), .RST(rst), .Q(sreg[1363]) );
  DFF \sreg_reg[1362]  ( .D(c[1366]), .CLK(clk), .RST(rst), .Q(sreg[1362]) );
  DFF \sreg_reg[1361]  ( .D(c[1365]), .CLK(clk), .RST(rst), .Q(sreg[1361]) );
  DFF \sreg_reg[1360]  ( .D(c[1364]), .CLK(clk), .RST(rst), .Q(sreg[1360]) );
  DFF \sreg_reg[1359]  ( .D(c[1363]), .CLK(clk), .RST(rst), .Q(sreg[1359]) );
  DFF \sreg_reg[1358]  ( .D(c[1362]), .CLK(clk), .RST(rst), .Q(sreg[1358]) );
  DFF \sreg_reg[1357]  ( .D(c[1361]), .CLK(clk), .RST(rst), .Q(sreg[1357]) );
  DFF \sreg_reg[1356]  ( .D(c[1360]), .CLK(clk), .RST(rst), .Q(sreg[1356]) );
  DFF \sreg_reg[1355]  ( .D(c[1359]), .CLK(clk), .RST(rst), .Q(sreg[1355]) );
  DFF \sreg_reg[1354]  ( .D(c[1358]), .CLK(clk), .RST(rst), .Q(sreg[1354]) );
  DFF \sreg_reg[1353]  ( .D(c[1357]), .CLK(clk), .RST(rst), .Q(sreg[1353]) );
  DFF \sreg_reg[1352]  ( .D(c[1356]), .CLK(clk), .RST(rst), .Q(sreg[1352]) );
  DFF \sreg_reg[1351]  ( .D(c[1355]), .CLK(clk), .RST(rst), .Q(sreg[1351]) );
  DFF \sreg_reg[1350]  ( .D(c[1354]), .CLK(clk), .RST(rst), .Q(sreg[1350]) );
  DFF \sreg_reg[1349]  ( .D(c[1353]), .CLK(clk), .RST(rst), .Q(sreg[1349]) );
  DFF \sreg_reg[1348]  ( .D(c[1352]), .CLK(clk), .RST(rst), .Q(sreg[1348]) );
  DFF \sreg_reg[1347]  ( .D(c[1351]), .CLK(clk), .RST(rst), .Q(sreg[1347]) );
  DFF \sreg_reg[1346]  ( .D(c[1350]), .CLK(clk), .RST(rst), .Q(sreg[1346]) );
  DFF \sreg_reg[1345]  ( .D(c[1349]), .CLK(clk), .RST(rst), .Q(sreg[1345]) );
  DFF \sreg_reg[1344]  ( .D(c[1348]), .CLK(clk), .RST(rst), .Q(sreg[1344]) );
  DFF \sreg_reg[1343]  ( .D(c[1347]), .CLK(clk), .RST(rst), .Q(sreg[1343]) );
  DFF \sreg_reg[1342]  ( .D(c[1346]), .CLK(clk), .RST(rst), .Q(sreg[1342]) );
  DFF \sreg_reg[1341]  ( .D(c[1345]), .CLK(clk), .RST(rst), .Q(sreg[1341]) );
  DFF \sreg_reg[1340]  ( .D(c[1344]), .CLK(clk), .RST(rst), .Q(sreg[1340]) );
  DFF \sreg_reg[1339]  ( .D(c[1343]), .CLK(clk), .RST(rst), .Q(sreg[1339]) );
  DFF \sreg_reg[1338]  ( .D(c[1342]), .CLK(clk), .RST(rst), .Q(sreg[1338]) );
  DFF \sreg_reg[1337]  ( .D(c[1341]), .CLK(clk), .RST(rst), .Q(sreg[1337]) );
  DFF \sreg_reg[1336]  ( .D(c[1340]), .CLK(clk), .RST(rst), .Q(sreg[1336]) );
  DFF \sreg_reg[1335]  ( .D(c[1339]), .CLK(clk), .RST(rst), .Q(sreg[1335]) );
  DFF \sreg_reg[1334]  ( .D(c[1338]), .CLK(clk), .RST(rst), .Q(sreg[1334]) );
  DFF \sreg_reg[1333]  ( .D(c[1337]), .CLK(clk), .RST(rst), .Q(sreg[1333]) );
  DFF \sreg_reg[1332]  ( .D(c[1336]), .CLK(clk), .RST(rst), .Q(sreg[1332]) );
  DFF \sreg_reg[1331]  ( .D(c[1335]), .CLK(clk), .RST(rst), .Q(sreg[1331]) );
  DFF \sreg_reg[1330]  ( .D(c[1334]), .CLK(clk), .RST(rst), .Q(sreg[1330]) );
  DFF \sreg_reg[1329]  ( .D(c[1333]), .CLK(clk), .RST(rst), .Q(sreg[1329]) );
  DFF \sreg_reg[1328]  ( .D(c[1332]), .CLK(clk), .RST(rst), .Q(sreg[1328]) );
  DFF \sreg_reg[1327]  ( .D(c[1331]), .CLK(clk), .RST(rst), .Q(sreg[1327]) );
  DFF \sreg_reg[1326]  ( .D(c[1330]), .CLK(clk), .RST(rst), .Q(sreg[1326]) );
  DFF \sreg_reg[1325]  ( .D(c[1329]), .CLK(clk), .RST(rst), .Q(sreg[1325]) );
  DFF \sreg_reg[1324]  ( .D(c[1328]), .CLK(clk), .RST(rst), .Q(sreg[1324]) );
  DFF \sreg_reg[1323]  ( .D(c[1327]), .CLK(clk), .RST(rst), .Q(sreg[1323]) );
  DFF \sreg_reg[1322]  ( .D(c[1326]), .CLK(clk), .RST(rst), .Q(sreg[1322]) );
  DFF \sreg_reg[1321]  ( .D(c[1325]), .CLK(clk), .RST(rst), .Q(sreg[1321]) );
  DFF \sreg_reg[1320]  ( .D(c[1324]), .CLK(clk), .RST(rst), .Q(sreg[1320]) );
  DFF \sreg_reg[1319]  ( .D(c[1323]), .CLK(clk), .RST(rst), .Q(sreg[1319]) );
  DFF \sreg_reg[1318]  ( .D(c[1322]), .CLK(clk), .RST(rst), .Q(sreg[1318]) );
  DFF \sreg_reg[1317]  ( .D(c[1321]), .CLK(clk), .RST(rst), .Q(sreg[1317]) );
  DFF \sreg_reg[1316]  ( .D(c[1320]), .CLK(clk), .RST(rst), .Q(sreg[1316]) );
  DFF \sreg_reg[1315]  ( .D(c[1319]), .CLK(clk), .RST(rst), .Q(sreg[1315]) );
  DFF \sreg_reg[1314]  ( .D(c[1318]), .CLK(clk), .RST(rst), .Q(sreg[1314]) );
  DFF \sreg_reg[1313]  ( .D(c[1317]), .CLK(clk), .RST(rst), .Q(sreg[1313]) );
  DFF \sreg_reg[1312]  ( .D(c[1316]), .CLK(clk), .RST(rst), .Q(sreg[1312]) );
  DFF \sreg_reg[1311]  ( .D(c[1315]), .CLK(clk), .RST(rst), .Q(sreg[1311]) );
  DFF \sreg_reg[1310]  ( .D(c[1314]), .CLK(clk), .RST(rst), .Q(sreg[1310]) );
  DFF \sreg_reg[1309]  ( .D(c[1313]), .CLK(clk), .RST(rst), .Q(sreg[1309]) );
  DFF \sreg_reg[1308]  ( .D(c[1312]), .CLK(clk), .RST(rst), .Q(sreg[1308]) );
  DFF \sreg_reg[1307]  ( .D(c[1311]), .CLK(clk), .RST(rst), .Q(sreg[1307]) );
  DFF \sreg_reg[1306]  ( .D(c[1310]), .CLK(clk), .RST(rst), .Q(sreg[1306]) );
  DFF \sreg_reg[1305]  ( .D(c[1309]), .CLK(clk), .RST(rst), .Q(sreg[1305]) );
  DFF \sreg_reg[1304]  ( .D(c[1308]), .CLK(clk), .RST(rst), .Q(sreg[1304]) );
  DFF \sreg_reg[1303]  ( .D(c[1307]), .CLK(clk), .RST(rst), .Q(sreg[1303]) );
  DFF \sreg_reg[1302]  ( .D(c[1306]), .CLK(clk), .RST(rst), .Q(sreg[1302]) );
  DFF \sreg_reg[1301]  ( .D(c[1305]), .CLK(clk), .RST(rst), .Q(sreg[1301]) );
  DFF \sreg_reg[1300]  ( .D(c[1304]), .CLK(clk), .RST(rst), .Q(sreg[1300]) );
  DFF \sreg_reg[1299]  ( .D(c[1303]), .CLK(clk), .RST(rst), .Q(sreg[1299]) );
  DFF \sreg_reg[1298]  ( .D(c[1302]), .CLK(clk), .RST(rst), .Q(sreg[1298]) );
  DFF \sreg_reg[1297]  ( .D(c[1301]), .CLK(clk), .RST(rst), .Q(sreg[1297]) );
  DFF \sreg_reg[1296]  ( .D(c[1300]), .CLK(clk), .RST(rst), .Q(sreg[1296]) );
  DFF \sreg_reg[1295]  ( .D(c[1299]), .CLK(clk), .RST(rst), .Q(sreg[1295]) );
  DFF \sreg_reg[1294]  ( .D(c[1298]), .CLK(clk), .RST(rst), .Q(sreg[1294]) );
  DFF \sreg_reg[1293]  ( .D(c[1297]), .CLK(clk), .RST(rst), .Q(sreg[1293]) );
  DFF \sreg_reg[1292]  ( .D(c[1296]), .CLK(clk), .RST(rst), .Q(sreg[1292]) );
  DFF \sreg_reg[1291]  ( .D(c[1295]), .CLK(clk), .RST(rst), .Q(sreg[1291]) );
  DFF \sreg_reg[1290]  ( .D(c[1294]), .CLK(clk), .RST(rst), .Q(sreg[1290]) );
  DFF \sreg_reg[1289]  ( .D(c[1293]), .CLK(clk), .RST(rst), .Q(sreg[1289]) );
  DFF \sreg_reg[1288]  ( .D(c[1292]), .CLK(clk), .RST(rst), .Q(sreg[1288]) );
  DFF \sreg_reg[1287]  ( .D(c[1291]), .CLK(clk), .RST(rst), .Q(sreg[1287]) );
  DFF \sreg_reg[1286]  ( .D(c[1290]), .CLK(clk), .RST(rst), .Q(sreg[1286]) );
  DFF \sreg_reg[1285]  ( .D(c[1289]), .CLK(clk), .RST(rst), .Q(sreg[1285]) );
  DFF \sreg_reg[1284]  ( .D(c[1288]), .CLK(clk), .RST(rst), .Q(sreg[1284]) );
  DFF \sreg_reg[1283]  ( .D(c[1287]), .CLK(clk), .RST(rst), .Q(sreg[1283]) );
  DFF \sreg_reg[1282]  ( .D(c[1286]), .CLK(clk), .RST(rst), .Q(sreg[1282]) );
  DFF \sreg_reg[1281]  ( .D(c[1285]), .CLK(clk), .RST(rst), .Q(sreg[1281]) );
  DFF \sreg_reg[1280]  ( .D(c[1284]), .CLK(clk), .RST(rst), .Q(sreg[1280]) );
  DFF \sreg_reg[1279]  ( .D(c[1283]), .CLK(clk), .RST(rst), .Q(sreg[1279]) );
  DFF \sreg_reg[1278]  ( .D(c[1282]), .CLK(clk), .RST(rst), .Q(sreg[1278]) );
  DFF \sreg_reg[1277]  ( .D(c[1281]), .CLK(clk), .RST(rst), .Q(sreg[1277]) );
  DFF \sreg_reg[1276]  ( .D(c[1280]), .CLK(clk), .RST(rst), .Q(sreg[1276]) );
  DFF \sreg_reg[1275]  ( .D(c[1279]), .CLK(clk), .RST(rst), .Q(sreg[1275]) );
  DFF \sreg_reg[1274]  ( .D(c[1278]), .CLK(clk), .RST(rst), .Q(sreg[1274]) );
  DFF \sreg_reg[1273]  ( .D(c[1277]), .CLK(clk), .RST(rst), .Q(sreg[1273]) );
  DFF \sreg_reg[1272]  ( .D(c[1276]), .CLK(clk), .RST(rst), .Q(sreg[1272]) );
  DFF \sreg_reg[1271]  ( .D(c[1275]), .CLK(clk), .RST(rst), .Q(sreg[1271]) );
  DFF \sreg_reg[1270]  ( .D(c[1274]), .CLK(clk), .RST(rst), .Q(sreg[1270]) );
  DFF \sreg_reg[1269]  ( .D(c[1273]), .CLK(clk), .RST(rst), .Q(sreg[1269]) );
  DFF \sreg_reg[1268]  ( .D(c[1272]), .CLK(clk), .RST(rst), .Q(sreg[1268]) );
  DFF \sreg_reg[1267]  ( .D(c[1271]), .CLK(clk), .RST(rst), .Q(sreg[1267]) );
  DFF \sreg_reg[1266]  ( .D(c[1270]), .CLK(clk), .RST(rst), .Q(sreg[1266]) );
  DFF \sreg_reg[1265]  ( .D(c[1269]), .CLK(clk), .RST(rst), .Q(sreg[1265]) );
  DFF \sreg_reg[1264]  ( .D(c[1268]), .CLK(clk), .RST(rst), .Q(sreg[1264]) );
  DFF \sreg_reg[1263]  ( .D(c[1267]), .CLK(clk), .RST(rst), .Q(sreg[1263]) );
  DFF \sreg_reg[1262]  ( .D(c[1266]), .CLK(clk), .RST(rst), .Q(sreg[1262]) );
  DFF \sreg_reg[1261]  ( .D(c[1265]), .CLK(clk), .RST(rst), .Q(sreg[1261]) );
  DFF \sreg_reg[1260]  ( .D(c[1264]), .CLK(clk), .RST(rst), .Q(sreg[1260]) );
  DFF \sreg_reg[1259]  ( .D(c[1263]), .CLK(clk), .RST(rst), .Q(sreg[1259]) );
  DFF \sreg_reg[1258]  ( .D(c[1262]), .CLK(clk), .RST(rst), .Q(sreg[1258]) );
  DFF \sreg_reg[1257]  ( .D(c[1261]), .CLK(clk), .RST(rst), .Q(sreg[1257]) );
  DFF \sreg_reg[1256]  ( .D(c[1260]), .CLK(clk), .RST(rst), .Q(sreg[1256]) );
  DFF \sreg_reg[1255]  ( .D(c[1259]), .CLK(clk), .RST(rst), .Q(sreg[1255]) );
  DFF \sreg_reg[1254]  ( .D(c[1258]), .CLK(clk), .RST(rst), .Q(sreg[1254]) );
  DFF \sreg_reg[1253]  ( .D(c[1257]), .CLK(clk), .RST(rst), .Q(sreg[1253]) );
  DFF \sreg_reg[1252]  ( .D(c[1256]), .CLK(clk), .RST(rst), .Q(sreg[1252]) );
  DFF \sreg_reg[1251]  ( .D(c[1255]), .CLK(clk), .RST(rst), .Q(sreg[1251]) );
  DFF \sreg_reg[1250]  ( .D(c[1254]), .CLK(clk), .RST(rst), .Q(sreg[1250]) );
  DFF \sreg_reg[1249]  ( .D(c[1253]), .CLK(clk), .RST(rst), .Q(sreg[1249]) );
  DFF \sreg_reg[1248]  ( .D(c[1252]), .CLK(clk), .RST(rst), .Q(sreg[1248]) );
  DFF \sreg_reg[1247]  ( .D(c[1251]), .CLK(clk), .RST(rst), .Q(sreg[1247]) );
  DFF \sreg_reg[1246]  ( .D(c[1250]), .CLK(clk), .RST(rst), .Q(sreg[1246]) );
  DFF \sreg_reg[1245]  ( .D(c[1249]), .CLK(clk), .RST(rst), .Q(sreg[1245]) );
  DFF \sreg_reg[1244]  ( .D(c[1248]), .CLK(clk), .RST(rst), .Q(sreg[1244]) );
  DFF \sreg_reg[1243]  ( .D(c[1247]), .CLK(clk), .RST(rst), .Q(sreg[1243]) );
  DFF \sreg_reg[1242]  ( .D(c[1246]), .CLK(clk), .RST(rst), .Q(sreg[1242]) );
  DFF \sreg_reg[1241]  ( .D(c[1245]), .CLK(clk), .RST(rst), .Q(sreg[1241]) );
  DFF \sreg_reg[1240]  ( .D(c[1244]), .CLK(clk), .RST(rst), .Q(sreg[1240]) );
  DFF \sreg_reg[1239]  ( .D(c[1243]), .CLK(clk), .RST(rst), .Q(sreg[1239]) );
  DFF \sreg_reg[1238]  ( .D(c[1242]), .CLK(clk), .RST(rst), .Q(sreg[1238]) );
  DFF \sreg_reg[1237]  ( .D(c[1241]), .CLK(clk), .RST(rst), .Q(sreg[1237]) );
  DFF \sreg_reg[1236]  ( .D(c[1240]), .CLK(clk), .RST(rst), .Q(sreg[1236]) );
  DFF \sreg_reg[1235]  ( .D(c[1239]), .CLK(clk), .RST(rst), .Q(sreg[1235]) );
  DFF \sreg_reg[1234]  ( .D(c[1238]), .CLK(clk), .RST(rst), .Q(sreg[1234]) );
  DFF \sreg_reg[1233]  ( .D(c[1237]), .CLK(clk), .RST(rst), .Q(sreg[1233]) );
  DFF \sreg_reg[1232]  ( .D(c[1236]), .CLK(clk), .RST(rst), .Q(sreg[1232]) );
  DFF \sreg_reg[1231]  ( .D(c[1235]), .CLK(clk), .RST(rst), .Q(sreg[1231]) );
  DFF \sreg_reg[1230]  ( .D(c[1234]), .CLK(clk), .RST(rst), .Q(sreg[1230]) );
  DFF \sreg_reg[1229]  ( .D(c[1233]), .CLK(clk), .RST(rst), .Q(sreg[1229]) );
  DFF \sreg_reg[1228]  ( .D(c[1232]), .CLK(clk), .RST(rst), .Q(sreg[1228]) );
  DFF \sreg_reg[1227]  ( .D(c[1231]), .CLK(clk), .RST(rst), .Q(sreg[1227]) );
  DFF \sreg_reg[1226]  ( .D(c[1230]), .CLK(clk), .RST(rst), .Q(sreg[1226]) );
  DFF \sreg_reg[1225]  ( .D(c[1229]), .CLK(clk), .RST(rst), .Q(sreg[1225]) );
  DFF \sreg_reg[1224]  ( .D(c[1228]), .CLK(clk), .RST(rst), .Q(sreg[1224]) );
  DFF \sreg_reg[1223]  ( .D(c[1227]), .CLK(clk), .RST(rst), .Q(sreg[1223]) );
  DFF \sreg_reg[1222]  ( .D(c[1226]), .CLK(clk), .RST(rst), .Q(sreg[1222]) );
  DFF \sreg_reg[1221]  ( .D(c[1225]), .CLK(clk), .RST(rst), .Q(sreg[1221]) );
  DFF \sreg_reg[1220]  ( .D(c[1224]), .CLK(clk), .RST(rst), .Q(sreg[1220]) );
  DFF \sreg_reg[1219]  ( .D(c[1223]), .CLK(clk), .RST(rst), .Q(sreg[1219]) );
  DFF \sreg_reg[1218]  ( .D(c[1222]), .CLK(clk), .RST(rst), .Q(sreg[1218]) );
  DFF \sreg_reg[1217]  ( .D(c[1221]), .CLK(clk), .RST(rst), .Q(sreg[1217]) );
  DFF \sreg_reg[1216]  ( .D(c[1220]), .CLK(clk), .RST(rst), .Q(sreg[1216]) );
  DFF \sreg_reg[1215]  ( .D(c[1219]), .CLK(clk), .RST(rst), .Q(sreg[1215]) );
  DFF \sreg_reg[1214]  ( .D(c[1218]), .CLK(clk), .RST(rst), .Q(sreg[1214]) );
  DFF \sreg_reg[1213]  ( .D(c[1217]), .CLK(clk), .RST(rst), .Q(sreg[1213]) );
  DFF \sreg_reg[1212]  ( .D(c[1216]), .CLK(clk), .RST(rst), .Q(sreg[1212]) );
  DFF \sreg_reg[1211]  ( .D(c[1215]), .CLK(clk), .RST(rst), .Q(sreg[1211]) );
  DFF \sreg_reg[1210]  ( .D(c[1214]), .CLK(clk), .RST(rst), .Q(sreg[1210]) );
  DFF \sreg_reg[1209]  ( .D(c[1213]), .CLK(clk), .RST(rst), .Q(sreg[1209]) );
  DFF \sreg_reg[1208]  ( .D(c[1212]), .CLK(clk), .RST(rst), .Q(sreg[1208]) );
  DFF \sreg_reg[1207]  ( .D(c[1211]), .CLK(clk), .RST(rst), .Q(sreg[1207]) );
  DFF \sreg_reg[1206]  ( .D(c[1210]), .CLK(clk), .RST(rst), .Q(sreg[1206]) );
  DFF \sreg_reg[1205]  ( .D(c[1209]), .CLK(clk), .RST(rst), .Q(sreg[1205]) );
  DFF \sreg_reg[1204]  ( .D(c[1208]), .CLK(clk), .RST(rst), .Q(sreg[1204]) );
  DFF \sreg_reg[1203]  ( .D(c[1207]), .CLK(clk), .RST(rst), .Q(sreg[1203]) );
  DFF \sreg_reg[1202]  ( .D(c[1206]), .CLK(clk), .RST(rst), .Q(sreg[1202]) );
  DFF \sreg_reg[1201]  ( .D(c[1205]), .CLK(clk), .RST(rst), .Q(sreg[1201]) );
  DFF \sreg_reg[1200]  ( .D(c[1204]), .CLK(clk), .RST(rst), .Q(sreg[1200]) );
  DFF \sreg_reg[1199]  ( .D(c[1203]), .CLK(clk), .RST(rst), .Q(sreg[1199]) );
  DFF \sreg_reg[1198]  ( .D(c[1202]), .CLK(clk), .RST(rst), .Q(sreg[1198]) );
  DFF \sreg_reg[1197]  ( .D(c[1201]), .CLK(clk), .RST(rst), .Q(sreg[1197]) );
  DFF \sreg_reg[1196]  ( .D(c[1200]), .CLK(clk), .RST(rst), .Q(sreg[1196]) );
  DFF \sreg_reg[1195]  ( .D(c[1199]), .CLK(clk), .RST(rst), .Q(sreg[1195]) );
  DFF \sreg_reg[1194]  ( .D(c[1198]), .CLK(clk), .RST(rst), .Q(sreg[1194]) );
  DFF \sreg_reg[1193]  ( .D(c[1197]), .CLK(clk), .RST(rst), .Q(sreg[1193]) );
  DFF \sreg_reg[1192]  ( .D(c[1196]), .CLK(clk), .RST(rst), .Q(sreg[1192]) );
  DFF \sreg_reg[1191]  ( .D(c[1195]), .CLK(clk), .RST(rst), .Q(sreg[1191]) );
  DFF \sreg_reg[1190]  ( .D(c[1194]), .CLK(clk), .RST(rst), .Q(sreg[1190]) );
  DFF \sreg_reg[1189]  ( .D(c[1193]), .CLK(clk), .RST(rst), .Q(sreg[1189]) );
  DFF \sreg_reg[1188]  ( .D(c[1192]), .CLK(clk), .RST(rst), .Q(sreg[1188]) );
  DFF \sreg_reg[1187]  ( .D(c[1191]), .CLK(clk), .RST(rst), .Q(sreg[1187]) );
  DFF \sreg_reg[1186]  ( .D(c[1190]), .CLK(clk), .RST(rst), .Q(sreg[1186]) );
  DFF \sreg_reg[1185]  ( .D(c[1189]), .CLK(clk), .RST(rst), .Q(sreg[1185]) );
  DFF \sreg_reg[1184]  ( .D(c[1188]), .CLK(clk), .RST(rst), .Q(sreg[1184]) );
  DFF \sreg_reg[1183]  ( .D(c[1187]), .CLK(clk), .RST(rst), .Q(sreg[1183]) );
  DFF \sreg_reg[1182]  ( .D(c[1186]), .CLK(clk), .RST(rst), .Q(sreg[1182]) );
  DFF \sreg_reg[1181]  ( .D(c[1185]), .CLK(clk), .RST(rst), .Q(sreg[1181]) );
  DFF \sreg_reg[1180]  ( .D(c[1184]), .CLK(clk), .RST(rst), .Q(sreg[1180]) );
  DFF \sreg_reg[1179]  ( .D(c[1183]), .CLK(clk), .RST(rst), .Q(sreg[1179]) );
  DFF \sreg_reg[1178]  ( .D(c[1182]), .CLK(clk), .RST(rst), .Q(sreg[1178]) );
  DFF \sreg_reg[1177]  ( .D(c[1181]), .CLK(clk), .RST(rst), .Q(sreg[1177]) );
  DFF \sreg_reg[1176]  ( .D(c[1180]), .CLK(clk), .RST(rst), .Q(sreg[1176]) );
  DFF \sreg_reg[1175]  ( .D(c[1179]), .CLK(clk), .RST(rst), .Q(sreg[1175]) );
  DFF \sreg_reg[1174]  ( .D(c[1178]), .CLK(clk), .RST(rst), .Q(sreg[1174]) );
  DFF \sreg_reg[1173]  ( .D(c[1177]), .CLK(clk), .RST(rst), .Q(sreg[1173]) );
  DFF \sreg_reg[1172]  ( .D(c[1176]), .CLK(clk), .RST(rst), .Q(sreg[1172]) );
  DFF \sreg_reg[1171]  ( .D(c[1175]), .CLK(clk), .RST(rst), .Q(sreg[1171]) );
  DFF \sreg_reg[1170]  ( .D(c[1174]), .CLK(clk), .RST(rst), .Q(sreg[1170]) );
  DFF \sreg_reg[1169]  ( .D(c[1173]), .CLK(clk), .RST(rst), .Q(sreg[1169]) );
  DFF \sreg_reg[1168]  ( .D(c[1172]), .CLK(clk), .RST(rst), .Q(sreg[1168]) );
  DFF \sreg_reg[1167]  ( .D(c[1171]), .CLK(clk), .RST(rst), .Q(sreg[1167]) );
  DFF \sreg_reg[1166]  ( .D(c[1170]), .CLK(clk), .RST(rst), .Q(sreg[1166]) );
  DFF \sreg_reg[1165]  ( .D(c[1169]), .CLK(clk), .RST(rst), .Q(sreg[1165]) );
  DFF \sreg_reg[1164]  ( .D(c[1168]), .CLK(clk), .RST(rst), .Q(sreg[1164]) );
  DFF \sreg_reg[1163]  ( .D(c[1167]), .CLK(clk), .RST(rst), .Q(sreg[1163]) );
  DFF \sreg_reg[1162]  ( .D(c[1166]), .CLK(clk), .RST(rst), .Q(sreg[1162]) );
  DFF \sreg_reg[1161]  ( .D(c[1165]), .CLK(clk), .RST(rst), .Q(sreg[1161]) );
  DFF \sreg_reg[1160]  ( .D(c[1164]), .CLK(clk), .RST(rst), .Q(sreg[1160]) );
  DFF \sreg_reg[1159]  ( .D(c[1163]), .CLK(clk), .RST(rst), .Q(sreg[1159]) );
  DFF \sreg_reg[1158]  ( .D(c[1162]), .CLK(clk), .RST(rst), .Q(sreg[1158]) );
  DFF \sreg_reg[1157]  ( .D(c[1161]), .CLK(clk), .RST(rst), .Q(sreg[1157]) );
  DFF \sreg_reg[1156]  ( .D(c[1160]), .CLK(clk), .RST(rst), .Q(sreg[1156]) );
  DFF \sreg_reg[1155]  ( .D(c[1159]), .CLK(clk), .RST(rst), .Q(sreg[1155]) );
  DFF \sreg_reg[1154]  ( .D(c[1158]), .CLK(clk), .RST(rst), .Q(sreg[1154]) );
  DFF \sreg_reg[1153]  ( .D(c[1157]), .CLK(clk), .RST(rst), .Q(sreg[1153]) );
  DFF \sreg_reg[1152]  ( .D(c[1156]), .CLK(clk), .RST(rst), .Q(sreg[1152]) );
  DFF \sreg_reg[1151]  ( .D(c[1155]), .CLK(clk), .RST(rst), .Q(sreg[1151]) );
  DFF \sreg_reg[1150]  ( .D(c[1154]), .CLK(clk), .RST(rst), .Q(sreg[1150]) );
  DFF \sreg_reg[1149]  ( .D(c[1153]), .CLK(clk), .RST(rst), .Q(sreg[1149]) );
  DFF \sreg_reg[1148]  ( .D(c[1152]), .CLK(clk), .RST(rst), .Q(sreg[1148]) );
  DFF \sreg_reg[1147]  ( .D(c[1151]), .CLK(clk), .RST(rst), .Q(sreg[1147]) );
  DFF \sreg_reg[1146]  ( .D(c[1150]), .CLK(clk), .RST(rst), .Q(sreg[1146]) );
  DFF \sreg_reg[1145]  ( .D(c[1149]), .CLK(clk), .RST(rst), .Q(sreg[1145]) );
  DFF \sreg_reg[1144]  ( .D(c[1148]), .CLK(clk), .RST(rst), .Q(sreg[1144]) );
  DFF \sreg_reg[1143]  ( .D(c[1147]), .CLK(clk), .RST(rst), .Q(sreg[1143]) );
  DFF \sreg_reg[1142]  ( .D(c[1146]), .CLK(clk), .RST(rst), .Q(sreg[1142]) );
  DFF \sreg_reg[1141]  ( .D(c[1145]), .CLK(clk), .RST(rst), .Q(sreg[1141]) );
  DFF \sreg_reg[1140]  ( .D(c[1144]), .CLK(clk), .RST(rst), .Q(sreg[1140]) );
  DFF \sreg_reg[1139]  ( .D(c[1143]), .CLK(clk), .RST(rst), .Q(sreg[1139]) );
  DFF \sreg_reg[1138]  ( .D(c[1142]), .CLK(clk), .RST(rst), .Q(sreg[1138]) );
  DFF \sreg_reg[1137]  ( .D(c[1141]), .CLK(clk), .RST(rst), .Q(sreg[1137]) );
  DFF \sreg_reg[1136]  ( .D(c[1140]), .CLK(clk), .RST(rst), .Q(sreg[1136]) );
  DFF \sreg_reg[1135]  ( .D(c[1139]), .CLK(clk), .RST(rst), .Q(sreg[1135]) );
  DFF \sreg_reg[1134]  ( .D(c[1138]), .CLK(clk), .RST(rst), .Q(sreg[1134]) );
  DFF \sreg_reg[1133]  ( .D(c[1137]), .CLK(clk), .RST(rst), .Q(sreg[1133]) );
  DFF \sreg_reg[1132]  ( .D(c[1136]), .CLK(clk), .RST(rst), .Q(sreg[1132]) );
  DFF \sreg_reg[1131]  ( .D(c[1135]), .CLK(clk), .RST(rst), .Q(sreg[1131]) );
  DFF \sreg_reg[1130]  ( .D(c[1134]), .CLK(clk), .RST(rst), .Q(sreg[1130]) );
  DFF \sreg_reg[1129]  ( .D(c[1133]), .CLK(clk), .RST(rst), .Q(sreg[1129]) );
  DFF \sreg_reg[1128]  ( .D(c[1132]), .CLK(clk), .RST(rst), .Q(sreg[1128]) );
  DFF \sreg_reg[1127]  ( .D(c[1131]), .CLK(clk), .RST(rst), .Q(sreg[1127]) );
  DFF \sreg_reg[1126]  ( .D(c[1130]), .CLK(clk), .RST(rst), .Q(sreg[1126]) );
  DFF \sreg_reg[1125]  ( .D(c[1129]), .CLK(clk), .RST(rst), .Q(sreg[1125]) );
  DFF \sreg_reg[1124]  ( .D(c[1128]), .CLK(clk), .RST(rst), .Q(sreg[1124]) );
  DFF \sreg_reg[1123]  ( .D(c[1127]), .CLK(clk), .RST(rst), .Q(sreg[1123]) );
  DFF \sreg_reg[1122]  ( .D(c[1126]), .CLK(clk), .RST(rst), .Q(sreg[1122]) );
  DFF \sreg_reg[1121]  ( .D(c[1125]), .CLK(clk), .RST(rst), .Q(sreg[1121]) );
  DFF \sreg_reg[1120]  ( .D(c[1124]), .CLK(clk), .RST(rst), .Q(sreg[1120]) );
  DFF \sreg_reg[1119]  ( .D(c[1123]), .CLK(clk), .RST(rst), .Q(sreg[1119]) );
  DFF \sreg_reg[1118]  ( .D(c[1122]), .CLK(clk), .RST(rst), .Q(sreg[1118]) );
  DFF \sreg_reg[1117]  ( .D(c[1121]), .CLK(clk), .RST(rst), .Q(sreg[1117]) );
  DFF \sreg_reg[1116]  ( .D(c[1120]), .CLK(clk), .RST(rst), .Q(sreg[1116]) );
  DFF \sreg_reg[1115]  ( .D(c[1119]), .CLK(clk), .RST(rst), .Q(sreg[1115]) );
  DFF \sreg_reg[1114]  ( .D(c[1118]), .CLK(clk), .RST(rst), .Q(sreg[1114]) );
  DFF \sreg_reg[1113]  ( .D(c[1117]), .CLK(clk), .RST(rst), .Q(sreg[1113]) );
  DFF \sreg_reg[1112]  ( .D(c[1116]), .CLK(clk), .RST(rst), .Q(sreg[1112]) );
  DFF \sreg_reg[1111]  ( .D(c[1115]), .CLK(clk), .RST(rst), .Q(sreg[1111]) );
  DFF \sreg_reg[1110]  ( .D(c[1114]), .CLK(clk), .RST(rst), .Q(sreg[1110]) );
  DFF \sreg_reg[1109]  ( .D(c[1113]), .CLK(clk), .RST(rst), .Q(sreg[1109]) );
  DFF \sreg_reg[1108]  ( .D(c[1112]), .CLK(clk), .RST(rst), .Q(sreg[1108]) );
  DFF \sreg_reg[1107]  ( .D(c[1111]), .CLK(clk), .RST(rst), .Q(sreg[1107]) );
  DFF \sreg_reg[1106]  ( .D(c[1110]), .CLK(clk), .RST(rst), .Q(sreg[1106]) );
  DFF \sreg_reg[1105]  ( .D(c[1109]), .CLK(clk), .RST(rst), .Q(sreg[1105]) );
  DFF \sreg_reg[1104]  ( .D(c[1108]), .CLK(clk), .RST(rst), .Q(sreg[1104]) );
  DFF \sreg_reg[1103]  ( .D(c[1107]), .CLK(clk), .RST(rst), .Q(sreg[1103]) );
  DFF \sreg_reg[1102]  ( .D(c[1106]), .CLK(clk), .RST(rst), .Q(sreg[1102]) );
  DFF \sreg_reg[1101]  ( .D(c[1105]), .CLK(clk), .RST(rst), .Q(sreg[1101]) );
  DFF \sreg_reg[1100]  ( .D(c[1104]), .CLK(clk), .RST(rst), .Q(sreg[1100]) );
  DFF \sreg_reg[1099]  ( .D(c[1103]), .CLK(clk), .RST(rst), .Q(sreg[1099]) );
  DFF \sreg_reg[1098]  ( .D(c[1102]), .CLK(clk), .RST(rst), .Q(sreg[1098]) );
  DFF \sreg_reg[1097]  ( .D(c[1101]), .CLK(clk), .RST(rst), .Q(sreg[1097]) );
  DFF \sreg_reg[1096]  ( .D(c[1100]), .CLK(clk), .RST(rst), .Q(sreg[1096]) );
  DFF \sreg_reg[1095]  ( .D(c[1099]), .CLK(clk), .RST(rst), .Q(sreg[1095]) );
  DFF \sreg_reg[1094]  ( .D(c[1098]), .CLK(clk), .RST(rst), .Q(sreg[1094]) );
  DFF \sreg_reg[1093]  ( .D(c[1097]), .CLK(clk), .RST(rst), .Q(sreg[1093]) );
  DFF \sreg_reg[1092]  ( .D(c[1096]), .CLK(clk), .RST(rst), .Q(sreg[1092]) );
  DFF \sreg_reg[1091]  ( .D(c[1095]), .CLK(clk), .RST(rst), .Q(sreg[1091]) );
  DFF \sreg_reg[1090]  ( .D(c[1094]), .CLK(clk), .RST(rst), .Q(sreg[1090]) );
  DFF \sreg_reg[1089]  ( .D(c[1093]), .CLK(clk), .RST(rst), .Q(sreg[1089]) );
  DFF \sreg_reg[1088]  ( .D(c[1092]), .CLK(clk), .RST(rst), .Q(sreg[1088]) );
  DFF \sreg_reg[1087]  ( .D(c[1091]), .CLK(clk), .RST(rst), .Q(sreg[1087]) );
  DFF \sreg_reg[1086]  ( .D(c[1090]), .CLK(clk), .RST(rst), .Q(sreg[1086]) );
  DFF \sreg_reg[1085]  ( .D(c[1089]), .CLK(clk), .RST(rst), .Q(sreg[1085]) );
  DFF \sreg_reg[1084]  ( .D(c[1088]), .CLK(clk), .RST(rst), .Q(sreg[1084]) );
  DFF \sreg_reg[1083]  ( .D(c[1087]), .CLK(clk), .RST(rst), .Q(sreg[1083]) );
  DFF \sreg_reg[1082]  ( .D(c[1086]), .CLK(clk), .RST(rst), .Q(sreg[1082]) );
  DFF \sreg_reg[1081]  ( .D(c[1085]), .CLK(clk), .RST(rst), .Q(sreg[1081]) );
  DFF \sreg_reg[1080]  ( .D(c[1084]), .CLK(clk), .RST(rst), .Q(sreg[1080]) );
  DFF \sreg_reg[1079]  ( .D(c[1083]), .CLK(clk), .RST(rst), .Q(sreg[1079]) );
  DFF \sreg_reg[1078]  ( .D(c[1082]), .CLK(clk), .RST(rst), .Q(sreg[1078]) );
  DFF \sreg_reg[1077]  ( .D(c[1081]), .CLK(clk), .RST(rst), .Q(sreg[1077]) );
  DFF \sreg_reg[1076]  ( .D(c[1080]), .CLK(clk), .RST(rst), .Q(sreg[1076]) );
  DFF \sreg_reg[1075]  ( .D(c[1079]), .CLK(clk), .RST(rst), .Q(sreg[1075]) );
  DFF \sreg_reg[1074]  ( .D(c[1078]), .CLK(clk), .RST(rst), .Q(sreg[1074]) );
  DFF \sreg_reg[1073]  ( .D(c[1077]), .CLK(clk), .RST(rst), .Q(sreg[1073]) );
  DFF \sreg_reg[1072]  ( .D(c[1076]), .CLK(clk), .RST(rst), .Q(sreg[1072]) );
  DFF \sreg_reg[1071]  ( .D(c[1075]), .CLK(clk), .RST(rst), .Q(sreg[1071]) );
  DFF \sreg_reg[1070]  ( .D(c[1074]), .CLK(clk), .RST(rst), .Q(sreg[1070]) );
  DFF \sreg_reg[1069]  ( .D(c[1073]), .CLK(clk), .RST(rst), .Q(sreg[1069]) );
  DFF \sreg_reg[1068]  ( .D(c[1072]), .CLK(clk), .RST(rst), .Q(sreg[1068]) );
  DFF \sreg_reg[1067]  ( .D(c[1071]), .CLK(clk), .RST(rst), .Q(sreg[1067]) );
  DFF \sreg_reg[1066]  ( .D(c[1070]), .CLK(clk), .RST(rst), .Q(sreg[1066]) );
  DFF \sreg_reg[1065]  ( .D(c[1069]), .CLK(clk), .RST(rst), .Q(sreg[1065]) );
  DFF \sreg_reg[1064]  ( .D(c[1068]), .CLK(clk), .RST(rst), .Q(sreg[1064]) );
  DFF \sreg_reg[1063]  ( .D(c[1067]), .CLK(clk), .RST(rst), .Q(sreg[1063]) );
  DFF \sreg_reg[1062]  ( .D(c[1066]), .CLK(clk), .RST(rst), .Q(sreg[1062]) );
  DFF \sreg_reg[1061]  ( .D(c[1065]), .CLK(clk), .RST(rst), .Q(sreg[1061]) );
  DFF \sreg_reg[1060]  ( .D(c[1064]), .CLK(clk), .RST(rst), .Q(sreg[1060]) );
  DFF \sreg_reg[1059]  ( .D(c[1063]), .CLK(clk), .RST(rst), .Q(sreg[1059]) );
  DFF \sreg_reg[1058]  ( .D(c[1062]), .CLK(clk), .RST(rst), .Q(sreg[1058]) );
  DFF \sreg_reg[1057]  ( .D(c[1061]), .CLK(clk), .RST(rst), .Q(sreg[1057]) );
  DFF \sreg_reg[1056]  ( .D(c[1060]), .CLK(clk), .RST(rst), .Q(sreg[1056]) );
  DFF \sreg_reg[1055]  ( .D(c[1059]), .CLK(clk), .RST(rst), .Q(sreg[1055]) );
  DFF \sreg_reg[1054]  ( .D(c[1058]), .CLK(clk), .RST(rst), .Q(sreg[1054]) );
  DFF \sreg_reg[1053]  ( .D(c[1057]), .CLK(clk), .RST(rst), .Q(sreg[1053]) );
  DFF \sreg_reg[1052]  ( .D(c[1056]), .CLK(clk), .RST(rst), .Q(sreg[1052]) );
  DFF \sreg_reg[1051]  ( .D(c[1055]), .CLK(clk), .RST(rst), .Q(sreg[1051]) );
  DFF \sreg_reg[1050]  ( .D(c[1054]), .CLK(clk), .RST(rst), .Q(sreg[1050]) );
  DFF \sreg_reg[1049]  ( .D(c[1053]), .CLK(clk), .RST(rst), .Q(sreg[1049]) );
  DFF \sreg_reg[1048]  ( .D(c[1052]), .CLK(clk), .RST(rst), .Q(sreg[1048]) );
  DFF \sreg_reg[1047]  ( .D(c[1051]), .CLK(clk), .RST(rst), .Q(sreg[1047]) );
  DFF \sreg_reg[1046]  ( .D(c[1050]), .CLK(clk), .RST(rst), .Q(sreg[1046]) );
  DFF \sreg_reg[1045]  ( .D(c[1049]), .CLK(clk), .RST(rst), .Q(sreg[1045]) );
  DFF \sreg_reg[1044]  ( .D(c[1048]), .CLK(clk), .RST(rst), .Q(sreg[1044]) );
  DFF \sreg_reg[1043]  ( .D(c[1047]), .CLK(clk), .RST(rst), .Q(sreg[1043]) );
  DFF \sreg_reg[1042]  ( .D(c[1046]), .CLK(clk), .RST(rst), .Q(sreg[1042]) );
  DFF \sreg_reg[1041]  ( .D(c[1045]), .CLK(clk), .RST(rst), .Q(sreg[1041]) );
  DFF \sreg_reg[1040]  ( .D(c[1044]), .CLK(clk), .RST(rst), .Q(sreg[1040]) );
  DFF \sreg_reg[1039]  ( .D(c[1043]), .CLK(clk), .RST(rst), .Q(sreg[1039]) );
  DFF \sreg_reg[1038]  ( .D(c[1042]), .CLK(clk), .RST(rst), .Q(sreg[1038]) );
  DFF \sreg_reg[1037]  ( .D(c[1041]), .CLK(clk), .RST(rst), .Q(sreg[1037]) );
  DFF \sreg_reg[1036]  ( .D(c[1040]), .CLK(clk), .RST(rst), .Q(sreg[1036]) );
  DFF \sreg_reg[1035]  ( .D(c[1039]), .CLK(clk), .RST(rst), .Q(sreg[1035]) );
  DFF \sreg_reg[1034]  ( .D(c[1038]), .CLK(clk), .RST(rst), .Q(sreg[1034]) );
  DFF \sreg_reg[1033]  ( .D(c[1037]), .CLK(clk), .RST(rst), .Q(sreg[1033]) );
  DFF \sreg_reg[1032]  ( .D(c[1036]), .CLK(clk), .RST(rst), .Q(sreg[1032]) );
  DFF \sreg_reg[1031]  ( .D(c[1035]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1030]  ( .D(c[1034]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1029]  ( .D(c[1033]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1028]  ( .D(c[1032]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1027]  ( .D(c[1031]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1026]  ( .D(c[1030]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1025]  ( .D(c[1029]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1024]  ( .D(c[1028]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1023]  ( .D(c[1027]), .CLK(clk), .RST(rst), .Q(sreg[1023]) );
  DFF \sreg_reg[1022]  ( .D(c[1026]), .CLK(clk), .RST(rst), .Q(sreg[1022]) );
  DFF \sreg_reg[1021]  ( .D(c[1025]), .CLK(clk), .RST(rst), .Q(sreg[1021]) );
  DFF \sreg_reg[1020]  ( .D(c[1024]), .CLK(clk), .RST(rst), .Q(sreg[1020]) );
  DFF \sreg_reg[1019]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1019]) );
  DFF \sreg_reg[1018]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1018]) );
  DFF \sreg_reg[1017]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1017]) );
  DFF \sreg_reg[1016]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1016]) );
  DFF \sreg_reg[1015]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1014]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1013]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1012]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1011]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1010]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1009]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1008]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1007]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1006]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1005]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1004]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1003]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1002]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1001]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1000]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[999]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[998]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[997]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[996]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[995]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[994]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[993]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[992]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[991]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[990]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[989]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[988]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[987]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[986]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[985]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[984]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[983]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[982]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[981]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[980]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[979]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[978]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[977]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[976]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[975]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[974]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[973]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[972]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[971]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[970]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[969]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[968]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[967]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[966]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[965]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[964]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[963]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[962]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[961]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[960]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[959]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[958]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[957]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[956]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[955]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[954]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[953]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[952]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[951]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[950]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[949]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[948]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[947]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[946]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[945]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[944]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[943]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[942]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[941]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[940]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[939]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[938]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[937]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[936]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[935]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[934]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[933]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[932]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[931]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[930]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[929]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[928]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[927]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[926]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[925]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[924]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[923]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[922]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[921]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[920]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[919]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[918]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[917]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[916]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[915]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[914]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[913]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[912]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[911]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[910]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[909]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[908]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[907]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[906]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[905]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[904]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[903]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[902]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[901]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[900]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[899]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[898]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[897]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[896]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[895]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[894]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[893]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[892]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[891]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[890]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[889]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[888]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[887]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[886]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[885]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[884]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[883]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[882]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[881]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[880]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[879]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[878]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[877]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[876]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[875]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[874]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[873]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[872]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[871]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[870]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[869]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[868]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[867]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[866]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[865]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[864]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[863]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[862]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[861]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[860]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[859]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[858]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[857]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[856]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[855]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[854]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[853]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[852]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[851]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[850]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[849]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[848]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[847]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[846]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[845]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[844]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[843]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[842]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[841]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[840]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[839]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[838]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[837]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[836]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[835]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[834]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[833]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[832]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[831]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[830]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[829]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[828]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[827]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[826]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[825]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[824]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[823]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[822]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[821]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[820]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[819]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[818]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[817]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[816]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[815]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[814]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[813]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[812]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[811]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[810]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[809]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[808]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[807]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[806]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[805]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[804]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[803]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[802]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[801]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[800]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[799]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[798]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[797]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[796]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[795]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[794]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[793]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[792]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[791]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[790]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[789]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[788]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[787]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[786]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[785]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[784]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[783]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[782]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[781]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[780]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[779]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[778]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[777]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[776]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[775]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[774]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[773]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[772]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[771]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[770]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[769]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[768]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[767]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[766]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[765]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[764]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[763]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[762]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[761]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[760]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[759]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[758]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[757]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[756]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[755]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[754]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[753]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[752]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[751]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[750]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[749]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[748]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[747]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[746]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[745]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[744]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[743]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[742]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[741]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[740]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[739]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[738]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[737]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[736]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[735]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[734]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[733]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[732]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[731]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[730]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[729]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[728]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[727]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[726]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[725]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[724]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[723]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[722]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[721]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[720]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[719]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[718]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[717]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[716]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[715]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[714]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[713]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[712]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[711]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[710]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[709]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[708]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[707]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[706]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[705]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[704]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[703]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[702]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[701]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[700]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[699]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[698]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[697]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[696]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[695]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[694]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[693]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[692]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[691]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[690]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[689]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[688]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[687]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[686]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[685]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[684]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[683]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[682]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[681]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[680]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[679]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[678]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[677]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[676]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[675]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[674]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[673]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[672]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[671]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[670]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[669]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[668]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[667]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[666]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[665]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[664]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[663]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[662]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[661]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[660]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[659]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[658]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[657]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[656]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[655]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[654]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[653]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[652]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[651]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[650]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[649]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[648]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[647]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[646]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[645]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[644]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[643]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[642]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[641]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[640]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[639]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[638]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[637]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[636]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[635]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[634]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[633]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[632]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[631]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[630]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[629]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[628]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[627]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[626]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[625]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[624]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[623]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[622]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[621]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[620]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[619]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[618]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[617]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[616]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[615]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[614]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[613]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[612]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[611]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[610]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[609]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[608]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[607]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[606]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[605]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[604]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[603]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[602]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[601]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[600]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[599]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[598]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[597]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[596]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[595]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[594]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[593]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[592]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[591]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[590]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[589]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[588]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[587]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[586]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[585]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[584]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[583]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[582]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[581]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[580]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[579]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[578]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[577]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[576]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[575]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[574]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[573]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[572]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[571]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[570]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[569]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[568]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[567]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[566]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[565]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[564]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[563]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[562]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[561]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[560]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[559]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[558]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[557]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[556]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[555]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[554]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[553]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[552]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[551]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[550]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[549]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[548]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[547]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[546]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[545]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[544]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[543]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[542]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[541]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[540]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[539]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[538]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[537]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[536]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[535]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[534]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[533]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[532]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[531]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[530]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[529]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[528]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[527]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[526]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[525]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[524]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[523]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[522]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[521]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[520]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[519]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[518]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[517]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[516]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[515]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[514]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[513]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[512]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[511]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[510]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[509]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[508]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[507]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[506]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[505]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[504]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[503]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[502]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[501]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[500]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[499]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[498]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[497]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[496]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[495]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[494]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[493]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[492]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[491]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[490]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[489]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[488]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[487]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[486]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[485]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[484]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[483]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[482]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[481]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[480]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[479]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[478]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[477]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[476]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[475]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[474]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[473]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[472]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[471]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[470]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[469]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[468]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[467]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[466]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[465]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[464]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[463]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[462]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[461]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[460]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[459]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[458]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[457]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[456]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[455]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[454]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[453]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[452]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[451]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[450]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[449]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[448]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[447]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[446]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[445]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[444]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[443]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[442]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[441]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[440]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[439]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[438]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[437]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[436]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[435]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[434]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[433]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[432]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[431]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[430]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[429]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[428]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[427]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[426]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[425]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[424]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[423]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[422]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[421]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[420]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[419]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[418]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[417]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[416]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[415]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[414]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[413]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[412]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[411]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[410]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[409]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[408]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[407]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[406]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[405]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[404]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[403]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[402]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[401]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[400]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[399]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[398]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[397]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[396]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[395]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[394]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[393]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[392]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[391]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[390]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[389]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[388]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[387]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[386]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[385]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[384]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[383]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[382]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[381]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[380]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[379]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[378]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[377]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[376]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[375]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[374]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[373]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[372]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[371]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[370]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[369]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[368]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[367]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[366]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[365]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[364]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[363]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[362]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[361]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[360]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[359]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[358]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[357]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[356]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[355]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[354]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[353]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[352]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[351]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[350]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[349]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[348]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[347]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[346]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[345]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[344]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[343]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[342]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[341]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[340]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[339]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[338]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[337]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[336]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[335]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[334]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[333]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[332]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[331]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[330]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[329]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[328]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[327]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[326]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[325]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[324]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[323]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[322]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[321]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[320]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[319]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[318]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[317]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[316]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[315]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[314]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[313]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[312]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[311]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[310]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[309]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[308]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[307]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[306]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[305]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[304]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[303]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[302]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[301]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[300]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[299]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[298]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[297]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[296]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[295]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[294]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[293]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[292]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[291]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[290]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[289]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[288]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[287]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[286]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[285]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[284]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[283]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[282]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[281]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[280]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[279]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[278]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[277]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[276]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[275]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[274]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[273]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[272]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[271]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[270]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[269]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[268]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[267]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[266]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[265]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[264]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[263]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[262]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[261]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[260]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[259]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[258]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[257]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[256]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[255]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[254]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NANDN U7 ( .A(n2604), .B(n2173), .Z(n1) );
  NANDN U8 ( .A(n2583), .B(n2174), .Z(n2) );
  AND U9 ( .A(n1), .B(n2), .Z(n2610) );
  NANDN U10 ( .A(n2898), .B(n2173), .Z(n3) );
  NANDN U11 ( .A(n2877), .B(n2174), .Z(n4) );
  AND U12 ( .A(n3), .B(n4), .Z(n2904) );
  NANDN U13 ( .A(n3192), .B(n2173), .Z(n5) );
  NANDN U14 ( .A(n3171), .B(n2174), .Z(n6) );
  AND U15 ( .A(n5), .B(n6), .Z(n3198) );
  NANDN U16 ( .A(n3486), .B(n2173), .Z(n7) );
  NANDN U17 ( .A(n3465), .B(n2174), .Z(n8) );
  AND U18 ( .A(n7), .B(n8), .Z(n3492) );
  NANDN U19 ( .A(n3780), .B(n2173), .Z(n9) );
  NANDN U20 ( .A(n3759), .B(n2174), .Z(n10) );
  AND U21 ( .A(n9), .B(n10), .Z(n3786) );
  NANDN U22 ( .A(n4074), .B(n2173), .Z(n11) );
  NANDN U23 ( .A(n4053), .B(n2174), .Z(n12) );
  AND U24 ( .A(n11), .B(n12), .Z(n4080) );
  NANDN U25 ( .A(n4368), .B(n2173), .Z(n13) );
  NANDN U26 ( .A(n4347), .B(n2174), .Z(n14) );
  AND U27 ( .A(n13), .B(n14), .Z(n4374) );
  NANDN U28 ( .A(n4658), .B(n2173), .Z(n15) );
  NANDN U29 ( .A(n4637), .B(n2174), .Z(n16) );
  AND U30 ( .A(n15), .B(n16), .Z(n4664) );
  NANDN U31 ( .A(n4952), .B(n2173), .Z(n17) );
  NANDN U32 ( .A(n4931), .B(n2174), .Z(n18) );
  AND U33 ( .A(n17), .B(n18), .Z(n4958) );
  NANDN U34 ( .A(n5246), .B(n2173), .Z(n19) );
  NANDN U35 ( .A(n5225), .B(n2174), .Z(n20) );
  AND U36 ( .A(n19), .B(n20), .Z(n5252) );
  NANDN U37 ( .A(n5540), .B(n2173), .Z(n21) );
  NANDN U38 ( .A(n5519), .B(n2174), .Z(n22) );
  AND U39 ( .A(n21), .B(n22), .Z(n5546) );
  NANDN U40 ( .A(n5834), .B(n2173), .Z(n23) );
  NANDN U41 ( .A(n5813), .B(n2174), .Z(n24) );
  AND U42 ( .A(n23), .B(n24), .Z(n5840) );
  NANDN U43 ( .A(n6128), .B(n2173), .Z(n25) );
  NANDN U44 ( .A(n6107), .B(n2174), .Z(n26) );
  AND U45 ( .A(n25), .B(n26), .Z(n6134) );
  NANDN U46 ( .A(n6420), .B(n2173), .Z(n27) );
  NANDN U47 ( .A(n6401), .B(n2174), .Z(n28) );
  AND U48 ( .A(n27), .B(n28), .Z(n6427) );
  NANDN U49 ( .A(n6712), .B(n2173), .Z(n29) );
  NANDN U50 ( .A(n6691), .B(n2174), .Z(n30) );
  AND U51 ( .A(n29), .B(n30), .Z(n6718) );
  NANDN U52 ( .A(n6998), .B(n2173), .Z(n31) );
  NANDN U53 ( .A(n6977), .B(n2174), .Z(n32) );
  AND U54 ( .A(n31), .B(n32), .Z(n7004) );
  NANDN U55 ( .A(n7288), .B(n2173), .Z(n33) );
  NANDN U56 ( .A(n7267), .B(n2174), .Z(n34) );
  AND U57 ( .A(n33), .B(n34), .Z(n7294) );
  NANDN U58 ( .A(n7578), .B(n2173), .Z(n35) );
  NANDN U59 ( .A(n7557), .B(n2174), .Z(n36) );
  AND U60 ( .A(n35), .B(n36), .Z(n7584) );
  NANDN U61 ( .A(n7868), .B(n2173), .Z(n37) );
  NANDN U62 ( .A(n7847), .B(n2174), .Z(n38) );
  AND U63 ( .A(n37), .B(n38), .Z(n7874) );
  NANDN U64 ( .A(n8158), .B(n2173), .Z(n39) );
  NANDN U65 ( .A(n8137), .B(n2174), .Z(n40) );
  AND U66 ( .A(n39), .B(n40), .Z(n8164) );
  NANDN U67 ( .A(n8448), .B(n2173), .Z(n41) );
  NANDN U68 ( .A(n8427), .B(n2174), .Z(n42) );
  AND U69 ( .A(n41), .B(n42), .Z(n8454) );
  NANDN U70 ( .A(n8742), .B(n2173), .Z(n43) );
  NANDN U71 ( .A(n8721), .B(n2174), .Z(n44) );
  AND U72 ( .A(n43), .B(n44), .Z(n8748) );
  NANDN U73 ( .A(n9036), .B(n2173), .Z(n45) );
  NANDN U74 ( .A(n9015), .B(n2174), .Z(n46) );
  AND U75 ( .A(n45), .B(n46), .Z(n9042) );
  NANDN U76 ( .A(n9322), .B(n2173), .Z(n47) );
  NANDN U77 ( .A(n9301), .B(n2174), .Z(n48) );
  AND U78 ( .A(n47), .B(n48), .Z(n9328) );
  NANDN U79 ( .A(n9616), .B(n2173), .Z(n49) );
  NANDN U80 ( .A(n9595), .B(n2174), .Z(n50) );
  AND U81 ( .A(n49), .B(n50), .Z(n9622) );
  NANDN U82 ( .A(n9910), .B(n2173), .Z(n51) );
  NANDN U83 ( .A(n9889), .B(n2174), .Z(n52) );
  AND U84 ( .A(n51), .B(n52), .Z(n9916) );
  NANDN U85 ( .A(n10204), .B(n2173), .Z(n53) );
  NANDN U86 ( .A(n10183), .B(n2174), .Z(n54) );
  AND U87 ( .A(n53), .B(n54), .Z(n10210) );
  NANDN U88 ( .A(n10498), .B(n2173), .Z(n55) );
  NANDN U89 ( .A(n10477), .B(n2174), .Z(n56) );
  AND U90 ( .A(n55), .B(n56), .Z(n10504) );
  NANDN U91 ( .A(n10792), .B(n2173), .Z(n57) );
  NANDN U92 ( .A(n10771), .B(n2174), .Z(n58) );
  AND U93 ( .A(n57), .B(n58), .Z(n10798) );
  NANDN U94 ( .A(n11086), .B(n2173), .Z(n59) );
  NANDN U95 ( .A(n11065), .B(n2174), .Z(n60) );
  AND U96 ( .A(n59), .B(n60), .Z(n11092) );
  NANDN U97 ( .A(n11380), .B(n2173), .Z(n61) );
  NANDN U98 ( .A(n11359), .B(n2174), .Z(n62) );
  AND U99 ( .A(n61), .B(n62), .Z(n11386) );
  NANDN U100 ( .A(n11674), .B(n2173), .Z(n63) );
  NANDN U101 ( .A(n11653), .B(n2174), .Z(n64) );
  AND U102 ( .A(n63), .B(n64), .Z(n11680) );
  NANDN U103 ( .A(n11960), .B(n2173), .Z(n65) );
  NANDN U104 ( .A(n11939), .B(n2174), .Z(n66) );
  AND U105 ( .A(n65), .B(n66), .Z(n11966) );
  NANDN U106 ( .A(n12254), .B(n2173), .Z(n67) );
  NANDN U107 ( .A(n12233), .B(n2174), .Z(n68) );
  AND U108 ( .A(n67), .B(n68), .Z(n12260) );
  NANDN U109 ( .A(n12548), .B(n2173), .Z(n69) );
  NANDN U110 ( .A(n12527), .B(n2174), .Z(n70) );
  AND U111 ( .A(n69), .B(n70), .Z(n12554) );
  NANDN U112 ( .A(n12838), .B(n2173), .Z(n71) );
  NANDN U113 ( .A(n12817), .B(n2174), .Z(n72) );
  AND U114 ( .A(n71), .B(n72), .Z(n12844) );
  NANDN U115 ( .A(n13132), .B(n2173), .Z(n73) );
  NANDN U116 ( .A(n13111), .B(n2174), .Z(n74) );
  AND U117 ( .A(n73), .B(n74), .Z(n13138) );
  NANDN U118 ( .A(n13426), .B(n2173), .Z(n75) );
  NANDN U119 ( .A(n13405), .B(n2174), .Z(n76) );
  AND U120 ( .A(n75), .B(n76), .Z(n13432) );
  NANDN U121 ( .A(n13720), .B(n2173), .Z(n77) );
  NANDN U122 ( .A(n13699), .B(n2174), .Z(n78) );
  AND U123 ( .A(n77), .B(n78), .Z(n13726) );
  NANDN U124 ( .A(n14010), .B(n2173), .Z(n79) );
  NANDN U125 ( .A(n13989), .B(n2174), .Z(n80) );
  AND U126 ( .A(n79), .B(n80), .Z(n14016) );
  NANDN U127 ( .A(n14304), .B(n2173), .Z(n81) );
  NANDN U128 ( .A(n14283), .B(n2174), .Z(n82) );
  AND U129 ( .A(n81), .B(n82), .Z(n14310) );
  NANDN U130 ( .A(n14598), .B(n2173), .Z(n83) );
  NANDN U131 ( .A(n14577), .B(n2174), .Z(n84) );
  AND U132 ( .A(n83), .B(n84), .Z(n14604) );
  NANDN U133 ( .A(n14888), .B(n2173), .Z(n85) );
  NANDN U134 ( .A(n14867), .B(n2174), .Z(n86) );
  AND U135 ( .A(n85), .B(n86), .Z(n14894) );
  NANDN U136 ( .A(n15182), .B(n2173), .Z(n87) );
  NANDN U137 ( .A(n15161), .B(n2174), .Z(n88) );
  AND U138 ( .A(n87), .B(n88), .Z(n15188) );
  NANDN U139 ( .A(n15476), .B(n2173), .Z(n89) );
  NANDN U140 ( .A(n15455), .B(n2174), .Z(n90) );
  AND U141 ( .A(n89), .B(n90), .Z(n15482) );
  NANDN U142 ( .A(n15766), .B(n2173), .Z(n91) );
  NANDN U143 ( .A(n15745), .B(n2174), .Z(n92) );
  AND U144 ( .A(n91), .B(n92), .Z(n15772) );
  NANDN U145 ( .A(n16060), .B(n2173), .Z(n93) );
  NANDN U146 ( .A(n16039), .B(n2174), .Z(n94) );
  AND U147 ( .A(n93), .B(n94), .Z(n16066) );
  NANDN U148 ( .A(n16354), .B(n2173), .Z(n95) );
  NANDN U149 ( .A(n16333), .B(n2174), .Z(n96) );
  AND U150 ( .A(n95), .B(n96), .Z(n16360) );
  NANDN U151 ( .A(n16648), .B(n2173), .Z(n97) );
  NANDN U152 ( .A(n16627), .B(n2174), .Z(n98) );
  AND U153 ( .A(n97), .B(n98), .Z(n16654) );
  NANDN U154 ( .A(n16942), .B(n2173), .Z(n99) );
  NANDN U155 ( .A(n16921), .B(n2174), .Z(n100) );
  AND U156 ( .A(n99), .B(n100), .Z(n16948) );
  NANDN U157 ( .A(n17236), .B(n2173), .Z(n101) );
  NANDN U158 ( .A(n17215), .B(n2174), .Z(n102) );
  AND U159 ( .A(n101), .B(n102), .Z(n17242) );
  NANDN U160 ( .A(n17530), .B(n2173), .Z(n103) );
  NANDN U161 ( .A(n17509), .B(n2174), .Z(n104) );
  AND U162 ( .A(n103), .B(n104), .Z(n17536) );
  NANDN U163 ( .A(n17816), .B(n2173), .Z(n105) );
  NANDN U164 ( .A(n17795), .B(n2174), .Z(n106) );
  AND U165 ( .A(n105), .B(n106), .Z(n17822) );
  NANDN U166 ( .A(n18108), .B(n2173), .Z(n107) );
  NANDN U167 ( .A(n18089), .B(n2174), .Z(n108) );
  AND U168 ( .A(n107), .B(n108), .Z(n18115) );
  NANDN U169 ( .A(n18400), .B(n2173), .Z(n109) );
  NANDN U170 ( .A(n18379), .B(n2174), .Z(n110) );
  AND U171 ( .A(n109), .B(n110), .Z(n18406) );
  NANDN U172 ( .A(n18694), .B(n2173), .Z(n111) );
  NANDN U173 ( .A(n18673), .B(n2174), .Z(n112) );
  AND U174 ( .A(n111), .B(n112), .Z(n18700) );
  NANDN U175 ( .A(n18988), .B(n2173), .Z(n113) );
  NANDN U176 ( .A(n18967), .B(n2174), .Z(n114) );
  AND U177 ( .A(n113), .B(n114), .Z(n18994) );
  NANDN U178 ( .A(n19282), .B(n2173), .Z(n115) );
  NANDN U179 ( .A(n19261), .B(n2174), .Z(n116) );
  AND U180 ( .A(n115), .B(n116), .Z(n19288) );
  NANDN U181 ( .A(n19576), .B(n2173), .Z(n117) );
  NANDN U182 ( .A(n19555), .B(n2174), .Z(n118) );
  AND U183 ( .A(n117), .B(n118), .Z(n19582) );
  NANDN U184 ( .A(n19866), .B(n2173), .Z(n119) );
  NANDN U185 ( .A(n19845), .B(n2174), .Z(n120) );
  AND U186 ( .A(n119), .B(n120), .Z(n19872) );
  NANDN U187 ( .A(n20156), .B(n2173), .Z(n121) );
  NANDN U188 ( .A(n20137), .B(n2174), .Z(n122) );
  AND U189 ( .A(n121), .B(n122), .Z(n20162) );
  NANDN U190 ( .A(n20450), .B(n2173), .Z(n123) );
  NANDN U191 ( .A(n20429), .B(n2174), .Z(n124) );
  AND U192 ( .A(n123), .B(n124), .Z(n20456) );
  NANDN U193 ( .A(n20744), .B(n2173), .Z(n125) );
  NANDN U194 ( .A(n20723), .B(n2174), .Z(n126) );
  AND U195 ( .A(n125), .B(n126), .Z(n20750) );
  NANDN U196 ( .A(n21036), .B(n2173), .Z(n127) );
  NANDN U197 ( .A(n21017), .B(n2174), .Z(n128) );
  AND U198 ( .A(n127), .B(n128), .Z(n21043) );
  NANDN U199 ( .A(n21324), .B(n2173), .Z(n129) );
  NANDN U200 ( .A(n21303), .B(n2174), .Z(n130) );
  AND U201 ( .A(n129), .B(n130), .Z(n21330) );
  NANDN U202 ( .A(n21618), .B(n2173), .Z(n131) );
  NANDN U203 ( .A(n21597), .B(n2174), .Z(n132) );
  AND U204 ( .A(n131), .B(n132), .Z(n21624) );
  NANDN U205 ( .A(n21912), .B(n2173), .Z(n133) );
  NANDN U206 ( .A(n21891), .B(n2174), .Z(n134) );
  AND U207 ( .A(n133), .B(n134), .Z(n21918) );
  NANDN U208 ( .A(n22206), .B(n2173), .Z(n135) );
  NANDN U209 ( .A(n22185), .B(n2174), .Z(n136) );
  AND U210 ( .A(n135), .B(n136), .Z(n22212) );
  NANDN U211 ( .A(n22496), .B(n2173), .Z(n137) );
  NANDN U212 ( .A(n22475), .B(n2174), .Z(n138) );
  AND U213 ( .A(n137), .B(n138), .Z(n22502) );
  NANDN U214 ( .A(n22790), .B(n2173), .Z(n139) );
  NANDN U215 ( .A(n22769), .B(n2174), .Z(n140) );
  AND U216 ( .A(n139), .B(n140), .Z(n22796) );
  NANDN U217 ( .A(n23084), .B(n2173), .Z(n141) );
  NANDN U218 ( .A(n23063), .B(n2174), .Z(n142) );
  AND U219 ( .A(n141), .B(n142), .Z(n23090) );
  NANDN U220 ( .A(n23378), .B(n2173), .Z(n143) );
  NANDN U221 ( .A(n23357), .B(n2174), .Z(n144) );
  AND U222 ( .A(n143), .B(n144), .Z(n23384) );
  NANDN U223 ( .A(n2457), .B(n2173), .Z(n145) );
  NANDN U224 ( .A(n2436), .B(n2174), .Z(n146) );
  AND U225 ( .A(n145), .B(n146), .Z(n2463) );
  NANDN U226 ( .A(n2751), .B(n2173), .Z(n147) );
  NANDN U227 ( .A(n2730), .B(n2174), .Z(n148) );
  AND U228 ( .A(n147), .B(n148), .Z(n2757) );
  NANDN U229 ( .A(n3045), .B(n2173), .Z(n149) );
  NANDN U230 ( .A(n3024), .B(n2174), .Z(n150) );
  AND U231 ( .A(n149), .B(n150), .Z(n3051) );
  NANDN U232 ( .A(n3339), .B(n2173), .Z(n151) );
  NANDN U233 ( .A(n3318), .B(n2174), .Z(n152) );
  AND U234 ( .A(n151), .B(n152), .Z(n3345) );
  NANDN U235 ( .A(n3633), .B(n2173), .Z(n153) );
  NANDN U236 ( .A(n3612), .B(n2174), .Z(n154) );
  AND U237 ( .A(n153), .B(n154), .Z(n3639) );
  NANDN U238 ( .A(n3927), .B(n2173), .Z(n155) );
  NANDN U239 ( .A(n3906), .B(n2174), .Z(n156) );
  AND U240 ( .A(n155), .B(n156), .Z(n3933) );
  NANDN U241 ( .A(n4221), .B(n2173), .Z(n157) );
  NANDN U242 ( .A(n4200), .B(n2174), .Z(n158) );
  AND U243 ( .A(n157), .B(n158), .Z(n4227) );
  NANDN U244 ( .A(n4511), .B(n2173), .Z(n159) );
  NANDN U245 ( .A(n4490), .B(n2174), .Z(n160) );
  AND U246 ( .A(n159), .B(n160), .Z(n4517) );
  NANDN U247 ( .A(n4805), .B(n2173), .Z(n161) );
  NANDN U248 ( .A(n4784), .B(n2174), .Z(n162) );
  AND U249 ( .A(n161), .B(n162), .Z(n4811) );
  NANDN U250 ( .A(n5099), .B(n2173), .Z(n163) );
  NANDN U251 ( .A(n5078), .B(n2174), .Z(n164) );
  AND U252 ( .A(n163), .B(n164), .Z(n5105) );
  NANDN U253 ( .A(n5393), .B(n2173), .Z(n165) );
  NANDN U254 ( .A(n5372), .B(n2174), .Z(n166) );
  AND U255 ( .A(n165), .B(n166), .Z(n5399) );
  NANDN U256 ( .A(n5687), .B(n2173), .Z(n167) );
  NANDN U257 ( .A(n5666), .B(n2174), .Z(n168) );
  AND U258 ( .A(n167), .B(n168), .Z(n5693) );
  NANDN U259 ( .A(n5981), .B(n2173), .Z(n169) );
  NANDN U260 ( .A(n5960), .B(n2174), .Z(n170) );
  AND U261 ( .A(n169), .B(n170), .Z(n5987) );
  NANDN U262 ( .A(n6275), .B(n2173), .Z(n171) );
  NANDN U263 ( .A(n6254), .B(n2174), .Z(n172) );
  AND U264 ( .A(n171), .B(n172), .Z(n6281) );
  NANDN U265 ( .A(n6565), .B(n2173), .Z(n173) );
  NANDN U266 ( .A(n6544), .B(n2174), .Z(n174) );
  AND U267 ( .A(n173), .B(n174), .Z(n6571) );
  NANDN U268 ( .A(n6855), .B(n2173), .Z(n175) );
  NANDN U269 ( .A(n6836), .B(n2174), .Z(n176) );
  AND U270 ( .A(n175), .B(n176), .Z(n6861) );
  NANDN U271 ( .A(n7141), .B(n2173), .Z(n177) );
  NANDN U272 ( .A(n7120), .B(n2174), .Z(n178) );
  AND U273 ( .A(n177), .B(n178), .Z(n7147) );
  NANDN U274 ( .A(n7435), .B(n2173), .Z(n179) );
  NANDN U275 ( .A(n7414), .B(n2174), .Z(n180) );
  AND U276 ( .A(n179), .B(n180), .Z(n7441) );
  NANDN U277 ( .A(n7725), .B(n2173), .Z(n181) );
  NANDN U278 ( .A(n7704), .B(n2174), .Z(n182) );
  AND U279 ( .A(n181), .B(n182), .Z(n7731) );
  NANDN U280 ( .A(n8011), .B(n2173), .Z(n183) );
  NANDN U281 ( .A(n7990), .B(n2174), .Z(n184) );
  AND U282 ( .A(n183), .B(n184), .Z(n8017) );
  NANDN U283 ( .A(n8301), .B(n2173), .Z(n185) );
  NANDN U284 ( .A(n8280), .B(n2174), .Z(n186) );
  AND U285 ( .A(n185), .B(n186), .Z(n8307) );
  NANDN U286 ( .A(n8595), .B(n2173), .Z(n187) );
  NANDN U287 ( .A(n8574), .B(n2174), .Z(n188) );
  AND U288 ( .A(n187), .B(n188), .Z(n8601) );
  NANDN U289 ( .A(n8889), .B(n2173), .Z(n189) );
  NANDN U290 ( .A(n8868), .B(n2174), .Z(n190) );
  AND U291 ( .A(n189), .B(n190), .Z(n8895) );
  NANDN U292 ( .A(n9179), .B(n2173), .Z(n191) );
  NANDN U293 ( .A(n9158), .B(n2174), .Z(n192) );
  AND U294 ( .A(n191), .B(n192), .Z(n9185) );
  NANDN U295 ( .A(n9469), .B(n2173), .Z(n193) );
  NANDN U296 ( .A(n9448), .B(n2174), .Z(n194) );
  AND U297 ( .A(n193), .B(n194), .Z(n9475) );
  NANDN U298 ( .A(n9763), .B(n2173), .Z(n195) );
  NANDN U299 ( .A(n9742), .B(n2174), .Z(n196) );
  AND U300 ( .A(n195), .B(n196), .Z(n9769) );
  NANDN U301 ( .A(n10057), .B(n2173), .Z(n197) );
  NANDN U302 ( .A(n10036), .B(n2174), .Z(n198) );
  AND U303 ( .A(n197), .B(n198), .Z(n10063) );
  NANDN U304 ( .A(n10351), .B(n2173), .Z(n199) );
  NANDN U305 ( .A(n10330), .B(n2174), .Z(n200) );
  AND U306 ( .A(n199), .B(n200), .Z(n10357) );
  NANDN U307 ( .A(n10645), .B(n2173), .Z(n201) );
  NANDN U308 ( .A(n10624), .B(n2174), .Z(n202) );
  AND U309 ( .A(n201), .B(n202), .Z(n10651) );
  NANDN U310 ( .A(n10939), .B(n2173), .Z(n203) );
  NANDN U311 ( .A(n10918), .B(n2174), .Z(n204) );
  AND U312 ( .A(n203), .B(n204), .Z(n10945) );
  NANDN U313 ( .A(n11233), .B(n2173), .Z(n205) );
  NANDN U314 ( .A(n11212), .B(n2174), .Z(n206) );
  AND U315 ( .A(n205), .B(n206), .Z(n11239) );
  NANDN U316 ( .A(n11527), .B(n2173), .Z(n207) );
  NANDN U317 ( .A(n11506), .B(n2174), .Z(n208) );
  AND U318 ( .A(n207), .B(n208), .Z(n11533) );
  NANDN U319 ( .A(n11813), .B(n2173), .Z(n209) );
  NANDN U320 ( .A(n11794), .B(n2174), .Z(n210) );
  AND U321 ( .A(n209), .B(n210), .Z(n11819) );
  NANDN U322 ( .A(n12107), .B(n2173), .Z(n211) );
  NANDN U323 ( .A(n12086), .B(n2174), .Z(n212) );
  AND U324 ( .A(n211), .B(n212), .Z(n12113) );
  NANDN U325 ( .A(n12401), .B(n2173), .Z(n213) );
  NANDN U326 ( .A(n12380), .B(n2174), .Z(n214) );
  AND U327 ( .A(n213), .B(n214), .Z(n12407) );
  NANDN U328 ( .A(n12691), .B(n2173), .Z(n215) );
  NANDN U329 ( .A(n12670), .B(n2174), .Z(n216) );
  AND U330 ( .A(n215), .B(n216), .Z(n12697) );
  NANDN U331 ( .A(n12985), .B(n2173), .Z(n217) );
  NANDN U332 ( .A(n12964), .B(n2174), .Z(n218) );
  AND U333 ( .A(n217), .B(n218), .Z(n12991) );
  NANDN U334 ( .A(n13279), .B(n2173), .Z(n219) );
  NANDN U335 ( .A(n13258), .B(n2174), .Z(n220) );
  AND U336 ( .A(n219), .B(n220), .Z(n13285) );
  NANDN U337 ( .A(n13573), .B(n2173), .Z(n221) );
  NANDN U338 ( .A(n13552), .B(n2174), .Z(n222) );
  AND U339 ( .A(n221), .B(n222), .Z(n13579) );
  NANDN U340 ( .A(n13863), .B(n2173), .Z(n223) );
  NANDN U341 ( .A(n13842), .B(n2174), .Z(n224) );
  AND U342 ( .A(n223), .B(n224), .Z(n13869) );
  NANDN U343 ( .A(n14157), .B(n2173), .Z(n225) );
  NANDN U344 ( .A(n14136), .B(n2174), .Z(n226) );
  AND U345 ( .A(n225), .B(n226), .Z(n14163) );
  NANDN U346 ( .A(n14451), .B(n2173), .Z(n227) );
  NANDN U347 ( .A(n14430), .B(n2174), .Z(n228) );
  AND U348 ( .A(n227), .B(n228), .Z(n14457) );
  NANDN U349 ( .A(n14745), .B(n2173), .Z(n229) );
  NANDN U350 ( .A(n14724), .B(n2174), .Z(n230) );
  AND U351 ( .A(n229), .B(n230), .Z(n14751) );
  NANDN U352 ( .A(n15035), .B(n2173), .Z(n231) );
  NANDN U353 ( .A(n15014), .B(n2174), .Z(n232) );
  AND U354 ( .A(n231), .B(n232), .Z(n15041) );
  NANDN U355 ( .A(n15329), .B(n2173), .Z(n233) );
  NANDN U356 ( .A(n15308), .B(n2174), .Z(n234) );
  AND U357 ( .A(n233), .B(n234), .Z(n15335) );
  NANDN U358 ( .A(n15621), .B(n2173), .Z(n235) );
  NANDN U359 ( .A(n15602), .B(n2174), .Z(n236) );
  AND U360 ( .A(n235), .B(n236), .Z(n15628) );
  NANDN U361 ( .A(n15913), .B(n2173), .Z(n237) );
  NANDN U362 ( .A(n15892), .B(n2174), .Z(n238) );
  AND U363 ( .A(n237), .B(n238), .Z(n15919) );
  NANDN U364 ( .A(n16207), .B(n2173), .Z(n239) );
  NANDN U365 ( .A(n16186), .B(n2174), .Z(n240) );
  AND U366 ( .A(n239), .B(n240), .Z(n16213) );
  NANDN U367 ( .A(n16501), .B(n2173), .Z(n241) );
  NANDN U368 ( .A(n16480), .B(n2174), .Z(n242) );
  AND U369 ( .A(n241), .B(n242), .Z(n16507) );
  NANDN U370 ( .A(n16795), .B(n2173), .Z(n243) );
  NANDN U371 ( .A(n16774), .B(n2174), .Z(n244) );
  AND U372 ( .A(n243), .B(n244), .Z(n16801) );
  NANDN U373 ( .A(n17089), .B(n2173), .Z(n245) );
  NANDN U374 ( .A(n17068), .B(n2174), .Z(n246) );
  AND U375 ( .A(n245), .B(n246), .Z(n17095) );
  NANDN U376 ( .A(n17383), .B(n2173), .Z(n247) );
  NANDN U377 ( .A(n17362), .B(n2174), .Z(n248) );
  AND U378 ( .A(n247), .B(n248), .Z(n17389) );
  NANDN U379 ( .A(n17677), .B(n2173), .Z(n249) );
  NANDN U380 ( .A(n17656), .B(n2174), .Z(n250) );
  AND U381 ( .A(n249), .B(n250), .Z(n17683) );
  NANDN U382 ( .A(n17963), .B(n2173), .Z(n251) );
  NANDN U383 ( .A(n17942), .B(n2174), .Z(n252) );
  AND U384 ( .A(n251), .B(n252), .Z(n17969) );
  NANDN U385 ( .A(n18253), .B(n2173), .Z(n253) );
  NANDN U386 ( .A(n18232), .B(n2174), .Z(n254) );
  AND U387 ( .A(n253), .B(n254), .Z(n18259) );
  NANDN U388 ( .A(n18547), .B(n2173), .Z(n255) );
  NANDN U389 ( .A(n18526), .B(n2174), .Z(n256) );
  AND U390 ( .A(n255), .B(n256), .Z(n18553) );
  NANDN U391 ( .A(n18841), .B(n2173), .Z(n257) );
  NANDN U392 ( .A(n18820), .B(n2174), .Z(n258) );
  AND U393 ( .A(n257), .B(n258), .Z(n18847) );
  NANDN U394 ( .A(n19135), .B(n2173), .Z(n259) );
  NANDN U395 ( .A(n19114), .B(n2174), .Z(n260) );
  AND U396 ( .A(n259), .B(n260), .Z(n19141) );
  NANDN U397 ( .A(n19429), .B(n2173), .Z(n261) );
  NANDN U398 ( .A(n19408), .B(n2174), .Z(n262) );
  AND U399 ( .A(n261), .B(n262), .Z(n19435) );
  NANDN U400 ( .A(n19719), .B(n2173), .Z(n263) );
  NANDN U401 ( .A(n19700), .B(n2174), .Z(n264) );
  AND U402 ( .A(n263), .B(n264), .Z(n19725) );
  NANDN U403 ( .A(n20013), .B(n2173), .Z(n265) );
  NANDN U404 ( .A(n19992), .B(n2174), .Z(n266) );
  AND U405 ( .A(n265), .B(n266), .Z(n20019) );
  NANDN U406 ( .A(n20303), .B(n2173), .Z(n267) );
  NANDN U407 ( .A(n20282), .B(n2174), .Z(n268) );
  AND U408 ( .A(n267), .B(n268), .Z(n20309) );
  NANDN U409 ( .A(n20597), .B(n2173), .Z(n269) );
  NANDN U410 ( .A(n20576), .B(n2174), .Z(n270) );
  AND U411 ( .A(n269), .B(n270), .Z(n20603) );
  NANDN U412 ( .A(n20891), .B(n2173), .Z(n271) );
  NANDN U413 ( .A(n20870), .B(n2174), .Z(n272) );
  AND U414 ( .A(n271), .B(n272), .Z(n20897) );
  NANDN U415 ( .A(n21181), .B(n2173), .Z(n273) );
  NANDN U416 ( .A(n21160), .B(n2174), .Z(n274) );
  AND U417 ( .A(n273), .B(n274), .Z(n21187) );
  NANDN U418 ( .A(n21471), .B(n2173), .Z(n275) );
  NANDN U419 ( .A(n21450), .B(n2174), .Z(n276) );
  AND U420 ( .A(n275), .B(n276), .Z(n21477) );
  NANDN U421 ( .A(n21765), .B(n2173), .Z(n277) );
  NANDN U422 ( .A(n21744), .B(n2174), .Z(n278) );
  AND U423 ( .A(n277), .B(n278), .Z(n21771) );
  NANDN U424 ( .A(n22059), .B(n2173), .Z(n279) );
  NANDN U425 ( .A(n22038), .B(n2174), .Z(n280) );
  AND U426 ( .A(n279), .B(n280), .Z(n22065) );
  NANDN U427 ( .A(n22349), .B(n2173), .Z(n281) );
  NANDN U428 ( .A(n22330), .B(n2174), .Z(n282) );
  AND U429 ( .A(n281), .B(n282), .Z(n22355) );
  NANDN U430 ( .A(n22643), .B(n2173), .Z(n283) );
  NANDN U431 ( .A(n22622), .B(n2174), .Z(n284) );
  AND U432 ( .A(n283), .B(n284), .Z(n22649) );
  NANDN U433 ( .A(n22937), .B(n2173), .Z(n285) );
  NANDN U434 ( .A(n22916), .B(n2174), .Z(n286) );
  AND U435 ( .A(n285), .B(n286), .Z(n22943) );
  NANDN U436 ( .A(n23231), .B(n2173), .Z(n287) );
  NANDN U437 ( .A(n23210), .B(n2174), .Z(n288) );
  AND U438 ( .A(n287), .B(n288), .Z(n23237) );
  NANDN U439 ( .A(n23525), .B(n2173), .Z(n289) );
  NANDN U440 ( .A(n23504), .B(n2174), .Z(n290) );
  AND U441 ( .A(n289), .B(n290), .Z(n23531) );
  NANDN U442 ( .A(n2478), .B(n2173), .Z(n291) );
  NANDN U443 ( .A(n2457), .B(n2174), .Z(n292) );
  AND U444 ( .A(n291), .B(n292), .Z(n2484) );
  NANDN U445 ( .A(n2625), .B(n2173), .Z(n293) );
  NANDN U446 ( .A(n2604), .B(n2174), .Z(n294) );
  AND U447 ( .A(n293), .B(n294), .Z(n2631) );
  NANDN U448 ( .A(n2772), .B(n2173), .Z(n295) );
  NANDN U449 ( .A(n2751), .B(n2174), .Z(n296) );
  AND U450 ( .A(n295), .B(n296), .Z(n2778) );
  NANDN U451 ( .A(n2919), .B(n2173), .Z(n297) );
  NANDN U452 ( .A(n2898), .B(n2174), .Z(n298) );
  AND U453 ( .A(n297), .B(n298), .Z(n2925) );
  NANDN U454 ( .A(n3066), .B(n2173), .Z(n299) );
  NANDN U455 ( .A(n3045), .B(n2174), .Z(n300) );
  AND U456 ( .A(n299), .B(n300), .Z(n3072) );
  NANDN U457 ( .A(n3213), .B(n2173), .Z(n301) );
  NANDN U458 ( .A(n3192), .B(n2174), .Z(n302) );
  AND U459 ( .A(n301), .B(n302), .Z(n3219) );
  NANDN U460 ( .A(n3360), .B(n2173), .Z(n303) );
  NANDN U461 ( .A(n3339), .B(n2174), .Z(n304) );
  AND U462 ( .A(n303), .B(n304), .Z(n3366) );
  NANDN U463 ( .A(n3507), .B(n2173), .Z(n305) );
  NANDN U464 ( .A(n3486), .B(n2174), .Z(n306) );
  AND U465 ( .A(n305), .B(n306), .Z(n3513) );
  NANDN U466 ( .A(n3654), .B(n2173), .Z(n307) );
  NANDN U467 ( .A(n3633), .B(n2174), .Z(n308) );
  AND U468 ( .A(n307), .B(n308), .Z(n3660) );
  NANDN U469 ( .A(n3801), .B(n2173), .Z(n309) );
  NANDN U470 ( .A(n3780), .B(n2174), .Z(n310) );
  AND U471 ( .A(n309), .B(n310), .Z(n3807) );
  NANDN U472 ( .A(n3948), .B(n2173), .Z(n311) );
  NANDN U473 ( .A(n3927), .B(n2174), .Z(n312) );
  AND U474 ( .A(n311), .B(n312), .Z(n3954) );
  NANDN U475 ( .A(n4095), .B(n2173), .Z(n313) );
  NANDN U476 ( .A(n4074), .B(n2174), .Z(n314) );
  AND U477 ( .A(n313), .B(n314), .Z(n4101) );
  NANDN U478 ( .A(n4242), .B(n2173), .Z(n315) );
  NANDN U479 ( .A(n4221), .B(n2174), .Z(n316) );
  AND U480 ( .A(n315), .B(n316), .Z(n4248) );
  NANDN U481 ( .A(n4389), .B(n2173), .Z(n317) );
  NANDN U482 ( .A(n4368), .B(n2174), .Z(n318) );
  AND U483 ( .A(n317), .B(n318), .Z(n4395) );
  NANDN U484 ( .A(n4532), .B(n2173), .Z(n319) );
  NANDN U485 ( .A(n4511), .B(n2174), .Z(n320) );
  AND U486 ( .A(n319), .B(n320), .Z(n4538) );
  NANDN U487 ( .A(n4679), .B(n2173), .Z(n321) );
  NANDN U488 ( .A(n4658), .B(n2174), .Z(n322) );
  AND U489 ( .A(n321), .B(n322), .Z(n4685) );
  NANDN U490 ( .A(n4826), .B(n2173), .Z(n323) );
  NANDN U491 ( .A(n4805), .B(n2174), .Z(n324) );
  AND U492 ( .A(n323), .B(n324), .Z(n4832) );
  NANDN U493 ( .A(n4973), .B(n2173), .Z(n325) );
  NANDN U494 ( .A(n4952), .B(n2174), .Z(n326) );
  AND U495 ( .A(n325), .B(n326), .Z(n4979) );
  NANDN U496 ( .A(n5120), .B(n2173), .Z(n327) );
  NANDN U497 ( .A(n5099), .B(n2174), .Z(n328) );
  AND U498 ( .A(n327), .B(n328), .Z(n5126) );
  NANDN U499 ( .A(n5267), .B(n2173), .Z(n329) );
  NANDN U500 ( .A(n5246), .B(n2174), .Z(n330) );
  AND U501 ( .A(n329), .B(n330), .Z(n5273) );
  NANDN U502 ( .A(n5414), .B(n2173), .Z(n331) );
  NANDN U503 ( .A(n5393), .B(n2174), .Z(n332) );
  AND U504 ( .A(n331), .B(n332), .Z(n5420) );
  NANDN U505 ( .A(n5561), .B(n2173), .Z(n333) );
  NANDN U506 ( .A(n5540), .B(n2174), .Z(n334) );
  AND U507 ( .A(n333), .B(n334), .Z(n5567) );
  NANDN U508 ( .A(n5708), .B(n2173), .Z(n335) );
  NANDN U509 ( .A(n5687), .B(n2174), .Z(n336) );
  AND U510 ( .A(n335), .B(n336), .Z(n5714) );
  NANDN U511 ( .A(n5855), .B(n2173), .Z(n337) );
  NANDN U512 ( .A(n5834), .B(n2174), .Z(n338) );
  AND U513 ( .A(n337), .B(n338), .Z(n5861) );
  NANDN U514 ( .A(n6002), .B(n2173), .Z(n339) );
  NANDN U515 ( .A(n5981), .B(n2174), .Z(n340) );
  AND U516 ( .A(n339), .B(n340), .Z(n6008) );
  NANDN U517 ( .A(n6149), .B(n2173), .Z(n341) );
  NANDN U518 ( .A(n6128), .B(n2174), .Z(n342) );
  AND U519 ( .A(n341), .B(n342), .Z(n6155) );
  NANDN U520 ( .A(n6296), .B(n2173), .Z(n343) );
  NANDN U521 ( .A(n6275), .B(n2174), .Z(n344) );
  AND U522 ( .A(n343), .B(n344), .Z(n6302) );
  NANDN U523 ( .A(n6439), .B(n2173), .Z(n345) );
  NANDN U524 ( .A(n6420), .B(n2174), .Z(n346) );
  AND U525 ( .A(n345), .B(n346), .Z(n6445) );
  NANDN U526 ( .A(n6586), .B(n2173), .Z(n347) );
  NANDN U527 ( .A(n6565), .B(n2174), .Z(n348) );
  AND U528 ( .A(n347), .B(n348), .Z(n6592) );
  NANDN U529 ( .A(n6733), .B(n2173), .Z(n349) );
  NANDN U530 ( .A(n6712), .B(n2174), .Z(n350) );
  AND U531 ( .A(n349), .B(n350), .Z(n6739) );
  NANDN U532 ( .A(n6876), .B(n2173), .Z(n351) );
  NANDN U533 ( .A(n6855), .B(n2174), .Z(n352) );
  AND U534 ( .A(n351), .B(n352), .Z(n6882) );
  NANDN U535 ( .A(n7019), .B(n2173), .Z(n353) );
  NANDN U536 ( .A(n6998), .B(n2174), .Z(n354) );
  AND U537 ( .A(n353), .B(n354), .Z(n7025) );
  NANDN U538 ( .A(n7162), .B(n2173), .Z(n355) );
  NANDN U539 ( .A(n7141), .B(n2174), .Z(n356) );
  AND U540 ( .A(n355), .B(n356), .Z(n7168) );
  NANDN U541 ( .A(n7309), .B(n2173), .Z(n357) );
  NANDN U542 ( .A(n7288), .B(n2174), .Z(n358) );
  AND U543 ( .A(n357), .B(n358), .Z(n7315) );
  NANDN U544 ( .A(n7456), .B(n2173), .Z(n359) );
  NANDN U545 ( .A(n7435), .B(n2174), .Z(n360) );
  AND U546 ( .A(n359), .B(n360), .Z(n7462) );
  NANDN U547 ( .A(n7599), .B(n2173), .Z(n361) );
  NANDN U548 ( .A(n7578), .B(n2174), .Z(n362) );
  AND U549 ( .A(n361), .B(n362), .Z(n7605) );
  NANDN U550 ( .A(n7746), .B(n2173), .Z(n363) );
  NANDN U551 ( .A(n7725), .B(n2174), .Z(n364) );
  AND U552 ( .A(n363), .B(n364), .Z(n7752) );
  NANDN U553 ( .A(n7889), .B(n2173), .Z(n365) );
  NANDN U554 ( .A(n7868), .B(n2174), .Z(n366) );
  AND U555 ( .A(n365), .B(n366), .Z(n7895) );
  NANDN U556 ( .A(n8032), .B(n2173), .Z(n367) );
  NANDN U557 ( .A(n8011), .B(n2174), .Z(n368) );
  AND U558 ( .A(n367), .B(n368), .Z(n8038) );
  NANDN U559 ( .A(n8179), .B(n2173), .Z(n369) );
  NANDN U560 ( .A(n8158), .B(n2174), .Z(n370) );
  AND U561 ( .A(n369), .B(n370), .Z(n8185) );
  NANDN U562 ( .A(n8322), .B(n2173), .Z(n371) );
  NANDN U563 ( .A(n8301), .B(n2174), .Z(n372) );
  AND U564 ( .A(n371), .B(n372), .Z(n8328) );
  NANDN U565 ( .A(n8469), .B(n2173), .Z(n373) );
  NANDN U566 ( .A(n8448), .B(n2174), .Z(n374) );
  AND U567 ( .A(n373), .B(n374), .Z(n8475) );
  NANDN U568 ( .A(n8616), .B(n2173), .Z(n375) );
  NANDN U569 ( .A(n8595), .B(n2174), .Z(n376) );
  AND U570 ( .A(n375), .B(n376), .Z(n8622) );
  NANDN U571 ( .A(n8763), .B(n2173), .Z(n377) );
  NANDN U572 ( .A(n8742), .B(n2174), .Z(n378) );
  AND U573 ( .A(n377), .B(n378), .Z(n8769) );
  NANDN U574 ( .A(n8910), .B(n2173), .Z(n379) );
  NANDN U575 ( .A(n8889), .B(n2174), .Z(n380) );
  AND U576 ( .A(n379), .B(n380), .Z(n8916) );
  NANDN U577 ( .A(n9055), .B(n2173), .Z(n381) );
  NANDN U578 ( .A(n9036), .B(n2174), .Z(n382) );
  AND U579 ( .A(n381), .B(n382), .Z(n9062) );
  NANDN U580 ( .A(n9198), .B(n2173), .Z(n383) );
  NANDN U581 ( .A(n9179), .B(n2174), .Z(n384) );
  AND U582 ( .A(n383), .B(n384), .Z(n9205) );
  NANDN U583 ( .A(n9343), .B(n2173), .Z(n385) );
  NANDN U584 ( .A(n9322), .B(n2174), .Z(n386) );
  AND U585 ( .A(n385), .B(n386), .Z(n9349) );
  NANDN U586 ( .A(n9490), .B(n2173), .Z(n387) );
  NANDN U587 ( .A(n9469), .B(n2174), .Z(n388) );
  AND U588 ( .A(n387), .B(n388), .Z(n9496) );
  NANDN U589 ( .A(n9637), .B(n2173), .Z(n389) );
  NANDN U590 ( .A(n9616), .B(n2174), .Z(n390) );
  AND U591 ( .A(n389), .B(n390), .Z(n9643) );
  NANDN U592 ( .A(n9784), .B(n2173), .Z(n391) );
  NANDN U593 ( .A(n9763), .B(n2174), .Z(n392) );
  AND U594 ( .A(n391), .B(n392), .Z(n9790) );
  NANDN U595 ( .A(n9931), .B(n2173), .Z(n393) );
  NANDN U596 ( .A(n9910), .B(n2174), .Z(n394) );
  AND U597 ( .A(n393), .B(n394), .Z(n9937) );
  NANDN U598 ( .A(n10078), .B(n2173), .Z(n395) );
  NANDN U599 ( .A(n10057), .B(n2174), .Z(n396) );
  AND U600 ( .A(n395), .B(n396), .Z(n10084) );
  NANDN U601 ( .A(n10225), .B(n2173), .Z(n397) );
  NANDN U602 ( .A(n10204), .B(n2174), .Z(n398) );
  AND U603 ( .A(n397), .B(n398), .Z(n10231) );
  NANDN U604 ( .A(n10372), .B(n2173), .Z(n399) );
  NANDN U605 ( .A(n10351), .B(n2174), .Z(n400) );
  AND U606 ( .A(n399), .B(n400), .Z(n10378) );
  NANDN U607 ( .A(n10519), .B(n2173), .Z(n401) );
  NANDN U608 ( .A(n10498), .B(n2174), .Z(n402) );
  AND U609 ( .A(n401), .B(n402), .Z(n10525) );
  NANDN U610 ( .A(n10666), .B(n2173), .Z(n403) );
  NANDN U611 ( .A(n10645), .B(n2174), .Z(n404) );
  AND U612 ( .A(n403), .B(n404), .Z(n10672) );
  NANDN U613 ( .A(n10813), .B(n2173), .Z(n405) );
  NANDN U614 ( .A(n10792), .B(n2174), .Z(n406) );
  AND U615 ( .A(n405), .B(n406), .Z(n10819) );
  NANDN U616 ( .A(n10960), .B(n2173), .Z(n407) );
  NANDN U617 ( .A(n10939), .B(n2174), .Z(n408) );
  AND U618 ( .A(n407), .B(n408), .Z(n10966) );
  NANDN U619 ( .A(n11107), .B(n2173), .Z(n409) );
  NANDN U620 ( .A(n11086), .B(n2174), .Z(n410) );
  AND U621 ( .A(n409), .B(n410), .Z(n11113) );
  NANDN U622 ( .A(n11254), .B(n2173), .Z(n411) );
  NANDN U623 ( .A(n11233), .B(n2174), .Z(n412) );
  AND U624 ( .A(n411), .B(n412), .Z(n11260) );
  NANDN U625 ( .A(n11401), .B(n2173), .Z(n413) );
  NANDN U626 ( .A(n11380), .B(n2174), .Z(n414) );
  AND U627 ( .A(n413), .B(n414), .Z(n11407) );
  NANDN U628 ( .A(n11548), .B(n2173), .Z(n415) );
  NANDN U629 ( .A(n11527), .B(n2174), .Z(n416) );
  AND U630 ( .A(n415), .B(n416), .Z(n11554) );
  NANDN U631 ( .A(n11695), .B(n2173), .Z(n417) );
  NANDN U632 ( .A(n11674), .B(n2174), .Z(n418) );
  AND U633 ( .A(n417), .B(n418), .Z(n11701) );
  NANDN U634 ( .A(n11834), .B(n2173), .Z(n419) );
  NANDN U635 ( .A(n11813), .B(n2174), .Z(n420) );
  AND U636 ( .A(n419), .B(n420), .Z(n11840) );
  NANDN U637 ( .A(n11981), .B(n2173), .Z(n421) );
  NANDN U638 ( .A(n11960), .B(n2174), .Z(n422) );
  AND U639 ( .A(n421), .B(n422), .Z(n11987) );
  NANDN U640 ( .A(n12128), .B(n2173), .Z(n423) );
  NANDN U641 ( .A(n12107), .B(n2174), .Z(n424) );
  AND U642 ( .A(n423), .B(n424), .Z(n12134) );
  NANDN U643 ( .A(n12275), .B(n2173), .Z(n425) );
  NANDN U644 ( .A(n12254), .B(n2174), .Z(n426) );
  AND U645 ( .A(n425), .B(n426), .Z(n12281) );
  NANDN U646 ( .A(n12422), .B(n2173), .Z(n427) );
  NANDN U647 ( .A(n12401), .B(n2174), .Z(n428) );
  AND U648 ( .A(n427), .B(n428), .Z(n12428) );
  NANDN U649 ( .A(n12569), .B(n2173), .Z(n429) );
  NANDN U650 ( .A(n12548), .B(n2174), .Z(n430) );
  AND U651 ( .A(n429), .B(n430), .Z(n12575) );
  NANDN U652 ( .A(n12712), .B(n2173), .Z(n431) );
  NANDN U653 ( .A(n12691), .B(n2174), .Z(n432) );
  AND U654 ( .A(n431), .B(n432), .Z(n12718) );
  NANDN U655 ( .A(n12859), .B(n2173), .Z(n433) );
  NANDN U656 ( .A(n12838), .B(n2174), .Z(n434) );
  AND U657 ( .A(n433), .B(n434), .Z(n12865) );
  NANDN U658 ( .A(n13006), .B(n2173), .Z(n435) );
  NANDN U659 ( .A(n12985), .B(n2174), .Z(n436) );
  AND U660 ( .A(n435), .B(n436), .Z(n13012) );
  NANDN U661 ( .A(n13153), .B(n2173), .Z(n437) );
  NANDN U662 ( .A(n13132), .B(n2174), .Z(n438) );
  AND U663 ( .A(n437), .B(n438), .Z(n13159) );
  NANDN U664 ( .A(n13300), .B(n2173), .Z(n439) );
  NANDN U665 ( .A(n13279), .B(n2174), .Z(n440) );
  AND U666 ( .A(n439), .B(n440), .Z(n13306) );
  NANDN U667 ( .A(n13447), .B(n2173), .Z(n441) );
  NANDN U668 ( .A(n13426), .B(n2174), .Z(n442) );
  AND U669 ( .A(n441), .B(n442), .Z(n13453) );
  NANDN U670 ( .A(n13594), .B(n2173), .Z(n443) );
  NANDN U671 ( .A(n13573), .B(n2174), .Z(n444) );
  AND U672 ( .A(n443), .B(n444), .Z(n13600) );
  NANDN U673 ( .A(n13741), .B(n2173), .Z(n445) );
  NANDN U674 ( .A(n13720), .B(n2174), .Z(n446) );
  AND U675 ( .A(n445), .B(n446), .Z(n13747) );
  NANDN U676 ( .A(n13884), .B(n2173), .Z(n447) );
  NANDN U677 ( .A(n13863), .B(n2174), .Z(n448) );
  AND U678 ( .A(n447), .B(n448), .Z(n13890) );
  NANDN U679 ( .A(n14031), .B(n2173), .Z(n449) );
  NANDN U680 ( .A(n14010), .B(n2174), .Z(n450) );
  AND U681 ( .A(n449), .B(n450), .Z(n14037) );
  NANDN U682 ( .A(n14178), .B(n2173), .Z(n451) );
  NANDN U683 ( .A(n14157), .B(n2174), .Z(n452) );
  AND U684 ( .A(n451), .B(n452), .Z(n14184) );
  NANDN U685 ( .A(n14325), .B(n2173), .Z(n453) );
  NANDN U686 ( .A(n14304), .B(n2174), .Z(n454) );
  AND U687 ( .A(n453), .B(n454), .Z(n14331) );
  NANDN U688 ( .A(n14472), .B(n2173), .Z(n455) );
  NANDN U689 ( .A(n14451), .B(n2174), .Z(n456) );
  AND U690 ( .A(n455), .B(n456), .Z(n14478) );
  NANDN U691 ( .A(n14619), .B(n2173), .Z(n457) );
  NANDN U692 ( .A(n14598), .B(n2174), .Z(n458) );
  AND U693 ( .A(n457), .B(n458), .Z(n14625) );
  NANDN U694 ( .A(n14764), .B(n2173), .Z(n459) );
  NANDN U695 ( .A(n14745), .B(n2174), .Z(n460) );
  AND U696 ( .A(n459), .B(n460), .Z(n14771) );
  NANDN U697 ( .A(n14909), .B(n2173), .Z(n461) );
  NANDN U698 ( .A(n14888), .B(n2174), .Z(n462) );
  AND U699 ( .A(n461), .B(n462), .Z(n14915) );
  NANDN U700 ( .A(n15056), .B(n2173), .Z(n463) );
  NANDN U701 ( .A(n15035), .B(n2174), .Z(n464) );
  AND U702 ( .A(n463), .B(n464), .Z(n15062) );
  NANDN U703 ( .A(n15203), .B(n2173), .Z(n465) );
  NANDN U704 ( .A(n15182), .B(n2174), .Z(n466) );
  AND U705 ( .A(n465), .B(n466), .Z(n15209) );
  NANDN U706 ( .A(n15350), .B(n2173), .Z(n467) );
  NANDN U707 ( .A(n15329), .B(n2174), .Z(n468) );
  AND U708 ( .A(n467), .B(n468), .Z(n15356) );
  NANDN U709 ( .A(n15497), .B(n2173), .Z(n469) );
  NANDN U710 ( .A(n15476), .B(n2174), .Z(n470) );
  AND U711 ( .A(n469), .B(n470), .Z(n15503) );
  NANDN U712 ( .A(n15640), .B(n2173), .Z(n471) );
  NANDN U713 ( .A(n15621), .B(n2174), .Z(n472) );
  AND U714 ( .A(n471), .B(n472), .Z(n15646) );
  NANDN U715 ( .A(n15787), .B(n2173), .Z(n473) );
  NANDN U716 ( .A(n15766), .B(n2174), .Z(n474) );
  AND U717 ( .A(n473), .B(n474), .Z(n15793) );
  NANDN U718 ( .A(n15934), .B(n2173), .Z(n475) );
  NANDN U719 ( .A(n15913), .B(n2174), .Z(n476) );
  AND U720 ( .A(n475), .B(n476), .Z(n15940) );
  NANDN U721 ( .A(n16081), .B(n2173), .Z(n477) );
  NANDN U722 ( .A(n16060), .B(n2174), .Z(n478) );
  AND U723 ( .A(n477), .B(n478), .Z(n16087) );
  NANDN U724 ( .A(n16228), .B(n2173), .Z(n479) );
  NANDN U725 ( .A(n16207), .B(n2174), .Z(n480) );
  AND U726 ( .A(n479), .B(n480), .Z(n16234) );
  NANDN U727 ( .A(n16375), .B(n2173), .Z(n481) );
  NANDN U728 ( .A(n16354), .B(n2174), .Z(n482) );
  AND U729 ( .A(n481), .B(n482), .Z(n16381) );
  NANDN U730 ( .A(n16522), .B(n2173), .Z(n483) );
  NANDN U731 ( .A(n16501), .B(n2174), .Z(n484) );
  AND U732 ( .A(n483), .B(n484), .Z(n16528) );
  NANDN U733 ( .A(n16669), .B(n2173), .Z(n485) );
  NANDN U734 ( .A(n16648), .B(n2174), .Z(n486) );
  AND U735 ( .A(n485), .B(n486), .Z(n16675) );
  NANDN U736 ( .A(n16816), .B(n2173), .Z(n487) );
  NANDN U737 ( .A(n16795), .B(n2174), .Z(n488) );
  AND U738 ( .A(n487), .B(n488), .Z(n16822) );
  NANDN U739 ( .A(n16963), .B(n2173), .Z(n489) );
  NANDN U740 ( .A(n16942), .B(n2174), .Z(n490) );
  AND U741 ( .A(n489), .B(n490), .Z(n16969) );
  NANDN U742 ( .A(n17110), .B(n2173), .Z(n491) );
  NANDN U743 ( .A(n17089), .B(n2174), .Z(n492) );
  AND U744 ( .A(n491), .B(n492), .Z(n17116) );
  NANDN U745 ( .A(n17257), .B(n2173), .Z(n493) );
  NANDN U746 ( .A(n17236), .B(n2174), .Z(n494) );
  AND U747 ( .A(n493), .B(n494), .Z(n17263) );
  NANDN U748 ( .A(n17404), .B(n2173), .Z(n495) );
  NANDN U749 ( .A(n17383), .B(n2174), .Z(n496) );
  AND U750 ( .A(n495), .B(n496), .Z(n17410) );
  NANDN U751 ( .A(n17551), .B(n2173), .Z(n497) );
  NANDN U752 ( .A(n17530), .B(n2174), .Z(n498) );
  AND U753 ( .A(n497), .B(n498), .Z(n17557) );
  NANDN U754 ( .A(n17698), .B(n2173), .Z(n499) );
  NANDN U755 ( .A(n17677), .B(n2174), .Z(n500) );
  AND U756 ( .A(n499), .B(n500), .Z(n17704) );
  NANDN U757 ( .A(n17837), .B(n2173), .Z(n501) );
  NANDN U758 ( .A(n17816), .B(n2174), .Z(n502) );
  AND U759 ( .A(n501), .B(n502), .Z(n17843) );
  NANDN U760 ( .A(n17984), .B(n2173), .Z(n503) );
  NANDN U761 ( .A(n17963), .B(n2174), .Z(n504) );
  AND U762 ( .A(n503), .B(n504), .Z(n17990) );
  NANDN U763 ( .A(n18127), .B(n2173), .Z(n505) );
  NANDN U764 ( .A(n18108), .B(n2174), .Z(n506) );
  AND U765 ( .A(n505), .B(n506), .Z(n18133) );
  NANDN U766 ( .A(n18274), .B(n2173), .Z(n507) );
  NANDN U767 ( .A(n18253), .B(n2174), .Z(n508) );
  AND U768 ( .A(n507), .B(n508), .Z(n18280) );
  NANDN U769 ( .A(n18421), .B(n2173), .Z(n509) );
  NANDN U770 ( .A(n18400), .B(n2174), .Z(n510) );
  AND U771 ( .A(n509), .B(n510), .Z(n18427) );
  NANDN U772 ( .A(n18568), .B(n2173), .Z(n511) );
  NANDN U773 ( .A(n18547), .B(n2174), .Z(n512) );
  AND U774 ( .A(n511), .B(n512), .Z(n18574) );
  NANDN U775 ( .A(n18715), .B(n2173), .Z(n513) );
  NANDN U776 ( .A(n18694), .B(n2174), .Z(n514) );
  AND U777 ( .A(n513), .B(n514), .Z(n18721) );
  NANDN U778 ( .A(n18862), .B(n2173), .Z(n515) );
  NANDN U779 ( .A(n18841), .B(n2174), .Z(n516) );
  AND U780 ( .A(n515), .B(n516), .Z(n18868) );
  NANDN U781 ( .A(n19009), .B(n2173), .Z(n517) );
  NANDN U782 ( .A(n18988), .B(n2174), .Z(n518) );
  AND U783 ( .A(n517), .B(n518), .Z(n19015) );
  NANDN U784 ( .A(n19156), .B(n2173), .Z(n519) );
  NANDN U785 ( .A(n19135), .B(n2174), .Z(n520) );
  AND U786 ( .A(n519), .B(n520), .Z(n19162) );
  NANDN U787 ( .A(n19303), .B(n2173), .Z(n521) );
  NANDN U788 ( .A(n19282), .B(n2174), .Z(n522) );
  AND U789 ( .A(n521), .B(n522), .Z(n19309) );
  NANDN U790 ( .A(n19450), .B(n2173), .Z(n523) );
  NANDN U791 ( .A(n19429), .B(n2174), .Z(n524) );
  AND U792 ( .A(n523), .B(n524), .Z(n19456) );
  NANDN U793 ( .A(n19597), .B(n2173), .Z(n525) );
  NANDN U794 ( .A(n19576), .B(n2174), .Z(n526) );
  AND U795 ( .A(n525), .B(n526), .Z(n19603) );
  NANDN U796 ( .A(n19740), .B(n2173), .Z(n527) );
  NANDN U797 ( .A(n19719), .B(n2174), .Z(n528) );
  AND U798 ( .A(n527), .B(n528), .Z(n19746) );
  NANDN U799 ( .A(n19887), .B(n2173), .Z(n529) );
  NANDN U800 ( .A(n19866), .B(n2174), .Z(n530) );
  AND U801 ( .A(n529), .B(n530), .Z(n19893) );
  NANDN U802 ( .A(n20034), .B(n2173), .Z(n531) );
  NANDN U803 ( .A(n20013), .B(n2174), .Z(n532) );
  AND U804 ( .A(n531), .B(n532), .Z(n20040) );
  NANDN U805 ( .A(n20177), .B(n2173), .Z(n533) );
  NANDN U806 ( .A(n20156), .B(n2174), .Z(n534) );
  AND U807 ( .A(n533), .B(n534), .Z(n20183) );
  NANDN U808 ( .A(n20324), .B(n2173), .Z(n535) );
  NANDN U809 ( .A(n20303), .B(n2174), .Z(n536) );
  AND U810 ( .A(n535), .B(n536), .Z(n20330) );
  NANDN U811 ( .A(n20471), .B(n2173), .Z(n537) );
  NANDN U812 ( .A(n20450), .B(n2174), .Z(n538) );
  AND U813 ( .A(n537), .B(n538), .Z(n20477) );
  NANDN U814 ( .A(n20618), .B(n2173), .Z(n539) );
  NANDN U815 ( .A(n20597), .B(n2174), .Z(n540) );
  AND U816 ( .A(n539), .B(n540), .Z(n20624) );
  NANDN U817 ( .A(n20765), .B(n2173), .Z(n541) );
  NANDN U818 ( .A(n20744), .B(n2174), .Z(n542) );
  AND U819 ( .A(n541), .B(n542), .Z(n20771) );
  NANDN U820 ( .A(n20912), .B(n2173), .Z(n543) );
  NANDN U821 ( .A(n20891), .B(n2174), .Z(n544) );
  AND U822 ( .A(n543), .B(n544), .Z(n20918) );
  NANDN U823 ( .A(n21055), .B(n2173), .Z(n545) );
  NANDN U824 ( .A(n21036), .B(n2174), .Z(n546) );
  AND U825 ( .A(n545), .B(n546), .Z(n21061) );
  NANDN U826 ( .A(n21202), .B(n2173), .Z(n547) );
  NANDN U827 ( .A(n21181), .B(n2174), .Z(n548) );
  AND U828 ( .A(n547), .B(n548), .Z(n21208) );
  NANDN U829 ( .A(n21345), .B(n2173), .Z(n549) );
  NANDN U830 ( .A(n21324), .B(n2174), .Z(n550) );
  AND U831 ( .A(n549), .B(n550), .Z(n21351) );
  NANDN U832 ( .A(n21492), .B(n2173), .Z(n551) );
  NANDN U833 ( .A(n21471), .B(n2174), .Z(n552) );
  AND U834 ( .A(n551), .B(n552), .Z(n21498) );
  NANDN U835 ( .A(n21639), .B(n2173), .Z(n553) );
  NANDN U836 ( .A(n21618), .B(n2174), .Z(n554) );
  AND U837 ( .A(n553), .B(n554), .Z(n21645) );
  NANDN U838 ( .A(n21786), .B(n2173), .Z(n555) );
  NANDN U839 ( .A(n21765), .B(n2174), .Z(n556) );
  AND U840 ( .A(n555), .B(n556), .Z(n21792) );
  NANDN U841 ( .A(n21933), .B(n2173), .Z(n557) );
  NANDN U842 ( .A(n21912), .B(n2174), .Z(n558) );
  AND U843 ( .A(n557), .B(n558), .Z(n21939) );
  NANDN U844 ( .A(n22080), .B(n2173), .Z(n559) );
  NANDN U845 ( .A(n22059), .B(n2174), .Z(n560) );
  AND U846 ( .A(n559), .B(n560), .Z(n22086) );
  NANDN U847 ( .A(n22227), .B(n2173), .Z(n561) );
  NANDN U848 ( .A(n22206), .B(n2174), .Z(n562) );
  AND U849 ( .A(n561), .B(n562), .Z(n22233) );
  NANDN U850 ( .A(n22370), .B(n2173), .Z(n563) );
  NANDN U851 ( .A(n22349), .B(n2174), .Z(n564) );
  AND U852 ( .A(n563), .B(n564), .Z(n22376) );
  NANDN U853 ( .A(n22517), .B(n2173), .Z(n565) );
  NANDN U854 ( .A(n22496), .B(n2174), .Z(n566) );
  AND U855 ( .A(n565), .B(n566), .Z(n22523) );
  NANDN U856 ( .A(n22664), .B(n2173), .Z(n567) );
  NANDN U857 ( .A(n22643), .B(n2174), .Z(n568) );
  AND U858 ( .A(n567), .B(n568), .Z(n22670) );
  NANDN U859 ( .A(n22811), .B(n2173), .Z(n569) );
  NANDN U860 ( .A(n22790), .B(n2174), .Z(n570) );
  AND U861 ( .A(n569), .B(n570), .Z(n22817) );
  NANDN U862 ( .A(n22958), .B(n2173), .Z(n571) );
  NANDN U863 ( .A(n22937), .B(n2174), .Z(n572) );
  AND U864 ( .A(n571), .B(n572), .Z(n22964) );
  NANDN U865 ( .A(n23105), .B(n2173), .Z(n573) );
  NANDN U866 ( .A(n23084), .B(n2174), .Z(n574) );
  AND U867 ( .A(n573), .B(n574), .Z(n23111) );
  NANDN U868 ( .A(n23252), .B(n2173), .Z(n575) );
  NANDN U869 ( .A(n23231), .B(n2174), .Z(n576) );
  AND U870 ( .A(n575), .B(n576), .Z(n23258) );
  NANDN U871 ( .A(n23399), .B(n2173), .Z(n577) );
  NANDN U872 ( .A(n23378), .B(n2174), .Z(n578) );
  AND U873 ( .A(n577), .B(n578), .Z(n23405) );
  NANDN U874 ( .A(n23546), .B(n2173), .Z(n579) );
  NANDN U875 ( .A(n23525), .B(n2174), .Z(n580) );
  AND U876 ( .A(n579), .B(n580), .Z(n23552) );
  NANDN U877 ( .A(n2499), .B(n2173), .Z(n581) );
  NANDN U878 ( .A(n2478), .B(n2174), .Z(n582) );
  AND U879 ( .A(n581), .B(n582), .Z(n2505) );
  NANDN U880 ( .A(n2646), .B(n2173), .Z(n583) );
  NANDN U881 ( .A(n2625), .B(n2174), .Z(n584) );
  AND U882 ( .A(n583), .B(n584), .Z(n2652) );
  NANDN U883 ( .A(n2793), .B(n2173), .Z(n585) );
  NANDN U884 ( .A(n2772), .B(n2174), .Z(n586) );
  AND U885 ( .A(n585), .B(n586), .Z(n2799) );
  NANDN U886 ( .A(n2940), .B(n2173), .Z(n587) );
  NANDN U887 ( .A(n2919), .B(n2174), .Z(n588) );
  AND U888 ( .A(n587), .B(n588), .Z(n2946) );
  NANDN U889 ( .A(n3087), .B(n2173), .Z(n589) );
  NANDN U890 ( .A(n3066), .B(n2174), .Z(n590) );
  AND U891 ( .A(n589), .B(n590), .Z(n3093) );
  NANDN U892 ( .A(n3234), .B(n2173), .Z(n591) );
  NANDN U893 ( .A(n3213), .B(n2174), .Z(n592) );
  AND U894 ( .A(n591), .B(n592), .Z(n3240) );
  NANDN U895 ( .A(n3381), .B(n2173), .Z(n593) );
  NANDN U896 ( .A(n3360), .B(n2174), .Z(n594) );
  AND U897 ( .A(n593), .B(n594), .Z(n3387) );
  NANDN U898 ( .A(n3528), .B(n2173), .Z(n595) );
  NANDN U899 ( .A(n3507), .B(n2174), .Z(n596) );
  AND U900 ( .A(n595), .B(n596), .Z(n3534) );
  NANDN U901 ( .A(n3675), .B(n2173), .Z(n597) );
  NANDN U902 ( .A(n3654), .B(n2174), .Z(n598) );
  AND U903 ( .A(n597), .B(n598), .Z(n3681) );
  NANDN U904 ( .A(n3822), .B(n2173), .Z(n599) );
  NANDN U905 ( .A(n3801), .B(n2174), .Z(n600) );
  AND U906 ( .A(n599), .B(n600), .Z(n3828) );
  NANDN U907 ( .A(n3969), .B(n2173), .Z(n601) );
  NANDN U908 ( .A(n3948), .B(n2174), .Z(n602) );
  AND U909 ( .A(n601), .B(n602), .Z(n3975) );
  NANDN U910 ( .A(n4116), .B(n2173), .Z(n603) );
  NANDN U911 ( .A(n4095), .B(n2174), .Z(n604) );
  AND U912 ( .A(n603), .B(n604), .Z(n4122) );
  NANDN U913 ( .A(n4263), .B(n2173), .Z(n605) );
  NANDN U914 ( .A(n4242), .B(n2174), .Z(n606) );
  AND U915 ( .A(n605), .B(n606), .Z(n4269) );
  NANDN U916 ( .A(n4408), .B(n2173), .Z(n607) );
  NANDN U917 ( .A(n4389), .B(n2174), .Z(n608) );
  AND U918 ( .A(n607), .B(n608), .Z(n4415) );
  NANDN U919 ( .A(n4553), .B(n2173), .Z(n609) );
  NANDN U920 ( .A(n4532), .B(n2174), .Z(n610) );
  AND U921 ( .A(n609), .B(n610), .Z(n4559) );
  NANDN U922 ( .A(n4700), .B(n2173), .Z(n611) );
  NANDN U923 ( .A(n4679), .B(n2174), .Z(n612) );
  AND U924 ( .A(n611), .B(n612), .Z(n4706) );
  NANDN U925 ( .A(n4847), .B(n2173), .Z(n613) );
  NANDN U926 ( .A(n4826), .B(n2174), .Z(n614) );
  AND U927 ( .A(n613), .B(n614), .Z(n4853) );
  NANDN U928 ( .A(n4994), .B(n2173), .Z(n615) );
  NANDN U929 ( .A(n4973), .B(n2174), .Z(n616) );
  AND U930 ( .A(n615), .B(n616), .Z(n5000) );
  NANDN U931 ( .A(n5141), .B(n2173), .Z(n617) );
  NANDN U932 ( .A(n5120), .B(n2174), .Z(n618) );
  AND U933 ( .A(n617), .B(n618), .Z(n5147) );
  NANDN U934 ( .A(n5288), .B(n2173), .Z(n619) );
  NANDN U935 ( .A(n5267), .B(n2174), .Z(n620) );
  AND U936 ( .A(n619), .B(n620), .Z(n5294) );
  NANDN U937 ( .A(n5435), .B(n2173), .Z(n621) );
  NANDN U938 ( .A(n5414), .B(n2174), .Z(n622) );
  AND U939 ( .A(n621), .B(n622), .Z(n5441) );
  NANDN U940 ( .A(n5582), .B(n2173), .Z(n623) );
  NANDN U941 ( .A(n5561), .B(n2174), .Z(n624) );
  AND U942 ( .A(n623), .B(n624), .Z(n5588) );
  NANDN U943 ( .A(n5729), .B(n2173), .Z(n625) );
  NANDN U944 ( .A(n5708), .B(n2174), .Z(n626) );
  AND U945 ( .A(n625), .B(n626), .Z(n5735) );
  NANDN U946 ( .A(n5876), .B(n2173), .Z(n627) );
  NANDN U947 ( .A(n5855), .B(n2174), .Z(n628) );
  AND U948 ( .A(n627), .B(n628), .Z(n5882) );
  NANDN U949 ( .A(n6023), .B(n2173), .Z(n629) );
  NANDN U950 ( .A(n6002), .B(n2174), .Z(n630) );
  AND U951 ( .A(n629), .B(n630), .Z(n6029) );
  NANDN U952 ( .A(n6170), .B(n2173), .Z(n631) );
  NANDN U953 ( .A(n6149), .B(n2174), .Z(n632) );
  AND U954 ( .A(n631), .B(n632), .Z(n6176) );
  NANDN U955 ( .A(n6317), .B(n2173), .Z(n633) );
  NANDN U956 ( .A(n6296), .B(n2174), .Z(n634) );
  AND U957 ( .A(n633), .B(n634), .Z(n6323) );
  NANDN U958 ( .A(n6460), .B(n2173), .Z(n635) );
  NANDN U959 ( .A(n6439), .B(n2174), .Z(n636) );
  AND U960 ( .A(n635), .B(n636), .Z(n6466) );
  NANDN U961 ( .A(n6607), .B(n2173), .Z(n637) );
  NANDN U962 ( .A(n6586), .B(n2174), .Z(n638) );
  AND U963 ( .A(n637), .B(n638), .Z(n6613) );
  NANDN U964 ( .A(n6754), .B(n2173), .Z(n639) );
  NANDN U965 ( .A(n6733), .B(n2174), .Z(n640) );
  AND U966 ( .A(n639), .B(n640), .Z(n6760) );
  NANDN U967 ( .A(n6897), .B(n2173), .Z(n641) );
  NANDN U968 ( .A(n6876), .B(n2174), .Z(n642) );
  AND U969 ( .A(n641), .B(n642), .Z(n6903) );
  NANDN U970 ( .A(n7040), .B(n2173), .Z(n643) );
  NANDN U971 ( .A(n7019), .B(n2174), .Z(n644) );
  AND U972 ( .A(n643), .B(n644), .Z(n7046) );
  NANDN U973 ( .A(n7183), .B(n2173), .Z(n645) );
  NANDN U974 ( .A(n7162), .B(n2174), .Z(n646) );
  AND U975 ( .A(n645), .B(n646), .Z(n7189) );
  NANDN U976 ( .A(n7330), .B(n2173), .Z(n647) );
  NANDN U977 ( .A(n7309), .B(n2174), .Z(n648) );
  AND U978 ( .A(n647), .B(n648), .Z(n7336) );
  NANDN U979 ( .A(n7477), .B(n2173), .Z(n649) );
  NANDN U980 ( .A(n7456), .B(n2174), .Z(n650) );
  AND U981 ( .A(n649), .B(n650), .Z(n7483) );
  NANDN U982 ( .A(n7620), .B(n2173), .Z(n651) );
  NANDN U983 ( .A(n7599), .B(n2174), .Z(n652) );
  AND U984 ( .A(n651), .B(n652), .Z(n7626) );
  NANDN U985 ( .A(n7767), .B(n2173), .Z(n653) );
  NANDN U986 ( .A(n7746), .B(n2174), .Z(n654) );
  AND U987 ( .A(n653), .B(n654), .Z(n7773) );
  NANDN U988 ( .A(n7910), .B(n2173), .Z(n655) );
  NANDN U989 ( .A(n7889), .B(n2174), .Z(n656) );
  AND U990 ( .A(n655), .B(n656), .Z(n7916) );
  NANDN U991 ( .A(n8053), .B(n2173), .Z(n657) );
  NANDN U992 ( .A(n8032), .B(n2174), .Z(n658) );
  AND U993 ( .A(n657), .B(n658), .Z(n8059) );
  NANDN U994 ( .A(n8198), .B(n2173), .Z(n659) );
  NANDN U995 ( .A(n8179), .B(n2174), .Z(n660) );
  AND U996 ( .A(n659), .B(n660), .Z(n8205) );
  NANDN U997 ( .A(n8343), .B(n2173), .Z(n661) );
  NANDN U998 ( .A(n8322), .B(n2174), .Z(n662) );
  AND U999 ( .A(n661), .B(n662), .Z(n8349) );
  NANDN U1000 ( .A(n8490), .B(n2173), .Z(n663) );
  NANDN U1001 ( .A(n8469), .B(n2174), .Z(n664) );
  AND U1002 ( .A(n663), .B(n664), .Z(n8496) );
  NANDN U1003 ( .A(n8637), .B(n2173), .Z(n665) );
  NANDN U1004 ( .A(n8616), .B(n2174), .Z(n666) );
  AND U1005 ( .A(n665), .B(n666), .Z(n8643) );
  NANDN U1006 ( .A(n8784), .B(n2173), .Z(n667) );
  NANDN U1007 ( .A(n8763), .B(n2174), .Z(n668) );
  AND U1008 ( .A(n667), .B(n668), .Z(n8790) );
  NANDN U1009 ( .A(n8931), .B(n2173), .Z(n669) );
  NANDN U1010 ( .A(n8910), .B(n2174), .Z(n670) );
  AND U1011 ( .A(n669), .B(n670), .Z(n8937) );
  NANDN U1012 ( .A(n9074), .B(n2173), .Z(n671) );
  NANDN U1013 ( .A(n9055), .B(n2174), .Z(n672) );
  AND U1014 ( .A(n671), .B(n672), .Z(n9080) );
  NANDN U1015 ( .A(n9217), .B(n2173), .Z(n673) );
  NANDN U1016 ( .A(n9198), .B(n2174), .Z(n674) );
  AND U1017 ( .A(n673), .B(n674), .Z(n9223) );
  NANDN U1018 ( .A(n9364), .B(n2173), .Z(n675) );
  NANDN U1019 ( .A(n9343), .B(n2174), .Z(n676) );
  AND U1020 ( .A(n675), .B(n676), .Z(n9370) );
  NANDN U1021 ( .A(n9511), .B(n2173), .Z(n677) );
  NANDN U1022 ( .A(n9490), .B(n2174), .Z(n678) );
  AND U1023 ( .A(n677), .B(n678), .Z(n9517) );
  NANDN U1024 ( .A(n9658), .B(n2173), .Z(n679) );
  NANDN U1025 ( .A(n9637), .B(n2174), .Z(n680) );
  AND U1026 ( .A(n679), .B(n680), .Z(n9664) );
  NANDN U1027 ( .A(n9805), .B(n2173), .Z(n681) );
  NANDN U1028 ( .A(n9784), .B(n2174), .Z(n682) );
  AND U1029 ( .A(n681), .B(n682), .Z(n9811) );
  NANDN U1030 ( .A(n9952), .B(n2173), .Z(n683) );
  NANDN U1031 ( .A(n9931), .B(n2174), .Z(n684) );
  AND U1032 ( .A(n683), .B(n684), .Z(n9958) );
  NANDN U1033 ( .A(n10099), .B(n2173), .Z(n685) );
  NANDN U1034 ( .A(n10078), .B(n2174), .Z(n686) );
  AND U1035 ( .A(n685), .B(n686), .Z(n10105) );
  NANDN U1036 ( .A(n10246), .B(n2173), .Z(n687) );
  NANDN U1037 ( .A(n10225), .B(n2174), .Z(n688) );
  AND U1038 ( .A(n687), .B(n688), .Z(n10252) );
  NANDN U1039 ( .A(n10393), .B(n2173), .Z(n689) );
  NANDN U1040 ( .A(n10372), .B(n2174), .Z(n690) );
  AND U1041 ( .A(n689), .B(n690), .Z(n10399) );
  NANDN U1042 ( .A(n10540), .B(n2173), .Z(n691) );
  NANDN U1043 ( .A(n10519), .B(n2174), .Z(n692) );
  AND U1044 ( .A(n691), .B(n692), .Z(n10546) );
  NANDN U1045 ( .A(n10687), .B(n2173), .Z(n693) );
  NANDN U1046 ( .A(n10666), .B(n2174), .Z(n694) );
  AND U1047 ( .A(n693), .B(n694), .Z(n10693) );
  NANDN U1048 ( .A(n10834), .B(n2173), .Z(n695) );
  NANDN U1049 ( .A(n10813), .B(n2174), .Z(n696) );
  AND U1050 ( .A(n695), .B(n696), .Z(n10840) );
  NANDN U1051 ( .A(n10981), .B(n2173), .Z(n697) );
  NANDN U1052 ( .A(n10960), .B(n2174), .Z(n698) );
  AND U1053 ( .A(n697), .B(n698), .Z(n10987) );
  NANDN U1054 ( .A(n11128), .B(n2173), .Z(n699) );
  NANDN U1055 ( .A(n11107), .B(n2174), .Z(n700) );
  AND U1056 ( .A(n699), .B(n700), .Z(n11134) );
  NANDN U1057 ( .A(n11275), .B(n2173), .Z(n701) );
  NANDN U1058 ( .A(n11254), .B(n2174), .Z(n702) );
  AND U1059 ( .A(n701), .B(n702), .Z(n11281) );
  NANDN U1060 ( .A(n11422), .B(n2173), .Z(n703) );
  NANDN U1061 ( .A(n11401), .B(n2174), .Z(n704) );
  AND U1062 ( .A(n703), .B(n704), .Z(n11428) );
  NANDN U1063 ( .A(n11569), .B(n2173), .Z(n705) );
  NANDN U1064 ( .A(n11548), .B(n2174), .Z(n706) );
  AND U1065 ( .A(n705), .B(n706), .Z(n11575) );
  NANDN U1066 ( .A(n11716), .B(n2173), .Z(n707) );
  NANDN U1067 ( .A(n11695), .B(n2174), .Z(n708) );
  AND U1068 ( .A(n707), .B(n708), .Z(n11722) );
  NANDN U1069 ( .A(n11855), .B(n2173), .Z(n709) );
  NANDN U1070 ( .A(n11834), .B(n2174), .Z(n710) );
  AND U1071 ( .A(n709), .B(n710), .Z(n11861) );
  NANDN U1072 ( .A(n12002), .B(n2173), .Z(n711) );
  NANDN U1073 ( .A(n11981), .B(n2174), .Z(n712) );
  AND U1074 ( .A(n711), .B(n712), .Z(n12008) );
  NANDN U1075 ( .A(n12149), .B(n2173), .Z(n713) );
  NANDN U1076 ( .A(n12128), .B(n2174), .Z(n714) );
  AND U1077 ( .A(n713), .B(n714), .Z(n12155) );
  NANDN U1078 ( .A(n12296), .B(n2173), .Z(n715) );
  NANDN U1079 ( .A(n12275), .B(n2174), .Z(n716) );
  AND U1080 ( .A(n715), .B(n716), .Z(n12302) );
  NANDN U1081 ( .A(n12443), .B(n2173), .Z(n717) );
  NANDN U1082 ( .A(n12422), .B(n2174), .Z(n718) );
  AND U1083 ( .A(n717), .B(n718), .Z(n12449) );
  NANDN U1084 ( .A(n12590), .B(n2173), .Z(n719) );
  NANDN U1085 ( .A(n12569), .B(n2174), .Z(n720) );
  AND U1086 ( .A(n719), .B(n720), .Z(n12596) );
  NANDN U1087 ( .A(n12733), .B(n2173), .Z(n721) );
  NANDN U1088 ( .A(n12712), .B(n2174), .Z(n722) );
  AND U1089 ( .A(n721), .B(n722), .Z(n12739) );
  NANDN U1090 ( .A(n12880), .B(n2173), .Z(n723) );
  NANDN U1091 ( .A(n12859), .B(n2174), .Z(n724) );
  AND U1092 ( .A(n723), .B(n724), .Z(n12886) );
  NANDN U1093 ( .A(n13027), .B(n2173), .Z(n725) );
  NANDN U1094 ( .A(n13006), .B(n2174), .Z(n726) );
  AND U1095 ( .A(n725), .B(n726), .Z(n13033) );
  NANDN U1096 ( .A(n13174), .B(n2173), .Z(n727) );
  NANDN U1097 ( .A(n13153), .B(n2174), .Z(n728) );
  AND U1098 ( .A(n727), .B(n728), .Z(n13180) );
  NANDN U1099 ( .A(n13321), .B(n2173), .Z(n729) );
  NANDN U1100 ( .A(n13300), .B(n2174), .Z(n730) );
  AND U1101 ( .A(n729), .B(n730), .Z(n13327) );
  NANDN U1102 ( .A(n13468), .B(n2173), .Z(n731) );
  NANDN U1103 ( .A(n13447), .B(n2174), .Z(n732) );
  AND U1104 ( .A(n731), .B(n732), .Z(n13474) );
  NANDN U1105 ( .A(n13615), .B(n2173), .Z(n733) );
  NANDN U1106 ( .A(n13594), .B(n2174), .Z(n734) );
  AND U1107 ( .A(n733), .B(n734), .Z(n13621) );
  NANDN U1108 ( .A(n13762), .B(n2173), .Z(n735) );
  NANDN U1109 ( .A(n13741), .B(n2174), .Z(n736) );
  AND U1110 ( .A(n735), .B(n736), .Z(n13768) );
  NANDN U1111 ( .A(n13905), .B(n2173), .Z(n737) );
  NANDN U1112 ( .A(n13884), .B(n2174), .Z(n738) );
  AND U1113 ( .A(n737), .B(n738), .Z(n13911) );
  NANDN U1114 ( .A(n14052), .B(n2173), .Z(n739) );
  NANDN U1115 ( .A(n14031), .B(n2174), .Z(n740) );
  AND U1116 ( .A(n739), .B(n740), .Z(n14058) );
  NANDN U1117 ( .A(n14199), .B(n2173), .Z(n741) );
  NANDN U1118 ( .A(n14178), .B(n2174), .Z(n742) );
  AND U1119 ( .A(n741), .B(n742), .Z(n14205) );
  NANDN U1120 ( .A(n14346), .B(n2173), .Z(n743) );
  NANDN U1121 ( .A(n14325), .B(n2174), .Z(n744) );
  AND U1122 ( .A(n743), .B(n744), .Z(n14352) );
  NANDN U1123 ( .A(n14493), .B(n2173), .Z(n745) );
  NANDN U1124 ( .A(n14472), .B(n2174), .Z(n746) );
  AND U1125 ( .A(n745), .B(n746), .Z(n14499) );
  NANDN U1126 ( .A(n14640), .B(n2173), .Z(n747) );
  NANDN U1127 ( .A(n14619), .B(n2174), .Z(n748) );
  AND U1128 ( .A(n747), .B(n748), .Z(n14646) );
  NANDN U1129 ( .A(n14783), .B(n2173), .Z(n749) );
  NANDN U1130 ( .A(n14764), .B(n2174), .Z(n750) );
  AND U1131 ( .A(n749), .B(n750), .Z(n14789) );
  NANDN U1132 ( .A(n14930), .B(n2173), .Z(n751) );
  NANDN U1133 ( .A(n14909), .B(n2174), .Z(n752) );
  AND U1134 ( .A(n751), .B(n752), .Z(n14936) );
  NANDN U1135 ( .A(n15077), .B(n2173), .Z(n753) );
  NANDN U1136 ( .A(n15056), .B(n2174), .Z(n754) );
  AND U1137 ( .A(n753), .B(n754), .Z(n15083) );
  NANDN U1138 ( .A(n15224), .B(n2173), .Z(n755) );
  NANDN U1139 ( .A(n15203), .B(n2174), .Z(n756) );
  AND U1140 ( .A(n755), .B(n756), .Z(n15230) );
  NANDN U1141 ( .A(n15371), .B(n2173), .Z(n757) );
  NANDN U1142 ( .A(n15350), .B(n2174), .Z(n758) );
  AND U1143 ( .A(n757), .B(n758), .Z(n15377) );
  NANDN U1144 ( .A(n15518), .B(n2173), .Z(n759) );
  NANDN U1145 ( .A(n15497), .B(n2174), .Z(n760) );
  AND U1146 ( .A(n759), .B(n760), .Z(n15524) );
  NANDN U1147 ( .A(n15661), .B(n2173), .Z(n761) );
  NANDN U1148 ( .A(n15640), .B(n2174), .Z(n762) );
  AND U1149 ( .A(n761), .B(n762), .Z(n15667) );
  NANDN U1150 ( .A(n15808), .B(n2173), .Z(n763) );
  NANDN U1151 ( .A(n15787), .B(n2174), .Z(n764) );
  AND U1152 ( .A(n763), .B(n764), .Z(n15814) );
  NANDN U1153 ( .A(n15955), .B(n2173), .Z(n765) );
  NANDN U1154 ( .A(n15934), .B(n2174), .Z(n766) );
  AND U1155 ( .A(n765), .B(n766), .Z(n15961) );
  NANDN U1156 ( .A(n16102), .B(n2173), .Z(n767) );
  NANDN U1157 ( .A(n16081), .B(n2174), .Z(n768) );
  AND U1158 ( .A(n767), .B(n768), .Z(n16108) );
  NANDN U1159 ( .A(n16249), .B(n2173), .Z(n769) );
  NANDN U1160 ( .A(n16228), .B(n2174), .Z(n770) );
  AND U1161 ( .A(n769), .B(n770), .Z(n16255) );
  NANDN U1162 ( .A(n16396), .B(n2173), .Z(n771) );
  NANDN U1163 ( .A(n16375), .B(n2174), .Z(n772) );
  AND U1164 ( .A(n771), .B(n772), .Z(n16402) );
  NANDN U1165 ( .A(n16543), .B(n2173), .Z(n773) );
  NANDN U1166 ( .A(n16522), .B(n2174), .Z(n774) );
  AND U1167 ( .A(n773), .B(n774), .Z(n16549) );
  NANDN U1168 ( .A(n16690), .B(n2173), .Z(n775) );
  NANDN U1169 ( .A(n16669), .B(n2174), .Z(n776) );
  AND U1170 ( .A(n775), .B(n776), .Z(n16696) );
  NANDN U1171 ( .A(n16837), .B(n2173), .Z(n777) );
  NANDN U1172 ( .A(n16816), .B(n2174), .Z(n778) );
  AND U1173 ( .A(n777), .B(n778), .Z(n16843) );
  NANDN U1174 ( .A(n16984), .B(n2173), .Z(n779) );
  NANDN U1175 ( .A(n16963), .B(n2174), .Z(n780) );
  AND U1176 ( .A(n779), .B(n780), .Z(n16990) );
  NANDN U1177 ( .A(n17131), .B(n2173), .Z(n781) );
  NANDN U1178 ( .A(n17110), .B(n2174), .Z(n782) );
  AND U1179 ( .A(n781), .B(n782), .Z(n17137) );
  NANDN U1180 ( .A(n17278), .B(n2173), .Z(n783) );
  NANDN U1181 ( .A(n17257), .B(n2174), .Z(n784) );
  AND U1182 ( .A(n783), .B(n784), .Z(n17284) );
  NANDN U1183 ( .A(n17425), .B(n2173), .Z(n785) );
  NANDN U1184 ( .A(n17404), .B(n2174), .Z(n786) );
  AND U1185 ( .A(n785), .B(n786), .Z(n17431) );
  NANDN U1186 ( .A(n17572), .B(n2173), .Z(n787) );
  NANDN U1187 ( .A(n17551), .B(n2174), .Z(n788) );
  AND U1188 ( .A(n787), .B(n788), .Z(n17578) );
  NANDN U1189 ( .A(n17719), .B(n2173), .Z(n789) );
  NANDN U1190 ( .A(n17698), .B(n2174), .Z(n790) );
  AND U1191 ( .A(n789), .B(n790), .Z(n17725) );
  NANDN U1192 ( .A(n17858), .B(n2173), .Z(n791) );
  NANDN U1193 ( .A(n17837), .B(n2174), .Z(n792) );
  AND U1194 ( .A(n791), .B(n792), .Z(n17864) );
  NANDN U1195 ( .A(n18005), .B(n2173), .Z(n793) );
  NANDN U1196 ( .A(n17984), .B(n2174), .Z(n794) );
  AND U1197 ( .A(n793), .B(n794), .Z(n18011) );
  NANDN U1198 ( .A(n18148), .B(n2173), .Z(n795) );
  NANDN U1199 ( .A(n18127), .B(n2174), .Z(n796) );
  AND U1200 ( .A(n795), .B(n796), .Z(n18154) );
  NANDN U1201 ( .A(n18295), .B(n2173), .Z(n797) );
  NANDN U1202 ( .A(n18274), .B(n2174), .Z(n798) );
  AND U1203 ( .A(n797), .B(n798), .Z(n18301) );
  NANDN U1204 ( .A(n18442), .B(n2173), .Z(n799) );
  NANDN U1205 ( .A(n18421), .B(n2174), .Z(n800) );
  AND U1206 ( .A(n799), .B(n800), .Z(n18448) );
  NANDN U1207 ( .A(n18589), .B(n2173), .Z(n801) );
  NANDN U1208 ( .A(n18568), .B(n2174), .Z(n802) );
  AND U1209 ( .A(n801), .B(n802), .Z(n18595) );
  NANDN U1210 ( .A(n18736), .B(n2173), .Z(n803) );
  NANDN U1211 ( .A(n18715), .B(n2174), .Z(n804) );
  AND U1212 ( .A(n803), .B(n804), .Z(n18742) );
  NANDN U1213 ( .A(n18883), .B(n2173), .Z(n805) );
  NANDN U1214 ( .A(n18862), .B(n2174), .Z(n806) );
  AND U1215 ( .A(n805), .B(n806), .Z(n18889) );
  NANDN U1216 ( .A(n19030), .B(n2173), .Z(n807) );
  NANDN U1217 ( .A(n19009), .B(n2174), .Z(n808) );
  AND U1218 ( .A(n807), .B(n808), .Z(n19036) );
  NANDN U1219 ( .A(n19177), .B(n2173), .Z(n809) );
  NANDN U1220 ( .A(n19156), .B(n2174), .Z(n810) );
  AND U1221 ( .A(n809), .B(n810), .Z(n19183) );
  NANDN U1222 ( .A(n19324), .B(n2173), .Z(n811) );
  NANDN U1223 ( .A(n19303), .B(n2174), .Z(n812) );
  AND U1224 ( .A(n811), .B(n812), .Z(n19330) );
  NANDN U1225 ( .A(n19471), .B(n2173), .Z(n813) );
  NANDN U1226 ( .A(n19450), .B(n2174), .Z(n814) );
  AND U1227 ( .A(n813), .B(n814), .Z(n19477) );
  NANDN U1228 ( .A(n19618), .B(n2173), .Z(n815) );
  NANDN U1229 ( .A(n19597), .B(n2174), .Z(n816) );
  AND U1230 ( .A(n815), .B(n816), .Z(n19624) );
  NANDN U1231 ( .A(n19761), .B(n2173), .Z(n817) );
  NANDN U1232 ( .A(n19740), .B(n2174), .Z(n818) );
  AND U1233 ( .A(n817), .B(n818), .Z(n19767) );
  NANDN U1234 ( .A(n19908), .B(n2173), .Z(n819) );
  NANDN U1235 ( .A(n19887), .B(n2174), .Z(n820) );
  AND U1236 ( .A(n819), .B(n820), .Z(n19914) );
  NANDN U1237 ( .A(n20055), .B(n2173), .Z(n821) );
  NANDN U1238 ( .A(n20034), .B(n2174), .Z(n822) );
  AND U1239 ( .A(n821), .B(n822), .Z(n20061) );
  NANDN U1240 ( .A(n20198), .B(n2173), .Z(n823) );
  NANDN U1241 ( .A(n20177), .B(n2174), .Z(n824) );
  AND U1242 ( .A(n823), .B(n824), .Z(n20204) );
  NANDN U1243 ( .A(n20345), .B(n2173), .Z(n825) );
  NANDN U1244 ( .A(n20324), .B(n2174), .Z(n826) );
  AND U1245 ( .A(n825), .B(n826), .Z(n20351) );
  NANDN U1246 ( .A(n20492), .B(n2173), .Z(n827) );
  NANDN U1247 ( .A(n20471), .B(n2174), .Z(n828) );
  AND U1248 ( .A(n827), .B(n828), .Z(n20498) );
  NANDN U1249 ( .A(n20639), .B(n2173), .Z(n829) );
  NANDN U1250 ( .A(n20618), .B(n2174), .Z(n830) );
  AND U1251 ( .A(n829), .B(n830), .Z(n20645) );
  NANDN U1252 ( .A(n20786), .B(n2173), .Z(n831) );
  NANDN U1253 ( .A(n20765), .B(n2174), .Z(n832) );
  AND U1254 ( .A(n831), .B(n832), .Z(n20792) );
  NANDN U1255 ( .A(n20933), .B(n2173), .Z(n833) );
  NANDN U1256 ( .A(n20912), .B(n2174), .Z(n834) );
  AND U1257 ( .A(n833), .B(n834), .Z(n20939) );
  NANDN U1258 ( .A(n21076), .B(n2173), .Z(n835) );
  NANDN U1259 ( .A(n21055), .B(n2174), .Z(n836) );
  AND U1260 ( .A(n835), .B(n836), .Z(n21082) );
  NANDN U1261 ( .A(n21223), .B(n2173), .Z(n837) );
  NANDN U1262 ( .A(n21202), .B(n2174), .Z(n838) );
  AND U1263 ( .A(n837), .B(n838), .Z(n21229) );
  NANDN U1264 ( .A(n21366), .B(n2173), .Z(n839) );
  NANDN U1265 ( .A(n21345), .B(n2174), .Z(n840) );
  AND U1266 ( .A(n839), .B(n840), .Z(n21372) );
  NANDN U1267 ( .A(n21513), .B(n2173), .Z(n841) );
  NANDN U1268 ( .A(n21492), .B(n2174), .Z(n842) );
  AND U1269 ( .A(n841), .B(n842), .Z(n21519) );
  NANDN U1270 ( .A(n21660), .B(n2173), .Z(n843) );
  NANDN U1271 ( .A(n21639), .B(n2174), .Z(n844) );
  AND U1272 ( .A(n843), .B(n844), .Z(n21666) );
  NANDN U1273 ( .A(n21807), .B(n2173), .Z(n845) );
  NANDN U1274 ( .A(n21786), .B(n2174), .Z(n846) );
  AND U1275 ( .A(n845), .B(n846), .Z(n21813) );
  NANDN U1276 ( .A(n21954), .B(n2173), .Z(n847) );
  NANDN U1277 ( .A(n21933), .B(n2174), .Z(n848) );
  AND U1278 ( .A(n847), .B(n848), .Z(n21960) );
  NANDN U1279 ( .A(n22101), .B(n2173), .Z(n849) );
  NANDN U1280 ( .A(n22080), .B(n2174), .Z(n850) );
  AND U1281 ( .A(n849), .B(n850), .Z(n22107) );
  NANDN U1282 ( .A(n22248), .B(n2173), .Z(n851) );
  NANDN U1283 ( .A(n22227), .B(n2174), .Z(n852) );
  AND U1284 ( .A(n851), .B(n852), .Z(n22254) );
  NANDN U1285 ( .A(n22391), .B(n2173), .Z(n853) );
  NANDN U1286 ( .A(n22370), .B(n2174), .Z(n854) );
  AND U1287 ( .A(n853), .B(n854), .Z(n22397) );
  NANDN U1288 ( .A(n22538), .B(n2173), .Z(n855) );
  NANDN U1289 ( .A(n22517), .B(n2174), .Z(n856) );
  AND U1290 ( .A(n855), .B(n856), .Z(n22544) );
  NANDN U1291 ( .A(n22685), .B(n2173), .Z(n857) );
  NANDN U1292 ( .A(n22664), .B(n2174), .Z(n858) );
  AND U1293 ( .A(n857), .B(n858), .Z(n22691) );
  NANDN U1294 ( .A(n22832), .B(n2173), .Z(n859) );
  NANDN U1295 ( .A(n22811), .B(n2174), .Z(n860) );
  AND U1296 ( .A(n859), .B(n860), .Z(n22838) );
  NANDN U1297 ( .A(n22979), .B(n2173), .Z(n861) );
  NANDN U1298 ( .A(n22958), .B(n2174), .Z(n862) );
  AND U1299 ( .A(n861), .B(n862), .Z(n22985) );
  NANDN U1300 ( .A(n23126), .B(n2173), .Z(n863) );
  NANDN U1301 ( .A(n23105), .B(n2174), .Z(n864) );
  AND U1302 ( .A(n863), .B(n864), .Z(n23132) );
  NANDN U1303 ( .A(n23273), .B(n2173), .Z(n865) );
  NANDN U1304 ( .A(n23252), .B(n2174), .Z(n866) );
  AND U1305 ( .A(n865), .B(n866), .Z(n23279) );
  NANDN U1306 ( .A(n23420), .B(n2173), .Z(n867) );
  NANDN U1307 ( .A(n23399), .B(n2174), .Z(n868) );
  AND U1308 ( .A(n867), .B(n868), .Z(n23426) );
  NANDN U1309 ( .A(n23567), .B(n2173), .Z(n869) );
  NANDN U1310 ( .A(n23546), .B(n2174), .Z(n870) );
  AND U1311 ( .A(n869), .B(n870), .Z(n23573) );
  NANDN U1312 ( .A(n2520), .B(n2173), .Z(n871) );
  NANDN U1313 ( .A(n2499), .B(n2174), .Z(n872) );
  AND U1314 ( .A(n871), .B(n872), .Z(n2526) );
  NANDN U1315 ( .A(n2667), .B(n2173), .Z(n873) );
  NANDN U1316 ( .A(n2646), .B(n2174), .Z(n874) );
  AND U1317 ( .A(n873), .B(n874), .Z(n2673) );
  NANDN U1318 ( .A(n2814), .B(n2173), .Z(n875) );
  NANDN U1319 ( .A(n2793), .B(n2174), .Z(n876) );
  AND U1320 ( .A(n875), .B(n876), .Z(n2820) );
  NANDN U1321 ( .A(n2961), .B(n2173), .Z(n877) );
  NANDN U1322 ( .A(n2940), .B(n2174), .Z(n878) );
  AND U1323 ( .A(n877), .B(n878), .Z(n2967) );
  NANDN U1324 ( .A(n3108), .B(n2173), .Z(n879) );
  NANDN U1325 ( .A(n3087), .B(n2174), .Z(n880) );
  AND U1326 ( .A(n879), .B(n880), .Z(n3114) );
  NANDN U1327 ( .A(n3255), .B(n2173), .Z(n881) );
  NANDN U1328 ( .A(n3234), .B(n2174), .Z(n882) );
  AND U1329 ( .A(n881), .B(n882), .Z(n3261) );
  NANDN U1330 ( .A(n3402), .B(n2173), .Z(n883) );
  NANDN U1331 ( .A(n3381), .B(n2174), .Z(n884) );
  AND U1332 ( .A(n883), .B(n884), .Z(n3408) );
  NANDN U1333 ( .A(n3549), .B(n2173), .Z(n885) );
  NANDN U1334 ( .A(n3528), .B(n2174), .Z(n886) );
  AND U1335 ( .A(n885), .B(n886), .Z(n3555) );
  NANDN U1336 ( .A(n3696), .B(n2173), .Z(n887) );
  NANDN U1337 ( .A(n3675), .B(n2174), .Z(n888) );
  AND U1338 ( .A(n887), .B(n888), .Z(n3702) );
  NANDN U1339 ( .A(n3843), .B(n2173), .Z(n889) );
  NANDN U1340 ( .A(n3822), .B(n2174), .Z(n890) );
  AND U1341 ( .A(n889), .B(n890), .Z(n3849) );
  NANDN U1342 ( .A(n3990), .B(n2173), .Z(n891) );
  NANDN U1343 ( .A(n3969), .B(n2174), .Z(n892) );
  AND U1344 ( .A(n891), .B(n892), .Z(n3996) );
  NANDN U1345 ( .A(n4137), .B(n2173), .Z(n893) );
  NANDN U1346 ( .A(n4116), .B(n2174), .Z(n894) );
  AND U1347 ( .A(n893), .B(n894), .Z(n4143) );
  NANDN U1348 ( .A(n4284), .B(n2173), .Z(n895) );
  NANDN U1349 ( .A(n4263), .B(n2174), .Z(n896) );
  AND U1350 ( .A(n895), .B(n896), .Z(n4290) );
  NANDN U1351 ( .A(n4427), .B(n2173), .Z(n897) );
  NANDN U1352 ( .A(n4408), .B(n2174), .Z(n898) );
  AND U1353 ( .A(n897), .B(n898), .Z(n4433) );
  NANDN U1354 ( .A(n4574), .B(n2173), .Z(n899) );
  NANDN U1355 ( .A(n4553), .B(n2174), .Z(n900) );
  AND U1356 ( .A(n899), .B(n900), .Z(n4580) );
  NANDN U1357 ( .A(n4721), .B(n2173), .Z(n901) );
  NANDN U1358 ( .A(n4700), .B(n2174), .Z(n902) );
  AND U1359 ( .A(n901), .B(n902), .Z(n4727) );
  NANDN U1360 ( .A(n4868), .B(n2173), .Z(n903) );
  NANDN U1361 ( .A(n4847), .B(n2174), .Z(n904) );
  AND U1362 ( .A(n903), .B(n904), .Z(n4874) );
  NANDN U1363 ( .A(n5015), .B(n2173), .Z(n905) );
  NANDN U1364 ( .A(n4994), .B(n2174), .Z(n906) );
  AND U1365 ( .A(n905), .B(n906), .Z(n5021) );
  NANDN U1366 ( .A(n5162), .B(n2173), .Z(n907) );
  NANDN U1367 ( .A(n5141), .B(n2174), .Z(n908) );
  AND U1368 ( .A(n907), .B(n908), .Z(n5168) );
  NANDN U1369 ( .A(n5309), .B(n2173), .Z(n909) );
  NANDN U1370 ( .A(n5288), .B(n2174), .Z(n910) );
  AND U1371 ( .A(n909), .B(n910), .Z(n5315) );
  NANDN U1372 ( .A(n5456), .B(n2173), .Z(n911) );
  NANDN U1373 ( .A(n5435), .B(n2174), .Z(n912) );
  AND U1374 ( .A(n911), .B(n912), .Z(n5462) );
  NANDN U1375 ( .A(n5603), .B(n2173), .Z(n913) );
  NANDN U1376 ( .A(n5582), .B(n2174), .Z(n914) );
  AND U1377 ( .A(n913), .B(n914), .Z(n5609) );
  NANDN U1378 ( .A(n5750), .B(n2173), .Z(n915) );
  NANDN U1379 ( .A(n5729), .B(n2174), .Z(n916) );
  AND U1380 ( .A(n915), .B(n916), .Z(n5756) );
  NANDN U1381 ( .A(n5897), .B(n2173), .Z(n917) );
  NANDN U1382 ( .A(n5876), .B(n2174), .Z(n918) );
  AND U1383 ( .A(n917), .B(n918), .Z(n5903) );
  NANDN U1384 ( .A(n6044), .B(n2173), .Z(n919) );
  NANDN U1385 ( .A(n6023), .B(n2174), .Z(n920) );
  AND U1386 ( .A(n919), .B(n920), .Z(n6050) );
  NANDN U1387 ( .A(n6191), .B(n2173), .Z(n921) );
  NANDN U1388 ( .A(n6170), .B(n2174), .Z(n922) );
  AND U1389 ( .A(n921), .B(n922), .Z(n6197) );
  NANDN U1390 ( .A(n6338), .B(n2173), .Z(n923) );
  NANDN U1391 ( .A(n6317), .B(n2174), .Z(n924) );
  AND U1392 ( .A(n923), .B(n924), .Z(n6344) );
  NANDN U1393 ( .A(n6481), .B(n2173), .Z(n925) );
  NANDN U1394 ( .A(n6460), .B(n2174), .Z(n926) );
  AND U1395 ( .A(n925), .B(n926), .Z(n6487) );
  NANDN U1396 ( .A(n6628), .B(n2173), .Z(n927) );
  NANDN U1397 ( .A(n6607), .B(n2174), .Z(n928) );
  AND U1398 ( .A(n927), .B(n928), .Z(n6634) );
  NANDN U1399 ( .A(n6775), .B(n2173), .Z(n929) );
  NANDN U1400 ( .A(n6754), .B(n2174), .Z(n930) );
  AND U1401 ( .A(n929), .B(n930), .Z(n6781) );
  NANDN U1402 ( .A(n6918), .B(n2173), .Z(n931) );
  NANDN U1403 ( .A(n6897), .B(n2174), .Z(n932) );
  AND U1404 ( .A(n931), .B(n932), .Z(n6924) );
  NANDN U1405 ( .A(n7082), .B(n2173), .Z(n933) );
  NANDN U1406 ( .A(n7061), .B(n2174), .Z(n934) );
  AND U1407 ( .A(n933), .B(n934), .Z(n7088) );
  NANDN U1408 ( .A(n7204), .B(n2173), .Z(n935) );
  NANDN U1409 ( .A(n7183), .B(n2174), .Z(n936) );
  AND U1410 ( .A(n935), .B(n936), .Z(n7210) );
  NANDN U1411 ( .A(n7351), .B(n2173), .Z(n937) );
  NANDN U1412 ( .A(n7330), .B(n2174), .Z(n938) );
  AND U1413 ( .A(n937), .B(n938), .Z(n7357) );
  NANDN U1414 ( .A(n7519), .B(n2173), .Z(n939) );
  NANDN U1415 ( .A(n7498), .B(n2174), .Z(n940) );
  AND U1416 ( .A(n939), .B(n940), .Z(n7525) );
  NANDN U1417 ( .A(n7641), .B(n2173), .Z(n941) );
  NANDN U1418 ( .A(n7620), .B(n2174), .Z(n942) );
  AND U1419 ( .A(n941), .B(n942), .Z(n7647) );
  NANDN U1420 ( .A(n7788), .B(n2173), .Z(n943) );
  NANDN U1421 ( .A(n7767), .B(n2174), .Z(n944) );
  AND U1422 ( .A(n943), .B(n944), .Z(n7794) );
  NANDN U1423 ( .A(n7929), .B(n2173), .Z(n945) );
  NANDN U1424 ( .A(n7910), .B(n2174), .Z(n946) );
  AND U1425 ( .A(n945), .B(n946), .Z(n7936) );
  NANDN U1426 ( .A(n8074), .B(n2173), .Z(n947) );
  NANDN U1427 ( .A(n8053), .B(n2174), .Z(n948) );
  AND U1428 ( .A(n947), .B(n948), .Z(n8080) );
  NANDN U1429 ( .A(n8217), .B(n2173), .Z(n949) );
  NANDN U1430 ( .A(n8198), .B(n2174), .Z(n950) );
  AND U1431 ( .A(n949), .B(n950), .Z(n8223) );
  NANDN U1432 ( .A(n8364), .B(n2173), .Z(n951) );
  NANDN U1433 ( .A(n8343), .B(n2174), .Z(n952) );
  AND U1434 ( .A(n951), .B(n952), .Z(n8370) );
  NANDN U1435 ( .A(n8511), .B(n2173), .Z(n953) );
  NANDN U1436 ( .A(n8490), .B(n2174), .Z(n954) );
  AND U1437 ( .A(n953), .B(n954), .Z(n8517) );
  NANDN U1438 ( .A(n8658), .B(n2173), .Z(n955) );
  NANDN U1439 ( .A(n8637), .B(n2174), .Z(n956) );
  AND U1440 ( .A(n955), .B(n956), .Z(n8664) );
  NANDN U1441 ( .A(n8805), .B(n2173), .Z(n957) );
  NANDN U1442 ( .A(n8784), .B(n2174), .Z(n958) );
  AND U1443 ( .A(n957), .B(n958), .Z(n8811) );
  NANDN U1444 ( .A(n8952), .B(n2173), .Z(n959) );
  NANDN U1445 ( .A(n8931), .B(n2174), .Z(n960) );
  AND U1446 ( .A(n959), .B(n960), .Z(n8958) );
  NANDN U1447 ( .A(n9095), .B(n2173), .Z(n961) );
  NANDN U1448 ( .A(n9074), .B(n2174), .Z(n962) );
  AND U1449 ( .A(n961), .B(n962), .Z(n9101) );
  NANDN U1450 ( .A(n9238), .B(n2173), .Z(n963) );
  NANDN U1451 ( .A(n9217), .B(n2174), .Z(n964) );
  AND U1452 ( .A(n963), .B(n964), .Z(n9244) );
  NANDN U1453 ( .A(n9385), .B(n2173), .Z(n965) );
  NANDN U1454 ( .A(n9364), .B(n2174), .Z(n966) );
  AND U1455 ( .A(n965), .B(n966), .Z(n9391) );
  NANDN U1456 ( .A(n9532), .B(n2173), .Z(n967) );
  NANDN U1457 ( .A(n9511), .B(n2174), .Z(n968) );
  AND U1458 ( .A(n967), .B(n968), .Z(n9538) );
  NANDN U1459 ( .A(n9679), .B(n2173), .Z(n969) );
  NANDN U1460 ( .A(n9658), .B(n2174), .Z(n970) );
  AND U1461 ( .A(n969), .B(n970), .Z(n9685) );
  NANDN U1462 ( .A(n9826), .B(n2173), .Z(n971) );
  NANDN U1463 ( .A(n9805), .B(n2174), .Z(n972) );
  AND U1464 ( .A(n971), .B(n972), .Z(n9832) );
  NANDN U1465 ( .A(n9973), .B(n2173), .Z(n973) );
  NANDN U1466 ( .A(n9952), .B(n2174), .Z(n974) );
  AND U1467 ( .A(n973), .B(n974), .Z(n9979) );
  NANDN U1468 ( .A(n10120), .B(n2173), .Z(n975) );
  NANDN U1469 ( .A(n10099), .B(n2174), .Z(n976) );
  AND U1470 ( .A(n975), .B(n976), .Z(n10126) );
  NANDN U1471 ( .A(n10267), .B(n2173), .Z(n977) );
  NANDN U1472 ( .A(n10246), .B(n2174), .Z(n978) );
  AND U1473 ( .A(n977), .B(n978), .Z(n10273) );
  NANDN U1474 ( .A(n10414), .B(n2173), .Z(n979) );
  NANDN U1475 ( .A(n10393), .B(n2174), .Z(n980) );
  AND U1476 ( .A(n979), .B(n980), .Z(n10420) );
  NANDN U1477 ( .A(n10561), .B(n2173), .Z(n981) );
  NANDN U1478 ( .A(n10540), .B(n2174), .Z(n982) );
  AND U1479 ( .A(n981), .B(n982), .Z(n10567) );
  NANDN U1480 ( .A(n10708), .B(n2173), .Z(n983) );
  NANDN U1481 ( .A(n10687), .B(n2174), .Z(n984) );
  AND U1482 ( .A(n983), .B(n984), .Z(n10714) );
  NANDN U1483 ( .A(n10855), .B(n2173), .Z(n985) );
  NANDN U1484 ( .A(n10834), .B(n2174), .Z(n986) );
  AND U1485 ( .A(n985), .B(n986), .Z(n10861) );
  NANDN U1486 ( .A(n11002), .B(n2173), .Z(n987) );
  NANDN U1487 ( .A(n10981), .B(n2174), .Z(n988) );
  AND U1488 ( .A(n987), .B(n988), .Z(n11008) );
  NANDN U1489 ( .A(n11149), .B(n2173), .Z(n989) );
  NANDN U1490 ( .A(n11128), .B(n2174), .Z(n990) );
  AND U1491 ( .A(n989), .B(n990), .Z(n11155) );
  NANDN U1492 ( .A(n11296), .B(n2173), .Z(n991) );
  NANDN U1493 ( .A(n11275), .B(n2174), .Z(n992) );
  AND U1494 ( .A(n991), .B(n992), .Z(n11302) );
  NANDN U1495 ( .A(n11443), .B(n2173), .Z(n993) );
  NANDN U1496 ( .A(n11422), .B(n2174), .Z(n994) );
  AND U1497 ( .A(n993), .B(n994), .Z(n11449) );
  NANDN U1498 ( .A(n11590), .B(n2173), .Z(n995) );
  NANDN U1499 ( .A(n11569), .B(n2174), .Z(n996) );
  AND U1500 ( .A(n995), .B(n996), .Z(n11596) );
  NANDN U1501 ( .A(n11737), .B(n2173), .Z(n997) );
  NANDN U1502 ( .A(n11716), .B(n2174), .Z(n998) );
  AND U1503 ( .A(n997), .B(n998), .Z(n11743) );
  NANDN U1504 ( .A(n11876), .B(n2173), .Z(n999) );
  NANDN U1505 ( .A(n11855), .B(n2174), .Z(n1000) );
  AND U1506 ( .A(n999), .B(n1000), .Z(n11882) );
  NANDN U1507 ( .A(n12023), .B(n2173), .Z(n1001) );
  NANDN U1508 ( .A(n12002), .B(n2174), .Z(n1002) );
  AND U1509 ( .A(n1001), .B(n1002), .Z(n12029) );
  NANDN U1510 ( .A(n12170), .B(n2173), .Z(n1003) );
  NANDN U1511 ( .A(n12149), .B(n2174), .Z(n1004) );
  AND U1512 ( .A(n1003), .B(n1004), .Z(n12176) );
  NANDN U1513 ( .A(n12317), .B(n2173), .Z(n1005) );
  NANDN U1514 ( .A(n12296), .B(n2174), .Z(n1006) );
  AND U1515 ( .A(n1005), .B(n1006), .Z(n12323) );
  NANDN U1516 ( .A(n12464), .B(n2173), .Z(n1007) );
  NANDN U1517 ( .A(n12443), .B(n2174), .Z(n1008) );
  AND U1518 ( .A(n1007), .B(n1008), .Z(n12470) );
  NANDN U1519 ( .A(n12632), .B(n2173), .Z(n1009) );
  NANDN U1520 ( .A(n12611), .B(n2174), .Z(n1010) );
  AND U1521 ( .A(n1009), .B(n1010), .Z(n12638) );
  NANDN U1522 ( .A(n12754), .B(n2173), .Z(n1011) );
  NANDN U1523 ( .A(n12733), .B(n2174), .Z(n1012) );
  AND U1524 ( .A(n1011), .B(n1012), .Z(n12760) );
  NANDN U1525 ( .A(n12901), .B(n2173), .Z(n1013) );
  NANDN U1526 ( .A(n12880), .B(n2174), .Z(n1014) );
  AND U1527 ( .A(n1013), .B(n1014), .Z(n12907) );
  NANDN U1528 ( .A(n13048), .B(n2173), .Z(n1015) );
  NANDN U1529 ( .A(n13027), .B(n2174), .Z(n1016) );
  AND U1530 ( .A(n1015), .B(n1016), .Z(n13054) );
  NANDN U1531 ( .A(n13195), .B(n2173), .Z(n1017) );
  NANDN U1532 ( .A(n13174), .B(n2174), .Z(n1018) );
  AND U1533 ( .A(n1017), .B(n1018), .Z(n13201) );
  NANDN U1534 ( .A(n13342), .B(n2173), .Z(n1019) );
  NANDN U1535 ( .A(n13321), .B(n2174), .Z(n1020) );
  AND U1536 ( .A(n1019), .B(n1020), .Z(n13348) );
  NANDN U1537 ( .A(n13489), .B(n2173), .Z(n1021) );
  NANDN U1538 ( .A(n13468), .B(n2174), .Z(n1022) );
  AND U1539 ( .A(n1021), .B(n1022), .Z(n13495) );
  NANDN U1540 ( .A(n13636), .B(n2173), .Z(n1023) );
  NANDN U1541 ( .A(n13615), .B(n2174), .Z(n1024) );
  AND U1542 ( .A(n1023), .B(n1024), .Z(n13642) );
  NANDN U1543 ( .A(n13804), .B(n2173), .Z(n1025) );
  NANDN U1544 ( .A(n13783), .B(n2174), .Z(n1026) );
  AND U1545 ( .A(n1025), .B(n1026), .Z(n13810) );
  NANDN U1546 ( .A(n13926), .B(n2173), .Z(n1027) );
  NANDN U1547 ( .A(n13905), .B(n2174), .Z(n1028) );
  AND U1548 ( .A(n1027), .B(n1028), .Z(n13932) );
  NANDN U1549 ( .A(n14073), .B(n2173), .Z(n1029) );
  NANDN U1550 ( .A(n14052), .B(n2174), .Z(n1030) );
  AND U1551 ( .A(n1029), .B(n1030), .Z(n14079) );
  NANDN U1552 ( .A(n14220), .B(n2173), .Z(n1031) );
  NANDN U1553 ( .A(n14199), .B(n2174), .Z(n1032) );
  AND U1554 ( .A(n1031), .B(n1032), .Z(n14226) );
  NANDN U1555 ( .A(n14367), .B(n2173), .Z(n1033) );
  NANDN U1556 ( .A(n14346), .B(n2174), .Z(n1034) );
  AND U1557 ( .A(n1033), .B(n1034), .Z(n14373) );
  NANDN U1558 ( .A(n14514), .B(n2173), .Z(n1035) );
  NANDN U1559 ( .A(n14493), .B(n2174), .Z(n1036) );
  AND U1560 ( .A(n1035), .B(n1036), .Z(n14520) );
  NANDN U1561 ( .A(n14661), .B(n2173), .Z(n1037) );
  NANDN U1562 ( .A(n14640), .B(n2174), .Z(n1038) );
  AND U1563 ( .A(n1037), .B(n1038), .Z(n14667) );
  NANDN U1564 ( .A(n14804), .B(n2173), .Z(n1039) );
  NANDN U1565 ( .A(n14783), .B(n2174), .Z(n1040) );
  AND U1566 ( .A(n1039), .B(n1040), .Z(n14810) );
  NANDN U1567 ( .A(n14951), .B(n2173), .Z(n1041) );
  NANDN U1568 ( .A(n14930), .B(n2174), .Z(n1042) );
  AND U1569 ( .A(n1041), .B(n1042), .Z(n14957) );
  NANDN U1570 ( .A(n15098), .B(n2173), .Z(n1043) );
  NANDN U1571 ( .A(n15077), .B(n2174), .Z(n1044) );
  AND U1572 ( .A(n1043), .B(n1044), .Z(n15104) );
  NANDN U1573 ( .A(n15245), .B(n2173), .Z(n1045) );
  NANDN U1574 ( .A(n15224), .B(n2174), .Z(n1046) );
  AND U1575 ( .A(n1045), .B(n1046), .Z(n15251) );
  NANDN U1576 ( .A(n15392), .B(n2173), .Z(n1047) );
  NANDN U1577 ( .A(n15371), .B(n2174), .Z(n1048) );
  AND U1578 ( .A(n1047), .B(n1048), .Z(n15398) );
  NANDN U1579 ( .A(n15539), .B(n2173), .Z(n1049) );
  NANDN U1580 ( .A(n15518), .B(n2174), .Z(n1050) );
  AND U1581 ( .A(n1049), .B(n1050), .Z(n15545) );
  NANDN U1582 ( .A(n15682), .B(n2173), .Z(n1051) );
  NANDN U1583 ( .A(n15661), .B(n2174), .Z(n1052) );
  AND U1584 ( .A(n1051), .B(n1052), .Z(n15688) );
  NANDN U1585 ( .A(n15829), .B(n2173), .Z(n1053) );
  NANDN U1586 ( .A(n15808), .B(n2174), .Z(n1054) );
  AND U1587 ( .A(n1053), .B(n1054), .Z(n15835) );
  NANDN U1588 ( .A(n15976), .B(n2173), .Z(n1055) );
  NANDN U1589 ( .A(n15955), .B(n2174), .Z(n1056) );
  AND U1590 ( .A(n1055), .B(n1056), .Z(n15982) );
  NANDN U1591 ( .A(n16123), .B(n2173), .Z(n1057) );
  NANDN U1592 ( .A(n16102), .B(n2174), .Z(n1058) );
  AND U1593 ( .A(n1057), .B(n1058), .Z(n16129) );
  NANDN U1594 ( .A(n16270), .B(n2173), .Z(n1059) );
  NANDN U1595 ( .A(n16249), .B(n2174), .Z(n1060) );
  AND U1596 ( .A(n1059), .B(n1060), .Z(n16276) );
  NANDN U1597 ( .A(n16417), .B(n2173), .Z(n1061) );
  NANDN U1598 ( .A(n16396), .B(n2174), .Z(n1062) );
  AND U1599 ( .A(n1061), .B(n1062), .Z(n16423) );
  NANDN U1600 ( .A(n16564), .B(n2173), .Z(n1063) );
  NANDN U1601 ( .A(n16543), .B(n2174), .Z(n1064) );
  AND U1602 ( .A(n1063), .B(n1064), .Z(n16570) );
  NANDN U1603 ( .A(n16711), .B(n2173), .Z(n1065) );
  NANDN U1604 ( .A(n16690), .B(n2174), .Z(n1066) );
  AND U1605 ( .A(n1065), .B(n1066), .Z(n16717) );
  NANDN U1606 ( .A(n16858), .B(n2173), .Z(n1067) );
  NANDN U1607 ( .A(n16837), .B(n2174), .Z(n1068) );
  AND U1608 ( .A(n1067), .B(n1068), .Z(n16864) );
  NANDN U1609 ( .A(n17005), .B(n2173), .Z(n1069) );
  NANDN U1610 ( .A(n16984), .B(n2174), .Z(n1070) );
  AND U1611 ( .A(n1069), .B(n1070), .Z(n17011) );
  NANDN U1612 ( .A(n17152), .B(n2173), .Z(n1071) );
  NANDN U1613 ( .A(n17131), .B(n2174), .Z(n1072) );
  AND U1614 ( .A(n1071), .B(n1072), .Z(n17158) );
  NANDN U1615 ( .A(n17299), .B(n2173), .Z(n1073) );
  NANDN U1616 ( .A(n17278), .B(n2174), .Z(n1074) );
  AND U1617 ( .A(n1073), .B(n1074), .Z(n17305) );
  NANDN U1618 ( .A(n17446), .B(n2173), .Z(n1075) );
  NANDN U1619 ( .A(n17425), .B(n2174), .Z(n1076) );
  AND U1620 ( .A(n1075), .B(n1076), .Z(n17452) );
  NANDN U1621 ( .A(n17593), .B(n2173), .Z(n1077) );
  NANDN U1622 ( .A(n17572), .B(n2174), .Z(n1078) );
  AND U1623 ( .A(n1077), .B(n1078), .Z(n17599) );
  NANDN U1624 ( .A(n17757), .B(n2173), .Z(n1079) );
  NANDN U1625 ( .A(n17738), .B(n2174), .Z(n1080) );
  AND U1626 ( .A(n1079), .B(n1080), .Z(n17763) );
  NANDN U1627 ( .A(n17879), .B(n2173), .Z(n1081) );
  NANDN U1628 ( .A(n17858), .B(n2174), .Z(n1082) );
  AND U1629 ( .A(n1081), .B(n1082), .Z(n17885) );
  NANDN U1630 ( .A(n18026), .B(n2173), .Z(n1083) );
  NANDN U1631 ( .A(n18005), .B(n2174), .Z(n1084) );
  AND U1632 ( .A(n1083), .B(n1084), .Z(n18032) );
  NANDN U1633 ( .A(n18169), .B(n2173), .Z(n1085) );
  NANDN U1634 ( .A(n18148), .B(n2174), .Z(n1086) );
  AND U1635 ( .A(n1085), .B(n1086), .Z(n18175) );
  NANDN U1636 ( .A(n18316), .B(n2173), .Z(n1087) );
  NANDN U1637 ( .A(n18295), .B(n2174), .Z(n1088) );
  AND U1638 ( .A(n1087), .B(n1088), .Z(n18322) );
  NANDN U1639 ( .A(n18463), .B(n2173), .Z(n1089) );
  NANDN U1640 ( .A(n18442), .B(n2174), .Z(n1090) );
  AND U1641 ( .A(n1089), .B(n1090), .Z(n18469) );
  NANDN U1642 ( .A(n18610), .B(n2173), .Z(n1091) );
  NANDN U1643 ( .A(n18589), .B(n2174), .Z(n1092) );
  AND U1644 ( .A(n1091), .B(n1092), .Z(n18616) );
  NANDN U1645 ( .A(n18757), .B(n2173), .Z(n1093) );
  NANDN U1646 ( .A(n18736), .B(n2174), .Z(n1094) );
  AND U1647 ( .A(n1093), .B(n1094), .Z(n18763) );
  NANDN U1648 ( .A(n18904), .B(n2173), .Z(n1095) );
  NANDN U1649 ( .A(n18883), .B(n2174), .Z(n1096) );
  AND U1650 ( .A(n1095), .B(n1096), .Z(n18910) );
  NANDN U1651 ( .A(n19051), .B(n2173), .Z(n1097) );
  NANDN U1652 ( .A(n19030), .B(n2174), .Z(n1098) );
  AND U1653 ( .A(n1097), .B(n1098), .Z(n19057) );
  NANDN U1654 ( .A(n19198), .B(n2173), .Z(n1099) );
  NANDN U1655 ( .A(n19177), .B(n2174), .Z(n1100) );
  AND U1656 ( .A(n1099), .B(n1100), .Z(n19204) );
  NANDN U1657 ( .A(n19345), .B(n2173), .Z(n1101) );
  NANDN U1658 ( .A(n19324), .B(n2174), .Z(n1102) );
  AND U1659 ( .A(n1101), .B(n1102), .Z(n19351) );
  NANDN U1660 ( .A(n19492), .B(n2173), .Z(n1103) );
  NANDN U1661 ( .A(n19471), .B(n2174), .Z(n1104) );
  AND U1662 ( .A(n1103), .B(n1104), .Z(n19498) );
  NANDN U1663 ( .A(n19639), .B(n2173), .Z(n1105) );
  NANDN U1664 ( .A(n19618), .B(n2174), .Z(n1106) );
  AND U1665 ( .A(n1105), .B(n1106), .Z(n19645) );
  NANDN U1666 ( .A(n19782), .B(n2173), .Z(n1107) );
  NANDN U1667 ( .A(n19761), .B(n2174), .Z(n1108) );
  AND U1668 ( .A(n1107), .B(n1108), .Z(n19788) );
  NANDN U1669 ( .A(n19929), .B(n2173), .Z(n1109) );
  NANDN U1670 ( .A(n19908), .B(n2174), .Z(n1110) );
  AND U1671 ( .A(n1109), .B(n1110), .Z(n19935) );
  NANDN U1672 ( .A(n20076), .B(n2173), .Z(n1111) );
  NANDN U1673 ( .A(n20055), .B(n2174), .Z(n1112) );
  AND U1674 ( .A(n1111), .B(n1112), .Z(n20082) );
  NANDN U1675 ( .A(n20219), .B(n2173), .Z(n1113) );
  NANDN U1676 ( .A(n20198), .B(n2174), .Z(n1114) );
  AND U1677 ( .A(n1113), .B(n1114), .Z(n20225) );
  NANDN U1678 ( .A(n20366), .B(n2173), .Z(n1115) );
  NANDN U1679 ( .A(n20345), .B(n2174), .Z(n1116) );
  AND U1680 ( .A(n1115), .B(n1116), .Z(n20372) );
  NANDN U1681 ( .A(n20513), .B(n2173), .Z(n1117) );
  NANDN U1682 ( .A(n20492), .B(n2174), .Z(n1118) );
  AND U1683 ( .A(n1117), .B(n1118), .Z(n20519) );
  NANDN U1684 ( .A(n20660), .B(n2173), .Z(n1119) );
  NANDN U1685 ( .A(n20639), .B(n2174), .Z(n1120) );
  AND U1686 ( .A(n1119), .B(n1120), .Z(n20666) );
  NANDN U1687 ( .A(n20807), .B(n2173), .Z(n1121) );
  NANDN U1688 ( .A(n20786), .B(n2174), .Z(n1122) );
  AND U1689 ( .A(n1121), .B(n1122), .Z(n20813) );
  NANDN U1690 ( .A(n20954), .B(n2173), .Z(n1123) );
  NANDN U1691 ( .A(n20933), .B(n2174), .Z(n1124) );
  AND U1692 ( .A(n1123), .B(n1124), .Z(n20960) );
  NANDN U1693 ( .A(n21097), .B(n2173), .Z(n1125) );
  NANDN U1694 ( .A(n21076), .B(n2174), .Z(n1126) );
  AND U1695 ( .A(n1125), .B(n1126), .Z(n21103) );
  NANDN U1696 ( .A(n21265), .B(n2173), .Z(n1127) );
  NANDN U1697 ( .A(n21244), .B(n2174), .Z(n1128) );
  AND U1698 ( .A(n1127), .B(n1128), .Z(n21271) );
  NANDN U1699 ( .A(n21387), .B(n2173), .Z(n1129) );
  NANDN U1700 ( .A(n21366), .B(n2174), .Z(n1130) );
  AND U1701 ( .A(n1129), .B(n1130), .Z(n21393) );
  NANDN U1702 ( .A(n21534), .B(n2173), .Z(n1131) );
  NANDN U1703 ( .A(n21513), .B(n2174), .Z(n1132) );
  AND U1704 ( .A(n1131), .B(n1132), .Z(n21540) );
  NANDN U1705 ( .A(n21681), .B(n2173), .Z(n1133) );
  NANDN U1706 ( .A(n21660), .B(n2174), .Z(n1134) );
  AND U1707 ( .A(n1133), .B(n1134), .Z(n21687) );
  NANDN U1708 ( .A(n21828), .B(n2173), .Z(n1135) );
  NANDN U1709 ( .A(n21807), .B(n2174), .Z(n1136) );
  AND U1710 ( .A(n1135), .B(n1136), .Z(n21834) );
  NANDN U1711 ( .A(n21975), .B(n2173), .Z(n1137) );
  NANDN U1712 ( .A(n21954), .B(n2174), .Z(n1138) );
  AND U1713 ( .A(n1137), .B(n1138), .Z(n21981) );
  NANDN U1714 ( .A(n22122), .B(n2173), .Z(n1139) );
  NANDN U1715 ( .A(n22101), .B(n2174), .Z(n1140) );
  AND U1716 ( .A(n1139), .B(n1140), .Z(n22128) );
  NANDN U1717 ( .A(n22269), .B(n2173), .Z(n1141) );
  NANDN U1718 ( .A(n22248), .B(n2174), .Z(n1142) );
  AND U1719 ( .A(n1141), .B(n1142), .Z(n22275) );
  NANDN U1720 ( .A(n22412), .B(n2173), .Z(n1143) );
  NANDN U1721 ( .A(n22391), .B(n2174), .Z(n1144) );
  AND U1722 ( .A(n1143), .B(n1144), .Z(n22418) );
  NANDN U1723 ( .A(n22559), .B(n2173), .Z(n1145) );
  NANDN U1724 ( .A(n22538), .B(n2174), .Z(n1146) );
  AND U1725 ( .A(n1145), .B(n1146), .Z(n22565) );
  NANDN U1726 ( .A(n22706), .B(n2173), .Z(n1147) );
  NANDN U1727 ( .A(n22685), .B(n2174), .Z(n1148) );
  AND U1728 ( .A(n1147), .B(n1148), .Z(n22712) );
  NANDN U1729 ( .A(n22853), .B(n2173), .Z(n1149) );
  NANDN U1730 ( .A(n22832), .B(n2174), .Z(n1150) );
  AND U1731 ( .A(n1149), .B(n1150), .Z(n22859) );
  NANDN U1732 ( .A(n23000), .B(n2173), .Z(n1151) );
  NANDN U1733 ( .A(n22979), .B(n2174), .Z(n1152) );
  AND U1734 ( .A(n1151), .B(n1152), .Z(n23006) );
  NANDN U1735 ( .A(n23147), .B(n2173), .Z(n1153) );
  NANDN U1736 ( .A(n23126), .B(n2174), .Z(n1154) );
  AND U1737 ( .A(n1153), .B(n1154), .Z(n23153) );
  NANDN U1738 ( .A(n23294), .B(n2173), .Z(n1155) );
  NANDN U1739 ( .A(n23273), .B(n2174), .Z(n1156) );
  AND U1740 ( .A(n1155), .B(n1156), .Z(n23300) );
  NANDN U1741 ( .A(n23441), .B(n2173), .Z(n1157) );
  NANDN U1742 ( .A(n23420), .B(n2174), .Z(n1158) );
  AND U1743 ( .A(n1157), .B(n1158), .Z(n23447) );
  NANDN U1744 ( .A(n23586), .B(n2173), .Z(n1159) );
  NANDN U1745 ( .A(n23567), .B(n2174), .Z(n1160) );
  AND U1746 ( .A(n1159), .B(n1160), .Z(n23594) );
  NANDN U1747 ( .A(n2394), .B(n2173), .Z(n1161) );
  NANDN U1748 ( .A(n2378), .B(n2174), .Z(n1162) );
  AND U1749 ( .A(n1161), .B(n1162), .Z(n2400) );
  NANDN U1750 ( .A(n2541), .B(n2173), .Z(n1163) );
  NANDN U1751 ( .A(n2520), .B(n2174), .Z(n1164) );
  AND U1752 ( .A(n1163), .B(n1164), .Z(n2547) );
  NANDN U1753 ( .A(n2688), .B(n2173), .Z(n1165) );
  NANDN U1754 ( .A(n2667), .B(n2174), .Z(n1166) );
  AND U1755 ( .A(n1165), .B(n1166), .Z(n2694) );
  NANDN U1756 ( .A(n2835), .B(n2173), .Z(n1167) );
  NANDN U1757 ( .A(n2814), .B(n2174), .Z(n1168) );
  AND U1758 ( .A(n1167), .B(n1168), .Z(n2841) );
  NANDN U1759 ( .A(n2982), .B(n2173), .Z(n1169) );
  NANDN U1760 ( .A(n2961), .B(n2174), .Z(n1170) );
  AND U1761 ( .A(n1169), .B(n1170), .Z(n2988) );
  NANDN U1762 ( .A(n3129), .B(n2173), .Z(n1171) );
  NANDN U1763 ( .A(n3108), .B(n2174), .Z(n1172) );
  AND U1764 ( .A(n1171), .B(n1172), .Z(n3135) );
  NANDN U1765 ( .A(n3276), .B(n2173), .Z(n1173) );
  NANDN U1766 ( .A(n3255), .B(n2174), .Z(n1174) );
  AND U1767 ( .A(n1173), .B(n1174), .Z(n3282) );
  NANDN U1768 ( .A(n3423), .B(n2173), .Z(n1175) );
  NANDN U1769 ( .A(n3402), .B(n2174), .Z(n1176) );
  AND U1770 ( .A(n1175), .B(n1176), .Z(n3429) );
  NANDN U1771 ( .A(n3570), .B(n2173), .Z(n1177) );
  NANDN U1772 ( .A(n3549), .B(n2174), .Z(n1178) );
  AND U1773 ( .A(n1177), .B(n1178), .Z(n3576) );
  NANDN U1774 ( .A(n3717), .B(n2173), .Z(n1179) );
  NANDN U1775 ( .A(n3696), .B(n2174), .Z(n1180) );
  AND U1776 ( .A(n1179), .B(n1180), .Z(n3723) );
  NANDN U1777 ( .A(n3864), .B(n2173), .Z(n1181) );
  NANDN U1778 ( .A(n3843), .B(n2174), .Z(n1182) );
  AND U1779 ( .A(n1181), .B(n1182), .Z(n3870) );
  NANDN U1780 ( .A(n4011), .B(n2173), .Z(n1183) );
  NANDN U1781 ( .A(n3990), .B(n2174), .Z(n1184) );
  AND U1782 ( .A(n1183), .B(n1184), .Z(n4017) );
  NANDN U1783 ( .A(n4158), .B(n2173), .Z(n1185) );
  NANDN U1784 ( .A(n4137), .B(n2174), .Z(n1186) );
  AND U1785 ( .A(n1185), .B(n1186), .Z(n4164) );
  NANDN U1786 ( .A(n4305), .B(n2173), .Z(n1187) );
  NANDN U1787 ( .A(n4284), .B(n2174), .Z(n1188) );
  AND U1788 ( .A(n1187), .B(n1188), .Z(n4311) );
  NANDN U1789 ( .A(n4448), .B(n2173), .Z(n1189) );
  NANDN U1790 ( .A(n4427), .B(n2174), .Z(n1190) );
  AND U1791 ( .A(n1189), .B(n1190), .Z(n4454) );
  NANDN U1792 ( .A(n4595), .B(n2173), .Z(n1191) );
  NANDN U1793 ( .A(n4574), .B(n2174), .Z(n1192) );
  AND U1794 ( .A(n1191), .B(n1192), .Z(n4601) );
  NANDN U1795 ( .A(n4742), .B(n2173), .Z(n1193) );
  NANDN U1796 ( .A(n4721), .B(n2174), .Z(n1194) );
  AND U1797 ( .A(n1193), .B(n1194), .Z(n4748) );
  NANDN U1798 ( .A(n4889), .B(n2173), .Z(n1195) );
  NANDN U1799 ( .A(n4868), .B(n2174), .Z(n1196) );
  AND U1800 ( .A(n1195), .B(n1196), .Z(n4895) );
  NANDN U1801 ( .A(n5036), .B(n2173), .Z(n1197) );
  NANDN U1802 ( .A(n5015), .B(n2174), .Z(n1198) );
  AND U1803 ( .A(n1197), .B(n1198), .Z(n5042) );
  NANDN U1804 ( .A(n5183), .B(n2173), .Z(n1199) );
  NANDN U1805 ( .A(n5162), .B(n2174), .Z(n1200) );
  AND U1806 ( .A(n1199), .B(n1200), .Z(n5189) );
  NANDN U1807 ( .A(n5330), .B(n2173), .Z(n1201) );
  NANDN U1808 ( .A(n5309), .B(n2174), .Z(n1202) );
  AND U1809 ( .A(n1201), .B(n1202), .Z(n5336) );
  NANDN U1810 ( .A(n5477), .B(n2173), .Z(n1203) );
  NANDN U1811 ( .A(n5456), .B(n2174), .Z(n1204) );
  AND U1812 ( .A(n1203), .B(n1204), .Z(n5483) );
  NANDN U1813 ( .A(n5624), .B(n2173), .Z(n1205) );
  NANDN U1814 ( .A(n5603), .B(n2174), .Z(n1206) );
  AND U1815 ( .A(n1205), .B(n1206), .Z(n5630) );
  NANDN U1816 ( .A(n5771), .B(n2173), .Z(n1207) );
  NANDN U1817 ( .A(n5750), .B(n2174), .Z(n1208) );
  AND U1818 ( .A(n1207), .B(n1208), .Z(n5777) );
  NANDN U1819 ( .A(n5918), .B(n2173), .Z(n1209) );
  NANDN U1820 ( .A(n5897), .B(n2174), .Z(n1210) );
  AND U1821 ( .A(n1209), .B(n1210), .Z(n5924) );
  NANDN U1822 ( .A(n6065), .B(n2173), .Z(n1211) );
  NANDN U1823 ( .A(n6044), .B(n2174), .Z(n1212) );
  AND U1824 ( .A(n1211), .B(n1212), .Z(n6071) );
  NANDN U1825 ( .A(n6212), .B(n2173), .Z(n1213) );
  NANDN U1826 ( .A(n6191), .B(n2174), .Z(n1214) );
  AND U1827 ( .A(n1213), .B(n1214), .Z(n6218) );
  NANDN U1828 ( .A(n6359), .B(n2173), .Z(n1215) );
  NANDN U1829 ( .A(n6338), .B(n2174), .Z(n1216) );
  AND U1830 ( .A(n1215), .B(n1216), .Z(n6365) );
  NANDN U1831 ( .A(n6502), .B(n2173), .Z(n1217) );
  NANDN U1832 ( .A(n6481), .B(n2174), .Z(n1218) );
  AND U1833 ( .A(n1217), .B(n1218), .Z(n6508) );
  NANDN U1834 ( .A(n6649), .B(n2173), .Z(n1219) );
  NANDN U1835 ( .A(n6628), .B(n2174), .Z(n1220) );
  AND U1836 ( .A(n1219), .B(n1220), .Z(n6655) );
  NANDN U1837 ( .A(n6817), .B(n2173), .Z(n1221) );
  NANDN U1838 ( .A(n6796), .B(n2174), .Z(n1222) );
  AND U1839 ( .A(n1221), .B(n1222), .Z(n6823) );
  NANDN U1840 ( .A(n6937), .B(n2173), .Z(n1223) );
  NANDN U1841 ( .A(n6918), .B(n2174), .Z(n1224) );
  AND U1842 ( .A(n1223), .B(n1224), .Z(n6944) );
  NANDN U1843 ( .A(n7101), .B(n2173), .Z(n1225) );
  NANDN U1844 ( .A(n7082), .B(n2174), .Z(n1226) );
  AND U1845 ( .A(n1225), .B(n1226), .Z(n7108) );
  NANDN U1846 ( .A(n7225), .B(n2173), .Z(n1227) );
  NANDN U1847 ( .A(n7204), .B(n2174), .Z(n1228) );
  AND U1848 ( .A(n1227), .B(n1228), .Z(n7231) );
  NANDN U1849 ( .A(n7372), .B(n2173), .Z(n1229) );
  NANDN U1850 ( .A(n7351), .B(n2174), .Z(n1230) );
  AND U1851 ( .A(n1229), .B(n1230), .Z(n7378) );
  NANDN U1852 ( .A(n7538), .B(n2173), .Z(n1231) );
  NANDN U1853 ( .A(n7519), .B(n2174), .Z(n1232) );
  AND U1854 ( .A(n1231), .B(n1232), .Z(n7545) );
  NANDN U1855 ( .A(n7662), .B(n2173), .Z(n1233) );
  NANDN U1856 ( .A(n7641), .B(n2174), .Z(n1234) );
  AND U1857 ( .A(n1233), .B(n1234), .Z(n7668) );
  NANDN U1858 ( .A(n7807), .B(n2173), .Z(n1235) );
  NANDN U1859 ( .A(n7788), .B(n2174), .Z(n1236) );
  AND U1860 ( .A(n1235), .B(n1236), .Z(n7814) );
  NANDN U1861 ( .A(n7948), .B(n2173), .Z(n1237) );
  NANDN U1862 ( .A(n7929), .B(n2174), .Z(n1238) );
  AND U1863 ( .A(n1237), .B(n1238), .Z(n7954) );
  NANDN U1864 ( .A(n8095), .B(n2173), .Z(n1239) );
  NANDN U1865 ( .A(n8074), .B(n2174), .Z(n1240) );
  AND U1866 ( .A(n1239), .B(n1240), .Z(n8101) );
  NANDN U1867 ( .A(n8238), .B(n2173), .Z(n1241) );
  NANDN U1868 ( .A(n8217), .B(n2174), .Z(n1242) );
  AND U1869 ( .A(n1241), .B(n1242), .Z(n8244) );
  NANDN U1870 ( .A(n8385), .B(n2173), .Z(n1243) );
  NANDN U1871 ( .A(n8364), .B(n2174), .Z(n1244) );
  AND U1872 ( .A(n1243), .B(n1244), .Z(n8391) );
  NANDN U1873 ( .A(n8532), .B(n2173), .Z(n1245) );
  NANDN U1874 ( .A(n8511), .B(n2174), .Z(n1246) );
  AND U1875 ( .A(n1245), .B(n1246), .Z(n8538) );
  NANDN U1876 ( .A(n8679), .B(n2173), .Z(n1247) );
  NANDN U1877 ( .A(n8658), .B(n2174), .Z(n1248) );
  AND U1878 ( .A(n1247), .B(n1248), .Z(n8685) );
  NANDN U1879 ( .A(n8826), .B(n2173), .Z(n1249) );
  NANDN U1880 ( .A(n8805), .B(n2174), .Z(n1250) );
  AND U1881 ( .A(n1249), .B(n1250), .Z(n8832) );
  NANDN U1882 ( .A(n8973), .B(n2173), .Z(n1251) );
  NANDN U1883 ( .A(n8952), .B(n2174), .Z(n1252) );
  AND U1884 ( .A(n1251), .B(n1252), .Z(n8979) );
  NANDN U1885 ( .A(n9116), .B(n2173), .Z(n1253) );
  NANDN U1886 ( .A(n9095), .B(n2174), .Z(n1254) );
  AND U1887 ( .A(n1253), .B(n1254), .Z(n9122) );
  NANDN U1888 ( .A(n9259), .B(n2173), .Z(n1255) );
  NANDN U1889 ( .A(n9238), .B(n2174), .Z(n1256) );
  AND U1890 ( .A(n1255), .B(n1256), .Z(n9265) );
  NANDN U1891 ( .A(n9406), .B(n2173), .Z(n1257) );
  NANDN U1892 ( .A(n9385), .B(n2174), .Z(n1258) );
  AND U1893 ( .A(n1257), .B(n1258), .Z(n9412) );
  NANDN U1894 ( .A(n9553), .B(n2173), .Z(n1259) );
  NANDN U1895 ( .A(n9532), .B(n2174), .Z(n1260) );
  AND U1896 ( .A(n1259), .B(n1260), .Z(n9559) );
  NANDN U1897 ( .A(n9700), .B(n2173), .Z(n1261) );
  NANDN U1898 ( .A(n9679), .B(n2174), .Z(n1262) );
  AND U1899 ( .A(n1261), .B(n1262), .Z(n9706) );
  NANDN U1900 ( .A(n9847), .B(n2173), .Z(n1263) );
  NANDN U1901 ( .A(n9826), .B(n2174), .Z(n1264) );
  AND U1902 ( .A(n1263), .B(n1264), .Z(n9853) );
  NANDN U1903 ( .A(n9994), .B(n2173), .Z(n1265) );
  NANDN U1904 ( .A(n9973), .B(n2174), .Z(n1266) );
  AND U1905 ( .A(n1265), .B(n1266), .Z(n10000) );
  NANDN U1906 ( .A(n10141), .B(n2173), .Z(n1267) );
  NANDN U1907 ( .A(n10120), .B(n2174), .Z(n1268) );
  AND U1908 ( .A(n1267), .B(n1268), .Z(n10147) );
  NANDN U1909 ( .A(n10288), .B(n2173), .Z(n1269) );
  NANDN U1910 ( .A(n10267), .B(n2174), .Z(n1270) );
  AND U1911 ( .A(n1269), .B(n1270), .Z(n10294) );
  NANDN U1912 ( .A(n10435), .B(n2173), .Z(n1271) );
  NANDN U1913 ( .A(n10414), .B(n2174), .Z(n1272) );
  AND U1914 ( .A(n1271), .B(n1272), .Z(n10441) );
  NANDN U1915 ( .A(n10582), .B(n2173), .Z(n1273) );
  NANDN U1916 ( .A(n10561), .B(n2174), .Z(n1274) );
  AND U1917 ( .A(n1273), .B(n1274), .Z(n10588) );
  NANDN U1918 ( .A(n10729), .B(n2173), .Z(n1275) );
  NANDN U1919 ( .A(n10708), .B(n2174), .Z(n1276) );
  AND U1920 ( .A(n1275), .B(n1276), .Z(n10735) );
  NANDN U1921 ( .A(n10876), .B(n2173), .Z(n1277) );
  NANDN U1922 ( .A(n10855), .B(n2174), .Z(n1278) );
  AND U1923 ( .A(n1277), .B(n1278), .Z(n10882) );
  NANDN U1924 ( .A(n11023), .B(n2173), .Z(n1279) );
  NANDN U1925 ( .A(n11002), .B(n2174), .Z(n1280) );
  AND U1926 ( .A(n1279), .B(n1280), .Z(n11029) );
  NANDN U1927 ( .A(n11170), .B(n2173), .Z(n1281) );
  NANDN U1928 ( .A(n11149), .B(n2174), .Z(n1282) );
  AND U1929 ( .A(n1281), .B(n1282), .Z(n11176) );
  NANDN U1930 ( .A(n11317), .B(n2173), .Z(n1283) );
  NANDN U1931 ( .A(n11296), .B(n2174), .Z(n1284) );
  AND U1932 ( .A(n1283), .B(n1284), .Z(n11323) );
  NANDN U1933 ( .A(n11464), .B(n2173), .Z(n1285) );
  NANDN U1934 ( .A(n11443), .B(n2174), .Z(n1286) );
  AND U1935 ( .A(n1285), .B(n1286), .Z(n11470) );
  NANDN U1936 ( .A(n11611), .B(n2173), .Z(n1287) );
  NANDN U1937 ( .A(n11590), .B(n2174), .Z(n1288) );
  AND U1938 ( .A(n1287), .B(n1288), .Z(n11617) );
  NANDN U1939 ( .A(n11775), .B(n2173), .Z(n1289) );
  NANDN U1940 ( .A(n11756), .B(n2174), .Z(n1290) );
  AND U1941 ( .A(n1289), .B(n1290), .Z(n11781) );
  NANDN U1942 ( .A(n11897), .B(n2173), .Z(n1291) );
  NANDN U1943 ( .A(n11876), .B(n2174), .Z(n1292) );
  AND U1944 ( .A(n1291), .B(n1292), .Z(n11903) );
  NANDN U1945 ( .A(n12044), .B(n2173), .Z(n1293) );
  NANDN U1946 ( .A(n12023), .B(n2174), .Z(n1294) );
  AND U1947 ( .A(n1293), .B(n1294), .Z(n12050) );
  NANDN U1948 ( .A(n12191), .B(n2173), .Z(n1295) );
  NANDN U1949 ( .A(n12170), .B(n2174), .Z(n1296) );
  AND U1950 ( .A(n1295), .B(n1296), .Z(n12197) );
  NANDN U1951 ( .A(n12338), .B(n2173), .Z(n1297) );
  NANDN U1952 ( .A(n12317), .B(n2174), .Z(n1298) );
  AND U1953 ( .A(n1297), .B(n1298), .Z(n12344) );
  NANDN U1954 ( .A(n12485), .B(n2173), .Z(n1299) );
  NANDN U1955 ( .A(n12464), .B(n2174), .Z(n1300) );
  AND U1956 ( .A(n1299), .B(n1300), .Z(n12491) );
  NANDN U1957 ( .A(n12651), .B(n2173), .Z(n1301) );
  NANDN U1958 ( .A(n12632), .B(n2174), .Z(n1302) );
  AND U1959 ( .A(n1301), .B(n1302), .Z(n12658) );
  NANDN U1960 ( .A(n12775), .B(n2173), .Z(n1303) );
  NANDN U1961 ( .A(n12754), .B(n2174), .Z(n1304) );
  AND U1962 ( .A(n1303), .B(n1304), .Z(n12781) );
  NANDN U1963 ( .A(n12922), .B(n2173), .Z(n1305) );
  NANDN U1964 ( .A(n12901), .B(n2174), .Z(n1306) );
  AND U1965 ( .A(n1305), .B(n1306), .Z(n12928) );
  NANDN U1966 ( .A(n13069), .B(n2173), .Z(n1307) );
  NANDN U1967 ( .A(n13048), .B(n2174), .Z(n1308) );
  AND U1968 ( .A(n1307), .B(n1308), .Z(n13075) );
  NANDN U1969 ( .A(n13216), .B(n2173), .Z(n1309) );
  NANDN U1970 ( .A(n13195), .B(n2174), .Z(n1310) );
  AND U1971 ( .A(n1309), .B(n1310), .Z(n13222) );
  NANDN U1972 ( .A(n13363), .B(n2173), .Z(n1311) );
  NANDN U1973 ( .A(n13342), .B(n2174), .Z(n1312) );
  AND U1974 ( .A(n1311), .B(n1312), .Z(n13369) );
  NANDN U1975 ( .A(n13510), .B(n2173), .Z(n1313) );
  NANDN U1976 ( .A(n13489), .B(n2174), .Z(n1314) );
  AND U1977 ( .A(n1313), .B(n1314), .Z(n13516) );
  NANDN U1978 ( .A(n13657), .B(n2173), .Z(n1315) );
  NANDN U1979 ( .A(n13636), .B(n2174), .Z(n1316) );
  AND U1980 ( .A(n1315), .B(n1316), .Z(n13663) );
  NANDN U1981 ( .A(n13823), .B(n2173), .Z(n1317) );
  NANDN U1982 ( .A(n13804), .B(n2174), .Z(n1318) );
  AND U1983 ( .A(n1317), .B(n1318), .Z(n13830) );
  NANDN U1984 ( .A(n13947), .B(n2173), .Z(n1319) );
  NANDN U1985 ( .A(n13926), .B(n2174), .Z(n1320) );
  AND U1986 ( .A(n1319), .B(n1320), .Z(n13953) );
  NANDN U1987 ( .A(n14094), .B(n2173), .Z(n1321) );
  NANDN U1988 ( .A(n14073), .B(n2174), .Z(n1322) );
  AND U1989 ( .A(n1321), .B(n1322), .Z(n14100) );
  NANDN U1990 ( .A(n14241), .B(n2173), .Z(n1323) );
  NANDN U1991 ( .A(n14220), .B(n2174), .Z(n1324) );
  AND U1992 ( .A(n1323), .B(n1324), .Z(n14247) );
  NANDN U1993 ( .A(n14388), .B(n2173), .Z(n1325) );
  NANDN U1994 ( .A(n14367), .B(n2174), .Z(n1326) );
  AND U1995 ( .A(n1325), .B(n1326), .Z(n14394) );
  NANDN U1996 ( .A(n14535), .B(n2173), .Z(n1327) );
  NANDN U1997 ( .A(n14514), .B(n2174), .Z(n1328) );
  AND U1998 ( .A(n1327), .B(n1328), .Z(n14541) );
  NANDN U1999 ( .A(n14682), .B(n2173), .Z(n1329) );
  NANDN U2000 ( .A(n14661), .B(n2174), .Z(n1330) );
  AND U2001 ( .A(n1329), .B(n1330), .Z(n14688) );
  NANDN U2002 ( .A(n14825), .B(n2173), .Z(n1331) );
  NANDN U2003 ( .A(n14804), .B(n2174), .Z(n1332) );
  AND U2004 ( .A(n1331), .B(n1332), .Z(n14831) );
  NANDN U2005 ( .A(n14972), .B(n2173), .Z(n1333) );
  NANDN U2006 ( .A(n14951), .B(n2174), .Z(n1334) );
  AND U2007 ( .A(n1333), .B(n1334), .Z(n14978) );
  NANDN U2008 ( .A(n15119), .B(n2173), .Z(n1335) );
  NANDN U2009 ( .A(n15098), .B(n2174), .Z(n1336) );
  AND U2010 ( .A(n1335), .B(n1336), .Z(n15125) );
  NANDN U2011 ( .A(n15266), .B(n2173), .Z(n1337) );
  NANDN U2012 ( .A(n15245), .B(n2174), .Z(n1338) );
  AND U2013 ( .A(n1337), .B(n1338), .Z(n15272) );
  NANDN U2014 ( .A(n15413), .B(n2173), .Z(n1339) );
  NANDN U2015 ( .A(n15392), .B(n2174), .Z(n1340) );
  AND U2016 ( .A(n1339), .B(n1340), .Z(n15419) );
  NANDN U2017 ( .A(n15560), .B(n2173), .Z(n1341) );
  NANDN U2018 ( .A(n15539), .B(n2174), .Z(n1342) );
  AND U2019 ( .A(n1341), .B(n1342), .Z(n15566) );
  NANDN U2020 ( .A(n15703), .B(n2173), .Z(n1343) );
  NANDN U2021 ( .A(n15682), .B(n2174), .Z(n1344) );
  AND U2022 ( .A(n1343), .B(n1344), .Z(n15709) );
  NANDN U2023 ( .A(n15850), .B(n2173), .Z(n1345) );
  NANDN U2024 ( .A(n15829), .B(n2174), .Z(n1346) );
  AND U2025 ( .A(n1345), .B(n1346), .Z(n15856) );
  NANDN U2026 ( .A(n15997), .B(n2173), .Z(n1347) );
  NANDN U2027 ( .A(n15976), .B(n2174), .Z(n1348) );
  AND U2028 ( .A(n1347), .B(n1348), .Z(n16003) );
  NANDN U2029 ( .A(n16144), .B(n2173), .Z(n1349) );
  NANDN U2030 ( .A(n16123), .B(n2174), .Z(n1350) );
  AND U2031 ( .A(n1349), .B(n1350), .Z(n16150) );
  NANDN U2032 ( .A(n16291), .B(n2173), .Z(n1351) );
  NANDN U2033 ( .A(n16270), .B(n2174), .Z(n1352) );
  AND U2034 ( .A(n1351), .B(n1352), .Z(n16297) );
  NANDN U2035 ( .A(n16438), .B(n2173), .Z(n1353) );
  NANDN U2036 ( .A(n16417), .B(n2174), .Z(n1354) );
  AND U2037 ( .A(n1353), .B(n1354), .Z(n16444) );
  NANDN U2038 ( .A(n16585), .B(n2173), .Z(n1355) );
  NANDN U2039 ( .A(n16564), .B(n2174), .Z(n1356) );
  AND U2040 ( .A(n1355), .B(n1356), .Z(n16591) );
  NANDN U2041 ( .A(n16732), .B(n2173), .Z(n1357) );
  NANDN U2042 ( .A(n16711), .B(n2174), .Z(n1358) );
  AND U2043 ( .A(n1357), .B(n1358), .Z(n16738) );
  NANDN U2044 ( .A(n16879), .B(n2173), .Z(n1359) );
  NANDN U2045 ( .A(n16858), .B(n2174), .Z(n1360) );
  AND U2046 ( .A(n1359), .B(n1360), .Z(n16885) );
  NANDN U2047 ( .A(n17026), .B(n2173), .Z(n1361) );
  NANDN U2048 ( .A(n17005), .B(n2174), .Z(n1362) );
  AND U2049 ( .A(n1361), .B(n1362), .Z(n17032) );
  NANDN U2050 ( .A(n17173), .B(n2173), .Z(n1363) );
  NANDN U2051 ( .A(n17152), .B(n2174), .Z(n1364) );
  AND U2052 ( .A(n1363), .B(n1364), .Z(n17179) );
  NANDN U2053 ( .A(n17320), .B(n2173), .Z(n1365) );
  NANDN U2054 ( .A(n17299), .B(n2174), .Z(n1366) );
  AND U2055 ( .A(n1365), .B(n1366), .Z(n17326) );
  NANDN U2056 ( .A(n17467), .B(n2173), .Z(n1367) );
  NANDN U2057 ( .A(n17446), .B(n2174), .Z(n1368) );
  AND U2058 ( .A(n1367), .B(n1368), .Z(n17473) );
  NANDN U2059 ( .A(n17614), .B(n2173), .Z(n1369) );
  NANDN U2060 ( .A(n17593), .B(n2174), .Z(n1370) );
  AND U2061 ( .A(n1369), .B(n1370), .Z(n17620) );
  NANDN U2062 ( .A(n17776), .B(n2173), .Z(n1371) );
  NANDN U2063 ( .A(n17757), .B(n2174), .Z(n1372) );
  AND U2064 ( .A(n1371), .B(n1372), .Z(n17783) );
  NANDN U2065 ( .A(n17900), .B(n2173), .Z(n1373) );
  NANDN U2066 ( .A(n17879), .B(n2174), .Z(n1374) );
  AND U2067 ( .A(n1373), .B(n1374), .Z(n17906) );
  NANDN U2068 ( .A(n18047), .B(n2173), .Z(n1375) );
  NANDN U2069 ( .A(n18026), .B(n2174), .Z(n1376) );
  AND U2070 ( .A(n1375), .B(n1376), .Z(n18053) );
  NANDN U2071 ( .A(n18190), .B(n2173), .Z(n1377) );
  NANDN U2072 ( .A(n18169), .B(n2174), .Z(n1378) );
  AND U2073 ( .A(n1377), .B(n1378), .Z(n18196) );
  NANDN U2074 ( .A(n18337), .B(n2173), .Z(n1379) );
  NANDN U2075 ( .A(n18316), .B(n2174), .Z(n1380) );
  AND U2076 ( .A(n1379), .B(n1380), .Z(n18343) );
  NANDN U2077 ( .A(n18484), .B(n2173), .Z(n1381) );
  NANDN U2078 ( .A(n18463), .B(n2174), .Z(n1382) );
  AND U2079 ( .A(n1381), .B(n1382), .Z(n18490) );
  NANDN U2080 ( .A(n18631), .B(n2173), .Z(n1383) );
  NANDN U2081 ( .A(n18610), .B(n2174), .Z(n1384) );
  AND U2082 ( .A(n1383), .B(n1384), .Z(n18637) );
  NANDN U2083 ( .A(n18778), .B(n2173), .Z(n1385) );
  NANDN U2084 ( .A(n18757), .B(n2174), .Z(n1386) );
  AND U2085 ( .A(n1385), .B(n1386), .Z(n18784) );
  NANDN U2086 ( .A(n18925), .B(n2173), .Z(n1387) );
  NANDN U2087 ( .A(n18904), .B(n2174), .Z(n1388) );
  AND U2088 ( .A(n1387), .B(n1388), .Z(n18931) );
  NANDN U2089 ( .A(n19072), .B(n2173), .Z(n1389) );
  NANDN U2090 ( .A(n19051), .B(n2174), .Z(n1390) );
  AND U2091 ( .A(n1389), .B(n1390), .Z(n19078) );
  NANDN U2092 ( .A(n19219), .B(n2173), .Z(n1391) );
  NANDN U2093 ( .A(n19198), .B(n2174), .Z(n1392) );
  AND U2094 ( .A(n1391), .B(n1392), .Z(n19225) );
  NANDN U2095 ( .A(n19366), .B(n2173), .Z(n1393) );
  NANDN U2096 ( .A(n19345), .B(n2174), .Z(n1394) );
  AND U2097 ( .A(n1393), .B(n1394), .Z(n19372) );
  NANDN U2098 ( .A(n19513), .B(n2173), .Z(n1395) );
  NANDN U2099 ( .A(n19492), .B(n2174), .Z(n1396) );
  AND U2100 ( .A(n1395), .B(n1396), .Z(n19519) );
  NANDN U2101 ( .A(n19681), .B(n2173), .Z(n1397) );
  NANDN U2102 ( .A(n19660), .B(n2174), .Z(n1398) );
  AND U2103 ( .A(n1397), .B(n1398), .Z(n19687) );
  NANDN U2104 ( .A(n19803), .B(n2173), .Z(n1399) );
  NANDN U2105 ( .A(n19782), .B(n2174), .Z(n1400) );
  AND U2106 ( .A(n1399), .B(n1400), .Z(n19809) );
  NANDN U2107 ( .A(n19950), .B(n2173), .Z(n1401) );
  NANDN U2108 ( .A(n19929), .B(n2174), .Z(n1402) );
  AND U2109 ( .A(n1401), .B(n1402), .Z(n19956) );
  NANDN U2110 ( .A(n20118), .B(n2173), .Z(n1403) );
  NANDN U2111 ( .A(n20097), .B(n2174), .Z(n1404) );
  AND U2112 ( .A(n1403), .B(n1404), .Z(n20124) );
  NANDN U2113 ( .A(n20240), .B(n2173), .Z(n1405) );
  NANDN U2114 ( .A(n20219), .B(n2174), .Z(n1406) );
  AND U2115 ( .A(n1405), .B(n1406), .Z(n20246) );
  NANDN U2116 ( .A(n20387), .B(n2173), .Z(n1407) );
  NANDN U2117 ( .A(n20366), .B(n2174), .Z(n1408) );
  AND U2118 ( .A(n1407), .B(n1408), .Z(n20393) );
  NANDN U2119 ( .A(n20534), .B(n2173), .Z(n1409) );
  NANDN U2120 ( .A(n20513), .B(n2174), .Z(n1410) );
  AND U2121 ( .A(n1409), .B(n1410), .Z(n20540) );
  NANDN U2122 ( .A(n20681), .B(n2173), .Z(n1411) );
  NANDN U2123 ( .A(n20660), .B(n2174), .Z(n1412) );
  AND U2124 ( .A(n1411), .B(n1412), .Z(n20687) );
  NANDN U2125 ( .A(n20828), .B(n2173), .Z(n1413) );
  NANDN U2126 ( .A(n20807), .B(n2174), .Z(n1414) );
  AND U2127 ( .A(n1413), .B(n1414), .Z(n20834) );
  NANDN U2128 ( .A(n20975), .B(n2173), .Z(n1415) );
  NANDN U2129 ( .A(n20954), .B(n2174), .Z(n1416) );
  AND U2130 ( .A(n1415), .B(n1416), .Z(n20981) );
  NANDN U2131 ( .A(n21118), .B(n2173), .Z(n1417) );
  NANDN U2132 ( .A(n21097), .B(n2174), .Z(n1418) );
  AND U2133 ( .A(n1417), .B(n1418), .Z(n21124) );
  NANDN U2134 ( .A(n21284), .B(n2173), .Z(n1419) );
  NANDN U2135 ( .A(n21265), .B(n2174), .Z(n1420) );
  AND U2136 ( .A(n1419), .B(n1420), .Z(n21291) );
  NANDN U2137 ( .A(n21408), .B(n2173), .Z(n1421) );
  NANDN U2138 ( .A(n21387), .B(n2174), .Z(n1422) );
  AND U2139 ( .A(n1421), .B(n1422), .Z(n21414) );
  NANDN U2140 ( .A(n21555), .B(n2173), .Z(n1423) );
  NANDN U2141 ( .A(n21534), .B(n2174), .Z(n1424) );
  AND U2142 ( .A(n1423), .B(n1424), .Z(n21561) );
  NANDN U2143 ( .A(n21702), .B(n2173), .Z(n1425) );
  NANDN U2144 ( .A(n21681), .B(n2174), .Z(n1426) );
  AND U2145 ( .A(n1425), .B(n1426), .Z(n21708) );
  NANDN U2146 ( .A(n21849), .B(n2173), .Z(n1427) );
  NANDN U2147 ( .A(n21828), .B(n2174), .Z(n1428) );
  AND U2148 ( .A(n1427), .B(n1428), .Z(n21855) );
  NANDN U2149 ( .A(n21996), .B(n2173), .Z(n1429) );
  NANDN U2150 ( .A(n21975), .B(n2174), .Z(n1430) );
  AND U2151 ( .A(n1429), .B(n1430), .Z(n22002) );
  NANDN U2152 ( .A(n22143), .B(n2173), .Z(n1431) );
  NANDN U2153 ( .A(n22122), .B(n2174), .Z(n1432) );
  AND U2154 ( .A(n1431), .B(n1432), .Z(n22149) );
  NANDN U2155 ( .A(n22311), .B(n2173), .Z(n1433) );
  NANDN U2156 ( .A(n22290), .B(n2174), .Z(n1434) );
  AND U2157 ( .A(n1433), .B(n1434), .Z(n22317) );
  NANDN U2158 ( .A(n22433), .B(n2173), .Z(n1435) );
  NANDN U2159 ( .A(n22412), .B(n2174), .Z(n1436) );
  AND U2160 ( .A(n1435), .B(n1436), .Z(n22439) );
  NANDN U2161 ( .A(n22580), .B(n2173), .Z(n1437) );
  NANDN U2162 ( .A(n22559), .B(n2174), .Z(n1438) );
  AND U2163 ( .A(n1437), .B(n1438), .Z(n22586) );
  NANDN U2164 ( .A(n22727), .B(n2173), .Z(n1439) );
  NANDN U2165 ( .A(n22706), .B(n2174), .Z(n1440) );
  AND U2166 ( .A(n1439), .B(n1440), .Z(n22733) );
  NANDN U2167 ( .A(n22874), .B(n2173), .Z(n1441) );
  NANDN U2168 ( .A(n22853), .B(n2174), .Z(n1442) );
  AND U2169 ( .A(n1441), .B(n1442), .Z(n22880) );
  NANDN U2170 ( .A(n23021), .B(n2173), .Z(n1443) );
  NANDN U2171 ( .A(n23000), .B(n2174), .Z(n1444) );
  AND U2172 ( .A(n1443), .B(n1444), .Z(n23027) );
  NANDN U2173 ( .A(n23168), .B(n2173), .Z(n1445) );
  NANDN U2174 ( .A(n23147), .B(n2174), .Z(n1446) );
  AND U2175 ( .A(n1445), .B(n1446), .Z(n23174) );
  NANDN U2176 ( .A(n23315), .B(n2173), .Z(n1447) );
  NANDN U2177 ( .A(n23294), .B(n2174), .Z(n1448) );
  AND U2178 ( .A(n1447), .B(n1448), .Z(n23321) );
  NANDN U2179 ( .A(n23462), .B(n2173), .Z(n1449) );
  NANDN U2180 ( .A(n23441), .B(n2174), .Z(n1450) );
  AND U2181 ( .A(n1449), .B(n1450), .Z(n23468) );
  NANDN U2182 ( .A(n23604), .B(n2173), .Z(n1451) );
  NANDN U2183 ( .A(n23586), .B(n2174), .Z(n1452) );
  AND U2184 ( .A(n1451), .B(n1452), .Z(n23611) );
  NANDN U2185 ( .A(n11752), .B(n11753), .Z(n1453) );
  NANDN U2186 ( .A(n11755), .B(n11754), .Z(n1454) );
  AND U2187 ( .A(n1453), .B(n1454), .Z(n11771) );
  NANDN U2188 ( .A(n17734), .B(n17735), .Z(n1455) );
  NANDN U2189 ( .A(n17737), .B(n17736), .Z(n1456) );
  AND U2190 ( .A(n1455), .B(n1456), .Z(n17753) );
  NANDN U2191 ( .A(n23582), .B(n23583), .Z(n1457) );
  NANDN U2192 ( .A(n23585), .B(n23584), .Z(n1458) );
  AND U2193 ( .A(n1457), .B(n1458), .Z(n23603) );
  NANDN U2194 ( .A(n2415), .B(n2173), .Z(n1459) );
  NANDN U2195 ( .A(n2394), .B(n2174), .Z(n1460) );
  AND U2196 ( .A(n1459), .B(n1460), .Z(n2421) );
  NANDN U2197 ( .A(n2562), .B(n2173), .Z(n1461) );
  NANDN U2198 ( .A(n2541), .B(n2174), .Z(n1462) );
  AND U2199 ( .A(n1461), .B(n1462), .Z(n2568) );
  NANDN U2200 ( .A(n2709), .B(n2173), .Z(n1463) );
  NANDN U2201 ( .A(n2688), .B(n2174), .Z(n1464) );
  AND U2202 ( .A(n1463), .B(n1464), .Z(n2715) );
  NANDN U2203 ( .A(n2856), .B(n2173), .Z(n1465) );
  NANDN U2204 ( .A(n2835), .B(n2174), .Z(n1466) );
  AND U2205 ( .A(n1465), .B(n1466), .Z(n2862) );
  NANDN U2206 ( .A(n3003), .B(n2173), .Z(n1467) );
  NANDN U2207 ( .A(n2982), .B(n2174), .Z(n1468) );
  AND U2208 ( .A(n1467), .B(n1468), .Z(n3009) );
  NANDN U2209 ( .A(n3150), .B(n2173), .Z(n1469) );
  NANDN U2210 ( .A(n3129), .B(n2174), .Z(n1470) );
  AND U2211 ( .A(n1469), .B(n1470), .Z(n3156) );
  NANDN U2212 ( .A(n3297), .B(n2173), .Z(n1471) );
  NANDN U2213 ( .A(n3276), .B(n2174), .Z(n1472) );
  AND U2214 ( .A(n1471), .B(n1472), .Z(n3303) );
  NANDN U2215 ( .A(n3444), .B(n2173), .Z(n1473) );
  NANDN U2216 ( .A(n3423), .B(n2174), .Z(n1474) );
  AND U2217 ( .A(n1473), .B(n1474), .Z(n3450) );
  NANDN U2218 ( .A(n3591), .B(n2173), .Z(n1475) );
  NANDN U2219 ( .A(n3570), .B(n2174), .Z(n1476) );
  AND U2220 ( .A(n1475), .B(n1476), .Z(n3597) );
  NANDN U2221 ( .A(n3738), .B(n2173), .Z(n1477) );
  NANDN U2222 ( .A(n3717), .B(n2174), .Z(n1478) );
  AND U2223 ( .A(n1477), .B(n1478), .Z(n3744) );
  NANDN U2224 ( .A(n3885), .B(n2173), .Z(n1479) );
  NANDN U2225 ( .A(n3864), .B(n2174), .Z(n1480) );
  AND U2226 ( .A(n1479), .B(n1480), .Z(n3891) );
  NANDN U2227 ( .A(n4032), .B(n2173), .Z(n1481) );
  NANDN U2228 ( .A(n4011), .B(n2174), .Z(n1482) );
  AND U2229 ( .A(n1481), .B(n1482), .Z(n4038) );
  NANDN U2230 ( .A(n4179), .B(n2173), .Z(n1483) );
  NANDN U2231 ( .A(n4158), .B(n2174), .Z(n1484) );
  AND U2232 ( .A(n1483), .B(n1484), .Z(n4185) );
  NANDN U2233 ( .A(n4326), .B(n2173), .Z(n1485) );
  NANDN U2234 ( .A(n4305), .B(n2174), .Z(n1486) );
  AND U2235 ( .A(n1485), .B(n1486), .Z(n4332) );
  NANDN U2236 ( .A(n4469), .B(n2173), .Z(n1487) );
  NANDN U2237 ( .A(n4448), .B(n2174), .Z(n1488) );
  AND U2238 ( .A(n1487), .B(n1488), .Z(n4475) );
  NANDN U2239 ( .A(n4616), .B(n2173), .Z(n1489) );
  NANDN U2240 ( .A(n4595), .B(n2174), .Z(n1490) );
  AND U2241 ( .A(n1489), .B(n1490), .Z(n4622) );
  NANDN U2242 ( .A(n4763), .B(n2173), .Z(n1491) );
  NANDN U2243 ( .A(n4742), .B(n2174), .Z(n1492) );
  AND U2244 ( .A(n1491), .B(n1492), .Z(n4769) );
  NANDN U2245 ( .A(n4910), .B(n2173), .Z(n1493) );
  NANDN U2246 ( .A(n4889), .B(n2174), .Z(n1494) );
  AND U2247 ( .A(n1493), .B(n1494), .Z(n4916) );
  NANDN U2248 ( .A(n5057), .B(n2173), .Z(n1495) );
  NANDN U2249 ( .A(n5036), .B(n2174), .Z(n1496) );
  AND U2250 ( .A(n1495), .B(n1496), .Z(n5063) );
  NANDN U2251 ( .A(n5204), .B(n2173), .Z(n1497) );
  NANDN U2252 ( .A(n5183), .B(n2174), .Z(n1498) );
  AND U2253 ( .A(n1497), .B(n1498), .Z(n5210) );
  NANDN U2254 ( .A(n5351), .B(n2173), .Z(n1499) );
  NANDN U2255 ( .A(n5330), .B(n2174), .Z(n1500) );
  AND U2256 ( .A(n1499), .B(n1500), .Z(n5357) );
  NANDN U2257 ( .A(n5498), .B(n2173), .Z(n1501) );
  NANDN U2258 ( .A(n5477), .B(n2174), .Z(n1502) );
  AND U2259 ( .A(n1501), .B(n1502), .Z(n5504) );
  NANDN U2260 ( .A(n5645), .B(n2173), .Z(n1503) );
  NANDN U2261 ( .A(n5624), .B(n2174), .Z(n1504) );
  AND U2262 ( .A(n1503), .B(n1504), .Z(n5651) );
  NANDN U2263 ( .A(n5792), .B(n2173), .Z(n1505) );
  NANDN U2264 ( .A(n5771), .B(n2174), .Z(n1506) );
  AND U2265 ( .A(n1505), .B(n1506), .Z(n5798) );
  NANDN U2266 ( .A(n5939), .B(n2173), .Z(n1507) );
  NANDN U2267 ( .A(n5918), .B(n2174), .Z(n1508) );
  AND U2268 ( .A(n1507), .B(n1508), .Z(n5945) );
  NANDN U2269 ( .A(n6086), .B(n2173), .Z(n1509) );
  NANDN U2270 ( .A(n6065), .B(n2174), .Z(n1510) );
  AND U2271 ( .A(n1509), .B(n1510), .Z(n6092) );
  NANDN U2272 ( .A(n6233), .B(n2173), .Z(n1511) );
  NANDN U2273 ( .A(n6212), .B(n2174), .Z(n1512) );
  AND U2274 ( .A(n1511), .B(n1512), .Z(n6239) );
  NANDN U2275 ( .A(n6380), .B(n2173), .Z(n1513) );
  NANDN U2276 ( .A(n6359), .B(n2174), .Z(n1514) );
  AND U2277 ( .A(n1513), .B(n1514), .Z(n6386) );
  NANDN U2278 ( .A(n6523), .B(n2173), .Z(n1515) );
  NANDN U2279 ( .A(n6502), .B(n2174), .Z(n1516) );
  AND U2280 ( .A(n1515), .B(n1516), .Z(n6529) );
  NANDN U2281 ( .A(n6670), .B(n2173), .Z(n1517) );
  NANDN U2282 ( .A(n6649), .B(n2174), .Z(n1518) );
  AND U2283 ( .A(n1517), .B(n1518), .Z(n6676) );
  NANDN U2284 ( .A(n6796), .B(n2173), .Z(n1519) );
  NANDN U2285 ( .A(n6775), .B(n2174), .Z(n1520) );
  AND U2286 ( .A(n1519), .B(n1520), .Z(n6802) );
  NANDN U2287 ( .A(n6956), .B(n2173), .Z(n1521) );
  NANDN U2288 ( .A(n6937), .B(n2174), .Z(n1522) );
  AND U2289 ( .A(n1521), .B(n1522), .Z(n6962) );
  NANDN U2290 ( .A(n7061), .B(n2173), .Z(n1523) );
  NANDN U2291 ( .A(n7040), .B(n2174), .Z(n1524) );
  AND U2292 ( .A(n1523), .B(n1524), .Z(n7067) );
  NANDN U2293 ( .A(n7246), .B(n2173), .Z(n1525) );
  NANDN U2294 ( .A(n7225), .B(n2174), .Z(n1526) );
  AND U2295 ( .A(n1525), .B(n1526), .Z(n7252) );
  NANDN U2296 ( .A(n7393), .B(n2173), .Z(n1527) );
  NANDN U2297 ( .A(n7372), .B(n2174), .Z(n1528) );
  AND U2298 ( .A(n1527), .B(n1528), .Z(n7399) );
  NANDN U2299 ( .A(n7498), .B(n2173), .Z(n1529) );
  NANDN U2300 ( .A(n7477), .B(n2174), .Z(n1530) );
  AND U2301 ( .A(n1529), .B(n1530), .Z(n7504) );
  NANDN U2302 ( .A(n7683), .B(n2173), .Z(n1531) );
  NANDN U2303 ( .A(n7662), .B(n2174), .Z(n1532) );
  AND U2304 ( .A(n1531), .B(n1532), .Z(n7689) );
  NANDN U2305 ( .A(n7826), .B(n2173), .Z(n1533) );
  NANDN U2306 ( .A(n7807), .B(n2174), .Z(n1534) );
  AND U2307 ( .A(n1533), .B(n1534), .Z(n7832) );
  NANDN U2308 ( .A(n7969), .B(n2173), .Z(n1535) );
  NANDN U2309 ( .A(n7948), .B(n2174), .Z(n1536) );
  AND U2310 ( .A(n1535), .B(n1536), .Z(n7975) );
  NANDN U2311 ( .A(n8116), .B(n2173), .Z(n1537) );
  NANDN U2312 ( .A(n8095), .B(n2174), .Z(n1538) );
  AND U2313 ( .A(n1537), .B(n1538), .Z(n8122) );
  NANDN U2314 ( .A(n8259), .B(n2173), .Z(n1539) );
  NANDN U2315 ( .A(n8238), .B(n2174), .Z(n1540) );
  AND U2316 ( .A(n1539), .B(n1540), .Z(n8265) );
  NANDN U2317 ( .A(n8406), .B(n2173), .Z(n1541) );
  NANDN U2318 ( .A(n8385), .B(n2174), .Z(n1542) );
  AND U2319 ( .A(n1541), .B(n1542), .Z(n8412) );
  NANDN U2320 ( .A(n8553), .B(n2173), .Z(n1543) );
  NANDN U2321 ( .A(n8532), .B(n2174), .Z(n1544) );
  AND U2322 ( .A(n1543), .B(n1544), .Z(n8559) );
  NANDN U2323 ( .A(n8700), .B(n2173), .Z(n1545) );
  NANDN U2324 ( .A(n8679), .B(n2174), .Z(n1546) );
  AND U2325 ( .A(n1545), .B(n1546), .Z(n8706) );
  NANDN U2326 ( .A(n8847), .B(n2173), .Z(n1547) );
  NANDN U2327 ( .A(n8826), .B(n2174), .Z(n1548) );
  AND U2328 ( .A(n1547), .B(n1548), .Z(n8853) );
  NANDN U2329 ( .A(n8994), .B(n2173), .Z(n1549) );
  NANDN U2330 ( .A(n8973), .B(n2174), .Z(n1550) );
  AND U2331 ( .A(n1549), .B(n1550), .Z(n9000) );
  NANDN U2332 ( .A(n9137), .B(n2173), .Z(n1551) );
  NANDN U2333 ( .A(n9116), .B(n2174), .Z(n1552) );
  AND U2334 ( .A(n1551), .B(n1552), .Z(n9143) );
  NANDN U2335 ( .A(n9280), .B(n2173), .Z(n1553) );
  NANDN U2336 ( .A(n9259), .B(n2174), .Z(n1554) );
  AND U2337 ( .A(n1553), .B(n1554), .Z(n9286) );
  NANDN U2338 ( .A(n9427), .B(n2173), .Z(n1555) );
  NANDN U2339 ( .A(n9406), .B(n2174), .Z(n1556) );
  AND U2340 ( .A(n1555), .B(n1556), .Z(n9433) );
  NANDN U2341 ( .A(n9574), .B(n2173), .Z(n1557) );
  NANDN U2342 ( .A(n9553), .B(n2174), .Z(n1558) );
  AND U2343 ( .A(n1557), .B(n1558), .Z(n9580) );
  NANDN U2344 ( .A(n9721), .B(n2173), .Z(n1559) );
  NANDN U2345 ( .A(n9700), .B(n2174), .Z(n1560) );
  AND U2346 ( .A(n1559), .B(n1560), .Z(n9727) );
  NANDN U2347 ( .A(n9868), .B(n2173), .Z(n1561) );
  NANDN U2348 ( .A(n9847), .B(n2174), .Z(n1562) );
  AND U2349 ( .A(n1561), .B(n1562), .Z(n9874) );
  NANDN U2350 ( .A(n10015), .B(n2173), .Z(n1563) );
  NANDN U2351 ( .A(n9994), .B(n2174), .Z(n1564) );
  AND U2352 ( .A(n1563), .B(n1564), .Z(n10021) );
  NANDN U2353 ( .A(n10162), .B(n2173), .Z(n1565) );
  NANDN U2354 ( .A(n10141), .B(n2174), .Z(n1566) );
  AND U2355 ( .A(n1565), .B(n1566), .Z(n10168) );
  NANDN U2356 ( .A(n10309), .B(n2173), .Z(n1567) );
  NANDN U2357 ( .A(n10288), .B(n2174), .Z(n1568) );
  AND U2358 ( .A(n1567), .B(n1568), .Z(n10315) );
  NANDN U2359 ( .A(n10456), .B(n2173), .Z(n1569) );
  NANDN U2360 ( .A(n10435), .B(n2174), .Z(n1570) );
  AND U2361 ( .A(n1569), .B(n1570), .Z(n10462) );
  NANDN U2362 ( .A(n10603), .B(n2173), .Z(n1571) );
  NANDN U2363 ( .A(n10582), .B(n2174), .Z(n1572) );
  AND U2364 ( .A(n1571), .B(n1572), .Z(n10609) );
  NANDN U2365 ( .A(n10750), .B(n2173), .Z(n1573) );
  NANDN U2366 ( .A(n10729), .B(n2174), .Z(n1574) );
  AND U2367 ( .A(n1573), .B(n1574), .Z(n10756) );
  NANDN U2368 ( .A(n10897), .B(n2173), .Z(n1575) );
  NANDN U2369 ( .A(n10876), .B(n2174), .Z(n1576) );
  AND U2370 ( .A(n1575), .B(n1576), .Z(n10903) );
  NANDN U2371 ( .A(n11044), .B(n2173), .Z(n1577) );
  NANDN U2372 ( .A(n11023), .B(n2174), .Z(n1578) );
  AND U2373 ( .A(n1577), .B(n1578), .Z(n11050) );
  NANDN U2374 ( .A(n11191), .B(n2173), .Z(n1579) );
  NANDN U2375 ( .A(n11170), .B(n2174), .Z(n1580) );
  AND U2376 ( .A(n1579), .B(n1580), .Z(n11197) );
  NANDN U2377 ( .A(n11338), .B(n2173), .Z(n1581) );
  NANDN U2378 ( .A(n11317), .B(n2174), .Z(n1582) );
  AND U2379 ( .A(n1581), .B(n1582), .Z(n11344) );
  NANDN U2380 ( .A(n11485), .B(n2173), .Z(n1583) );
  NANDN U2381 ( .A(n11464), .B(n2174), .Z(n1584) );
  AND U2382 ( .A(n1583), .B(n1584), .Z(n11491) );
  NANDN U2383 ( .A(n11632), .B(n2173), .Z(n1585) );
  NANDN U2384 ( .A(n11611), .B(n2174), .Z(n1586) );
  AND U2385 ( .A(n1585), .B(n1586), .Z(n11638) );
  NANDN U2386 ( .A(n11756), .B(n2173), .Z(n1587) );
  NANDN U2387 ( .A(n11737), .B(n2174), .Z(n1588) );
  AND U2388 ( .A(n1587), .B(n1588), .Z(n11763) );
  NANDN U2389 ( .A(n11918), .B(n2173), .Z(n1589) );
  NANDN U2390 ( .A(n11897), .B(n2174), .Z(n1590) );
  AND U2391 ( .A(n1589), .B(n1590), .Z(n11924) );
  NANDN U2392 ( .A(n12065), .B(n2173), .Z(n1591) );
  NANDN U2393 ( .A(n12044), .B(n2174), .Z(n1592) );
  AND U2394 ( .A(n1591), .B(n1592), .Z(n12071) );
  NANDN U2395 ( .A(n12212), .B(n2173), .Z(n1593) );
  NANDN U2396 ( .A(n12191), .B(n2174), .Z(n1594) );
  AND U2397 ( .A(n1593), .B(n1594), .Z(n12218) );
  NANDN U2398 ( .A(n12359), .B(n2173), .Z(n1595) );
  NANDN U2399 ( .A(n12338), .B(n2174), .Z(n1596) );
  AND U2400 ( .A(n1595), .B(n1596), .Z(n12365) );
  NANDN U2401 ( .A(n12506), .B(n2173), .Z(n1597) );
  NANDN U2402 ( .A(n12485), .B(n2174), .Z(n1598) );
  AND U2403 ( .A(n1597), .B(n1598), .Z(n12512) );
  NANDN U2404 ( .A(n12611), .B(n2173), .Z(n1599) );
  NANDN U2405 ( .A(n12590), .B(n2174), .Z(n1600) );
  AND U2406 ( .A(n1599), .B(n1600), .Z(n12617) );
  NANDN U2407 ( .A(n12796), .B(n2173), .Z(n1601) );
  NANDN U2408 ( .A(n12775), .B(n2174), .Z(n1602) );
  AND U2409 ( .A(n1601), .B(n1602), .Z(n12802) );
  NANDN U2410 ( .A(n12943), .B(n2173), .Z(n1603) );
  NANDN U2411 ( .A(n12922), .B(n2174), .Z(n1604) );
  AND U2412 ( .A(n1603), .B(n1604), .Z(n12949) );
  NANDN U2413 ( .A(n13090), .B(n2173), .Z(n1605) );
  NANDN U2414 ( .A(n13069), .B(n2174), .Z(n1606) );
  AND U2415 ( .A(n1605), .B(n1606), .Z(n13096) );
  NANDN U2416 ( .A(n13237), .B(n2173), .Z(n1607) );
  NANDN U2417 ( .A(n13216), .B(n2174), .Z(n1608) );
  AND U2418 ( .A(n1607), .B(n1608), .Z(n13243) );
  NANDN U2419 ( .A(n13384), .B(n2173), .Z(n1609) );
  NANDN U2420 ( .A(n13363), .B(n2174), .Z(n1610) );
  AND U2421 ( .A(n1609), .B(n1610), .Z(n13390) );
  NANDN U2422 ( .A(n13531), .B(n2173), .Z(n1611) );
  NANDN U2423 ( .A(n13510), .B(n2174), .Z(n1612) );
  AND U2424 ( .A(n1611), .B(n1612), .Z(n13537) );
  NANDN U2425 ( .A(n13678), .B(n2173), .Z(n1613) );
  NANDN U2426 ( .A(n13657), .B(n2174), .Z(n1614) );
  AND U2427 ( .A(n1613), .B(n1614), .Z(n13684) );
  NANDN U2428 ( .A(n13783), .B(n2173), .Z(n1615) );
  NANDN U2429 ( .A(n13762), .B(n2174), .Z(n1616) );
  AND U2430 ( .A(n1615), .B(n1616), .Z(n13789) );
  NANDN U2431 ( .A(n13968), .B(n2173), .Z(n1617) );
  NANDN U2432 ( .A(n13947), .B(n2174), .Z(n1618) );
  AND U2433 ( .A(n1617), .B(n1618), .Z(n13974) );
  NANDN U2434 ( .A(n14115), .B(n2173), .Z(n1619) );
  NANDN U2435 ( .A(n14094), .B(n2174), .Z(n1620) );
  AND U2436 ( .A(n1619), .B(n1620), .Z(n14121) );
  NANDN U2437 ( .A(n14262), .B(n2173), .Z(n1621) );
  NANDN U2438 ( .A(n14241), .B(n2174), .Z(n1622) );
  AND U2439 ( .A(n1621), .B(n1622), .Z(n14268) );
  NANDN U2440 ( .A(n14409), .B(n2173), .Z(n1623) );
  NANDN U2441 ( .A(n14388), .B(n2174), .Z(n1624) );
  AND U2442 ( .A(n1623), .B(n1624), .Z(n14415) );
  NANDN U2443 ( .A(n14556), .B(n2173), .Z(n1625) );
  NANDN U2444 ( .A(n14535), .B(n2174), .Z(n1626) );
  AND U2445 ( .A(n1625), .B(n1626), .Z(n14562) );
  NANDN U2446 ( .A(n14703), .B(n2173), .Z(n1627) );
  NANDN U2447 ( .A(n14682), .B(n2174), .Z(n1628) );
  AND U2448 ( .A(n1627), .B(n1628), .Z(n14709) );
  NANDN U2449 ( .A(n14846), .B(n2173), .Z(n1629) );
  NANDN U2450 ( .A(n14825), .B(n2174), .Z(n1630) );
  AND U2451 ( .A(n1629), .B(n1630), .Z(n14852) );
  NANDN U2452 ( .A(n14993), .B(n2173), .Z(n1631) );
  NANDN U2453 ( .A(n14972), .B(n2174), .Z(n1632) );
  AND U2454 ( .A(n1631), .B(n1632), .Z(n14999) );
  NANDN U2455 ( .A(n15140), .B(n2173), .Z(n1633) );
  NANDN U2456 ( .A(n15119), .B(n2174), .Z(n1634) );
  AND U2457 ( .A(n1633), .B(n1634), .Z(n15146) );
  NANDN U2458 ( .A(n15287), .B(n2173), .Z(n1635) );
  NANDN U2459 ( .A(n15266), .B(n2174), .Z(n1636) );
  AND U2460 ( .A(n1635), .B(n1636), .Z(n15293) );
  NANDN U2461 ( .A(n15434), .B(n2173), .Z(n1637) );
  NANDN U2462 ( .A(n15413), .B(n2174), .Z(n1638) );
  AND U2463 ( .A(n1637), .B(n1638), .Z(n15440) );
  NANDN U2464 ( .A(n15581), .B(n2173), .Z(n1639) );
  NANDN U2465 ( .A(n15560), .B(n2174), .Z(n1640) );
  AND U2466 ( .A(n1639), .B(n1640), .Z(n15587) );
  NANDN U2467 ( .A(n15724), .B(n2173), .Z(n1641) );
  NANDN U2468 ( .A(n15703), .B(n2174), .Z(n1642) );
  AND U2469 ( .A(n1641), .B(n1642), .Z(n15730) );
  NANDN U2470 ( .A(n15871), .B(n2173), .Z(n1643) );
  NANDN U2471 ( .A(n15850), .B(n2174), .Z(n1644) );
  AND U2472 ( .A(n1643), .B(n1644), .Z(n15877) );
  NANDN U2473 ( .A(n16018), .B(n2173), .Z(n1645) );
  NANDN U2474 ( .A(n15997), .B(n2174), .Z(n1646) );
  AND U2475 ( .A(n1645), .B(n1646), .Z(n16024) );
  NANDN U2476 ( .A(n16165), .B(n2173), .Z(n1647) );
  NANDN U2477 ( .A(n16144), .B(n2174), .Z(n1648) );
  AND U2478 ( .A(n1647), .B(n1648), .Z(n16171) );
  NANDN U2479 ( .A(n16312), .B(n2173), .Z(n1649) );
  NANDN U2480 ( .A(n16291), .B(n2174), .Z(n1650) );
  AND U2481 ( .A(n1649), .B(n1650), .Z(n16318) );
  NANDN U2482 ( .A(n16459), .B(n2173), .Z(n1651) );
  NANDN U2483 ( .A(n16438), .B(n2174), .Z(n1652) );
  AND U2484 ( .A(n1651), .B(n1652), .Z(n16465) );
  NANDN U2485 ( .A(n16606), .B(n2173), .Z(n1653) );
  NANDN U2486 ( .A(n16585), .B(n2174), .Z(n1654) );
  AND U2487 ( .A(n1653), .B(n1654), .Z(n16612) );
  NANDN U2488 ( .A(n16753), .B(n2173), .Z(n1655) );
  NANDN U2489 ( .A(n16732), .B(n2174), .Z(n1656) );
  AND U2490 ( .A(n1655), .B(n1656), .Z(n16759) );
  NANDN U2491 ( .A(n16900), .B(n2173), .Z(n1657) );
  NANDN U2492 ( .A(n16879), .B(n2174), .Z(n1658) );
  AND U2493 ( .A(n1657), .B(n1658), .Z(n16906) );
  NANDN U2494 ( .A(n17047), .B(n2173), .Z(n1659) );
  NANDN U2495 ( .A(n17026), .B(n2174), .Z(n1660) );
  AND U2496 ( .A(n1659), .B(n1660), .Z(n17053) );
  NANDN U2497 ( .A(n17194), .B(n2173), .Z(n1661) );
  NANDN U2498 ( .A(n17173), .B(n2174), .Z(n1662) );
  AND U2499 ( .A(n1661), .B(n1662), .Z(n17200) );
  NANDN U2500 ( .A(n17341), .B(n2173), .Z(n1663) );
  NANDN U2501 ( .A(n17320), .B(n2174), .Z(n1664) );
  AND U2502 ( .A(n1663), .B(n1664), .Z(n17347) );
  NANDN U2503 ( .A(n17488), .B(n2173), .Z(n1665) );
  NANDN U2504 ( .A(n17467), .B(n2174), .Z(n1666) );
  AND U2505 ( .A(n1665), .B(n1666), .Z(n17494) );
  NANDN U2506 ( .A(n17635), .B(n2173), .Z(n1667) );
  NANDN U2507 ( .A(n17614), .B(n2174), .Z(n1668) );
  AND U2508 ( .A(n1667), .B(n1668), .Z(n17641) );
  NANDN U2509 ( .A(n17738), .B(n2173), .Z(n1669) );
  NANDN U2510 ( .A(n17719), .B(n2174), .Z(n1670) );
  AND U2511 ( .A(n1669), .B(n1670), .Z(n17745) );
  NANDN U2512 ( .A(n17921), .B(n2173), .Z(n1671) );
  NANDN U2513 ( .A(n17900), .B(n2174), .Z(n1672) );
  AND U2514 ( .A(n1671), .B(n1672), .Z(n17927) );
  NANDN U2515 ( .A(n18068), .B(n2173), .Z(n1673) );
  NANDN U2516 ( .A(n18047), .B(n2174), .Z(n1674) );
  AND U2517 ( .A(n1673), .B(n1674), .Z(n18074) );
  NANDN U2518 ( .A(n18211), .B(n2173), .Z(n1675) );
  NANDN U2519 ( .A(n18190), .B(n2174), .Z(n1676) );
  AND U2520 ( .A(n1675), .B(n1676), .Z(n18217) );
  NANDN U2521 ( .A(n18358), .B(n2173), .Z(n1677) );
  NANDN U2522 ( .A(n18337), .B(n2174), .Z(n1678) );
  AND U2523 ( .A(n1677), .B(n1678), .Z(n18364) );
  NANDN U2524 ( .A(n18505), .B(n2173), .Z(n1679) );
  NANDN U2525 ( .A(n18484), .B(n2174), .Z(n1680) );
  AND U2526 ( .A(n1679), .B(n1680), .Z(n18511) );
  NANDN U2527 ( .A(n18652), .B(n2173), .Z(n1681) );
  NANDN U2528 ( .A(n18631), .B(n2174), .Z(n1682) );
  AND U2529 ( .A(n1681), .B(n1682), .Z(n18658) );
  NANDN U2530 ( .A(n18799), .B(n2173), .Z(n1683) );
  NANDN U2531 ( .A(n18778), .B(n2174), .Z(n1684) );
  AND U2532 ( .A(n1683), .B(n1684), .Z(n18805) );
  NANDN U2533 ( .A(n18946), .B(n2173), .Z(n1685) );
  NANDN U2534 ( .A(n18925), .B(n2174), .Z(n1686) );
  AND U2535 ( .A(n1685), .B(n1686), .Z(n18952) );
  NANDN U2536 ( .A(n19093), .B(n2173), .Z(n1687) );
  NANDN U2537 ( .A(n19072), .B(n2174), .Z(n1688) );
  AND U2538 ( .A(n1687), .B(n1688), .Z(n19099) );
  NANDN U2539 ( .A(n19240), .B(n2173), .Z(n1689) );
  NANDN U2540 ( .A(n19219), .B(n2174), .Z(n1690) );
  AND U2541 ( .A(n1689), .B(n1690), .Z(n19246) );
  NANDN U2542 ( .A(n19387), .B(n2173), .Z(n1691) );
  NANDN U2543 ( .A(n19366), .B(n2174), .Z(n1692) );
  AND U2544 ( .A(n1691), .B(n1692), .Z(n19393) );
  NANDN U2545 ( .A(n19534), .B(n2173), .Z(n1693) );
  NANDN U2546 ( .A(n19513), .B(n2174), .Z(n1694) );
  AND U2547 ( .A(n1693), .B(n1694), .Z(n19540) );
  NANDN U2548 ( .A(n19660), .B(n2173), .Z(n1695) );
  NANDN U2549 ( .A(n19639), .B(n2174), .Z(n1696) );
  AND U2550 ( .A(n1695), .B(n1696), .Z(n19666) );
  NANDN U2551 ( .A(n19824), .B(n2173), .Z(n1697) );
  NANDN U2552 ( .A(n19803), .B(n2174), .Z(n1698) );
  AND U2553 ( .A(n1697), .B(n1698), .Z(n19830) );
  NANDN U2554 ( .A(n19971), .B(n2173), .Z(n1699) );
  NANDN U2555 ( .A(n19950), .B(n2174), .Z(n1700) );
  AND U2556 ( .A(n1699), .B(n1700), .Z(n19977) );
  NANDN U2557 ( .A(n20097), .B(n2173), .Z(n1701) );
  NANDN U2558 ( .A(n20076), .B(n2174), .Z(n1702) );
  AND U2559 ( .A(n1701), .B(n1702), .Z(n20103) );
  NANDN U2560 ( .A(n20261), .B(n2173), .Z(n1703) );
  NANDN U2561 ( .A(n20240), .B(n2174), .Z(n1704) );
  AND U2562 ( .A(n1703), .B(n1704), .Z(n20267) );
  NANDN U2563 ( .A(n20408), .B(n2173), .Z(n1705) );
  NANDN U2564 ( .A(n20387), .B(n2174), .Z(n1706) );
  AND U2565 ( .A(n1705), .B(n1706), .Z(n20414) );
  NANDN U2566 ( .A(n20555), .B(n2173), .Z(n1707) );
  NANDN U2567 ( .A(n20534), .B(n2174), .Z(n1708) );
  AND U2568 ( .A(n1707), .B(n1708), .Z(n20561) );
  NANDN U2569 ( .A(n20702), .B(n2173), .Z(n1709) );
  NANDN U2570 ( .A(n20681), .B(n2174), .Z(n1710) );
  AND U2571 ( .A(n1709), .B(n1710), .Z(n20708) );
  NANDN U2572 ( .A(n20849), .B(n2173), .Z(n1711) );
  NANDN U2573 ( .A(n20828), .B(n2174), .Z(n1712) );
  AND U2574 ( .A(n1711), .B(n1712), .Z(n20855) );
  NANDN U2575 ( .A(n20996), .B(n2173), .Z(n1713) );
  NANDN U2576 ( .A(n20975), .B(n2174), .Z(n1714) );
  AND U2577 ( .A(n1713), .B(n1714), .Z(n21002) );
  NANDN U2578 ( .A(n21139), .B(n2173), .Z(n1715) );
  NANDN U2579 ( .A(n21118), .B(n2174), .Z(n1716) );
  AND U2580 ( .A(n1715), .B(n1716), .Z(n21145) );
  NANDN U2581 ( .A(n21244), .B(n2173), .Z(n1717) );
  NANDN U2582 ( .A(n21223), .B(n2174), .Z(n1718) );
  AND U2583 ( .A(n1717), .B(n1718), .Z(n21250) );
  NANDN U2584 ( .A(n21429), .B(n2173), .Z(n1719) );
  NANDN U2585 ( .A(n21408), .B(n2174), .Z(n1720) );
  AND U2586 ( .A(n1719), .B(n1720), .Z(n21435) );
  NANDN U2587 ( .A(n21576), .B(n2173), .Z(n1721) );
  NANDN U2588 ( .A(n21555), .B(n2174), .Z(n1722) );
  AND U2589 ( .A(n1721), .B(n1722), .Z(n21582) );
  NANDN U2590 ( .A(n21723), .B(n2173), .Z(n1723) );
  NANDN U2591 ( .A(n21702), .B(n2174), .Z(n1724) );
  AND U2592 ( .A(n1723), .B(n1724), .Z(n21729) );
  NANDN U2593 ( .A(n21870), .B(n2173), .Z(n1725) );
  NANDN U2594 ( .A(n21849), .B(n2174), .Z(n1726) );
  AND U2595 ( .A(n1725), .B(n1726), .Z(n21876) );
  NANDN U2596 ( .A(n22017), .B(n2173), .Z(n1727) );
  NANDN U2597 ( .A(n21996), .B(n2174), .Z(n1728) );
  AND U2598 ( .A(n1727), .B(n1728), .Z(n22023) );
  NANDN U2599 ( .A(n22164), .B(n2173), .Z(n1729) );
  NANDN U2600 ( .A(n22143), .B(n2174), .Z(n1730) );
  AND U2601 ( .A(n1729), .B(n1730), .Z(n22170) );
  NANDN U2602 ( .A(n22290), .B(n2173), .Z(n1731) );
  NANDN U2603 ( .A(n22269), .B(n2174), .Z(n1732) );
  AND U2604 ( .A(n1731), .B(n1732), .Z(n22296) );
  NANDN U2605 ( .A(n22454), .B(n2173), .Z(n1733) );
  NANDN U2606 ( .A(n22433), .B(n2174), .Z(n1734) );
  AND U2607 ( .A(n1733), .B(n1734), .Z(n22460) );
  NANDN U2608 ( .A(n22601), .B(n2173), .Z(n1735) );
  NANDN U2609 ( .A(n22580), .B(n2174), .Z(n1736) );
  AND U2610 ( .A(n1735), .B(n1736), .Z(n22607) );
  NANDN U2611 ( .A(n22748), .B(n2173), .Z(n1737) );
  NANDN U2612 ( .A(n22727), .B(n2174), .Z(n1738) );
  AND U2613 ( .A(n1737), .B(n1738), .Z(n22754) );
  NANDN U2614 ( .A(n22895), .B(n2173), .Z(n1739) );
  NANDN U2615 ( .A(n22874), .B(n2174), .Z(n1740) );
  AND U2616 ( .A(n1739), .B(n1740), .Z(n22901) );
  NANDN U2617 ( .A(n23042), .B(n2173), .Z(n1741) );
  NANDN U2618 ( .A(n23021), .B(n2174), .Z(n1742) );
  AND U2619 ( .A(n1741), .B(n1742), .Z(n23048) );
  NANDN U2620 ( .A(n23189), .B(n2173), .Z(n1743) );
  NANDN U2621 ( .A(n23168), .B(n2174), .Z(n1744) );
  AND U2622 ( .A(n1743), .B(n1744), .Z(n23195) );
  NANDN U2623 ( .A(n23336), .B(n2173), .Z(n1745) );
  NANDN U2624 ( .A(n23315), .B(n2174), .Z(n1746) );
  AND U2625 ( .A(n1745), .B(n1746), .Z(n23342) );
  NANDN U2626 ( .A(n23483), .B(n2173), .Z(n1747) );
  NANDN U2627 ( .A(n23462), .B(n2174), .Z(n1748) );
  AND U2628 ( .A(n1747), .B(n1748), .Z(n23489) );
  OR U2629 ( .A(n2171), .B(n23644), .Z(n1749) );
  NANDN U2630 ( .A(n23623), .B(n2174), .Z(n1750) );
  AND U2631 ( .A(n1749), .B(n1750), .Z(n23652) );
  NANDN U2632 ( .A(n4404), .B(n4405), .Z(n1751) );
  NANDN U2633 ( .A(n4407), .B(n4406), .Z(n1752) );
  AND U2634 ( .A(n1751), .B(n1752), .Z(n4423) );
  NANDN U2635 ( .A(n6416), .B(n6417), .Z(n1753) );
  NANDN U2636 ( .A(n6419), .B(n6418), .Z(n1754) );
  AND U2637 ( .A(n1753), .B(n1754), .Z(n6435) );
  NANDN U2638 ( .A(n6832), .B(n6833), .Z(n1755) );
  NANDN U2639 ( .A(n6835), .B(n6834), .Z(n1756) );
  AND U2640 ( .A(n1755), .B(n1756), .Z(n6851) );
  NANDN U2641 ( .A(n6933), .B(n6934), .Z(n1757) );
  NANDN U2642 ( .A(n6936), .B(n6935), .Z(n1758) );
  AND U2643 ( .A(n1757), .B(n1758), .Z(n6952) );
  NANDN U2644 ( .A(n7097), .B(n7098), .Z(n1759) );
  NANDN U2645 ( .A(n7100), .B(n7099), .Z(n1760) );
  AND U2646 ( .A(n1759), .B(n1760), .Z(n7116) );
  NANDN U2647 ( .A(n7534), .B(n7535), .Z(n1761) );
  NANDN U2648 ( .A(n7537), .B(n7536), .Z(n1762) );
  AND U2649 ( .A(n1761), .B(n1762), .Z(n7553) );
  NANDN U2650 ( .A(n7803), .B(n7804), .Z(n1763) );
  NANDN U2651 ( .A(n7806), .B(n7805), .Z(n1764) );
  AND U2652 ( .A(n1763), .B(n1764), .Z(n7822) );
  NANDN U2653 ( .A(n7925), .B(n7926), .Z(n1765) );
  NANDN U2654 ( .A(n7928), .B(n7927), .Z(n1766) );
  AND U2655 ( .A(n1765), .B(n1766), .Z(n7944) );
  NANDN U2656 ( .A(n8194), .B(n8195), .Z(n1767) );
  NANDN U2657 ( .A(n8197), .B(n8196), .Z(n1768) );
  AND U2658 ( .A(n1767), .B(n1768), .Z(n8213) );
  NANDN U2659 ( .A(n9051), .B(n9052), .Z(n1769) );
  NANDN U2660 ( .A(n9054), .B(n9053), .Z(n1770) );
  AND U2661 ( .A(n1769), .B(n1770), .Z(n9070) );
  NANDN U2662 ( .A(n9194), .B(n9195), .Z(n1771) );
  NANDN U2663 ( .A(n9197), .B(n9196), .Z(n1772) );
  AND U2664 ( .A(n1771), .B(n1772), .Z(n9213) );
  NANDN U2665 ( .A(n11790), .B(n11791), .Z(n1773) );
  NANDN U2666 ( .A(n11793), .B(n11792), .Z(n1774) );
  AND U2667 ( .A(n1773), .B(n1774), .Z(n11809) );
  NANDN U2668 ( .A(n12647), .B(n12648), .Z(n1775) );
  NANDN U2669 ( .A(n12650), .B(n12649), .Z(n1776) );
  AND U2670 ( .A(n1775), .B(n1776), .Z(n12666) );
  NANDN U2671 ( .A(n13819), .B(n13820), .Z(n1777) );
  NANDN U2672 ( .A(n13822), .B(n13821), .Z(n1778) );
  AND U2673 ( .A(n1777), .B(n1778), .Z(n13838) );
  NANDN U2674 ( .A(n14760), .B(n14761), .Z(n1779) );
  NANDN U2675 ( .A(n14763), .B(n14762), .Z(n1780) );
  AND U2676 ( .A(n1779), .B(n1780), .Z(n14779) );
  NANDN U2677 ( .A(n15617), .B(n15618), .Z(n1781) );
  NANDN U2678 ( .A(n15620), .B(n15619), .Z(n1782) );
  AND U2679 ( .A(n1781), .B(n1782), .Z(n15636) );
  NANDN U2680 ( .A(n17772), .B(n17773), .Z(n1783) );
  NANDN U2681 ( .A(n17775), .B(n17774), .Z(n1784) );
  AND U2682 ( .A(n1783), .B(n1784), .Z(n17791) );
  NANDN U2683 ( .A(n18104), .B(n18105), .Z(n1785) );
  NANDN U2684 ( .A(n18107), .B(n18106), .Z(n1786) );
  AND U2685 ( .A(n1785), .B(n1786), .Z(n18123) );
  NANDN U2686 ( .A(n19696), .B(n19697), .Z(n1787) );
  NANDN U2687 ( .A(n19699), .B(n19698), .Z(n1788) );
  AND U2688 ( .A(n1787), .B(n1788), .Z(n19715) );
  NANDN U2689 ( .A(n20133), .B(n20134), .Z(n1789) );
  NANDN U2690 ( .A(n20136), .B(n20135), .Z(n1790) );
  AND U2691 ( .A(n1789), .B(n1790), .Z(n20152) );
  NANDN U2692 ( .A(n21032), .B(n21033), .Z(n1791) );
  NANDN U2693 ( .A(n21035), .B(n21034), .Z(n1792) );
  AND U2694 ( .A(n1791), .B(n1792), .Z(n21051) );
  NANDN U2695 ( .A(n21280), .B(n21281), .Z(n1793) );
  NANDN U2696 ( .A(n21283), .B(n21282), .Z(n1794) );
  AND U2697 ( .A(n1793), .B(n1794), .Z(n21299) );
  NANDN U2698 ( .A(n22326), .B(n22327), .Z(n1795) );
  NANDN U2699 ( .A(n22329), .B(n22328), .Z(n1796) );
  AND U2700 ( .A(n1795), .B(n1796), .Z(n22345) );
  NANDN U2701 ( .A(n23600), .B(n23601), .Z(n1797) );
  NANDN U2702 ( .A(n23603), .B(n23602), .Z(n1798) );
  AND U2703 ( .A(n1797), .B(n1798), .Z(n23619) );
  NANDN U2704 ( .A(n23687), .B(n23688), .Z(n1799) );
  NANDN U2705 ( .A(n23689), .B(n23690), .Z(n1800) );
  AND U2706 ( .A(n1799), .B(n1800), .Z(n23695) );
  XOR U2707 ( .A(n2368), .B(sreg[1023]), .Z(n1801) );
  NAND U2708 ( .A(n1801), .B(n2367), .Z(n1802) );
  NAND U2709 ( .A(n2368), .B(sreg[1023]), .Z(n1803) );
  AND U2710 ( .A(n1802), .B(n1803), .Z(n2370) );
  NAND U2711 ( .A(n11768), .B(n11767), .Z(n1804) );
  NANDN U2712 ( .A(n11766), .B(sreg[1473]), .Z(n1805) );
  NAND U2713 ( .A(n1804), .B(n1805), .Z(n11786) );
  NAND U2714 ( .A(n17750), .B(n17749), .Z(n1806) );
  NANDN U2715 ( .A(n17748), .B(sreg[1759]), .Z(n1807) );
  NAND U2716 ( .A(n1806), .B(n1807), .Z(n17768) );
  NAND U2717 ( .A(n23599), .B(n23598), .Z(n1808) );
  NANDN U2718 ( .A(n23597), .B(sreg[2039]), .Z(n1809) );
  NAND U2719 ( .A(n1808), .B(n1809), .Z(n23615) );
  NAND U2720 ( .A(n23678), .B(n23677), .Z(n1810) );
  NANDN U2721 ( .A(n23676), .B(sreg[2043]), .Z(n1811) );
  NAND U2722 ( .A(n1810), .B(n1811), .Z(n23679) );
  NANDN U2723 ( .A(n2436), .B(n2173), .Z(n1812) );
  NANDN U2724 ( .A(n2415), .B(n2174), .Z(n1813) );
  AND U2725 ( .A(n1812), .B(n1813), .Z(n2442) );
  NANDN U2726 ( .A(n2583), .B(n2173), .Z(n1814) );
  NANDN U2727 ( .A(n2562), .B(n2174), .Z(n1815) );
  AND U2728 ( .A(n1814), .B(n1815), .Z(n2589) );
  NANDN U2729 ( .A(n2730), .B(n2173), .Z(n1816) );
  NANDN U2730 ( .A(n2709), .B(n2174), .Z(n1817) );
  AND U2731 ( .A(n1816), .B(n1817), .Z(n2736) );
  NANDN U2732 ( .A(n2877), .B(n2173), .Z(n1818) );
  NANDN U2733 ( .A(n2856), .B(n2174), .Z(n1819) );
  AND U2734 ( .A(n1818), .B(n1819), .Z(n2883) );
  NANDN U2735 ( .A(n3024), .B(n2173), .Z(n1820) );
  NANDN U2736 ( .A(n3003), .B(n2174), .Z(n1821) );
  AND U2737 ( .A(n1820), .B(n1821), .Z(n3030) );
  NANDN U2738 ( .A(n3171), .B(n2173), .Z(n1822) );
  NANDN U2739 ( .A(n3150), .B(n2174), .Z(n1823) );
  AND U2740 ( .A(n1822), .B(n1823), .Z(n3177) );
  NANDN U2741 ( .A(n3318), .B(n2173), .Z(n1824) );
  NANDN U2742 ( .A(n3297), .B(n2174), .Z(n1825) );
  AND U2743 ( .A(n1824), .B(n1825), .Z(n3324) );
  NANDN U2744 ( .A(n3465), .B(n2173), .Z(n1826) );
  NANDN U2745 ( .A(n3444), .B(n2174), .Z(n1827) );
  AND U2746 ( .A(n1826), .B(n1827), .Z(n3471) );
  NANDN U2747 ( .A(n3612), .B(n2173), .Z(n1828) );
  NANDN U2748 ( .A(n3591), .B(n2174), .Z(n1829) );
  AND U2749 ( .A(n1828), .B(n1829), .Z(n3618) );
  NANDN U2750 ( .A(n3759), .B(n2173), .Z(n1830) );
  NANDN U2751 ( .A(n3738), .B(n2174), .Z(n1831) );
  AND U2752 ( .A(n1830), .B(n1831), .Z(n3765) );
  NANDN U2753 ( .A(n3906), .B(n2173), .Z(n1832) );
  NANDN U2754 ( .A(n3885), .B(n2174), .Z(n1833) );
  AND U2755 ( .A(n1832), .B(n1833), .Z(n3912) );
  NANDN U2756 ( .A(n4053), .B(n2173), .Z(n1834) );
  NANDN U2757 ( .A(n4032), .B(n2174), .Z(n1835) );
  AND U2758 ( .A(n1834), .B(n1835), .Z(n4059) );
  NANDN U2759 ( .A(n4200), .B(n2173), .Z(n1836) );
  NANDN U2760 ( .A(n4179), .B(n2174), .Z(n1837) );
  AND U2761 ( .A(n1836), .B(n1837), .Z(n4206) );
  NANDN U2762 ( .A(n4347), .B(n2173), .Z(n1838) );
  NANDN U2763 ( .A(n4326), .B(n2174), .Z(n1839) );
  AND U2764 ( .A(n1838), .B(n1839), .Z(n4353) );
  NANDN U2765 ( .A(n4490), .B(n2173), .Z(n1840) );
  NANDN U2766 ( .A(n4469), .B(n2174), .Z(n1841) );
  AND U2767 ( .A(n1840), .B(n1841), .Z(n4496) );
  NANDN U2768 ( .A(n4637), .B(n2173), .Z(n1842) );
  NANDN U2769 ( .A(n4616), .B(n2174), .Z(n1843) );
  AND U2770 ( .A(n1842), .B(n1843), .Z(n4643) );
  NANDN U2771 ( .A(n4784), .B(n2173), .Z(n1844) );
  NANDN U2772 ( .A(n4763), .B(n2174), .Z(n1845) );
  AND U2773 ( .A(n1844), .B(n1845), .Z(n4790) );
  NANDN U2774 ( .A(n4931), .B(n2173), .Z(n1846) );
  NANDN U2775 ( .A(n4910), .B(n2174), .Z(n1847) );
  AND U2776 ( .A(n1846), .B(n1847), .Z(n4937) );
  NANDN U2777 ( .A(n5078), .B(n2173), .Z(n1848) );
  NANDN U2778 ( .A(n5057), .B(n2174), .Z(n1849) );
  AND U2779 ( .A(n1848), .B(n1849), .Z(n5084) );
  NANDN U2780 ( .A(n5225), .B(n2173), .Z(n1850) );
  NANDN U2781 ( .A(n5204), .B(n2174), .Z(n1851) );
  AND U2782 ( .A(n1850), .B(n1851), .Z(n5231) );
  NANDN U2783 ( .A(n5372), .B(n2173), .Z(n1852) );
  NANDN U2784 ( .A(n5351), .B(n2174), .Z(n1853) );
  AND U2785 ( .A(n1852), .B(n1853), .Z(n5378) );
  NANDN U2786 ( .A(n5519), .B(n2173), .Z(n1854) );
  NANDN U2787 ( .A(n5498), .B(n2174), .Z(n1855) );
  AND U2788 ( .A(n1854), .B(n1855), .Z(n5525) );
  NANDN U2789 ( .A(n5666), .B(n2173), .Z(n1856) );
  NANDN U2790 ( .A(n5645), .B(n2174), .Z(n1857) );
  AND U2791 ( .A(n1856), .B(n1857), .Z(n5672) );
  NANDN U2792 ( .A(n5813), .B(n2173), .Z(n1858) );
  NANDN U2793 ( .A(n5792), .B(n2174), .Z(n1859) );
  AND U2794 ( .A(n1858), .B(n1859), .Z(n5819) );
  NANDN U2795 ( .A(n5960), .B(n2173), .Z(n1860) );
  NANDN U2796 ( .A(n5939), .B(n2174), .Z(n1861) );
  AND U2797 ( .A(n1860), .B(n1861), .Z(n5966) );
  NANDN U2798 ( .A(n6107), .B(n2173), .Z(n1862) );
  NANDN U2799 ( .A(n6086), .B(n2174), .Z(n1863) );
  AND U2800 ( .A(n1862), .B(n1863), .Z(n6113) );
  NANDN U2801 ( .A(n6254), .B(n2173), .Z(n1864) );
  NANDN U2802 ( .A(n6233), .B(n2174), .Z(n1865) );
  AND U2803 ( .A(n1864), .B(n1865), .Z(n6260) );
  NANDN U2804 ( .A(n6401), .B(n2173), .Z(n1866) );
  NANDN U2805 ( .A(n6380), .B(n2174), .Z(n1867) );
  AND U2806 ( .A(n1866), .B(n1867), .Z(n6407) );
  NANDN U2807 ( .A(n6544), .B(n2173), .Z(n1868) );
  NANDN U2808 ( .A(n6523), .B(n2174), .Z(n1869) );
  AND U2809 ( .A(n1868), .B(n1869), .Z(n6550) );
  NANDN U2810 ( .A(n6691), .B(n2173), .Z(n1870) );
  NANDN U2811 ( .A(n6670), .B(n2174), .Z(n1871) );
  AND U2812 ( .A(n1870), .B(n1871), .Z(n6697) );
  NANDN U2813 ( .A(n6836), .B(n2173), .Z(n1872) );
  NANDN U2814 ( .A(n6817), .B(n2174), .Z(n1873) );
  AND U2815 ( .A(n1872), .B(n1873), .Z(n6843) );
  NANDN U2816 ( .A(n6977), .B(n2173), .Z(n1874) );
  NANDN U2817 ( .A(n6956), .B(n2174), .Z(n1875) );
  AND U2818 ( .A(n1874), .B(n1875), .Z(n6983) );
  NANDN U2819 ( .A(n7120), .B(n2173), .Z(n1876) );
  NANDN U2820 ( .A(n7101), .B(n2174), .Z(n1877) );
  AND U2821 ( .A(n1876), .B(n1877), .Z(n7126) );
  NANDN U2822 ( .A(n7267), .B(n2173), .Z(n1878) );
  NANDN U2823 ( .A(n7246), .B(n2174), .Z(n1879) );
  AND U2824 ( .A(n1878), .B(n1879), .Z(n7273) );
  NANDN U2825 ( .A(n7414), .B(n2173), .Z(n1880) );
  NANDN U2826 ( .A(n7393), .B(n2174), .Z(n1881) );
  AND U2827 ( .A(n1880), .B(n1881), .Z(n7420) );
  NANDN U2828 ( .A(n7557), .B(n2173), .Z(n1882) );
  NANDN U2829 ( .A(n7538), .B(n2174), .Z(n1883) );
  AND U2830 ( .A(n1882), .B(n1883), .Z(n7563) );
  NANDN U2831 ( .A(n7704), .B(n2173), .Z(n1884) );
  NANDN U2832 ( .A(n7683), .B(n2174), .Z(n1885) );
  AND U2833 ( .A(n1884), .B(n1885), .Z(n7710) );
  NANDN U2834 ( .A(n7847), .B(n2173), .Z(n1886) );
  NANDN U2835 ( .A(n7826), .B(n2174), .Z(n1887) );
  AND U2836 ( .A(n1886), .B(n1887), .Z(n7853) );
  NANDN U2837 ( .A(n7990), .B(n2173), .Z(n1888) );
  NANDN U2838 ( .A(n7969), .B(n2174), .Z(n1889) );
  AND U2839 ( .A(n1888), .B(n1889), .Z(n7996) );
  NANDN U2840 ( .A(n8137), .B(n2173), .Z(n1890) );
  NANDN U2841 ( .A(n8116), .B(n2174), .Z(n1891) );
  AND U2842 ( .A(n1890), .B(n1891), .Z(n8143) );
  NANDN U2843 ( .A(n8280), .B(n2173), .Z(n1892) );
  NANDN U2844 ( .A(n8259), .B(n2174), .Z(n1893) );
  AND U2845 ( .A(n1892), .B(n1893), .Z(n8286) );
  NANDN U2846 ( .A(n8427), .B(n2173), .Z(n1894) );
  NANDN U2847 ( .A(n8406), .B(n2174), .Z(n1895) );
  AND U2848 ( .A(n1894), .B(n1895), .Z(n8433) );
  NANDN U2849 ( .A(n8574), .B(n2173), .Z(n1896) );
  NANDN U2850 ( .A(n8553), .B(n2174), .Z(n1897) );
  AND U2851 ( .A(n1896), .B(n1897), .Z(n8580) );
  NANDN U2852 ( .A(n8721), .B(n2173), .Z(n1898) );
  NANDN U2853 ( .A(n8700), .B(n2174), .Z(n1899) );
  AND U2854 ( .A(n1898), .B(n1899), .Z(n8727) );
  NANDN U2855 ( .A(n8868), .B(n2173), .Z(n1900) );
  NANDN U2856 ( .A(n8847), .B(n2174), .Z(n1901) );
  AND U2857 ( .A(n1900), .B(n1901), .Z(n8874) );
  NANDN U2858 ( .A(n9015), .B(n2173), .Z(n1902) );
  NANDN U2859 ( .A(n8994), .B(n2174), .Z(n1903) );
  AND U2860 ( .A(n1902), .B(n1903), .Z(n9021) );
  NANDN U2861 ( .A(n9158), .B(n2173), .Z(n1904) );
  NANDN U2862 ( .A(n9137), .B(n2174), .Z(n1905) );
  AND U2863 ( .A(n1904), .B(n1905), .Z(n9164) );
  NANDN U2864 ( .A(n9301), .B(n2173), .Z(n1906) );
  NANDN U2865 ( .A(n9280), .B(n2174), .Z(n1907) );
  AND U2866 ( .A(n1906), .B(n1907), .Z(n9307) );
  NANDN U2867 ( .A(n9448), .B(n2173), .Z(n1908) );
  NANDN U2868 ( .A(n9427), .B(n2174), .Z(n1909) );
  AND U2869 ( .A(n1908), .B(n1909), .Z(n9454) );
  NANDN U2870 ( .A(n9595), .B(n2173), .Z(n1910) );
  NANDN U2871 ( .A(n9574), .B(n2174), .Z(n1911) );
  AND U2872 ( .A(n1910), .B(n1911), .Z(n9601) );
  NANDN U2873 ( .A(n9742), .B(n2173), .Z(n1912) );
  NANDN U2874 ( .A(n9721), .B(n2174), .Z(n1913) );
  AND U2875 ( .A(n1912), .B(n1913), .Z(n9748) );
  NANDN U2876 ( .A(n9889), .B(n2173), .Z(n1914) );
  NANDN U2877 ( .A(n9868), .B(n2174), .Z(n1915) );
  AND U2878 ( .A(n1914), .B(n1915), .Z(n9895) );
  NANDN U2879 ( .A(n10036), .B(n2173), .Z(n1916) );
  NANDN U2880 ( .A(n10015), .B(n2174), .Z(n1917) );
  AND U2881 ( .A(n1916), .B(n1917), .Z(n10042) );
  NANDN U2882 ( .A(n10183), .B(n2173), .Z(n1918) );
  NANDN U2883 ( .A(n10162), .B(n2174), .Z(n1919) );
  AND U2884 ( .A(n1918), .B(n1919), .Z(n10189) );
  NANDN U2885 ( .A(n10330), .B(n2173), .Z(n1920) );
  NANDN U2886 ( .A(n10309), .B(n2174), .Z(n1921) );
  AND U2887 ( .A(n1920), .B(n1921), .Z(n10336) );
  NANDN U2888 ( .A(n10477), .B(n2173), .Z(n1922) );
  NANDN U2889 ( .A(n10456), .B(n2174), .Z(n1923) );
  AND U2890 ( .A(n1922), .B(n1923), .Z(n10483) );
  NANDN U2891 ( .A(n10624), .B(n2173), .Z(n1924) );
  NANDN U2892 ( .A(n10603), .B(n2174), .Z(n1925) );
  AND U2893 ( .A(n1924), .B(n1925), .Z(n10630) );
  NANDN U2894 ( .A(n10771), .B(n2173), .Z(n1926) );
  NANDN U2895 ( .A(n10750), .B(n2174), .Z(n1927) );
  AND U2896 ( .A(n1926), .B(n1927), .Z(n10777) );
  NANDN U2897 ( .A(n10918), .B(n2173), .Z(n1928) );
  NANDN U2898 ( .A(n10897), .B(n2174), .Z(n1929) );
  AND U2899 ( .A(n1928), .B(n1929), .Z(n10924) );
  NANDN U2900 ( .A(n11065), .B(n2173), .Z(n1930) );
  NANDN U2901 ( .A(n11044), .B(n2174), .Z(n1931) );
  AND U2902 ( .A(n1930), .B(n1931), .Z(n11071) );
  NANDN U2903 ( .A(n11212), .B(n2173), .Z(n1932) );
  NANDN U2904 ( .A(n11191), .B(n2174), .Z(n1933) );
  AND U2905 ( .A(n1932), .B(n1933), .Z(n11218) );
  NANDN U2906 ( .A(n11359), .B(n2173), .Z(n1934) );
  NANDN U2907 ( .A(n11338), .B(n2174), .Z(n1935) );
  AND U2908 ( .A(n1934), .B(n1935), .Z(n11365) );
  NANDN U2909 ( .A(n11506), .B(n2173), .Z(n1936) );
  NANDN U2910 ( .A(n11485), .B(n2174), .Z(n1937) );
  AND U2911 ( .A(n1936), .B(n1937), .Z(n11512) );
  NANDN U2912 ( .A(n11653), .B(n2173), .Z(n1938) );
  NANDN U2913 ( .A(n11632), .B(n2174), .Z(n1939) );
  AND U2914 ( .A(n1938), .B(n1939), .Z(n11659) );
  NANDN U2915 ( .A(n11794), .B(n2173), .Z(n1940) );
  NANDN U2916 ( .A(n11775), .B(n2174), .Z(n1941) );
  AND U2917 ( .A(n1940), .B(n1941), .Z(n11801) );
  NANDN U2918 ( .A(n11939), .B(n2173), .Z(n1942) );
  NANDN U2919 ( .A(n11918), .B(n2174), .Z(n1943) );
  AND U2920 ( .A(n1942), .B(n1943), .Z(n11945) );
  NANDN U2921 ( .A(n12086), .B(n2173), .Z(n1944) );
  NANDN U2922 ( .A(n12065), .B(n2174), .Z(n1945) );
  AND U2923 ( .A(n1944), .B(n1945), .Z(n12092) );
  NANDN U2924 ( .A(n12233), .B(n2173), .Z(n1946) );
  NANDN U2925 ( .A(n12212), .B(n2174), .Z(n1947) );
  AND U2926 ( .A(n1946), .B(n1947), .Z(n12239) );
  NANDN U2927 ( .A(n12380), .B(n2173), .Z(n1948) );
  NANDN U2928 ( .A(n12359), .B(n2174), .Z(n1949) );
  AND U2929 ( .A(n1948), .B(n1949), .Z(n12386) );
  NANDN U2930 ( .A(n12527), .B(n2173), .Z(n1950) );
  NANDN U2931 ( .A(n12506), .B(n2174), .Z(n1951) );
  AND U2932 ( .A(n1950), .B(n1951), .Z(n12533) );
  NANDN U2933 ( .A(n12670), .B(n2173), .Z(n1952) );
  NANDN U2934 ( .A(n12651), .B(n2174), .Z(n1953) );
  AND U2935 ( .A(n1952), .B(n1953), .Z(n12676) );
  NANDN U2936 ( .A(n12817), .B(n2173), .Z(n1954) );
  NANDN U2937 ( .A(n12796), .B(n2174), .Z(n1955) );
  AND U2938 ( .A(n1954), .B(n1955), .Z(n12823) );
  NANDN U2939 ( .A(n12964), .B(n2173), .Z(n1956) );
  NANDN U2940 ( .A(n12943), .B(n2174), .Z(n1957) );
  AND U2941 ( .A(n1956), .B(n1957), .Z(n12970) );
  NANDN U2942 ( .A(n13111), .B(n2173), .Z(n1958) );
  NANDN U2943 ( .A(n13090), .B(n2174), .Z(n1959) );
  AND U2944 ( .A(n1958), .B(n1959), .Z(n13117) );
  NANDN U2945 ( .A(n13258), .B(n2173), .Z(n1960) );
  NANDN U2946 ( .A(n13237), .B(n2174), .Z(n1961) );
  AND U2947 ( .A(n1960), .B(n1961), .Z(n13264) );
  NANDN U2948 ( .A(n13405), .B(n2173), .Z(n1962) );
  NANDN U2949 ( .A(n13384), .B(n2174), .Z(n1963) );
  AND U2950 ( .A(n1962), .B(n1963), .Z(n13411) );
  NANDN U2951 ( .A(n13552), .B(n2173), .Z(n1964) );
  NANDN U2952 ( .A(n13531), .B(n2174), .Z(n1965) );
  AND U2953 ( .A(n1964), .B(n1965), .Z(n13558) );
  NANDN U2954 ( .A(n13699), .B(n2173), .Z(n1966) );
  NANDN U2955 ( .A(n13678), .B(n2174), .Z(n1967) );
  AND U2956 ( .A(n1966), .B(n1967), .Z(n13705) );
  NANDN U2957 ( .A(n13842), .B(n2173), .Z(n1968) );
  NANDN U2958 ( .A(n13823), .B(n2174), .Z(n1969) );
  AND U2959 ( .A(n1968), .B(n1969), .Z(n13848) );
  NANDN U2960 ( .A(n13989), .B(n2173), .Z(n1970) );
  NANDN U2961 ( .A(n13968), .B(n2174), .Z(n1971) );
  AND U2962 ( .A(n1970), .B(n1971), .Z(n13995) );
  NANDN U2963 ( .A(n14136), .B(n2173), .Z(n1972) );
  NANDN U2964 ( .A(n14115), .B(n2174), .Z(n1973) );
  AND U2965 ( .A(n1972), .B(n1973), .Z(n14142) );
  NANDN U2966 ( .A(n14283), .B(n2173), .Z(n1974) );
  NANDN U2967 ( .A(n14262), .B(n2174), .Z(n1975) );
  AND U2968 ( .A(n1974), .B(n1975), .Z(n14289) );
  NANDN U2969 ( .A(n14430), .B(n2173), .Z(n1976) );
  NANDN U2970 ( .A(n14409), .B(n2174), .Z(n1977) );
  AND U2971 ( .A(n1976), .B(n1977), .Z(n14436) );
  NANDN U2972 ( .A(n14577), .B(n2173), .Z(n1978) );
  NANDN U2973 ( .A(n14556), .B(n2174), .Z(n1979) );
  AND U2974 ( .A(n1978), .B(n1979), .Z(n14583) );
  NANDN U2975 ( .A(n14724), .B(n2173), .Z(n1980) );
  NANDN U2976 ( .A(n14703), .B(n2174), .Z(n1981) );
  AND U2977 ( .A(n1980), .B(n1981), .Z(n14730) );
  NANDN U2978 ( .A(n14867), .B(n2173), .Z(n1982) );
  NANDN U2979 ( .A(n14846), .B(n2174), .Z(n1983) );
  AND U2980 ( .A(n1982), .B(n1983), .Z(n14873) );
  NANDN U2981 ( .A(n15014), .B(n2173), .Z(n1984) );
  NANDN U2982 ( .A(n14993), .B(n2174), .Z(n1985) );
  AND U2983 ( .A(n1984), .B(n1985), .Z(n15020) );
  NANDN U2984 ( .A(n15161), .B(n2173), .Z(n1986) );
  NANDN U2985 ( .A(n15140), .B(n2174), .Z(n1987) );
  AND U2986 ( .A(n1986), .B(n1987), .Z(n15167) );
  NANDN U2987 ( .A(n15308), .B(n2173), .Z(n1988) );
  NANDN U2988 ( .A(n15287), .B(n2174), .Z(n1989) );
  AND U2989 ( .A(n1988), .B(n1989), .Z(n15314) );
  NANDN U2990 ( .A(n15455), .B(n2173), .Z(n1990) );
  NANDN U2991 ( .A(n15434), .B(n2174), .Z(n1991) );
  AND U2992 ( .A(n1990), .B(n1991), .Z(n15461) );
  NANDN U2993 ( .A(n15602), .B(n2173), .Z(n1992) );
  NANDN U2994 ( .A(n15581), .B(n2174), .Z(n1993) );
  AND U2995 ( .A(n1992), .B(n1993), .Z(n15608) );
  NANDN U2996 ( .A(n15745), .B(n2173), .Z(n1994) );
  NANDN U2997 ( .A(n15724), .B(n2174), .Z(n1995) );
  AND U2998 ( .A(n1994), .B(n1995), .Z(n15751) );
  NANDN U2999 ( .A(n15892), .B(n2173), .Z(n1996) );
  NANDN U3000 ( .A(n15871), .B(n2174), .Z(n1997) );
  AND U3001 ( .A(n1996), .B(n1997), .Z(n15898) );
  NANDN U3002 ( .A(n16039), .B(n2173), .Z(n1998) );
  NANDN U3003 ( .A(n16018), .B(n2174), .Z(n1999) );
  AND U3004 ( .A(n1998), .B(n1999), .Z(n16045) );
  NANDN U3005 ( .A(n16186), .B(n2173), .Z(n2000) );
  NANDN U3006 ( .A(n16165), .B(n2174), .Z(n2001) );
  AND U3007 ( .A(n2000), .B(n2001), .Z(n16192) );
  NANDN U3008 ( .A(n16333), .B(n2173), .Z(n2002) );
  NANDN U3009 ( .A(n16312), .B(n2174), .Z(n2003) );
  AND U3010 ( .A(n2002), .B(n2003), .Z(n16339) );
  NANDN U3011 ( .A(n16480), .B(n2173), .Z(n2004) );
  NANDN U3012 ( .A(n16459), .B(n2174), .Z(n2005) );
  AND U3013 ( .A(n2004), .B(n2005), .Z(n16486) );
  NANDN U3014 ( .A(n16627), .B(n2173), .Z(n2006) );
  NANDN U3015 ( .A(n16606), .B(n2174), .Z(n2007) );
  AND U3016 ( .A(n2006), .B(n2007), .Z(n16633) );
  NANDN U3017 ( .A(n16774), .B(n2173), .Z(n2008) );
  NANDN U3018 ( .A(n16753), .B(n2174), .Z(n2009) );
  AND U3019 ( .A(n2008), .B(n2009), .Z(n16780) );
  NANDN U3020 ( .A(n16921), .B(n2173), .Z(n2010) );
  NANDN U3021 ( .A(n16900), .B(n2174), .Z(n2011) );
  AND U3022 ( .A(n2010), .B(n2011), .Z(n16927) );
  NANDN U3023 ( .A(n17068), .B(n2173), .Z(n2012) );
  NANDN U3024 ( .A(n17047), .B(n2174), .Z(n2013) );
  AND U3025 ( .A(n2012), .B(n2013), .Z(n17074) );
  NANDN U3026 ( .A(n17215), .B(n2173), .Z(n2014) );
  NANDN U3027 ( .A(n17194), .B(n2174), .Z(n2015) );
  AND U3028 ( .A(n2014), .B(n2015), .Z(n17221) );
  NANDN U3029 ( .A(n17362), .B(n2173), .Z(n2016) );
  NANDN U3030 ( .A(n17341), .B(n2174), .Z(n2017) );
  AND U3031 ( .A(n2016), .B(n2017), .Z(n17368) );
  NANDN U3032 ( .A(n17509), .B(n2173), .Z(n2018) );
  NANDN U3033 ( .A(n17488), .B(n2174), .Z(n2019) );
  AND U3034 ( .A(n2018), .B(n2019), .Z(n17515) );
  NANDN U3035 ( .A(n17656), .B(n2173), .Z(n2020) );
  NANDN U3036 ( .A(n17635), .B(n2174), .Z(n2021) );
  AND U3037 ( .A(n2020), .B(n2021), .Z(n17662) );
  NANDN U3038 ( .A(n17795), .B(n2173), .Z(n2022) );
  NANDN U3039 ( .A(n17776), .B(n2174), .Z(n2023) );
  AND U3040 ( .A(n2022), .B(n2023), .Z(n17801) );
  NANDN U3041 ( .A(n17942), .B(n2173), .Z(n2024) );
  NANDN U3042 ( .A(n17921), .B(n2174), .Z(n2025) );
  AND U3043 ( .A(n2024), .B(n2025), .Z(n17948) );
  NANDN U3044 ( .A(n18089), .B(n2173), .Z(n2026) );
  NANDN U3045 ( .A(n18068), .B(n2174), .Z(n2027) );
  AND U3046 ( .A(n2026), .B(n2027), .Z(n18095) );
  NANDN U3047 ( .A(n18232), .B(n2173), .Z(n2028) );
  NANDN U3048 ( .A(n18211), .B(n2174), .Z(n2029) );
  AND U3049 ( .A(n2028), .B(n2029), .Z(n18238) );
  NANDN U3050 ( .A(n18379), .B(n2173), .Z(n2030) );
  NANDN U3051 ( .A(n18358), .B(n2174), .Z(n2031) );
  AND U3052 ( .A(n2030), .B(n2031), .Z(n18385) );
  NANDN U3053 ( .A(n18526), .B(n2173), .Z(n2032) );
  NANDN U3054 ( .A(n18505), .B(n2174), .Z(n2033) );
  AND U3055 ( .A(n2032), .B(n2033), .Z(n18532) );
  NANDN U3056 ( .A(n18673), .B(n2173), .Z(n2034) );
  NANDN U3057 ( .A(n18652), .B(n2174), .Z(n2035) );
  AND U3058 ( .A(n2034), .B(n2035), .Z(n18679) );
  NANDN U3059 ( .A(n18820), .B(n2173), .Z(n2036) );
  NANDN U3060 ( .A(n18799), .B(n2174), .Z(n2037) );
  AND U3061 ( .A(n2036), .B(n2037), .Z(n18826) );
  NANDN U3062 ( .A(n18967), .B(n2173), .Z(n2038) );
  NANDN U3063 ( .A(n18946), .B(n2174), .Z(n2039) );
  AND U3064 ( .A(n2038), .B(n2039), .Z(n18973) );
  NANDN U3065 ( .A(n19114), .B(n2173), .Z(n2040) );
  NANDN U3066 ( .A(n19093), .B(n2174), .Z(n2041) );
  AND U3067 ( .A(n2040), .B(n2041), .Z(n19120) );
  NANDN U3068 ( .A(n19261), .B(n2173), .Z(n2042) );
  NANDN U3069 ( .A(n19240), .B(n2174), .Z(n2043) );
  AND U3070 ( .A(n2042), .B(n2043), .Z(n19267) );
  NANDN U3071 ( .A(n19408), .B(n2173), .Z(n2044) );
  NANDN U3072 ( .A(n19387), .B(n2174), .Z(n2045) );
  AND U3073 ( .A(n2044), .B(n2045), .Z(n19414) );
  NANDN U3074 ( .A(n19555), .B(n2173), .Z(n2046) );
  NANDN U3075 ( .A(n19534), .B(n2174), .Z(n2047) );
  AND U3076 ( .A(n2046), .B(n2047), .Z(n19561) );
  NANDN U3077 ( .A(n19700), .B(n2173), .Z(n2048) );
  NANDN U3078 ( .A(n19681), .B(n2174), .Z(n2049) );
  AND U3079 ( .A(n2048), .B(n2049), .Z(n19707) );
  NANDN U3080 ( .A(n19845), .B(n2173), .Z(n2050) );
  NANDN U3081 ( .A(n19824), .B(n2174), .Z(n2051) );
  AND U3082 ( .A(n2050), .B(n2051), .Z(n19851) );
  NANDN U3083 ( .A(n19992), .B(n2173), .Z(n2052) );
  NANDN U3084 ( .A(n19971), .B(n2174), .Z(n2053) );
  AND U3085 ( .A(n2052), .B(n2053), .Z(n19998) );
  NANDN U3086 ( .A(n20137), .B(n2173), .Z(n2054) );
  NANDN U3087 ( .A(n20118), .B(n2174), .Z(n2055) );
  AND U3088 ( .A(n2054), .B(n2055), .Z(n20144) );
  NANDN U3089 ( .A(n20282), .B(n2173), .Z(n2056) );
  NANDN U3090 ( .A(n20261), .B(n2174), .Z(n2057) );
  AND U3091 ( .A(n2056), .B(n2057), .Z(n20288) );
  NANDN U3092 ( .A(n20429), .B(n2173), .Z(n2058) );
  NANDN U3093 ( .A(n20408), .B(n2174), .Z(n2059) );
  AND U3094 ( .A(n2058), .B(n2059), .Z(n20435) );
  NANDN U3095 ( .A(n20576), .B(n2173), .Z(n2060) );
  NANDN U3096 ( .A(n20555), .B(n2174), .Z(n2061) );
  AND U3097 ( .A(n2060), .B(n2061), .Z(n20582) );
  NANDN U3098 ( .A(n20723), .B(n2173), .Z(n2062) );
  NANDN U3099 ( .A(n20702), .B(n2174), .Z(n2063) );
  AND U3100 ( .A(n2062), .B(n2063), .Z(n20729) );
  NANDN U3101 ( .A(n20870), .B(n2173), .Z(n2064) );
  NANDN U3102 ( .A(n20849), .B(n2174), .Z(n2065) );
  AND U3103 ( .A(n2064), .B(n2065), .Z(n20876) );
  NANDN U3104 ( .A(n21017), .B(n2173), .Z(n2066) );
  NANDN U3105 ( .A(n20996), .B(n2174), .Z(n2067) );
  AND U3106 ( .A(n2066), .B(n2067), .Z(n21023) );
  NANDN U3107 ( .A(n21160), .B(n2173), .Z(n2068) );
  NANDN U3108 ( .A(n21139), .B(n2174), .Z(n2069) );
  AND U3109 ( .A(n2068), .B(n2069), .Z(n21166) );
  NANDN U3110 ( .A(n21303), .B(n2173), .Z(n2070) );
  NANDN U3111 ( .A(n21284), .B(n2174), .Z(n2071) );
  AND U3112 ( .A(n2070), .B(n2071), .Z(n21309) );
  NANDN U3113 ( .A(n21450), .B(n2173), .Z(n2072) );
  NANDN U3114 ( .A(n21429), .B(n2174), .Z(n2073) );
  AND U3115 ( .A(n2072), .B(n2073), .Z(n21456) );
  NANDN U3116 ( .A(n21597), .B(n2173), .Z(n2074) );
  NANDN U3117 ( .A(n21576), .B(n2174), .Z(n2075) );
  AND U3118 ( .A(n2074), .B(n2075), .Z(n21603) );
  NANDN U3119 ( .A(n21744), .B(n2173), .Z(n2076) );
  NANDN U3120 ( .A(n21723), .B(n2174), .Z(n2077) );
  AND U3121 ( .A(n2076), .B(n2077), .Z(n21750) );
  NANDN U3122 ( .A(n21891), .B(n2173), .Z(n2078) );
  NANDN U3123 ( .A(n21870), .B(n2174), .Z(n2079) );
  AND U3124 ( .A(n2078), .B(n2079), .Z(n21897) );
  NANDN U3125 ( .A(n22038), .B(n2173), .Z(n2080) );
  NANDN U3126 ( .A(n22017), .B(n2174), .Z(n2081) );
  AND U3127 ( .A(n2080), .B(n2081), .Z(n22044) );
  NANDN U3128 ( .A(n22185), .B(n2173), .Z(n2082) );
  NANDN U3129 ( .A(n22164), .B(n2174), .Z(n2083) );
  AND U3130 ( .A(n2082), .B(n2083), .Z(n22191) );
  NANDN U3131 ( .A(n22330), .B(n2173), .Z(n2084) );
  NANDN U3132 ( .A(n22311), .B(n2174), .Z(n2085) );
  AND U3133 ( .A(n2084), .B(n2085), .Z(n22337) );
  NANDN U3134 ( .A(n22475), .B(n2173), .Z(n2086) );
  NANDN U3135 ( .A(n22454), .B(n2174), .Z(n2087) );
  AND U3136 ( .A(n2086), .B(n2087), .Z(n22481) );
  NANDN U3137 ( .A(n22622), .B(n2173), .Z(n2088) );
  NANDN U3138 ( .A(n22601), .B(n2174), .Z(n2089) );
  AND U3139 ( .A(n2088), .B(n2089), .Z(n22628) );
  NANDN U3140 ( .A(n22769), .B(n2173), .Z(n2090) );
  NANDN U3141 ( .A(n22748), .B(n2174), .Z(n2091) );
  AND U3142 ( .A(n2090), .B(n2091), .Z(n22775) );
  NANDN U3143 ( .A(n22916), .B(n2173), .Z(n2092) );
  NANDN U3144 ( .A(n22895), .B(n2174), .Z(n2093) );
  AND U3145 ( .A(n2092), .B(n2093), .Z(n22922) );
  NANDN U3146 ( .A(n23063), .B(n2173), .Z(n2094) );
  NANDN U3147 ( .A(n23042), .B(n2174), .Z(n2095) );
  AND U3148 ( .A(n2094), .B(n2095), .Z(n23069) );
  NANDN U3149 ( .A(n23210), .B(n2173), .Z(n2096) );
  NANDN U3150 ( .A(n23189), .B(n2174), .Z(n2097) );
  AND U3151 ( .A(n2096), .B(n2097), .Z(n23216) );
  NANDN U3152 ( .A(n23357), .B(n2173), .Z(n2098) );
  NANDN U3153 ( .A(n23336), .B(n2174), .Z(n2099) );
  AND U3154 ( .A(n2098), .B(n2099), .Z(n23363) );
  NANDN U3155 ( .A(n23504), .B(n2173), .Z(n2100) );
  NANDN U3156 ( .A(n23483), .B(n2174), .Z(n2101) );
  AND U3157 ( .A(n2100), .B(n2101), .Z(n23510) );
  NANDN U3158 ( .A(n23623), .B(n2173), .Z(n2102) );
  NANDN U3159 ( .A(n23604), .B(n2174), .Z(n2103) );
  AND U3160 ( .A(n2102), .B(n2103), .Z(n23629) );
  NANDN U3161 ( .A(n23664), .B(n23663), .Z(n2104) );
  NANDN U3162 ( .A(n23661), .B(n23662), .Z(n2105) );
  NAND U3163 ( .A(n2104), .B(n2105), .Z(n23683) );
  NAND U3164 ( .A(n2371), .B(n2370), .Z(n2106) );
  XOR U3165 ( .A(n2371), .B(n2370), .Z(n2107) );
  NANDN U3166 ( .A(sreg[1024]), .B(n2107), .Z(n2108) );
  NAND U3167 ( .A(n2106), .B(n2108), .Z(n2406) );
  NAND U3168 ( .A(n4420), .B(n4419), .Z(n2109) );
  NANDN U3169 ( .A(n4418), .B(sreg[1121]), .Z(n2110) );
  NAND U3170 ( .A(n2109), .B(n2110), .Z(n4438) );
  NAND U3171 ( .A(n6432), .B(n6431), .Z(n2111) );
  NANDN U3172 ( .A(n6430), .B(sreg[1217]), .Z(n2112) );
  NAND U3173 ( .A(n2111), .B(n2112), .Z(n6450) );
  NAND U3174 ( .A(n6848), .B(n6847), .Z(n2113) );
  NANDN U3175 ( .A(n6846), .B(sreg[1237]), .Z(n2114) );
  NAND U3176 ( .A(n2113), .B(n2114), .Z(n6866) );
  NAND U3177 ( .A(n6949), .B(n6948), .Z(n2115) );
  NANDN U3178 ( .A(n6947), .B(sreg[1242]), .Z(n2116) );
  NAND U3179 ( .A(n2115), .B(n2116), .Z(n6967) );
  NAND U3180 ( .A(n7113), .B(n7112), .Z(n2117) );
  NANDN U3181 ( .A(n7111), .B(sreg[1250]), .Z(n2118) );
  NAND U3182 ( .A(n2117), .B(n2118), .Z(n7131) );
  NAND U3183 ( .A(n7550), .B(n7549), .Z(n2119) );
  NANDN U3184 ( .A(n7548), .B(sreg[1271]), .Z(n2120) );
  NAND U3185 ( .A(n2119), .B(n2120), .Z(n7568) );
  NAND U3186 ( .A(n7819), .B(n7818), .Z(n2121) );
  NANDN U3187 ( .A(n7817), .B(sreg[1284]), .Z(n2122) );
  NAND U3188 ( .A(n2121), .B(n2122), .Z(n7837) );
  NAND U3189 ( .A(n7941), .B(n7940), .Z(n2123) );
  NANDN U3190 ( .A(n7939), .B(sreg[1290]), .Z(n2124) );
  NAND U3191 ( .A(n2123), .B(n2124), .Z(n7959) );
  NAND U3192 ( .A(n8210), .B(n8209), .Z(n2125) );
  NANDN U3193 ( .A(n8208), .B(sreg[1303]), .Z(n2126) );
  NAND U3194 ( .A(n2125), .B(n2126), .Z(n8228) );
  NAND U3195 ( .A(n9067), .B(n9066), .Z(n2127) );
  NANDN U3196 ( .A(n9065), .B(sreg[1344]), .Z(n2128) );
  NAND U3197 ( .A(n2127), .B(n2128), .Z(n9085) );
  NAND U3198 ( .A(n9210), .B(n9209), .Z(n2129) );
  NANDN U3199 ( .A(n9208), .B(sreg[1351]), .Z(n2130) );
  NAND U3200 ( .A(n2129), .B(n2130), .Z(n9228) );
  NAND U3201 ( .A(n11806), .B(n11805), .Z(n2131) );
  NANDN U3202 ( .A(n11804), .B(sreg[1475]), .Z(n2132) );
  NAND U3203 ( .A(n2131), .B(n2132), .Z(n11824) );
  NAND U3204 ( .A(n12663), .B(n12662), .Z(n2133) );
  NANDN U3205 ( .A(n12661), .B(sreg[1516]), .Z(n2134) );
  NAND U3206 ( .A(n2133), .B(n2134), .Z(n12681) );
  NAND U3207 ( .A(n13835), .B(n13834), .Z(n2135) );
  NANDN U3208 ( .A(n13833), .B(sreg[1572]), .Z(n2136) );
  NAND U3209 ( .A(n2135), .B(n2136), .Z(n13853) );
  NAND U3210 ( .A(n14776), .B(n14775), .Z(n2137) );
  NANDN U3211 ( .A(n14774), .B(sreg[1617]), .Z(n2138) );
  NAND U3212 ( .A(n2137), .B(n2138), .Z(n14794) );
  NAND U3213 ( .A(n15633), .B(n15632), .Z(n2139) );
  NANDN U3214 ( .A(n15631), .B(sreg[1658]), .Z(n2140) );
  NAND U3215 ( .A(n2139), .B(n2140), .Z(n15651) );
  NAND U3216 ( .A(n17788), .B(n17787), .Z(n2141) );
  NANDN U3217 ( .A(n17786), .B(sreg[1761]), .Z(n2142) );
  NAND U3218 ( .A(n2141), .B(n2142), .Z(n17806) );
  NAND U3219 ( .A(n18120), .B(n18119), .Z(n2143) );
  NANDN U3220 ( .A(n18118), .B(sreg[1777]), .Z(n2144) );
  NAND U3221 ( .A(n2143), .B(n2144), .Z(n18138) );
  NAND U3222 ( .A(n19712), .B(n19711), .Z(n2145) );
  NANDN U3223 ( .A(n19710), .B(sreg[1853]), .Z(n2146) );
  NAND U3224 ( .A(n2145), .B(n2146), .Z(n19730) );
  NAND U3225 ( .A(n20149), .B(n20148), .Z(n2147) );
  NANDN U3226 ( .A(n20147), .B(sreg[1874]), .Z(n2148) );
  NAND U3227 ( .A(n2147), .B(n2148), .Z(n20167) );
  NAND U3228 ( .A(n21048), .B(n21047), .Z(n2149) );
  NANDN U3229 ( .A(n21046), .B(sreg[1917]), .Z(n2150) );
  NAND U3230 ( .A(n2149), .B(n2150), .Z(n21066) );
  NAND U3231 ( .A(n21296), .B(n21295), .Z(n2151) );
  NANDN U3232 ( .A(n21294), .B(sreg[1929]), .Z(n2152) );
  NAND U3233 ( .A(n2151), .B(n2152), .Z(n21314) );
  NAND U3234 ( .A(n22342), .B(n22341), .Z(n2153) );
  NANDN U3235 ( .A(n22340), .B(sreg[1979]), .Z(n2154) );
  NAND U3236 ( .A(n2153), .B(n2154), .Z(n22360) );
  NAND U3237 ( .A(n23616), .B(n23615), .Z(n2155) );
  NANDN U3238 ( .A(n23614), .B(sreg[2040]), .Z(n2156) );
  NAND U3239 ( .A(n2155), .B(n2156), .Z(n23634) );
  XNOR U3240 ( .A(n23712), .B(n23713), .Z(n2157) );
  NAND U3241 ( .A(n23714), .B(n2157), .Z(n2158) );
  NANDN U3242 ( .A(n23712), .B(n23713), .Z(n2159) );
  AND U3243 ( .A(n2158), .B(n2159), .Z(n2160) );
  XOR U3244 ( .A(n23714), .B(n2157), .Z(n2161) );
  NAND U3245 ( .A(n2161), .B(n23715), .Z(n2162) );
  NAND U3246 ( .A(n2160), .B(n2162), .Z(n2163) );
  NANDN U3247 ( .A(n23716), .B(n23717), .Z(n2164) );
  NANDN U3248 ( .A(n23718), .B(n23719), .Z(n2165) );
  AND U3249 ( .A(n2164), .B(n2165), .Z(n2166) );
  XNOR U3250 ( .A(a[1021]), .B(a[1023]), .Z(n2167) );
  XNOR U3251 ( .A(n23720), .B(n2167), .Z(n2168) );
  AND U3252 ( .A(n2168), .B(b[3]), .Z(n2169) );
  XNOR U3253 ( .A(n2163), .B(n2166), .Z(n2170) );
  XNOR U3254 ( .A(n2169), .B(n2170), .Z(c[2047]) );
  XNOR U3255 ( .A(b[1]), .B(b[2]), .Z(n2171) );
  NAND U3256 ( .A(n2344), .B(n2171), .Z(n2172) );
  IV U3257 ( .A(n2171), .Z(n2173) );
  IV U3258 ( .A(n2172), .Z(n2174) );
  IV U3259 ( .A(b[1]), .Z(n2175) );
  IV U3260 ( .A(b[3]), .Z(n2176) );
  IV U3261 ( .A(b[3]), .Z(n2177) );
  IV U3262 ( .A(b[3]), .Z(n2178) );
  IV U3263 ( .A(b[3]), .Z(n2179) );
  IV U3264 ( .A(b[3]), .Z(n2180) );
  IV U3265 ( .A(b[3]), .Z(n2181) );
  IV U3266 ( .A(b[3]), .Z(n2182) );
  IV U3267 ( .A(b[3]), .Z(n2183) );
  IV U3268 ( .A(b[3]), .Z(n2184) );
  IV U3269 ( .A(b[3]), .Z(n2185) );
  IV U3270 ( .A(b[3]), .Z(n2186) );
  IV U3271 ( .A(b[3]), .Z(n2187) );
  IV U3272 ( .A(b[3]), .Z(n2188) );
  IV U3273 ( .A(b[3]), .Z(n2189) );
  IV U3274 ( .A(b[3]), .Z(n2190) );
  IV U3275 ( .A(b[3]), .Z(n2191) );
  IV U3276 ( .A(b[3]), .Z(n2192) );
  IV U3277 ( .A(b[3]), .Z(n2193) );
  IV U3278 ( .A(b[3]), .Z(n2194) );
  IV U3279 ( .A(b[3]), .Z(n2195) );
  IV U3280 ( .A(b[3]), .Z(n2196) );
  IV U3281 ( .A(b[3]), .Z(n2197) );
  IV U3282 ( .A(b[3]), .Z(n2198) );
  IV U3283 ( .A(b[3]), .Z(n2199) );
  IV U3284 ( .A(b[3]), .Z(n2200) );
  IV U3285 ( .A(b[3]), .Z(n2201) );
  IV U3286 ( .A(b[3]), .Z(n2202) );
  IV U3287 ( .A(b[3]), .Z(n2203) );
  IV U3288 ( .A(b[3]), .Z(n2204) );
  IV U3289 ( .A(b[3]), .Z(n2205) );
  IV U3290 ( .A(b[3]), .Z(n2206) );
  IV U3291 ( .A(b[3]), .Z(n2207) );
  IV U3292 ( .A(b[3]), .Z(n2208) );
  IV U3293 ( .A(b[3]), .Z(n2209) );
  IV U3294 ( .A(b[3]), .Z(n2210) );
  IV U3295 ( .A(b[3]), .Z(n2211) );
  IV U3296 ( .A(b[3]), .Z(n2212) );
  IV U3297 ( .A(b[3]), .Z(n2213) );
  IV U3298 ( .A(b[3]), .Z(n2214) );
  IV U3299 ( .A(b[3]), .Z(n2215) );
  IV U3300 ( .A(b[3]), .Z(n2216) );
  IV U3301 ( .A(b[3]), .Z(n2217) );
  IV U3302 ( .A(b[3]), .Z(n2218) );
  IV U3303 ( .A(b[3]), .Z(n2219) );
  IV U3304 ( .A(b[3]), .Z(n2220) );
  IV U3305 ( .A(b[3]), .Z(n2221) );
  IV U3306 ( .A(b[3]), .Z(n2222) );
  IV U3307 ( .A(b[3]), .Z(n2223) );
  IV U3308 ( .A(b[3]), .Z(n2224) );
  IV U3309 ( .A(b[3]), .Z(n2225) );
  IV U3310 ( .A(b[3]), .Z(n2226) );
  IV U3311 ( .A(b[3]), .Z(n2227) );
  IV U3312 ( .A(b[3]), .Z(n2228) );
  IV U3313 ( .A(b[3]), .Z(n2229) );
  IV U3314 ( .A(b[3]), .Z(n2230) );
  IV U3315 ( .A(b[3]), .Z(n2231) );
  IV U3316 ( .A(b[3]), .Z(n2232) );
  IV U3317 ( .A(b[3]), .Z(n2233) );
  IV U3318 ( .A(b[3]), .Z(n2234) );
  IV U3319 ( .A(b[3]), .Z(n2235) );
  IV U3320 ( .A(b[3]), .Z(n2236) );
  IV U3321 ( .A(b[3]), .Z(n2237) );
  IV U3322 ( .A(b[3]), .Z(n2238) );
  IV U3323 ( .A(b[3]), .Z(n2239) );
  IV U3324 ( .A(b[3]), .Z(n2240) );
  IV U3325 ( .A(b[3]), .Z(n2241) );
  IV U3326 ( .A(b[3]), .Z(n2242) );
  IV U3327 ( .A(b[3]), .Z(n2243) );
  IV U3328 ( .A(b[3]), .Z(n2244) );
  IV U3329 ( .A(b[3]), .Z(n2245) );
  IV U3330 ( .A(b[3]), .Z(n2246) );
  IV U3331 ( .A(b[3]), .Z(n2247) );
  IV U3332 ( .A(b[3]), .Z(n2248) );
  IV U3333 ( .A(b[3]), .Z(n2249) );
  IV U3334 ( .A(b[3]), .Z(n2250) );
  IV U3335 ( .A(b[3]), .Z(n2251) );
  IV U3336 ( .A(b[3]), .Z(n2252) );
  IV U3337 ( .A(b[3]), .Z(n2253) );
  IV U3338 ( .A(b[3]), .Z(n2254) );
  IV U3339 ( .A(b[3]), .Z(n2255) );
  IV U3340 ( .A(b[3]), .Z(n2256) );
  IV U3341 ( .A(b[3]), .Z(n2257) );
  IV U3342 ( .A(b[3]), .Z(n2258) );
  IV U3343 ( .A(b[3]), .Z(n2259) );
  IV U3344 ( .A(b[3]), .Z(n2260) );
  IV U3345 ( .A(b[3]), .Z(n2261) );
  IV U3346 ( .A(b[3]), .Z(n2262) );
  IV U3347 ( .A(b[3]), .Z(n2263) );
  IV U3348 ( .A(b[3]), .Z(n2264) );
  IV U3349 ( .A(b[3]), .Z(n2265) );
  IV U3350 ( .A(b[3]), .Z(n2266) );
  IV U3351 ( .A(b[3]), .Z(n2267) );
  IV U3352 ( .A(b[3]), .Z(n2268) );
  IV U3353 ( .A(b[3]), .Z(n2269) );
  IV U3354 ( .A(b[3]), .Z(n2270) );
  IV U3355 ( .A(b[3]), .Z(n2271) );
  IV U3356 ( .A(b[3]), .Z(n2272) );
  IV U3357 ( .A(b[3]), .Z(n2273) );
  IV U3358 ( .A(b[3]), .Z(n2274) );
  IV U3359 ( .A(b[3]), .Z(n2275) );
  IV U3360 ( .A(b[3]), .Z(n2276) );
  IV U3361 ( .A(b[3]), .Z(n2277) );
  IV U3362 ( .A(b[3]), .Z(n2278) );
  IV U3363 ( .A(b[3]), .Z(n2279) );
  IV U3364 ( .A(b[3]), .Z(n2280) );
  IV U3365 ( .A(b[3]), .Z(n2281) );
  IV U3366 ( .A(b[3]), .Z(n2282) );
  IV U3367 ( .A(b[3]), .Z(n2283) );
  IV U3368 ( .A(b[3]), .Z(n2284) );
  IV U3369 ( .A(b[3]), .Z(n2285) );
  IV U3370 ( .A(b[3]), .Z(n2286) );
  IV U3371 ( .A(b[3]), .Z(n2287) );
  IV U3372 ( .A(b[3]), .Z(n2288) );
  IV U3373 ( .A(b[3]), .Z(n2289) );
  IV U3374 ( .A(b[3]), .Z(n2290) );
  IV U3375 ( .A(b[3]), .Z(n2291) );
  IV U3376 ( .A(b[3]), .Z(n2292) );
  IV U3377 ( .A(b[3]), .Z(n2293) );
  IV U3378 ( .A(b[3]), .Z(n2294) );
  IV U3379 ( .A(b[3]), .Z(n2295) );
  IV U3380 ( .A(b[3]), .Z(n2296) );
  IV U3381 ( .A(b[3]), .Z(n2297) );
  IV U3382 ( .A(b[3]), .Z(n2298) );
  IV U3383 ( .A(b[3]), .Z(n2299) );
  IV U3384 ( .A(b[3]), .Z(n2300) );
  IV U3385 ( .A(b[3]), .Z(n2301) );
  IV U3386 ( .A(b[3]), .Z(n2302) );
  IV U3387 ( .A(b[3]), .Z(n2303) );
  IV U3388 ( .A(b[3]), .Z(n2304) );
  IV U3389 ( .A(b[3]), .Z(n2305) );
  IV U3390 ( .A(b[3]), .Z(n2306) );
  IV U3391 ( .A(b[3]), .Z(n2307) );
  IV U3392 ( .A(b[3]), .Z(n2308) );
  IV U3393 ( .A(b[3]), .Z(n2309) );
  IV U3394 ( .A(b[3]), .Z(n2310) );
  IV U3395 ( .A(b[3]), .Z(n2311) );
  IV U3396 ( .A(b[3]), .Z(n2312) );
  IV U3397 ( .A(b[3]), .Z(n2313) );
  IV U3398 ( .A(b[3]), .Z(n2314) );
  IV U3399 ( .A(b[3]), .Z(n2315) );
  IV U3400 ( .A(b[3]), .Z(n2316) );
  IV U3401 ( .A(b[3]), .Z(n2317) );
  IV U3402 ( .A(b[3]), .Z(n2318) );
  IV U3403 ( .A(b[3]), .Z(n2319) );
  IV U3404 ( .A(b[3]), .Z(n2320) );
  IV U3405 ( .A(b[3]), .Z(n2321) );
  AND U3406 ( .A(b[0]), .B(a[0]), .Z(n2323) );
  XOR U3407 ( .A(n2323), .B(sreg[1020]), .Z(c[1020]) );
  AND U3408 ( .A(b[0]), .B(a[1]), .Z(n2330) );
  NAND U3409 ( .A(b[1]), .B(a[0]), .Z(n2322) );
  XOR U3410 ( .A(n2330), .B(n2322), .Z(n2324) );
  XNOR U3411 ( .A(sreg[1021]), .B(n2324), .Z(n2326) );
  AND U3412 ( .A(n2323), .B(sreg[1020]), .Z(n2325) );
  XOR U3413 ( .A(n2326), .B(n2325), .Z(c[1021]) );
  NANDN U3414 ( .A(n2324), .B(sreg[1021]), .Z(n2328) );
  NAND U3415 ( .A(n2326), .B(n2325), .Z(n2327) );
  AND U3416 ( .A(n2328), .B(n2327), .Z(n2336) );
  XNOR U3417 ( .A(n2336), .B(sreg[1022]), .Z(n2338) );
  AND U3418 ( .A(b[2]), .B(a[0]), .Z(n2329) );
  XNOR U3419 ( .A(n2329), .B(n2175), .Z(n2332) );
  NANDN U3420 ( .A(a[0]), .B(n2330), .Z(n2331) );
  NAND U3421 ( .A(n2332), .B(n2331), .Z(n2351) );
  AND U3422 ( .A(a[2]), .B(b[0]), .Z(n2333) );
  XNOR U3423 ( .A(n2333), .B(n2175), .Z(n2335) );
  NANDN U3424 ( .A(b[0]), .B(a[1]), .Z(n2334) );
  NAND U3425 ( .A(n2335), .B(n2334), .Z(n2350) );
  XOR U3426 ( .A(n2351), .B(n2350), .Z(n2337) );
  XOR U3427 ( .A(n2338), .B(n2337), .Z(c[1022]) );
  NANDN U3428 ( .A(n2336), .B(sreg[1022]), .Z(n2340) );
  NAND U3429 ( .A(n2338), .B(n2337), .Z(n2339) );
  NAND U3430 ( .A(n2340), .B(n2339), .Z(n2368) );
  AND U3431 ( .A(a[3]), .B(b[0]), .Z(n2341) );
  XNOR U3432 ( .A(n2341), .B(n2175), .Z(n2343) );
  NANDN U3433 ( .A(b[0]), .B(a[2]), .Z(n2342) );
  NAND U3434 ( .A(n2343), .B(n2342), .Z(n2366) );
  XNOR U3435 ( .A(a[1]), .B(n2176), .Z(n2359) );
  AND U3436 ( .A(n2359), .B(n2173), .Z(n2347) );
  XOR U3437 ( .A(b[2]), .B(b[3]), .Z(n2344) );
  XOR U3438 ( .A(a[0]), .B(b[3]), .Z(n2345) );
  NAND U3439 ( .A(n2174), .B(n2345), .Z(n2346) );
  NANDN U3440 ( .A(n2347), .B(n2346), .Z(n2365) );
  XNOR U3441 ( .A(n2366), .B(n2365), .Z(n2353) );
  NAND U3442 ( .A(b[1]), .B(b[2]), .Z(n23720) );
  AND U3443 ( .A(n23720), .B(b[3]), .Z(n2349) );
  NAND U3444 ( .A(n2173), .B(a[0]), .Z(n2348) );
  NAND U3445 ( .A(n2349), .B(n2348), .Z(n2354) );
  XNOR U3446 ( .A(n2353), .B(n2354), .Z(n2355) );
  OR U3447 ( .A(n2351), .B(n2350), .Z(n2356) );
  XNOR U3448 ( .A(n2355), .B(n2356), .Z(n2367) );
  XNOR U3449 ( .A(n2367), .B(sreg[1023]), .Z(n2352) );
  XNOR U3450 ( .A(n2368), .B(n2352), .Z(c[1023]) );
  NANDN U3451 ( .A(n2354), .B(n2353), .Z(n2358) );
  NANDN U3452 ( .A(n2356), .B(n2355), .Z(n2357) );
  AND U3453 ( .A(n2358), .B(n2357), .Z(n2374) );
  XOR U3454 ( .A(a[2]), .B(n2176), .Z(n2378) );
  NANDN U3455 ( .A(n2378), .B(n2173), .Z(n2361) );
  NAND U3456 ( .A(n2174), .B(n2359), .Z(n2360) );
  AND U3457 ( .A(n2361), .B(n2360), .Z(n2385) );
  AND U3458 ( .A(a[4]), .B(b[0]), .Z(n2362) );
  XNOR U3459 ( .A(n2362), .B(n2175), .Z(n2364) );
  NANDN U3460 ( .A(b[0]), .B(a[3]), .Z(n2363) );
  NAND U3461 ( .A(n2364), .B(n2363), .Z(n2383) );
  AND U3462 ( .A(a[0]), .B(b[3]), .Z(n2382) );
  XNOR U3463 ( .A(n2383), .B(n2382), .Z(n2384) );
  XNOR U3464 ( .A(n2385), .B(n2384), .Z(n2372) );
  NANDN U3465 ( .A(n2366), .B(n2365), .Z(n2373) );
  XOR U3466 ( .A(n2372), .B(n2373), .Z(n2375) );
  XNOR U3467 ( .A(n2374), .B(n2375), .Z(n2371) );
  XNOR U3468 ( .A(n2370), .B(sreg[1024]), .Z(n2369) );
  XNOR U3469 ( .A(n2371), .B(n2369), .Z(c[1024]) );
  NANDN U3470 ( .A(n2373), .B(n2372), .Z(n2377) );
  OR U3471 ( .A(n2375), .B(n2374), .Z(n2376) );
  AND U3472 ( .A(n2377), .B(n2376), .Z(n2391) );
  XOR U3473 ( .A(a[3]), .B(n2176), .Z(n2394) );
  AND U3474 ( .A(a[1]), .B(b[3]), .Z(n2398) );
  AND U3475 ( .A(a[5]), .B(b[0]), .Z(n2379) );
  XNOR U3476 ( .A(n2379), .B(n2175), .Z(n2381) );
  NANDN U3477 ( .A(b[0]), .B(a[4]), .Z(n2380) );
  NAND U3478 ( .A(n2381), .B(n2380), .Z(n2399) );
  XOR U3479 ( .A(n2398), .B(n2399), .Z(n2401) );
  XOR U3480 ( .A(n2400), .B(n2401), .Z(n2389) );
  NANDN U3481 ( .A(n2383), .B(n2382), .Z(n2387) );
  NANDN U3482 ( .A(n2385), .B(n2384), .Z(n2386) );
  AND U3483 ( .A(n2387), .B(n2386), .Z(n2388) );
  XNOR U3484 ( .A(n2389), .B(n2388), .Z(n2390) );
  XOR U3485 ( .A(n2391), .B(n2390), .Z(n2404) );
  XNOR U3486 ( .A(n2404), .B(sreg[1025]), .Z(n2405) );
  XNOR U3487 ( .A(n2406), .B(n2405), .Z(c[1025]) );
  NANDN U3488 ( .A(n2389), .B(n2388), .Z(n2393) );
  NAND U3489 ( .A(n2391), .B(n2390), .Z(n2392) );
  AND U3490 ( .A(n2393), .B(n2392), .Z(n2411) );
  XOR U3491 ( .A(a[4]), .B(n2176), .Z(n2415) );
  AND U3492 ( .A(a[6]), .B(b[0]), .Z(n2395) );
  XNOR U3493 ( .A(n2395), .B(n2175), .Z(n2397) );
  NANDN U3494 ( .A(b[0]), .B(a[5]), .Z(n2396) );
  NAND U3495 ( .A(n2397), .B(n2396), .Z(n2420) );
  AND U3496 ( .A(a[2]), .B(b[3]), .Z(n2419) );
  XOR U3497 ( .A(n2420), .B(n2419), .Z(n2422) );
  XOR U3498 ( .A(n2421), .B(n2422), .Z(n2410) );
  NANDN U3499 ( .A(n2399), .B(n2398), .Z(n2403) );
  OR U3500 ( .A(n2401), .B(n2400), .Z(n2402) );
  AND U3501 ( .A(n2403), .B(n2402), .Z(n2409) );
  XOR U3502 ( .A(n2410), .B(n2409), .Z(n2412) );
  XOR U3503 ( .A(n2411), .B(n2412), .Z(n2425) );
  XNOR U3504 ( .A(n2425), .B(sreg[1026]), .Z(n2427) );
  NANDN U3505 ( .A(n2404), .B(sreg[1025]), .Z(n2408) );
  NANDN U3506 ( .A(n2406), .B(n2405), .Z(n2407) );
  NAND U3507 ( .A(n2408), .B(n2407), .Z(n2426) );
  XOR U3508 ( .A(n2427), .B(n2426), .Z(c[1026]) );
  NANDN U3509 ( .A(n2410), .B(n2409), .Z(n2414) );
  OR U3510 ( .A(n2412), .B(n2411), .Z(n2413) );
  AND U3511 ( .A(n2414), .B(n2413), .Z(n2432) );
  XOR U3512 ( .A(a[5]), .B(n2176), .Z(n2436) );
  AND U3513 ( .A(a[3]), .B(b[3]), .Z(n2440) );
  AND U3514 ( .A(a[7]), .B(b[0]), .Z(n2416) );
  XNOR U3515 ( .A(n2416), .B(n2175), .Z(n2418) );
  NANDN U3516 ( .A(b[0]), .B(a[6]), .Z(n2417) );
  NAND U3517 ( .A(n2418), .B(n2417), .Z(n2441) );
  XOR U3518 ( .A(n2440), .B(n2441), .Z(n2443) );
  XOR U3519 ( .A(n2442), .B(n2443), .Z(n2431) );
  NANDN U3520 ( .A(n2420), .B(n2419), .Z(n2424) );
  OR U3521 ( .A(n2422), .B(n2421), .Z(n2423) );
  AND U3522 ( .A(n2424), .B(n2423), .Z(n2430) );
  XOR U3523 ( .A(n2431), .B(n2430), .Z(n2433) );
  XOR U3524 ( .A(n2432), .B(n2433), .Z(n2446) );
  XNOR U3525 ( .A(n2446), .B(sreg[1027]), .Z(n2448) );
  NANDN U3526 ( .A(n2425), .B(sreg[1026]), .Z(n2429) );
  NAND U3527 ( .A(n2427), .B(n2426), .Z(n2428) );
  NAND U3528 ( .A(n2429), .B(n2428), .Z(n2447) );
  XOR U3529 ( .A(n2448), .B(n2447), .Z(c[1027]) );
  NANDN U3530 ( .A(n2431), .B(n2430), .Z(n2435) );
  OR U3531 ( .A(n2433), .B(n2432), .Z(n2434) );
  AND U3532 ( .A(n2435), .B(n2434), .Z(n2453) );
  XOR U3533 ( .A(a[6]), .B(n2177), .Z(n2457) );
  AND U3534 ( .A(a[8]), .B(b[0]), .Z(n2437) );
  XNOR U3535 ( .A(n2437), .B(n2175), .Z(n2439) );
  NANDN U3536 ( .A(b[0]), .B(a[7]), .Z(n2438) );
  NAND U3537 ( .A(n2439), .B(n2438), .Z(n2462) );
  AND U3538 ( .A(a[4]), .B(b[3]), .Z(n2461) );
  XOR U3539 ( .A(n2462), .B(n2461), .Z(n2464) );
  XOR U3540 ( .A(n2463), .B(n2464), .Z(n2452) );
  NANDN U3541 ( .A(n2441), .B(n2440), .Z(n2445) );
  OR U3542 ( .A(n2443), .B(n2442), .Z(n2444) );
  AND U3543 ( .A(n2445), .B(n2444), .Z(n2451) );
  XOR U3544 ( .A(n2452), .B(n2451), .Z(n2454) );
  XOR U3545 ( .A(n2453), .B(n2454), .Z(n2467) );
  XNOR U3546 ( .A(n2467), .B(sreg[1028]), .Z(n2469) );
  NANDN U3547 ( .A(n2446), .B(sreg[1027]), .Z(n2450) );
  NAND U3548 ( .A(n2448), .B(n2447), .Z(n2449) );
  NAND U3549 ( .A(n2450), .B(n2449), .Z(n2468) );
  XOR U3550 ( .A(n2469), .B(n2468), .Z(c[1028]) );
  NANDN U3551 ( .A(n2452), .B(n2451), .Z(n2456) );
  OR U3552 ( .A(n2454), .B(n2453), .Z(n2455) );
  AND U3553 ( .A(n2456), .B(n2455), .Z(n2474) );
  XOR U3554 ( .A(a[7]), .B(n2177), .Z(n2478) );
  AND U3555 ( .A(a[5]), .B(b[3]), .Z(n2482) );
  AND U3556 ( .A(a[9]), .B(b[0]), .Z(n2458) );
  XNOR U3557 ( .A(n2458), .B(n2175), .Z(n2460) );
  NANDN U3558 ( .A(b[0]), .B(a[8]), .Z(n2459) );
  NAND U3559 ( .A(n2460), .B(n2459), .Z(n2483) );
  XOR U3560 ( .A(n2482), .B(n2483), .Z(n2485) );
  XOR U3561 ( .A(n2484), .B(n2485), .Z(n2473) );
  NANDN U3562 ( .A(n2462), .B(n2461), .Z(n2466) );
  OR U3563 ( .A(n2464), .B(n2463), .Z(n2465) );
  AND U3564 ( .A(n2466), .B(n2465), .Z(n2472) );
  XOR U3565 ( .A(n2473), .B(n2472), .Z(n2475) );
  XOR U3566 ( .A(n2474), .B(n2475), .Z(n2488) );
  XNOR U3567 ( .A(n2488), .B(sreg[1029]), .Z(n2490) );
  NANDN U3568 ( .A(n2467), .B(sreg[1028]), .Z(n2471) );
  NAND U3569 ( .A(n2469), .B(n2468), .Z(n2470) );
  NAND U3570 ( .A(n2471), .B(n2470), .Z(n2489) );
  XOR U3571 ( .A(n2490), .B(n2489), .Z(c[1029]) );
  NANDN U3572 ( .A(n2473), .B(n2472), .Z(n2477) );
  OR U3573 ( .A(n2475), .B(n2474), .Z(n2476) );
  AND U3574 ( .A(n2477), .B(n2476), .Z(n2495) );
  XOR U3575 ( .A(a[8]), .B(n2177), .Z(n2499) );
  AND U3576 ( .A(a[6]), .B(b[3]), .Z(n2503) );
  AND U3577 ( .A(a[10]), .B(b[0]), .Z(n2479) );
  XNOR U3578 ( .A(n2479), .B(n2175), .Z(n2481) );
  NANDN U3579 ( .A(b[0]), .B(a[9]), .Z(n2480) );
  NAND U3580 ( .A(n2481), .B(n2480), .Z(n2504) );
  XOR U3581 ( .A(n2503), .B(n2504), .Z(n2506) );
  XOR U3582 ( .A(n2505), .B(n2506), .Z(n2494) );
  NANDN U3583 ( .A(n2483), .B(n2482), .Z(n2487) );
  OR U3584 ( .A(n2485), .B(n2484), .Z(n2486) );
  AND U3585 ( .A(n2487), .B(n2486), .Z(n2493) );
  XOR U3586 ( .A(n2494), .B(n2493), .Z(n2496) );
  XOR U3587 ( .A(n2495), .B(n2496), .Z(n2509) );
  XNOR U3588 ( .A(n2509), .B(sreg[1030]), .Z(n2511) );
  NANDN U3589 ( .A(n2488), .B(sreg[1029]), .Z(n2492) );
  NAND U3590 ( .A(n2490), .B(n2489), .Z(n2491) );
  NAND U3591 ( .A(n2492), .B(n2491), .Z(n2510) );
  XOR U3592 ( .A(n2511), .B(n2510), .Z(c[1030]) );
  NANDN U3593 ( .A(n2494), .B(n2493), .Z(n2498) );
  OR U3594 ( .A(n2496), .B(n2495), .Z(n2497) );
  AND U3595 ( .A(n2498), .B(n2497), .Z(n2516) );
  XOR U3596 ( .A(a[9]), .B(n2177), .Z(n2520) );
  AND U3597 ( .A(a[11]), .B(b[0]), .Z(n2500) );
  XNOR U3598 ( .A(n2500), .B(n2175), .Z(n2502) );
  NANDN U3599 ( .A(b[0]), .B(a[10]), .Z(n2501) );
  NAND U3600 ( .A(n2502), .B(n2501), .Z(n2525) );
  AND U3601 ( .A(a[7]), .B(b[3]), .Z(n2524) );
  XOR U3602 ( .A(n2525), .B(n2524), .Z(n2527) );
  XOR U3603 ( .A(n2526), .B(n2527), .Z(n2515) );
  NANDN U3604 ( .A(n2504), .B(n2503), .Z(n2508) );
  OR U3605 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U3606 ( .A(n2508), .B(n2507), .Z(n2514) );
  XOR U3607 ( .A(n2515), .B(n2514), .Z(n2517) );
  XOR U3608 ( .A(n2516), .B(n2517), .Z(n2530) );
  XNOR U3609 ( .A(n2530), .B(sreg[1031]), .Z(n2532) );
  NANDN U3610 ( .A(n2509), .B(sreg[1030]), .Z(n2513) );
  NAND U3611 ( .A(n2511), .B(n2510), .Z(n2512) );
  NAND U3612 ( .A(n2513), .B(n2512), .Z(n2531) );
  XOR U3613 ( .A(n2532), .B(n2531), .Z(c[1031]) );
  NANDN U3614 ( .A(n2515), .B(n2514), .Z(n2519) );
  OR U3615 ( .A(n2517), .B(n2516), .Z(n2518) );
  AND U3616 ( .A(n2519), .B(n2518), .Z(n2537) );
  XOR U3617 ( .A(a[10]), .B(n2177), .Z(n2541) );
  AND U3618 ( .A(a[12]), .B(b[0]), .Z(n2521) );
  XNOR U3619 ( .A(n2521), .B(n2175), .Z(n2523) );
  NANDN U3620 ( .A(b[0]), .B(a[11]), .Z(n2522) );
  NAND U3621 ( .A(n2523), .B(n2522), .Z(n2546) );
  AND U3622 ( .A(a[8]), .B(b[3]), .Z(n2545) );
  XOR U3623 ( .A(n2546), .B(n2545), .Z(n2548) );
  XOR U3624 ( .A(n2547), .B(n2548), .Z(n2536) );
  NANDN U3625 ( .A(n2525), .B(n2524), .Z(n2529) );
  OR U3626 ( .A(n2527), .B(n2526), .Z(n2528) );
  AND U3627 ( .A(n2529), .B(n2528), .Z(n2535) );
  XOR U3628 ( .A(n2536), .B(n2535), .Z(n2538) );
  XOR U3629 ( .A(n2537), .B(n2538), .Z(n2551) );
  XNOR U3630 ( .A(n2551), .B(sreg[1032]), .Z(n2553) );
  NANDN U3631 ( .A(n2530), .B(sreg[1031]), .Z(n2534) );
  NAND U3632 ( .A(n2532), .B(n2531), .Z(n2533) );
  NAND U3633 ( .A(n2534), .B(n2533), .Z(n2552) );
  XOR U3634 ( .A(n2553), .B(n2552), .Z(c[1032]) );
  NANDN U3635 ( .A(n2536), .B(n2535), .Z(n2540) );
  OR U3636 ( .A(n2538), .B(n2537), .Z(n2539) );
  AND U3637 ( .A(n2540), .B(n2539), .Z(n2558) );
  XOR U3638 ( .A(a[11]), .B(n2177), .Z(n2562) );
  AND U3639 ( .A(a[13]), .B(b[0]), .Z(n2542) );
  XNOR U3640 ( .A(n2542), .B(n2175), .Z(n2544) );
  NANDN U3641 ( .A(b[0]), .B(a[12]), .Z(n2543) );
  NAND U3642 ( .A(n2544), .B(n2543), .Z(n2567) );
  AND U3643 ( .A(a[9]), .B(b[3]), .Z(n2566) );
  XOR U3644 ( .A(n2567), .B(n2566), .Z(n2569) );
  XOR U3645 ( .A(n2568), .B(n2569), .Z(n2557) );
  NANDN U3646 ( .A(n2546), .B(n2545), .Z(n2550) );
  OR U3647 ( .A(n2548), .B(n2547), .Z(n2549) );
  AND U3648 ( .A(n2550), .B(n2549), .Z(n2556) );
  XOR U3649 ( .A(n2557), .B(n2556), .Z(n2559) );
  XOR U3650 ( .A(n2558), .B(n2559), .Z(n2572) );
  XNOR U3651 ( .A(n2572), .B(sreg[1033]), .Z(n2574) );
  NANDN U3652 ( .A(n2551), .B(sreg[1032]), .Z(n2555) );
  NAND U3653 ( .A(n2553), .B(n2552), .Z(n2554) );
  NAND U3654 ( .A(n2555), .B(n2554), .Z(n2573) );
  XOR U3655 ( .A(n2574), .B(n2573), .Z(c[1033]) );
  NANDN U3656 ( .A(n2557), .B(n2556), .Z(n2561) );
  OR U3657 ( .A(n2559), .B(n2558), .Z(n2560) );
  AND U3658 ( .A(n2561), .B(n2560), .Z(n2579) );
  XOR U3659 ( .A(a[12]), .B(n2177), .Z(n2583) );
  AND U3660 ( .A(a[10]), .B(b[3]), .Z(n2587) );
  AND U3661 ( .A(a[14]), .B(b[0]), .Z(n2563) );
  XNOR U3662 ( .A(n2563), .B(n2175), .Z(n2565) );
  NANDN U3663 ( .A(b[0]), .B(a[13]), .Z(n2564) );
  NAND U3664 ( .A(n2565), .B(n2564), .Z(n2588) );
  XOR U3665 ( .A(n2587), .B(n2588), .Z(n2590) );
  XOR U3666 ( .A(n2589), .B(n2590), .Z(n2578) );
  NANDN U3667 ( .A(n2567), .B(n2566), .Z(n2571) );
  OR U3668 ( .A(n2569), .B(n2568), .Z(n2570) );
  AND U3669 ( .A(n2571), .B(n2570), .Z(n2577) );
  XOR U3670 ( .A(n2578), .B(n2577), .Z(n2580) );
  XOR U3671 ( .A(n2579), .B(n2580), .Z(n2593) );
  XNOR U3672 ( .A(n2593), .B(sreg[1034]), .Z(n2595) );
  NANDN U3673 ( .A(n2572), .B(sreg[1033]), .Z(n2576) );
  NAND U3674 ( .A(n2574), .B(n2573), .Z(n2575) );
  NAND U3675 ( .A(n2576), .B(n2575), .Z(n2594) );
  XOR U3676 ( .A(n2595), .B(n2594), .Z(c[1034]) );
  NANDN U3677 ( .A(n2578), .B(n2577), .Z(n2582) );
  OR U3678 ( .A(n2580), .B(n2579), .Z(n2581) );
  AND U3679 ( .A(n2582), .B(n2581), .Z(n2600) );
  XOR U3680 ( .A(a[13]), .B(n2178), .Z(n2604) );
  AND U3681 ( .A(a[11]), .B(b[3]), .Z(n2608) );
  AND U3682 ( .A(a[15]), .B(b[0]), .Z(n2584) );
  XNOR U3683 ( .A(n2584), .B(n2175), .Z(n2586) );
  NANDN U3684 ( .A(b[0]), .B(a[14]), .Z(n2585) );
  NAND U3685 ( .A(n2586), .B(n2585), .Z(n2609) );
  XOR U3686 ( .A(n2608), .B(n2609), .Z(n2611) );
  XOR U3687 ( .A(n2610), .B(n2611), .Z(n2599) );
  NANDN U3688 ( .A(n2588), .B(n2587), .Z(n2592) );
  OR U3689 ( .A(n2590), .B(n2589), .Z(n2591) );
  AND U3690 ( .A(n2592), .B(n2591), .Z(n2598) );
  XOR U3691 ( .A(n2599), .B(n2598), .Z(n2601) );
  XOR U3692 ( .A(n2600), .B(n2601), .Z(n2614) );
  XNOR U3693 ( .A(n2614), .B(sreg[1035]), .Z(n2616) );
  NANDN U3694 ( .A(n2593), .B(sreg[1034]), .Z(n2597) );
  NAND U3695 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U3696 ( .A(n2597), .B(n2596), .Z(n2615) );
  XOR U3697 ( .A(n2616), .B(n2615), .Z(c[1035]) );
  NANDN U3698 ( .A(n2599), .B(n2598), .Z(n2603) );
  OR U3699 ( .A(n2601), .B(n2600), .Z(n2602) );
  AND U3700 ( .A(n2603), .B(n2602), .Z(n2621) );
  XOR U3701 ( .A(a[14]), .B(n2178), .Z(n2625) );
  AND U3702 ( .A(a[12]), .B(b[3]), .Z(n2629) );
  AND U3703 ( .A(a[16]), .B(b[0]), .Z(n2605) );
  XNOR U3704 ( .A(n2605), .B(n2175), .Z(n2607) );
  NANDN U3705 ( .A(b[0]), .B(a[15]), .Z(n2606) );
  NAND U3706 ( .A(n2607), .B(n2606), .Z(n2630) );
  XOR U3707 ( .A(n2629), .B(n2630), .Z(n2632) );
  XOR U3708 ( .A(n2631), .B(n2632), .Z(n2620) );
  NANDN U3709 ( .A(n2609), .B(n2608), .Z(n2613) );
  OR U3710 ( .A(n2611), .B(n2610), .Z(n2612) );
  AND U3711 ( .A(n2613), .B(n2612), .Z(n2619) );
  XOR U3712 ( .A(n2620), .B(n2619), .Z(n2622) );
  XOR U3713 ( .A(n2621), .B(n2622), .Z(n2635) );
  XNOR U3714 ( .A(n2635), .B(sreg[1036]), .Z(n2637) );
  NANDN U3715 ( .A(n2614), .B(sreg[1035]), .Z(n2618) );
  NAND U3716 ( .A(n2616), .B(n2615), .Z(n2617) );
  NAND U3717 ( .A(n2618), .B(n2617), .Z(n2636) );
  XOR U3718 ( .A(n2637), .B(n2636), .Z(c[1036]) );
  NANDN U3719 ( .A(n2620), .B(n2619), .Z(n2624) );
  OR U3720 ( .A(n2622), .B(n2621), .Z(n2623) );
  AND U3721 ( .A(n2624), .B(n2623), .Z(n2642) );
  XOR U3722 ( .A(a[15]), .B(n2178), .Z(n2646) );
  AND U3723 ( .A(a[17]), .B(b[0]), .Z(n2626) );
  XNOR U3724 ( .A(n2626), .B(n2175), .Z(n2628) );
  NANDN U3725 ( .A(b[0]), .B(a[16]), .Z(n2627) );
  NAND U3726 ( .A(n2628), .B(n2627), .Z(n2651) );
  AND U3727 ( .A(a[13]), .B(b[3]), .Z(n2650) );
  XOR U3728 ( .A(n2651), .B(n2650), .Z(n2653) );
  XOR U3729 ( .A(n2652), .B(n2653), .Z(n2641) );
  NANDN U3730 ( .A(n2630), .B(n2629), .Z(n2634) );
  OR U3731 ( .A(n2632), .B(n2631), .Z(n2633) );
  AND U3732 ( .A(n2634), .B(n2633), .Z(n2640) );
  XOR U3733 ( .A(n2641), .B(n2640), .Z(n2643) );
  XOR U3734 ( .A(n2642), .B(n2643), .Z(n2656) );
  XNOR U3735 ( .A(n2656), .B(sreg[1037]), .Z(n2658) );
  NANDN U3736 ( .A(n2635), .B(sreg[1036]), .Z(n2639) );
  NAND U3737 ( .A(n2637), .B(n2636), .Z(n2638) );
  NAND U3738 ( .A(n2639), .B(n2638), .Z(n2657) );
  XOR U3739 ( .A(n2658), .B(n2657), .Z(c[1037]) );
  NANDN U3740 ( .A(n2641), .B(n2640), .Z(n2645) );
  OR U3741 ( .A(n2643), .B(n2642), .Z(n2644) );
  AND U3742 ( .A(n2645), .B(n2644), .Z(n2663) );
  XOR U3743 ( .A(a[16]), .B(n2178), .Z(n2667) );
  AND U3744 ( .A(a[18]), .B(b[0]), .Z(n2647) );
  XNOR U3745 ( .A(n2647), .B(n2175), .Z(n2649) );
  NANDN U3746 ( .A(b[0]), .B(a[17]), .Z(n2648) );
  NAND U3747 ( .A(n2649), .B(n2648), .Z(n2672) );
  AND U3748 ( .A(a[14]), .B(b[3]), .Z(n2671) );
  XOR U3749 ( .A(n2672), .B(n2671), .Z(n2674) );
  XOR U3750 ( .A(n2673), .B(n2674), .Z(n2662) );
  NANDN U3751 ( .A(n2651), .B(n2650), .Z(n2655) );
  OR U3752 ( .A(n2653), .B(n2652), .Z(n2654) );
  AND U3753 ( .A(n2655), .B(n2654), .Z(n2661) );
  XOR U3754 ( .A(n2662), .B(n2661), .Z(n2664) );
  XOR U3755 ( .A(n2663), .B(n2664), .Z(n2677) );
  XNOR U3756 ( .A(n2677), .B(sreg[1038]), .Z(n2679) );
  NANDN U3757 ( .A(n2656), .B(sreg[1037]), .Z(n2660) );
  NAND U3758 ( .A(n2658), .B(n2657), .Z(n2659) );
  NAND U3759 ( .A(n2660), .B(n2659), .Z(n2678) );
  XOR U3760 ( .A(n2679), .B(n2678), .Z(c[1038]) );
  NANDN U3761 ( .A(n2662), .B(n2661), .Z(n2666) );
  OR U3762 ( .A(n2664), .B(n2663), .Z(n2665) );
  AND U3763 ( .A(n2666), .B(n2665), .Z(n2684) );
  XOR U3764 ( .A(a[17]), .B(n2178), .Z(n2688) );
  AND U3765 ( .A(a[15]), .B(b[3]), .Z(n2692) );
  AND U3766 ( .A(a[19]), .B(b[0]), .Z(n2668) );
  XNOR U3767 ( .A(n2668), .B(n2175), .Z(n2670) );
  NANDN U3768 ( .A(b[0]), .B(a[18]), .Z(n2669) );
  NAND U3769 ( .A(n2670), .B(n2669), .Z(n2693) );
  XOR U3770 ( .A(n2692), .B(n2693), .Z(n2695) );
  XOR U3771 ( .A(n2694), .B(n2695), .Z(n2683) );
  NANDN U3772 ( .A(n2672), .B(n2671), .Z(n2676) );
  OR U3773 ( .A(n2674), .B(n2673), .Z(n2675) );
  AND U3774 ( .A(n2676), .B(n2675), .Z(n2682) );
  XOR U3775 ( .A(n2683), .B(n2682), .Z(n2685) );
  XOR U3776 ( .A(n2684), .B(n2685), .Z(n2698) );
  XNOR U3777 ( .A(n2698), .B(sreg[1039]), .Z(n2700) );
  NANDN U3778 ( .A(n2677), .B(sreg[1038]), .Z(n2681) );
  NAND U3779 ( .A(n2679), .B(n2678), .Z(n2680) );
  NAND U3780 ( .A(n2681), .B(n2680), .Z(n2699) );
  XOR U3781 ( .A(n2700), .B(n2699), .Z(c[1039]) );
  NANDN U3782 ( .A(n2683), .B(n2682), .Z(n2687) );
  OR U3783 ( .A(n2685), .B(n2684), .Z(n2686) );
  AND U3784 ( .A(n2687), .B(n2686), .Z(n2705) );
  XOR U3785 ( .A(a[18]), .B(n2178), .Z(n2709) );
  AND U3786 ( .A(a[20]), .B(b[0]), .Z(n2689) );
  XNOR U3787 ( .A(n2689), .B(n2175), .Z(n2691) );
  NANDN U3788 ( .A(b[0]), .B(a[19]), .Z(n2690) );
  NAND U3789 ( .A(n2691), .B(n2690), .Z(n2714) );
  AND U3790 ( .A(a[16]), .B(b[3]), .Z(n2713) );
  XOR U3791 ( .A(n2714), .B(n2713), .Z(n2716) );
  XOR U3792 ( .A(n2715), .B(n2716), .Z(n2704) );
  NANDN U3793 ( .A(n2693), .B(n2692), .Z(n2697) );
  OR U3794 ( .A(n2695), .B(n2694), .Z(n2696) );
  AND U3795 ( .A(n2697), .B(n2696), .Z(n2703) );
  XOR U3796 ( .A(n2704), .B(n2703), .Z(n2706) );
  XOR U3797 ( .A(n2705), .B(n2706), .Z(n2719) );
  XNOR U3798 ( .A(n2719), .B(sreg[1040]), .Z(n2721) );
  NANDN U3799 ( .A(n2698), .B(sreg[1039]), .Z(n2702) );
  NAND U3800 ( .A(n2700), .B(n2699), .Z(n2701) );
  NAND U3801 ( .A(n2702), .B(n2701), .Z(n2720) );
  XOR U3802 ( .A(n2721), .B(n2720), .Z(c[1040]) );
  NANDN U3803 ( .A(n2704), .B(n2703), .Z(n2708) );
  OR U3804 ( .A(n2706), .B(n2705), .Z(n2707) );
  AND U3805 ( .A(n2708), .B(n2707), .Z(n2726) );
  XOR U3806 ( .A(a[19]), .B(n2178), .Z(n2730) );
  AND U3807 ( .A(a[21]), .B(b[0]), .Z(n2710) );
  XNOR U3808 ( .A(n2710), .B(n2175), .Z(n2712) );
  NANDN U3809 ( .A(b[0]), .B(a[20]), .Z(n2711) );
  NAND U3810 ( .A(n2712), .B(n2711), .Z(n2735) );
  AND U3811 ( .A(a[17]), .B(b[3]), .Z(n2734) );
  XOR U3812 ( .A(n2735), .B(n2734), .Z(n2737) );
  XOR U3813 ( .A(n2736), .B(n2737), .Z(n2725) );
  NANDN U3814 ( .A(n2714), .B(n2713), .Z(n2718) );
  OR U3815 ( .A(n2716), .B(n2715), .Z(n2717) );
  AND U3816 ( .A(n2718), .B(n2717), .Z(n2724) );
  XOR U3817 ( .A(n2725), .B(n2724), .Z(n2727) );
  XOR U3818 ( .A(n2726), .B(n2727), .Z(n2740) );
  XNOR U3819 ( .A(n2740), .B(sreg[1041]), .Z(n2742) );
  NANDN U3820 ( .A(n2719), .B(sreg[1040]), .Z(n2723) );
  NAND U3821 ( .A(n2721), .B(n2720), .Z(n2722) );
  NAND U3822 ( .A(n2723), .B(n2722), .Z(n2741) );
  XOR U3823 ( .A(n2742), .B(n2741), .Z(c[1041]) );
  NANDN U3824 ( .A(n2725), .B(n2724), .Z(n2729) );
  OR U3825 ( .A(n2727), .B(n2726), .Z(n2728) );
  AND U3826 ( .A(n2729), .B(n2728), .Z(n2747) );
  XOR U3827 ( .A(a[20]), .B(n2179), .Z(n2751) );
  AND U3828 ( .A(a[22]), .B(b[0]), .Z(n2731) );
  XNOR U3829 ( .A(n2731), .B(n2175), .Z(n2733) );
  NANDN U3830 ( .A(b[0]), .B(a[21]), .Z(n2732) );
  NAND U3831 ( .A(n2733), .B(n2732), .Z(n2756) );
  AND U3832 ( .A(a[18]), .B(b[3]), .Z(n2755) );
  XOR U3833 ( .A(n2756), .B(n2755), .Z(n2758) );
  XOR U3834 ( .A(n2757), .B(n2758), .Z(n2746) );
  NANDN U3835 ( .A(n2735), .B(n2734), .Z(n2739) );
  OR U3836 ( .A(n2737), .B(n2736), .Z(n2738) );
  AND U3837 ( .A(n2739), .B(n2738), .Z(n2745) );
  XOR U3838 ( .A(n2746), .B(n2745), .Z(n2748) );
  XOR U3839 ( .A(n2747), .B(n2748), .Z(n2761) );
  XNOR U3840 ( .A(n2761), .B(sreg[1042]), .Z(n2763) );
  NANDN U3841 ( .A(n2740), .B(sreg[1041]), .Z(n2744) );
  NAND U3842 ( .A(n2742), .B(n2741), .Z(n2743) );
  NAND U3843 ( .A(n2744), .B(n2743), .Z(n2762) );
  XOR U3844 ( .A(n2763), .B(n2762), .Z(c[1042]) );
  NANDN U3845 ( .A(n2746), .B(n2745), .Z(n2750) );
  OR U3846 ( .A(n2748), .B(n2747), .Z(n2749) );
  AND U3847 ( .A(n2750), .B(n2749), .Z(n2768) );
  XOR U3848 ( .A(a[21]), .B(n2179), .Z(n2772) );
  AND U3849 ( .A(a[23]), .B(b[0]), .Z(n2752) );
  XNOR U3850 ( .A(n2752), .B(n2175), .Z(n2754) );
  NANDN U3851 ( .A(b[0]), .B(a[22]), .Z(n2753) );
  NAND U3852 ( .A(n2754), .B(n2753), .Z(n2777) );
  AND U3853 ( .A(a[19]), .B(b[3]), .Z(n2776) );
  XOR U3854 ( .A(n2777), .B(n2776), .Z(n2779) );
  XOR U3855 ( .A(n2778), .B(n2779), .Z(n2767) );
  NANDN U3856 ( .A(n2756), .B(n2755), .Z(n2760) );
  OR U3857 ( .A(n2758), .B(n2757), .Z(n2759) );
  AND U3858 ( .A(n2760), .B(n2759), .Z(n2766) );
  XOR U3859 ( .A(n2767), .B(n2766), .Z(n2769) );
  XOR U3860 ( .A(n2768), .B(n2769), .Z(n2782) );
  XNOR U3861 ( .A(n2782), .B(sreg[1043]), .Z(n2784) );
  NANDN U3862 ( .A(n2761), .B(sreg[1042]), .Z(n2765) );
  NAND U3863 ( .A(n2763), .B(n2762), .Z(n2764) );
  NAND U3864 ( .A(n2765), .B(n2764), .Z(n2783) );
  XOR U3865 ( .A(n2784), .B(n2783), .Z(c[1043]) );
  NANDN U3866 ( .A(n2767), .B(n2766), .Z(n2771) );
  OR U3867 ( .A(n2769), .B(n2768), .Z(n2770) );
  AND U3868 ( .A(n2771), .B(n2770), .Z(n2789) );
  XOR U3869 ( .A(a[22]), .B(n2179), .Z(n2793) );
  AND U3870 ( .A(a[24]), .B(b[0]), .Z(n2773) );
  XNOR U3871 ( .A(n2773), .B(n2175), .Z(n2775) );
  NANDN U3872 ( .A(b[0]), .B(a[23]), .Z(n2774) );
  NAND U3873 ( .A(n2775), .B(n2774), .Z(n2798) );
  AND U3874 ( .A(a[20]), .B(b[3]), .Z(n2797) );
  XOR U3875 ( .A(n2798), .B(n2797), .Z(n2800) );
  XOR U3876 ( .A(n2799), .B(n2800), .Z(n2788) );
  NANDN U3877 ( .A(n2777), .B(n2776), .Z(n2781) );
  OR U3878 ( .A(n2779), .B(n2778), .Z(n2780) );
  AND U3879 ( .A(n2781), .B(n2780), .Z(n2787) );
  XOR U3880 ( .A(n2788), .B(n2787), .Z(n2790) );
  XOR U3881 ( .A(n2789), .B(n2790), .Z(n2803) );
  XNOR U3882 ( .A(n2803), .B(sreg[1044]), .Z(n2805) );
  NANDN U3883 ( .A(n2782), .B(sreg[1043]), .Z(n2786) );
  NAND U3884 ( .A(n2784), .B(n2783), .Z(n2785) );
  NAND U3885 ( .A(n2786), .B(n2785), .Z(n2804) );
  XOR U3886 ( .A(n2805), .B(n2804), .Z(c[1044]) );
  NANDN U3887 ( .A(n2788), .B(n2787), .Z(n2792) );
  OR U3888 ( .A(n2790), .B(n2789), .Z(n2791) );
  AND U3889 ( .A(n2792), .B(n2791), .Z(n2810) );
  XOR U3890 ( .A(a[23]), .B(n2179), .Z(n2814) );
  AND U3891 ( .A(a[21]), .B(b[3]), .Z(n2818) );
  AND U3892 ( .A(a[25]), .B(b[0]), .Z(n2794) );
  XNOR U3893 ( .A(n2794), .B(n2175), .Z(n2796) );
  NANDN U3894 ( .A(b[0]), .B(a[24]), .Z(n2795) );
  NAND U3895 ( .A(n2796), .B(n2795), .Z(n2819) );
  XOR U3896 ( .A(n2818), .B(n2819), .Z(n2821) );
  XOR U3897 ( .A(n2820), .B(n2821), .Z(n2809) );
  NANDN U3898 ( .A(n2798), .B(n2797), .Z(n2802) );
  OR U3899 ( .A(n2800), .B(n2799), .Z(n2801) );
  AND U3900 ( .A(n2802), .B(n2801), .Z(n2808) );
  XOR U3901 ( .A(n2809), .B(n2808), .Z(n2811) );
  XOR U3902 ( .A(n2810), .B(n2811), .Z(n2824) );
  XNOR U3903 ( .A(n2824), .B(sreg[1045]), .Z(n2826) );
  NANDN U3904 ( .A(n2803), .B(sreg[1044]), .Z(n2807) );
  NAND U3905 ( .A(n2805), .B(n2804), .Z(n2806) );
  NAND U3906 ( .A(n2807), .B(n2806), .Z(n2825) );
  XOR U3907 ( .A(n2826), .B(n2825), .Z(c[1045]) );
  NANDN U3908 ( .A(n2809), .B(n2808), .Z(n2813) );
  OR U3909 ( .A(n2811), .B(n2810), .Z(n2812) );
  AND U3910 ( .A(n2813), .B(n2812), .Z(n2831) );
  XOR U3911 ( .A(a[24]), .B(n2179), .Z(n2835) );
  AND U3912 ( .A(a[26]), .B(b[0]), .Z(n2815) );
  XNOR U3913 ( .A(n2815), .B(n2175), .Z(n2817) );
  NANDN U3914 ( .A(b[0]), .B(a[25]), .Z(n2816) );
  NAND U3915 ( .A(n2817), .B(n2816), .Z(n2840) );
  AND U3916 ( .A(a[22]), .B(b[3]), .Z(n2839) );
  XOR U3917 ( .A(n2840), .B(n2839), .Z(n2842) );
  XOR U3918 ( .A(n2841), .B(n2842), .Z(n2830) );
  NANDN U3919 ( .A(n2819), .B(n2818), .Z(n2823) );
  OR U3920 ( .A(n2821), .B(n2820), .Z(n2822) );
  AND U3921 ( .A(n2823), .B(n2822), .Z(n2829) );
  XOR U3922 ( .A(n2830), .B(n2829), .Z(n2832) );
  XOR U3923 ( .A(n2831), .B(n2832), .Z(n2845) );
  XNOR U3924 ( .A(n2845), .B(sreg[1046]), .Z(n2847) );
  NANDN U3925 ( .A(n2824), .B(sreg[1045]), .Z(n2828) );
  NAND U3926 ( .A(n2826), .B(n2825), .Z(n2827) );
  NAND U3927 ( .A(n2828), .B(n2827), .Z(n2846) );
  XOR U3928 ( .A(n2847), .B(n2846), .Z(c[1046]) );
  NANDN U3929 ( .A(n2830), .B(n2829), .Z(n2834) );
  OR U3930 ( .A(n2832), .B(n2831), .Z(n2833) );
  AND U3931 ( .A(n2834), .B(n2833), .Z(n2852) );
  XOR U3932 ( .A(a[25]), .B(n2179), .Z(n2856) );
  AND U3933 ( .A(a[27]), .B(b[0]), .Z(n2836) );
  XNOR U3934 ( .A(n2836), .B(n2175), .Z(n2838) );
  NANDN U3935 ( .A(b[0]), .B(a[26]), .Z(n2837) );
  NAND U3936 ( .A(n2838), .B(n2837), .Z(n2861) );
  AND U3937 ( .A(a[23]), .B(b[3]), .Z(n2860) );
  XOR U3938 ( .A(n2861), .B(n2860), .Z(n2863) );
  XOR U3939 ( .A(n2862), .B(n2863), .Z(n2851) );
  NANDN U3940 ( .A(n2840), .B(n2839), .Z(n2844) );
  OR U3941 ( .A(n2842), .B(n2841), .Z(n2843) );
  AND U3942 ( .A(n2844), .B(n2843), .Z(n2850) );
  XOR U3943 ( .A(n2851), .B(n2850), .Z(n2853) );
  XOR U3944 ( .A(n2852), .B(n2853), .Z(n2866) );
  XNOR U3945 ( .A(n2866), .B(sreg[1047]), .Z(n2868) );
  NANDN U3946 ( .A(n2845), .B(sreg[1046]), .Z(n2849) );
  NAND U3947 ( .A(n2847), .B(n2846), .Z(n2848) );
  NAND U3948 ( .A(n2849), .B(n2848), .Z(n2867) );
  XOR U3949 ( .A(n2868), .B(n2867), .Z(c[1047]) );
  NANDN U3950 ( .A(n2851), .B(n2850), .Z(n2855) );
  OR U3951 ( .A(n2853), .B(n2852), .Z(n2854) );
  AND U3952 ( .A(n2855), .B(n2854), .Z(n2873) );
  XOR U3953 ( .A(a[26]), .B(n2179), .Z(n2877) );
  AND U3954 ( .A(a[24]), .B(b[3]), .Z(n2881) );
  AND U3955 ( .A(a[28]), .B(b[0]), .Z(n2857) );
  XNOR U3956 ( .A(n2857), .B(n2175), .Z(n2859) );
  NANDN U3957 ( .A(b[0]), .B(a[27]), .Z(n2858) );
  NAND U3958 ( .A(n2859), .B(n2858), .Z(n2882) );
  XOR U3959 ( .A(n2881), .B(n2882), .Z(n2884) );
  XOR U3960 ( .A(n2883), .B(n2884), .Z(n2872) );
  NANDN U3961 ( .A(n2861), .B(n2860), .Z(n2865) );
  OR U3962 ( .A(n2863), .B(n2862), .Z(n2864) );
  AND U3963 ( .A(n2865), .B(n2864), .Z(n2871) );
  XOR U3964 ( .A(n2872), .B(n2871), .Z(n2874) );
  XOR U3965 ( .A(n2873), .B(n2874), .Z(n2887) );
  XNOR U3966 ( .A(n2887), .B(sreg[1048]), .Z(n2889) );
  NANDN U3967 ( .A(n2866), .B(sreg[1047]), .Z(n2870) );
  NAND U3968 ( .A(n2868), .B(n2867), .Z(n2869) );
  NAND U3969 ( .A(n2870), .B(n2869), .Z(n2888) );
  XOR U3970 ( .A(n2889), .B(n2888), .Z(c[1048]) );
  NANDN U3971 ( .A(n2872), .B(n2871), .Z(n2876) );
  OR U3972 ( .A(n2874), .B(n2873), .Z(n2875) );
  AND U3973 ( .A(n2876), .B(n2875), .Z(n2894) );
  XOR U3974 ( .A(a[27]), .B(n2180), .Z(n2898) );
  AND U3975 ( .A(a[29]), .B(b[0]), .Z(n2878) );
  XNOR U3976 ( .A(n2878), .B(n2175), .Z(n2880) );
  NANDN U3977 ( .A(b[0]), .B(a[28]), .Z(n2879) );
  NAND U3978 ( .A(n2880), .B(n2879), .Z(n2903) );
  AND U3979 ( .A(a[25]), .B(b[3]), .Z(n2902) );
  XOR U3980 ( .A(n2903), .B(n2902), .Z(n2905) );
  XOR U3981 ( .A(n2904), .B(n2905), .Z(n2893) );
  NANDN U3982 ( .A(n2882), .B(n2881), .Z(n2886) );
  OR U3983 ( .A(n2884), .B(n2883), .Z(n2885) );
  AND U3984 ( .A(n2886), .B(n2885), .Z(n2892) );
  XOR U3985 ( .A(n2893), .B(n2892), .Z(n2895) );
  XOR U3986 ( .A(n2894), .B(n2895), .Z(n2908) );
  XNOR U3987 ( .A(n2908), .B(sreg[1049]), .Z(n2910) );
  NANDN U3988 ( .A(n2887), .B(sreg[1048]), .Z(n2891) );
  NAND U3989 ( .A(n2889), .B(n2888), .Z(n2890) );
  NAND U3990 ( .A(n2891), .B(n2890), .Z(n2909) );
  XOR U3991 ( .A(n2910), .B(n2909), .Z(c[1049]) );
  NANDN U3992 ( .A(n2893), .B(n2892), .Z(n2897) );
  OR U3993 ( .A(n2895), .B(n2894), .Z(n2896) );
  AND U3994 ( .A(n2897), .B(n2896), .Z(n2915) );
  XOR U3995 ( .A(a[28]), .B(n2180), .Z(n2919) );
  AND U3996 ( .A(a[30]), .B(b[0]), .Z(n2899) );
  XNOR U3997 ( .A(n2899), .B(n2175), .Z(n2901) );
  NANDN U3998 ( .A(b[0]), .B(a[29]), .Z(n2900) );
  NAND U3999 ( .A(n2901), .B(n2900), .Z(n2924) );
  AND U4000 ( .A(a[26]), .B(b[3]), .Z(n2923) );
  XOR U4001 ( .A(n2924), .B(n2923), .Z(n2926) );
  XOR U4002 ( .A(n2925), .B(n2926), .Z(n2914) );
  NANDN U4003 ( .A(n2903), .B(n2902), .Z(n2907) );
  OR U4004 ( .A(n2905), .B(n2904), .Z(n2906) );
  AND U4005 ( .A(n2907), .B(n2906), .Z(n2913) );
  XOR U4006 ( .A(n2914), .B(n2913), .Z(n2916) );
  XOR U4007 ( .A(n2915), .B(n2916), .Z(n2929) );
  XNOR U4008 ( .A(n2929), .B(sreg[1050]), .Z(n2931) );
  NANDN U4009 ( .A(n2908), .B(sreg[1049]), .Z(n2912) );
  NAND U4010 ( .A(n2910), .B(n2909), .Z(n2911) );
  NAND U4011 ( .A(n2912), .B(n2911), .Z(n2930) );
  XOR U4012 ( .A(n2931), .B(n2930), .Z(c[1050]) );
  NANDN U4013 ( .A(n2914), .B(n2913), .Z(n2918) );
  OR U4014 ( .A(n2916), .B(n2915), .Z(n2917) );
  AND U4015 ( .A(n2918), .B(n2917), .Z(n2936) );
  XOR U4016 ( .A(a[29]), .B(n2180), .Z(n2940) );
  AND U4017 ( .A(a[27]), .B(b[3]), .Z(n2944) );
  AND U4018 ( .A(a[31]), .B(b[0]), .Z(n2920) );
  XNOR U4019 ( .A(n2920), .B(n2175), .Z(n2922) );
  NANDN U4020 ( .A(b[0]), .B(a[30]), .Z(n2921) );
  NAND U4021 ( .A(n2922), .B(n2921), .Z(n2945) );
  XOR U4022 ( .A(n2944), .B(n2945), .Z(n2947) );
  XOR U4023 ( .A(n2946), .B(n2947), .Z(n2935) );
  NANDN U4024 ( .A(n2924), .B(n2923), .Z(n2928) );
  OR U4025 ( .A(n2926), .B(n2925), .Z(n2927) );
  AND U4026 ( .A(n2928), .B(n2927), .Z(n2934) );
  XOR U4027 ( .A(n2935), .B(n2934), .Z(n2937) );
  XOR U4028 ( .A(n2936), .B(n2937), .Z(n2950) );
  XNOR U4029 ( .A(n2950), .B(sreg[1051]), .Z(n2952) );
  NANDN U4030 ( .A(n2929), .B(sreg[1050]), .Z(n2933) );
  NAND U4031 ( .A(n2931), .B(n2930), .Z(n2932) );
  NAND U4032 ( .A(n2933), .B(n2932), .Z(n2951) );
  XOR U4033 ( .A(n2952), .B(n2951), .Z(c[1051]) );
  NANDN U4034 ( .A(n2935), .B(n2934), .Z(n2939) );
  OR U4035 ( .A(n2937), .B(n2936), .Z(n2938) );
  AND U4036 ( .A(n2939), .B(n2938), .Z(n2957) );
  XOR U4037 ( .A(a[30]), .B(n2180), .Z(n2961) );
  AND U4038 ( .A(a[32]), .B(b[0]), .Z(n2941) );
  XNOR U4039 ( .A(n2941), .B(n2175), .Z(n2943) );
  NANDN U4040 ( .A(b[0]), .B(a[31]), .Z(n2942) );
  NAND U4041 ( .A(n2943), .B(n2942), .Z(n2966) );
  AND U4042 ( .A(a[28]), .B(b[3]), .Z(n2965) );
  XOR U4043 ( .A(n2966), .B(n2965), .Z(n2968) );
  XOR U4044 ( .A(n2967), .B(n2968), .Z(n2956) );
  NANDN U4045 ( .A(n2945), .B(n2944), .Z(n2949) );
  OR U4046 ( .A(n2947), .B(n2946), .Z(n2948) );
  AND U4047 ( .A(n2949), .B(n2948), .Z(n2955) );
  XOR U4048 ( .A(n2956), .B(n2955), .Z(n2958) );
  XOR U4049 ( .A(n2957), .B(n2958), .Z(n2971) );
  XNOR U4050 ( .A(n2971), .B(sreg[1052]), .Z(n2973) );
  NANDN U4051 ( .A(n2950), .B(sreg[1051]), .Z(n2954) );
  NAND U4052 ( .A(n2952), .B(n2951), .Z(n2953) );
  NAND U4053 ( .A(n2954), .B(n2953), .Z(n2972) );
  XOR U4054 ( .A(n2973), .B(n2972), .Z(c[1052]) );
  NANDN U4055 ( .A(n2956), .B(n2955), .Z(n2960) );
  OR U4056 ( .A(n2958), .B(n2957), .Z(n2959) );
  AND U4057 ( .A(n2960), .B(n2959), .Z(n2978) );
  XOR U4058 ( .A(a[31]), .B(n2180), .Z(n2982) );
  AND U4059 ( .A(a[29]), .B(b[3]), .Z(n2986) );
  AND U4060 ( .A(a[33]), .B(b[0]), .Z(n2962) );
  XNOR U4061 ( .A(n2962), .B(n2175), .Z(n2964) );
  NANDN U4062 ( .A(b[0]), .B(a[32]), .Z(n2963) );
  NAND U4063 ( .A(n2964), .B(n2963), .Z(n2987) );
  XOR U4064 ( .A(n2986), .B(n2987), .Z(n2989) );
  XOR U4065 ( .A(n2988), .B(n2989), .Z(n2977) );
  NANDN U4066 ( .A(n2966), .B(n2965), .Z(n2970) );
  OR U4067 ( .A(n2968), .B(n2967), .Z(n2969) );
  AND U4068 ( .A(n2970), .B(n2969), .Z(n2976) );
  XOR U4069 ( .A(n2977), .B(n2976), .Z(n2979) );
  XOR U4070 ( .A(n2978), .B(n2979), .Z(n2992) );
  XNOR U4071 ( .A(n2992), .B(sreg[1053]), .Z(n2994) );
  NANDN U4072 ( .A(n2971), .B(sreg[1052]), .Z(n2975) );
  NAND U4073 ( .A(n2973), .B(n2972), .Z(n2974) );
  NAND U4074 ( .A(n2975), .B(n2974), .Z(n2993) );
  XOR U4075 ( .A(n2994), .B(n2993), .Z(c[1053]) );
  NANDN U4076 ( .A(n2977), .B(n2976), .Z(n2981) );
  OR U4077 ( .A(n2979), .B(n2978), .Z(n2980) );
  AND U4078 ( .A(n2981), .B(n2980), .Z(n2999) );
  XOR U4079 ( .A(a[32]), .B(n2180), .Z(n3003) );
  AND U4080 ( .A(a[34]), .B(b[0]), .Z(n2983) );
  XNOR U4081 ( .A(n2983), .B(n2175), .Z(n2985) );
  NANDN U4082 ( .A(b[0]), .B(a[33]), .Z(n2984) );
  NAND U4083 ( .A(n2985), .B(n2984), .Z(n3008) );
  AND U4084 ( .A(a[30]), .B(b[3]), .Z(n3007) );
  XOR U4085 ( .A(n3008), .B(n3007), .Z(n3010) );
  XOR U4086 ( .A(n3009), .B(n3010), .Z(n2998) );
  NANDN U4087 ( .A(n2987), .B(n2986), .Z(n2991) );
  OR U4088 ( .A(n2989), .B(n2988), .Z(n2990) );
  AND U4089 ( .A(n2991), .B(n2990), .Z(n2997) );
  XOR U4090 ( .A(n2998), .B(n2997), .Z(n3000) );
  XOR U4091 ( .A(n2999), .B(n3000), .Z(n3013) );
  XNOR U4092 ( .A(n3013), .B(sreg[1054]), .Z(n3015) );
  NANDN U4093 ( .A(n2992), .B(sreg[1053]), .Z(n2996) );
  NAND U4094 ( .A(n2994), .B(n2993), .Z(n2995) );
  NAND U4095 ( .A(n2996), .B(n2995), .Z(n3014) );
  XOR U4096 ( .A(n3015), .B(n3014), .Z(c[1054]) );
  NANDN U4097 ( .A(n2998), .B(n2997), .Z(n3002) );
  OR U4098 ( .A(n3000), .B(n2999), .Z(n3001) );
  AND U4099 ( .A(n3002), .B(n3001), .Z(n3020) );
  XOR U4100 ( .A(a[33]), .B(n2180), .Z(n3024) );
  AND U4101 ( .A(a[31]), .B(b[3]), .Z(n3028) );
  AND U4102 ( .A(a[35]), .B(b[0]), .Z(n3004) );
  XNOR U4103 ( .A(n3004), .B(n2175), .Z(n3006) );
  NANDN U4104 ( .A(b[0]), .B(a[34]), .Z(n3005) );
  NAND U4105 ( .A(n3006), .B(n3005), .Z(n3029) );
  XOR U4106 ( .A(n3028), .B(n3029), .Z(n3031) );
  XOR U4107 ( .A(n3030), .B(n3031), .Z(n3019) );
  NANDN U4108 ( .A(n3008), .B(n3007), .Z(n3012) );
  OR U4109 ( .A(n3010), .B(n3009), .Z(n3011) );
  AND U4110 ( .A(n3012), .B(n3011), .Z(n3018) );
  XOR U4111 ( .A(n3019), .B(n3018), .Z(n3021) );
  XOR U4112 ( .A(n3020), .B(n3021), .Z(n3034) );
  XNOR U4113 ( .A(n3034), .B(sreg[1055]), .Z(n3036) );
  NANDN U4114 ( .A(n3013), .B(sreg[1054]), .Z(n3017) );
  NAND U4115 ( .A(n3015), .B(n3014), .Z(n3016) );
  NAND U4116 ( .A(n3017), .B(n3016), .Z(n3035) );
  XOR U4117 ( .A(n3036), .B(n3035), .Z(c[1055]) );
  NANDN U4118 ( .A(n3019), .B(n3018), .Z(n3023) );
  OR U4119 ( .A(n3021), .B(n3020), .Z(n3022) );
  AND U4120 ( .A(n3023), .B(n3022), .Z(n3041) );
  XOR U4121 ( .A(a[34]), .B(n2181), .Z(n3045) );
  AND U4122 ( .A(a[32]), .B(b[3]), .Z(n3049) );
  AND U4123 ( .A(a[36]), .B(b[0]), .Z(n3025) );
  XNOR U4124 ( .A(n3025), .B(n2175), .Z(n3027) );
  NANDN U4125 ( .A(b[0]), .B(a[35]), .Z(n3026) );
  NAND U4126 ( .A(n3027), .B(n3026), .Z(n3050) );
  XOR U4127 ( .A(n3049), .B(n3050), .Z(n3052) );
  XOR U4128 ( .A(n3051), .B(n3052), .Z(n3040) );
  NANDN U4129 ( .A(n3029), .B(n3028), .Z(n3033) );
  OR U4130 ( .A(n3031), .B(n3030), .Z(n3032) );
  AND U4131 ( .A(n3033), .B(n3032), .Z(n3039) );
  XOR U4132 ( .A(n3040), .B(n3039), .Z(n3042) );
  XOR U4133 ( .A(n3041), .B(n3042), .Z(n3055) );
  XNOR U4134 ( .A(n3055), .B(sreg[1056]), .Z(n3057) );
  NANDN U4135 ( .A(n3034), .B(sreg[1055]), .Z(n3038) );
  NAND U4136 ( .A(n3036), .B(n3035), .Z(n3037) );
  NAND U4137 ( .A(n3038), .B(n3037), .Z(n3056) );
  XOR U4138 ( .A(n3057), .B(n3056), .Z(c[1056]) );
  NANDN U4139 ( .A(n3040), .B(n3039), .Z(n3044) );
  OR U4140 ( .A(n3042), .B(n3041), .Z(n3043) );
  AND U4141 ( .A(n3044), .B(n3043), .Z(n3062) );
  XOR U4142 ( .A(a[35]), .B(n2181), .Z(n3066) );
  AND U4143 ( .A(a[33]), .B(b[3]), .Z(n3070) );
  AND U4144 ( .A(a[37]), .B(b[0]), .Z(n3046) );
  XNOR U4145 ( .A(n3046), .B(n2175), .Z(n3048) );
  NANDN U4146 ( .A(b[0]), .B(a[36]), .Z(n3047) );
  NAND U4147 ( .A(n3048), .B(n3047), .Z(n3071) );
  XOR U4148 ( .A(n3070), .B(n3071), .Z(n3073) );
  XOR U4149 ( .A(n3072), .B(n3073), .Z(n3061) );
  NANDN U4150 ( .A(n3050), .B(n3049), .Z(n3054) );
  OR U4151 ( .A(n3052), .B(n3051), .Z(n3053) );
  AND U4152 ( .A(n3054), .B(n3053), .Z(n3060) );
  XOR U4153 ( .A(n3061), .B(n3060), .Z(n3063) );
  XOR U4154 ( .A(n3062), .B(n3063), .Z(n3076) );
  XNOR U4155 ( .A(n3076), .B(sreg[1057]), .Z(n3078) );
  NANDN U4156 ( .A(n3055), .B(sreg[1056]), .Z(n3059) );
  NAND U4157 ( .A(n3057), .B(n3056), .Z(n3058) );
  NAND U4158 ( .A(n3059), .B(n3058), .Z(n3077) );
  XOR U4159 ( .A(n3078), .B(n3077), .Z(c[1057]) );
  NANDN U4160 ( .A(n3061), .B(n3060), .Z(n3065) );
  OR U4161 ( .A(n3063), .B(n3062), .Z(n3064) );
  AND U4162 ( .A(n3065), .B(n3064), .Z(n3083) );
  XOR U4163 ( .A(a[36]), .B(n2181), .Z(n3087) );
  AND U4164 ( .A(a[38]), .B(b[0]), .Z(n3067) );
  XNOR U4165 ( .A(n3067), .B(n2175), .Z(n3069) );
  NANDN U4166 ( .A(b[0]), .B(a[37]), .Z(n3068) );
  NAND U4167 ( .A(n3069), .B(n3068), .Z(n3092) );
  AND U4168 ( .A(a[34]), .B(b[3]), .Z(n3091) );
  XOR U4169 ( .A(n3092), .B(n3091), .Z(n3094) );
  XOR U4170 ( .A(n3093), .B(n3094), .Z(n3082) );
  NANDN U4171 ( .A(n3071), .B(n3070), .Z(n3075) );
  OR U4172 ( .A(n3073), .B(n3072), .Z(n3074) );
  AND U4173 ( .A(n3075), .B(n3074), .Z(n3081) );
  XOR U4174 ( .A(n3082), .B(n3081), .Z(n3084) );
  XOR U4175 ( .A(n3083), .B(n3084), .Z(n3097) );
  XNOR U4176 ( .A(n3097), .B(sreg[1058]), .Z(n3099) );
  NANDN U4177 ( .A(n3076), .B(sreg[1057]), .Z(n3080) );
  NAND U4178 ( .A(n3078), .B(n3077), .Z(n3079) );
  NAND U4179 ( .A(n3080), .B(n3079), .Z(n3098) );
  XOR U4180 ( .A(n3099), .B(n3098), .Z(c[1058]) );
  NANDN U4181 ( .A(n3082), .B(n3081), .Z(n3086) );
  OR U4182 ( .A(n3084), .B(n3083), .Z(n3085) );
  AND U4183 ( .A(n3086), .B(n3085), .Z(n3104) );
  XOR U4184 ( .A(a[37]), .B(n2181), .Z(n3108) );
  AND U4185 ( .A(a[35]), .B(b[3]), .Z(n3112) );
  AND U4186 ( .A(a[39]), .B(b[0]), .Z(n3088) );
  XNOR U4187 ( .A(n3088), .B(n2175), .Z(n3090) );
  NANDN U4188 ( .A(b[0]), .B(a[38]), .Z(n3089) );
  NAND U4189 ( .A(n3090), .B(n3089), .Z(n3113) );
  XOR U4190 ( .A(n3112), .B(n3113), .Z(n3115) );
  XOR U4191 ( .A(n3114), .B(n3115), .Z(n3103) );
  NANDN U4192 ( .A(n3092), .B(n3091), .Z(n3096) );
  OR U4193 ( .A(n3094), .B(n3093), .Z(n3095) );
  AND U4194 ( .A(n3096), .B(n3095), .Z(n3102) );
  XOR U4195 ( .A(n3103), .B(n3102), .Z(n3105) );
  XOR U4196 ( .A(n3104), .B(n3105), .Z(n3118) );
  XNOR U4197 ( .A(n3118), .B(sreg[1059]), .Z(n3120) );
  NANDN U4198 ( .A(n3097), .B(sreg[1058]), .Z(n3101) );
  NAND U4199 ( .A(n3099), .B(n3098), .Z(n3100) );
  NAND U4200 ( .A(n3101), .B(n3100), .Z(n3119) );
  XOR U4201 ( .A(n3120), .B(n3119), .Z(c[1059]) );
  NANDN U4202 ( .A(n3103), .B(n3102), .Z(n3107) );
  OR U4203 ( .A(n3105), .B(n3104), .Z(n3106) );
  AND U4204 ( .A(n3107), .B(n3106), .Z(n3125) );
  XOR U4205 ( .A(a[38]), .B(n2181), .Z(n3129) );
  AND U4206 ( .A(a[40]), .B(b[0]), .Z(n3109) );
  XNOR U4207 ( .A(n3109), .B(n2175), .Z(n3111) );
  NANDN U4208 ( .A(b[0]), .B(a[39]), .Z(n3110) );
  NAND U4209 ( .A(n3111), .B(n3110), .Z(n3134) );
  AND U4210 ( .A(a[36]), .B(b[3]), .Z(n3133) );
  XOR U4211 ( .A(n3134), .B(n3133), .Z(n3136) );
  XOR U4212 ( .A(n3135), .B(n3136), .Z(n3124) );
  NANDN U4213 ( .A(n3113), .B(n3112), .Z(n3117) );
  OR U4214 ( .A(n3115), .B(n3114), .Z(n3116) );
  AND U4215 ( .A(n3117), .B(n3116), .Z(n3123) );
  XOR U4216 ( .A(n3124), .B(n3123), .Z(n3126) );
  XOR U4217 ( .A(n3125), .B(n3126), .Z(n3139) );
  XNOR U4218 ( .A(n3139), .B(sreg[1060]), .Z(n3141) );
  NANDN U4219 ( .A(n3118), .B(sreg[1059]), .Z(n3122) );
  NAND U4220 ( .A(n3120), .B(n3119), .Z(n3121) );
  NAND U4221 ( .A(n3122), .B(n3121), .Z(n3140) );
  XOR U4222 ( .A(n3141), .B(n3140), .Z(c[1060]) );
  NANDN U4223 ( .A(n3124), .B(n3123), .Z(n3128) );
  OR U4224 ( .A(n3126), .B(n3125), .Z(n3127) );
  AND U4225 ( .A(n3128), .B(n3127), .Z(n3146) );
  XOR U4226 ( .A(a[39]), .B(n2181), .Z(n3150) );
  AND U4227 ( .A(a[41]), .B(b[0]), .Z(n3130) );
  XNOR U4228 ( .A(n3130), .B(n2175), .Z(n3132) );
  NANDN U4229 ( .A(b[0]), .B(a[40]), .Z(n3131) );
  NAND U4230 ( .A(n3132), .B(n3131), .Z(n3155) );
  AND U4231 ( .A(a[37]), .B(b[3]), .Z(n3154) );
  XOR U4232 ( .A(n3155), .B(n3154), .Z(n3157) );
  XOR U4233 ( .A(n3156), .B(n3157), .Z(n3145) );
  NANDN U4234 ( .A(n3134), .B(n3133), .Z(n3138) );
  OR U4235 ( .A(n3136), .B(n3135), .Z(n3137) );
  AND U4236 ( .A(n3138), .B(n3137), .Z(n3144) );
  XOR U4237 ( .A(n3145), .B(n3144), .Z(n3147) );
  XOR U4238 ( .A(n3146), .B(n3147), .Z(n3160) );
  XNOR U4239 ( .A(n3160), .B(sreg[1061]), .Z(n3162) );
  NANDN U4240 ( .A(n3139), .B(sreg[1060]), .Z(n3143) );
  NAND U4241 ( .A(n3141), .B(n3140), .Z(n3142) );
  NAND U4242 ( .A(n3143), .B(n3142), .Z(n3161) );
  XOR U4243 ( .A(n3162), .B(n3161), .Z(c[1061]) );
  NANDN U4244 ( .A(n3145), .B(n3144), .Z(n3149) );
  OR U4245 ( .A(n3147), .B(n3146), .Z(n3148) );
  AND U4246 ( .A(n3149), .B(n3148), .Z(n3167) );
  XOR U4247 ( .A(a[40]), .B(n2181), .Z(n3171) );
  AND U4248 ( .A(a[42]), .B(b[0]), .Z(n3151) );
  XNOR U4249 ( .A(n3151), .B(n2175), .Z(n3153) );
  NANDN U4250 ( .A(b[0]), .B(a[41]), .Z(n3152) );
  NAND U4251 ( .A(n3153), .B(n3152), .Z(n3176) );
  AND U4252 ( .A(a[38]), .B(b[3]), .Z(n3175) );
  XOR U4253 ( .A(n3176), .B(n3175), .Z(n3178) );
  XOR U4254 ( .A(n3177), .B(n3178), .Z(n3166) );
  NANDN U4255 ( .A(n3155), .B(n3154), .Z(n3159) );
  OR U4256 ( .A(n3157), .B(n3156), .Z(n3158) );
  AND U4257 ( .A(n3159), .B(n3158), .Z(n3165) );
  XOR U4258 ( .A(n3166), .B(n3165), .Z(n3168) );
  XOR U4259 ( .A(n3167), .B(n3168), .Z(n3181) );
  XNOR U4260 ( .A(n3181), .B(sreg[1062]), .Z(n3183) );
  NANDN U4261 ( .A(n3160), .B(sreg[1061]), .Z(n3164) );
  NAND U4262 ( .A(n3162), .B(n3161), .Z(n3163) );
  NAND U4263 ( .A(n3164), .B(n3163), .Z(n3182) );
  XOR U4264 ( .A(n3183), .B(n3182), .Z(c[1062]) );
  NANDN U4265 ( .A(n3166), .B(n3165), .Z(n3170) );
  OR U4266 ( .A(n3168), .B(n3167), .Z(n3169) );
  AND U4267 ( .A(n3170), .B(n3169), .Z(n3188) );
  XOR U4268 ( .A(a[41]), .B(n2182), .Z(n3192) );
  AND U4269 ( .A(a[43]), .B(b[0]), .Z(n3172) );
  XNOR U4270 ( .A(n3172), .B(n2175), .Z(n3174) );
  NANDN U4271 ( .A(b[0]), .B(a[42]), .Z(n3173) );
  NAND U4272 ( .A(n3174), .B(n3173), .Z(n3197) );
  AND U4273 ( .A(a[39]), .B(b[3]), .Z(n3196) );
  XOR U4274 ( .A(n3197), .B(n3196), .Z(n3199) );
  XOR U4275 ( .A(n3198), .B(n3199), .Z(n3187) );
  NANDN U4276 ( .A(n3176), .B(n3175), .Z(n3180) );
  OR U4277 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U4278 ( .A(n3180), .B(n3179), .Z(n3186) );
  XOR U4279 ( .A(n3187), .B(n3186), .Z(n3189) );
  XOR U4280 ( .A(n3188), .B(n3189), .Z(n3202) );
  XNOR U4281 ( .A(n3202), .B(sreg[1063]), .Z(n3204) );
  NANDN U4282 ( .A(n3181), .B(sreg[1062]), .Z(n3185) );
  NAND U4283 ( .A(n3183), .B(n3182), .Z(n3184) );
  NAND U4284 ( .A(n3185), .B(n3184), .Z(n3203) );
  XOR U4285 ( .A(n3204), .B(n3203), .Z(c[1063]) );
  NANDN U4286 ( .A(n3187), .B(n3186), .Z(n3191) );
  OR U4287 ( .A(n3189), .B(n3188), .Z(n3190) );
  AND U4288 ( .A(n3191), .B(n3190), .Z(n3209) );
  XOR U4289 ( .A(a[42]), .B(n2182), .Z(n3213) );
  AND U4290 ( .A(a[40]), .B(b[3]), .Z(n3217) );
  AND U4291 ( .A(a[44]), .B(b[0]), .Z(n3193) );
  XNOR U4292 ( .A(n3193), .B(n2175), .Z(n3195) );
  NANDN U4293 ( .A(b[0]), .B(a[43]), .Z(n3194) );
  NAND U4294 ( .A(n3195), .B(n3194), .Z(n3218) );
  XOR U4295 ( .A(n3217), .B(n3218), .Z(n3220) );
  XOR U4296 ( .A(n3219), .B(n3220), .Z(n3208) );
  NANDN U4297 ( .A(n3197), .B(n3196), .Z(n3201) );
  OR U4298 ( .A(n3199), .B(n3198), .Z(n3200) );
  AND U4299 ( .A(n3201), .B(n3200), .Z(n3207) );
  XOR U4300 ( .A(n3208), .B(n3207), .Z(n3210) );
  XOR U4301 ( .A(n3209), .B(n3210), .Z(n3223) );
  XNOR U4302 ( .A(n3223), .B(sreg[1064]), .Z(n3225) );
  NANDN U4303 ( .A(n3202), .B(sreg[1063]), .Z(n3206) );
  NAND U4304 ( .A(n3204), .B(n3203), .Z(n3205) );
  NAND U4305 ( .A(n3206), .B(n3205), .Z(n3224) );
  XOR U4306 ( .A(n3225), .B(n3224), .Z(c[1064]) );
  NANDN U4307 ( .A(n3208), .B(n3207), .Z(n3212) );
  OR U4308 ( .A(n3210), .B(n3209), .Z(n3211) );
  AND U4309 ( .A(n3212), .B(n3211), .Z(n3230) );
  XOR U4310 ( .A(a[43]), .B(n2182), .Z(n3234) );
  AND U4311 ( .A(a[41]), .B(b[3]), .Z(n3238) );
  AND U4312 ( .A(a[45]), .B(b[0]), .Z(n3214) );
  XNOR U4313 ( .A(n3214), .B(n2175), .Z(n3216) );
  NANDN U4314 ( .A(b[0]), .B(a[44]), .Z(n3215) );
  NAND U4315 ( .A(n3216), .B(n3215), .Z(n3239) );
  XOR U4316 ( .A(n3238), .B(n3239), .Z(n3241) );
  XOR U4317 ( .A(n3240), .B(n3241), .Z(n3229) );
  NANDN U4318 ( .A(n3218), .B(n3217), .Z(n3222) );
  OR U4319 ( .A(n3220), .B(n3219), .Z(n3221) );
  AND U4320 ( .A(n3222), .B(n3221), .Z(n3228) );
  XOR U4321 ( .A(n3229), .B(n3228), .Z(n3231) );
  XOR U4322 ( .A(n3230), .B(n3231), .Z(n3244) );
  XNOR U4323 ( .A(n3244), .B(sreg[1065]), .Z(n3246) );
  NANDN U4324 ( .A(n3223), .B(sreg[1064]), .Z(n3227) );
  NAND U4325 ( .A(n3225), .B(n3224), .Z(n3226) );
  NAND U4326 ( .A(n3227), .B(n3226), .Z(n3245) );
  XOR U4327 ( .A(n3246), .B(n3245), .Z(c[1065]) );
  NANDN U4328 ( .A(n3229), .B(n3228), .Z(n3233) );
  OR U4329 ( .A(n3231), .B(n3230), .Z(n3232) );
  AND U4330 ( .A(n3233), .B(n3232), .Z(n3251) );
  XOR U4331 ( .A(a[44]), .B(n2182), .Z(n3255) );
  AND U4332 ( .A(a[42]), .B(b[3]), .Z(n3259) );
  AND U4333 ( .A(a[46]), .B(b[0]), .Z(n3235) );
  XNOR U4334 ( .A(n3235), .B(n2175), .Z(n3237) );
  NANDN U4335 ( .A(b[0]), .B(a[45]), .Z(n3236) );
  NAND U4336 ( .A(n3237), .B(n3236), .Z(n3260) );
  XOR U4337 ( .A(n3259), .B(n3260), .Z(n3262) );
  XOR U4338 ( .A(n3261), .B(n3262), .Z(n3250) );
  NANDN U4339 ( .A(n3239), .B(n3238), .Z(n3243) );
  OR U4340 ( .A(n3241), .B(n3240), .Z(n3242) );
  AND U4341 ( .A(n3243), .B(n3242), .Z(n3249) );
  XOR U4342 ( .A(n3250), .B(n3249), .Z(n3252) );
  XOR U4343 ( .A(n3251), .B(n3252), .Z(n3265) );
  XNOR U4344 ( .A(n3265), .B(sreg[1066]), .Z(n3267) );
  NANDN U4345 ( .A(n3244), .B(sreg[1065]), .Z(n3248) );
  NAND U4346 ( .A(n3246), .B(n3245), .Z(n3247) );
  NAND U4347 ( .A(n3248), .B(n3247), .Z(n3266) );
  XOR U4348 ( .A(n3267), .B(n3266), .Z(c[1066]) );
  NANDN U4349 ( .A(n3250), .B(n3249), .Z(n3254) );
  OR U4350 ( .A(n3252), .B(n3251), .Z(n3253) );
  AND U4351 ( .A(n3254), .B(n3253), .Z(n3272) );
  XOR U4352 ( .A(a[45]), .B(n2182), .Z(n3276) );
  AND U4353 ( .A(a[47]), .B(b[0]), .Z(n3256) );
  XNOR U4354 ( .A(n3256), .B(n2175), .Z(n3258) );
  NANDN U4355 ( .A(b[0]), .B(a[46]), .Z(n3257) );
  NAND U4356 ( .A(n3258), .B(n3257), .Z(n3281) );
  AND U4357 ( .A(a[43]), .B(b[3]), .Z(n3280) );
  XOR U4358 ( .A(n3281), .B(n3280), .Z(n3283) );
  XOR U4359 ( .A(n3282), .B(n3283), .Z(n3271) );
  NANDN U4360 ( .A(n3260), .B(n3259), .Z(n3264) );
  OR U4361 ( .A(n3262), .B(n3261), .Z(n3263) );
  AND U4362 ( .A(n3264), .B(n3263), .Z(n3270) );
  XOR U4363 ( .A(n3271), .B(n3270), .Z(n3273) );
  XOR U4364 ( .A(n3272), .B(n3273), .Z(n3286) );
  XNOR U4365 ( .A(n3286), .B(sreg[1067]), .Z(n3288) );
  NANDN U4366 ( .A(n3265), .B(sreg[1066]), .Z(n3269) );
  NAND U4367 ( .A(n3267), .B(n3266), .Z(n3268) );
  NAND U4368 ( .A(n3269), .B(n3268), .Z(n3287) );
  XOR U4369 ( .A(n3288), .B(n3287), .Z(c[1067]) );
  NANDN U4370 ( .A(n3271), .B(n3270), .Z(n3275) );
  OR U4371 ( .A(n3273), .B(n3272), .Z(n3274) );
  AND U4372 ( .A(n3275), .B(n3274), .Z(n3293) );
  XOR U4373 ( .A(a[46]), .B(n2182), .Z(n3297) );
  AND U4374 ( .A(a[48]), .B(b[0]), .Z(n3277) );
  XNOR U4375 ( .A(n3277), .B(n2175), .Z(n3279) );
  NANDN U4376 ( .A(b[0]), .B(a[47]), .Z(n3278) );
  NAND U4377 ( .A(n3279), .B(n3278), .Z(n3302) );
  AND U4378 ( .A(a[44]), .B(b[3]), .Z(n3301) );
  XOR U4379 ( .A(n3302), .B(n3301), .Z(n3304) );
  XOR U4380 ( .A(n3303), .B(n3304), .Z(n3292) );
  NANDN U4381 ( .A(n3281), .B(n3280), .Z(n3285) );
  OR U4382 ( .A(n3283), .B(n3282), .Z(n3284) );
  AND U4383 ( .A(n3285), .B(n3284), .Z(n3291) );
  XOR U4384 ( .A(n3292), .B(n3291), .Z(n3294) );
  XOR U4385 ( .A(n3293), .B(n3294), .Z(n3307) );
  XNOR U4386 ( .A(n3307), .B(sreg[1068]), .Z(n3309) );
  NANDN U4387 ( .A(n3286), .B(sreg[1067]), .Z(n3290) );
  NAND U4388 ( .A(n3288), .B(n3287), .Z(n3289) );
  NAND U4389 ( .A(n3290), .B(n3289), .Z(n3308) );
  XOR U4390 ( .A(n3309), .B(n3308), .Z(c[1068]) );
  NANDN U4391 ( .A(n3292), .B(n3291), .Z(n3296) );
  OR U4392 ( .A(n3294), .B(n3293), .Z(n3295) );
  AND U4393 ( .A(n3296), .B(n3295), .Z(n3314) );
  XOR U4394 ( .A(a[47]), .B(n2182), .Z(n3318) );
  AND U4395 ( .A(a[49]), .B(b[0]), .Z(n3298) );
  XNOR U4396 ( .A(n3298), .B(n2175), .Z(n3300) );
  NANDN U4397 ( .A(b[0]), .B(a[48]), .Z(n3299) );
  NAND U4398 ( .A(n3300), .B(n3299), .Z(n3323) );
  AND U4399 ( .A(a[45]), .B(b[3]), .Z(n3322) );
  XOR U4400 ( .A(n3323), .B(n3322), .Z(n3325) );
  XOR U4401 ( .A(n3324), .B(n3325), .Z(n3313) );
  NANDN U4402 ( .A(n3302), .B(n3301), .Z(n3306) );
  OR U4403 ( .A(n3304), .B(n3303), .Z(n3305) );
  AND U4404 ( .A(n3306), .B(n3305), .Z(n3312) );
  XOR U4405 ( .A(n3313), .B(n3312), .Z(n3315) );
  XOR U4406 ( .A(n3314), .B(n3315), .Z(n3328) );
  XNOR U4407 ( .A(n3328), .B(sreg[1069]), .Z(n3330) );
  NANDN U4408 ( .A(n3307), .B(sreg[1068]), .Z(n3311) );
  NAND U4409 ( .A(n3309), .B(n3308), .Z(n3310) );
  NAND U4410 ( .A(n3311), .B(n3310), .Z(n3329) );
  XOR U4411 ( .A(n3330), .B(n3329), .Z(c[1069]) );
  NANDN U4412 ( .A(n3313), .B(n3312), .Z(n3317) );
  OR U4413 ( .A(n3315), .B(n3314), .Z(n3316) );
  AND U4414 ( .A(n3317), .B(n3316), .Z(n3335) );
  XOR U4415 ( .A(a[48]), .B(n2183), .Z(n3339) );
  AND U4416 ( .A(a[50]), .B(b[0]), .Z(n3319) );
  XNOR U4417 ( .A(n3319), .B(n2175), .Z(n3321) );
  NANDN U4418 ( .A(b[0]), .B(a[49]), .Z(n3320) );
  NAND U4419 ( .A(n3321), .B(n3320), .Z(n3344) );
  AND U4420 ( .A(a[46]), .B(b[3]), .Z(n3343) );
  XOR U4421 ( .A(n3344), .B(n3343), .Z(n3346) );
  XOR U4422 ( .A(n3345), .B(n3346), .Z(n3334) );
  NANDN U4423 ( .A(n3323), .B(n3322), .Z(n3327) );
  OR U4424 ( .A(n3325), .B(n3324), .Z(n3326) );
  AND U4425 ( .A(n3327), .B(n3326), .Z(n3333) );
  XOR U4426 ( .A(n3334), .B(n3333), .Z(n3336) );
  XOR U4427 ( .A(n3335), .B(n3336), .Z(n3349) );
  XNOR U4428 ( .A(n3349), .B(sreg[1070]), .Z(n3351) );
  NANDN U4429 ( .A(n3328), .B(sreg[1069]), .Z(n3332) );
  NAND U4430 ( .A(n3330), .B(n3329), .Z(n3331) );
  NAND U4431 ( .A(n3332), .B(n3331), .Z(n3350) );
  XOR U4432 ( .A(n3351), .B(n3350), .Z(c[1070]) );
  NANDN U4433 ( .A(n3334), .B(n3333), .Z(n3338) );
  OR U4434 ( .A(n3336), .B(n3335), .Z(n3337) );
  AND U4435 ( .A(n3338), .B(n3337), .Z(n3356) );
  XOR U4436 ( .A(a[49]), .B(n2183), .Z(n3360) );
  AND U4437 ( .A(a[51]), .B(b[0]), .Z(n3340) );
  XNOR U4438 ( .A(n3340), .B(n2175), .Z(n3342) );
  NANDN U4439 ( .A(b[0]), .B(a[50]), .Z(n3341) );
  NAND U4440 ( .A(n3342), .B(n3341), .Z(n3365) );
  AND U4441 ( .A(a[47]), .B(b[3]), .Z(n3364) );
  XOR U4442 ( .A(n3365), .B(n3364), .Z(n3367) );
  XOR U4443 ( .A(n3366), .B(n3367), .Z(n3355) );
  NANDN U4444 ( .A(n3344), .B(n3343), .Z(n3348) );
  OR U4445 ( .A(n3346), .B(n3345), .Z(n3347) );
  AND U4446 ( .A(n3348), .B(n3347), .Z(n3354) );
  XOR U4447 ( .A(n3355), .B(n3354), .Z(n3357) );
  XOR U4448 ( .A(n3356), .B(n3357), .Z(n3370) );
  XNOR U4449 ( .A(n3370), .B(sreg[1071]), .Z(n3372) );
  NANDN U4450 ( .A(n3349), .B(sreg[1070]), .Z(n3353) );
  NAND U4451 ( .A(n3351), .B(n3350), .Z(n3352) );
  NAND U4452 ( .A(n3353), .B(n3352), .Z(n3371) );
  XOR U4453 ( .A(n3372), .B(n3371), .Z(c[1071]) );
  NANDN U4454 ( .A(n3355), .B(n3354), .Z(n3359) );
  OR U4455 ( .A(n3357), .B(n3356), .Z(n3358) );
  AND U4456 ( .A(n3359), .B(n3358), .Z(n3377) );
  XOR U4457 ( .A(a[50]), .B(n2183), .Z(n3381) );
  AND U4458 ( .A(a[52]), .B(b[0]), .Z(n3361) );
  XNOR U4459 ( .A(n3361), .B(n2175), .Z(n3363) );
  NANDN U4460 ( .A(b[0]), .B(a[51]), .Z(n3362) );
  NAND U4461 ( .A(n3363), .B(n3362), .Z(n3386) );
  AND U4462 ( .A(a[48]), .B(b[3]), .Z(n3385) );
  XOR U4463 ( .A(n3386), .B(n3385), .Z(n3388) );
  XOR U4464 ( .A(n3387), .B(n3388), .Z(n3376) );
  NANDN U4465 ( .A(n3365), .B(n3364), .Z(n3369) );
  OR U4466 ( .A(n3367), .B(n3366), .Z(n3368) );
  AND U4467 ( .A(n3369), .B(n3368), .Z(n3375) );
  XOR U4468 ( .A(n3376), .B(n3375), .Z(n3378) );
  XOR U4469 ( .A(n3377), .B(n3378), .Z(n3391) );
  XNOR U4470 ( .A(n3391), .B(sreg[1072]), .Z(n3393) );
  NANDN U4471 ( .A(n3370), .B(sreg[1071]), .Z(n3374) );
  NAND U4472 ( .A(n3372), .B(n3371), .Z(n3373) );
  NAND U4473 ( .A(n3374), .B(n3373), .Z(n3392) );
  XOR U4474 ( .A(n3393), .B(n3392), .Z(c[1072]) );
  NANDN U4475 ( .A(n3376), .B(n3375), .Z(n3380) );
  OR U4476 ( .A(n3378), .B(n3377), .Z(n3379) );
  AND U4477 ( .A(n3380), .B(n3379), .Z(n3398) );
  XOR U4478 ( .A(a[51]), .B(n2183), .Z(n3402) );
  AND U4479 ( .A(a[53]), .B(b[0]), .Z(n3382) );
  XNOR U4480 ( .A(n3382), .B(n2175), .Z(n3384) );
  NANDN U4481 ( .A(b[0]), .B(a[52]), .Z(n3383) );
  NAND U4482 ( .A(n3384), .B(n3383), .Z(n3407) );
  AND U4483 ( .A(a[49]), .B(b[3]), .Z(n3406) );
  XOR U4484 ( .A(n3407), .B(n3406), .Z(n3409) );
  XOR U4485 ( .A(n3408), .B(n3409), .Z(n3397) );
  NANDN U4486 ( .A(n3386), .B(n3385), .Z(n3390) );
  OR U4487 ( .A(n3388), .B(n3387), .Z(n3389) );
  AND U4488 ( .A(n3390), .B(n3389), .Z(n3396) );
  XOR U4489 ( .A(n3397), .B(n3396), .Z(n3399) );
  XOR U4490 ( .A(n3398), .B(n3399), .Z(n3412) );
  XNOR U4491 ( .A(n3412), .B(sreg[1073]), .Z(n3414) );
  NANDN U4492 ( .A(n3391), .B(sreg[1072]), .Z(n3395) );
  NAND U4493 ( .A(n3393), .B(n3392), .Z(n3394) );
  NAND U4494 ( .A(n3395), .B(n3394), .Z(n3413) );
  XOR U4495 ( .A(n3414), .B(n3413), .Z(c[1073]) );
  NANDN U4496 ( .A(n3397), .B(n3396), .Z(n3401) );
  OR U4497 ( .A(n3399), .B(n3398), .Z(n3400) );
  AND U4498 ( .A(n3401), .B(n3400), .Z(n3419) );
  XOR U4499 ( .A(a[52]), .B(n2183), .Z(n3423) );
  AND U4500 ( .A(a[54]), .B(b[0]), .Z(n3403) );
  XNOR U4501 ( .A(n3403), .B(n2175), .Z(n3405) );
  NANDN U4502 ( .A(b[0]), .B(a[53]), .Z(n3404) );
  NAND U4503 ( .A(n3405), .B(n3404), .Z(n3428) );
  AND U4504 ( .A(a[50]), .B(b[3]), .Z(n3427) );
  XOR U4505 ( .A(n3428), .B(n3427), .Z(n3430) );
  XOR U4506 ( .A(n3429), .B(n3430), .Z(n3418) );
  NANDN U4507 ( .A(n3407), .B(n3406), .Z(n3411) );
  OR U4508 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U4509 ( .A(n3411), .B(n3410), .Z(n3417) );
  XOR U4510 ( .A(n3418), .B(n3417), .Z(n3420) );
  XOR U4511 ( .A(n3419), .B(n3420), .Z(n3433) );
  XNOR U4512 ( .A(n3433), .B(sreg[1074]), .Z(n3435) );
  NANDN U4513 ( .A(n3412), .B(sreg[1073]), .Z(n3416) );
  NAND U4514 ( .A(n3414), .B(n3413), .Z(n3415) );
  NAND U4515 ( .A(n3416), .B(n3415), .Z(n3434) );
  XOR U4516 ( .A(n3435), .B(n3434), .Z(c[1074]) );
  NANDN U4517 ( .A(n3418), .B(n3417), .Z(n3422) );
  OR U4518 ( .A(n3420), .B(n3419), .Z(n3421) );
  AND U4519 ( .A(n3422), .B(n3421), .Z(n3440) );
  XOR U4520 ( .A(a[53]), .B(n2183), .Z(n3444) );
  AND U4521 ( .A(a[55]), .B(b[0]), .Z(n3424) );
  XNOR U4522 ( .A(n3424), .B(n2175), .Z(n3426) );
  NANDN U4523 ( .A(b[0]), .B(a[54]), .Z(n3425) );
  NAND U4524 ( .A(n3426), .B(n3425), .Z(n3449) );
  AND U4525 ( .A(a[51]), .B(b[3]), .Z(n3448) );
  XOR U4526 ( .A(n3449), .B(n3448), .Z(n3451) );
  XOR U4527 ( .A(n3450), .B(n3451), .Z(n3439) );
  NANDN U4528 ( .A(n3428), .B(n3427), .Z(n3432) );
  OR U4529 ( .A(n3430), .B(n3429), .Z(n3431) );
  AND U4530 ( .A(n3432), .B(n3431), .Z(n3438) );
  XOR U4531 ( .A(n3439), .B(n3438), .Z(n3441) );
  XOR U4532 ( .A(n3440), .B(n3441), .Z(n3454) );
  XNOR U4533 ( .A(n3454), .B(sreg[1075]), .Z(n3456) );
  NANDN U4534 ( .A(n3433), .B(sreg[1074]), .Z(n3437) );
  NAND U4535 ( .A(n3435), .B(n3434), .Z(n3436) );
  NAND U4536 ( .A(n3437), .B(n3436), .Z(n3455) );
  XOR U4537 ( .A(n3456), .B(n3455), .Z(c[1075]) );
  NANDN U4538 ( .A(n3439), .B(n3438), .Z(n3443) );
  OR U4539 ( .A(n3441), .B(n3440), .Z(n3442) );
  AND U4540 ( .A(n3443), .B(n3442), .Z(n3461) );
  XOR U4541 ( .A(a[54]), .B(n2183), .Z(n3465) );
  AND U4542 ( .A(a[52]), .B(b[3]), .Z(n3469) );
  AND U4543 ( .A(a[56]), .B(b[0]), .Z(n3445) );
  XNOR U4544 ( .A(n3445), .B(n2175), .Z(n3447) );
  NANDN U4545 ( .A(b[0]), .B(a[55]), .Z(n3446) );
  NAND U4546 ( .A(n3447), .B(n3446), .Z(n3470) );
  XOR U4547 ( .A(n3469), .B(n3470), .Z(n3472) );
  XOR U4548 ( .A(n3471), .B(n3472), .Z(n3460) );
  NANDN U4549 ( .A(n3449), .B(n3448), .Z(n3453) );
  OR U4550 ( .A(n3451), .B(n3450), .Z(n3452) );
  AND U4551 ( .A(n3453), .B(n3452), .Z(n3459) );
  XOR U4552 ( .A(n3460), .B(n3459), .Z(n3462) );
  XOR U4553 ( .A(n3461), .B(n3462), .Z(n3475) );
  XNOR U4554 ( .A(n3475), .B(sreg[1076]), .Z(n3477) );
  NANDN U4555 ( .A(n3454), .B(sreg[1075]), .Z(n3458) );
  NAND U4556 ( .A(n3456), .B(n3455), .Z(n3457) );
  NAND U4557 ( .A(n3458), .B(n3457), .Z(n3476) );
  XOR U4558 ( .A(n3477), .B(n3476), .Z(c[1076]) );
  NANDN U4559 ( .A(n3460), .B(n3459), .Z(n3464) );
  OR U4560 ( .A(n3462), .B(n3461), .Z(n3463) );
  AND U4561 ( .A(n3464), .B(n3463), .Z(n3482) );
  XOR U4562 ( .A(a[55]), .B(n2184), .Z(n3486) );
  AND U4563 ( .A(a[57]), .B(b[0]), .Z(n3466) );
  XNOR U4564 ( .A(n3466), .B(n2175), .Z(n3468) );
  NANDN U4565 ( .A(b[0]), .B(a[56]), .Z(n3467) );
  NAND U4566 ( .A(n3468), .B(n3467), .Z(n3491) );
  AND U4567 ( .A(a[53]), .B(b[3]), .Z(n3490) );
  XOR U4568 ( .A(n3491), .B(n3490), .Z(n3493) );
  XOR U4569 ( .A(n3492), .B(n3493), .Z(n3481) );
  NANDN U4570 ( .A(n3470), .B(n3469), .Z(n3474) );
  OR U4571 ( .A(n3472), .B(n3471), .Z(n3473) );
  AND U4572 ( .A(n3474), .B(n3473), .Z(n3480) );
  XOR U4573 ( .A(n3481), .B(n3480), .Z(n3483) );
  XOR U4574 ( .A(n3482), .B(n3483), .Z(n3496) );
  XNOR U4575 ( .A(n3496), .B(sreg[1077]), .Z(n3498) );
  NANDN U4576 ( .A(n3475), .B(sreg[1076]), .Z(n3479) );
  NAND U4577 ( .A(n3477), .B(n3476), .Z(n3478) );
  NAND U4578 ( .A(n3479), .B(n3478), .Z(n3497) );
  XOR U4579 ( .A(n3498), .B(n3497), .Z(c[1077]) );
  NANDN U4580 ( .A(n3481), .B(n3480), .Z(n3485) );
  OR U4581 ( .A(n3483), .B(n3482), .Z(n3484) );
  AND U4582 ( .A(n3485), .B(n3484), .Z(n3503) );
  XOR U4583 ( .A(a[56]), .B(n2184), .Z(n3507) );
  AND U4584 ( .A(a[54]), .B(b[3]), .Z(n3511) );
  AND U4585 ( .A(a[58]), .B(b[0]), .Z(n3487) );
  XNOR U4586 ( .A(n3487), .B(n2175), .Z(n3489) );
  NANDN U4587 ( .A(b[0]), .B(a[57]), .Z(n3488) );
  NAND U4588 ( .A(n3489), .B(n3488), .Z(n3512) );
  XOR U4589 ( .A(n3511), .B(n3512), .Z(n3514) );
  XOR U4590 ( .A(n3513), .B(n3514), .Z(n3502) );
  NANDN U4591 ( .A(n3491), .B(n3490), .Z(n3495) );
  OR U4592 ( .A(n3493), .B(n3492), .Z(n3494) );
  AND U4593 ( .A(n3495), .B(n3494), .Z(n3501) );
  XOR U4594 ( .A(n3502), .B(n3501), .Z(n3504) );
  XOR U4595 ( .A(n3503), .B(n3504), .Z(n3517) );
  XNOR U4596 ( .A(n3517), .B(sreg[1078]), .Z(n3519) );
  NANDN U4597 ( .A(n3496), .B(sreg[1077]), .Z(n3500) );
  NAND U4598 ( .A(n3498), .B(n3497), .Z(n3499) );
  NAND U4599 ( .A(n3500), .B(n3499), .Z(n3518) );
  XOR U4600 ( .A(n3519), .B(n3518), .Z(c[1078]) );
  NANDN U4601 ( .A(n3502), .B(n3501), .Z(n3506) );
  OR U4602 ( .A(n3504), .B(n3503), .Z(n3505) );
  AND U4603 ( .A(n3506), .B(n3505), .Z(n3524) );
  XOR U4604 ( .A(a[57]), .B(n2184), .Z(n3528) );
  AND U4605 ( .A(a[59]), .B(b[0]), .Z(n3508) );
  XNOR U4606 ( .A(n3508), .B(n2175), .Z(n3510) );
  NANDN U4607 ( .A(b[0]), .B(a[58]), .Z(n3509) );
  NAND U4608 ( .A(n3510), .B(n3509), .Z(n3533) );
  AND U4609 ( .A(a[55]), .B(b[3]), .Z(n3532) );
  XOR U4610 ( .A(n3533), .B(n3532), .Z(n3535) );
  XOR U4611 ( .A(n3534), .B(n3535), .Z(n3523) );
  NANDN U4612 ( .A(n3512), .B(n3511), .Z(n3516) );
  OR U4613 ( .A(n3514), .B(n3513), .Z(n3515) );
  AND U4614 ( .A(n3516), .B(n3515), .Z(n3522) );
  XOR U4615 ( .A(n3523), .B(n3522), .Z(n3525) );
  XOR U4616 ( .A(n3524), .B(n3525), .Z(n3538) );
  XNOR U4617 ( .A(n3538), .B(sreg[1079]), .Z(n3540) );
  NANDN U4618 ( .A(n3517), .B(sreg[1078]), .Z(n3521) );
  NAND U4619 ( .A(n3519), .B(n3518), .Z(n3520) );
  NAND U4620 ( .A(n3521), .B(n3520), .Z(n3539) );
  XOR U4621 ( .A(n3540), .B(n3539), .Z(c[1079]) );
  NANDN U4622 ( .A(n3523), .B(n3522), .Z(n3527) );
  OR U4623 ( .A(n3525), .B(n3524), .Z(n3526) );
  AND U4624 ( .A(n3527), .B(n3526), .Z(n3545) );
  XOR U4625 ( .A(a[58]), .B(n2184), .Z(n3549) );
  AND U4626 ( .A(a[60]), .B(b[0]), .Z(n3529) );
  XNOR U4627 ( .A(n3529), .B(n2175), .Z(n3531) );
  NANDN U4628 ( .A(b[0]), .B(a[59]), .Z(n3530) );
  NAND U4629 ( .A(n3531), .B(n3530), .Z(n3554) );
  AND U4630 ( .A(a[56]), .B(b[3]), .Z(n3553) );
  XOR U4631 ( .A(n3554), .B(n3553), .Z(n3556) );
  XOR U4632 ( .A(n3555), .B(n3556), .Z(n3544) );
  NANDN U4633 ( .A(n3533), .B(n3532), .Z(n3537) );
  OR U4634 ( .A(n3535), .B(n3534), .Z(n3536) );
  AND U4635 ( .A(n3537), .B(n3536), .Z(n3543) );
  XOR U4636 ( .A(n3544), .B(n3543), .Z(n3546) );
  XOR U4637 ( .A(n3545), .B(n3546), .Z(n3559) );
  XNOR U4638 ( .A(n3559), .B(sreg[1080]), .Z(n3561) );
  NANDN U4639 ( .A(n3538), .B(sreg[1079]), .Z(n3542) );
  NAND U4640 ( .A(n3540), .B(n3539), .Z(n3541) );
  NAND U4641 ( .A(n3542), .B(n3541), .Z(n3560) );
  XOR U4642 ( .A(n3561), .B(n3560), .Z(c[1080]) );
  NANDN U4643 ( .A(n3544), .B(n3543), .Z(n3548) );
  OR U4644 ( .A(n3546), .B(n3545), .Z(n3547) );
  AND U4645 ( .A(n3548), .B(n3547), .Z(n3566) );
  XOR U4646 ( .A(a[59]), .B(n2184), .Z(n3570) );
  AND U4647 ( .A(a[57]), .B(b[3]), .Z(n3574) );
  AND U4648 ( .A(a[61]), .B(b[0]), .Z(n3550) );
  XNOR U4649 ( .A(n3550), .B(n2175), .Z(n3552) );
  NANDN U4650 ( .A(b[0]), .B(a[60]), .Z(n3551) );
  NAND U4651 ( .A(n3552), .B(n3551), .Z(n3575) );
  XOR U4652 ( .A(n3574), .B(n3575), .Z(n3577) );
  XOR U4653 ( .A(n3576), .B(n3577), .Z(n3565) );
  NANDN U4654 ( .A(n3554), .B(n3553), .Z(n3558) );
  OR U4655 ( .A(n3556), .B(n3555), .Z(n3557) );
  AND U4656 ( .A(n3558), .B(n3557), .Z(n3564) );
  XOR U4657 ( .A(n3565), .B(n3564), .Z(n3567) );
  XOR U4658 ( .A(n3566), .B(n3567), .Z(n3580) );
  XNOR U4659 ( .A(n3580), .B(sreg[1081]), .Z(n3582) );
  NANDN U4660 ( .A(n3559), .B(sreg[1080]), .Z(n3563) );
  NAND U4661 ( .A(n3561), .B(n3560), .Z(n3562) );
  NAND U4662 ( .A(n3563), .B(n3562), .Z(n3581) );
  XOR U4663 ( .A(n3582), .B(n3581), .Z(c[1081]) );
  NANDN U4664 ( .A(n3565), .B(n3564), .Z(n3569) );
  OR U4665 ( .A(n3567), .B(n3566), .Z(n3568) );
  AND U4666 ( .A(n3569), .B(n3568), .Z(n3587) );
  XOR U4667 ( .A(a[60]), .B(n2184), .Z(n3591) );
  AND U4668 ( .A(a[58]), .B(b[3]), .Z(n3595) );
  AND U4669 ( .A(a[62]), .B(b[0]), .Z(n3571) );
  XNOR U4670 ( .A(n3571), .B(n2175), .Z(n3573) );
  NANDN U4671 ( .A(b[0]), .B(a[61]), .Z(n3572) );
  NAND U4672 ( .A(n3573), .B(n3572), .Z(n3596) );
  XOR U4673 ( .A(n3595), .B(n3596), .Z(n3598) );
  XOR U4674 ( .A(n3597), .B(n3598), .Z(n3586) );
  NANDN U4675 ( .A(n3575), .B(n3574), .Z(n3579) );
  OR U4676 ( .A(n3577), .B(n3576), .Z(n3578) );
  AND U4677 ( .A(n3579), .B(n3578), .Z(n3585) );
  XOR U4678 ( .A(n3586), .B(n3585), .Z(n3588) );
  XOR U4679 ( .A(n3587), .B(n3588), .Z(n3601) );
  XNOR U4680 ( .A(n3601), .B(sreg[1082]), .Z(n3603) );
  NANDN U4681 ( .A(n3580), .B(sreg[1081]), .Z(n3584) );
  NAND U4682 ( .A(n3582), .B(n3581), .Z(n3583) );
  NAND U4683 ( .A(n3584), .B(n3583), .Z(n3602) );
  XOR U4684 ( .A(n3603), .B(n3602), .Z(c[1082]) );
  NANDN U4685 ( .A(n3586), .B(n3585), .Z(n3590) );
  OR U4686 ( .A(n3588), .B(n3587), .Z(n3589) );
  AND U4687 ( .A(n3590), .B(n3589), .Z(n3608) );
  XOR U4688 ( .A(a[61]), .B(n2184), .Z(n3612) );
  AND U4689 ( .A(a[63]), .B(b[0]), .Z(n3592) );
  XNOR U4690 ( .A(n3592), .B(n2175), .Z(n3594) );
  NANDN U4691 ( .A(b[0]), .B(a[62]), .Z(n3593) );
  NAND U4692 ( .A(n3594), .B(n3593), .Z(n3617) );
  AND U4693 ( .A(a[59]), .B(b[3]), .Z(n3616) );
  XOR U4694 ( .A(n3617), .B(n3616), .Z(n3619) );
  XOR U4695 ( .A(n3618), .B(n3619), .Z(n3607) );
  NANDN U4696 ( .A(n3596), .B(n3595), .Z(n3600) );
  OR U4697 ( .A(n3598), .B(n3597), .Z(n3599) );
  AND U4698 ( .A(n3600), .B(n3599), .Z(n3606) );
  XOR U4699 ( .A(n3607), .B(n3606), .Z(n3609) );
  XOR U4700 ( .A(n3608), .B(n3609), .Z(n3622) );
  XNOR U4701 ( .A(n3622), .B(sreg[1083]), .Z(n3624) );
  NANDN U4702 ( .A(n3601), .B(sreg[1082]), .Z(n3605) );
  NAND U4703 ( .A(n3603), .B(n3602), .Z(n3604) );
  NAND U4704 ( .A(n3605), .B(n3604), .Z(n3623) );
  XOR U4705 ( .A(n3624), .B(n3623), .Z(c[1083]) );
  NANDN U4706 ( .A(n3607), .B(n3606), .Z(n3611) );
  OR U4707 ( .A(n3609), .B(n3608), .Z(n3610) );
  AND U4708 ( .A(n3611), .B(n3610), .Z(n3629) );
  XOR U4709 ( .A(a[62]), .B(n2185), .Z(n3633) );
  AND U4710 ( .A(a[64]), .B(b[0]), .Z(n3613) );
  XNOR U4711 ( .A(n3613), .B(n2175), .Z(n3615) );
  NANDN U4712 ( .A(b[0]), .B(a[63]), .Z(n3614) );
  NAND U4713 ( .A(n3615), .B(n3614), .Z(n3638) );
  AND U4714 ( .A(a[60]), .B(b[3]), .Z(n3637) );
  XOR U4715 ( .A(n3638), .B(n3637), .Z(n3640) );
  XOR U4716 ( .A(n3639), .B(n3640), .Z(n3628) );
  NANDN U4717 ( .A(n3617), .B(n3616), .Z(n3621) );
  OR U4718 ( .A(n3619), .B(n3618), .Z(n3620) );
  AND U4719 ( .A(n3621), .B(n3620), .Z(n3627) );
  XOR U4720 ( .A(n3628), .B(n3627), .Z(n3630) );
  XOR U4721 ( .A(n3629), .B(n3630), .Z(n3643) );
  XNOR U4722 ( .A(n3643), .B(sreg[1084]), .Z(n3645) );
  NANDN U4723 ( .A(n3622), .B(sreg[1083]), .Z(n3626) );
  NAND U4724 ( .A(n3624), .B(n3623), .Z(n3625) );
  NAND U4725 ( .A(n3626), .B(n3625), .Z(n3644) );
  XOR U4726 ( .A(n3645), .B(n3644), .Z(c[1084]) );
  NANDN U4727 ( .A(n3628), .B(n3627), .Z(n3632) );
  OR U4728 ( .A(n3630), .B(n3629), .Z(n3631) );
  AND U4729 ( .A(n3632), .B(n3631), .Z(n3650) );
  XOR U4730 ( .A(a[63]), .B(n2185), .Z(n3654) );
  AND U4731 ( .A(a[61]), .B(b[3]), .Z(n3658) );
  AND U4732 ( .A(a[65]), .B(b[0]), .Z(n3634) );
  XNOR U4733 ( .A(n3634), .B(n2175), .Z(n3636) );
  NANDN U4734 ( .A(b[0]), .B(a[64]), .Z(n3635) );
  NAND U4735 ( .A(n3636), .B(n3635), .Z(n3659) );
  XOR U4736 ( .A(n3658), .B(n3659), .Z(n3661) );
  XOR U4737 ( .A(n3660), .B(n3661), .Z(n3649) );
  NANDN U4738 ( .A(n3638), .B(n3637), .Z(n3642) );
  OR U4739 ( .A(n3640), .B(n3639), .Z(n3641) );
  AND U4740 ( .A(n3642), .B(n3641), .Z(n3648) );
  XOR U4741 ( .A(n3649), .B(n3648), .Z(n3651) );
  XOR U4742 ( .A(n3650), .B(n3651), .Z(n3664) );
  XNOR U4743 ( .A(n3664), .B(sreg[1085]), .Z(n3666) );
  NANDN U4744 ( .A(n3643), .B(sreg[1084]), .Z(n3647) );
  NAND U4745 ( .A(n3645), .B(n3644), .Z(n3646) );
  NAND U4746 ( .A(n3647), .B(n3646), .Z(n3665) );
  XOR U4747 ( .A(n3666), .B(n3665), .Z(c[1085]) );
  NANDN U4748 ( .A(n3649), .B(n3648), .Z(n3653) );
  OR U4749 ( .A(n3651), .B(n3650), .Z(n3652) );
  AND U4750 ( .A(n3653), .B(n3652), .Z(n3671) );
  XOR U4751 ( .A(a[64]), .B(n2185), .Z(n3675) );
  AND U4752 ( .A(a[66]), .B(b[0]), .Z(n3655) );
  XNOR U4753 ( .A(n3655), .B(n2175), .Z(n3657) );
  NANDN U4754 ( .A(b[0]), .B(a[65]), .Z(n3656) );
  NAND U4755 ( .A(n3657), .B(n3656), .Z(n3680) );
  AND U4756 ( .A(a[62]), .B(b[3]), .Z(n3679) );
  XOR U4757 ( .A(n3680), .B(n3679), .Z(n3682) );
  XOR U4758 ( .A(n3681), .B(n3682), .Z(n3670) );
  NANDN U4759 ( .A(n3659), .B(n3658), .Z(n3663) );
  OR U4760 ( .A(n3661), .B(n3660), .Z(n3662) );
  AND U4761 ( .A(n3663), .B(n3662), .Z(n3669) );
  XOR U4762 ( .A(n3670), .B(n3669), .Z(n3672) );
  XOR U4763 ( .A(n3671), .B(n3672), .Z(n3685) );
  XNOR U4764 ( .A(n3685), .B(sreg[1086]), .Z(n3687) );
  NANDN U4765 ( .A(n3664), .B(sreg[1085]), .Z(n3668) );
  NAND U4766 ( .A(n3666), .B(n3665), .Z(n3667) );
  NAND U4767 ( .A(n3668), .B(n3667), .Z(n3686) );
  XOR U4768 ( .A(n3687), .B(n3686), .Z(c[1086]) );
  NANDN U4769 ( .A(n3670), .B(n3669), .Z(n3674) );
  OR U4770 ( .A(n3672), .B(n3671), .Z(n3673) );
  AND U4771 ( .A(n3674), .B(n3673), .Z(n3692) );
  XOR U4772 ( .A(a[65]), .B(n2185), .Z(n3696) );
  AND U4773 ( .A(a[63]), .B(b[3]), .Z(n3700) );
  AND U4774 ( .A(a[67]), .B(b[0]), .Z(n3676) );
  XNOR U4775 ( .A(n3676), .B(n2175), .Z(n3678) );
  NANDN U4776 ( .A(b[0]), .B(a[66]), .Z(n3677) );
  NAND U4777 ( .A(n3678), .B(n3677), .Z(n3701) );
  XOR U4778 ( .A(n3700), .B(n3701), .Z(n3703) );
  XOR U4779 ( .A(n3702), .B(n3703), .Z(n3691) );
  NANDN U4780 ( .A(n3680), .B(n3679), .Z(n3684) );
  OR U4781 ( .A(n3682), .B(n3681), .Z(n3683) );
  AND U4782 ( .A(n3684), .B(n3683), .Z(n3690) );
  XOR U4783 ( .A(n3691), .B(n3690), .Z(n3693) );
  XOR U4784 ( .A(n3692), .B(n3693), .Z(n3706) );
  XNOR U4785 ( .A(n3706), .B(sreg[1087]), .Z(n3708) );
  NANDN U4786 ( .A(n3685), .B(sreg[1086]), .Z(n3689) );
  NAND U4787 ( .A(n3687), .B(n3686), .Z(n3688) );
  NAND U4788 ( .A(n3689), .B(n3688), .Z(n3707) );
  XOR U4789 ( .A(n3708), .B(n3707), .Z(c[1087]) );
  NANDN U4790 ( .A(n3691), .B(n3690), .Z(n3695) );
  OR U4791 ( .A(n3693), .B(n3692), .Z(n3694) );
  AND U4792 ( .A(n3695), .B(n3694), .Z(n3713) );
  XOR U4793 ( .A(a[66]), .B(n2185), .Z(n3717) );
  AND U4794 ( .A(a[68]), .B(b[0]), .Z(n3697) );
  XNOR U4795 ( .A(n3697), .B(n2175), .Z(n3699) );
  NANDN U4796 ( .A(b[0]), .B(a[67]), .Z(n3698) );
  NAND U4797 ( .A(n3699), .B(n3698), .Z(n3722) );
  AND U4798 ( .A(a[64]), .B(b[3]), .Z(n3721) );
  XOR U4799 ( .A(n3722), .B(n3721), .Z(n3724) );
  XOR U4800 ( .A(n3723), .B(n3724), .Z(n3712) );
  NANDN U4801 ( .A(n3701), .B(n3700), .Z(n3705) );
  OR U4802 ( .A(n3703), .B(n3702), .Z(n3704) );
  AND U4803 ( .A(n3705), .B(n3704), .Z(n3711) );
  XOR U4804 ( .A(n3712), .B(n3711), .Z(n3714) );
  XOR U4805 ( .A(n3713), .B(n3714), .Z(n3727) );
  XNOR U4806 ( .A(n3727), .B(sreg[1088]), .Z(n3729) );
  NANDN U4807 ( .A(n3706), .B(sreg[1087]), .Z(n3710) );
  NAND U4808 ( .A(n3708), .B(n3707), .Z(n3709) );
  NAND U4809 ( .A(n3710), .B(n3709), .Z(n3728) );
  XOR U4810 ( .A(n3729), .B(n3728), .Z(c[1088]) );
  NANDN U4811 ( .A(n3712), .B(n3711), .Z(n3716) );
  OR U4812 ( .A(n3714), .B(n3713), .Z(n3715) );
  AND U4813 ( .A(n3716), .B(n3715), .Z(n3734) );
  XOR U4814 ( .A(a[67]), .B(n2185), .Z(n3738) );
  AND U4815 ( .A(a[69]), .B(b[0]), .Z(n3718) );
  XNOR U4816 ( .A(n3718), .B(n2175), .Z(n3720) );
  NANDN U4817 ( .A(b[0]), .B(a[68]), .Z(n3719) );
  NAND U4818 ( .A(n3720), .B(n3719), .Z(n3743) );
  AND U4819 ( .A(a[65]), .B(b[3]), .Z(n3742) );
  XOR U4820 ( .A(n3743), .B(n3742), .Z(n3745) );
  XOR U4821 ( .A(n3744), .B(n3745), .Z(n3733) );
  NANDN U4822 ( .A(n3722), .B(n3721), .Z(n3726) );
  OR U4823 ( .A(n3724), .B(n3723), .Z(n3725) );
  AND U4824 ( .A(n3726), .B(n3725), .Z(n3732) );
  XOR U4825 ( .A(n3733), .B(n3732), .Z(n3735) );
  XOR U4826 ( .A(n3734), .B(n3735), .Z(n3748) );
  XNOR U4827 ( .A(n3748), .B(sreg[1089]), .Z(n3750) );
  NANDN U4828 ( .A(n3727), .B(sreg[1088]), .Z(n3731) );
  NAND U4829 ( .A(n3729), .B(n3728), .Z(n3730) );
  NAND U4830 ( .A(n3731), .B(n3730), .Z(n3749) );
  XOR U4831 ( .A(n3750), .B(n3749), .Z(c[1089]) );
  NANDN U4832 ( .A(n3733), .B(n3732), .Z(n3737) );
  OR U4833 ( .A(n3735), .B(n3734), .Z(n3736) );
  AND U4834 ( .A(n3737), .B(n3736), .Z(n3755) );
  XOR U4835 ( .A(a[68]), .B(n2185), .Z(n3759) );
  AND U4836 ( .A(a[66]), .B(b[3]), .Z(n3763) );
  AND U4837 ( .A(a[70]), .B(b[0]), .Z(n3739) );
  XNOR U4838 ( .A(n3739), .B(n2175), .Z(n3741) );
  NANDN U4839 ( .A(b[0]), .B(a[69]), .Z(n3740) );
  NAND U4840 ( .A(n3741), .B(n3740), .Z(n3764) );
  XOR U4841 ( .A(n3763), .B(n3764), .Z(n3766) );
  XOR U4842 ( .A(n3765), .B(n3766), .Z(n3754) );
  NANDN U4843 ( .A(n3743), .B(n3742), .Z(n3747) );
  OR U4844 ( .A(n3745), .B(n3744), .Z(n3746) );
  AND U4845 ( .A(n3747), .B(n3746), .Z(n3753) );
  XOR U4846 ( .A(n3754), .B(n3753), .Z(n3756) );
  XOR U4847 ( .A(n3755), .B(n3756), .Z(n3769) );
  XNOR U4848 ( .A(n3769), .B(sreg[1090]), .Z(n3771) );
  NANDN U4849 ( .A(n3748), .B(sreg[1089]), .Z(n3752) );
  NAND U4850 ( .A(n3750), .B(n3749), .Z(n3751) );
  NAND U4851 ( .A(n3752), .B(n3751), .Z(n3770) );
  XOR U4852 ( .A(n3771), .B(n3770), .Z(c[1090]) );
  NANDN U4853 ( .A(n3754), .B(n3753), .Z(n3758) );
  OR U4854 ( .A(n3756), .B(n3755), .Z(n3757) );
  AND U4855 ( .A(n3758), .B(n3757), .Z(n3776) );
  XOR U4856 ( .A(a[69]), .B(n2186), .Z(n3780) );
  AND U4857 ( .A(a[71]), .B(b[0]), .Z(n3760) );
  XNOR U4858 ( .A(n3760), .B(n2175), .Z(n3762) );
  NANDN U4859 ( .A(b[0]), .B(a[70]), .Z(n3761) );
  NAND U4860 ( .A(n3762), .B(n3761), .Z(n3785) );
  AND U4861 ( .A(a[67]), .B(b[3]), .Z(n3784) );
  XOR U4862 ( .A(n3785), .B(n3784), .Z(n3787) );
  XOR U4863 ( .A(n3786), .B(n3787), .Z(n3775) );
  NANDN U4864 ( .A(n3764), .B(n3763), .Z(n3768) );
  OR U4865 ( .A(n3766), .B(n3765), .Z(n3767) );
  AND U4866 ( .A(n3768), .B(n3767), .Z(n3774) );
  XOR U4867 ( .A(n3775), .B(n3774), .Z(n3777) );
  XOR U4868 ( .A(n3776), .B(n3777), .Z(n3790) );
  XNOR U4869 ( .A(n3790), .B(sreg[1091]), .Z(n3792) );
  NANDN U4870 ( .A(n3769), .B(sreg[1090]), .Z(n3773) );
  NAND U4871 ( .A(n3771), .B(n3770), .Z(n3772) );
  NAND U4872 ( .A(n3773), .B(n3772), .Z(n3791) );
  XOR U4873 ( .A(n3792), .B(n3791), .Z(c[1091]) );
  NANDN U4874 ( .A(n3775), .B(n3774), .Z(n3779) );
  OR U4875 ( .A(n3777), .B(n3776), .Z(n3778) );
  AND U4876 ( .A(n3779), .B(n3778), .Z(n3797) );
  XOR U4877 ( .A(a[70]), .B(n2186), .Z(n3801) );
  AND U4878 ( .A(a[72]), .B(b[0]), .Z(n3781) );
  XNOR U4879 ( .A(n3781), .B(n2175), .Z(n3783) );
  NANDN U4880 ( .A(b[0]), .B(a[71]), .Z(n3782) );
  NAND U4881 ( .A(n3783), .B(n3782), .Z(n3806) );
  AND U4882 ( .A(a[68]), .B(b[3]), .Z(n3805) );
  XOR U4883 ( .A(n3806), .B(n3805), .Z(n3808) );
  XOR U4884 ( .A(n3807), .B(n3808), .Z(n3796) );
  NANDN U4885 ( .A(n3785), .B(n3784), .Z(n3789) );
  OR U4886 ( .A(n3787), .B(n3786), .Z(n3788) );
  AND U4887 ( .A(n3789), .B(n3788), .Z(n3795) );
  XOR U4888 ( .A(n3796), .B(n3795), .Z(n3798) );
  XOR U4889 ( .A(n3797), .B(n3798), .Z(n3811) );
  XNOR U4890 ( .A(n3811), .B(sreg[1092]), .Z(n3813) );
  NANDN U4891 ( .A(n3790), .B(sreg[1091]), .Z(n3794) );
  NAND U4892 ( .A(n3792), .B(n3791), .Z(n3793) );
  NAND U4893 ( .A(n3794), .B(n3793), .Z(n3812) );
  XOR U4894 ( .A(n3813), .B(n3812), .Z(c[1092]) );
  NANDN U4895 ( .A(n3796), .B(n3795), .Z(n3800) );
  OR U4896 ( .A(n3798), .B(n3797), .Z(n3799) );
  AND U4897 ( .A(n3800), .B(n3799), .Z(n3818) );
  XOR U4898 ( .A(a[71]), .B(n2186), .Z(n3822) );
  AND U4899 ( .A(a[69]), .B(b[3]), .Z(n3826) );
  AND U4900 ( .A(a[73]), .B(b[0]), .Z(n3802) );
  XNOR U4901 ( .A(n3802), .B(n2175), .Z(n3804) );
  NANDN U4902 ( .A(b[0]), .B(a[72]), .Z(n3803) );
  NAND U4903 ( .A(n3804), .B(n3803), .Z(n3827) );
  XOR U4904 ( .A(n3826), .B(n3827), .Z(n3829) );
  XOR U4905 ( .A(n3828), .B(n3829), .Z(n3817) );
  NANDN U4906 ( .A(n3806), .B(n3805), .Z(n3810) );
  OR U4907 ( .A(n3808), .B(n3807), .Z(n3809) );
  AND U4908 ( .A(n3810), .B(n3809), .Z(n3816) );
  XOR U4909 ( .A(n3817), .B(n3816), .Z(n3819) );
  XOR U4910 ( .A(n3818), .B(n3819), .Z(n3832) );
  XNOR U4911 ( .A(n3832), .B(sreg[1093]), .Z(n3834) );
  NANDN U4912 ( .A(n3811), .B(sreg[1092]), .Z(n3815) );
  NAND U4913 ( .A(n3813), .B(n3812), .Z(n3814) );
  NAND U4914 ( .A(n3815), .B(n3814), .Z(n3833) );
  XOR U4915 ( .A(n3834), .B(n3833), .Z(c[1093]) );
  NANDN U4916 ( .A(n3817), .B(n3816), .Z(n3821) );
  OR U4917 ( .A(n3819), .B(n3818), .Z(n3820) );
  AND U4918 ( .A(n3821), .B(n3820), .Z(n3839) );
  XOR U4919 ( .A(a[72]), .B(n2186), .Z(n3843) );
  AND U4920 ( .A(a[74]), .B(b[0]), .Z(n3823) );
  XNOR U4921 ( .A(n3823), .B(n2175), .Z(n3825) );
  NANDN U4922 ( .A(b[0]), .B(a[73]), .Z(n3824) );
  NAND U4923 ( .A(n3825), .B(n3824), .Z(n3848) );
  AND U4924 ( .A(a[70]), .B(b[3]), .Z(n3847) );
  XOR U4925 ( .A(n3848), .B(n3847), .Z(n3850) );
  XOR U4926 ( .A(n3849), .B(n3850), .Z(n3838) );
  NANDN U4927 ( .A(n3827), .B(n3826), .Z(n3831) );
  OR U4928 ( .A(n3829), .B(n3828), .Z(n3830) );
  AND U4929 ( .A(n3831), .B(n3830), .Z(n3837) );
  XOR U4930 ( .A(n3838), .B(n3837), .Z(n3840) );
  XOR U4931 ( .A(n3839), .B(n3840), .Z(n3853) );
  XNOR U4932 ( .A(n3853), .B(sreg[1094]), .Z(n3855) );
  NANDN U4933 ( .A(n3832), .B(sreg[1093]), .Z(n3836) );
  NAND U4934 ( .A(n3834), .B(n3833), .Z(n3835) );
  NAND U4935 ( .A(n3836), .B(n3835), .Z(n3854) );
  XOR U4936 ( .A(n3855), .B(n3854), .Z(c[1094]) );
  NANDN U4937 ( .A(n3838), .B(n3837), .Z(n3842) );
  OR U4938 ( .A(n3840), .B(n3839), .Z(n3841) );
  AND U4939 ( .A(n3842), .B(n3841), .Z(n3860) );
  XOR U4940 ( .A(a[73]), .B(n2186), .Z(n3864) );
  AND U4941 ( .A(a[75]), .B(b[0]), .Z(n3844) );
  XNOR U4942 ( .A(n3844), .B(n2175), .Z(n3846) );
  NANDN U4943 ( .A(b[0]), .B(a[74]), .Z(n3845) );
  NAND U4944 ( .A(n3846), .B(n3845), .Z(n3869) );
  AND U4945 ( .A(a[71]), .B(b[3]), .Z(n3868) );
  XOR U4946 ( .A(n3869), .B(n3868), .Z(n3871) );
  XOR U4947 ( .A(n3870), .B(n3871), .Z(n3859) );
  NANDN U4948 ( .A(n3848), .B(n3847), .Z(n3852) );
  OR U4949 ( .A(n3850), .B(n3849), .Z(n3851) );
  AND U4950 ( .A(n3852), .B(n3851), .Z(n3858) );
  XOR U4951 ( .A(n3859), .B(n3858), .Z(n3861) );
  XOR U4952 ( .A(n3860), .B(n3861), .Z(n3874) );
  XNOR U4953 ( .A(n3874), .B(sreg[1095]), .Z(n3876) );
  NANDN U4954 ( .A(n3853), .B(sreg[1094]), .Z(n3857) );
  NAND U4955 ( .A(n3855), .B(n3854), .Z(n3856) );
  NAND U4956 ( .A(n3857), .B(n3856), .Z(n3875) );
  XOR U4957 ( .A(n3876), .B(n3875), .Z(c[1095]) );
  NANDN U4958 ( .A(n3859), .B(n3858), .Z(n3863) );
  OR U4959 ( .A(n3861), .B(n3860), .Z(n3862) );
  AND U4960 ( .A(n3863), .B(n3862), .Z(n3881) );
  XOR U4961 ( .A(a[74]), .B(n2186), .Z(n3885) );
  AND U4962 ( .A(a[72]), .B(b[3]), .Z(n3889) );
  AND U4963 ( .A(a[76]), .B(b[0]), .Z(n3865) );
  XNOR U4964 ( .A(n3865), .B(n2175), .Z(n3867) );
  NANDN U4965 ( .A(b[0]), .B(a[75]), .Z(n3866) );
  NAND U4966 ( .A(n3867), .B(n3866), .Z(n3890) );
  XOR U4967 ( .A(n3889), .B(n3890), .Z(n3892) );
  XOR U4968 ( .A(n3891), .B(n3892), .Z(n3880) );
  NANDN U4969 ( .A(n3869), .B(n3868), .Z(n3873) );
  OR U4970 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U4971 ( .A(n3873), .B(n3872), .Z(n3879) );
  XOR U4972 ( .A(n3880), .B(n3879), .Z(n3882) );
  XOR U4973 ( .A(n3881), .B(n3882), .Z(n3895) );
  XNOR U4974 ( .A(n3895), .B(sreg[1096]), .Z(n3897) );
  NANDN U4975 ( .A(n3874), .B(sreg[1095]), .Z(n3878) );
  NAND U4976 ( .A(n3876), .B(n3875), .Z(n3877) );
  NAND U4977 ( .A(n3878), .B(n3877), .Z(n3896) );
  XOR U4978 ( .A(n3897), .B(n3896), .Z(c[1096]) );
  NANDN U4979 ( .A(n3880), .B(n3879), .Z(n3884) );
  OR U4980 ( .A(n3882), .B(n3881), .Z(n3883) );
  AND U4981 ( .A(n3884), .B(n3883), .Z(n3902) );
  XOR U4982 ( .A(a[75]), .B(n2186), .Z(n3906) );
  AND U4983 ( .A(a[77]), .B(b[0]), .Z(n3886) );
  XNOR U4984 ( .A(n3886), .B(n2175), .Z(n3888) );
  NANDN U4985 ( .A(b[0]), .B(a[76]), .Z(n3887) );
  NAND U4986 ( .A(n3888), .B(n3887), .Z(n3911) );
  AND U4987 ( .A(a[73]), .B(b[3]), .Z(n3910) );
  XOR U4988 ( .A(n3911), .B(n3910), .Z(n3913) );
  XOR U4989 ( .A(n3912), .B(n3913), .Z(n3901) );
  NANDN U4990 ( .A(n3890), .B(n3889), .Z(n3894) );
  OR U4991 ( .A(n3892), .B(n3891), .Z(n3893) );
  AND U4992 ( .A(n3894), .B(n3893), .Z(n3900) );
  XOR U4993 ( .A(n3901), .B(n3900), .Z(n3903) );
  XOR U4994 ( .A(n3902), .B(n3903), .Z(n3916) );
  XNOR U4995 ( .A(n3916), .B(sreg[1097]), .Z(n3918) );
  NANDN U4996 ( .A(n3895), .B(sreg[1096]), .Z(n3899) );
  NAND U4997 ( .A(n3897), .B(n3896), .Z(n3898) );
  NAND U4998 ( .A(n3899), .B(n3898), .Z(n3917) );
  XOR U4999 ( .A(n3918), .B(n3917), .Z(c[1097]) );
  NANDN U5000 ( .A(n3901), .B(n3900), .Z(n3905) );
  OR U5001 ( .A(n3903), .B(n3902), .Z(n3904) );
  AND U5002 ( .A(n3905), .B(n3904), .Z(n3923) );
  XOR U5003 ( .A(a[76]), .B(n2187), .Z(n3927) );
  AND U5004 ( .A(a[78]), .B(b[0]), .Z(n3907) );
  XNOR U5005 ( .A(n3907), .B(n2175), .Z(n3909) );
  NANDN U5006 ( .A(b[0]), .B(a[77]), .Z(n3908) );
  NAND U5007 ( .A(n3909), .B(n3908), .Z(n3932) );
  AND U5008 ( .A(a[74]), .B(b[3]), .Z(n3931) );
  XOR U5009 ( .A(n3932), .B(n3931), .Z(n3934) );
  XOR U5010 ( .A(n3933), .B(n3934), .Z(n3922) );
  NANDN U5011 ( .A(n3911), .B(n3910), .Z(n3915) );
  OR U5012 ( .A(n3913), .B(n3912), .Z(n3914) );
  AND U5013 ( .A(n3915), .B(n3914), .Z(n3921) );
  XOR U5014 ( .A(n3922), .B(n3921), .Z(n3924) );
  XOR U5015 ( .A(n3923), .B(n3924), .Z(n3937) );
  XNOR U5016 ( .A(n3937), .B(sreg[1098]), .Z(n3939) );
  NANDN U5017 ( .A(n3916), .B(sreg[1097]), .Z(n3920) );
  NAND U5018 ( .A(n3918), .B(n3917), .Z(n3919) );
  NAND U5019 ( .A(n3920), .B(n3919), .Z(n3938) );
  XOR U5020 ( .A(n3939), .B(n3938), .Z(c[1098]) );
  NANDN U5021 ( .A(n3922), .B(n3921), .Z(n3926) );
  OR U5022 ( .A(n3924), .B(n3923), .Z(n3925) );
  AND U5023 ( .A(n3926), .B(n3925), .Z(n3944) );
  XOR U5024 ( .A(a[77]), .B(n2187), .Z(n3948) );
  AND U5025 ( .A(a[79]), .B(b[0]), .Z(n3928) );
  XNOR U5026 ( .A(n3928), .B(n2175), .Z(n3930) );
  NANDN U5027 ( .A(b[0]), .B(a[78]), .Z(n3929) );
  NAND U5028 ( .A(n3930), .B(n3929), .Z(n3953) );
  AND U5029 ( .A(a[75]), .B(b[3]), .Z(n3952) );
  XOR U5030 ( .A(n3953), .B(n3952), .Z(n3955) );
  XOR U5031 ( .A(n3954), .B(n3955), .Z(n3943) );
  NANDN U5032 ( .A(n3932), .B(n3931), .Z(n3936) );
  OR U5033 ( .A(n3934), .B(n3933), .Z(n3935) );
  AND U5034 ( .A(n3936), .B(n3935), .Z(n3942) );
  XOR U5035 ( .A(n3943), .B(n3942), .Z(n3945) );
  XOR U5036 ( .A(n3944), .B(n3945), .Z(n3958) );
  XNOR U5037 ( .A(n3958), .B(sreg[1099]), .Z(n3960) );
  NANDN U5038 ( .A(n3937), .B(sreg[1098]), .Z(n3941) );
  NAND U5039 ( .A(n3939), .B(n3938), .Z(n3940) );
  NAND U5040 ( .A(n3941), .B(n3940), .Z(n3959) );
  XOR U5041 ( .A(n3960), .B(n3959), .Z(c[1099]) );
  NANDN U5042 ( .A(n3943), .B(n3942), .Z(n3947) );
  OR U5043 ( .A(n3945), .B(n3944), .Z(n3946) );
  AND U5044 ( .A(n3947), .B(n3946), .Z(n3965) );
  XOR U5045 ( .A(a[78]), .B(n2187), .Z(n3969) );
  AND U5046 ( .A(a[76]), .B(b[3]), .Z(n3973) );
  AND U5047 ( .A(a[80]), .B(b[0]), .Z(n3949) );
  XNOR U5048 ( .A(n3949), .B(n2175), .Z(n3951) );
  NANDN U5049 ( .A(b[0]), .B(a[79]), .Z(n3950) );
  NAND U5050 ( .A(n3951), .B(n3950), .Z(n3974) );
  XOR U5051 ( .A(n3973), .B(n3974), .Z(n3976) );
  XOR U5052 ( .A(n3975), .B(n3976), .Z(n3964) );
  NANDN U5053 ( .A(n3953), .B(n3952), .Z(n3957) );
  OR U5054 ( .A(n3955), .B(n3954), .Z(n3956) );
  AND U5055 ( .A(n3957), .B(n3956), .Z(n3963) );
  XOR U5056 ( .A(n3964), .B(n3963), .Z(n3966) );
  XOR U5057 ( .A(n3965), .B(n3966), .Z(n3979) );
  XNOR U5058 ( .A(n3979), .B(sreg[1100]), .Z(n3981) );
  NANDN U5059 ( .A(n3958), .B(sreg[1099]), .Z(n3962) );
  NAND U5060 ( .A(n3960), .B(n3959), .Z(n3961) );
  NAND U5061 ( .A(n3962), .B(n3961), .Z(n3980) );
  XOR U5062 ( .A(n3981), .B(n3980), .Z(c[1100]) );
  NANDN U5063 ( .A(n3964), .B(n3963), .Z(n3968) );
  OR U5064 ( .A(n3966), .B(n3965), .Z(n3967) );
  AND U5065 ( .A(n3968), .B(n3967), .Z(n3986) );
  XOR U5066 ( .A(a[79]), .B(n2187), .Z(n3990) );
  AND U5067 ( .A(a[81]), .B(b[0]), .Z(n3970) );
  XNOR U5068 ( .A(n3970), .B(n2175), .Z(n3972) );
  NANDN U5069 ( .A(b[0]), .B(a[80]), .Z(n3971) );
  NAND U5070 ( .A(n3972), .B(n3971), .Z(n3995) );
  AND U5071 ( .A(a[77]), .B(b[3]), .Z(n3994) );
  XOR U5072 ( .A(n3995), .B(n3994), .Z(n3997) );
  XOR U5073 ( .A(n3996), .B(n3997), .Z(n3985) );
  NANDN U5074 ( .A(n3974), .B(n3973), .Z(n3978) );
  OR U5075 ( .A(n3976), .B(n3975), .Z(n3977) );
  AND U5076 ( .A(n3978), .B(n3977), .Z(n3984) );
  XOR U5077 ( .A(n3985), .B(n3984), .Z(n3987) );
  XOR U5078 ( .A(n3986), .B(n3987), .Z(n4000) );
  XNOR U5079 ( .A(n4000), .B(sreg[1101]), .Z(n4002) );
  NANDN U5080 ( .A(n3979), .B(sreg[1100]), .Z(n3983) );
  NAND U5081 ( .A(n3981), .B(n3980), .Z(n3982) );
  NAND U5082 ( .A(n3983), .B(n3982), .Z(n4001) );
  XOR U5083 ( .A(n4002), .B(n4001), .Z(c[1101]) );
  NANDN U5084 ( .A(n3985), .B(n3984), .Z(n3989) );
  OR U5085 ( .A(n3987), .B(n3986), .Z(n3988) );
  AND U5086 ( .A(n3989), .B(n3988), .Z(n4007) );
  XOR U5087 ( .A(a[80]), .B(n2187), .Z(n4011) );
  AND U5088 ( .A(a[82]), .B(b[0]), .Z(n3991) );
  XNOR U5089 ( .A(n3991), .B(n2175), .Z(n3993) );
  NANDN U5090 ( .A(b[0]), .B(a[81]), .Z(n3992) );
  NAND U5091 ( .A(n3993), .B(n3992), .Z(n4016) );
  AND U5092 ( .A(a[78]), .B(b[3]), .Z(n4015) );
  XOR U5093 ( .A(n4016), .B(n4015), .Z(n4018) );
  XOR U5094 ( .A(n4017), .B(n4018), .Z(n4006) );
  NANDN U5095 ( .A(n3995), .B(n3994), .Z(n3999) );
  OR U5096 ( .A(n3997), .B(n3996), .Z(n3998) );
  AND U5097 ( .A(n3999), .B(n3998), .Z(n4005) );
  XOR U5098 ( .A(n4006), .B(n4005), .Z(n4008) );
  XOR U5099 ( .A(n4007), .B(n4008), .Z(n4021) );
  XNOR U5100 ( .A(n4021), .B(sreg[1102]), .Z(n4023) );
  NANDN U5101 ( .A(n4000), .B(sreg[1101]), .Z(n4004) );
  NAND U5102 ( .A(n4002), .B(n4001), .Z(n4003) );
  NAND U5103 ( .A(n4004), .B(n4003), .Z(n4022) );
  XOR U5104 ( .A(n4023), .B(n4022), .Z(c[1102]) );
  NANDN U5105 ( .A(n4006), .B(n4005), .Z(n4010) );
  OR U5106 ( .A(n4008), .B(n4007), .Z(n4009) );
  AND U5107 ( .A(n4010), .B(n4009), .Z(n4028) );
  XOR U5108 ( .A(a[81]), .B(n2187), .Z(n4032) );
  AND U5109 ( .A(a[83]), .B(b[0]), .Z(n4012) );
  XNOR U5110 ( .A(n4012), .B(n2175), .Z(n4014) );
  NANDN U5111 ( .A(b[0]), .B(a[82]), .Z(n4013) );
  NAND U5112 ( .A(n4014), .B(n4013), .Z(n4037) );
  AND U5113 ( .A(a[79]), .B(b[3]), .Z(n4036) );
  XOR U5114 ( .A(n4037), .B(n4036), .Z(n4039) );
  XOR U5115 ( .A(n4038), .B(n4039), .Z(n4027) );
  NANDN U5116 ( .A(n4016), .B(n4015), .Z(n4020) );
  OR U5117 ( .A(n4018), .B(n4017), .Z(n4019) );
  AND U5118 ( .A(n4020), .B(n4019), .Z(n4026) );
  XOR U5119 ( .A(n4027), .B(n4026), .Z(n4029) );
  XOR U5120 ( .A(n4028), .B(n4029), .Z(n4042) );
  XNOR U5121 ( .A(n4042), .B(sreg[1103]), .Z(n4044) );
  NANDN U5122 ( .A(n4021), .B(sreg[1102]), .Z(n4025) );
  NAND U5123 ( .A(n4023), .B(n4022), .Z(n4024) );
  NAND U5124 ( .A(n4025), .B(n4024), .Z(n4043) );
  XOR U5125 ( .A(n4044), .B(n4043), .Z(c[1103]) );
  NANDN U5126 ( .A(n4027), .B(n4026), .Z(n4031) );
  OR U5127 ( .A(n4029), .B(n4028), .Z(n4030) );
  AND U5128 ( .A(n4031), .B(n4030), .Z(n4049) );
  XOR U5129 ( .A(a[82]), .B(n2187), .Z(n4053) );
  AND U5130 ( .A(a[84]), .B(b[0]), .Z(n4033) );
  XNOR U5131 ( .A(n4033), .B(n2175), .Z(n4035) );
  NANDN U5132 ( .A(b[0]), .B(a[83]), .Z(n4034) );
  NAND U5133 ( .A(n4035), .B(n4034), .Z(n4058) );
  AND U5134 ( .A(a[80]), .B(b[3]), .Z(n4057) );
  XOR U5135 ( .A(n4058), .B(n4057), .Z(n4060) );
  XOR U5136 ( .A(n4059), .B(n4060), .Z(n4048) );
  NANDN U5137 ( .A(n4037), .B(n4036), .Z(n4041) );
  OR U5138 ( .A(n4039), .B(n4038), .Z(n4040) );
  AND U5139 ( .A(n4041), .B(n4040), .Z(n4047) );
  XOR U5140 ( .A(n4048), .B(n4047), .Z(n4050) );
  XOR U5141 ( .A(n4049), .B(n4050), .Z(n4063) );
  XNOR U5142 ( .A(n4063), .B(sreg[1104]), .Z(n4065) );
  NANDN U5143 ( .A(n4042), .B(sreg[1103]), .Z(n4046) );
  NAND U5144 ( .A(n4044), .B(n4043), .Z(n4045) );
  NAND U5145 ( .A(n4046), .B(n4045), .Z(n4064) );
  XOR U5146 ( .A(n4065), .B(n4064), .Z(c[1104]) );
  NANDN U5147 ( .A(n4048), .B(n4047), .Z(n4052) );
  OR U5148 ( .A(n4050), .B(n4049), .Z(n4051) );
  AND U5149 ( .A(n4052), .B(n4051), .Z(n4070) );
  XOR U5150 ( .A(a[83]), .B(n2188), .Z(n4074) );
  AND U5151 ( .A(a[85]), .B(b[0]), .Z(n4054) );
  XNOR U5152 ( .A(n4054), .B(n2175), .Z(n4056) );
  NANDN U5153 ( .A(b[0]), .B(a[84]), .Z(n4055) );
  NAND U5154 ( .A(n4056), .B(n4055), .Z(n4079) );
  AND U5155 ( .A(a[81]), .B(b[3]), .Z(n4078) );
  XOR U5156 ( .A(n4079), .B(n4078), .Z(n4081) );
  XOR U5157 ( .A(n4080), .B(n4081), .Z(n4069) );
  NANDN U5158 ( .A(n4058), .B(n4057), .Z(n4062) );
  OR U5159 ( .A(n4060), .B(n4059), .Z(n4061) );
  AND U5160 ( .A(n4062), .B(n4061), .Z(n4068) );
  XOR U5161 ( .A(n4069), .B(n4068), .Z(n4071) );
  XOR U5162 ( .A(n4070), .B(n4071), .Z(n4084) );
  XNOR U5163 ( .A(n4084), .B(sreg[1105]), .Z(n4086) );
  NANDN U5164 ( .A(n4063), .B(sreg[1104]), .Z(n4067) );
  NAND U5165 ( .A(n4065), .B(n4064), .Z(n4066) );
  NAND U5166 ( .A(n4067), .B(n4066), .Z(n4085) );
  XOR U5167 ( .A(n4086), .B(n4085), .Z(c[1105]) );
  NANDN U5168 ( .A(n4069), .B(n4068), .Z(n4073) );
  OR U5169 ( .A(n4071), .B(n4070), .Z(n4072) );
  AND U5170 ( .A(n4073), .B(n4072), .Z(n4091) );
  XOR U5171 ( .A(a[84]), .B(n2188), .Z(n4095) );
  AND U5172 ( .A(a[86]), .B(b[0]), .Z(n4075) );
  XNOR U5173 ( .A(n4075), .B(n2175), .Z(n4077) );
  NANDN U5174 ( .A(b[0]), .B(a[85]), .Z(n4076) );
  NAND U5175 ( .A(n4077), .B(n4076), .Z(n4100) );
  AND U5176 ( .A(a[82]), .B(b[3]), .Z(n4099) );
  XOR U5177 ( .A(n4100), .B(n4099), .Z(n4102) );
  XOR U5178 ( .A(n4101), .B(n4102), .Z(n4090) );
  NANDN U5179 ( .A(n4079), .B(n4078), .Z(n4083) );
  OR U5180 ( .A(n4081), .B(n4080), .Z(n4082) );
  AND U5181 ( .A(n4083), .B(n4082), .Z(n4089) );
  XOR U5182 ( .A(n4090), .B(n4089), .Z(n4092) );
  XOR U5183 ( .A(n4091), .B(n4092), .Z(n4105) );
  XNOR U5184 ( .A(n4105), .B(sreg[1106]), .Z(n4107) );
  NANDN U5185 ( .A(n4084), .B(sreg[1105]), .Z(n4088) );
  NAND U5186 ( .A(n4086), .B(n4085), .Z(n4087) );
  NAND U5187 ( .A(n4088), .B(n4087), .Z(n4106) );
  XOR U5188 ( .A(n4107), .B(n4106), .Z(c[1106]) );
  NANDN U5189 ( .A(n4090), .B(n4089), .Z(n4094) );
  OR U5190 ( .A(n4092), .B(n4091), .Z(n4093) );
  AND U5191 ( .A(n4094), .B(n4093), .Z(n4112) );
  XOR U5192 ( .A(a[85]), .B(n2188), .Z(n4116) );
  AND U5193 ( .A(a[87]), .B(b[0]), .Z(n4096) );
  XNOR U5194 ( .A(n4096), .B(n2175), .Z(n4098) );
  NANDN U5195 ( .A(b[0]), .B(a[86]), .Z(n4097) );
  NAND U5196 ( .A(n4098), .B(n4097), .Z(n4121) );
  AND U5197 ( .A(a[83]), .B(b[3]), .Z(n4120) );
  XOR U5198 ( .A(n4121), .B(n4120), .Z(n4123) );
  XOR U5199 ( .A(n4122), .B(n4123), .Z(n4111) );
  NANDN U5200 ( .A(n4100), .B(n4099), .Z(n4104) );
  OR U5201 ( .A(n4102), .B(n4101), .Z(n4103) );
  AND U5202 ( .A(n4104), .B(n4103), .Z(n4110) );
  XOR U5203 ( .A(n4111), .B(n4110), .Z(n4113) );
  XOR U5204 ( .A(n4112), .B(n4113), .Z(n4126) );
  XNOR U5205 ( .A(n4126), .B(sreg[1107]), .Z(n4128) );
  NANDN U5206 ( .A(n4105), .B(sreg[1106]), .Z(n4109) );
  NAND U5207 ( .A(n4107), .B(n4106), .Z(n4108) );
  NAND U5208 ( .A(n4109), .B(n4108), .Z(n4127) );
  XOR U5209 ( .A(n4128), .B(n4127), .Z(c[1107]) );
  NANDN U5210 ( .A(n4111), .B(n4110), .Z(n4115) );
  OR U5211 ( .A(n4113), .B(n4112), .Z(n4114) );
  AND U5212 ( .A(n4115), .B(n4114), .Z(n4133) );
  XOR U5213 ( .A(a[86]), .B(n2188), .Z(n4137) );
  AND U5214 ( .A(a[88]), .B(b[0]), .Z(n4117) );
  XNOR U5215 ( .A(n4117), .B(n2175), .Z(n4119) );
  NANDN U5216 ( .A(b[0]), .B(a[87]), .Z(n4118) );
  NAND U5217 ( .A(n4119), .B(n4118), .Z(n4142) );
  AND U5218 ( .A(a[84]), .B(b[3]), .Z(n4141) );
  XOR U5219 ( .A(n4142), .B(n4141), .Z(n4144) );
  XOR U5220 ( .A(n4143), .B(n4144), .Z(n4132) );
  NANDN U5221 ( .A(n4121), .B(n4120), .Z(n4125) );
  OR U5222 ( .A(n4123), .B(n4122), .Z(n4124) );
  AND U5223 ( .A(n4125), .B(n4124), .Z(n4131) );
  XOR U5224 ( .A(n4132), .B(n4131), .Z(n4134) );
  XOR U5225 ( .A(n4133), .B(n4134), .Z(n4147) );
  XNOR U5226 ( .A(n4147), .B(sreg[1108]), .Z(n4149) );
  NANDN U5227 ( .A(n4126), .B(sreg[1107]), .Z(n4130) );
  NAND U5228 ( .A(n4128), .B(n4127), .Z(n4129) );
  NAND U5229 ( .A(n4130), .B(n4129), .Z(n4148) );
  XOR U5230 ( .A(n4149), .B(n4148), .Z(c[1108]) );
  NANDN U5231 ( .A(n4132), .B(n4131), .Z(n4136) );
  OR U5232 ( .A(n4134), .B(n4133), .Z(n4135) );
  AND U5233 ( .A(n4136), .B(n4135), .Z(n4154) );
  XOR U5234 ( .A(a[87]), .B(n2188), .Z(n4158) );
  AND U5235 ( .A(a[89]), .B(b[0]), .Z(n4138) );
  XNOR U5236 ( .A(n4138), .B(n2175), .Z(n4140) );
  NANDN U5237 ( .A(b[0]), .B(a[88]), .Z(n4139) );
  NAND U5238 ( .A(n4140), .B(n4139), .Z(n4163) );
  AND U5239 ( .A(a[85]), .B(b[3]), .Z(n4162) );
  XOR U5240 ( .A(n4163), .B(n4162), .Z(n4165) );
  XOR U5241 ( .A(n4164), .B(n4165), .Z(n4153) );
  NANDN U5242 ( .A(n4142), .B(n4141), .Z(n4146) );
  OR U5243 ( .A(n4144), .B(n4143), .Z(n4145) );
  AND U5244 ( .A(n4146), .B(n4145), .Z(n4152) );
  XOR U5245 ( .A(n4153), .B(n4152), .Z(n4155) );
  XOR U5246 ( .A(n4154), .B(n4155), .Z(n4168) );
  XNOR U5247 ( .A(n4168), .B(sreg[1109]), .Z(n4170) );
  NANDN U5248 ( .A(n4147), .B(sreg[1108]), .Z(n4151) );
  NAND U5249 ( .A(n4149), .B(n4148), .Z(n4150) );
  NAND U5250 ( .A(n4151), .B(n4150), .Z(n4169) );
  XOR U5251 ( .A(n4170), .B(n4169), .Z(c[1109]) );
  NANDN U5252 ( .A(n4153), .B(n4152), .Z(n4157) );
  OR U5253 ( .A(n4155), .B(n4154), .Z(n4156) );
  AND U5254 ( .A(n4157), .B(n4156), .Z(n4175) );
  XOR U5255 ( .A(a[88]), .B(n2188), .Z(n4179) );
  AND U5256 ( .A(a[90]), .B(b[0]), .Z(n4159) );
  XNOR U5257 ( .A(n4159), .B(n2175), .Z(n4161) );
  NANDN U5258 ( .A(b[0]), .B(a[89]), .Z(n4160) );
  NAND U5259 ( .A(n4161), .B(n4160), .Z(n4184) );
  AND U5260 ( .A(a[86]), .B(b[3]), .Z(n4183) );
  XOR U5261 ( .A(n4184), .B(n4183), .Z(n4186) );
  XOR U5262 ( .A(n4185), .B(n4186), .Z(n4174) );
  NANDN U5263 ( .A(n4163), .B(n4162), .Z(n4167) );
  OR U5264 ( .A(n4165), .B(n4164), .Z(n4166) );
  AND U5265 ( .A(n4167), .B(n4166), .Z(n4173) );
  XOR U5266 ( .A(n4174), .B(n4173), .Z(n4176) );
  XOR U5267 ( .A(n4175), .B(n4176), .Z(n4189) );
  XNOR U5268 ( .A(n4189), .B(sreg[1110]), .Z(n4191) );
  NANDN U5269 ( .A(n4168), .B(sreg[1109]), .Z(n4172) );
  NAND U5270 ( .A(n4170), .B(n4169), .Z(n4171) );
  NAND U5271 ( .A(n4172), .B(n4171), .Z(n4190) );
  XOR U5272 ( .A(n4191), .B(n4190), .Z(c[1110]) );
  NANDN U5273 ( .A(n4174), .B(n4173), .Z(n4178) );
  OR U5274 ( .A(n4176), .B(n4175), .Z(n4177) );
  AND U5275 ( .A(n4178), .B(n4177), .Z(n4196) );
  XOR U5276 ( .A(a[89]), .B(n2188), .Z(n4200) );
  AND U5277 ( .A(a[91]), .B(b[0]), .Z(n4180) );
  XNOR U5278 ( .A(n4180), .B(n2175), .Z(n4182) );
  NANDN U5279 ( .A(b[0]), .B(a[90]), .Z(n4181) );
  NAND U5280 ( .A(n4182), .B(n4181), .Z(n4205) );
  AND U5281 ( .A(a[87]), .B(b[3]), .Z(n4204) );
  XOR U5282 ( .A(n4205), .B(n4204), .Z(n4207) );
  XOR U5283 ( .A(n4206), .B(n4207), .Z(n4195) );
  NANDN U5284 ( .A(n4184), .B(n4183), .Z(n4188) );
  OR U5285 ( .A(n4186), .B(n4185), .Z(n4187) );
  AND U5286 ( .A(n4188), .B(n4187), .Z(n4194) );
  XOR U5287 ( .A(n4195), .B(n4194), .Z(n4197) );
  XOR U5288 ( .A(n4196), .B(n4197), .Z(n4210) );
  XNOR U5289 ( .A(n4210), .B(sreg[1111]), .Z(n4212) );
  NANDN U5290 ( .A(n4189), .B(sreg[1110]), .Z(n4193) );
  NAND U5291 ( .A(n4191), .B(n4190), .Z(n4192) );
  NAND U5292 ( .A(n4193), .B(n4192), .Z(n4211) );
  XOR U5293 ( .A(n4212), .B(n4211), .Z(c[1111]) );
  NANDN U5294 ( .A(n4195), .B(n4194), .Z(n4199) );
  OR U5295 ( .A(n4197), .B(n4196), .Z(n4198) );
  AND U5296 ( .A(n4199), .B(n4198), .Z(n4217) );
  XOR U5297 ( .A(a[90]), .B(n2189), .Z(n4221) );
  AND U5298 ( .A(a[92]), .B(b[0]), .Z(n4201) );
  XNOR U5299 ( .A(n4201), .B(n2175), .Z(n4203) );
  NANDN U5300 ( .A(b[0]), .B(a[91]), .Z(n4202) );
  NAND U5301 ( .A(n4203), .B(n4202), .Z(n4226) );
  AND U5302 ( .A(a[88]), .B(b[3]), .Z(n4225) );
  XOR U5303 ( .A(n4226), .B(n4225), .Z(n4228) );
  XOR U5304 ( .A(n4227), .B(n4228), .Z(n4216) );
  NANDN U5305 ( .A(n4205), .B(n4204), .Z(n4209) );
  OR U5306 ( .A(n4207), .B(n4206), .Z(n4208) );
  AND U5307 ( .A(n4209), .B(n4208), .Z(n4215) );
  XOR U5308 ( .A(n4216), .B(n4215), .Z(n4218) );
  XOR U5309 ( .A(n4217), .B(n4218), .Z(n4231) );
  XNOR U5310 ( .A(n4231), .B(sreg[1112]), .Z(n4233) );
  NANDN U5311 ( .A(n4210), .B(sreg[1111]), .Z(n4214) );
  NAND U5312 ( .A(n4212), .B(n4211), .Z(n4213) );
  NAND U5313 ( .A(n4214), .B(n4213), .Z(n4232) );
  XOR U5314 ( .A(n4233), .B(n4232), .Z(c[1112]) );
  NANDN U5315 ( .A(n4216), .B(n4215), .Z(n4220) );
  OR U5316 ( .A(n4218), .B(n4217), .Z(n4219) );
  AND U5317 ( .A(n4220), .B(n4219), .Z(n4238) );
  XOR U5318 ( .A(a[91]), .B(n2189), .Z(n4242) );
  AND U5319 ( .A(a[93]), .B(b[0]), .Z(n4222) );
  XNOR U5320 ( .A(n4222), .B(n2175), .Z(n4224) );
  NANDN U5321 ( .A(b[0]), .B(a[92]), .Z(n4223) );
  NAND U5322 ( .A(n4224), .B(n4223), .Z(n4247) );
  AND U5323 ( .A(a[89]), .B(b[3]), .Z(n4246) );
  XOR U5324 ( .A(n4247), .B(n4246), .Z(n4249) );
  XOR U5325 ( .A(n4248), .B(n4249), .Z(n4237) );
  NANDN U5326 ( .A(n4226), .B(n4225), .Z(n4230) );
  OR U5327 ( .A(n4228), .B(n4227), .Z(n4229) );
  AND U5328 ( .A(n4230), .B(n4229), .Z(n4236) );
  XOR U5329 ( .A(n4237), .B(n4236), .Z(n4239) );
  XOR U5330 ( .A(n4238), .B(n4239), .Z(n4252) );
  XNOR U5331 ( .A(n4252), .B(sreg[1113]), .Z(n4254) );
  NANDN U5332 ( .A(n4231), .B(sreg[1112]), .Z(n4235) );
  NAND U5333 ( .A(n4233), .B(n4232), .Z(n4234) );
  NAND U5334 ( .A(n4235), .B(n4234), .Z(n4253) );
  XOR U5335 ( .A(n4254), .B(n4253), .Z(c[1113]) );
  NANDN U5336 ( .A(n4237), .B(n4236), .Z(n4241) );
  OR U5337 ( .A(n4239), .B(n4238), .Z(n4240) );
  AND U5338 ( .A(n4241), .B(n4240), .Z(n4259) );
  XOR U5339 ( .A(a[92]), .B(n2189), .Z(n4263) );
  AND U5340 ( .A(a[94]), .B(b[0]), .Z(n4243) );
  XNOR U5341 ( .A(n4243), .B(n2175), .Z(n4245) );
  NANDN U5342 ( .A(b[0]), .B(a[93]), .Z(n4244) );
  NAND U5343 ( .A(n4245), .B(n4244), .Z(n4268) );
  AND U5344 ( .A(a[90]), .B(b[3]), .Z(n4267) );
  XOR U5345 ( .A(n4268), .B(n4267), .Z(n4270) );
  XOR U5346 ( .A(n4269), .B(n4270), .Z(n4258) );
  NANDN U5347 ( .A(n4247), .B(n4246), .Z(n4251) );
  OR U5348 ( .A(n4249), .B(n4248), .Z(n4250) );
  AND U5349 ( .A(n4251), .B(n4250), .Z(n4257) );
  XOR U5350 ( .A(n4258), .B(n4257), .Z(n4260) );
  XOR U5351 ( .A(n4259), .B(n4260), .Z(n4273) );
  XNOR U5352 ( .A(n4273), .B(sreg[1114]), .Z(n4275) );
  NANDN U5353 ( .A(n4252), .B(sreg[1113]), .Z(n4256) );
  NAND U5354 ( .A(n4254), .B(n4253), .Z(n4255) );
  NAND U5355 ( .A(n4256), .B(n4255), .Z(n4274) );
  XOR U5356 ( .A(n4275), .B(n4274), .Z(c[1114]) );
  NANDN U5357 ( .A(n4258), .B(n4257), .Z(n4262) );
  OR U5358 ( .A(n4260), .B(n4259), .Z(n4261) );
  AND U5359 ( .A(n4262), .B(n4261), .Z(n4280) );
  XOR U5360 ( .A(a[93]), .B(n2189), .Z(n4284) );
  AND U5361 ( .A(a[95]), .B(b[0]), .Z(n4264) );
  XNOR U5362 ( .A(n4264), .B(n2175), .Z(n4266) );
  NANDN U5363 ( .A(b[0]), .B(a[94]), .Z(n4265) );
  NAND U5364 ( .A(n4266), .B(n4265), .Z(n4289) );
  AND U5365 ( .A(a[91]), .B(b[3]), .Z(n4288) );
  XOR U5366 ( .A(n4289), .B(n4288), .Z(n4291) );
  XOR U5367 ( .A(n4290), .B(n4291), .Z(n4279) );
  NANDN U5368 ( .A(n4268), .B(n4267), .Z(n4272) );
  OR U5369 ( .A(n4270), .B(n4269), .Z(n4271) );
  AND U5370 ( .A(n4272), .B(n4271), .Z(n4278) );
  XOR U5371 ( .A(n4279), .B(n4278), .Z(n4281) );
  XOR U5372 ( .A(n4280), .B(n4281), .Z(n4294) );
  XNOR U5373 ( .A(n4294), .B(sreg[1115]), .Z(n4296) );
  NANDN U5374 ( .A(n4273), .B(sreg[1114]), .Z(n4277) );
  NAND U5375 ( .A(n4275), .B(n4274), .Z(n4276) );
  NAND U5376 ( .A(n4277), .B(n4276), .Z(n4295) );
  XOR U5377 ( .A(n4296), .B(n4295), .Z(c[1115]) );
  NANDN U5378 ( .A(n4279), .B(n4278), .Z(n4283) );
  OR U5379 ( .A(n4281), .B(n4280), .Z(n4282) );
  AND U5380 ( .A(n4283), .B(n4282), .Z(n4301) );
  XOR U5381 ( .A(a[94]), .B(n2189), .Z(n4305) );
  AND U5382 ( .A(a[92]), .B(b[3]), .Z(n4309) );
  AND U5383 ( .A(a[96]), .B(b[0]), .Z(n4285) );
  XNOR U5384 ( .A(n4285), .B(n2175), .Z(n4287) );
  NANDN U5385 ( .A(b[0]), .B(a[95]), .Z(n4286) );
  NAND U5386 ( .A(n4287), .B(n4286), .Z(n4310) );
  XOR U5387 ( .A(n4309), .B(n4310), .Z(n4312) );
  XOR U5388 ( .A(n4311), .B(n4312), .Z(n4300) );
  NANDN U5389 ( .A(n4289), .B(n4288), .Z(n4293) );
  OR U5390 ( .A(n4291), .B(n4290), .Z(n4292) );
  AND U5391 ( .A(n4293), .B(n4292), .Z(n4299) );
  XOR U5392 ( .A(n4300), .B(n4299), .Z(n4302) );
  XOR U5393 ( .A(n4301), .B(n4302), .Z(n4315) );
  XNOR U5394 ( .A(n4315), .B(sreg[1116]), .Z(n4317) );
  NANDN U5395 ( .A(n4294), .B(sreg[1115]), .Z(n4298) );
  NAND U5396 ( .A(n4296), .B(n4295), .Z(n4297) );
  NAND U5397 ( .A(n4298), .B(n4297), .Z(n4316) );
  XOR U5398 ( .A(n4317), .B(n4316), .Z(c[1116]) );
  NANDN U5399 ( .A(n4300), .B(n4299), .Z(n4304) );
  OR U5400 ( .A(n4302), .B(n4301), .Z(n4303) );
  AND U5401 ( .A(n4304), .B(n4303), .Z(n4322) );
  XOR U5402 ( .A(a[95]), .B(n2189), .Z(n4326) );
  AND U5403 ( .A(a[97]), .B(b[0]), .Z(n4306) );
  XNOR U5404 ( .A(n4306), .B(n2175), .Z(n4308) );
  NANDN U5405 ( .A(b[0]), .B(a[96]), .Z(n4307) );
  NAND U5406 ( .A(n4308), .B(n4307), .Z(n4331) );
  AND U5407 ( .A(a[93]), .B(b[3]), .Z(n4330) );
  XOR U5408 ( .A(n4331), .B(n4330), .Z(n4333) );
  XOR U5409 ( .A(n4332), .B(n4333), .Z(n4321) );
  NANDN U5410 ( .A(n4310), .B(n4309), .Z(n4314) );
  OR U5411 ( .A(n4312), .B(n4311), .Z(n4313) );
  AND U5412 ( .A(n4314), .B(n4313), .Z(n4320) );
  XOR U5413 ( .A(n4321), .B(n4320), .Z(n4323) );
  XOR U5414 ( .A(n4322), .B(n4323), .Z(n4336) );
  XNOR U5415 ( .A(n4336), .B(sreg[1117]), .Z(n4338) );
  NANDN U5416 ( .A(n4315), .B(sreg[1116]), .Z(n4319) );
  NAND U5417 ( .A(n4317), .B(n4316), .Z(n4318) );
  NAND U5418 ( .A(n4319), .B(n4318), .Z(n4337) );
  XOR U5419 ( .A(n4338), .B(n4337), .Z(c[1117]) );
  NANDN U5420 ( .A(n4321), .B(n4320), .Z(n4325) );
  OR U5421 ( .A(n4323), .B(n4322), .Z(n4324) );
  AND U5422 ( .A(n4325), .B(n4324), .Z(n4343) );
  XOR U5423 ( .A(a[96]), .B(n2189), .Z(n4347) );
  AND U5424 ( .A(a[98]), .B(b[0]), .Z(n4327) );
  XNOR U5425 ( .A(n4327), .B(n2175), .Z(n4329) );
  NANDN U5426 ( .A(b[0]), .B(a[97]), .Z(n4328) );
  NAND U5427 ( .A(n4329), .B(n4328), .Z(n4352) );
  AND U5428 ( .A(a[94]), .B(b[3]), .Z(n4351) );
  XOR U5429 ( .A(n4352), .B(n4351), .Z(n4354) );
  XOR U5430 ( .A(n4353), .B(n4354), .Z(n4342) );
  NANDN U5431 ( .A(n4331), .B(n4330), .Z(n4335) );
  OR U5432 ( .A(n4333), .B(n4332), .Z(n4334) );
  AND U5433 ( .A(n4335), .B(n4334), .Z(n4341) );
  XOR U5434 ( .A(n4342), .B(n4341), .Z(n4344) );
  XOR U5435 ( .A(n4343), .B(n4344), .Z(n4357) );
  XNOR U5436 ( .A(n4357), .B(sreg[1118]), .Z(n4359) );
  NANDN U5437 ( .A(n4336), .B(sreg[1117]), .Z(n4340) );
  NAND U5438 ( .A(n4338), .B(n4337), .Z(n4339) );
  NAND U5439 ( .A(n4340), .B(n4339), .Z(n4358) );
  XOR U5440 ( .A(n4359), .B(n4358), .Z(c[1118]) );
  NANDN U5441 ( .A(n4342), .B(n4341), .Z(n4346) );
  OR U5442 ( .A(n4344), .B(n4343), .Z(n4345) );
  AND U5443 ( .A(n4346), .B(n4345), .Z(n4364) );
  XOR U5444 ( .A(a[97]), .B(n2190), .Z(n4368) );
  AND U5445 ( .A(a[95]), .B(b[3]), .Z(n4372) );
  AND U5446 ( .A(a[99]), .B(b[0]), .Z(n4348) );
  XNOR U5447 ( .A(n4348), .B(n2175), .Z(n4350) );
  NANDN U5448 ( .A(b[0]), .B(a[98]), .Z(n4349) );
  NAND U5449 ( .A(n4350), .B(n4349), .Z(n4373) );
  XOR U5450 ( .A(n4372), .B(n4373), .Z(n4375) );
  XOR U5451 ( .A(n4374), .B(n4375), .Z(n4363) );
  NANDN U5452 ( .A(n4352), .B(n4351), .Z(n4356) );
  OR U5453 ( .A(n4354), .B(n4353), .Z(n4355) );
  AND U5454 ( .A(n4356), .B(n4355), .Z(n4362) );
  XOR U5455 ( .A(n4363), .B(n4362), .Z(n4365) );
  XOR U5456 ( .A(n4364), .B(n4365), .Z(n4378) );
  XNOR U5457 ( .A(n4378), .B(sreg[1119]), .Z(n4380) );
  NANDN U5458 ( .A(n4357), .B(sreg[1118]), .Z(n4361) );
  NAND U5459 ( .A(n4359), .B(n4358), .Z(n4360) );
  NAND U5460 ( .A(n4361), .B(n4360), .Z(n4379) );
  XOR U5461 ( .A(n4380), .B(n4379), .Z(c[1119]) );
  NANDN U5462 ( .A(n4363), .B(n4362), .Z(n4367) );
  OR U5463 ( .A(n4365), .B(n4364), .Z(n4366) );
  AND U5464 ( .A(n4367), .B(n4366), .Z(n4385) );
  XOR U5465 ( .A(a[98]), .B(n2190), .Z(n4389) );
  AND U5466 ( .A(a[100]), .B(b[0]), .Z(n4369) );
  XNOR U5467 ( .A(n4369), .B(n2175), .Z(n4371) );
  NANDN U5468 ( .A(b[0]), .B(a[99]), .Z(n4370) );
  NAND U5469 ( .A(n4371), .B(n4370), .Z(n4394) );
  AND U5470 ( .A(a[96]), .B(b[3]), .Z(n4393) );
  XOR U5471 ( .A(n4394), .B(n4393), .Z(n4396) );
  XOR U5472 ( .A(n4395), .B(n4396), .Z(n4384) );
  NANDN U5473 ( .A(n4373), .B(n4372), .Z(n4377) );
  OR U5474 ( .A(n4375), .B(n4374), .Z(n4376) );
  AND U5475 ( .A(n4377), .B(n4376), .Z(n4383) );
  XOR U5476 ( .A(n4384), .B(n4383), .Z(n4386) );
  XOR U5477 ( .A(n4385), .B(n4386), .Z(n4399) );
  XNOR U5478 ( .A(n4399), .B(sreg[1120]), .Z(n4401) );
  NANDN U5479 ( .A(n4378), .B(sreg[1119]), .Z(n4382) );
  NAND U5480 ( .A(n4380), .B(n4379), .Z(n4381) );
  NAND U5481 ( .A(n4382), .B(n4381), .Z(n4400) );
  XOR U5482 ( .A(n4401), .B(n4400), .Z(c[1120]) );
  NANDN U5483 ( .A(n4384), .B(n4383), .Z(n4388) );
  OR U5484 ( .A(n4386), .B(n4385), .Z(n4387) );
  AND U5485 ( .A(n4388), .B(n4387), .Z(n4407) );
  XOR U5486 ( .A(a[99]), .B(n2190), .Z(n4408) );
  AND U5487 ( .A(b[0]), .B(a[101]), .Z(n4390) );
  XOR U5488 ( .A(b[1]), .B(n4390), .Z(n4392) );
  NANDN U5489 ( .A(b[0]), .B(a[100]), .Z(n4391) );
  AND U5490 ( .A(n4392), .B(n4391), .Z(n4412) );
  AND U5491 ( .A(a[97]), .B(b[3]), .Z(n4413) );
  XOR U5492 ( .A(n4412), .B(n4413), .Z(n4414) );
  XNOR U5493 ( .A(n4415), .B(n4414), .Z(n4404) );
  NANDN U5494 ( .A(n4394), .B(n4393), .Z(n4398) );
  OR U5495 ( .A(n4396), .B(n4395), .Z(n4397) );
  AND U5496 ( .A(n4398), .B(n4397), .Z(n4405) );
  XNOR U5497 ( .A(n4404), .B(n4405), .Z(n4406) );
  XNOR U5498 ( .A(n4407), .B(n4406), .Z(n4418) );
  XNOR U5499 ( .A(n4418), .B(sreg[1121]), .Z(n4420) );
  NANDN U5500 ( .A(n4399), .B(sreg[1120]), .Z(n4403) );
  NAND U5501 ( .A(n4401), .B(n4400), .Z(n4402) );
  NAND U5502 ( .A(n4403), .B(n4402), .Z(n4419) );
  XOR U5503 ( .A(n4420), .B(n4419), .Z(c[1121]) );
  XOR U5504 ( .A(a[100]), .B(n2190), .Z(n4427) );
  AND U5505 ( .A(a[102]), .B(b[0]), .Z(n4409) );
  XNOR U5506 ( .A(n4409), .B(n2175), .Z(n4411) );
  NANDN U5507 ( .A(b[0]), .B(a[101]), .Z(n4410) );
  NAND U5508 ( .A(n4411), .B(n4410), .Z(n4432) );
  AND U5509 ( .A(a[98]), .B(b[3]), .Z(n4431) );
  XOR U5510 ( .A(n4432), .B(n4431), .Z(n4434) );
  XOR U5511 ( .A(n4433), .B(n4434), .Z(n4422) );
  NAND U5512 ( .A(n4413), .B(n4412), .Z(n4417) );
  NANDN U5513 ( .A(n4415), .B(n4414), .Z(n4416) );
  AND U5514 ( .A(n4417), .B(n4416), .Z(n4421) );
  XOR U5515 ( .A(n4422), .B(n4421), .Z(n4424) );
  XOR U5516 ( .A(n4423), .B(n4424), .Z(n4437) );
  XNOR U5517 ( .A(n4437), .B(sreg[1122]), .Z(n4439) );
  XOR U5518 ( .A(n4439), .B(n4438), .Z(c[1122]) );
  NANDN U5519 ( .A(n4422), .B(n4421), .Z(n4426) );
  OR U5520 ( .A(n4424), .B(n4423), .Z(n4425) );
  AND U5521 ( .A(n4426), .B(n4425), .Z(n4444) );
  XOR U5522 ( .A(a[101]), .B(n2190), .Z(n4448) );
  AND U5523 ( .A(a[99]), .B(b[3]), .Z(n4452) );
  AND U5524 ( .A(a[103]), .B(b[0]), .Z(n4428) );
  XNOR U5525 ( .A(n4428), .B(n2175), .Z(n4430) );
  NANDN U5526 ( .A(b[0]), .B(a[102]), .Z(n4429) );
  NAND U5527 ( .A(n4430), .B(n4429), .Z(n4453) );
  XOR U5528 ( .A(n4452), .B(n4453), .Z(n4455) );
  XOR U5529 ( .A(n4454), .B(n4455), .Z(n4443) );
  NANDN U5530 ( .A(n4432), .B(n4431), .Z(n4436) );
  OR U5531 ( .A(n4434), .B(n4433), .Z(n4435) );
  AND U5532 ( .A(n4436), .B(n4435), .Z(n4442) );
  XOR U5533 ( .A(n4443), .B(n4442), .Z(n4445) );
  XOR U5534 ( .A(n4444), .B(n4445), .Z(n4458) );
  XNOR U5535 ( .A(n4458), .B(sreg[1123]), .Z(n4460) );
  NANDN U5536 ( .A(n4437), .B(sreg[1122]), .Z(n4441) );
  NAND U5537 ( .A(n4439), .B(n4438), .Z(n4440) );
  NAND U5538 ( .A(n4441), .B(n4440), .Z(n4459) );
  XOR U5539 ( .A(n4460), .B(n4459), .Z(c[1123]) );
  NANDN U5540 ( .A(n4443), .B(n4442), .Z(n4447) );
  OR U5541 ( .A(n4445), .B(n4444), .Z(n4446) );
  AND U5542 ( .A(n4447), .B(n4446), .Z(n4465) );
  XOR U5543 ( .A(a[102]), .B(n2190), .Z(n4469) );
  AND U5544 ( .A(a[104]), .B(b[0]), .Z(n4449) );
  XNOR U5545 ( .A(n4449), .B(n2175), .Z(n4451) );
  NANDN U5546 ( .A(b[0]), .B(a[103]), .Z(n4450) );
  NAND U5547 ( .A(n4451), .B(n4450), .Z(n4474) );
  AND U5548 ( .A(a[100]), .B(b[3]), .Z(n4473) );
  XOR U5549 ( .A(n4474), .B(n4473), .Z(n4476) );
  XOR U5550 ( .A(n4475), .B(n4476), .Z(n4464) );
  NANDN U5551 ( .A(n4453), .B(n4452), .Z(n4457) );
  OR U5552 ( .A(n4455), .B(n4454), .Z(n4456) );
  AND U5553 ( .A(n4457), .B(n4456), .Z(n4463) );
  XOR U5554 ( .A(n4464), .B(n4463), .Z(n4466) );
  XOR U5555 ( .A(n4465), .B(n4466), .Z(n4479) );
  XNOR U5556 ( .A(n4479), .B(sreg[1124]), .Z(n4481) );
  NANDN U5557 ( .A(n4458), .B(sreg[1123]), .Z(n4462) );
  NAND U5558 ( .A(n4460), .B(n4459), .Z(n4461) );
  NAND U5559 ( .A(n4462), .B(n4461), .Z(n4480) );
  XOR U5560 ( .A(n4481), .B(n4480), .Z(c[1124]) );
  NANDN U5561 ( .A(n4464), .B(n4463), .Z(n4468) );
  OR U5562 ( .A(n4466), .B(n4465), .Z(n4467) );
  AND U5563 ( .A(n4468), .B(n4467), .Z(n4486) );
  XOR U5564 ( .A(a[103]), .B(n2190), .Z(n4490) );
  AND U5565 ( .A(a[101]), .B(b[3]), .Z(n4494) );
  AND U5566 ( .A(a[105]), .B(b[0]), .Z(n4470) );
  XNOR U5567 ( .A(n4470), .B(n2175), .Z(n4472) );
  NANDN U5568 ( .A(b[0]), .B(a[104]), .Z(n4471) );
  NAND U5569 ( .A(n4472), .B(n4471), .Z(n4495) );
  XOR U5570 ( .A(n4494), .B(n4495), .Z(n4497) );
  XOR U5571 ( .A(n4496), .B(n4497), .Z(n4485) );
  NANDN U5572 ( .A(n4474), .B(n4473), .Z(n4478) );
  OR U5573 ( .A(n4476), .B(n4475), .Z(n4477) );
  AND U5574 ( .A(n4478), .B(n4477), .Z(n4484) );
  XOR U5575 ( .A(n4485), .B(n4484), .Z(n4487) );
  XOR U5576 ( .A(n4486), .B(n4487), .Z(n4500) );
  XNOR U5577 ( .A(n4500), .B(sreg[1125]), .Z(n4502) );
  NANDN U5578 ( .A(n4479), .B(sreg[1124]), .Z(n4483) );
  NAND U5579 ( .A(n4481), .B(n4480), .Z(n4482) );
  NAND U5580 ( .A(n4483), .B(n4482), .Z(n4501) );
  XOR U5581 ( .A(n4502), .B(n4501), .Z(c[1125]) );
  NANDN U5582 ( .A(n4485), .B(n4484), .Z(n4489) );
  OR U5583 ( .A(n4487), .B(n4486), .Z(n4488) );
  AND U5584 ( .A(n4489), .B(n4488), .Z(n4507) );
  XOR U5585 ( .A(a[104]), .B(n2191), .Z(n4511) );
  AND U5586 ( .A(a[106]), .B(b[0]), .Z(n4491) );
  XNOR U5587 ( .A(n4491), .B(n2175), .Z(n4493) );
  NANDN U5588 ( .A(b[0]), .B(a[105]), .Z(n4492) );
  NAND U5589 ( .A(n4493), .B(n4492), .Z(n4516) );
  AND U5590 ( .A(a[102]), .B(b[3]), .Z(n4515) );
  XOR U5591 ( .A(n4516), .B(n4515), .Z(n4518) );
  XOR U5592 ( .A(n4517), .B(n4518), .Z(n4506) );
  NANDN U5593 ( .A(n4495), .B(n4494), .Z(n4499) );
  OR U5594 ( .A(n4497), .B(n4496), .Z(n4498) );
  AND U5595 ( .A(n4499), .B(n4498), .Z(n4505) );
  XOR U5596 ( .A(n4506), .B(n4505), .Z(n4508) );
  XOR U5597 ( .A(n4507), .B(n4508), .Z(n4521) );
  XNOR U5598 ( .A(n4521), .B(sreg[1126]), .Z(n4523) );
  NANDN U5599 ( .A(n4500), .B(sreg[1125]), .Z(n4504) );
  NAND U5600 ( .A(n4502), .B(n4501), .Z(n4503) );
  NAND U5601 ( .A(n4504), .B(n4503), .Z(n4522) );
  XOR U5602 ( .A(n4523), .B(n4522), .Z(c[1126]) );
  NANDN U5603 ( .A(n4506), .B(n4505), .Z(n4510) );
  OR U5604 ( .A(n4508), .B(n4507), .Z(n4509) );
  AND U5605 ( .A(n4510), .B(n4509), .Z(n4528) );
  XOR U5606 ( .A(a[105]), .B(n2191), .Z(n4532) );
  AND U5607 ( .A(a[107]), .B(b[0]), .Z(n4512) );
  XNOR U5608 ( .A(n4512), .B(n2175), .Z(n4514) );
  NANDN U5609 ( .A(b[0]), .B(a[106]), .Z(n4513) );
  NAND U5610 ( .A(n4514), .B(n4513), .Z(n4537) );
  AND U5611 ( .A(a[103]), .B(b[3]), .Z(n4536) );
  XOR U5612 ( .A(n4537), .B(n4536), .Z(n4539) );
  XOR U5613 ( .A(n4538), .B(n4539), .Z(n4527) );
  NANDN U5614 ( .A(n4516), .B(n4515), .Z(n4520) );
  OR U5615 ( .A(n4518), .B(n4517), .Z(n4519) );
  AND U5616 ( .A(n4520), .B(n4519), .Z(n4526) );
  XOR U5617 ( .A(n4527), .B(n4526), .Z(n4529) );
  XOR U5618 ( .A(n4528), .B(n4529), .Z(n4542) );
  XNOR U5619 ( .A(n4542), .B(sreg[1127]), .Z(n4544) );
  NANDN U5620 ( .A(n4521), .B(sreg[1126]), .Z(n4525) );
  NAND U5621 ( .A(n4523), .B(n4522), .Z(n4524) );
  NAND U5622 ( .A(n4525), .B(n4524), .Z(n4543) );
  XOR U5623 ( .A(n4544), .B(n4543), .Z(c[1127]) );
  NANDN U5624 ( .A(n4527), .B(n4526), .Z(n4531) );
  OR U5625 ( .A(n4529), .B(n4528), .Z(n4530) );
  AND U5626 ( .A(n4531), .B(n4530), .Z(n4549) );
  XOR U5627 ( .A(a[106]), .B(n2191), .Z(n4553) );
  AND U5628 ( .A(a[108]), .B(b[0]), .Z(n4533) );
  XNOR U5629 ( .A(n4533), .B(n2175), .Z(n4535) );
  NANDN U5630 ( .A(b[0]), .B(a[107]), .Z(n4534) );
  NAND U5631 ( .A(n4535), .B(n4534), .Z(n4558) );
  AND U5632 ( .A(a[104]), .B(b[3]), .Z(n4557) );
  XOR U5633 ( .A(n4558), .B(n4557), .Z(n4560) );
  XOR U5634 ( .A(n4559), .B(n4560), .Z(n4548) );
  NANDN U5635 ( .A(n4537), .B(n4536), .Z(n4541) );
  OR U5636 ( .A(n4539), .B(n4538), .Z(n4540) );
  AND U5637 ( .A(n4541), .B(n4540), .Z(n4547) );
  XOR U5638 ( .A(n4548), .B(n4547), .Z(n4550) );
  XOR U5639 ( .A(n4549), .B(n4550), .Z(n4563) );
  XNOR U5640 ( .A(n4563), .B(sreg[1128]), .Z(n4565) );
  NANDN U5641 ( .A(n4542), .B(sreg[1127]), .Z(n4546) );
  NAND U5642 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U5643 ( .A(n4546), .B(n4545), .Z(n4564) );
  XOR U5644 ( .A(n4565), .B(n4564), .Z(c[1128]) );
  NANDN U5645 ( .A(n4548), .B(n4547), .Z(n4552) );
  OR U5646 ( .A(n4550), .B(n4549), .Z(n4551) );
  AND U5647 ( .A(n4552), .B(n4551), .Z(n4570) );
  XOR U5648 ( .A(a[107]), .B(n2191), .Z(n4574) );
  AND U5649 ( .A(a[105]), .B(b[3]), .Z(n4578) );
  AND U5650 ( .A(a[109]), .B(b[0]), .Z(n4554) );
  XNOR U5651 ( .A(n4554), .B(n2175), .Z(n4556) );
  NANDN U5652 ( .A(b[0]), .B(a[108]), .Z(n4555) );
  NAND U5653 ( .A(n4556), .B(n4555), .Z(n4579) );
  XOR U5654 ( .A(n4578), .B(n4579), .Z(n4581) );
  XOR U5655 ( .A(n4580), .B(n4581), .Z(n4569) );
  NANDN U5656 ( .A(n4558), .B(n4557), .Z(n4562) );
  OR U5657 ( .A(n4560), .B(n4559), .Z(n4561) );
  AND U5658 ( .A(n4562), .B(n4561), .Z(n4568) );
  XOR U5659 ( .A(n4569), .B(n4568), .Z(n4571) );
  XOR U5660 ( .A(n4570), .B(n4571), .Z(n4584) );
  XNOR U5661 ( .A(n4584), .B(sreg[1129]), .Z(n4586) );
  NANDN U5662 ( .A(n4563), .B(sreg[1128]), .Z(n4567) );
  NAND U5663 ( .A(n4565), .B(n4564), .Z(n4566) );
  NAND U5664 ( .A(n4567), .B(n4566), .Z(n4585) );
  XOR U5665 ( .A(n4586), .B(n4585), .Z(c[1129]) );
  NANDN U5666 ( .A(n4569), .B(n4568), .Z(n4573) );
  OR U5667 ( .A(n4571), .B(n4570), .Z(n4572) );
  AND U5668 ( .A(n4573), .B(n4572), .Z(n4591) );
  XOR U5669 ( .A(a[108]), .B(n2191), .Z(n4595) );
  AND U5670 ( .A(a[110]), .B(b[0]), .Z(n4575) );
  XNOR U5671 ( .A(n4575), .B(n2175), .Z(n4577) );
  NANDN U5672 ( .A(b[0]), .B(a[109]), .Z(n4576) );
  NAND U5673 ( .A(n4577), .B(n4576), .Z(n4600) );
  AND U5674 ( .A(a[106]), .B(b[3]), .Z(n4599) );
  XOR U5675 ( .A(n4600), .B(n4599), .Z(n4602) );
  XOR U5676 ( .A(n4601), .B(n4602), .Z(n4590) );
  NANDN U5677 ( .A(n4579), .B(n4578), .Z(n4583) );
  OR U5678 ( .A(n4581), .B(n4580), .Z(n4582) );
  AND U5679 ( .A(n4583), .B(n4582), .Z(n4589) );
  XOR U5680 ( .A(n4590), .B(n4589), .Z(n4592) );
  XOR U5681 ( .A(n4591), .B(n4592), .Z(n4605) );
  XNOR U5682 ( .A(n4605), .B(sreg[1130]), .Z(n4607) );
  NANDN U5683 ( .A(n4584), .B(sreg[1129]), .Z(n4588) );
  NAND U5684 ( .A(n4586), .B(n4585), .Z(n4587) );
  NAND U5685 ( .A(n4588), .B(n4587), .Z(n4606) );
  XOR U5686 ( .A(n4607), .B(n4606), .Z(c[1130]) );
  NANDN U5687 ( .A(n4590), .B(n4589), .Z(n4594) );
  OR U5688 ( .A(n4592), .B(n4591), .Z(n4593) );
  AND U5689 ( .A(n4594), .B(n4593), .Z(n4612) );
  XOR U5690 ( .A(a[109]), .B(n2191), .Z(n4616) );
  AND U5691 ( .A(a[111]), .B(b[0]), .Z(n4596) );
  XNOR U5692 ( .A(n4596), .B(n2175), .Z(n4598) );
  NANDN U5693 ( .A(b[0]), .B(a[110]), .Z(n4597) );
  NAND U5694 ( .A(n4598), .B(n4597), .Z(n4621) );
  AND U5695 ( .A(a[107]), .B(b[3]), .Z(n4620) );
  XOR U5696 ( .A(n4621), .B(n4620), .Z(n4623) );
  XOR U5697 ( .A(n4622), .B(n4623), .Z(n4611) );
  NANDN U5698 ( .A(n4600), .B(n4599), .Z(n4604) );
  OR U5699 ( .A(n4602), .B(n4601), .Z(n4603) );
  AND U5700 ( .A(n4604), .B(n4603), .Z(n4610) );
  XOR U5701 ( .A(n4611), .B(n4610), .Z(n4613) );
  XOR U5702 ( .A(n4612), .B(n4613), .Z(n4626) );
  XNOR U5703 ( .A(n4626), .B(sreg[1131]), .Z(n4628) );
  NANDN U5704 ( .A(n4605), .B(sreg[1130]), .Z(n4609) );
  NAND U5705 ( .A(n4607), .B(n4606), .Z(n4608) );
  NAND U5706 ( .A(n4609), .B(n4608), .Z(n4627) );
  XOR U5707 ( .A(n4628), .B(n4627), .Z(c[1131]) );
  NANDN U5708 ( .A(n4611), .B(n4610), .Z(n4615) );
  OR U5709 ( .A(n4613), .B(n4612), .Z(n4614) );
  AND U5710 ( .A(n4615), .B(n4614), .Z(n4633) );
  XOR U5711 ( .A(a[110]), .B(n2191), .Z(n4637) );
  AND U5712 ( .A(a[112]), .B(b[0]), .Z(n4617) );
  XNOR U5713 ( .A(n4617), .B(n2175), .Z(n4619) );
  NANDN U5714 ( .A(b[0]), .B(a[111]), .Z(n4618) );
  NAND U5715 ( .A(n4619), .B(n4618), .Z(n4642) );
  AND U5716 ( .A(a[108]), .B(b[3]), .Z(n4641) );
  XOR U5717 ( .A(n4642), .B(n4641), .Z(n4644) );
  XOR U5718 ( .A(n4643), .B(n4644), .Z(n4632) );
  NANDN U5719 ( .A(n4621), .B(n4620), .Z(n4625) );
  OR U5720 ( .A(n4623), .B(n4622), .Z(n4624) );
  AND U5721 ( .A(n4625), .B(n4624), .Z(n4631) );
  XOR U5722 ( .A(n4632), .B(n4631), .Z(n4634) );
  XOR U5723 ( .A(n4633), .B(n4634), .Z(n4647) );
  XNOR U5724 ( .A(n4647), .B(sreg[1132]), .Z(n4649) );
  NANDN U5725 ( .A(n4626), .B(sreg[1131]), .Z(n4630) );
  NAND U5726 ( .A(n4628), .B(n4627), .Z(n4629) );
  NAND U5727 ( .A(n4630), .B(n4629), .Z(n4648) );
  XOR U5728 ( .A(n4649), .B(n4648), .Z(c[1132]) );
  NANDN U5729 ( .A(n4632), .B(n4631), .Z(n4636) );
  OR U5730 ( .A(n4634), .B(n4633), .Z(n4635) );
  AND U5731 ( .A(n4636), .B(n4635), .Z(n4654) );
  XOR U5732 ( .A(a[111]), .B(n2192), .Z(n4658) );
  AND U5733 ( .A(a[109]), .B(b[3]), .Z(n4662) );
  AND U5734 ( .A(a[113]), .B(b[0]), .Z(n4638) );
  XNOR U5735 ( .A(n4638), .B(n2175), .Z(n4640) );
  NANDN U5736 ( .A(b[0]), .B(a[112]), .Z(n4639) );
  NAND U5737 ( .A(n4640), .B(n4639), .Z(n4663) );
  XOR U5738 ( .A(n4662), .B(n4663), .Z(n4665) );
  XOR U5739 ( .A(n4664), .B(n4665), .Z(n4653) );
  NANDN U5740 ( .A(n4642), .B(n4641), .Z(n4646) );
  OR U5741 ( .A(n4644), .B(n4643), .Z(n4645) );
  AND U5742 ( .A(n4646), .B(n4645), .Z(n4652) );
  XOR U5743 ( .A(n4653), .B(n4652), .Z(n4655) );
  XOR U5744 ( .A(n4654), .B(n4655), .Z(n4668) );
  XNOR U5745 ( .A(n4668), .B(sreg[1133]), .Z(n4670) );
  NANDN U5746 ( .A(n4647), .B(sreg[1132]), .Z(n4651) );
  NAND U5747 ( .A(n4649), .B(n4648), .Z(n4650) );
  NAND U5748 ( .A(n4651), .B(n4650), .Z(n4669) );
  XOR U5749 ( .A(n4670), .B(n4669), .Z(c[1133]) );
  NANDN U5750 ( .A(n4653), .B(n4652), .Z(n4657) );
  OR U5751 ( .A(n4655), .B(n4654), .Z(n4656) );
  AND U5752 ( .A(n4657), .B(n4656), .Z(n4675) );
  XOR U5753 ( .A(a[112]), .B(n2192), .Z(n4679) );
  AND U5754 ( .A(a[114]), .B(b[0]), .Z(n4659) );
  XNOR U5755 ( .A(n4659), .B(n2175), .Z(n4661) );
  NANDN U5756 ( .A(b[0]), .B(a[113]), .Z(n4660) );
  NAND U5757 ( .A(n4661), .B(n4660), .Z(n4684) );
  AND U5758 ( .A(a[110]), .B(b[3]), .Z(n4683) );
  XOR U5759 ( .A(n4684), .B(n4683), .Z(n4686) );
  XOR U5760 ( .A(n4685), .B(n4686), .Z(n4674) );
  NANDN U5761 ( .A(n4663), .B(n4662), .Z(n4667) );
  OR U5762 ( .A(n4665), .B(n4664), .Z(n4666) );
  AND U5763 ( .A(n4667), .B(n4666), .Z(n4673) );
  XOR U5764 ( .A(n4674), .B(n4673), .Z(n4676) );
  XOR U5765 ( .A(n4675), .B(n4676), .Z(n4689) );
  XNOR U5766 ( .A(n4689), .B(sreg[1134]), .Z(n4691) );
  NANDN U5767 ( .A(n4668), .B(sreg[1133]), .Z(n4672) );
  NAND U5768 ( .A(n4670), .B(n4669), .Z(n4671) );
  NAND U5769 ( .A(n4672), .B(n4671), .Z(n4690) );
  XOR U5770 ( .A(n4691), .B(n4690), .Z(c[1134]) );
  NANDN U5771 ( .A(n4674), .B(n4673), .Z(n4678) );
  OR U5772 ( .A(n4676), .B(n4675), .Z(n4677) );
  AND U5773 ( .A(n4678), .B(n4677), .Z(n4696) );
  XOR U5774 ( .A(a[113]), .B(n2192), .Z(n4700) );
  AND U5775 ( .A(a[115]), .B(b[0]), .Z(n4680) );
  XNOR U5776 ( .A(n4680), .B(n2175), .Z(n4682) );
  NANDN U5777 ( .A(b[0]), .B(a[114]), .Z(n4681) );
  NAND U5778 ( .A(n4682), .B(n4681), .Z(n4705) );
  AND U5779 ( .A(a[111]), .B(b[3]), .Z(n4704) );
  XOR U5780 ( .A(n4705), .B(n4704), .Z(n4707) );
  XOR U5781 ( .A(n4706), .B(n4707), .Z(n4695) );
  NANDN U5782 ( .A(n4684), .B(n4683), .Z(n4688) );
  OR U5783 ( .A(n4686), .B(n4685), .Z(n4687) );
  AND U5784 ( .A(n4688), .B(n4687), .Z(n4694) );
  XOR U5785 ( .A(n4695), .B(n4694), .Z(n4697) );
  XOR U5786 ( .A(n4696), .B(n4697), .Z(n4710) );
  XNOR U5787 ( .A(n4710), .B(sreg[1135]), .Z(n4712) );
  NANDN U5788 ( .A(n4689), .B(sreg[1134]), .Z(n4693) );
  NAND U5789 ( .A(n4691), .B(n4690), .Z(n4692) );
  NAND U5790 ( .A(n4693), .B(n4692), .Z(n4711) );
  XOR U5791 ( .A(n4712), .B(n4711), .Z(c[1135]) );
  NANDN U5792 ( .A(n4695), .B(n4694), .Z(n4699) );
  OR U5793 ( .A(n4697), .B(n4696), .Z(n4698) );
  AND U5794 ( .A(n4699), .B(n4698), .Z(n4717) );
  XOR U5795 ( .A(a[114]), .B(n2192), .Z(n4721) );
  AND U5796 ( .A(a[112]), .B(b[3]), .Z(n4725) );
  AND U5797 ( .A(a[116]), .B(b[0]), .Z(n4701) );
  XNOR U5798 ( .A(n4701), .B(n2175), .Z(n4703) );
  NANDN U5799 ( .A(b[0]), .B(a[115]), .Z(n4702) );
  NAND U5800 ( .A(n4703), .B(n4702), .Z(n4726) );
  XOR U5801 ( .A(n4725), .B(n4726), .Z(n4728) );
  XOR U5802 ( .A(n4727), .B(n4728), .Z(n4716) );
  NANDN U5803 ( .A(n4705), .B(n4704), .Z(n4709) );
  OR U5804 ( .A(n4707), .B(n4706), .Z(n4708) );
  AND U5805 ( .A(n4709), .B(n4708), .Z(n4715) );
  XOR U5806 ( .A(n4716), .B(n4715), .Z(n4718) );
  XOR U5807 ( .A(n4717), .B(n4718), .Z(n4731) );
  XNOR U5808 ( .A(n4731), .B(sreg[1136]), .Z(n4733) );
  NANDN U5809 ( .A(n4710), .B(sreg[1135]), .Z(n4714) );
  NAND U5810 ( .A(n4712), .B(n4711), .Z(n4713) );
  NAND U5811 ( .A(n4714), .B(n4713), .Z(n4732) );
  XOR U5812 ( .A(n4733), .B(n4732), .Z(c[1136]) );
  NANDN U5813 ( .A(n4716), .B(n4715), .Z(n4720) );
  OR U5814 ( .A(n4718), .B(n4717), .Z(n4719) );
  AND U5815 ( .A(n4720), .B(n4719), .Z(n4738) );
  XOR U5816 ( .A(a[115]), .B(n2192), .Z(n4742) );
  AND U5817 ( .A(a[117]), .B(b[0]), .Z(n4722) );
  XNOR U5818 ( .A(n4722), .B(n2175), .Z(n4724) );
  NANDN U5819 ( .A(b[0]), .B(a[116]), .Z(n4723) );
  NAND U5820 ( .A(n4724), .B(n4723), .Z(n4747) );
  AND U5821 ( .A(a[113]), .B(b[3]), .Z(n4746) );
  XOR U5822 ( .A(n4747), .B(n4746), .Z(n4749) );
  XOR U5823 ( .A(n4748), .B(n4749), .Z(n4737) );
  NANDN U5824 ( .A(n4726), .B(n4725), .Z(n4730) );
  OR U5825 ( .A(n4728), .B(n4727), .Z(n4729) );
  AND U5826 ( .A(n4730), .B(n4729), .Z(n4736) );
  XOR U5827 ( .A(n4737), .B(n4736), .Z(n4739) );
  XOR U5828 ( .A(n4738), .B(n4739), .Z(n4752) );
  XNOR U5829 ( .A(n4752), .B(sreg[1137]), .Z(n4754) );
  NANDN U5830 ( .A(n4731), .B(sreg[1136]), .Z(n4735) );
  NAND U5831 ( .A(n4733), .B(n4732), .Z(n4734) );
  NAND U5832 ( .A(n4735), .B(n4734), .Z(n4753) );
  XOR U5833 ( .A(n4754), .B(n4753), .Z(c[1137]) );
  NANDN U5834 ( .A(n4737), .B(n4736), .Z(n4741) );
  OR U5835 ( .A(n4739), .B(n4738), .Z(n4740) );
  AND U5836 ( .A(n4741), .B(n4740), .Z(n4759) );
  XOR U5837 ( .A(a[116]), .B(n2192), .Z(n4763) );
  AND U5838 ( .A(a[118]), .B(b[0]), .Z(n4743) );
  XNOR U5839 ( .A(n4743), .B(n2175), .Z(n4745) );
  NANDN U5840 ( .A(b[0]), .B(a[117]), .Z(n4744) );
  NAND U5841 ( .A(n4745), .B(n4744), .Z(n4768) );
  AND U5842 ( .A(a[114]), .B(b[3]), .Z(n4767) );
  XOR U5843 ( .A(n4768), .B(n4767), .Z(n4770) );
  XOR U5844 ( .A(n4769), .B(n4770), .Z(n4758) );
  NANDN U5845 ( .A(n4747), .B(n4746), .Z(n4751) );
  OR U5846 ( .A(n4749), .B(n4748), .Z(n4750) );
  AND U5847 ( .A(n4751), .B(n4750), .Z(n4757) );
  XOR U5848 ( .A(n4758), .B(n4757), .Z(n4760) );
  XOR U5849 ( .A(n4759), .B(n4760), .Z(n4773) );
  XNOR U5850 ( .A(n4773), .B(sreg[1138]), .Z(n4775) );
  NANDN U5851 ( .A(n4752), .B(sreg[1137]), .Z(n4756) );
  NAND U5852 ( .A(n4754), .B(n4753), .Z(n4755) );
  NAND U5853 ( .A(n4756), .B(n4755), .Z(n4774) );
  XOR U5854 ( .A(n4775), .B(n4774), .Z(c[1138]) );
  NANDN U5855 ( .A(n4758), .B(n4757), .Z(n4762) );
  OR U5856 ( .A(n4760), .B(n4759), .Z(n4761) );
  AND U5857 ( .A(n4762), .B(n4761), .Z(n4780) );
  XOR U5858 ( .A(a[117]), .B(n2192), .Z(n4784) );
  AND U5859 ( .A(a[119]), .B(b[0]), .Z(n4764) );
  XNOR U5860 ( .A(n4764), .B(n2175), .Z(n4766) );
  NANDN U5861 ( .A(b[0]), .B(a[118]), .Z(n4765) );
  NAND U5862 ( .A(n4766), .B(n4765), .Z(n4789) );
  AND U5863 ( .A(a[115]), .B(b[3]), .Z(n4788) );
  XOR U5864 ( .A(n4789), .B(n4788), .Z(n4791) );
  XOR U5865 ( .A(n4790), .B(n4791), .Z(n4779) );
  NANDN U5866 ( .A(n4768), .B(n4767), .Z(n4772) );
  OR U5867 ( .A(n4770), .B(n4769), .Z(n4771) );
  AND U5868 ( .A(n4772), .B(n4771), .Z(n4778) );
  XOR U5869 ( .A(n4779), .B(n4778), .Z(n4781) );
  XOR U5870 ( .A(n4780), .B(n4781), .Z(n4794) );
  XNOR U5871 ( .A(n4794), .B(sreg[1139]), .Z(n4796) );
  NANDN U5872 ( .A(n4773), .B(sreg[1138]), .Z(n4777) );
  NAND U5873 ( .A(n4775), .B(n4774), .Z(n4776) );
  NAND U5874 ( .A(n4777), .B(n4776), .Z(n4795) );
  XOR U5875 ( .A(n4796), .B(n4795), .Z(c[1139]) );
  NANDN U5876 ( .A(n4779), .B(n4778), .Z(n4783) );
  OR U5877 ( .A(n4781), .B(n4780), .Z(n4782) );
  AND U5878 ( .A(n4783), .B(n4782), .Z(n4801) );
  XOR U5879 ( .A(a[118]), .B(n2193), .Z(n4805) );
  AND U5880 ( .A(a[120]), .B(b[0]), .Z(n4785) );
  XNOR U5881 ( .A(n4785), .B(n2175), .Z(n4787) );
  NANDN U5882 ( .A(b[0]), .B(a[119]), .Z(n4786) );
  NAND U5883 ( .A(n4787), .B(n4786), .Z(n4810) );
  AND U5884 ( .A(a[116]), .B(b[3]), .Z(n4809) );
  XOR U5885 ( .A(n4810), .B(n4809), .Z(n4812) );
  XOR U5886 ( .A(n4811), .B(n4812), .Z(n4800) );
  NANDN U5887 ( .A(n4789), .B(n4788), .Z(n4793) );
  OR U5888 ( .A(n4791), .B(n4790), .Z(n4792) );
  AND U5889 ( .A(n4793), .B(n4792), .Z(n4799) );
  XOR U5890 ( .A(n4800), .B(n4799), .Z(n4802) );
  XOR U5891 ( .A(n4801), .B(n4802), .Z(n4815) );
  XNOR U5892 ( .A(n4815), .B(sreg[1140]), .Z(n4817) );
  NANDN U5893 ( .A(n4794), .B(sreg[1139]), .Z(n4798) );
  NAND U5894 ( .A(n4796), .B(n4795), .Z(n4797) );
  NAND U5895 ( .A(n4798), .B(n4797), .Z(n4816) );
  XOR U5896 ( .A(n4817), .B(n4816), .Z(c[1140]) );
  NANDN U5897 ( .A(n4800), .B(n4799), .Z(n4804) );
  OR U5898 ( .A(n4802), .B(n4801), .Z(n4803) );
  AND U5899 ( .A(n4804), .B(n4803), .Z(n4822) );
  XOR U5900 ( .A(a[119]), .B(n2193), .Z(n4826) );
  AND U5901 ( .A(a[121]), .B(b[0]), .Z(n4806) );
  XNOR U5902 ( .A(n4806), .B(n2175), .Z(n4808) );
  NANDN U5903 ( .A(b[0]), .B(a[120]), .Z(n4807) );
  NAND U5904 ( .A(n4808), .B(n4807), .Z(n4831) );
  AND U5905 ( .A(a[117]), .B(b[3]), .Z(n4830) );
  XOR U5906 ( .A(n4831), .B(n4830), .Z(n4833) );
  XOR U5907 ( .A(n4832), .B(n4833), .Z(n4821) );
  NANDN U5908 ( .A(n4810), .B(n4809), .Z(n4814) );
  OR U5909 ( .A(n4812), .B(n4811), .Z(n4813) );
  AND U5910 ( .A(n4814), .B(n4813), .Z(n4820) );
  XOR U5911 ( .A(n4821), .B(n4820), .Z(n4823) );
  XOR U5912 ( .A(n4822), .B(n4823), .Z(n4836) );
  XNOR U5913 ( .A(n4836), .B(sreg[1141]), .Z(n4838) );
  NANDN U5914 ( .A(n4815), .B(sreg[1140]), .Z(n4819) );
  NAND U5915 ( .A(n4817), .B(n4816), .Z(n4818) );
  NAND U5916 ( .A(n4819), .B(n4818), .Z(n4837) );
  XOR U5917 ( .A(n4838), .B(n4837), .Z(c[1141]) );
  NANDN U5918 ( .A(n4821), .B(n4820), .Z(n4825) );
  OR U5919 ( .A(n4823), .B(n4822), .Z(n4824) );
  AND U5920 ( .A(n4825), .B(n4824), .Z(n4843) );
  XOR U5921 ( .A(a[120]), .B(n2193), .Z(n4847) );
  AND U5922 ( .A(a[122]), .B(b[0]), .Z(n4827) );
  XNOR U5923 ( .A(n4827), .B(n2175), .Z(n4829) );
  NANDN U5924 ( .A(b[0]), .B(a[121]), .Z(n4828) );
  NAND U5925 ( .A(n4829), .B(n4828), .Z(n4852) );
  AND U5926 ( .A(a[118]), .B(b[3]), .Z(n4851) );
  XOR U5927 ( .A(n4852), .B(n4851), .Z(n4854) );
  XOR U5928 ( .A(n4853), .B(n4854), .Z(n4842) );
  NANDN U5929 ( .A(n4831), .B(n4830), .Z(n4835) );
  OR U5930 ( .A(n4833), .B(n4832), .Z(n4834) );
  AND U5931 ( .A(n4835), .B(n4834), .Z(n4841) );
  XOR U5932 ( .A(n4842), .B(n4841), .Z(n4844) );
  XOR U5933 ( .A(n4843), .B(n4844), .Z(n4857) );
  XNOR U5934 ( .A(n4857), .B(sreg[1142]), .Z(n4859) );
  NANDN U5935 ( .A(n4836), .B(sreg[1141]), .Z(n4840) );
  NAND U5936 ( .A(n4838), .B(n4837), .Z(n4839) );
  NAND U5937 ( .A(n4840), .B(n4839), .Z(n4858) );
  XOR U5938 ( .A(n4859), .B(n4858), .Z(c[1142]) );
  NANDN U5939 ( .A(n4842), .B(n4841), .Z(n4846) );
  OR U5940 ( .A(n4844), .B(n4843), .Z(n4845) );
  AND U5941 ( .A(n4846), .B(n4845), .Z(n4864) );
  XOR U5942 ( .A(a[121]), .B(n2193), .Z(n4868) );
  AND U5943 ( .A(a[123]), .B(b[0]), .Z(n4848) );
  XNOR U5944 ( .A(n4848), .B(n2175), .Z(n4850) );
  NANDN U5945 ( .A(b[0]), .B(a[122]), .Z(n4849) );
  NAND U5946 ( .A(n4850), .B(n4849), .Z(n4873) );
  AND U5947 ( .A(a[119]), .B(b[3]), .Z(n4872) );
  XOR U5948 ( .A(n4873), .B(n4872), .Z(n4875) );
  XOR U5949 ( .A(n4874), .B(n4875), .Z(n4863) );
  NANDN U5950 ( .A(n4852), .B(n4851), .Z(n4856) );
  OR U5951 ( .A(n4854), .B(n4853), .Z(n4855) );
  AND U5952 ( .A(n4856), .B(n4855), .Z(n4862) );
  XOR U5953 ( .A(n4863), .B(n4862), .Z(n4865) );
  XOR U5954 ( .A(n4864), .B(n4865), .Z(n4878) );
  XNOR U5955 ( .A(n4878), .B(sreg[1143]), .Z(n4880) );
  NANDN U5956 ( .A(n4857), .B(sreg[1142]), .Z(n4861) );
  NAND U5957 ( .A(n4859), .B(n4858), .Z(n4860) );
  NAND U5958 ( .A(n4861), .B(n4860), .Z(n4879) );
  XOR U5959 ( .A(n4880), .B(n4879), .Z(c[1143]) );
  NANDN U5960 ( .A(n4863), .B(n4862), .Z(n4867) );
  OR U5961 ( .A(n4865), .B(n4864), .Z(n4866) );
  AND U5962 ( .A(n4867), .B(n4866), .Z(n4885) );
  XOR U5963 ( .A(a[122]), .B(n2193), .Z(n4889) );
  AND U5964 ( .A(a[120]), .B(b[3]), .Z(n4893) );
  AND U5965 ( .A(a[124]), .B(b[0]), .Z(n4869) );
  XNOR U5966 ( .A(n4869), .B(n2175), .Z(n4871) );
  NANDN U5967 ( .A(b[0]), .B(a[123]), .Z(n4870) );
  NAND U5968 ( .A(n4871), .B(n4870), .Z(n4894) );
  XOR U5969 ( .A(n4893), .B(n4894), .Z(n4896) );
  XOR U5970 ( .A(n4895), .B(n4896), .Z(n4884) );
  NANDN U5971 ( .A(n4873), .B(n4872), .Z(n4877) );
  OR U5972 ( .A(n4875), .B(n4874), .Z(n4876) );
  AND U5973 ( .A(n4877), .B(n4876), .Z(n4883) );
  XOR U5974 ( .A(n4884), .B(n4883), .Z(n4886) );
  XOR U5975 ( .A(n4885), .B(n4886), .Z(n4899) );
  XNOR U5976 ( .A(n4899), .B(sreg[1144]), .Z(n4901) );
  NANDN U5977 ( .A(n4878), .B(sreg[1143]), .Z(n4882) );
  NAND U5978 ( .A(n4880), .B(n4879), .Z(n4881) );
  NAND U5979 ( .A(n4882), .B(n4881), .Z(n4900) );
  XOR U5980 ( .A(n4901), .B(n4900), .Z(c[1144]) );
  NANDN U5981 ( .A(n4884), .B(n4883), .Z(n4888) );
  OR U5982 ( .A(n4886), .B(n4885), .Z(n4887) );
  AND U5983 ( .A(n4888), .B(n4887), .Z(n4906) );
  XOR U5984 ( .A(a[123]), .B(n2193), .Z(n4910) );
  AND U5985 ( .A(a[125]), .B(b[0]), .Z(n4890) );
  XNOR U5986 ( .A(n4890), .B(n2175), .Z(n4892) );
  NANDN U5987 ( .A(b[0]), .B(a[124]), .Z(n4891) );
  NAND U5988 ( .A(n4892), .B(n4891), .Z(n4915) );
  AND U5989 ( .A(a[121]), .B(b[3]), .Z(n4914) );
  XOR U5990 ( .A(n4915), .B(n4914), .Z(n4917) );
  XOR U5991 ( .A(n4916), .B(n4917), .Z(n4905) );
  NANDN U5992 ( .A(n4894), .B(n4893), .Z(n4898) );
  OR U5993 ( .A(n4896), .B(n4895), .Z(n4897) );
  AND U5994 ( .A(n4898), .B(n4897), .Z(n4904) );
  XOR U5995 ( .A(n4905), .B(n4904), .Z(n4907) );
  XOR U5996 ( .A(n4906), .B(n4907), .Z(n4920) );
  XNOR U5997 ( .A(n4920), .B(sreg[1145]), .Z(n4922) );
  NANDN U5998 ( .A(n4899), .B(sreg[1144]), .Z(n4903) );
  NAND U5999 ( .A(n4901), .B(n4900), .Z(n4902) );
  NAND U6000 ( .A(n4903), .B(n4902), .Z(n4921) );
  XOR U6001 ( .A(n4922), .B(n4921), .Z(c[1145]) );
  NANDN U6002 ( .A(n4905), .B(n4904), .Z(n4909) );
  OR U6003 ( .A(n4907), .B(n4906), .Z(n4908) );
  AND U6004 ( .A(n4909), .B(n4908), .Z(n4927) );
  XOR U6005 ( .A(a[124]), .B(n2193), .Z(n4931) );
  AND U6006 ( .A(a[122]), .B(b[3]), .Z(n4935) );
  AND U6007 ( .A(a[126]), .B(b[0]), .Z(n4911) );
  XNOR U6008 ( .A(n4911), .B(n2175), .Z(n4913) );
  NANDN U6009 ( .A(b[0]), .B(a[125]), .Z(n4912) );
  NAND U6010 ( .A(n4913), .B(n4912), .Z(n4936) );
  XOR U6011 ( .A(n4935), .B(n4936), .Z(n4938) );
  XOR U6012 ( .A(n4937), .B(n4938), .Z(n4926) );
  NANDN U6013 ( .A(n4915), .B(n4914), .Z(n4919) );
  OR U6014 ( .A(n4917), .B(n4916), .Z(n4918) );
  AND U6015 ( .A(n4919), .B(n4918), .Z(n4925) );
  XOR U6016 ( .A(n4926), .B(n4925), .Z(n4928) );
  XOR U6017 ( .A(n4927), .B(n4928), .Z(n4941) );
  XNOR U6018 ( .A(n4941), .B(sreg[1146]), .Z(n4943) );
  NANDN U6019 ( .A(n4920), .B(sreg[1145]), .Z(n4924) );
  NAND U6020 ( .A(n4922), .B(n4921), .Z(n4923) );
  NAND U6021 ( .A(n4924), .B(n4923), .Z(n4942) );
  XOR U6022 ( .A(n4943), .B(n4942), .Z(c[1146]) );
  NANDN U6023 ( .A(n4926), .B(n4925), .Z(n4930) );
  OR U6024 ( .A(n4928), .B(n4927), .Z(n4929) );
  AND U6025 ( .A(n4930), .B(n4929), .Z(n4948) );
  XOR U6026 ( .A(a[125]), .B(n2194), .Z(n4952) );
  AND U6027 ( .A(a[123]), .B(b[3]), .Z(n4956) );
  AND U6028 ( .A(a[127]), .B(b[0]), .Z(n4932) );
  XNOR U6029 ( .A(n4932), .B(n2175), .Z(n4934) );
  NANDN U6030 ( .A(b[0]), .B(a[126]), .Z(n4933) );
  NAND U6031 ( .A(n4934), .B(n4933), .Z(n4957) );
  XOR U6032 ( .A(n4956), .B(n4957), .Z(n4959) );
  XOR U6033 ( .A(n4958), .B(n4959), .Z(n4947) );
  NANDN U6034 ( .A(n4936), .B(n4935), .Z(n4940) );
  OR U6035 ( .A(n4938), .B(n4937), .Z(n4939) );
  AND U6036 ( .A(n4940), .B(n4939), .Z(n4946) );
  XOR U6037 ( .A(n4947), .B(n4946), .Z(n4949) );
  XOR U6038 ( .A(n4948), .B(n4949), .Z(n4962) );
  XNOR U6039 ( .A(n4962), .B(sreg[1147]), .Z(n4964) );
  NANDN U6040 ( .A(n4941), .B(sreg[1146]), .Z(n4945) );
  NAND U6041 ( .A(n4943), .B(n4942), .Z(n4944) );
  NAND U6042 ( .A(n4945), .B(n4944), .Z(n4963) );
  XOR U6043 ( .A(n4964), .B(n4963), .Z(c[1147]) );
  NANDN U6044 ( .A(n4947), .B(n4946), .Z(n4951) );
  OR U6045 ( .A(n4949), .B(n4948), .Z(n4950) );
  AND U6046 ( .A(n4951), .B(n4950), .Z(n4969) );
  XOR U6047 ( .A(a[126]), .B(n2194), .Z(n4973) );
  AND U6048 ( .A(a[124]), .B(b[3]), .Z(n4977) );
  AND U6049 ( .A(a[128]), .B(b[0]), .Z(n4953) );
  XNOR U6050 ( .A(n4953), .B(n2175), .Z(n4955) );
  NANDN U6051 ( .A(b[0]), .B(a[127]), .Z(n4954) );
  NAND U6052 ( .A(n4955), .B(n4954), .Z(n4978) );
  XOR U6053 ( .A(n4977), .B(n4978), .Z(n4980) );
  XOR U6054 ( .A(n4979), .B(n4980), .Z(n4968) );
  NANDN U6055 ( .A(n4957), .B(n4956), .Z(n4961) );
  OR U6056 ( .A(n4959), .B(n4958), .Z(n4960) );
  AND U6057 ( .A(n4961), .B(n4960), .Z(n4967) );
  XOR U6058 ( .A(n4968), .B(n4967), .Z(n4970) );
  XOR U6059 ( .A(n4969), .B(n4970), .Z(n4983) );
  XNOR U6060 ( .A(n4983), .B(sreg[1148]), .Z(n4985) );
  NANDN U6061 ( .A(n4962), .B(sreg[1147]), .Z(n4966) );
  NAND U6062 ( .A(n4964), .B(n4963), .Z(n4965) );
  NAND U6063 ( .A(n4966), .B(n4965), .Z(n4984) );
  XOR U6064 ( .A(n4985), .B(n4984), .Z(c[1148]) );
  NANDN U6065 ( .A(n4968), .B(n4967), .Z(n4972) );
  OR U6066 ( .A(n4970), .B(n4969), .Z(n4971) );
  AND U6067 ( .A(n4972), .B(n4971), .Z(n4990) );
  XOR U6068 ( .A(a[127]), .B(n2194), .Z(n4994) );
  AND U6069 ( .A(a[129]), .B(b[0]), .Z(n4974) );
  XNOR U6070 ( .A(n4974), .B(n2175), .Z(n4976) );
  NANDN U6071 ( .A(b[0]), .B(a[128]), .Z(n4975) );
  NAND U6072 ( .A(n4976), .B(n4975), .Z(n4999) );
  AND U6073 ( .A(a[125]), .B(b[3]), .Z(n4998) );
  XOR U6074 ( .A(n4999), .B(n4998), .Z(n5001) );
  XOR U6075 ( .A(n5000), .B(n5001), .Z(n4989) );
  NANDN U6076 ( .A(n4978), .B(n4977), .Z(n4982) );
  OR U6077 ( .A(n4980), .B(n4979), .Z(n4981) );
  AND U6078 ( .A(n4982), .B(n4981), .Z(n4988) );
  XOR U6079 ( .A(n4989), .B(n4988), .Z(n4991) );
  XOR U6080 ( .A(n4990), .B(n4991), .Z(n5004) );
  XNOR U6081 ( .A(n5004), .B(sreg[1149]), .Z(n5006) );
  NANDN U6082 ( .A(n4983), .B(sreg[1148]), .Z(n4987) );
  NAND U6083 ( .A(n4985), .B(n4984), .Z(n4986) );
  NAND U6084 ( .A(n4987), .B(n4986), .Z(n5005) );
  XOR U6085 ( .A(n5006), .B(n5005), .Z(c[1149]) );
  NANDN U6086 ( .A(n4989), .B(n4988), .Z(n4993) );
  OR U6087 ( .A(n4991), .B(n4990), .Z(n4992) );
  AND U6088 ( .A(n4993), .B(n4992), .Z(n5011) );
  XOR U6089 ( .A(a[128]), .B(n2194), .Z(n5015) );
  AND U6090 ( .A(a[130]), .B(b[0]), .Z(n4995) );
  XNOR U6091 ( .A(n4995), .B(n2175), .Z(n4997) );
  NANDN U6092 ( .A(b[0]), .B(a[129]), .Z(n4996) );
  NAND U6093 ( .A(n4997), .B(n4996), .Z(n5020) );
  AND U6094 ( .A(a[126]), .B(b[3]), .Z(n5019) );
  XOR U6095 ( .A(n5020), .B(n5019), .Z(n5022) );
  XOR U6096 ( .A(n5021), .B(n5022), .Z(n5010) );
  NANDN U6097 ( .A(n4999), .B(n4998), .Z(n5003) );
  OR U6098 ( .A(n5001), .B(n5000), .Z(n5002) );
  AND U6099 ( .A(n5003), .B(n5002), .Z(n5009) );
  XOR U6100 ( .A(n5010), .B(n5009), .Z(n5012) );
  XOR U6101 ( .A(n5011), .B(n5012), .Z(n5025) );
  XNOR U6102 ( .A(n5025), .B(sreg[1150]), .Z(n5027) );
  NANDN U6103 ( .A(n5004), .B(sreg[1149]), .Z(n5008) );
  NAND U6104 ( .A(n5006), .B(n5005), .Z(n5007) );
  NAND U6105 ( .A(n5008), .B(n5007), .Z(n5026) );
  XOR U6106 ( .A(n5027), .B(n5026), .Z(c[1150]) );
  NANDN U6107 ( .A(n5010), .B(n5009), .Z(n5014) );
  OR U6108 ( .A(n5012), .B(n5011), .Z(n5013) );
  AND U6109 ( .A(n5014), .B(n5013), .Z(n5032) );
  XOR U6110 ( .A(a[129]), .B(n2194), .Z(n5036) );
  AND U6111 ( .A(a[127]), .B(b[3]), .Z(n5040) );
  AND U6112 ( .A(a[131]), .B(b[0]), .Z(n5016) );
  XNOR U6113 ( .A(n5016), .B(n2175), .Z(n5018) );
  NANDN U6114 ( .A(b[0]), .B(a[130]), .Z(n5017) );
  NAND U6115 ( .A(n5018), .B(n5017), .Z(n5041) );
  XOR U6116 ( .A(n5040), .B(n5041), .Z(n5043) );
  XOR U6117 ( .A(n5042), .B(n5043), .Z(n5031) );
  NANDN U6118 ( .A(n5020), .B(n5019), .Z(n5024) );
  OR U6119 ( .A(n5022), .B(n5021), .Z(n5023) );
  AND U6120 ( .A(n5024), .B(n5023), .Z(n5030) );
  XOR U6121 ( .A(n5031), .B(n5030), .Z(n5033) );
  XOR U6122 ( .A(n5032), .B(n5033), .Z(n5046) );
  XNOR U6123 ( .A(n5046), .B(sreg[1151]), .Z(n5048) );
  NANDN U6124 ( .A(n5025), .B(sreg[1150]), .Z(n5029) );
  NAND U6125 ( .A(n5027), .B(n5026), .Z(n5028) );
  NAND U6126 ( .A(n5029), .B(n5028), .Z(n5047) );
  XOR U6127 ( .A(n5048), .B(n5047), .Z(c[1151]) );
  NANDN U6128 ( .A(n5031), .B(n5030), .Z(n5035) );
  OR U6129 ( .A(n5033), .B(n5032), .Z(n5034) );
  AND U6130 ( .A(n5035), .B(n5034), .Z(n5053) );
  XOR U6131 ( .A(a[130]), .B(n2194), .Z(n5057) );
  AND U6132 ( .A(a[132]), .B(b[0]), .Z(n5037) );
  XNOR U6133 ( .A(n5037), .B(n2175), .Z(n5039) );
  NANDN U6134 ( .A(b[0]), .B(a[131]), .Z(n5038) );
  NAND U6135 ( .A(n5039), .B(n5038), .Z(n5062) );
  AND U6136 ( .A(a[128]), .B(b[3]), .Z(n5061) );
  XOR U6137 ( .A(n5062), .B(n5061), .Z(n5064) );
  XOR U6138 ( .A(n5063), .B(n5064), .Z(n5052) );
  NANDN U6139 ( .A(n5041), .B(n5040), .Z(n5045) );
  OR U6140 ( .A(n5043), .B(n5042), .Z(n5044) );
  AND U6141 ( .A(n5045), .B(n5044), .Z(n5051) );
  XOR U6142 ( .A(n5052), .B(n5051), .Z(n5054) );
  XOR U6143 ( .A(n5053), .B(n5054), .Z(n5067) );
  XNOR U6144 ( .A(n5067), .B(sreg[1152]), .Z(n5069) );
  NANDN U6145 ( .A(n5046), .B(sreg[1151]), .Z(n5050) );
  NAND U6146 ( .A(n5048), .B(n5047), .Z(n5049) );
  NAND U6147 ( .A(n5050), .B(n5049), .Z(n5068) );
  XOR U6148 ( .A(n5069), .B(n5068), .Z(c[1152]) );
  NANDN U6149 ( .A(n5052), .B(n5051), .Z(n5056) );
  OR U6150 ( .A(n5054), .B(n5053), .Z(n5055) );
  AND U6151 ( .A(n5056), .B(n5055), .Z(n5074) );
  XOR U6152 ( .A(a[131]), .B(n2194), .Z(n5078) );
  AND U6153 ( .A(a[133]), .B(b[0]), .Z(n5058) );
  XNOR U6154 ( .A(n5058), .B(n2175), .Z(n5060) );
  NANDN U6155 ( .A(b[0]), .B(a[132]), .Z(n5059) );
  NAND U6156 ( .A(n5060), .B(n5059), .Z(n5083) );
  AND U6157 ( .A(a[129]), .B(b[3]), .Z(n5082) );
  XOR U6158 ( .A(n5083), .B(n5082), .Z(n5085) );
  XOR U6159 ( .A(n5084), .B(n5085), .Z(n5073) );
  NANDN U6160 ( .A(n5062), .B(n5061), .Z(n5066) );
  OR U6161 ( .A(n5064), .B(n5063), .Z(n5065) );
  AND U6162 ( .A(n5066), .B(n5065), .Z(n5072) );
  XOR U6163 ( .A(n5073), .B(n5072), .Z(n5075) );
  XOR U6164 ( .A(n5074), .B(n5075), .Z(n5088) );
  XNOR U6165 ( .A(n5088), .B(sreg[1153]), .Z(n5090) );
  NANDN U6166 ( .A(n5067), .B(sreg[1152]), .Z(n5071) );
  NAND U6167 ( .A(n5069), .B(n5068), .Z(n5070) );
  NAND U6168 ( .A(n5071), .B(n5070), .Z(n5089) );
  XOR U6169 ( .A(n5090), .B(n5089), .Z(c[1153]) );
  NANDN U6170 ( .A(n5073), .B(n5072), .Z(n5077) );
  OR U6171 ( .A(n5075), .B(n5074), .Z(n5076) );
  AND U6172 ( .A(n5077), .B(n5076), .Z(n5095) );
  XOR U6173 ( .A(a[132]), .B(n2195), .Z(n5099) );
  AND U6174 ( .A(a[134]), .B(b[0]), .Z(n5079) );
  XNOR U6175 ( .A(n5079), .B(n2175), .Z(n5081) );
  NANDN U6176 ( .A(b[0]), .B(a[133]), .Z(n5080) );
  NAND U6177 ( .A(n5081), .B(n5080), .Z(n5104) );
  AND U6178 ( .A(a[130]), .B(b[3]), .Z(n5103) );
  XOR U6179 ( .A(n5104), .B(n5103), .Z(n5106) );
  XOR U6180 ( .A(n5105), .B(n5106), .Z(n5094) );
  NANDN U6181 ( .A(n5083), .B(n5082), .Z(n5087) );
  OR U6182 ( .A(n5085), .B(n5084), .Z(n5086) );
  AND U6183 ( .A(n5087), .B(n5086), .Z(n5093) );
  XOR U6184 ( .A(n5094), .B(n5093), .Z(n5096) );
  XOR U6185 ( .A(n5095), .B(n5096), .Z(n5109) );
  XNOR U6186 ( .A(n5109), .B(sreg[1154]), .Z(n5111) );
  NANDN U6187 ( .A(n5088), .B(sreg[1153]), .Z(n5092) );
  NAND U6188 ( .A(n5090), .B(n5089), .Z(n5091) );
  NAND U6189 ( .A(n5092), .B(n5091), .Z(n5110) );
  XOR U6190 ( .A(n5111), .B(n5110), .Z(c[1154]) );
  NANDN U6191 ( .A(n5094), .B(n5093), .Z(n5098) );
  OR U6192 ( .A(n5096), .B(n5095), .Z(n5097) );
  AND U6193 ( .A(n5098), .B(n5097), .Z(n5116) );
  XOR U6194 ( .A(a[133]), .B(n2195), .Z(n5120) );
  AND U6195 ( .A(a[131]), .B(b[3]), .Z(n5124) );
  AND U6196 ( .A(a[135]), .B(b[0]), .Z(n5100) );
  XNOR U6197 ( .A(n5100), .B(n2175), .Z(n5102) );
  NANDN U6198 ( .A(b[0]), .B(a[134]), .Z(n5101) );
  NAND U6199 ( .A(n5102), .B(n5101), .Z(n5125) );
  XOR U6200 ( .A(n5124), .B(n5125), .Z(n5127) );
  XOR U6201 ( .A(n5126), .B(n5127), .Z(n5115) );
  NANDN U6202 ( .A(n5104), .B(n5103), .Z(n5108) );
  OR U6203 ( .A(n5106), .B(n5105), .Z(n5107) );
  AND U6204 ( .A(n5108), .B(n5107), .Z(n5114) );
  XOR U6205 ( .A(n5115), .B(n5114), .Z(n5117) );
  XOR U6206 ( .A(n5116), .B(n5117), .Z(n5130) );
  XNOR U6207 ( .A(n5130), .B(sreg[1155]), .Z(n5132) );
  NANDN U6208 ( .A(n5109), .B(sreg[1154]), .Z(n5113) );
  NAND U6209 ( .A(n5111), .B(n5110), .Z(n5112) );
  NAND U6210 ( .A(n5113), .B(n5112), .Z(n5131) );
  XOR U6211 ( .A(n5132), .B(n5131), .Z(c[1155]) );
  NANDN U6212 ( .A(n5115), .B(n5114), .Z(n5119) );
  OR U6213 ( .A(n5117), .B(n5116), .Z(n5118) );
  AND U6214 ( .A(n5119), .B(n5118), .Z(n5137) );
  XOR U6215 ( .A(a[134]), .B(n2195), .Z(n5141) );
  AND U6216 ( .A(a[136]), .B(b[0]), .Z(n5121) );
  XNOR U6217 ( .A(n5121), .B(n2175), .Z(n5123) );
  NANDN U6218 ( .A(b[0]), .B(a[135]), .Z(n5122) );
  NAND U6219 ( .A(n5123), .B(n5122), .Z(n5146) );
  AND U6220 ( .A(a[132]), .B(b[3]), .Z(n5145) );
  XOR U6221 ( .A(n5146), .B(n5145), .Z(n5148) );
  XOR U6222 ( .A(n5147), .B(n5148), .Z(n5136) );
  NANDN U6223 ( .A(n5125), .B(n5124), .Z(n5129) );
  OR U6224 ( .A(n5127), .B(n5126), .Z(n5128) );
  AND U6225 ( .A(n5129), .B(n5128), .Z(n5135) );
  XOR U6226 ( .A(n5136), .B(n5135), .Z(n5138) );
  XOR U6227 ( .A(n5137), .B(n5138), .Z(n5151) );
  XNOR U6228 ( .A(n5151), .B(sreg[1156]), .Z(n5153) );
  NANDN U6229 ( .A(n5130), .B(sreg[1155]), .Z(n5134) );
  NAND U6230 ( .A(n5132), .B(n5131), .Z(n5133) );
  NAND U6231 ( .A(n5134), .B(n5133), .Z(n5152) );
  XOR U6232 ( .A(n5153), .B(n5152), .Z(c[1156]) );
  NANDN U6233 ( .A(n5136), .B(n5135), .Z(n5140) );
  OR U6234 ( .A(n5138), .B(n5137), .Z(n5139) );
  AND U6235 ( .A(n5140), .B(n5139), .Z(n5158) );
  XOR U6236 ( .A(a[135]), .B(n2195), .Z(n5162) );
  AND U6237 ( .A(a[133]), .B(b[3]), .Z(n5166) );
  AND U6238 ( .A(a[137]), .B(b[0]), .Z(n5142) );
  XNOR U6239 ( .A(n5142), .B(n2175), .Z(n5144) );
  NANDN U6240 ( .A(b[0]), .B(a[136]), .Z(n5143) );
  NAND U6241 ( .A(n5144), .B(n5143), .Z(n5167) );
  XOR U6242 ( .A(n5166), .B(n5167), .Z(n5169) );
  XOR U6243 ( .A(n5168), .B(n5169), .Z(n5157) );
  NANDN U6244 ( .A(n5146), .B(n5145), .Z(n5150) );
  OR U6245 ( .A(n5148), .B(n5147), .Z(n5149) );
  AND U6246 ( .A(n5150), .B(n5149), .Z(n5156) );
  XOR U6247 ( .A(n5157), .B(n5156), .Z(n5159) );
  XOR U6248 ( .A(n5158), .B(n5159), .Z(n5172) );
  XNOR U6249 ( .A(n5172), .B(sreg[1157]), .Z(n5174) );
  NANDN U6250 ( .A(n5151), .B(sreg[1156]), .Z(n5155) );
  NAND U6251 ( .A(n5153), .B(n5152), .Z(n5154) );
  NAND U6252 ( .A(n5155), .B(n5154), .Z(n5173) );
  XOR U6253 ( .A(n5174), .B(n5173), .Z(c[1157]) );
  NANDN U6254 ( .A(n5157), .B(n5156), .Z(n5161) );
  OR U6255 ( .A(n5159), .B(n5158), .Z(n5160) );
  AND U6256 ( .A(n5161), .B(n5160), .Z(n5179) );
  XOR U6257 ( .A(a[136]), .B(n2195), .Z(n5183) );
  AND U6258 ( .A(a[134]), .B(b[3]), .Z(n5187) );
  AND U6259 ( .A(a[138]), .B(b[0]), .Z(n5163) );
  XNOR U6260 ( .A(n5163), .B(n2175), .Z(n5165) );
  NANDN U6261 ( .A(b[0]), .B(a[137]), .Z(n5164) );
  NAND U6262 ( .A(n5165), .B(n5164), .Z(n5188) );
  XOR U6263 ( .A(n5187), .B(n5188), .Z(n5190) );
  XOR U6264 ( .A(n5189), .B(n5190), .Z(n5178) );
  NANDN U6265 ( .A(n5167), .B(n5166), .Z(n5171) );
  OR U6266 ( .A(n5169), .B(n5168), .Z(n5170) );
  AND U6267 ( .A(n5171), .B(n5170), .Z(n5177) );
  XOR U6268 ( .A(n5178), .B(n5177), .Z(n5180) );
  XOR U6269 ( .A(n5179), .B(n5180), .Z(n5193) );
  XNOR U6270 ( .A(n5193), .B(sreg[1158]), .Z(n5195) );
  NANDN U6271 ( .A(n5172), .B(sreg[1157]), .Z(n5176) );
  NAND U6272 ( .A(n5174), .B(n5173), .Z(n5175) );
  NAND U6273 ( .A(n5176), .B(n5175), .Z(n5194) );
  XOR U6274 ( .A(n5195), .B(n5194), .Z(c[1158]) );
  NANDN U6275 ( .A(n5178), .B(n5177), .Z(n5182) );
  OR U6276 ( .A(n5180), .B(n5179), .Z(n5181) );
  AND U6277 ( .A(n5182), .B(n5181), .Z(n5200) );
  XOR U6278 ( .A(a[137]), .B(n2195), .Z(n5204) );
  AND U6279 ( .A(a[135]), .B(b[3]), .Z(n5208) );
  AND U6280 ( .A(a[139]), .B(b[0]), .Z(n5184) );
  XNOR U6281 ( .A(n5184), .B(n2175), .Z(n5186) );
  NANDN U6282 ( .A(b[0]), .B(a[138]), .Z(n5185) );
  NAND U6283 ( .A(n5186), .B(n5185), .Z(n5209) );
  XOR U6284 ( .A(n5208), .B(n5209), .Z(n5211) );
  XOR U6285 ( .A(n5210), .B(n5211), .Z(n5199) );
  NANDN U6286 ( .A(n5188), .B(n5187), .Z(n5192) );
  OR U6287 ( .A(n5190), .B(n5189), .Z(n5191) );
  AND U6288 ( .A(n5192), .B(n5191), .Z(n5198) );
  XOR U6289 ( .A(n5199), .B(n5198), .Z(n5201) );
  XOR U6290 ( .A(n5200), .B(n5201), .Z(n5214) );
  XNOR U6291 ( .A(n5214), .B(sreg[1159]), .Z(n5216) );
  NANDN U6292 ( .A(n5193), .B(sreg[1158]), .Z(n5197) );
  NAND U6293 ( .A(n5195), .B(n5194), .Z(n5196) );
  NAND U6294 ( .A(n5197), .B(n5196), .Z(n5215) );
  XOR U6295 ( .A(n5216), .B(n5215), .Z(c[1159]) );
  NANDN U6296 ( .A(n5199), .B(n5198), .Z(n5203) );
  OR U6297 ( .A(n5201), .B(n5200), .Z(n5202) );
  AND U6298 ( .A(n5203), .B(n5202), .Z(n5221) );
  XOR U6299 ( .A(a[138]), .B(n2195), .Z(n5225) );
  AND U6300 ( .A(a[140]), .B(b[0]), .Z(n5205) );
  XNOR U6301 ( .A(n5205), .B(n2175), .Z(n5207) );
  NANDN U6302 ( .A(b[0]), .B(a[139]), .Z(n5206) );
  NAND U6303 ( .A(n5207), .B(n5206), .Z(n5230) );
  AND U6304 ( .A(a[136]), .B(b[3]), .Z(n5229) );
  XOR U6305 ( .A(n5230), .B(n5229), .Z(n5232) );
  XOR U6306 ( .A(n5231), .B(n5232), .Z(n5220) );
  NANDN U6307 ( .A(n5209), .B(n5208), .Z(n5213) );
  OR U6308 ( .A(n5211), .B(n5210), .Z(n5212) );
  AND U6309 ( .A(n5213), .B(n5212), .Z(n5219) );
  XOR U6310 ( .A(n5220), .B(n5219), .Z(n5222) );
  XOR U6311 ( .A(n5221), .B(n5222), .Z(n5235) );
  XNOR U6312 ( .A(n5235), .B(sreg[1160]), .Z(n5237) );
  NANDN U6313 ( .A(n5214), .B(sreg[1159]), .Z(n5218) );
  NAND U6314 ( .A(n5216), .B(n5215), .Z(n5217) );
  NAND U6315 ( .A(n5218), .B(n5217), .Z(n5236) );
  XOR U6316 ( .A(n5237), .B(n5236), .Z(c[1160]) );
  NANDN U6317 ( .A(n5220), .B(n5219), .Z(n5224) );
  OR U6318 ( .A(n5222), .B(n5221), .Z(n5223) );
  AND U6319 ( .A(n5224), .B(n5223), .Z(n5242) );
  XOR U6320 ( .A(a[139]), .B(n2196), .Z(n5246) );
  AND U6321 ( .A(a[141]), .B(b[0]), .Z(n5226) );
  XNOR U6322 ( .A(n5226), .B(n2175), .Z(n5228) );
  NANDN U6323 ( .A(b[0]), .B(a[140]), .Z(n5227) );
  NAND U6324 ( .A(n5228), .B(n5227), .Z(n5251) );
  AND U6325 ( .A(a[137]), .B(b[3]), .Z(n5250) );
  XOR U6326 ( .A(n5251), .B(n5250), .Z(n5253) );
  XOR U6327 ( .A(n5252), .B(n5253), .Z(n5241) );
  NANDN U6328 ( .A(n5230), .B(n5229), .Z(n5234) );
  OR U6329 ( .A(n5232), .B(n5231), .Z(n5233) );
  AND U6330 ( .A(n5234), .B(n5233), .Z(n5240) );
  XOR U6331 ( .A(n5241), .B(n5240), .Z(n5243) );
  XOR U6332 ( .A(n5242), .B(n5243), .Z(n5256) );
  XNOR U6333 ( .A(n5256), .B(sreg[1161]), .Z(n5258) );
  NANDN U6334 ( .A(n5235), .B(sreg[1160]), .Z(n5239) );
  NAND U6335 ( .A(n5237), .B(n5236), .Z(n5238) );
  NAND U6336 ( .A(n5239), .B(n5238), .Z(n5257) );
  XOR U6337 ( .A(n5258), .B(n5257), .Z(c[1161]) );
  NANDN U6338 ( .A(n5241), .B(n5240), .Z(n5245) );
  OR U6339 ( .A(n5243), .B(n5242), .Z(n5244) );
  AND U6340 ( .A(n5245), .B(n5244), .Z(n5263) );
  XOR U6341 ( .A(a[140]), .B(n2196), .Z(n5267) );
  AND U6342 ( .A(a[138]), .B(b[3]), .Z(n5271) );
  AND U6343 ( .A(a[142]), .B(b[0]), .Z(n5247) );
  XNOR U6344 ( .A(n5247), .B(n2175), .Z(n5249) );
  NANDN U6345 ( .A(b[0]), .B(a[141]), .Z(n5248) );
  NAND U6346 ( .A(n5249), .B(n5248), .Z(n5272) );
  XOR U6347 ( .A(n5271), .B(n5272), .Z(n5274) );
  XOR U6348 ( .A(n5273), .B(n5274), .Z(n5262) );
  NANDN U6349 ( .A(n5251), .B(n5250), .Z(n5255) );
  OR U6350 ( .A(n5253), .B(n5252), .Z(n5254) );
  AND U6351 ( .A(n5255), .B(n5254), .Z(n5261) );
  XOR U6352 ( .A(n5262), .B(n5261), .Z(n5264) );
  XOR U6353 ( .A(n5263), .B(n5264), .Z(n5277) );
  XNOR U6354 ( .A(n5277), .B(sreg[1162]), .Z(n5279) );
  NANDN U6355 ( .A(n5256), .B(sreg[1161]), .Z(n5260) );
  NAND U6356 ( .A(n5258), .B(n5257), .Z(n5259) );
  NAND U6357 ( .A(n5260), .B(n5259), .Z(n5278) );
  XOR U6358 ( .A(n5279), .B(n5278), .Z(c[1162]) );
  NANDN U6359 ( .A(n5262), .B(n5261), .Z(n5266) );
  OR U6360 ( .A(n5264), .B(n5263), .Z(n5265) );
  AND U6361 ( .A(n5266), .B(n5265), .Z(n5284) );
  XOR U6362 ( .A(a[141]), .B(n2196), .Z(n5288) );
  AND U6363 ( .A(a[139]), .B(b[3]), .Z(n5292) );
  AND U6364 ( .A(a[143]), .B(b[0]), .Z(n5268) );
  XNOR U6365 ( .A(n5268), .B(n2175), .Z(n5270) );
  NANDN U6366 ( .A(b[0]), .B(a[142]), .Z(n5269) );
  NAND U6367 ( .A(n5270), .B(n5269), .Z(n5293) );
  XOR U6368 ( .A(n5292), .B(n5293), .Z(n5295) );
  XOR U6369 ( .A(n5294), .B(n5295), .Z(n5283) );
  NANDN U6370 ( .A(n5272), .B(n5271), .Z(n5276) );
  OR U6371 ( .A(n5274), .B(n5273), .Z(n5275) );
  AND U6372 ( .A(n5276), .B(n5275), .Z(n5282) );
  XOR U6373 ( .A(n5283), .B(n5282), .Z(n5285) );
  XOR U6374 ( .A(n5284), .B(n5285), .Z(n5298) );
  XNOR U6375 ( .A(n5298), .B(sreg[1163]), .Z(n5300) );
  NANDN U6376 ( .A(n5277), .B(sreg[1162]), .Z(n5281) );
  NAND U6377 ( .A(n5279), .B(n5278), .Z(n5280) );
  NAND U6378 ( .A(n5281), .B(n5280), .Z(n5299) );
  XOR U6379 ( .A(n5300), .B(n5299), .Z(c[1163]) );
  NANDN U6380 ( .A(n5283), .B(n5282), .Z(n5287) );
  OR U6381 ( .A(n5285), .B(n5284), .Z(n5286) );
  AND U6382 ( .A(n5287), .B(n5286), .Z(n5305) );
  XOR U6383 ( .A(a[142]), .B(n2196), .Z(n5309) );
  AND U6384 ( .A(a[144]), .B(b[0]), .Z(n5289) );
  XNOR U6385 ( .A(n5289), .B(n2175), .Z(n5291) );
  NANDN U6386 ( .A(b[0]), .B(a[143]), .Z(n5290) );
  NAND U6387 ( .A(n5291), .B(n5290), .Z(n5314) );
  AND U6388 ( .A(a[140]), .B(b[3]), .Z(n5313) );
  XOR U6389 ( .A(n5314), .B(n5313), .Z(n5316) );
  XOR U6390 ( .A(n5315), .B(n5316), .Z(n5304) );
  NANDN U6391 ( .A(n5293), .B(n5292), .Z(n5297) );
  OR U6392 ( .A(n5295), .B(n5294), .Z(n5296) );
  AND U6393 ( .A(n5297), .B(n5296), .Z(n5303) );
  XOR U6394 ( .A(n5304), .B(n5303), .Z(n5306) );
  XOR U6395 ( .A(n5305), .B(n5306), .Z(n5319) );
  XNOR U6396 ( .A(n5319), .B(sreg[1164]), .Z(n5321) );
  NANDN U6397 ( .A(n5298), .B(sreg[1163]), .Z(n5302) );
  NAND U6398 ( .A(n5300), .B(n5299), .Z(n5301) );
  NAND U6399 ( .A(n5302), .B(n5301), .Z(n5320) );
  XOR U6400 ( .A(n5321), .B(n5320), .Z(c[1164]) );
  NANDN U6401 ( .A(n5304), .B(n5303), .Z(n5308) );
  OR U6402 ( .A(n5306), .B(n5305), .Z(n5307) );
  AND U6403 ( .A(n5308), .B(n5307), .Z(n5326) );
  XOR U6404 ( .A(a[143]), .B(n2196), .Z(n5330) );
  AND U6405 ( .A(a[145]), .B(b[0]), .Z(n5310) );
  XNOR U6406 ( .A(n5310), .B(n2175), .Z(n5312) );
  NANDN U6407 ( .A(b[0]), .B(a[144]), .Z(n5311) );
  NAND U6408 ( .A(n5312), .B(n5311), .Z(n5335) );
  AND U6409 ( .A(a[141]), .B(b[3]), .Z(n5334) );
  XOR U6410 ( .A(n5335), .B(n5334), .Z(n5337) );
  XOR U6411 ( .A(n5336), .B(n5337), .Z(n5325) );
  NANDN U6412 ( .A(n5314), .B(n5313), .Z(n5318) );
  OR U6413 ( .A(n5316), .B(n5315), .Z(n5317) );
  AND U6414 ( .A(n5318), .B(n5317), .Z(n5324) );
  XOR U6415 ( .A(n5325), .B(n5324), .Z(n5327) );
  XOR U6416 ( .A(n5326), .B(n5327), .Z(n5340) );
  XNOR U6417 ( .A(n5340), .B(sreg[1165]), .Z(n5342) );
  NANDN U6418 ( .A(n5319), .B(sreg[1164]), .Z(n5323) );
  NAND U6419 ( .A(n5321), .B(n5320), .Z(n5322) );
  NAND U6420 ( .A(n5323), .B(n5322), .Z(n5341) );
  XOR U6421 ( .A(n5342), .B(n5341), .Z(c[1165]) );
  NANDN U6422 ( .A(n5325), .B(n5324), .Z(n5329) );
  OR U6423 ( .A(n5327), .B(n5326), .Z(n5328) );
  AND U6424 ( .A(n5329), .B(n5328), .Z(n5347) );
  XOR U6425 ( .A(a[144]), .B(n2196), .Z(n5351) );
  AND U6426 ( .A(a[146]), .B(b[0]), .Z(n5331) );
  XNOR U6427 ( .A(n5331), .B(n2175), .Z(n5333) );
  NANDN U6428 ( .A(b[0]), .B(a[145]), .Z(n5332) );
  NAND U6429 ( .A(n5333), .B(n5332), .Z(n5356) );
  AND U6430 ( .A(a[142]), .B(b[3]), .Z(n5355) );
  XOR U6431 ( .A(n5356), .B(n5355), .Z(n5358) );
  XOR U6432 ( .A(n5357), .B(n5358), .Z(n5346) );
  NANDN U6433 ( .A(n5335), .B(n5334), .Z(n5339) );
  OR U6434 ( .A(n5337), .B(n5336), .Z(n5338) );
  AND U6435 ( .A(n5339), .B(n5338), .Z(n5345) );
  XOR U6436 ( .A(n5346), .B(n5345), .Z(n5348) );
  XOR U6437 ( .A(n5347), .B(n5348), .Z(n5361) );
  XNOR U6438 ( .A(n5361), .B(sreg[1166]), .Z(n5363) );
  NANDN U6439 ( .A(n5340), .B(sreg[1165]), .Z(n5344) );
  NAND U6440 ( .A(n5342), .B(n5341), .Z(n5343) );
  NAND U6441 ( .A(n5344), .B(n5343), .Z(n5362) );
  XOR U6442 ( .A(n5363), .B(n5362), .Z(c[1166]) );
  NANDN U6443 ( .A(n5346), .B(n5345), .Z(n5350) );
  OR U6444 ( .A(n5348), .B(n5347), .Z(n5349) );
  AND U6445 ( .A(n5350), .B(n5349), .Z(n5368) );
  XOR U6446 ( .A(a[145]), .B(n2196), .Z(n5372) );
  AND U6447 ( .A(a[147]), .B(b[0]), .Z(n5352) );
  XNOR U6448 ( .A(n5352), .B(n2175), .Z(n5354) );
  NANDN U6449 ( .A(b[0]), .B(a[146]), .Z(n5353) );
  NAND U6450 ( .A(n5354), .B(n5353), .Z(n5377) );
  AND U6451 ( .A(a[143]), .B(b[3]), .Z(n5376) );
  XOR U6452 ( .A(n5377), .B(n5376), .Z(n5379) );
  XOR U6453 ( .A(n5378), .B(n5379), .Z(n5367) );
  NANDN U6454 ( .A(n5356), .B(n5355), .Z(n5360) );
  OR U6455 ( .A(n5358), .B(n5357), .Z(n5359) );
  AND U6456 ( .A(n5360), .B(n5359), .Z(n5366) );
  XOR U6457 ( .A(n5367), .B(n5366), .Z(n5369) );
  XOR U6458 ( .A(n5368), .B(n5369), .Z(n5382) );
  XNOR U6459 ( .A(n5382), .B(sreg[1167]), .Z(n5384) );
  NANDN U6460 ( .A(n5361), .B(sreg[1166]), .Z(n5365) );
  NAND U6461 ( .A(n5363), .B(n5362), .Z(n5364) );
  NAND U6462 ( .A(n5365), .B(n5364), .Z(n5383) );
  XOR U6463 ( .A(n5384), .B(n5383), .Z(c[1167]) );
  NANDN U6464 ( .A(n5367), .B(n5366), .Z(n5371) );
  OR U6465 ( .A(n5369), .B(n5368), .Z(n5370) );
  AND U6466 ( .A(n5371), .B(n5370), .Z(n5389) );
  XOR U6467 ( .A(a[146]), .B(n2197), .Z(n5393) );
  AND U6468 ( .A(a[148]), .B(b[0]), .Z(n5373) );
  XNOR U6469 ( .A(n5373), .B(n2175), .Z(n5375) );
  NANDN U6470 ( .A(b[0]), .B(a[147]), .Z(n5374) );
  NAND U6471 ( .A(n5375), .B(n5374), .Z(n5398) );
  AND U6472 ( .A(a[144]), .B(b[3]), .Z(n5397) );
  XOR U6473 ( .A(n5398), .B(n5397), .Z(n5400) );
  XOR U6474 ( .A(n5399), .B(n5400), .Z(n5388) );
  NANDN U6475 ( .A(n5377), .B(n5376), .Z(n5381) );
  OR U6476 ( .A(n5379), .B(n5378), .Z(n5380) );
  AND U6477 ( .A(n5381), .B(n5380), .Z(n5387) );
  XOR U6478 ( .A(n5388), .B(n5387), .Z(n5390) );
  XOR U6479 ( .A(n5389), .B(n5390), .Z(n5403) );
  XNOR U6480 ( .A(n5403), .B(sreg[1168]), .Z(n5405) );
  NANDN U6481 ( .A(n5382), .B(sreg[1167]), .Z(n5386) );
  NAND U6482 ( .A(n5384), .B(n5383), .Z(n5385) );
  NAND U6483 ( .A(n5386), .B(n5385), .Z(n5404) );
  XOR U6484 ( .A(n5405), .B(n5404), .Z(c[1168]) );
  NANDN U6485 ( .A(n5388), .B(n5387), .Z(n5392) );
  OR U6486 ( .A(n5390), .B(n5389), .Z(n5391) );
  AND U6487 ( .A(n5392), .B(n5391), .Z(n5410) );
  XOR U6488 ( .A(a[147]), .B(n2197), .Z(n5414) );
  AND U6489 ( .A(a[145]), .B(b[3]), .Z(n5418) );
  AND U6490 ( .A(a[149]), .B(b[0]), .Z(n5394) );
  XNOR U6491 ( .A(n5394), .B(n2175), .Z(n5396) );
  NANDN U6492 ( .A(b[0]), .B(a[148]), .Z(n5395) );
  NAND U6493 ( .A(n5396), .B(n5395), .Z(n5419) );
  XOR U6494 ( .A(n5418), .B(n5419), .Z(n5421) );
  XOR U6495 ( .A(n5420), .B(n5421), .Z(n5409) );
  NANDN U6496 ( .A(n5398), .B(n5397), .Z(n5402) );
  OR U6497 ( .A(n5400), .B(n5399), .Z(n5401) );
  AND U6498 ( .A(n5402), .B(n5401), .Z(n5408) );
  XOR U6499 ( .A(n5409), .B(n5408), .Z(n5411) );
  XOR U6500 ( .A(n5410), .B(n5411), .Z(n5424) );
  XNOR U6501 ( .A(n5424), .B(sreg[1169]), .Z(n5426) );
  NANDN U6502 ( .A(n5403), .B(sreg[1168]), .Z(n5407) );
  NAND U6503 ( .A(n5405), .B(n5404), .Z(n5406) );
  NAND U6504 ( .A(n5407), .B(n5406), .Z(n5425) );
  XOR U6505 ( .A(n5426), .B(n5425), .Z(c[1169]) );
  NANDN U6506 ( .A(n5409), .B(n5408), .Z(n5413) );
  OR U6507 ( .A(n5411), .B(n5410), .Z(n5412) );
  AND U6508 ( .A(n5413), .B(n5412), .Z(n5431) );
  XOR U6509 ( .A(a[148]), .B(n2197), .Z(n5435) );
  AND U6510 ( .A(a[150]), .B(b[0]), .Z(n5415) );
  XNOR U6511 ( .A(n5415), .B(n2175), .Z(n5417) );
  NANDN U6512 ( .A(b[0]), .B(a[149]), .Z(n5416) );
  NAND U6513 ( .A(n5417), .B(n5416), .Z(n5440) );
  AND U6514 ( .A(a[146]), .B(b[3]), .Z(n5439) );
  XOR U6515 ( .A(n5440), .B(n5439), .Z(n5442) );
  XOR U6516 ( .A(n5441), .B(n5442), .Z(n5430) );
  NANDN U6517 ( .A(n5419), .B(n5418), .Z(n5423) );
  OR U6518 ( .A(n5421), .B(n5420), .Z(n5422) );
  AND U6519 ( .A(n5423), .B(n5422), .Z(n5429) );
  XOR U6520 ( .A(n5430), .B(n5429), .Z(n5432) );
  XOR U6521 ( .A(n5431), .B(n5432), .Z(n5445) );
  XNOR U6522 ( .A(n5445), .B(sreg[1170]), .Z(n5447) );
  NANDN U6523 ( .A(n5424), .B(sreg[1169]), .Z(n5428) );
  NAND U6524 ( .A(n5426), .B(n5425), .Z(n5427) );
  NAND U6525 ( .A(n5428), .B(n5427), .Z(n5446) );
  XOR U6526 ( .A(n5447), .B(n5446), .Z(c[1170]) );
  NANDN U6527 ( .A(n5430), .B(n5429), .Z(n5434) );
  OR U6528 ( .A(n5432), .B(n5431), .Z(n5433) );
  AND U6529 ( .A(n5434), .B(n5433), .Z(n5452) );
  XOR U6530 ( .A(a[149]), .B(n2197), .Z(n5456) );
  AND U6531 ( .A(a[147]), .B(b[3]), .Z(n5460) );
  AND U6532 ( .A(a[151]), .B(b[0]), .Z(n5436) );
  XNOR U6533 ( .A(n5436), .B(n2175), .Z(n5438) );
  NANDN U6534 ( .A(b[0]), .B(a[150]), .Z(n5437) );
  NAND U6535 ( .A(n5438), .B(n5437), .Z(n5461) );
  XOR U6536 ( .A(n5460), .B(n5461), .Z(n5463) );
  XOR U6537 ( .A(n5462), .B(n5463), .Z(n5451) );
  NANDN U6538 ( .A(n5440), .B(n5439), .Z(n5444) );
  OR U6539 ( .A(n5442), .B(n5441), .Z(n5443) );
  AND U6540 ( .A(n5444), .B(n5443), .Z(n5450) );
  XOR U6541 ( .A(n5451), .B(n5450), .Z(n5453) );
  XOR U6542 ( .A(n5452), .B(n5453), .Z(n5466) );
  XNOR U6543 ( .A(n5466), .B(sreg[1171]), .Z(n5468) );
  NANDN U6544 ( .A(n5445), .B(sreg[1170]), .Z(n5449) );
  NAND U6545 ( .A(n5447), .B(n5446), .Z(n5448) );
  NAND U6546 ( .A(n5449), .B(n5448), .Z(n5467) );
  XOR U6547 ( .A(n5468), .B(n5467), .Z(c[1171]) );
  NANDN U6548 ( .A(n5451), .B(n5450), .Z(n5455) );
  OR U6549 ( .A(n5453), .B(n5452), .Z(n5454) );
  AND U6550 ( .A(n5455), .B(n5454), .Z(n5473) );
  XOR U6551 ( .A(a[150]), .B(n2197), .Z(n5477) );
  AND U6552 ( .A(a[152]), .B(b[0]), .Z(n5457) );
  XNOR U6553 ( .A(n5457), .B(n2175), .Z(n5459) );
  NANDN U6554 ( .A(b[0]), .B(a[151]), .Z(n5458) );
  NAND U6555 ( .A(n5459), .B(n5458), .Z(n5482) );
  AND U6556 ( .A(a[148]), .B(b[3]), .Z(n5481) );
  XOR U6557 ( .A(n5482), .B(n5481), .Z(n5484) );
  XOR U6558 ( .A(n5483), .B(n5484), .Z(n5472) );
  NANDN U6559 ( .A(n5461), .B(n5460), .Z(n5465) );
  OR U6560 ( .A(n5463), .B(n5462), .Z(n5464) );
  AND U6561 ( .A(n5465), .B(n5464), .Z(n5471) );
  XOR U6562 ( .A(n5472), .B(n5471), .Z(n5474) );
  XOR U6563 ( .A(n5473), .B(n5474), .Z(n5487) );
  XNOR U6564 ( .A(n5487), .B(sreg[1172]), .Z(n5489) );
  NANDN U6565 ( .A(n5466), .B(sreg[1171]), .Z(n5470) );
  NAND U6566 ( .A(n5468), .B(n5467), .Z(n5469) );
  NAND U6567 ( .A(n5470), .B(n5469), .Z(n5488) );
  XOR U6568 ( .A(n5489), .B(n5488), .Z(c[1172]) );
  NANDN U6569 ( .A(n5472), .B(n5471), .Z(n5476) );
  OR U6570 ( .A(n5474), .B(n5473), .Z(n5475) );
  AND U6571 ( .A(n5476), .B(n5475), .Z(n5494) );
  XOR U6572 ( .A(a[151]), .B(n2197), .Z(n5498) );
  AND U6573 ( .A(a[153]), .B(b[0]), .Z(n5478) );
  XNOR U6574 ( .A(n5478), .B(n2175), .Z(n5480) );
  NANDN U6575 ( .A(b[0]), .B(a[152]), .Z(n5479) );
  NAND U6576 ( .A(n5480), .B(n5479), .Z(n5503) );
  AND U6577 ( .A(a[149]), .B(b[3]), .Z(n5502) );
  XOR U6578 ( .A(n5503), .B(n5502), .Z(n5505) );
  XOR U6579 ( .A(n5504), .B(n5505), .Z(n5493) );
  NANDN U6580 ( .A(n5482), .B(n5481), .Z(n5486) );
  OR U6581 ( .A(n5484), .B(n5483), .Z(n5485) );
  AND U6582 ( .A(n5486), .B(n5485), .Z(n5492) );
  XOR U6583 ( .A(n5493), .B(n5492), .Z(n5495) );
  XOR U6584 ( .A(n5494), .B(n5495), .Z(n5508) );
  XNOR U6585 ( .A(n5508), .B(sreg[1173]), .Z(n5510) );
  NANDN U6586 ( .A(n5487), .B(sreg[1172]), .Z(n5491) );
  NAND U6587 ( .A(n5489), .B(n5488), .Z(n5490) );
  NAND U6588 ( .A(n5491), .B(n5490), .Z(n5509) );
  XOR U6589 ( .A(n5510), .B(n5509), .Z(c[1173]) );
  NANDN U6590 ( .A(n5493), .B(n5492), .Z(n5497) );
  OR U6591 ( .A(n5495), .B(n5494), .Z(n5496) );
  AND U6592 ( .A(n5497), .B(n5496), .Z(n5515) );
  XOR U6593 ( .A(a[152]), .B(n2197), .Z(n5519) );
  AND U6594 ( .A(a[154]), .B(b[0]), .Z(n5499) );
  XNOR U6595 ( .A(n5499), .B(n2175), .Z(n5501) );
  NANDN U6596 ( .A(b[0]), .B(a[153]), .Z(n5500) );
  NAND U6597 ( .A(n5501), .B(n5500), .Z(n5524) );
  AND U6598 ( .A(a[150]), .B(b[3]), .Z(n5523) );
  XOR U6599 ( .A(n5524), .B(n5523), .Z(n5526) );
  XOR U6600 ( .A(n5525), .B(n5526), .Z(n5514) );
  NANDN U6601 ( .A(n5503), .B(n5502), .Z(n5507) );
  OR U6602 ( .A(n5505), .B(n5504), .Z(n5506) );
  AND U6603 ( .A(n5507), .B(n5506), .Z(n5513) );
  XOR U6604 ( .A(n5514), .B(n5513), .Z(n5516) );
  XOR U6605 ( .A(n5515), .B(n5516), .Z(n5529) );
  XNOR U6606 ( .A(n5529), .B(sreg[1174]), .Z(n5531) );
  NANDN U6607 ( .A(n5508), .B(sreg[1173]), .Z(n5512) );
  NAND U6608 ( .A(n5510), .B(n5509), .Z(n5511) );
  NAND U6609 ( .A(n5512), .B(n5511), .Z(n5530) );
  XOR U6610 ( .A(n5531), .B(n5530), .Z(c[1174]) );
  NANDN U6611 ( .A(n5514), .B(n5513), .Z(n5518) );
  OR U6612 ( .A(n5516), .B(n5515), .Z(n5517) );
  AND U6613 ( .A(n5518), .B(n5517), .Z(n5536) );
  XOR U6614 ( .A(a[153]), .B(n2198), .Z(n5540) );
  AND U6615 ( .A(a[155]), .B(b[0]), .Z(n5520) );
  XNOR U6616 ( .A(n5520), .B(n2175), .Z(n5522) );
  NANDN U6617 ( .A(b[0]), .B(a[154]), .Z(n5521) );
  NAND U6618 ( .A(n5522), .B(n5521), .Z(n5545) );
  AND U6619 ( .A(a[151]), .B(b[3]), .Z(n5544) );
  XOR U6620 ( .A(n5545), .B(n5544), .Z(n5547) );
  XOR U6621 ( .A(n5546), .B(n5547), .Z(n5535) );
  NANDN U6622 ( .A(n5524), .B(n5523), .Z(n5528) );
  OR U6623 ( .A(n5526), .B(n5525), .Z(n5527) );
  AND U6624 ( .A(n5528), .B(n5527), .Z(n5534) );
  XOR U6625 ( .A(n5535), .B(n5534), .Z(n5537) );
  XOR U6626 ( .A(n5536), .B(n5537), .Z(n5550) );
  XNOR U6627 ( .A(n5550), .B(sreg[1175]), .Z(n5552) );
  NANDN U6628 ( .A(n5529), .B(sreg[1174]), .Z(n5533) );
  NAND U6629 ( .A(n5531), .B(n5530), .Z(n5532) );
  NAND U6630 ( .A(n5533), .B(n5532), .Z(n5551) );
  XOR U6631 ( .A(n5552), .B(n5551), .Z(c[1175]) );
  NANDN U6632 ( .A(n5535), .B(n5534), .Z(n5539) );
  OR U6633 ( .A(n5537), .B(n5536), .Z(n5538) );
  AND U6634 ( .A(n5539), .B(n5538), .Z(n5557) );
  XOR U6635 ( .A(a[154]), .B(n2198), .Z(n5561) );
  AND U6636 ( .A(a[152]), .B(b[3]), .Z(n5565) );
  AND U6637 ( .A(a[156]), .B(b[0]), .Z(n5541) );
  XNOR U6638 ( .A(n5541), .B(n2175), .Z(n5543) );
  NANDN U6639 ( .A(b[0]), .B(a[155]), .Z(n5542) );
  NAND U6640 ( .A(n5543), .B(n5542), .Z(n5566) );
  XOR U6641 ( .A(n5565), .B(n5566), .Z(n5568) );
  XOR U6642 ( .A(n5567), .B(n5568), .Z(n5556) );
  NANDN U6643 ( .A(n5545), .B(n5544), .Z(n5549) );
  OR U6644 ( .A(n5547), .B(n5546), .Z(n5548) );
  AND U6645 ( .A(n5549), .B(n5548), .Z(n5555) );
  XOR U6646 ( .A(n5556), .B(n5555), .Z(n5558) );
  XOR U6647 ( .A(n5557), .B(n5558), .Z(n5571) );
  XNOR U6648 ( .A(n5571), .B(sreg[1176]), .Z(n5573) );
  NANDN U6649 ( .A(n5550), .B(sreg[1175]), .Z(n5554) );
  NAND U6650 ( .A(n5552), .B(n5551), .Z(n5553) );
  NAND U6651 ( .A(n5554), .B(n5553), .Z(n5572) );
  XOR U6652 ( .A(n5573), .B(n5572), .Z(c[1176]) );
  NANDN U6653 ( .A(n5556), .B(n5555), .Z(n5560) );
  OR U6654 ( .A(n5558), .B(n5557), .Z(n5559) );
  AND U6655 ( .A(n5560), .B(n5559), .Z(n5578) );
  XOR U6656 ( .A(a[155]), .B(n2198), .Z(n5582) );
  AND U6657 ( .A(a[153]), .B(b[3]), .Z(n5586) );
  AND U6658 ( .A(a[157]), .B(b[0]), .Z(n5562) );
  XNOR U6659 ( .A(n5562), .B(n2175), .Z(n5564) );
  NANDN U6660 ( .A(b[0]), .B(a[156]), .Z(n5563) );
  NAND U6661 ( .A(n5564), .B(n5563), .Z(n5587) );
  XOR U6662 ( .A(n5586), .B(n5587), .Z(n5589) );
  XOR U6663 ( .A(n5588), .B(n5589), .Z(n5577) );
  NANDN U6664 ( .A(n5566), .B(n5565), .Z(n5570) );
  OR U6665 ( .A(n5568), .B(n5567), .Z(n5569) );
  AND U6666 ( .A(n5570), .B(n5569), .Z(n5576) );
  XOR U6667 ( .A(n5577), .B(n5576), .Z(n5579) );
  XOR U6668 ( .A(n5578), .B(n5579), .Z(n5592) );
  XNOR U6669 ( .A(n5592), .B(sreg[1177]), .Z(n5594) );
  NANDN U6670 ( .A(n5571), .B(sreg[1176]), .Z(n5575) );
  NAND U6671 ( .A(n5573), .B(n5572), .Z(n5574) );
  NAND U6672 ( .A(n5575), .B(n5574), .Z(n5593) );
  XOR U6673 ( .A(n5594), .B(n5593), .Z(c[1177]) );
  NANDN U6674 ( .A(n5577), .B(n5576), .Z(n5581) );
  OR U6675 ( .A(n5579), .B(n5578), .Z(n5580) );
  AND U6676 ( .A(n5581), .B(n5580), .Z(n5599) );
  XOR U6677 ( .A(a[156]), .B(n2198), .Z(n5603) );
  AND U6678 ( .A(a[158]), .B(b[0]), .Z(n5583) );
  XNOR U6679 ( .A(n5583), .B(n2175), .Z(n5585) );
  NANDN U6680 ( .A(b[0]), .B(a[157]), .Z(n5584) );
  NAND U6681 ( .A(n5585), .B(n5584), .Z(n5608) );
  AND U6682 ( .A(a[154]), .B(b[3]), .Z(n5607) );
  XOR U6683 ( .A(n5608), .B(n5607), .Z(n5610) );
  XOR U6684 ( .A(n5609), .B(n5610), .Z(n5598) );
  NANDN U6685 ( .A(n5587), .B(n5586), .Z(n5591) );
  OR U6686 ( .A(n5589), .B(n5588), .Z(n5590) );
  AND U6687 ( .A(n5591), .B(n5590), .Z(n5597) );
  XOR U6688 ( .A(n5598), .B(n5597), .Z(n5600) );
  XOR U6689 ( .A(n5599), .B(n5600), .Z(n5613) );
  XNOR U6690 ( .A(n5613), .B(sreg[1178]), .Z(n5615) );
  NANDN U6691 ( .A(n5592), .B(sreg[1177]), .Z(n5596) );
  NAND U6692 ( .A(n5594), .B(n5593), .Z(n5595) );
  NAND U6693 ( .A(n5596), .B(n5595), .Z(n5614) );
  XOR U6694 ( .A(n5615), .B(n5614), .Z(c[1178]) );
  NANDN U6695 ( .A(n5598), .B(n5597), .Z(n5602) );
  OR U6696 ( .A(n5600), .B(n5599), .Z(n5601) );
  AND U6697 ( .A(n5602), .B(n5601), .Z(n5620) );
  XOR U6698 ( .A(a[157]), .B(n2198), .Z(n5624) );
  AND U6699 ( .A(a[159]), .B(b[0]), .Z(n5604) );
  XNOR U6700 ( .A(n5604), .B(n2175), .Z(n5606) );
  NANDN U6701 ( .A(b[0]), .B(a[158]), .Z(n5605) );
  NAND U6702 ( .A(n5606), .B(n5605), .Z(n5629) );
  AND U6703 ( .A(a[155]), .B(b[3]), .Z(n5628) );
  XOR U6704 ( .A(n5629), .B(n5628), .Z(n5631) );
  XOR U6705 ( .A(n5630), .B(n5631), .Z(n5619) );
  NANDN U6706 ( .A(n5608), .B(n5607), .Z(n5612) );
  OR U6707 ( .A(n5610), .B(n5609), .Z(n5611) );
  AND U6708 ( .A(n5612), .B(n5611), .Z(n5618) );
  XOR U6709 ( .A(n5619), .B(n5618), .Z(n5621) );
  XOR U6710 ( .A(n5620), .B(n5621), .Z(n5634) );
  XNOR U6711 ( .A(n5634), .B(sreg[1179]), .Z(n5636) );
  NANDN U6712 ( .A(n5613), .B(sreg[1178]), .Z(n5617) );
  NAND U6713 ( .A(n5615), .B(n5614), .Z(n5616) );
  NAND U6714 ( .A(n5617), .B(n5616), .Z(n5635) );
  XOR U6715 ( .A(n5636), .B(n5635), .Z(c[1179]) );
  NANDN U6716 ( .A(n5619), .B(n5618), .Z(n5623) );
  OR U6717 ( .A(n5621), .B(n5620), .Z(n5622) );
  AND U6718 ( .A(n5623), .B(n5622), .Z(n5641) );
  XOR U6719 ( .A(a[158]), .B(n2198), .Z(n5645) );
  AND U6720 ( .A(a[160]), .B(b[0]), .Z(n5625) );
  XNOR U6721 ( .A(n5625), .B(n2175), .Z(n5627) );
  NANDN U6722 ( .A(b[0]), .B(a[159]), .Z(n5626) );
  NAND U6723 ( .A(n5627), .B(n5626), .Z(n5650) );
  AND U6724 ( .A(a[156]), .B(b[3]), .Z(n5649) );
  XOR U6725 ( .A(n5650), .B(n5649), .Z(n5652) );
  XOR U6726 ( .A(n5651), .B(n5652), .Z(n5640) );
  NANDN U6727 ( .A(n5629), .B(n5628), .Z(n5633) );
  OR U6728 ( .A(n5631), .B(n5630), .Z(n5632) );
  AND U6729 ( .A(n5633), .B(n5632), .Z(n5639) );
  XOR U6730 ( .A(n5640), .B(n5639), .Z(n5642) );
  XOR U6731 ( .A(n5641), .B(n5642), .Z(n5655) );
  XNOR U6732 ( .A(n5655), .B(sreg[1180]), .Z(n5657) );
  NANDN U6733 ( .A(n5634), .B(sreg[1179]), .Z(n5638) );
  NAND U6734 ( .A(n5636), .B(n5635), .Z(n5637) );
  NAND U6735 ( .A(n5638), .B(n5637), .Z(n5656) );
  XOR U6736 ( .A(n5657), .B(n5656), .Z(c[1180]) );
  NANDN U6737 ( .A(n5640), .B(n5639), .Z(n5644) );
  OR U6738 ( .A(n5642), .B(n5641), .Z(n5643) );
  AND U6739 ( .A(n5644), .B(n5643), .Z(n5662) );
  XOR U6740 ( .A(a[159]), .B(n2198), .Z(n5666) );
  AND U6741 ( .A(a[161]), .B(b[0]), .Z(n5646) );
  XNOR U6742 ( .A(n5646), .B(n2175), .Z(n5648) );
  NANDN U6743 ( .A(b[0]), .B(a[160]), .Z(n5647) );
  NAND U6744 ( .A(n5648), .B(n5647), .Z(n5671) );
  AND U6745 ( .A(a[157]), .B(b[3]), .Z(n5670) );
  XOR U6746 ( .A(n5671), .B(n5670), .Z(n5673) );
  XOR U6747 ( .A(n5672), .B(n5673), .Z(n5661) );
  NANDN U6748 ( .A(n5650), .B(n5649), .Z(n5654) );
  OR U6749 ( .A(n5652), .B(n5651), .Z(n5653) );
  AND U6750 ( .A(n5654), .B(n5653), .Z(n5660) );
  XOR U6751 ( .A(n5661), .B(n5660), .Z(n5663) );
  XOR U6752 ( .A(n5662), .B(n5663), .Z(n5676) );
  XNOR U6753 ( .A(n5676), .B(sreg[1181]), .Z(n5678) );
  NANDN U6754 ( .A(n5655), .B(sreg[1180]), .Z(n5659) );
  NAND U6755 ( .A(n5657), .B(n5656), .Z(n5658) );
  NAND U6756 ( .A(n5659), .B(n5658), .Z(n5677) );
  XOR U6757 ( .A(n5678), .B(n5677), .Z(c[1181]) );
  NANDN U6758 ( .A(n5661), .B(n5660), .Z(n5665) );
  OR U6759 ( .A(n5663), .B(n5662), .Z(n5664) );
  AND U6760 ( .A(n5665), .B(n5664), .Z(n5683) );
  XOR U6761 ( .A(a[160]), .B(n2199), .Z(n5687) );
  AND U6762 ( .A(a[162]), .B(b[0]), .Z(n5667) );
  XNOR U6763 ( .A(n5667), .B(n2175), .Z(n5669) );
  NANDN U6764 ( .A(b[0]), .B(a[161]), .Z(n5668) );
  NAND U6765 ( .A(n5669), .B(n5668), .Z(n5692) );
  AND U6766 ( .A(a[158]), .B(b[3]), .Z(n5691) );
  XOR U6767 ( .A(n5692), .B(n5691), .Z(n5694) );
  XOR U6768 ( .A(n5693), .B(n5694), .Z(n5682) );
  NANDN U6769 ( .A(n5671), .B(n5670), .Z(n5675) );
  OR U6770 ( .A(n5673), .B(n5672), .Z(n5674) );
  AND U6771 ( .A(n5675), .B(n5674), .Z(n5681) );
  XOR U6772 ( .A(n5682), .B(n5681), .Z(n5684) );
  XOR U6773 ( .A(n5683), .B(n5684), .Z(n5697) );
  XNOR U6774 ( .A(n5697), .B(sreg[1182]), .Z(n5699) );
  NANDN U6775 ( .A(n5676), .B(sreg[1181]), .Z(n5680) );
  NAND U6776 ( .A(n5678), .B(n5677), .Z(n5679) );
  NAND U6777 ( .A(n5680), .B(n5679), .Z(n5698) );
  XOR U6778 ( .A(n5699), .B(n5698), .Z(c[1182]) );
  NANDN U6779 ( .A(n5682), .B(n5681), .Z(n5686) );
  OR U6780 ( .A(n5684), .B(n5683), .Z(n5685) );
  AND U6781 ( .A(n5686), .B(n5685), .Z(n5704) );
  XOR U6782 ( .A(a[161]), .B(n2199), .Z(n5708) );
  AND U6783 ( .A(a[163]), .B(b[0]), .Z(n5688) );
  XNOR U6784 ( .A(n5688), .B(n2175), .Z(n5690) );
  NANDN U6785 ( .A(b[0]), .B(a[162]), .Z(n5689) );
  NAND U6786 ( .A(n5690), .B(n5689), .Z(n5713) );
  AND U6787 ( .A(a[159]), .B(b[3]), .Z(n5712) );
  XOR U6788 ( .A(n5713), .B(n5712), .Z(n5715) );
  XOR U6789 ( .A(n5714), .B(n5715), .Z(n5703) );
  NANDN U6790 ( .A(n5692), .B(n5691), .Z(n5696) );
  OR U6791 ( .A(n5694), .B(n5693), .Z(n5695) );
  AND U6792 ( .A(n5696), .B(n5695), .Z(n5702) );
  XOR U6793 ( .A(n5703), .B(n5702), .Z(n5705) );
  XOR U6794 ( .A(n5704), .B(n5705), .Z(n5718) );
  XNOR U6795 ( .A(n5718), .B(sreg[1183]), .Z(n5720) );
  NANDN U6796 ( .A(n5697), .B(sreg[1182]), .Z(n5701) );
  NAND U6797 ( .A(n5699), .B(n5698), .Z(n5700) );
  NAND U6798 ( .A(n5701), .B(n5700), .Z(n5719) );
  XOR U6799 ( .A(n5720), .B(n5719), .Z(c[1183]) );
  NANDN U6800 ( .A(n5703), .B(n5702), .Z(n5707) );
  OR U6801 ( .A(n5705), .B(n5704), .Z(n5706) );
  AND U6802 ( .A(n5707), .B(n5706), .Z(n5725) );
  XOR U6803 ( .A(a[162]), .B(n2199), .Z(n5729) );
  AND U6804 ( .A(a[164]), .B(b[0]), .Z(n5709) );
  XNOR U6805 ( .A(n5709), .B(n2175), .Z(n5711) );
  NANDN U6806 ( .A(b[0]), .B(a[163]), .Z(n5710) );
  NAND U6807 ( .A(n5711), .B(n5710), .Z(n5734) );
  AND U6808 ( .A(a[160]), .B(b[3]), .Z(n5733) );
  XOR U6809 ( .A(n5734), .B(n5733), .Z(n5736) );
  XOR U6810 ( .A(n5735), .B(n5736), .Z(n5724) );
  NANDN U6811 ( .A(n5713), .B(n5712), .Z(n5717) );
  OR U6812 ( .A(n5715), .B(n5714), .Z(n5716) );
  AND U6813 ( .A(n5717), .B(n5716), .Z(n5723) );
  XOR U6814 ( .A(n5724), .B(n5723), .Z(n5726) );
  XOR U6815 ( .A(n5725), .B(n5726), .Z(n5739) );
  XNOR U6816 ( .A(n5739), .B(sreg[1184]), .Z(n5741) );
  NANDN U6817 ( .A(n5718), .B(sreg[1183]), .Z(n5722) );
  NAND U6818 ( .A(n5720), .B(n5719), .Z(n5721) );
  NAND U6819 ( .A(n5722), .B(n5721), .Z(n5740) );
  XOR U6820 ( .A(n5741), .B(n5740), .Z(c[1184]) );
  NANDN U6821 ( .A(n5724), .B(n5723), .Z(n5728) );
  OR U6822 ( .A(n5726), .B(n5725), .Z(n5727) );
  AND U6823 ( .A(n5728), .B(n5727), .Z(n5746) );
  XOR U6824 ( .A(a[163]), .B(n2199), .Z(n5750) );
  AND U6825 ( .A(a[165]), .B(b[0]), .Z(n5730) );
  XNOR U6826 ( .A(n5730), .B(n2175), .Z(n5732) );
  NANDN U6827 ( .A(b[0]), .B(a[164]), .Z(n5731) );
  NAND U6828 ( .A(n5732), .B(n5731), .Z(n5755) );
  AND U6829 ( .A(a[161]), .B(b[3]), .Z(n5754) );
  XOR U6830 ( .A(n5755), .B(n5754), .Z(n5757) );
  XOR U6831 ( .A(n5756), .B(n5757), .Z(n5745) );
  NANDN U6832 ( .A(n5734), .B(n5733), .Z(n5738) );
  OR U6833 ( .A(n5736), .B(n5735), .Z(n5737) );
  AND U6834 ( .A(n5738), .B(n5737), .Z(n5744) );
  XOR U6835 ( .A(n5745), .B(n5744), .Z(n5747) );
  XOR U6836 ( .A(n5746), .B(n5747), .Z(n5760) );
  XNOR U6837 ( .A(n5760), .B(sreg[1185]), .Z(n5762) );
  NANDN U6838 ( .A(n5739), .B(sreg[1184]), .Z(n5743) );
  NAND U6839 ( .A(n5741), .B(n5740), .Z(n5742) );
  NAND U6840 ( .A(n5743), .B(n5742), .Z(n5761) );
  XOR U6841 ( .A(n5762), .B(n5761), .Z(c[1185]) );
  NANDN U6842 ( .A(n5745), .B(n5744), .Z(n5749) );
  OR U6843 ( .A(n5747), .B(n5746), .Z(n5748) );
  AND U6844 ( .A(n5749), .B(n5748), .Z(n5767) );
  XOR U6845 ( .A(a[164]), .B(n2199), .Z(n5771) );
  AND U6846 ( .A(a[166]), .B(b[0]), .Z(n5751) );
  XNOR U6847 ( .A(n5751), .B(n2175), .Z(n5753) );
  NANDN U6848 ( .A(b[0]), .B(a[165]), .Z(n5752) );
  NAND U6849 ( .A(n5753), .B(n5752), .Z(n5776) );
  AND U6850 ( .A(a[162]), .B(b[3]), .Z(n5775) );
  XOR U6851 ( .A(n5776), .B(n5775), .Z(n5778) );
  XOR U6852 ( .A(n5777), .B(n5778), .Z(n5766) );
  NANDN U6853 ( .A(n5755), .B(n5754), .Z(n5759) );
  OR U6854 ( .A(n5757), .B(n5756), .Z(n5758) );
  AND U6855 ( .A(n5759), .B(n5758), .Z(n5765) );
  XOR U6856 ( .A(n5766), .B(n5765), .Z(n5768) );
  XOR U6857 ( .A(n5767), .B(n5768), .Z(n5781) );
  XNOR U6858 ( .A(n5781), .B(sreg[1186]), .Z(n5783) );
  NANDN U6859 ( .A(n5760), .B(sreg[1185]), .Z(n5764) );
  NAND U6860 ( .A(n5762), .B(n5761), .Z(n5763) );
  NAND U6861 ( .A(n5764), .B(n5763), .Z(n5782) );
  XOR U6862 ( .A(n5783), .B(n5782), .Z(c[1186]) );
  NANDN U6863 ( .A(n5766), .B(n5765), .Z(n5770) );
  OR U6864 ( .A(n5768), .B(n5767), .Z(n5769) );
  AND U6865 ( .A(n5770), .B(n5769), .Z(n5788) );
  XOR U6866 ( .A(a[165]), .B(n2199), .Z(n5792) );
  AND U6867 ( .A(a[167]), .B(b[0]), .Z(n5772) );
  XNOR U6868 ( .A(n5772), .B(n2175), .Z(n5774) );
  NANDN U6869 ( .A(b[0]), .B(a[166]), .Z(n5773) );
  NAND U6870 ( .A(n5774), .B(n5773), .Z(n5797) );
  AND U6871 ( .A(a[163]), .B(b[3]), .Z(n5796) );
  XOR U6872 ( .A(n5797), .B(n5796), .Z(n5799) );
  XOR U6873 ( .A(n5798), .B(n5799), .Z(n5787) );
  NANDN U6874 ( .A(n5776), .B(n5775), .Z(n5780) );
  OR U6875 ( .A(n5778), .B(n5777), .Z(n5779) );
  AND U6876 ( .A(n5780), .B(n5779), .Z(n5786) );
  XOR U6877 ( .A(n5787), .B(n5786), .Z(n5789) );
  XOR U6878 ( .A(n5788), .B(n5789), .Z(n5802) );
  XNOR U6879 ( .A(n5802), .B(sreg[1187]), .Z(n5804) );
  NANDN U6880 ( .A(n5781), .B(sreg[1186]), .Z(n5785) );
  NAND U6881 ( .A(n5783), .B(n5782), .Z(n5784) );
  NAND U6882 ( .A(n5785), .B(n5784), .Z(n5803) );
  XOR U6883 ( .A(n5804), .B(n5803), .Z(c[1187]) );
  NANDN U6884 ( .A(n5787), .B(n5786), .Z(n5791) );
  OR U6885 ( .A(n5789), .B(n5788), .Z(n5790) );
  AND U6886 ( .A(n5791), .B(n5790), .Z(n5809) );
  XOR U6887 ( .A(a[166]), .B(n2199), .Z(n5813) );
  AND U6888 ( .A(a[168]), .B(b[0]), .Z(n5793) );
  XNOR U6889 ( .A(n5793), .B(n2175), .Z(n5795) );
  NANDN U6890 ( .A(b[0]), .B(a[167]), .Z(n5794) );
  NAND U6891 ( .A(n5795), .B(n5794), .Z(n5818) );
  AND U6892 ( .A(a[164]), .B(b[3]), .Z(n5817) );
  XOR U6893 ( .A(n5818), .B(n5817), .Z(n5820) );
  XOR U6894 ( .A(n5819), .B(n5820), .Z(n5808) );
  NANDN U6895 ( .A(n5797), .B(n5796), .Z(n5801) );
  OR U6896 ( .A(n5799), .B(n5798), .Z(n5800) );
  AND U6897 ( .A(n5801), .B(n5800), .Z(n5807) );
  XOR U6898 ( .A(n5808), .B(n5807), .Z(n5810) );
  XOR U6899 ( .A(n5809), .B(n5810), .Z(n5823) );
  XNOR U6900 ( .A(n5823), .B(sreg[1188]), .Z(n5825) );
  NANDN U6901 ( .A(n5802), .B(sreg[1187]), .Z(n5806) );
  NAND U6902 ( .A(n5804), .B(n5803), .Z(n5805) );
  NAND U6903 ( .A(n5806), .B(n5805), .Z(n5824) );
  XOR U6904 ( .A(n5825), .B(n5824), .Z(c[1188]) );
  NANDN U6905 ( .A(n5808), .B(n5807), .Z(n5812) );
  OR U6906 ( .A(n5810), .B(n5809), .Z(n5811) );
  AND U6907 ( .A(n5812), .B(n5811), .Z(n5830) );
  XOR U6908 ( .A(a[167]), .B(n2200), .Z(n5834) );
  AND U6909 ( .A(a[169]), .B(b[0]), .Z(n5814) );
  XNOR U6910 ( .A(n5814), .B(n2175), .Z(n5816) );
  NANDN U6911 ( .A(b[0]), .B(a[168]), .Z(n5815) );
  NAND U6912 ( .A(n5816), .B(n5815), .Z(n5839) );
  AND U6913 ( .A(a[165]), .B(b[3]), .Z(n5838) );
  XOR U6914 ( .A(n5839), .B(n5838), .Z(n5841) );
  XOR U6915 ( .A(n5840), .B(n5841), .Z(n5829) );
  NANDN U6916 ( .A(n5818), .B(n5817), .Z(n5822) );
  OR U6917 ( .A(n5820), .B(n5819), .Z(n5821) );
  AND U6918 ( .A(n5822), .B(n5821), .Z(n5828) );
  XOR U6919 ( .A(n5829), .B(n5828), .Z(n5831) );
  XOR U6920 ( .A(n5830), .B(n5831), .Z(n5844) );
  XNOR U6921 ( .A(n5844), .B(sreg[1189]), .Z(n5846) );
  NANDN U6922 ( .A(n5823), .B(sreg[1188]), .Z(n5827) );
  NAND U6923 ( .A(n5825), .B(n5824), .Z(n5826) );
  NAND U6924 ( .A(n5827), .B(n5826), .Z(n5845) );
  XOR U6925 ( .A(n5846), .B(n5845), .Z(c[1189]) );
  NANDN U6926 ( .A(n5829), .B(n5828), .Z(n5833) );
  OR U6927 ( .A(n5831), .B(n5830), .Z(n5832) );
  AND U6928 ( .A(n5833), .B(n5832), .Z(n5851) );
  XOR U6929 ( .A(a[168]), .B(n2200), .Z(n5855) );
  AND U6930 ( .A(a[170]), .B(b[0]), .Z(n5835) );
  XNOR U6931 ( .A(n5835), .B(n2175), .Z(n5837) );
  NANDN U6932 ( .A(b[0]), .B(a[169]), .Z(n5836) );
  NAND U6933 ( .A(n5837), .B(n5836), .Z(n5860) );
  AND U6934 ( .A(a[166]), .B(b[3]), .Z(n5859) );
  XOR U6935 ( .A(n5860), .B(n5859), .Z(n5862) );
  XOR U6936 ( .A(n5861), .B(n5862), .Z(n5850) );
  NANDN U6937 ( .A(n5839), .B(n5838), .Z(n5843) );
  OR U6938 ( .A(n5841), .B(n5840), .Z(n5842) );
  AND U6939 ( .A(n5843), .B(n5842), .Z(n5849) );
  XOR U6940 ( .A(n5850), .B(n5849), .Z(n5852) );
  XOR U6941 ( .A(n5851), .B(n5852), .Z(n5865) );
  XNOR U6942 ( .A(n5865), .B(sreg[1190]), .Z(n5867) );
  NANDN U6943 ( .A(n5844), .B(sreg[1189]), .Z(n5848) );
  NAND U6944 ( .A(n5846), .B(n5845), .Z(n5847) );
  NAND U6945 ( .A(n5848), .B(n5847), .Z(n5866) );
  XOR U6946 ( .A(n5867), .B(n5866), .Z(c[1190]) );
  NANDN U6947 ( .A(n5850), .B(n5849), .Z(n5854) );
  OR U6948 ( .A(n5852), .B(n5851), .Z(n5853) );
  AND U6949 ( .A(n5854), .B(n5853), .Z(n5872) );
  XOR U6950 ( .A(a[169]), .B(n2200), .Z(n5876) );
  AND U6951 ( .A(a[171]), .B(b[0]), .Z(n5856) );
  XNOR U6952 ( .A(n5856), .B(n2175), .Z(n5858) );
  NANDN U6953 ( .A(b[0]), .B(a[170]), .Z(n5857) );
  NAND U6954 ( .A(n5858), .B(n5857), .Z(n5881) );
  AND U6955 ( .A(a[167]), .B(b[3]), .Z(n5880) );
  XOR U6956 ( .A(n5881), .B(n5880), .Z(n5883) );
  XOR U6957 ( .A(n5882), .B(n5883), .Z(n5871) );
  NANDN U6958 ( .A(n5860), .B(n5859), .Z(n5864) );
  OR U6959 ( .A(n5862), .B(n5861), .Z(n5863) );
  AND U6960 ( .A(n5864), .B(n5863), .Z(n5870) );
  XOR U6961 ( .A(n5871), .B(n5870), .Z(n5873) );
  XOR U6962 ( .A(n5872), .B(n5873), .Z(n5886) );
  XNOR U6963 ( .A(n5886), .B(sreg[1191]), .Z(n5888) );
  NANDN U6964 ( .A(n5865), .B(sreg[1190]), .Z(n5869) );
  NAND U6965 ( .A(n5867), .B(n5866), .Z(n5868) );
  NAND U6966 ( .A(n5869), .B(n5868), .Z(n5887) );
  XOR U6967 ( .A(n5888), .B(n5887), .Z(c[1191]) );
  NANDN U6968 ( .A(n5871), .B(n5870), .Z(n5875) );
  OR U6969 ( .A(n5873), .B(n5872), .Z(n5874) );
  AND U6970 ( .A(n5875), .B(n5874), .Z(n5893) );
  XOR U6971 ( .A(a[170]), .B(n2200), .Z(n5897) );
  AND U6972 ( .A(a[172]), .B(b[0]), .Z(n5877) );
  XNOR U6973 ( .A(n5877), .B(n2175), .Z(n5879) );
  NANDN U6974 ( .A(b[0]), .B(a[171]), .Z(n5878) );
  NAND U6975 ( .A(n5879), .B(n5878), .Z(n5902) );
  AND U6976 ( .A(a[168]), .B(b[3]), .Z(n5901) );
  XOR U6977 ( .A(n5902), .B(n5901), .Z(n5904) );
  XOR U6978 ( .A(n5903), .B(n5904), .Z(n5892) );
  NANDN U6979 ( .A(n5881), .B(n5880), .Z(n5885) );
  OR U6980 ( .A(n5883), .B(n5882), .Z(n5884) );
  AND U6981 ( .A(n5885), .B(n5884), .Z(n5891) );
  XOR U6982 ( .A(n5892), .B(n5891), .Z(n5894) );
  XOR U6983 ( .A(n5893), .B(n5894), .Z(n5907) );
  XNOR U6984 ( .A(n5907), .B(sreg[1192]), .Z(n5909) );
  NANDN U6985 ( .A(n5886), .B(sreg[1191]), .Z(n5890) );
  NAND U6986 ( .A(n5888), .B(n5887), .Z(n5889) );
  NAND U6987 ( .A(n5890), .B(n5889), .Z(n5908) );
  XOR U6988 ( .A(n5909), .B(n5908), .Z(c[1192]) );
  NANDN U6989 ( .A(n5892), .B(n5891), .Z(n5896) );
  OR U6990 ( .A(n5894), .B(n5893), .Z(n5895) );
  AND U6991 ( .A(n5896), .B(n5895), .Z(n5914) );
  XOR U6992 ( .A(a[171]), .B(n2200), .Z(n5918) );
  AND U6993 ( .A(a[169]), .B(b[3]), .Z(n5922) );
  AND U6994 ( .A(a[173]), .B(b[0]), .Z(n5898) );
  XNOR U6995 ( .A(n5898), .B(n2175), .Z(n5900) );
  NANDN U6996 ( .A(b[0]), .B(a[172]), .Z(n5899) );
  NAND U6997 ( .A(n5900), .B(n5899), .Z(n5923) );
  XOR U6998 ( .A(n5922), .B(n5923), .Z(n5925) );
  XOR U6999 ( .A(n5924), .B(n5925), .Z(n5913) );
  NANDN U7000 ( .A(n5902), .B(n5901), .Z(n5906) );
  OR U7001 ( .A(n5904), .B(n5903), .Z(n5905) );
  AND U7002 ( .A(n5906), .B(n5905), .Z(n5912) );
  XOR U7003 ( .A(n5913), .B(n5912), .Z(n5915) );
  XOR U7004 ( .A(n5914), .B(n5915), .Z(n5928) );
  XNOR U7005 ( .A(n5928), .B(sreg[1193]), .Z(n5930) );
  NANDN U7006 ( .A(n5907), .B(sreg[1192]), .Z(n5911) );
  NAND U7007 ( .A(n5909), .B(n5908), .Z(n5910) );
  NAND U7008 ( .A(n5911), .B(n5910), .Z(n5929) );
  XOR U7009 ( .A(n5930), .B(n5929), .Z(c[1193]) );
  NANDN U7010 ( .A(n5913), .B(n5912), .Z(n5917) );
  OR U7011 ( .A(n5915), .B(n5914), .Z(n5916) );
  AND U7012 ( .A(n5917), .B(n5916), .Z(n5935) );
  XOR U7013 ( .A(a[172]), .B(n2200), .Z(n5939) );
  AND U7014 ( .A(a[174]), .B(b[0]), .Z(n5919) );
  XNOR U7015 ( .A(n5919), .B(n2175), .Z(n5921) );
  NANDN U7016 ( .A(b[0]), .B(a[173]), .Z(n5920) );
  NAND U7017 ( .A(n5921), .B(n5920), .Z(n5944) );
  AND U7018 ( .A(a[170]), .B(b[3]), .Z(n5943) );
  XOR U7019 ( .A(n5944), .B(n5943), .Z(n5946) );
  XOR U7020 ( .A(n5945), .B(n5946), .Z(n5934) );
  NANDN U7021 ( .A(n5923), .B(n5922), .Z(n5927) );
  OR U7022 ( .A(n5925), .B(n5924), .Z(n5926) );
  AND U7023 ( .A(n5927), .B(n5926), .Z(n5933) );
  XOR U7024 ( .A(n5934), .B(n5933), .Z(n5936) );
  XOR U7025 ( .A(n5935), .B(n5936), .Z(n5949) );
  XNOR U7026 ( .A(n5949), .B(sreg[1194]), .Z(n5951) );
  NANDN U7027 ( .A(n5928), .B(sreg[1193]), .Z(n5932) );
  NAND U7028 ( .A(n5930), .B(n5929), .Z(n5931) );
  NAND U7029 ( .A(n5932), .B(n5931), .Z(n5950) );
  XOR U7030 ( .A(n5951), .B(n5950), .Z(c[1194]) );
  NANDN U7031 ( .A(n5934), .B(n5933), .Z(n5938) );
  OR U7032 ( .A(n5936), .B(n5935), .Z(n5937) );
  AND U7033 ( .A(n5938), .B(n5937), .Z(n5956) );
  XOR U7034 ( .A(a[173]), .B(n2200), .Z(n5960) );
  AND U7035 ( .A(a[175]), .B(b[0]), .Z(n5940) );
  XNOR U7036 ( .A(n5940), .B(n2175), .Z(n5942) );
  NANDN U7037 ( .A(b[0]), .B(a[174]), .Z(n5941) );
  NAND U7038 ( .A(n5942), .B(n5941), .Z(n5965) );
  AND U7039 ( .A(a[171]), .B(b[3]), .Z(n5964) );
  XOR U7040 ( .A(n5965), .B(n5964), .Z(n5967) );
  XOR U7041 ( .A(n5966), .B(n5967), .Z(n5955) );
  NANDN U7042 ( .A(n5944), .B(n5943), .Z(n5948) );
  OR U7043 ( .A(n5946), .B(n5945), .Z(n5947) );
  AND U7044 ( .A(n5948), .B(n5947), .Z(n5954) );
  XOR U7045 ( .A(n5955), .B(n5954), .Z(n5957) );
  XOR U7046 ( .A(n5956), .B(n5957), .Z(n5970) );
  XNOR U7047 ( .A(n5970), .B(sreg[1195]), .Z(n5972) );
  NANDN U7048 ( .A(n5949), .B(sreg[1194]), .Z(n5953) );
  NAND U7049 ( .A(n5951), .B(n5950), .Z(n5952) );
  NAND U7050 ( .A(n5953), .B(n5952), .Z(n5971) );
  XOR U7051 ( .A(n5972), .B(n5971), .Z(c[1195]) );
  NANDN U7052 ( .A(n5955), .B(n5954), .Z(n5959) );
  OR U7053 ( .A(n5957), .B(n5956), .Z(n5958) );
  AND U7054 ( .A(n5959), .B(n5958), .Z(n5977) );
  XOR U7055 ( .A(a[174]), .B(n2201), .Z(n5981) );
  AND U7056 ( .A(a[172]), .B(b[3]), .Z(n5985) );
  AND U7057 ( .A(a[176]), .B(b[0]), .Z(n5961) );
  XNOR U7058 ( .A(n5961), .B(n2175), .Z(n5963) );
  NANDN U7059 ( .A(b[0]), .B(a[175]), .Z(n5962) );
  NAND U7060 ( .A(n5963), .B(n5962), .Z(n5986) );
  XOR U7061 ( .A(n5985), .B(n5986), .Z(n5988) );
  XOR U7062 ( .A(n5987), .B(n5988), .Z(n5976) );
  NANDN U7063 ( .A(n5965), .B(n5964), .Z(n5969) );
  OR U7064 ( .A(n5967), .B(n5966), .Z(n5968) );
  AND U7065 ( .A(n5969), .B(n5968), .Z(n5975) );
  XOR U7066 ( .A(n5976), .B(n5975), .Z(n5978) );
  XOR U7067 ( .A(n5977), .B(n5978), .Z(n5991) );
  XNOR U7068 ( .A(n5991), .B(sreg[1196]), .Z(n5993) );
  NANDN U7069 ( .A(n5970), .B(sreg[1195]), .Z(n5974) );
  NAND U7070 ( .A(n5972), .B(n5971), .Z(n5973) );
  NAND U7071 ( .A(n5974), .B(n5973), .Z(n5992) );
  XOR U7072 ( .A(n5993), .B(n5992), .Z(c[1196]) );
  NANDN U7073 ( .A(n5976), .B(n5975), .Z(n5980) );
  OR U7074 ( .A(n5978), .B(n5977), .Z(n5979) );
  AND U7075 ( .A(n5980), .B(n5979), .Z(n5998) );
  XOR U7076 ( .A(a[175]), .B(n2201), .Z(n6002) );
  AND U7077 ( .A(a[177]), .B(b[0]), .Z(n5982) );
  XNOR U7078 ( .A(n5982), .B(n2175), .Z(n5984) );
  NANDN U7079 ( .A(b[0]), .B(a[176]), .Z(n5983) );
  NAND U7080 ( .A(n5984), .B(n5983), .Z(n6007) );
  AND U7081 ( .A(a[173]), .B(b[3]), .Z(n6006) );
  XOR U7082 ( .A(n6007), .B(n6006), .Z(n6009) );
  XOR U7083 ( .A(n6008), .B(n6009), .Z(n5997) );
  NANDN U7084 ( .A(n5986), .B(n5985), .Z(n5990) );
  OR U7085 ( .A(n5988), .B(n5987), .Z(n5989) );
  AND U7086 ( .A(n5990), .B(n5989), .Z(n5996) );
  XOR U7087 ( .A(n5997), .B(n5996), .Z(n5999) );
  XOR U7088 ( .A(n5998), .B(n5999), .Z(n6012) );
  XNOR U7089 ( .A(n6012), .B(sreg[1197]), .Z(n6014) );
  NANDN U7090 ( .A(n5991), .B(sreg[1196]), .Z(n5995) );
  NAND U7091 ( .A(n5993), .B(n5992), .Z(n5994) );
  NAND U7092 ( .A(n5995), .B(n5994), .Z(n6013) );
  XOR U7093 ( .A(n6014), .B(n6013), .Z(c[1197]) );
  NANDN U7094 ( .A(n5997), .B(n5996), .Z(n6001) );
  OR U7095 ( .A(n5999), .B(n5998), .Z(n6000) );
  AND U7096 ( .A(n6001), .B(n6000), .Z(n6019) );
  XOR U7097 ( .A(a[176]), .B(n2201), .Z(n6023) );
  AND U7098 ( .A(a[174]), .B(b[3]), .Z(n6027) );
  AND U7099 ( .A(a[178]), .B(b[0]), .Z(n6003) );
  XNOR U7100 ( .A(n6003), .B(n2175), .Z(n6005) );
  NANDN U7101 ( .A(b[0]), .B(a[177]), .Z(n6004) );
  NAND U7102 ( .A(n6005), .B(n6004), .Z(n6028) );
  XOR U7103 ( .A(n6027), .B(n6028), .Z(n6030) );
  XOR U7104 ( .A(n6029), .B(n6030), .Z(n6018) );
  NANDN U7105 ( .A(n6007), .B(n6006), .Z(n6011) );
  OR U7106 ( .A(n6009), .B(n6008), .Z(n6010) );
  AND U7107 ( .A(n6011), .B(n6010), .Z(n6017) );
  XOR U7108 ( .A(n6018), .B(n6017), .Z(n6020) );
  XOR U7109 ( .A(n6019), .B(n6020), .Z(n6033) );
  XNOR U7110 ( .A(n6033), .B(sreg[1198]), .Z(n6035) );
  NANDN U7111 ( .A(n6012), .B(sreg[1197]), .Z(n6016) );
  NAND U7112 ( .A(n6014), .B(n6013), .Z(n6015) );
  NAND U7113 ( .A(n6016), .B(n6015), .Z(n6034) );
  XOR U7114 ( .A(n6035), .B(n6034), .Z(c[1198]) );
  NANDN U7115 ( .A(n6018), .B(n6017), .Z(n6022) );
  OR U7116 ( .A(n6020), .B(n6019), .Z(n6021) );
  AND U7117 ( .A(n6022), .B(n6021), .Z(n6040) );
  XOR U7118 ( .A(a[177]), .B(n2201), .Z(n6044) );
  AND U7119 ( .A(a[179]), .B(b[0]), .Z(n6024) );
  XNOR U7120 ( .A(n6024), .B(n2175), .Z(n6026) );
  NANDN U7121 ( .A(b[0]), .B(a[178]), .Z(n6025) );
  NAND U7122 ( .A(n6026), .B(n6025), .Z(n6049) );
  AND U7123 ( .A(a[175]), .B(b[3]), .Z(n6048) );
  XOR U7124 ( .A(n6049), .B(n6048), .Z(n6051) );
  XOR U7125 ( .A(n6050), .B(n6051), .Z(n6039) );
  NANDN U7126 ( .A(n6028), .B(n6027), .Z(n6032) );
  OR U7127 ( .A(n6030), .B(n6029), .Z(n6031) );
  AND U7128 ( .A(n6032), .B(n6031), .Z(n6038) );
  XOR U7129 ( .A(n6039), .B(n6038), .Z(n6041) );
  XOR U7130 ( .A(n6040), .B(n6041), .Z(n6054) );
  XNOR U7131 ( .A(n6054), .B(sreg[1199]), .Z(n6056) );
  NANDN U7132 ( .A(n6033), .B(sreg[1198]), .Z(n6037) );
  NAND U7133 ( .A(n6035), .B(n6034), .Z(n6036) );
  NAND U7134 ( .A(n6037), .B(n6036), .Z(n6055) );
  XOR U7135 ( .A(n6056), .B(n6055), .Z(c[1199]) );
  NANDN U7136 ( .A(n6039), .B(n6038), .Z(n6043) );
  OR U7137 ( .A(n6041), .B(n6040), .Z(n6042) );
  AND U7138 ( .A(n6043), .B(n6042), .Z(n6061) );
  XOR U7139 ( .A(a[178]), .B(n2201), .Z(n6065) );
  AND U7140 ( .A(a[176]), .B(b[3]), .Z(n6069) );
  AND U7141 ( .A(a[180]), .B(b[0]), .Z(n6045) );
  XNOR U7142 ( .A(n6045), .B(n2175), .Z(n6047) );
  NANDN U7143 ( .A(b[0]), .B(a[179]), .Z(n6046) );
  NAND U7144 ( .A(n6047), .B(n6046), .Z(n6070) );
  XOR U7145 ( .A(n6069), .B(n6070), .Z(n6072) );
  XOR U7146 ( .A(n6071), .B(n6072), .Z(n6060) );
  NANDN U7147 ( .A(n6049), .B(n6048), .Z(n6053) );
  OR U7148 ( .A(n6051), .B(n6050), .Z(n6052) );
  AND U7149 ( .A(n6053), .B(n6052), .Z(n6059) );
  XOR U7150 ( .A(n6060), .B(n6059), .Z(n6062) );
  XOR U7151 ( .A(n6061), .B(n6062), .Z(n6075) );
  XNOR U7152 ( .A(n6075), .B(sreg[1200]), .Z(n6077) );
  NANDN U7153 ( .A(n6054), .B(sreg[1199]), .Z(n6058) );
  NAND U7154 ( .A(n6056), .B(n6055), .Z(n6057) );
  NAND U7155 ( .A(n6058), .B(n6057), .Z(n6076) );
  XOR U7156 ( .A(n6077), .B(n6076), .Z(c[1200]) );
  NANDN U7157 ( .A(n6060), .B(n6059), .Z(n6064) );
  OR U7158 ( .A(n6062), .B(n6061), .Z(n6063) );
  AND U7159 ( .A(n6064), .B(n6063), .Z(n6082) );
  XOR U7160 ( .A(a[179]), .B(n2201), .Z(n6086) );
  AND U7161 ( .A(a[181]), .B(b[0]), .Z(n6066) );
  XNOR U7162 ( .A(n6066), .B(n2175), .Z(n6068) );
  NANDN U7163 ( .A(b[0]), .B(a[180]), .Z(n6067) );
  NAND U7164 ( .A(n6068), .B(n6067), .Z(n6091) );
  AND U7165 ( .A(a[177]), .B(b[3]), .Z(n6090) );
  XOR U7166 ( .A(n6091), .B(n6090), .Z(n6093) );
  XOR U7167 ( .A(n6092), .B(n6093), .Z(n6081) );
  NANDN U7168 ( .A(n6070), .B(n6069), .Z(n6074) );
  OR U7169 ( .A(n6072), .B(n6071), .Z(n6073) );
  AND U7170 ( .A(n6074), .B(n6073), .Z(n6080) );
  XOR U7171 ( .A(n6081), .B(n6080), .Z(n6083) );
  XOR U7172 ( .A(n6082), .B(n6083), .Z(n6096) );
  XNOR U7173 ( .A(n6096), .B(sreg[1201]), .Z(n6098) );
  NANDN U7174 ( .A(n6075), .B(sreg[1200]), .Z(n6079) );
  NAND U7175 ( .A(n6077), .B(n6076), .Z(n6078) );
  NAND U7176 ( .A(n6079), .B(n6078), .Z(n6097) );
  XOR U7177 ( .A(n6098), .B(n6097), .Z(c[1201]) );
  NANDN U7178 ( .A(n6081), .B(n6080), .Z(n6085) );
  OR U7179 ( .A(n6083), .B(n6082), .Z(n6084) );
  AND U7180 ( .A(n6085), .B(n6084), .Z(n6103) );
  XOR U7181 ( .A(a[180]), .B(n2201), .Z(n6107) );
  AND U7182 ( .A(a[182]), .B(b[0]), .Z(n6087) );
  XNOR U7183 ( .A(n6087), .B(n2175), .Z(n6089) );
  NANDN U7184 ( .A(b[0]), .B(a[181]), .Z(n6088) );
  NAND U7185 ( .A(n6089), .B(n6088), .Z(n6112) );
  AND U7186 ( .A(a[178]), .B(b[3]), .Z(n6111) );
  XOR U7187 ( .A(n6112), .B(n6111), .Z(n6114) );
  XOR U7188 ( .A(n6113), .B(n6114), .Z(n6102) );
  NANDN U7189 ( .A(n6091), .B(n6090), .Z(n6095) );
  OR U7190 ( .A(n6093), .B(n6092), .Z(n6094) );
  AND U7191 ( .A(n6095), .B(n6094), .Z(n6101) );
  XOR U7192 ( .A(n6102), .B(n6101), .Z(n6104) );
  XOR U7193 ( .A(n6103), .B(n6104), .Z(n6117) );
  XNOR U7194 ( .A(n6117), .B(sreg[1202]), .Z(n6119) );
  NANDN U7195 ( .A(n6096), .B(sreg[1201]), .Z(n6100) );
  NAND U7196 ( .A(n6098), .B(n6097), .Z(n6099) );
  NAND U7197 ( .A(n6100), .B(n6099), .Z(n6118) );
  XOR U7198 ( .A(n6119), .B(n6118), .Z(c[1202]) );
  NANDN U7199 ( .A(n6102), .B(n6101), .Z(n6106) );
  OR U7200 ( .A(n6104), .B(n6103), .Z(n6105) );
  AND U7201 ( .A(n6106), .B(n6105), .Z(n6124) );
  XOR U7202 ( .A(a[181]), .B(n2202), .Z(n6128) );
  AND U7203 ( .A(a[183]), .B(b[0]), .Z(n6108) );
  XNOR U7204 ( .A(n6108), .B(n2175), .Z(n6110) );
  NANDN U7205 ( .A(b[0]), .B(a[182]), .Z(n6109) );
  NAND U7206 ( .A(n6110), .B(n6109), .Z(n6133) );
  AND U7207 ( .A(a[179]), .B(b[3]), .Z(n6132) );
  XOR U7208 ( .A(n6133), .B(n6132), .Z(n6135) );
  XOR U7209 ( .A(n6134), .B(n6135), .Z(n6123) );
  NANDN U7210 ( .A(n6112), .B(n6111), .Z(n6116) );
  OR U7211 ( .A(n6114), .B(n6113), .Z(n6115) );
  AND U7212 ( .A(n6116), .B(n6115), .Z(n6122) );
  XOR U7213 ( .A(n6123), .B(n6122), .Z(n6125) );
  XOR U7214 ( .A(n6124), .B(n6125), .Z(n6138) );
  XNOR U7215 ( .A(n6138), .B(sreg[1203]), .Z(n6140) );
  NANDN U7216 ( .A(n6117), .B(sreg[1202]), .Z(n6121) );
  NAND U7217 ( .A(n6119), .B(n6118), .Z(n6120) );
  NAND U7218 ( .A(n6121), .B(n6120), .Z(n6139) );
  XOR U7219 ( .A(n6140), .B(n6139), .Z(c[1203]) );
  NANDN U7220 ( .A(n6123), .B(n6122), .Z(n6127) );
  OR U7221 ( .A(n6125), .B(n6124), .Z(n6126) );
  AND U7222 ( .A(n6127), .B(n6126), .Z(n6145) );
  XOR U7223 ( .A(a[182]), .B(n2202), .Z(n6149) );
  AND U7224 ( .A(a[180]), .B(b[3]), .Z(n6153) );
  AND U7225 ( .A(a[184]), .B(b[0]), .Z(n6129) );
  XNOR U7226 ( .A(n6129), .B(n2175), .Z(n6131) );
  NANDN U7227 ( .A(b[0]), .B(a[183]), .Z(n6130) );
  NAND U7228 ( .A(n6131), .B(n6130), .Z(n6154) );
  XOR U7229 ( .A(n6153), .B(n6154), .Z(n6156) );
  XOR U7230 ( .A(n6155), .B(n6156), .Z(n6144) );
  NANDN U7231 ( .A(n6133), .B(n6132), .Z(n6137) );
  OR U7232 ( .A(n6135), .B(n6134), .Z(n6136) );
  AND U7233 ( .A(n6137), .B(n6136), .Z(n6143) );
  XOR U7234 ( .A(n6144), .B(n6143), .Z(n6146) );
  XOR U7235 ( .A(n6145), .B(n6146), .Z(n6159) );
  XNOR U7236 ( .A(n6159), .B(sreg[1204]), .Z(n6161) );
  NANDN U7237 ( .A(n6138), .B(sreg[1203]), .Z(n6142) );
  NAND U7238 ( .A(n6140), .B(n6139), .Z(n6141) );
  NAND U7239 ( .A(n6142), .B(n6141), .Z(n6160) );
  XOR U7240 ( .A(n6161), .B(n6160), .Z(c[1204]) );
  NANDN U7241 ( .A(n6144), .B(n6143), .Z(n6148) );
  OR U7242 ( .A(n6146), .B(n6145), .Z(n6147) );
  AND U7243 ( .A(n6148), .B(n6147), .Z(n6166) );
  XOR U7244 ( .A(a[183]), .B(n2202), .Z(n6170) );
  AND U7245 ( .A(a[185]), .B(b[0]), .Z(n6150) );
  XNOR U7246 ( .A(n6150), .B(n2175), .Z(n6152) );
  NANDN U7247 ( .A(b[0]), .B(a[184]), .Z(n6151) );
  NAND U7248 ( .A(n6152), .B(n6151), .Z(n6175) );
  AND U7249 ( .A(a[181]), .B(b[3]), .Z(n6174) );
  XOR U7250 ( .A(n6175), .B(n6174), .Z(n6177) );
  XOR U7251 ( .A(n6176), .B(n6177), .Z(n6165) );
  NANDN U7252 ( .A(n6154), .B(n6153), .Z(n6158) );
  OR U7253 ( .A(n6156), .B(n6155), .Z(n6157) );
  AND U7254 ( .A(n6158), .B(n6157), .Z(n6164) );
  XOR U7255 ( .A(n6165), .B(n6164), .Z(n6167) );
  XOR U7256 ( .A(n6166), .B(n6167), .Z(n6180) );
  XNOR U7257 ( .A(n6180), .B(sreg[1205]), .Z(n6182) );
  NANDN U7258 ( .A(n6159), .B(sreg[1204]), .Z(n6163) );
  NAND U7259 ( .A(n6161), .B(n6160), .Z(n6162) );
  NAND U7260 ( .A(n6163), .B(n6162), .Z(n6181) );
  XOR U7261 ( .A(n6182), .B(n6181), .Z(c[1205]) );
  NANDN U7262 ( .A(n6165), .B(n6164), .Z(n6169) );
  OR U7263 ( .A(n6167), .B(n6166), .Z(n6168) );
  AND U7264 ( .A(n6169), .B(n6168), .Z(n6187) );
  XOR U7265 ( .A(a[184]), .B(n2202), .Z(n6191) );
  AND U7266 ( .A(a[186]), .B(b[0]), .Z(n6171) );
  XNOR U7267 ( .A(n6171), .B(n2175), .Z(n6173) );
  NANDN U7268 ( .A(b[0]), .B(a[185]), .Z(n6172) );
  NAND U7269 ( .A(n6173), .B(n6172), .Z(n6196) );
  AND U7270 ( .A(a[182]), .B(b[3]), .Z(n6195) );
  XOR U7271 ( .A(n6196), .B(n6195), .Z(n6198) );
  XOR U7272 ( .A(n6197), .B(n6198), .Z(n6186) );
  NANDN U7273 ( .A(n6175), .B(n6174), .Z(n6179) );
  OR U7274 ( .A(n6177), .B(n6176), .Z(n6178) );
  AND U7275 ( .A(n6179), .B(n6178), .Z(n6185) );
  XOR U7276 ( .A(n6186), .B(n6185), .Z(n6188) );
  XOR U7277 ( .A(n6187), .B(n6188), .Z(n6201) );
  XNOR U7278 ( .A(n6201), .B(sreg[1206]), .Z(n6203) );
  NANDN U7279 ( .A(n6180), .B(sreg[1205]), .Z(n6184) );
  NAND U7280 ( .A(n6182), .B(n6181), .Z(n6183) );
  NAND U7281 ( .A(n6184), .B(n6183), .Z(n6202) );
  XOR U7282 ( .A(n6203), .B(n6202), .Z(c[1206]) );
  NANDN U7283 ( .A(n6186), .B(n6185), .Z(n6190) );
  OR U7284 ( .A(n6188), .B(n6187), .Z(n6189) );
  AND U7285 ( .A(n6190), .B(n6189), .Z(n6208) );
  XOR U7286 ( .A(a[185]), .B(n2202), .Z(n6212) );
  AND U7287 ( .A(a[187]), .B(b[0]), .Z(n6192) );
  XNOR U7288 ( .A(n6192), .B(n2175), .Z(n6194) );
  NANDN U7289 ( .A(b[0]), .B(a[186]), .Z(n6193) );
  NAND U7290 ( .A(n6194), .B(n6193), .Z(n6217) );
  AND U7291 ( .A(a[183]), .B(b[3]), .Z(n6216) );
  XOR U7292 ( .A(n6217), .B(n6216), .Z(n6219) );
  XOR U7293 ( .A(n6218), .B(n6219), .Z(n6207) );
  NANDN U7294 ( .A(n6196), .B(n6195), .Z(n6200) );
  OR U7295 ( .A(n6198), .B(n6197), .Z(n6199) );
  AND U7296 ( .A(n6200), .B(n6199), .Z(n6206) );
  XOR U7297 ( .A(n6207), .B(n6206), .Z(n6209) );
  XOR U7298 ( .A(n6208), .B(n6209), .Z(n6222) );
  XNOR U7299 ( .A(n6222), .B(sreg[1207]), .Z(n6224) );
  NANDN U7300 ( .A(n6201), .B(sreg[1206]), .Z(n6205) );
  NAND U7301 ( .A(n6203), .B(n6202), .Z(n6204) );
  NAND U7302 ( .A(n6205), .B(n6204), .Z(n6223) );
  XOR U7303 ( .A(n6224), .B(n6223), .Z(c[1207]) );
  NANDN U7304 ( .A(n6207), .B(n6206), .Z(n6211) );
  OR U7305 ( .A(n6209), .B(n6208), .Z(n6210) );
  AND U7306 ( .A(n6211), .B(n6210), .Z(n6229) );
  XOR U7307 ( .A(a[186]), .B(n2202), .Z(n6233) );
  AND U7308 ( .A(a[188]), .B(b[0]), .Z(n6213) );
  XNOR U7309 ( .A(n6213), .B(n2175), .Z(n6215) );
  NANDN U7310 ( .A(b[0]), .B(a[187]), .Z(n6214) );
  NAND U7311 ( .A(n6215), .B(n6214), .Z(n6238) );
  AND U7312 ( .A(a[184]), .B(b[3]), .Z(n6237) );
  XOR U7313 ( .A(n6238), .B(n6237), .Z(n6240) );
  XOR U7314 ( .A(n6239), .B(n6240), .Z(n6228) );
  NANDN U7315 ( .A(n6217), .B(n6216), .Z(n6221) );
  OR U7316 ( .A(n6219), .B(n6218), .Z(n6220) );
  AND U7317 ( .A(n6221), .B(n6220), .Z(n6227) );
  XOR U7318 ( .A(n6228), .B(n6227), .Z(n6230) );
  XOR U7319 ( .A(n6229), .B(n6230), .Z(n6243) );
  XNOR U7320 ( .A(n6243), .B(sreg[1208]), .Z(n6245) );
  NANDN U7321 ( .A(n6222), .B(sreg[1207]), .Z(n6226) );
  NAND U7322 ( .A(n6224), .B(n6223), .Z(n6225) );
  NAND U7323 ( .A(n6226), .B(n6225), .Z(n6244) );
  XOR U7324 ( .A(n6245), .B(n6244), .Z(c[1208]) );
  NANDN U7325 ( .A(n6228), .B(n6227), .Z(n6232) );
  OR U7326 ( .A(n6230), .B(n6229), .Z(n6231) );
  AND U7327 ( .A(n6232), .B(n6231), .Z(n6250) );
  XOR U7328 ( .A(a[187]), .B(n2202), .Z(n6254) );
  AND U7329 ( .A(a[189]), .B(b[0]), .Z(n6234) );
  XNOR U7330 ( .A(n6234), .B(n2175), .Z(n6236) );
  NANDN U7331 ( .A(b[0]), .B(a[188]), .Z(n6235) );
  NAND U7332 ( .A(n6236), .B(n6235), .Z(n6259) );
  AND U7333 ( .A(a[185]), .B(b[3]), .Z(n6258) );
  XOR U7334 ( .A(n6259), .B(n6258), .Z(n6261) );
  XOR U7335 ( .A(n6260), .B(n6261), .Z(n6249) );
  NANDN U7336 ( .A(n6238), .B(n6237), .Z(n6242) );
  OR U7337 ( .A(n6240), .B(n6239), .Z(n6241) );
  AND U7338 ( .A(n6242), .B(n6241), .Z(n6248) );
  XOR U7339 ( .A(n6249), .B(n6248), .Z(n6251) );
  XOR U7340 ( .A(n6250), .B(n6251), .Z(n6264) );
  XNOR U7341 ( .A(n6264), .B(sreg[1209]), .Z(n6266) );
  NANDN U7342 ( .A(n6243), .B(sreg[1208]), .Z(n6247) );
  NAND U7343 ( .A(n6245), .B(n6244), .Z(n6246) );
  NAND U7344 ( .A(n6247), .B(n6246), .Z(n6265) );
  XOR U7345 ( .A(n6266), .B(n6265), .Z(c[1209]) );
  NANDN U7346 ( .A(n6249), .B(n6248), .Z(n6253) );
  OR U7347 ( .A(n6251), .B(n6250), .Z(n6252) );
  AND U7348 ( .A(n6253), .B(n6252), .Z(n6271) );
  XOR U7349 ( .A(a[188]), .B(n2203), .Z(n6275) );
  AND U7350 ( .A(a[186]), .B(b[3]), .Z(n6279) );
  AND U7351 ( .A(a[190]), .B(b[0]), .Z(n6255) );
  XNOR U7352 ( .A(n6255), .B(n2175), .Z(n6257) );
  NANDN U7353 ( .A(b[0]), .B(a[189]), .Z(n6256) );
  NAND U7354 ( .A(n6257), .B(n6256), .Z(n6280) );
  XOR U7355 ( .A(n6279), .B(n6280), .Z(n6282) );
  XOR U7356 ( .A(n6281), .B(n6282), .Z(n6270) );
  NANDN U7357 ( .A(n6259), .B(n6258), .Z(n6263) );
  OR U7358 ( .A(n6261), .B(n6260), .Z(n6262) );
  AND U7359 ( .A(n6263), .B(n6262), .Z(n6269) );
  XOR U7360 ( .A(n6270), .B(n6269), .Z(n6272) );
  XOR U7361 ( .A(n6271), .B(n6272), .Z(n6285) );
  XNOR U7362 ( .A(n6285), .B(sreg[1210]), .Z(n6287) );
  NANDN U7363 ( .A(n6264), .B(sreg[1209]), .Z(n6268) );
  NAND U7364 ( .A(n6266), .B(n6265), .Z(n6267) );
  NAND U7365 ( .A(n6268), .B(n6267), .Z(n6286) );
  XOR U7366 ( .A(n6287), .B(n6286), .Z(c[1210]) );
  NANDN U7367 ( .A(n6270), .B(n6269), .Z(n6274) );
  OR U7368 ( .A(n6272), .B(n6271), .Z(n6273) );
  AND U7369 ( .A(n6274), .B(n6273), .Z(n6292) );
  XOR U7370 ( .A(a[189]), .B(n2203), .Z(n6296) );
  AND U7371 ( .A(a[187]), .B(b[3]), .Z(n6300) );
  AND U7372 ( .A(a[191]), .B(b[0]), .Z(n6276) );
  XNOR U7373 ( .A(n6276), .B(n2175), .Z(n6278) );
  NANDN U7374 ( .A(b[0]), .B(a[190]), .Z(n6277) );
  NAND U7375 ( .A(n6278), .B(n6277), .Z(n6301) );
  XOR U7376 ( .A(n6300), .B(n6301), .Z(n6303) );
  XOR U7377 ( .A(n6302), .B(n6303), .Z(n6291) );
  NANDN U7378 ( .A(n6280), .B(n6279), .Z(n6284) );
  OR U7379 ( .A(n6282), .B(n6281), .Z(n6283) );
  AND U7380 ( .A(n6284), .B(n6283), .Z(n6290) );
  XOR U7381 ( .A(n6291), .B(n6290), .Z(n6293) );
  XOR U7382 ( .A(n6292), .B(n6293), .Z(n6306) );
  XNOR U7383 ( .A(n6306), .B(sreg[1211]), .Z(n6308) );
  NANDN U7384 ( .A(n6285), .B(sreg[1210]), .Z(n6289) );
  NAND U7385 ( .A(n6287), .B(n6286), .Z(n6288) );
  NAND U7386 ( .A(n6289), .B(n6288), .Z(n6307) );
  XOR U7387 ( .A(n6308), .B(n6307), .Z(c[1211]) );
  NANDN U7388 ( .A(n6291), .B(n6290), .Z(n6295) );
  OR U7389 ( .A(n6293), .B(n6292), .Z(n6294) );
  AND U7390 ( .A(n6295), .B(n6294), .Z(n6313) );
  XOR U7391 ( .A(a[190]), .B(n2203), .Z(n6317) );
  AND U7392 ( .A(a[192]), .B(b[0]), .Z(n6297) );
  XNOR U7393 ( .A(n6297), .B(n2175), .Z(n6299) );
  NANDN U7394 ( .A(b[0]), .B(a[191]), .Z(n6298) );
  NAND U7395 ( .A(n6299), .B(n6298), .Z(n6322) );
  AND U7396 ( .A(a[188]), .B(b[3]), .Z(n6321) );
  XOR U7397 ( .A(n6322), .B(n6321), .Z(n6324) );
  XOR U7398 ( .A(n6323), .B(n6324), .Z(n6312) );
  NANDN U7399 ( .A(n6301), .B(n6300), .Z(n6305) );
  OR U7400 ( .A(n6303), .B(n6302), .Z(n6304) );
  AND U7401 ( .A(n6305), .B(n6304), .Z(n6311) );
  XOR U7402 ( .A(n6312), .B(n6311), .Z(n6314) );
  XOR U7403 ( .A(n6313), .B(n6314), .Z(n6327) );
  XNOR U7404 ( .A(n6327), .B(sreg[1212]), .Z(n6329) );
  NANDN U7405 ( .A(n6306), .B(sreg[1211]), .Z(n6310) );
  NAND U7406 ( .A(n6308), .B(n6307), .Z(n6309) );
  NAND U7407 ( .A(n6310), .B(n6309), .Z(n6328) );
  XOR U7408 ( .A(n6329), .B(n6328), .Z(c[1212]) );
  NANDN U7409 ( .A(n6312), .B(n6311), .Z(n6316) );
  OR U7410 ( .A(n6314), .B(n6313), .Z(n6315) );
  AND U7411 ( .A(n6316), .B(n6315), .Z(n6334) );
  XOR U7412 ( .A(a[191]), .B(n2203), .Z(n6338) );
  AND U7413 ( .A(a[189]), .B(b[3]), .Z(n6342) );
  AND U7414 ( .A(a[193]), .B(b[0]), .Z(n6318) );
  XNOR U7415 ( .A(n6318), .B(n2175), .Z(n6320) );
  NANDN U7416 ( .A(b[0]), .B(a[192]), .Z(n6319) );
  NAND U7417 ( .A(n6320), .B(n6319), .Z(n6343) );
  XOR U7418 ( .A(n6342), .B(n6343), .Z(n6345) );
  XOR U7419 ( .A(n6344), .B(n6345), .Z(n6333) );
  NANDN U7420 ( .A(n6322), .B(n6321), .Z(n6326) );
  OR U7421 ( .A(n6324), .B(n6323), .Z(n6325) );
  AND U7422 ( .A(n6326), .B(n6325), .Z(n6332) );
  XOR U7423 ( .A(n6333), .B(n6332), .Z(n6335) );
  XOR U7424 ( .A(n6334), .B(n6335), .Z(n6348) );
  XNOR U7425 ( .A(n6348), .B(sreg[1213]), .Z(n6350) );
  NANDN U7426 ( .A(n6327), .B(sreg[1212]), .Z(n6331) );
  NAND U7427 ( .A(n6329), .B(n6328), .Z(n6330) );
  NAND U7428 ( .A(n6331), .B(n6330), .Z(n6349) );
  XOR U7429 ( .A(n6350), .B(n6349), .Z(c[1213]) );
  NANDN U7430 ( .A(n6333), .B(n6332), .Z(n6337) );
  OR U7431 ( .A(n6335), .B(n6334), .Z(n6336) );
  AND U7432 ( .A(n6337), .B(n6336), .Z(n6355) );
  XOR U7433 ( .A(a[192]), .B(n2203), .Z(n6359) );
  AND U7434 ( .A(a[194]), .B(b[0]), .Z(n6339) );
  XNOR U7435 ( .A(n6339), .B(n2175), .Z(n6341) );
  NANDN U7436 ( .A(b[0]), .B(a[193]), .Z(n6340) );
  NAND U7437 ( .A(n6341), .B(n6340), .Z(n6364) );
  AND U7438 ( .A(a[190]), .B(b[3]), .Z(n6363) );
  XOR U7439 ( .A(n6364), .B(n6363), .Z(n6366) );
  XOR U7440 ( .A(n6365), .B(n6366), .Z(n6354) );
  NANDN U7441 ( .A(n6343), .B(n6342), .Z(n6347) );
  OR U7442 ( .A(n6345), .B(n6344), .Z(n6346) );
  AND U7443 ( .A(n6347), .B(n6346), .Z(n6353) );
  XOR U7444 ( .A(n6354), .B(n6353), .Z(n6356) );
  XOR U7445 ( .A(n6355), .B(n6356), .Z(n6369) );
  XNOR U7446 ( .A(n6369), .B(sreg[1214]), .Z(n6371) );
  NANDN U7447 ( .A(n6348), .B(sreg[1213]), .Z(n6352) );
  NAND U7448 ( .A(n6350), .B(n6349), .Z(n6351) );
  NAND U7449 ( .A(n6352), .B(n6351), .Z(n6370) );
  XOR U7450 ( .A(n6371), .B(n6370), .Z(c[1214]) );
  NANDN U7451 ( .A(n6354), .B(n6353), .Z(n6358) );
  OR U7452 ( .A(n6356), .B(n6355), .Z(n6357) );
  AND U7453 ( .A(n6358), .B(n6357), .Z(n6376) );
  XOR U7454 ( .A(a[193]), .B(n2203), .Z(n6380) );
  AND U7455 ( .A(a[191]), .B(b[3]), .Z(n6384) );
  AND U7456 ( .A(a[195]), .B(b[0]), .Z(n6360) );
  XNOR U7457 ( .A(n6360), .B(n2175), .Z(n6362) );
  NANDN U7458 ( .A(b[0]), .B(a[194]), .Z(n6361) );
  NAND U7459 ( .A(n6362), .B(n6361), .Z(n6385) );
  XOR U7460 ( .A(n6384), .B(n6385), .Z(n6387) );
  XOR U7461 ( .A(n6386), .B(n6387), .Z(n6375) );
  NANDN U7462 ( .A(n6364), .B(n6363), .Z(n6368) );
  OR U7463 ( .A(n6366), .B(n6365), .Z(n6367) );
  AND U7464 ( .A(n6368), .B(n6367), .Z(n6374) );
  XOR U7465 ( .A(n6375), .B(n6374), .Z(n6377) );
  XOR U7466 ( .A(n6376), .B(n6377), .Z(n6390) );
  XNOR U7467 ( .A(n6390), .B(sreg[1215]), .Z(n6392) );
  NANDN U7468 ( .A(n6369), .B(sreg[1214]), .Z(n6373) );
  NAND U7469 ( .A(n6371), .B(n6370), .Z(n6372) );
  NAND U7470 ( .A(n6373), .B(n6372), .Z(n6391) );
  XOR U7471 ( .A(n6392), .B(n6391), .Z(c[1215]) );
  NANDN U7472 ( .A(n6375), .B(n6374), .Z(n6379) );
  OR U7473 ( .A(n6377), .B(n6376), .Z(n6378) );
  AND U7474 ( .A(n6379), .B(n6378), .Z(n6397) );
  XOR U7475 ( .A(a[194]), .B(n2203), .Z(n6401) );
  AND U7476 ( .A(a[192]), .B(b[3]), .Z(n6405) );
  AND U7477 ( .A(a[196]), .B(b[0]), .Z(n6381) );
  XNOR U7478 ( .A(n6381), .B(n2175), .Z(n6383) );
  NANDN U7479 ( .A(b[0]), .B(a[195]), .Z(n6382) );
  NAND U7480 ( .A(n6383), .B(n6382), .Z(n6406) );
  XOR U7481 ( .A(n6405), .B(n6406), .Z(n6408) );
  XOR U7482 ( .A(n6407), .B(n6408), .Z(n6396) );
  NANDN U7483 ( .A(n6385), .B(n6384), .Z(n6389) );
  OR U7484 ( .A(n6387), .B(n6386), .Z(n6388) );
  AND U7485 ( .A(n6389), .B(n6388), .Z(n6395) );
  XOR U7486 ( .A(n6396), .B(n6395), .Z(n6398) );
  XOR U7487 ( .A(n6397), .B(n6398), .Z(n6411) );
  XNOR U7488 ( .A(n6411), .B(sreg[1216]), .Z(n6413) );
  NANDN U7489 ( .A(n6390), .B(sreg[1215]), .Z(n6394) );
  NAND U7490 ( .A(n6392), .B(n6391), .Z(n6393) );
  NAND U7491 ( .A(n6394), .B(n6393), .Z(n6412) );
  XOR U7492 ( .A(n6413), .B(n6412), .Z(c[1216]) );
  NANDN U7493 ( .A(n6396), .B(n6395), .Z(n6400) );
  OR U7494 ( .A(n6398), .B(n6397), .Z(n6399) );
  AND U7495 ( .A(n6400), .B(n6399), .Z(n6419) );
  XOR U7496 ( .A(a[195]), .B(n2204), .Z(n6420) );
  AND U7497 ( .A(b[0]), .B(a[197]), .Z(n6402) );
  XOR U7498 ( .A(b[1]), .B(n6402), .Z(n6404) );
  NANDN U7499 ( .A(b[0]), .B(a[196]), .Z(n6403) );
  AND U7500 ( .A(n6404), .B(n6403), .Z(n6424) );
  AND U7501 ( .A(a[193]), .B(b[3]), .Z(n6425) );
  XOR U7502 ( .A(n6424), .B(n6425), .Z(n6426) );
  XNOR U7503 ( .A(n6427), .B(n6426), .Z(n6416) );
  NANDN U7504 ( .A(n6406), .B(n6405), .Z(n6410) );
  OR U7505 ( .A(n6408), .B(n6407), .Z(n6409) );
  AND U7506 ( .A(n6410), .B(n6409), .Z(n6417) );
  XNOR U7507 ( .A(n6416), .B(n6417), .Z(n6418) );
  XNOR U7508 ( .A(n6419), .B(n6418), .Z(n6430) );
  XNOR U7509 ( .A(n6430), .B(sreg[1217]), .Z(n6432) );
  NANDN U7510 ( .A(n6411), .B(sreg[1216]), .Z(n6415) );
  NAND U7511 ( .A(n6413), .B(n6412), .Z(n6414) );
  NAND U7512 ( .A(n6415), .B(n6414), .Z(n6431) );
  XOR U7513 ( .A(n6432), .B(n6431), .Z(c[1217]) );
  XOR U7514 ( .A(a[196]), .B(n2204), .Z(n6439) );
  AND U7515 ( .A(a[198]), .B(b[0]), .Z(n6421) );
  XNOR U7516 ( .A(n6421), .B(n2175), .Z(n6423) );
  NANDN U7517 ( .A(b[0]), .B(a[197]), .Z(n6422) );
  NAND U7518 ( .A(n6423), .B(n6422), .Z(n6444) );
  AND U7519 ( .A(a[194]), .B(b[3]), .Z(n6443) );
  XOR U7520 ( .A(n6444), .B(n6443), .Z(n6446) );
  XOR U7521 ( .A(n6445), .B(n6446), .Z(n6434) );
  NAND U7522 ( .A(n6425), .B(n6424), .Z(n6429) );
  NANDN U7523 ( .A(n6427), .B(n6426), .Z(n6428) );
  AND U7524 ( .A(n6429), .B(n6428), .Z(n6433) );
  XOR U7525 ( .A(n6434), .B(n6433), .Z(n6436) );
  XOR U7526 ( .A(n6435), .B(n6436), .Z(n6449) );
  XNOR U7527 ( .A(n6449), .B(sreg[1218]), .Z(n6451) );
  XOR U7528 ( .A(n6451), .B(n6450), .Z(c[1218]) );
  NANDN U7529 ( .A(n6434), .B(n6433), .Z(n6438) );
  OR U7530 ( .A(n6436), .B(n6435), .Z(n6437) );
  AND U7531 ( .A(n6438), .B(n6437), .Z(n6456) );
  XOR U7532 ( .A(a[197]), .B(n2204), .Z(n6460) );
  AND U7533 ( .A(a[199]), .B(b[0]), .Z(n6440) );
  XNOR U7534 ( .A(n6440), .B(n2175), .Z(n6442) );
  NANDN U7535 ( .A(b[0]), .B(a[198]), .Z(n6441) );
  NAND U7536 ( .A(n6442), .B(n6441), .Z(n6465) );
  AND U7537 ( .A(a[195]), .B(b[3]), .Z(n6464) );
  XOR U7538 ( .A(n6465), .B(n6464), .Z(n6467) );
  XOR U7539 ( .A(n6466), .B(n6467), .Z(n6455) );
  NANDN U7540 ( .A(n6444), .B(n6443), .Z(n6448) );
  OR U7541 ( .A(n6446), .B(n6445), .Z(n6447) );
  AND U7542 ( .A(n6448), .B(n6447), .Z(n6454) );
  XOR U7543 ( .A(n6455), .B(n6454), .Z(n6457) );
  XOR U7544 ( .A(n6456), .B(n6457), .Z(n6470) );
  XNOR U7545 ( .A(n6470), .B(sreg[1219]), .Z(n6472) );
  NANDN U7546 ( .A(n6449), .B(sreg[1218]), .Z(n6453) );
  NAND U7547 ( .A(n6451), .B(n6450), .Z(n6452) );
  NAND U7548 ( .A(n6453), .B(n6452), .Z(n6471) );
  XOR U7549 ( .A(n6472), .B(n6471), .Z(c[1219]) );
  NANDN U7550 ( .A(n6455), .B(n6454), .Z(n6459) );
  OR U7551 ( .A(n6457), .B(n6456), .Z(n6458) );
  AND U7552 ( .A(n6459), .B(n6458), .Z(n6477) );
  XOR U7553 ( .A(a[198]), .B(n2204), .Z(n6481) );
  AND U7554 ( .A(a[200]), .B(b[0]), .Z(n6461) );
  XNOR U7555 ( .A(n6461), .B(n2175), .Z(n6463) );
  NANDN U7556 ( .A(b[0]), .B(a[199]), .Z(n6462) );
  NAND U7557 ( .A(n6463), .B(n6462), .Z(n6486) );
  AND U7558 ( .A(a[196]), .B(b[3]), .Z(n6485) );
  XOR U7559 ( .A(n6486), .B(n6485), .Z(n6488) );
  XOR U7560 ( .A(n6487), .B(n6488), .Z(n6476) );
  NANDN U7561 ( .A(n6465), .B(n6464), .Z(n6469) );
  OR U7562 ( .A(n6467), .B(n6466), .Z(n6468) );
  AND U7563 ( .A(n6469), .B(n6468), .Z(n6475) );
  XOR U7564 ( .A(n6476), .B(n6475), .Z(n6478) );
  XOR U7565 ( .A(n6477), .B(n6478), .Z(n6491) );
  XNOR U7566 ( .A(n6491), .B(sreg[1220]), .Z(n6493) );
  NANDN U7567 ( .A(n6470), .B(sreg[1219]), .Z(n6474) );
  NAND U7568 ( .A(n6472), .B(n6471), .Z(n6473) );
  NAND U7569 ( .A(n6474), .B(n6473), .Z(n6492) );
  XOR U7570 ( .A(n6493), .B(n6492), .Z(c[1220]) );
  NANDN U7571 ( .A(n6476), .B(n6475), .Z(n6480) );
  OR U7572 ( .A(n6478), .B(n6477), .Z(n6479) );
  AND U7573 ( .A(n6480), .B(n6479), .Z(n6498) );
  XOR U7574 ( .A(a[199]), .B(n2204), .Z(n6502) );
  AND U7575 ( .A(a[201]), .B(b[0]), .Z(n6482) );
  XNOR U7576 ( .A(n6482), .B(n2175), .Z(n6484) );
  NANDN U7577 ( .A(b[0]), .B(a[200]), .Z(n6483) );
  NAND U7578 ( .A(n6484), .B(n6483), .Z(n6507) );
  AND U7579 ( .A(a[197]), .B(b[3]), .Z(n6506) );
  XOR U7580 ( .A(n6507), .B(n6506), .Z(n6509) );
  XOR U7581 ( .A(n6508), .B(n6509), .Z(n6497) );
  NANDN U7582 ( .A(n6486), .B(n6485), .Z(n6490) );
  OR U7583 ( .A(n6488), .B(n6487), .Z(n6489) );
  AND U7584 ( .A(n6490), .B(n6489), .Z(n6496) );
  XOR U7585 ( .A(n6497), .B(n6496), .Z(n6499) );
  XOR U7586 ( .A(n6498), .B(n6499), .Z(n6512) );
  XNOR U7587 ( .A(n6512), .B(sreg[1221]), .Z(n6514) );
  NANDN U7588 ( .A(n6491), .B(sreg[1220]), .Z(n6495) );
  NAND U7589 ( .A(n6493), .B(n6492), .Z(n6494) );
  NAND U7590 ( .A(n6495), .B(n6494), .Z(n6513) );
  XOR U7591 ( .A(n6514), .B(n6513), .Z(c[1221]) );
  NANDN U7592 ( .A(n6497), .B(n6496), .Z(n6501) );
  OR U7593 ( .A(n6499), .B(n6498), .Z(n6500) );
  AND U7594 ( .A(n6501), .B(n6500), .Z(n6519) );
  XOR U7595 ( .A(a[200]), .B(n2204), .Z(n6523) );
  AND U7596 ( .A(a[202]), .B(b[0]), .Z(n6503) );
  XNOR U7597 ( .A(n6503), .B(n2175), .Z(n6505) );
  NANDN U7598 ( .A(b[0]), .B(a[201]), .Z(n6504) );
  NAND U7599 ( .A(n6505), .B(n6504), .Z(n6528) );
  AND U7600 ( .A(a[198]), .B(b[3]), .Z(n6527) );
  XOR U7601 ( .A(n6528), .B(n6527), .Z(n6530) );
  XOR U7602 ( .A(n6529), .B(n6530), .Z(n6518) );
  NANDN U7603 ( .A(n6507), .B(n6506), .Z(n6511) );
  OR U7604 ( .A(n6509), .B(n6508), .Z(n6510) );
  AND U7605 ( .A(n6511), .B(n6510), .Z(n6517) );
  XOR U7606 ( .A(n6518), .B(n6517), .Z(n6520) );
  XOR U7607 ( .A(n6519), .B(n6520), .Z(n6533) );
  XNOR U7608 ( .A(n6533), .B(sreg[1222]), .Z(n6535) );
  NANDN U7609 ( .A(n6512), .B(sreg[1221]), .Z(n6516) );
  NAND U7610 ( .A(n6514), .B(n6513), .Z(n6515) );
  NAND U7611 ( .A(n6516), .B(n6515), .Z(n6534) );
  XOR U7612 ( .A(n6535), .B(n6534), .Z(c[1222]) );
  NANDN U7613 ( .A(n6518), .B(n6517), .Z(n6522) );
  OR U7614 ( .A(n6520), .B(n6519), .Z(n6521) );
  AND U7615 ( .A(n6522), .B(n6521), .Z(n6540) );
  XOR U7616 ( .A(a[201]), .B(n2204), .Z(n6544) );
  AND U7617 ( .A(a[199]), .B(b[3]), .Z(n6548) );
  AND U7618 ( .A(a[203]), .B(b[0]), .Z(n6524) );
  XNOR U7619 ( .A(n6524), .B(n2175), .Z(n6526) );
  NANDN U7620 ( .A(b[0]), .B(a[202]), .Z(n6525) );
  NAND U7621 ( .A(n6526), .B(n6525), .Z(n6549) );
  XOR U7622 ( .A(n6548), .B(n6549), .Z(n6551) );
  XOR U7623 ( .A(n6550), .B(n6551), .Z(n6539) );
  NANDN U7624 ( .A(n6528), .B(n6527), .Z(n6532) );
  OR U7625 ( .A(n6530), .B(n6529), .Z(n6531) );
  AND U7626 ( .A(n6532), .B(n6531), .Z(n6538) );
  XOR U7627 ( .A(n6539), .B(n6538), .Z(n6541) );
  XOR U7628 ( .A(n6540), .B(n6541), .Z(n6554) );
  XNOR U7629 ( .A(n6554), .B(sreg[1223]), .Z(n6556) );
  NANDN U7630 ( .A(n6533), .B(sreg[1222]), .Z(n6537) );
  NAND U7631 ( .A(n6535), .B(n6534), .Z(n6536) );
  NAND U7632 ( .A(n6537), .B(n6536), .Z(n6555) );
  XOR U7633 ( .A(n6556), .B(n6555), .Z(c[1223]) );
  NANDN U7634 ( .A(n6539), .B(n6538), .Z(n6543) );
  OR U7635 ( .A(n6541), .B(n6540), .Z(n6542) );
  AND U7636 ( .A(n6543), .B(n6542), .Z(n6561) );
  XOR U7637 ( .A(a[202]), .B(n2205), .Z(n6565) );
  AND U7638 ( .A(a[204]), .B(b[0]), .Z(n6545) );
  XNOR U7639 ( .A(n6545), .B(n2175), .Z(n6547) );
  NANDN U7640 ( .A(b[0]), .B(a[203]), .Z(n6546) );
  NAND U7641 ( .A(n6547), .B(n6546), .Z(n6570) );
  AND U7642 ( .A(a[200]), .B(b[3]), .Z(n6569) );
  XOR U7643 ( .A(n6570), .B(n6569), .Z(n6572) );
  XOR U7644 ( .A(n6571), .B(n6572), .Z(n6560) );
  NANDN U7645 ( .A(n6549), .B(n6548), .Z(n6553) );
  OR U7646 ( .A(n6551), .B(n6550), .Z(n6552) );
  AND U7647 ( .A(n6553), .B(n6552), .Z(n6559) );
  XOR U7648 ( .A(n6560), .B(n6559), .Z(n6562) );
  XOR U7649 ( .A(n6561), .B(n6562), .Z(n6575) );
  XNOR U7650 ( .A(n6575), .B(sreg[1224]), .Z(n6577) );
  NANDN U7651 ( .A(n6554), .B(sreg[1223]), .Z(n6558) );
  NAND U7652 ( .A(n6556), .B(n6555), .Z(n6557) );
  NAND U7653 ( .A(n6558), .B(n6557), .Z(n6576) );
  XOR U7654 ( .A(n6577), .B(n6576), .Z(c[1224]) );
  NANDN U7655 ( .A(n6560), .B(n6559), .Z(n6564) );
  OR U7656 ( .A(n6562), .B(n6561), .Z(n6563) );
  AND U7657 ( .A(n6564), .B(n6563), .Z(n6582) );
  XOR U7658 ( .A(a[203]), .B(n2205), .Z(n6586) );
  AND U7659 ( .A(a[205]), .B(b[0]), .Z(n6566) );
  XNOR U7660 ( .A(n6566), .B(n2175), .Z(n6568) );
  NANDN U7661 ( .A(b[0]), .B(a[204]), .Z(n6567) );
  NAND U7662 ( .A(n6568), .B(n6567), .Z(n6591) );
  AND U7663 ( .A(a[201]), .B(b[3]), .Z(n6590) );
  XOR U7664 ( .A(n6591), .B(n6590), .Z(n6593) );
  XOR U7665 ( .A(n6592), .B(n6593), .Z(n6581) );
  NANDN U7666 ( .A(n6570), .B(n6569), .Z(n6574) );
  OR U7667 ( .A(n6572), .B(n6571), .Z(n6573) );
  AND U7668 ( .A(n6574), .B(n6573), .Z(n6580) );
  XOR U7669 ( .A(n6581), .B(n6580), .Z(n6583) );
  XOR U7670 ( .A(n6582), .B(n6583), .Z(n6596) );
  XNOR U7671 ( .A(n6596), .B(sreg[1225]), .Z(n6598) );
  NANDN U7672 ( .A(n6575), .B(sreg[1224]), .Z(n6579) );
  NAND U7673 ( .A(n6577), .B(n6576), .Z(n6578) );
  NAND U7674 ( .A(n6579), .B(n6578), .Z(n6597) );
  XOR U7675 ( .A(n6598), .B(n6597), .Z(c[1225]) );
  NANDN U7676 ( .A(n6581), .B(n6580), .Z(n6585) );
  OR U7677 ( .A(n6583), .B(n6582), .Z(n6584) );
  AND U7678 ( .A(n6585), .B(n6584), .Z(n6603) );
  XOR U7679 ( .A(a[204]), .B(n2205), .Z(n6607) );
  AND U7680 ( .A(a[206]), .B(b[0]), .Z(n6587) );
  XNOR U7681 ( .A(n6587), .B(n2175), .Z(n6589) );
  NANDN U7682 ( .A(b[0]), .B(a[205]), .Z(n6588) );
  NAND U7683 ( .A(n6589), .B(n6588), .Z(n6612) );
  AND U7684 ( .A(a[202]), .B(b[3]), .Z(n6611) );
  XOR U7685 ( .A(n6612), .B(n6611), .Z(n6614) );
  XOR U7686 ( .A(n6613), .B(n6614), .Z(n6602) );
  NANDN U7687 ( .A(n6591), .B(n6590), .Z(n6595) );
  OR U7688 ( .A(n6593), .B(n6592), .Z(n6594) );
  AND U7689 ( .A(n6595), .B(n6594), .Z(n6601) );
  XOR U7690 ( .A(n6602), .B(n6601), .Z(n6604) );
  XOR U7691 ( .A(n6603), .B(n6604), .Z(n6617) );
  XNOR U7692 ( .A(n6617), .B(sreg[1226]), .Z(n6619) );
  NANDN U7693 ( .A(n6596), .B(sreg[1225]), .Z(n6600) );
  NAND U7694 ( .A(n6598), .B(n6597), .Z(n6599) );
  NAND U7695 ( .A(n6600), .B(n6599), .Z(n6618) );
  XOR U7696 ( .A(n6619), .B(n6618), .Z(c[1226]) );
  NANDN U7697 ( .A(n6602), .B(n6601), .Z(n6606) );
  OR U7698 ( .A(n6604), .B(n6603), .Z(n6605) );
  AND U7699 ( .A(n6606), .B(n6605), .Z(n6624) );
  XOR U7700 ( .A(a[205]), .B(n2205), .Z(n6628) );
  AND U7701 ( .A(a[207]), .B(b[0]), .Z(n6608) );
  XNOR U7702 ( .A(n6608), .B(n2175), .Z(n6610) );
  NANDN U7703 ( .A(b[0]), .B(a[206]), .Z(n6609) );
  NAND U7704 ( .A(n6610), .B(n6609), .Z(n6633) );
  AND U7705 ( .A(a[203]), .B(b[3]), .Z(n6632) );
  XOR U7706 ( .A(n6633), .B(n6632), .Z(n6635) );
  XOR U7707 ( .A(n6634), .B(n6635), .Z(n6623) );
  NANDN U7708 ( .A(n6612), .B(n6611), .Z(n6616) );
  OR U7709 ( .A(n6614), .B(n6613), .Z(n6615) );
  AND U7710 ( .A(n6616), .B(n6615), .Z(n6622) );
  XOR U7711 ( .A(n6623), .B(n6622), .Z(n6625) );
  XOR U7712 ( .A(n6624), .B(n6625), .Z(n6638) );
  XNOR U7713 ( .A(n6638), .B(sreg[1227]), .Z(n6640) );
  NANDN U7714 ( .A(n6617), .B(sreg[1226]), .Z(n6621) );
  NAND U7715 ( .A(n6619), .B(n6618), .Z(n6620) );
  NAND U7716 ( .A(n6621), .B(n6620), .Z(n6639) );
  XOR U7717 ( .A(n6640), .B(n6639), .Z(c[1227]) );
  NANDN U7718 ( .A(n6623), .B(n6622), .Z(n6627) );
  OR U7719 ( .A(n6625), .B(n6624), .Z(n6626) );
  AND U7720 ( .A(n6627), .B(n6626), .Z(n6645) );
  XOR U7721 ( .A(a[206]), .B(n2205), .Z(n6649) );
  AND U7722 ( .A(a[208]), .B(b[0]), .Z(n6629) );
  XNOR U7723 ( .A(n6629), .B(n2175), .Z(n6631) );
  NANDN U7724 ( .A(b[0]), .B(a[207]), .Z(n6630) );
  NAND U7725 ( .A(n6631), .B(n6630), .Z(n6654) );
  AND U7726 ( .A(a[204]), .B(b[3]), .Z(n6653) );
  XOR U7727 ( .A(n6654), .B(n6653), .Z(n6656) );
  XOR U7728 ( .A(n6655), .B(n6656), .Z(n6644) );
  NANDN U7729 ( .A(n6633), .B(n6632), .Z(n6637) );
  OR U7730 ( .A(n6635), .B(n6634), .Z(n6636) );
  AND U7731 ( .A(n6637), .B(n6636), .Z(n6643) );
  XOR U7732 ( .A(n6644), .B(n6643), .Z(n6646) );
  XOR U7733 ( .A(n6645), .B(n6646), .Z(n6659) );
  XNOR U7734 ( .A(n6659), .B(sreg[1228]), .Z(n6661) );
  NANDN U7735 ( .A(n6638), .B(sreg[1227]), .Z(n6642) );
  NAND U7736 ( .A(n6640), .B(n6639), .Z(n6641) );
  NAND U7737 ( .A(n6642), .B(n6641), .Z(n6660) );
  XOR U7738 ( .A(n6661), .B(n6660), .Z(c[1228]) );
  NANDN U7739 ( .A(n6644), .B(n6643), .Z(n6648) );
  OR U7740 ( .A(n6646), .B(n6645), .Z(n6647) );
  AND U7741 ( .A(n6648), .B(n6647), .Z(n6666) );
  XOR U7742 ( .A(a[207]), .B(n2205), .Z(n6670) );
  AND U7743 ( .A(a[205]), .B(b[3]), .Z(n6674) );
  AND U7744 ( .A(a[209]), .B(b[0]), .Z(n6650) );
  XNOR U7745 ( .A(n6650), .B(n2175), .Z(n6652) );
  NANDN U7746 ( .A(b[0]), .B(a[208]), .Z(n6651) );
  NAND U7747 ( .A(n6652), .B(n6651), .Z(n6675) );
  XOR U7748 ( .A(n6674), .B(n6675), .Z(n6677) );
  XOR U7749 ( .A(n6676), .B(n6677), .Z(n6665) );
  NANDN U7750 ( .A(n6654), .B(n6653), .Z(n6658) );
  OR U7751 ( .A(n6656), .B(n6655), .Z(n6657) );
  AND U7752 ( .A(n6658), .B(n6657), .Z(n6664) );
  XOR U7753 ( .A(n6665), .B(n6664), .Z(n6667) );
  XOR U7754 ( .A(n6666), .B(n6667), .Z(n6680) );
  XNOR U7755 ( .A(n6680), .B(sreg[1229]), .Z(n6682) );
  NANDN U7756 ( .A(n6659), .B(sreg[1228]), .Z(n6663) );
  NAND U7757 ( .A(n6661), .B(n6660), .Z(n6662) );
  NAND U7758 ( .A(n6663), .B(n6662), .Z(n6681) );
  XOR U7759 ( .A(n6682), .B(n6681), .Z(c[1229]) );
  NANDN U7760 ( .A(n6665), .B(n6664), .Z(n6669) );
  OR U7761 ( .A(n6667), .B(n6666), .Z(n6668) );
  AND U7762 ( .A(n6669), .B(n6668), .Z(n6687) );
  XOR U7763 ( .A(a[208]), .B(n2205), .Z(n6691) );
  AND U7764 ( .A(a[206]), .B(b[3]), .Z(n6695) );
  AND U7765 ( .A(a[210]), .B(b[0]), .Z(n6671) );
  XNOR U7766 ( .A(n6671), .B(n2175), .Z(n6673) );
  NANDN U7767 ( .A(b[0]), .B(a[209]), .Z(n6672) );
  NAND U7768 ( .A(n6673), .B(n6672), .Z(n6696) );
  XOR U7769 ( .A(n6695), .B(n6696), .Z(n6698) );
  XOR U7770 ( .A(n6697), .B(n6698), .Z(n6686) );
  NANDN U7771 ( .A(n6675), .B(n6674), .Z(n6679) );
  OR U7772 ( .A(n6677), .B(n6676), .Z(n6678) );
  AND U7773 ( .A(n6679), .B(n6678), .Z(n6685) );
  XOR U7774 ( .A(n6686), .B(n6685), .Z(n6688) );
  XOR U7775 ( .A(n6687), .B(n6688), .Z(n6701) );
  XNOR U7776 ( .A(n6701), .B(sreg[1230]), .Z(n6703) );
  NANDN U7777 ( .A(n6680), .B(sreg[1229]), .Z(n6684) );
  NAND U7778 ( .A(n6682), .B(n6681), .Z(n6683) );
  NAND U7779 ( .A(n6684), .B(n6683), .Z(n6702) );
  XOR U7780 ( .A(n6703), .B(n6702), .Z(c[1230]) );
  NANDN U7781 ( .A(n6686), .B(n6685), .Z(n6690) );
  OR U7782 ( .A(n6688), .B(n6687), .Z(n6689) );
  AND U7783 ( .A(n6690), .B(n6689), .Z(n6708) );
  XOR U7784 ( .A(a[209]), .B(n2206), .Z(n6712) );
  AND U7785 ( .A(a[211]), .B(b[0]), .Z(n6692) );
  XNOR U7786 ( .A(n6692), .B(n2175), .Z(n6694) );
  NANDN U7787 ( .A(b[0]), .B(a[210]), .Z(n6693) );
  NAND U7788 ( .A(n6694), .B(n6693), .Z(n6717) );
  AND U7789 ( .A(a[207]), .B(b[3]), .Z(n6716) );
  XOR U7790 ( .A(n6717), .B(n6716), .Z(n6719) );
  XOR U7791 ( .A(n6718), .B(n6719), .Z(n6707) );
  NANDN U7792 ( .A(n6696), .B(n6695), .Z(n6700) );
  OR U7793 ( .A(n6698), .B(n6697), .Z(n6699) );
  AND U7794 ( .A(n6700), .B(n6699), .Z(n6706) );
  XOR U7795 ( .A(n6707), .B(n6706), .Z(n6709) );
  XOR U7796 ( .A(n6708), .B(n6709), .Z(n6722) );
  XNOR U7797 ( .A(n6722), .B(sreg[1231]), .Z(n6724) );
  NANDN U7798 ( .A(n6701), .B(sreg[1230]), .Z(n6705) );
  NAND U7799 ( .A(n6703), .B(n6702), .Z(n6704) );
  NAND U7800 ( .A(n6705), .B(n6704), .Z(n6723) );
  XOR U7801 ( .A(n6724), .B(n6723), .Z(c[1231]) );
  NANDN U7802 ( .A(n6707), .B(n6706), .Z(n6711) );
  OR U7803 ( .A(n6709), .B(n6708), .Z(n6710) );
  AND U7804 ( .A(n6711), .B(n6710), .Z(n6729) );
  XOR U7805 ( .A(a[210]), .B(n2206), .Z(n6733) );
  AND U7806 ( .A(a[212]), .B(b[0]), .Z(n6713) );
  XNOR U7807 ( .A(n6713), .B(n2175), .Z(n6715) );
  NANDN U7808 ( .A(b[0]), .B(a[211]), .Z(n6714) );
  NAND U7809 ( .A(n6715), .B(n6714), .Z(n6738) );
  AND U7810 ( .A(a[208]), .B(b[3]), .Z(n6737) );
  XOR U7811 ( .A(n6738), .B(n6737), .Z(n6740) );
  XOR U7812 ( .A(n6739), .B(n6740), .Z(n6728) );
  NANDN U7813 ( .A(n6717), .B(n6716), .Z(n6721) );
  OR U7814 ( .A(n6719), .B(n6718), .Z(n6720) );
  AND U7815 ( .A(n6721), .B(n6720), .Z(n6727) );
  XOR U7816 ( .A(n6728), .B(n6727), .Z(n6730) );
  XOR U7817 ( .A(n6729), .B(n6730), .Z(n6743) );
  XNOR U7818 ( .A(n6743), .B(sreg[1232]), .Z(n6745) );
  NANDN U7819 ( .A(n6722), .B(sreg[1231]), .Z(n6726) );
  NAND U7820 ( .A(n6724), .B(n6723), .Z(n6725) );
  NAND U7821 ( .A(n6726), .B(n6725), .Z(n6744) );
  XOR U7822 ( .A(n6745), .B(n6744), .Z(c[1232]) );
  NANDN U7823 ( .A(n6728), .B(n6727), .Z(n6732) );
  OR U7824 ( .A(n6730), .B(n6729), .Z(n6731) );
  AND U7825 ( .A(n6732), .B(n6731), .Z(n6750) );
  XOR U7826 ( .A(a[211]), .B(n2206), .Z(n6754) );
  AND U7827 ( .A(a[209]), .B(b[3]), .Z(n6758) );
  AND U7828 ( .A(a[213]), .B(b[0]), .Z(n6734) );
  XNOR U7829 ( .A(n6734), .B(n2175), .Z(n6736) );
  NANDN U7830 ( .A(b[0]), .B(a[212]), .Z(n6735) );
  NAND U7831 ( .A(n6736), .B(n6735), .Z(n6759) );
  XOR U7832 ( .A(n6758), .B(n6759), .Z(n6761) );
  XOR U7833 ( .A(n6760), .B(n6761), .Z(n6749) );
  NANDN U7834 ( .A(n6738), .B(n6737), .Z(n6742) );
  OR U7835 ( .A(n6740), .B(n6739), .Z(n6741) );
  AND U7836 ( .A(n6742), .B(n6741), .Z(n6748) );
  XOR U7837 ( .A(n6749), .B(n6748), .Z(n6751) );
  XOR U7838 ( .A(n6750), .B(n6751), .Z(n6764) );
  XNOR U7839 ( .A(n6764), .B(sreg[1233]), .Z(n6766) );
  NANDN U7840 ( .A(n6743), .B(sreg[1232]), .Z(n6747) );
  NAND U7841 ( .A(n6745), .B(n6744), .Z(n6746) );
  NAND U7842 ( .A(n6747), .B(n6746), .Z(n6765) );
  XOR U7843 ( .A(n6766), .B(n6765), .Z(c[1233]) );
  NANDN U7844 ( .A(n6749), .B(n6748), .Z(n6753) );
  OR U7845 ( .A(n6751), .B(n6750), .Z(n6752) );
  AND U7846 ( .A(n6753), .B(n6752), .Z(n6771) );
  XOR U7847 ( .A(a[212]), .B(n2206), .Z(n6775) );
  AND U7848 ( .A(a[214]), .B(b[0]), .Z(n6755) );
  XNOR U7849 ( .A(n6755), .B(n2175), .Z(n6757) );
  NANDN U7850 ( .A(b[0]), .B(a[213]), .Z(n6756) );
  NAND U7851 ( .A(n6757), .B(n6756), .Z(n6780) );
  AND U7852 ( .A(a[210]), .B(b[3]), .Z(n6779) );
  XOR U7853 ( .A(n6780), .B(n6779), .Z(n6782) );
  XOR U7854 ( .A(n6781), .B(n6782), .Z(n6770) );
  NANDN U7855 ( .A(n6759), .B(n6758), .Z(n6763) );
  OR U7856 ( .A(n6761), .B(n6760), .Z(n6762) );
  AND U7857 ( .A(n6763), .B(n6762), .Z(n6769) );
  XOR U7858 ( .A(n6770), .B(n6769), .Z(n6772) );
  XOR U7859 ( .A(n6771), .B(n6772), .Z(n6785) );
  XNOR U7860 ( .A(n6785), .B(sreg[1234]), .Z(n6787) );
  NANDN U7861 ( .A(n6764), .B(sreg[1233]), .Z(n6768) );
  NAND U7862 ( .A(n6766), .B(n6765), .Z(n6767) );
  NAND U7863 ( .A(n6768), .B(n6767), .Z(n6786) );
  XOR U7864 ( .A(n6787), .B(n6786), .Z(c[1234]) );
  NANDN U7865 ( .A(n6770), .B(n6769), .Z(n6774) );
  OR U7866 ( .A(n6772), .B(n6771), .Z(n6773) );
  AND U7867 ( .A(n6774), .B(n6773), .Z(n6792) );
  XOR U7868 ( .A(a[213]), .B(n2206), .Z(n6796) );
  AND U7869 ( .A(a[215]), .B(b[0]), .Z(n6776) );
  XNOR U7870 ( .A(n6776), .B(n2175), .Z(n6778) );
  NANDN U7871 ( .A(b[0]), .B(a[214]), .Z(n6777) );
  NAND U7872 ( .A(n6778), .B(n6777), .Z(n6801) );
  AND U7873 ( .A(a[211]), .B(b[3]), .Z(n6800) );
  XOR U7874 ( .A(n6801), .B(n6800), .Z(n6803) );
  XOR U7875 ( .A(n6802), .B(n6803), .Z(n6791) );
  NANDN U7876 ( .A(n6780), .B(n6779), .Z(n6784) );
  OR U7877 ( .A(n6782), .B(n6781), .Z(n6783) );
  AND U7878 ( .A(n6784), .B(n6783), .Z(n6790) );
  XOR U7879 ( .A(n6791), .B(n6790), .Z(n6793) );
  XOR U7880 ( .A(n6792), .B(n6793), .Z(n6806) );
  XNOR U7881 ( .A(n6806), .B(sreg[1235]), .Z(n6808) );
  NANDN U7882 ( .A(n6785), .B(sreg[1234]), .Z(n6789) );
  NAND U7883 ( .A(n6787), .B(n6786), .Z(n6788) );
  NAND U7884 ( .A(n6789), .B(n6788), .Z(n6807) );
  XOR U7885 ( .A(n6808), .B(n6807), .Z(c[1235]) );
  NANDN U7886 ( .A(n6791), .B(n6790), .Z(n6795) );
  OR U7887 ( .A(n6793), .B(n6792), .Z(n6794) );
  AND U7888 ( .A(n6795), .B(n6794), .Z(n6813) );
  XOR U7889 ( .A(a[214]), .B(n2206), .Z(n6817) );
  AND U7890 ( .A(a[216]), .B(b[0]), .Z(n6797) );
  XNOR U7891 ( .A(n6797), .B(n2175), .Z(n6799) );
  NANDN U7892 ( .A(b[0]), .B(a[215]), .Z(n6798) );
  NAND U7893 ( .A(n6799), .B(n6798), .Z(n6822) );
  AND U7894 ( .A(a[212]), .B(b[3]), .Z(n6821) );
  XOR U7895 ( .A(n6822), .B(n6821), .Z(n6824) );
  XOR U7896 ( .A(n6823), .B(n6824), .Z(n6812) );
  NANDN U7897 ( .A(n6801), .B(n6800), .Z(n6805) );
  OR U7898 ( .A(n6803), .B(n6802), .Z(n6804) );
  AND U7899 ( .A(n6805), .B(n6804), .Z(n6811) );
  XOR U7900 ( .A(n6812), .B(n6811), .Z(n6814) );
  XOR U7901 ( .A(n6813), .B(n6814), .Z(n6827) );
  XNOR U7902 ( .A(n6827), .B(sreg[1236]), .Z(n6829) );
  NANDN U7903 ( .A(n6806), .B(sreg[1235]), .Z(n6810) );
  NAND U7904 ( .A(n6808), .B(n6807), .Z(n6809) );
  NAND U7905 ( .A(n6810), .B(n6809), .Z(n6828) );
  XOR U7906 ( .A(n6829), .B(n6828), .Z(c[1236]) );
  NANDN U7907 ( .A(n6812), .B(n6811), .Z(n6816) );
  OR U7908 ( .A(n6814), .B(n6813), .Z(n6815) );
  AND U7909 ( .A(n6816), .B(n6815), .Z(n6835) );
  XOR U7910 ( .A(a[215]), .B(n2206), .Z(n6836) );
  AND U7911 ( .A(b[0]), .B(a[217]), .Z(n6818) );
  XOR U7912 ( .A(b[1]), .B(n6818), .Z(n6820) );
  NANDN U7913 ( .A(b[0]), .B(a[216]), .Z(n6819) );
  AND U7914 ( .A(n6820), .B(n6819), .Z(n6840) );
  AND U7915 ( .A(a[213]), .B(b[3]), .Z(n6841) );
  XOR U7916 ( .A(n6840), .B(n6841), .Z(n6842) );
  XNOR U7917 ( .A(n6843), .B(n6842), .Z(n6832) );
  NANDN U7918 ( .A(n6822), .B(n6821), .Z(n6826) );
  OR U7919 ( .A(n6824), .B(n6823), .Z(n6825) );
  AND U7920 ( .A(n6826), .B(n6825), .Z(n6833) );
  XNOR U7921 ( .A(n6832), .B(n6833), .Z(n6834) );
  XNOR U7922 ( .A(n6835), .B(n6834), .Z(n6846) );
  XNOR U7923 ( .A(n6846), .B(sreg[1237]), .Z(n6848) );
  NANDN U7924 ( .A(n6827), .B(sreg[1236]), .Z(n6831) );
  NAND U7925 ( .A(n6829), .B(n6828), .Z(n6830) );
  NAND U7926 ( .A(n6831), .B(n6830), .Z(n6847) );
  XOR U7927 ( .A(n6848), .B(n6847), .Z(c[1237]) );
  XOR U7928 ( .A(a[216]), .B(n2207), .Z(n6855) );
  AND U7929 ( .A(a[218]), .B(b[0]), .Z(n6837) );
  XNOR U7930 ( .A(n6837), .B(n2175), .Z(n6839) );
  NANDN U7931 ( .A(b[0]), .B(a[217]), .Z(n6838) );
  NAND U7932 ( .A(n6839), .B(n6838), .Z(n6860) );
  AND U7933 ( .A(a[214]), .B(b[3]), .Z(n6859) );
  XOR U7934 ( .A(n6860), .B(n6859), .Z(n6862) );
  XOR U7935 ( .A(n6861), .B(n6862), .Z(n6850) );
  NAND U7936 ( .A(n6841), .B(n6840), .Z(n6845) );
  NANDN U7937 ( .A(n6843), .B(n6842), .Z(n6844) );
  AND U7938 ( .A(n6845), .B(n6844), .Z(n6849) );
  XOR U7939 ( .A(n6850), .B(n6849), .Z(n6852) );
  XOR U7940 ( .A(n6851), .B(n6852), .Z(n6865) );
  XNOR U7941 ( .A(n6865), .B(sreg[1238]), .Z(n6867) );
  XOR U7942 ( .A(n6867), .B(n6866), .Z(c[1238]) );
  NANDN U7943 ( .A(n6850), .B(n6849), .Z(n6854) );
  OR U7944 ( .A(n6852), .B(n6851), .Z(n6853) );
  AND U7945 ( .A(n6854), .B(n6853), .Z(n6872) );
  XOR U7946 ( .A(a[217]), .B(n2207), .Z(n6876) );
  AND U7947 ( .A(a[219]), .B(b[0]), .Z(n6856) );
  XNOR U7948 ( .A(n6856), .B(n2175), .Z(n6858) );
  NANDN U7949 ( .A(b[0]), .B(a[218]), .Z(n6857) );
  NAND U7950 ( .A(n6858), .B(n6857), .Z(n6881) );
  AND U7951 ( .A(a[215]), .B(b[3]), .Z(n6880) );
  XOR U7952 ( .A(n6881), .B(n6880), .Z(n6883) );
  XOR U7953 ( .A(n6882), .B(n6883), .Z(n6871) );
  NANDN U7954 ( .A(n6860), .B(n6859), .Z(n6864) );
  OR U7955 ( .A(n6862), .B(n6861), .Z(n6863) );
  AND U7956 ( .A(n6864), .B(n6863), .Z(n6870) );
  XOR U7957 ( .A(n6871), .B(n6870), .Z(n6873) );
  XOR U7958 ( .A(n6872), .B(n6873), .Z(n6886) );
  XNOR U7959 ( .A(n6886), .B(sreg[1239]), .Z(n6888) );
  NANDN U7960 ( .A(n6865), .B(sreg[1238]), .Z(n6869) );
  NAND U7961 ( .A(n6867), .B(n6866), .Z(n6868) );
  NAND U7962 ( .A(n6869), .B(n6868), .Z(n6887) );
  XOR U7963 ( .A(n6888), .B(n6887), .Z(c[1239]) );
  NANDN U7964 ( .A(n6871), .B(n6870), .Z(n6875) );
  OR U7965 ( .A(n6873), .B(n6872), .Z(n6874) );
  AND U7966 ( .A(n6875), .B(n6874), .Z(n6893) );
  XOR U7967 ( .A(a[218]), .B(n2207), .Z(n6897) );
  AND U7968 ( .A(a[220]), .B(b[0]), .Z(n6877) );
  XNOR U7969 ( .A(n6877), .B(n2175), .Z(n6879) );
  NANDN U7970 ( .A(b[0]), .B(a[219]), .Z(n6878) );
  NAND U7971 ( .A(n6879), .B(n6878), .Z(n6902) );
  AND U7972 ( .A(a[216]), .B(b[3]), .Z(n6901) );
  XOR U7973 ( .A(n6902), .B(n6901), .Z(n6904) );
  XOR U7974 ( .A(n6903), .B(n6904), .Z(n6892) );
  NANDN U7975 ( .A(n6881), .B(n6880), .Z(n6885) );
  OR U7976 ( .A(n6883), .B(n6882), .Z(n6884) );
  AND U7977 ( .A(n6885), .B(n6884), .Z(n6891) );
  XOR U7978 ( .A(n6892), .B(n6891), .Z(n6894) );
  XOR U7979 ( .A(n6893), .B(n6894), .Z(n6907) );
  XNOR U7980 ( .A(n6907), .B(sreg[1240]), .Z(n6909) );
  NANDN U7981 ( .A(n6886), .B(sreg[1239]), .Z(n6890) );
  NAND U7982 ( .A(n6888), .B(n6887), .Z(n6889) );
  NAND U7983 ( .A(n6890), .B(n6889), .Z(n6908) );
  XOR U7984 ( .A(n6909), .B(n6908), .Z(c[1240]) );
  NANDN U7985 ( .A(n6892), .B(n6891), .Z(n6896) );
  OR U7986 ( .A(n6894), .B(n6893), .Z(n6895) );
  AND U7987 ( .A(n6896), .B(n6895), .Z(n6914) );
  XOR U7988 ( .A(a[219]), .B(n2207), .Z(n6918) );
  AND U7989 ( .A(a[217]), .B(b[3]), .Z(n6922) );
  AND U7990 ( .A(a[221]), .B(b[0]), .Z(n6898) );
  XNOR U7991 ( .A(n6898), .B(n2175), .Z(n6900) );
  NANDN U7992 ( .A(b[0]), .B(a[220]), .Z(n6899) );
  NAND U7993 ( .A(n6900), .B(n6899), .Z(n6923) );
  XOR U7994 ( .A(n6922), .B(n6923), .Z(n6925) );
  XOR U7995 ( .A(n6924), .B(n6925), .Z(n6913) );
  NANDN U7996 ( .A(n6902), .B(n6901), .Z(n6906) );
  OR U7997 ( .A(n6904), .B(n6903), .Z(n6905) );
  AND U7998 ( .A(n6906), .B(n6905), .Z(n6912) );
  XOR U7999 ( .A(n6913), .B(n6912), .Z(n6915) );
  XOR U8000 ( .A(n6914), .B(n6915), .Z(n6928) );
  XNOR U8001 ( .A(n6928), .B(sreg[1241]), .Z(n6930) );
  NANDN U8002 ( .A(n6907), .B(sreg[1240]), .Z(n6911) );
  NAND U8003 ( .A(n6909), .B(n6908), .Z(n6910) );
  NAND U8004 ( .A(n6911), .B(n6910), .Z(n6929) );
  XOR U8005 ( .A(n6930), .B(n6929), .Z(c[1241]) );
  NANDN U8006 ( .A(n6913), .B(n6912), .Z(n6917) );
  OR U8007 ( .A(n6915), .B(n6914), .Z(n6916) );
  AND U8008 ( .A(n6917), .B(n6916), .Z(n6936) );
  XOR U8009 ( .A(a[220]), .B(n2207), .Z(n6937) );
  AND U8010 ( .A(b[0]), .B(a[222]), .Z(n6919) );
  XOR U8011 ( .A(b[1]), .B(n6919), .Z(n6921) );
  NANDN U8012 ( .A(b[0]), .B(a[221]), .Z(n6920) );
  AND U8013 ( .A(n6921), .B(n6920), .Z(n6941) );
  AND U8014 ( .A(a[218]), .B(b[3]), .Z(n6942) );
  XOR U8015 ( .A(n6941), .B(n6942), .Z(n6943) );
  XNOR U8016 ( .A(n6944), .B(n6943), .Z(n6933) );
  NANDN U8017 ( .A(n6923), .B(n6922), .Z(n6927) );
  OR U8018 ( .A(n6925), .B(n6924), .Z(n6926) );
  AND U8019 ( .A(n6927), .B(n6926), .Z(n6934) );
  XNOR U8020 ( .A(n6933), .B(n6934), .Z(n6935) );
  XNOR U8021 ( .A(n6936), .B(n6935), .Z(n6947) );
  XNOR U8022 ( .A(n6947), .B(sreg[1242]), .Z(n6949) );
  NANDN U8023 ( .A(n6928), .B(sreg[1241]), .Z(n6932) );
  NAND U8024 ( .A(n6930), .B(n6929), .Z(n6931) );
  NAND U8025 ( .A(n6932), .B(n6931), .Z(n6948) );
  XOR U8026 ( .A(n6949), .B(n6948), .Z(c[1242]) );
  XOR U8027 ( .A(a[221]), .B(n2207), .Z(n6956) );
  AND U8028 ( .A(a[223]), .B(b[0]), .Z(n6938) );
  XNOR U8029 ( .A(n6938), .B(n2175), .Z(n6940) );
  NANDN U8030 ( .A(b[0]), .B(a[222]), .Z(n6939) );
  NAND U8031 ( .A(n6940), .B(n6939), .Z(n6961) );
  AND U8032 ( .A(a[219]), .B(b[3]), .Z(n6960) );
  XOR U8033 ( .A(n6961), .B(n6960), .Z(n6963) );
  XOR U8034 ( .A(n6962), .B(n6963), .Z(n6951) );
  NAND U8035 ( .A(n6942), .B(n6941), .Z(n6946) );
  NANDN U8036 ( .A(n6944), .B(n6943), .Z(n6945) );
  AND U8037 ( .A(n6946), .B(n6945), .Z(n6950) );
  XOR U8038 ( .A(n6951), .B(n6950), .Z(n6953) );
  XOR U8039 ( .A(n6952), .B(n6953), .Z(n6966) );
  XNOR U8040 ( .A(n6966), .B(sreg[1243]), .Z(n6968) );
  XOR U8041 ( .A(n6968), .B(n6967), .Z(c[1243]) );
  NANDN U8042 ( .A(n6951), .B(n6950), .Z(n6955) );
  OR U8043 ( .A(n6953), .B(n6952), .Z(n6954) );
  AND U8044 ( .A(n6955), .B(n6954), .Z(n6973) );
  XOR U8045 ( .A(a[222]), .B(n2207), .Z(n6977) );
  AND U8046 ( .A(a[224]), .B(b[0]), .Z(n6957) );
  XNOR U8047 ( .A(n6957), .B(n2175), .Z(n6959) );
  NANDN U8048 ( .A(b[0]), .B(a[223]), .Z(n6958) );
  NAND U8049 ( .A(n6959), .B(n6958), .Z(n6982) );
  AND U8050 ( .A(a[220]), .B(b[3]), .Z(n6981) );
  XOR U8051 ( .A(n6982), .B(n6981), .Z(n6984) );
  XOR U8052 ( .A(n6983), .B(n6984), .Z(n6972) );
  NANDN U8053 ( .A(n6961), .B(n6960), .Z(n6965) );
  OR U8054 ( .A(n6963), .B(n6962), .Z(n6964) );
  AND U8055 ( .A(n6965), .B(n6964), .Z(n6971) );
  XOR U8056 ( .A(n6972), .B(n6971), .Z(n6974) );
  XOR U8057 ( .A(n6973), .B(n6974), .Z(n6987) );
  XNOR U8058 ( .A(n6987), .B(sreg[1244]), .Z(n6989) );
  NANDN U8059 ( .A(n6966), .B(sreg[1243]), .Z(n6970) );
  NAND U8060 ( .A(n6968), .B(n6967), .Z(n6969) );
  NAND U8061 ( .A(n6970), .B(n6969), .Z(n6988) );
  XOR U8062 ( .A(n6989), .B(n6988), .Z(c[1244]) );
  NANDN U8063 ( .A(n6972), .B(n6971), .Z(n6976) );
  OR U8064 ( .A(n6974), .B(n6973), .Z(n6975) );
  AND U8065 ( .A(n6976), .B(n6975), .Z(n6994) );
  XOR U8066 ( .A(a[223]), .B(n2208), .Z(n6998) );
  AND U8067 ( .A(a[225]), .B(b[0]), .Z(n6978) );
  XNOR U8068 ( .A(n6978), .B(n2175), .Z(n6980) );
  NANDN U8069 ( .A(b[0]), .B(a[224]), .Z(n6979) );
  NAND U8070 ( .A(n6980), .B(n6979), .Z(n7003) );
  AND U8071 ( .A(a[221]), .B(b[3]), .Z(n7002) );
  XOR U8072 ( .A(n7003), .B(n7002), .Z(n7005) );
  XOR U8073 ( .A(n7004), .B(n7005), .Z(n6993) );
  NANDN U8074 ( .A(n6982), .B(n6981), .Z(n6986) );
  OR U8075 ( .A(n6984), .B(n6983), .Z(n6985) );
  AND U8076 ( .A(n6986), .B(n6985), .Z(n6992) );
  XOR U8077 ( .A(n6993), .B(n6992), .Z(n6995) );
  XOR U8078 ( .A(n6994), .B(n6995), .Z(n7008) );
  XNOR U8079 ( .A(n7008), .B(sreg[1245]), .Z(n7010) );
  NANDN U8080 ( .A(n6987), .B(sreg[1244]), .Z(n6991) );
  NAND U8081 ( .A(n6989), .B(n6988), .Z(n6990) );
  NAND U8082 ( .A(n6991), .B(n6990), .Z(n7009) );
  XOR U8083 ( .A(n7010), .B(n7009), .Z(c[1245]) );
  NANDN U8084 ( .A(n6993), .B(n6992), .Z(n6997) );
  OR U8085 ( .A(n6995), .B(n6994), .Z(n6996) );
  AND U8086 ( .A(n6997), .B(n6996), .Z(n7015) );
  XOR U8087 ( .A(a[224]), .B(n2208), .Z(n7019) );
  AND U8088 ( .A(a[226]), .B(b[0]), .Z(n6999) );
  XNOR U8089 ( .A(n6999), .B(n2175), .Z(n7001) );
  NANDN U8090 ( .A(b[0]), .B(a[225]), .Z(n7000) );
  NAND U8091 ( .A(n7001), .B(n7000), .Z(n7024) );
  AND U8092 ( .A(a[222]), .B(b[3]), .Z(n7023) );
  XOR U8093 ( .A(n7024), .B(n7023), .Z(n7026) );
  XOR U8094 ( .A(n7025), .B(n7026), .Z(n7014) );
  NANDN U8095 ( .A(n7003), .B(n7002), .Z(n7007) );
  OR U8096 ( .A(n7005), .B(n7004), .Z(n7006) );
  AND U8097 ( .A(n7007), .B(n7006), .Z(n7013) );
  XOR U8098 ( .A(n7014), .B(n7013), .Z(n7016) );
  XOR U8099 ( .A(n7015), .B(n7016), .Z(n7029) );
  XNOR U8100 ( .A(n7029), .B(sreg[1246]), .Z(n7031) );
  NANDN U8101 ( .A(n7008), .B(sreg[1245]), .Z(n7012) );
  NAND U8102 ( .A(n7010), .B(n7009), .Z(n7011) );
  NAND U8103 ( .A(n7012), .B(n7011), .Z(n7030) );
  XOR U8104 ( .A(n7031), .B(n7030), .Z(c[1246]) );
  NANDN U8105 ( .A(n7014), .B(n7013), .Z(n7018) );
  OR U8106 ( .A(n7016), .B(n7015), .Z(n7017) );
  AND U8107 ( .A(n7018), .B(n7017), .Z(n7036) );
  XOR U8108 ( .A(a[225]), .B(n2208), .Z(n7040) );
  AND U8109 ( .A(a[227]), .B(b[0]), .Z(n7020) );
  XNOR U8110 ( .A(n7020), .B(n2175), .Z(n7022) );
  NANDN U8111 ( .A(b[0]), .B(a[226]), .Z(n7021) );
  NAND U8112 ( .A(n7022), .B(n7021), .Z(n7045) );
  AND U8113 ( .A(a[223]), .B(b[3]), .Z(n7044) );
  XOR U8114 ( .A(n7045), .B(n7044), .Z(n7047) );
  XOR U8115 ( .A(n7046), .B(n7047), .Z(n7035) );
  NANDN U8116 ( .A(n7024), .B(n7023), .Z(n7028) );
  OR U8117 ( .A(n7026), .B(n7025), .Z(n7027) );
  AND U8118 ( .A(n7028), .B(n7027), .Z(n7034) );
  XOR U8119 ( .A(n7035), .B(n7034), .Z(n7037) );
  XOR U8120 ( .A(n7036), .B(n7037), .Z(n7050) );
  XNOR U8121 ( .A(n7050), .B(sreg[1247]), .Z(n7052) );
  NANDN U8122 ( .A(n7029), .B(sreg[1246]), .Z(n7033) );
  NAND U8123 ( .A(n7031), .B(n7030), .Z(n7032) );
  NAND U8124 ( .A(n7033), .B(n7032), .Z(n7051) );
  XOR U8125 ( .A(n7052), .B(n7051), .Z(c[1247]) );
  NANDN U8126 ( .A(n7035), .B(n7034), .Z(n7039) );
  OR U8127 ( .A(n7037), .B(n7036), .Z(n7038) );
  AND U8128 ( .A(n7039), .B(n7038), .Z(n7057) );
  XOR U8129 ( .A(a[226]), .B(n2208), .Z(n7061) );
  AND U8130 ( .A(a[228]), .B(b[0]), .Z(n7041) );
  XNOR U8131 ( .A(n7041), .B(n2175), .Z(n7043) );
  NANDN U8132 ( .A(b[0]), .B(a[227]), .Z(n7042) );
  NAND U8133 ( .A(n7043), .B(n7042), .Z(n7066) );
  AND U8134 ( .A(a[224]), .B(b[3]), .Z(n7065) );
  XOR U8135 ( .A(n7066), .B(n7065), .Z(n7068) );
  XOR U8136 ( .A(n7067), .B(n7068), .Z(n7056) );
  NANDN U8137 ( .A(n7045), .B(n7044), .Z(n7049) );
  OR U8138 ( .A(n7047), .B(n7046), .Z(n7048) );
  AND U8139 ( .A(n7049), .B(n7048), .Z(n7055) );
  XOR U8140 ( .A(n7056), .B(n7055), .Z(n7058) );
  XOR U8141 ( .A(n7057), .B(n7058), .Z(n7071) );
  XNOR U8142 ( .A(n7071), .B(sreg[1248]), .Z(n7073) );
  NANDN U8143 ( .A(n7050), .B(sreg[1247]), .Z(n7054) );
  NAND U8144 ( .A(n7052), .B(n7051), .Z(n7053) );
  NAND U8145 ( .A(n7054), .B(n7053), .Z(n7072) );
  XOR U8146 ( .A(n7073), .B(n7072), .Z(c[1248]) );
  NANDN U8147 ( .A(n7056), .B(n7055), .Z(n7060) );
  OR U8148 ( .A(n7058), .B(n7057), .Z(n7059) );
  AND U8149 ( .A(n7060), .B(n7059), .Z(n7078) );
  XOR U8150 ( .A(a[227]), .B(n2208), .Z(n7082) );
  AND U8151 ( .A(a[225]), .B(b[3]), .Z(n7086) );
  AND U8152 ( .A(a[229]), .B(b[0]), .Z(n7062) );
  XNOR U8153 ( .A(n7062), .B(n2175), .Z(n7064) );
  NANDN U8154 ( .A(b[0]), .B(a[228]), .Z(n7063) );
  NAND U8155 ( .A(n7064), .B(n7063), .Z(n7087) );
  XOR U8156 ( .A(n7086), .B(n7087), .Z(n7089) );
  XOR U8157 ( .A(n7088), .B(n7089), .Z(n7077) );
  NANDN U8158 ( .A(n7066), .B(n7065), .Z(n7070) );
  OR U8159 ( .A(n7068), .B(n7067), .Z(n7069) );
  AND U8160 ( .A(n7070), .B(n7069), .Z(n7076) );
  XOR U8161 ( .A(n7077), .B(n7076), .Z(n7079) );
  XOR U8162 ( .A(n7078), .B(n7079), .Z(n7092) );
  XNOR U8163 ( .A(n7092), .B(sreg[1249]), .Z(n7094) );
  NANDN U8164 ( .A(n7071), .B(sreg[1248]), .Z(n7075) );
  NAND U8165 ( .A(n7073), .B(n7072), .Z(n7074) );
  NAND U8166 ( .A(n7075), .B(n7074), .Z(n7093) );
  XOR U8167 ( .A(n7094), .B(n7093), .Z(c[1249]) );
  NANDN U8168 ( .A(n7077), .B(n7076), .Z(n7081) );
  OR U8169 ( .A(n7079), .B(n7078), .Z(n7080) );
  AND U8170 ( .A(n7081), .B(n7080), .Z(n7100) );
  XOR U8171 ( .A(a[228]), .B(n2208), .Z(n7101) );
  AND U8172 ( .A(b[0]), .B(a[230]), .Z(n7083) );
  XOR U8173 ( .A(b[1]), .B(n7083), .Z(n7085) );
  NANDN U8174 ( .A(b[0]), .B(a[229]), .Z(n7084) );
  AND U8175 ( .A(n7085), .B(n7084), .Z(n7105) );
  AND U8176 ( .A(a[226]), .B(b[3]), .Z(n7106) );
  XOR U8177 ( .A(n7105), .B(n7106), .Z(n7107) );
  XNOR U8178 ( .A(n7108), .B(n7107), .Z(n7097) );
  NANDN U8179 ( .A(n7087), .B(n7086), .Z(n7091) );
  OR U8180 ( .A(n7089), .B(n7088), .Z(n7090) );
  AND U8181 ( .A(n7091), .B(n7090), .Z(n7098) );
  XNOR U8182 ( .A(n7097), .B(n7098), .Z(n7099) );
  XNOR U8183 ( .A(n7100), .B(n7099), .Z(n7111) );
  XNOR U8184 ( .A(n7111), .B(sreg[1250]), .Z(n7113) );
  NANDN U8185 ( .A(n7092), .B(sreg[1249]), .Z(n7096) );
  NAND U8186 ( .A(n7094), .B(n7093), .Z(n7095) );
  NAND U8187 ( .A(n7096), .B(n7095), .Z(n7112) );
  XOR U8188 ( .A(n7113), .B(n7112), .Z(c[1250]) );
  XOR U8189 ( .A(a[229]), .B(n2208), .Z(n7120) );
  AND U8190 ( .A(a[231]), .B(b[0]), .Z(n7102) );
  XNOR U8191 ( .A(n7102), .B(n2175), .Z(n7104) );
  NANDN U8192 ( .A(b[0]), .B(a[230]), .Z(n7103) );
  NAND U8193 ( .A(n7104), .B(n7103), .Z(n7125) );
  AND U8194 ( .A(a[227]), .B(b[3]), .Z(n7124) );
  XOR U8195 ( .A(n7125), .B(n7124), .Z(n7127) );
  XOR U8196 ( .A(n7126), .B(n7127), .Z(n7115) );
  NAND U8197 ( .A(n7106), .B(n7105), .Z(n7110) );
  NANDN U8198 ( .A(n7108), .B(n7107), .Z(n7109) );
  AND U8199 ( .A(n7110), .B(n7109), .Z(n7114) );
  XOR U8200 ( .A(n7115), .B(n7114), .Z(n7117) );
  XOR U8201 ( .A(n7116), .B(n7117), .Z(n7130) );
  XNOR U8202 ( .A(n7130), .B(sreg[1251]), .Z(n7132) );
  XOR U8203 ( .A(n7132), .B(n7131), .Z(c[1251]) );
  NANDN U8204 ( .A(n7115), .B(n7114), .Z(n7119) );
  OR U8205 ( .A(n7117), .B(n7116), .Z(n7118) );
  AND U8206 ( .A(n7119), .B(n7118), .Z(n7137) );
  XOR U8207 ( .A(a[230]), .B(n2209), .Z(n7141) );
  AND U8208 ( .A(a[228]), .B(b[3]), .Z(n7145) );
  AND U8209 ( .A(a[232]), .B(b[0]), .Z(n7121) );
  XNOR U8210 ( .A(n7121), .B(n2175), .Z(n7123) );
  NANDN U8211 ( .A(b[0]), .B(a[231]), .Z(n7122) );
  NAND U8212 ( .A(n7123), .B(n7122), .Z(n7146) );
  XOR U8213 ( .A(n7145), .B(n7146), .Z(n7148) );
  XOR U8214 ( .A(n7147), .B(n7148), .Z(n7136) );
  NANDN U8215 ( .A(n7125), .B(n7124), .Z(n7129) );
  OR U8216 ( .A(n7127), .B(n7126), .Z(n7128) );
  AND U8217 ( .A(n7129), .B(n7128), .Z(n7135) );
  XOR U8218 ( .A(n7136), .B(n7135), .Z(n7138) );
  XOR U8219 ( .A(n7137), .B(n7138), .Z(n7151) );
  XNOR U8220 ( .A(n7151), .B(sreg[1252]), .Z(n7153) );
  NANDN U8221 ( .A(n7130), .B(sreg[1251]), .Z(n7134) );
  NAND U8222 ( .A(n7132), .B(n7131), .Z(n7133) );
  NAND U8223 ( .A(n7134), .B(n7133), .Z(n7152) );
  XOR U8224 ( .A(n7153), .B(n7152), .Z(c[1252]) );
  NANDN U8225 ( .A(n7136), .B(n7135), .Z(n7140) );
  OR U8226 ( .A(n7138), .B(n7137), .Z(n7139) );
  AND U8227 ( .A(n7140), .B(n7139), .Z(n7158) );
  XOR U8228 ( .A(a[231]), .B(n2209), .Z(n7162) );
  AND U8229 ( .A(a[233]), .B(b[0]), .Z(n7142) );
  XNOR U8230 ( .A(n7142), .B(n2175), .Z(n7144) );
  NANDN U8231 ( .A(b[0]), .B(a[232]), .Z(n7143) );
  NAND U8232 ( .A(n7144), .B(n7143), .Z(n7167) );
  AND U8233 ( .A(a[229]), .B(b[3]), .Z(n7166) );
  XOR U8234 ( .A(n7167), .B(n7166), .Z(n7169) );
  XOR U8235 ( .A(n7168), .B(n7169), .Z(n7157) );
  NANDN U8236 ( .A(n7146), .B(n7145), .Z(n7150) );
  OR U8237 ( .A(n7148), .B(n7147), .Z(n7149) );
  AND U8238 ( .A(n7150), .B(n7149), .Z(n7156) );
  XOR U8239 ( .A(n7157), .B(n7156), .Z(n7159) );
  XOR U8240 ( .A(n7158), .B(n7159), .Z(n7172) );
  XNOR U8241 ( .A(n7172), .B(sreg[1253]), .Z(n7174) );
  NANDN U8242 ( .A(n7151), .B(sreg[1252]), .Z(n7155) );
  NAND U8243 ( .A(n7153), .B(n7152), .Z(n7154) );
  NAND U8244 ( .A(n7155), .B(n7154), .Z(n7173) );
  XOR U8245 ( .A(n7174), .B(n7173), .Z(c[1253]) );
  NANDN U8246 ( .A(n7157), .B(n7156), .Z(n7161) );
  OR U8247 ( .A(n7159), .B(n7158), .Z(n7160) );
  AND U8248 ( .A(n7161), .B(n7160), .Z(n7179) );
  XOR U8249 ( .A(a[232]), .B(n2209), .Z(n7183) );
  AND U8250 ( .A(a[230]), .B(b[3]), .Z(n7187) );
  AND U8251 ( .A(a[234]), .B(b[0]), .Z(n7163) );
  XNOR U8252 ( .A(n7163), .B(n2175), .Z(n7165) );
  NANDN U8253 ( .A(b[0]), .B(a[233]), .Z(n7164) );
  NAND U8254 ( .A(n7165), .B(n7164), .Z(n7188) );
  XOR U8255 ( .A(n7187), .B(n7188), .Z(n7190) );
  XOR U8256 ( .A(n7189), .B(n7190), .Z(n7178) );
  NANDN U8257 ( .A(n7167), .B(n7166), .Z(n7171) );
  OR U8258 ( .A(n7169), .B(n7168), .Z(n7170) );
  AND U8259 ( .A(n7171), .B(n7170), .Z(n7177) );
  XOR U8260 ( .A(n7178), .B(n7177), .Z(n7180) );
  XOR U8261 ( .A(n7179), .B(n7180), .Z(n7193) );
  XNOR U8262 ( .A(n7193), .B(sreg[1254]), .Z(n7195) );
  NANDN U8263 ( .A(n7172), .B(sreg[1253]), .Z(n7176) );
  NAND U8264 ( .A(n7174), .B(n7173), .Z(n7175) );
  NAND U8265 ( .A(n7176), .B(n7175), .Z(n7194) );
  XOR U8266 ( .A(n7195), .B(n7194), .Z(c[1254]) );
  NANDN U8267 ( .A(n7178), .B(n7177), .Z(n7182) );
  OR U8268 ( .A(n7180), .B(n7179), .Z(n7181) );
  AND U8269 ( .A(n7182), .B(n7181), .Z(n7200) );
  XOR U8270 ( .A(a[233]), .B(n2209), .Z(n7204) );
  AND U8271 ( .A(a[231]), .B(b[3]), .Z(n7208) );
  AND U8272 ( .A(a[235]), .B(b[0]), .Z(n7184) );
  XNOR U8273 ( .A(n7184), .B(n2175), .Z(n7186) );
  NANDN U8274 ( .A(b[0]), .B(a[234]), .Z(n7185) );
  NAND U8275 ( .A(n7186), .B(n7185), .Z(n7209) );
  XOR U8276 ( .A(n7208), .B(n7209), .Z(n7211) );
  XOR U8277 ( .A(n7210), .B(n7211), .Z(n7199) );
  NANDN U8278 ( .A(n7188), .B(n7187), .Z(n7192) );
  OR U8279 ( .A(n7190), .B(n7189), .Z(n7191) );
  AND U8280 ( .A(n7192), .B(n7191), .Z(n7198) );
  XOR U8281 ( .A(n7199), .B(n7198), .Z(n7201) );
  XOR U8282 ( .A(n7200), .B(n7201), .Z(n7214) );
  XNOR U8283 ( .A(n7214), .B(sreg[1255]), .Z(n7216) );
  NANDN U8284 ( .A(n7193), .B(sreg[1254]), .Z(n7197) );
  NAND U8285 ( .A(n7195), .B(n7194), .Z(n7196) );
  NAND U8286 ( .A(n7197), .B(n7196), .Z(n7215) );
  XOR U8287 ( .A(n7216), .B(n7215), .Z(c[1255]) );
  NANDN U8288 ( .A(n7199), .B(n7198), .Z(n7203) );
  OR U8289 ( .A(n7201), .B(n7200), .Z(n7202) );
  AND U8290 ( .A(n7203), .B(n7202), .Z(n7221) );
  XOR U8291 ( .A(a[234]), .B(n2209), .Z(n7225) );
  AND U8292 ( .A(a[236]), .B(b[0]), .Z(n7205) );
  XNOR U8293 ( .A(n7205), .B(n2175), .Z(n7207) );
  NANDN U8294 ( .A(b[0]), .B(a[235]), .Z(n7206) );
  NAND U8295 ( .A(n7207), .B(n7206), .Z(n7230) );
  AND U8296 ( .A(a[232]), .B(b[3]), .Z(n7229) );
  XOR U8297 ( .A(n7230), .B(n7229), .Z(n7232) );
  XOR U8298 ( .A(n7231), .B(n7232), .Z(n7220) );
  NANDN U8299 ( .A(n7209), .B(n7208), .Z(n7213) );
  OR U8300 ( .A(n7211), .B(n7210), .Z(n7212) );
  AND U8301 ( .A(n7213), .B(n7212), .Z(n7219) );
  XOR U8302 ( .A(n7220), .B(n7219), .Z(n7222) );
  XOR U8303 ( .A(n7221), .B(n7222), .Z(n7235) );
  XNOR U8304 ( .A(n7235), .B(sreg[1256]), .Z(n7237) );
  NANDN U8305 ( .A(n7214), .B(sreg[1255]), .Z(n7218) );
  NAND U8306 ( .A(n7216), .B(n7215), .Z(n7217) );
  NAND U8307 ( .A(n7218), .B(n7217), .Z(n7236) );
  XOR U8308 ( .A(n7237), .B(n7236), .Z(c[1256]) );
  NANDN U8309 ( .A(n7220), .B(n7219), .Z(n7224) );
  OR U8310 ( .A(n7222), .B(n7221), .Z(n7223) );
  AND U8311 ( .A(n7224), .B(n7223), .Z(n7242) );
  XOR U8312 ( .A(a[235]), .B(n2209), .Z(n7246) );
  AND U8313 ( .A(a[237]), .B(b[0]), .Z(n7226) );
  XNOR U8314 ( .A(n7226), .B(n2175), .Z(n7228) );
  NANDN U8315 ( .A(b[0]), .B(a[236]), .Z(n7227) );
  NAND U8316 ( .A(n7228), .B(n7227), .Z(n7251) );
  AND U8317 ( .A(a[233]), .B(b[3]), .Z(n7250) );
  XOR U8318 ( .A(n7251), .B(n7250), .Z(n7253) );
  XOR U8319 ( .A(n7252), .B(n7253), .Z(n7241) );
  NANDN U8320 ( .A(n7230), .B(n7229), .Z(n7234) );
  OR U8321 ( .A(n7232), .B(n7231), .Z(n7233) );
  AND U8322 ( .A(n7234), .B(n7233), .Z(n7240) );
  XOR U8323 ( .A(n7241), .B(n7240), .Z(n7243) );
  XOR U8324 ( .A(n7242), .B(n7243), .Z(n7256) );
  XNOR U8325 ( .A(n7256), .B(sreg[1257]), .Z(n7258) );
  NANDN U8326 ( .A(n7235), .B(sreg[1256]), .Z(n7239) );
  NAND U8327 ( .A(n7237), .B(n7236), .Z(n7238) );
  NAND U8328 ( .A(n7239), .B(n7238), .Z(n7257) );
  XOR U8329 ( .A(n7258), .B(n7257), .Z(c[1257]) );
  NANDN U8330 ( .A(n7241), .B(n7240), .Z(n7245) );
  OR U8331 ( .A(n7243), .B(n7242), .Z(n7244) );
  AND U8332 ( .A(n7245), .B(n7244), .Z(n7263) );
  XOR U8333 ( .A(a[236]), .B(n2209), .Z(n7267) );
  AND U8334 ( .A(a[238]), .B(b[0]), .Z(n7247) );
  XNOR U8335 ( .A(n7247), .B(n2175), .Z(n7249) );
  NANDN U8336 ( .A(b[0]), .B(a[237]), .Z(n7248) );
  NAND U8337 ( .A(n7249), .B(n7248), .Z(n7272) );
  AND U8338 ( .A(a[234]), .B(b[3]), .Z(n7271) );
  XOR U8339 ( .A(n7272), .B(n7271), .Z(n7274) );
  XOR U8340 ( .A(n7273), .B(n7274), .Z(n7262) );
  NANDN U8341 ( .A(n7251), .B(n7250), .Z(n7255) );
  OR U8342 ( .A(n7253), .B(n7252), .Z(n7254) );
  AND U8343 ( .A(n7255), .B(n7254), .Z(n7261) );
  XOR U8344 ( .A(n7262), .B(n7261), .Z(n7264) );
  XOR U8345 ( .A(n7263), .B(n7264), .Z(n7277) );
  XNOR U8346 ( .A(n7277), .B(sreg[1258]), .Z(n7279) );
  NANDN U8347 ( .A(n7256), .B(sreg[1257]), .Z(n7260) );
  NAND U8348 ( .A(n7258), .B(n7257), .Z(n7259) );
  NAND U8349 ( .A(n7260), .B(n7259), .Z(n7278) );
  XOR U8350 ( .A(n7279), .B(n7278), .Z(c[1258]) );
  NANDN U8351 ( .A(n7262), .B(n7261), .Z(n7266) );
  OR U8352 ( .A(n7264), .B(n7263), .Z(n7265) );
  AND U8353 ( .A(n7266), .B(n7265), .Z(n7284) );
  XOR U8354 ( .A(a[237]), .B(n2210), .Z(n7288) );
  AND U8355 ( .A(a[235]), .B(b[3]), .Z(n7292) );
  AND U8356 ( .A(a[239]), .B(b[0]), .Z(n7268) );
  XNOR U8357 ( .A(n7268), .B(n2175), .Z(n7270) );
  NANDN U8358 ( .A(b[0]), .B(a[238]), .Z(n7269) );
  NAND U8359 ( .A(n7270), .B(n7269), .Z(n7293) );
  XOR U8360 ( .A(n7292), .B(n7293), .Z(n7295) );
  XOR U8361 ( .A(n7294), .B(n7295), .Z(n7283) );
  NANDN U8362 ( .A(n7272), .B(n7271), .Z(n7276) );
  OR U8363 ( .A(n7274), .B(n7273), .Z(n7275) );
  AND U8364 ( .A(n7276), .B(n7275), .Z(n7282) );
  XOR U8365 ( .A(n7283), .B(n7282), .Z(n7285) );
  XOR U8366 ( .A(n7284), .B(n7285), .Z(n7298) );
  XNOR U8367 ( .A(n7298), .B(sreg[1259]), .Z(n7300) );
  NANDN U8368 ( .A(n7277), .B(sreg[1258]), .Z(n7281) );
  NAND U8369 ( .A(n7279), .B(n7278), .Z(n7280) );
  NAND U8370 ( .A(n7281), .B(n7280), .Z(n7299) );
  XOR U8371 ( .A(n7300), .B(n7299), .Z(c[1259]) );
  NANDN U8372 ( .A(n7283), .B(n7282), .Z(n7287) );
  OR U8373 ( .A(n7285), .B(n7284), .Z(n7286) );
  AND U8374 ( .A(n7287), .B(n7286), .Z(n7305) );
  XOR U8375 ( .A(a[238]), .B(n2210), .Z(n7309) );
  AND U8376 ( .A(a[240]), .B(b[0]), .Z(n7289) );
  XNOR U8377 ( .A(n7289), .B(n2175), .Z(n7291) );
  NANDN U8378 ( .A(b[0]), .B(a[239]), .Z(n7290) );
  NAND U8379 ( .A(n7291), .B(n7290), .Z(n7314) );
  AND U8380 ( .A(a[236]), .B(b[3]), .Z(n7313) );
  XOR U8381 ( .A(n7314), .B(n7313), .Z(n7316) );
  XOR U8382 ( .A(n7315), .B(n7316), .Z(n7304) );
  NANDN U8383 ( .A(n7293), .B(n7292), .Z(n7297) );
  OR U8384 ( .A(n7295), .B(n7294), .Z(n7296) );
  AND U8385 ( .A(n7297), .B(n7296), .Z(n7303) );
  XOR U8386 ( .A(n7304), .B(n7303), .Z(n7306) );
  XOR U8387 ( .A(n7305), .B(n7306), .Z(n7319) );
  XNOR U8388 ( .A(n7319), .B(sreg[1260]), .Z(n7321) );
  NANDN U8389 ( .A(n7298), .B(sreg[1259]), .Z(n7302) );
  NAND U8390 ( .A(n7300), .B(n7299), .Z(n7301) );
  NAND U8391 ( .A(n7302), .B(n7301), .Z(n7320) );
  XOR U8392 ( .A(n7321), .B(n7320), .Z(c[1260]) );
  NANDN U8393 ( .A(n7304), .B(n7303), .Z(n7308) );
  OR U8394 ( .A(n7306), .B(n7305), .Z(n7307) );
  AND U8395 ( .A(n7308), .B(n7307), .Z(n7326) );
  XOR U8396 ( .A(a[239]), .B(n2210), .Z(n7330) );
  AND U8397 ( .A(a[241]), .B(b[0]), .Z(n7310) );
  XNOR U8398 ( .A(n7310), .B(n2175), .Z(n7312) );
  NANDN U8399 ( .A(b[0]), .B(a[240]), .Z(n7311) );
  NAND U8400 ( .A(n7312), .B(n7311), .Z(n7335) );
  AND U8401 ( .A(a[237]), .B(b[3]), .Z(n7334) );
  XOR U8402 ( .A(n7335), .B(n7334), .Z(n7337) );
  XOR U8403 ( .A(n7336), .B(n7337), .Z(n7325) );
  NANDN U8404 ( .A(n7314), .B(n7313), .Z(n7318) );
  OR U8405 ( .A(n7316), .B(n7315), .Z(n7317) );
  AND U8406 ( .A(n7318), .B(n7317), .Z(n7324) );
  XOR U8407 ( .A(n7325), .B(n7324), .Z(n7327) );
  XOR U8408 ( .A(n7326), .B(n7327), .Z(n7340) );
  XNOR U8409 ( .A(n7340), .B(sreg[1261]), .Z(n7342) );
  NANDN U8410 ( .A(n7319), .B(sreg[1260]), .Z(n7323) );
  NAND U8411 ( .A(n7321), .B(n7320), .Z(n7322) );
  NAND U8412 ( .A(n7323), .B(n7322), .Z(n7341) );
  XOR U8413 ( .A(n7342), .B(n7341), .Z(c[1261]) );
  NANDN U8414 ( .A(n7325), .B(n7324), .Z(n7329) );
  OR U8415 ( .A(n7327), .B(n7326), .Z(n7328) );
  AND U8416 ( .A(n7329), .B(n7328), .Z(n7347) );
  XOR U8417 ( .A(a[240]), .B(n2210), .Z(n7351) );
  AND U8418 ( .A(a[242]), .B(b[0]), .Z(n7331) );
  XNOR U8419 ( .A(n7331), .B(n2175), .Z(n7333) );
  NANDN U8420 ( .A(b[0]), .B(a[241]), .Z(n7332) );
  NAND U8421 ( .A(n7333), .B(n7332), .Z(n7356) );
  AND U8422 ( .A(a[238]), .B(b[3]), .Z(n7355) );
  XOR U8423 ( .A(n7356), .B(n7355), .Z(n7358) );
  XOR U8424 ( .A(n7357), .B(n7358), .Z(n7346) );
  NANDN U8425 ( .A(n7335), .B(n7334), .Z(n7339) );
  OR U8426 ( .A(n7337), .B(n7336), .Z(n7338) );
  AND U8427 ( .A(n7339), .B(n7338), .Z(n7345) );
  XOR U8428 ( .A(n7346), .B(n7345), .Z(n7348) );
  XOR U8429 ( .A(n7347), .B(n7348), .Z(n7361) );
  XNOR U8430 ( .A(n7361), .B(sreg[1262]), .Z(n7363) );
  NANDN U8431 ( .A(n7340), .B(sreg[1261]), .Z(n7344) );
  NAND U8432 ( .A(n7342), .B(n7341), .Z(n7343) );
  NAND U8433 ( .A(n7344), .B(n7343), .Z(n7362) );
  XOR U8434 ( .A(n7363), .B(n7362), .Z(c[1262]) );
  NANDN U8435 ( .A(n7346), .B(n7345), .Z(n7350) );
  OR U8436 ( .A(n7348), .B(n7347), .Z(n7349) );
  AND U8437 ( .A(n7350), .B(n7349), .Z(n7368) );
  XOR U8438 ( .A(a[241]), .B(n2210), .Z(n7372) );
  AND U8439 ( .A(a[243]), .B(b[0]), .Z(n7352) );
  XNOR U8440 ( .A(n7352), .B(n2175), .Z(n7354) );
  NANDN U8441 ( .A(b[0]), .B(a[242]), .Z(n7353) );
  NAND U8442 ( .A(n7354), .B(n7353), .Z(n7377) );
  AND U8443 ( .A(a[239]), .B(b[3]), .Z(n7376) );
  XOR U8444 ( .A(n7377), .B(n7376), .Z(n7379) );
  XOR U8445 ( .A(n7378), .B(n7379), .Z(n7367) );
  NANDN U8446 ( .A(n7356), .B(n7355), .Z(n7360) );
  OR U8447 ( .A(n7358), .B(n7357), .Z(n7359) );
  AND U8448 ( .A(n7360), .B(n7359), .Z(n7366) );
  XOR U8449 ( .A(n7367), .B(n7366), .Z(n7369) );
  XOR U8450 ( .A(n7368), .B(n7369), .Z(n7382) );
  XNOR U8451 ( .A(n7382), .B(sreg[1263]), .Z(n7384) );
  NANDN U8452 ( .A(n7361), .B(sreg[1262]), .Z(n7365) );
  NAND U8453 ( .A(n7363), .B(n7362), .Z(n7364) );
  NAND U8454 ( .A(n7365), .B(n7364), .Z(n7383) );
  XOR U8455 ( .A(n7384), .B(n7383), .Z(c[1263]) );
  NANDN U8456 ( .A(n7367), .B(n7366), .Z(n7371) );
  OR U8457 ( .A(n7369), .B(n7368), .Z(n7370) );
  AND U8458 ( .A(n7371), .B(n7370), .Z(n7389) );
  XOR U8459 ( .A(a[242]), .B(n2210), .Z(n7393) );
  AND U8460 ( .A(a[240]), .B(b[3]), .Z(n7397) );
  AND U8461 ( .A(a[244]), .B(b[0]), .Z(n7373) );
  XNOR U8462 ( .A(n7373), .B(n2175), .Z(n7375) );
  NANDN U8463 ( .A(b[0]), .B(a[243]), .Z(n7374) );
  NAND U8464 ( .A(n7375), .B(n7374), .Z(n7398) );
  XOR U8465 ( .A(n7397), .B(n7398), .Z(n7400) );
  XOR U8466 ( .A(n7399), .B(n7400), .Z(n7388) );
  NANDN U8467 ( .A(n7377), .B(n7376), .Z(n7381) );
  OR U8468 ( .A(n7379), .B(n7378), .Z(n7380) );
  AND U8469 ( .A(n7381), .B(n7380), .Z(n7387) );
  XOR U8470 ( .A(n7388), .B(n7387), .Z(n7390) );
  XOR U8471 ( .A(n7389), .B(n7390), .Z(n7403) );
  XNOR U8472 ( .A(n7403), .B(sreg[1264]), .Z(n7405) );
  NANDN U8473 ( .A(n7382), .B(sreg[1263]), .Z(n7386) );
  NAND U8474 ( .A(n7384), .B(n7383), .Z(n7385) );
  NAND U8475 ( .A(n7386), .B(n7385), .Z(n7404) );
  XOR U8476 ( .A(n7405), .B(n7404), .Z(c[1264]) );
  NANDN U8477 ( .A(n7388), .B(n7387), .Z(n7392) );
  OR U8478 ( .A(n7390), .B(n7389), .Z(n7391) );
  AND U8479 ( .A(n7392), .B(n7391), .Z(n7410) );
  XOR U8480 ( .A(a[243]), .B(n2210), .Z(n7414) );
  AND U8481 ( .A(a[245]), .B(b[0]), .Z(n7394) );
  XNOR U8482 ( .A(n7394), .B(n2175), .Z(n7396) );
  NANDN U8483 ( .A(b[0]), .B(a[244]), .Z(n7395) );
  NAND U8484 ( .A(n7396), .B(n7395), .Z(n7419) );
  AND U8485 ( .A(a[241]), .B(b[3]), .Z(n7418) );
  XOR U8486 ( .A(n7419), .B(n7418), .Z(n7421) );
  XOR U8487 ( .A(n7420), .B(n7421), .Z(n7409) );
  NANDN U8488 ( .A(n7398), .B(n7397), .Z(n7402) );
  OR U8489 ( .A(n7400), .B(n7399), .Z(n7401) );
  AND U8490 ( .A(n7402), .B(n7401), .Z(n7408) );
  XOR U8491 ( .A(n7409), .B(n7408), .Z(n7411) );
  XOR U8492 ( .A(n7410), .B(n7411), .Z(n7424) );
  XNOR U8493 ( .A(n7424), .B(sreg[1265]), .Z(n7426) );
  NANDN U8494 ( .A(n7403), .B(sreg[1264]), .Z(n7407) );
  NAND U8495 ( .A(n7405), .B(n7404), .Z(n7406) );
  NAND U8496 ( .A(n7407), .B(n7406), .Z(n7425) );
  XOR U8497 ( .A(n7426), .B(n7425), .Z(c[1265]) );
  NANDN U8498 ( .A(n7409), .B(n7408), .Z(n7413) );
  OR U8499 ( .A(n7411), .B(n7410), .Z(n7412) );
  AND U8500 ( .A(n7413), .B(n7412), .Z(n7431) );
  XOR U8501 ( .A(a[244]), .B(n2211), .Z(n7435) );
  AND U8502 ( .A(a[242]), .B(b[3]), .Z(n7439) );
  AND U8503 ( .A(a[246]), .B(b[0]), .Z(n7415) );
  XNOR U8504 ( .A(n7415), .B(n2175), .Z(n7417) );
  NANDN U8505 ( .A(b[0]), .B(a[245]), .Z(n7416) );
  NAND U8506 ( .A(n7417), .B(n7416), .Z(n7440) );
  XOR U8507 ( .A(n7439), .B(n7440), .Z(n7442) );
  XOR U8508 ( .A(n7441), .B(n7442), .Z(n7430) );
  NANDN U8509 ( .A(n7419), .B(n7418), .Z(n7423) );
  OR U8510 ( .A(n7421), .B(n7420), .Z(n7422) );
  AND U8511 ( .A(n7423), .B(n7422), .Z(n7429) );
  XOR U8512 ( .A(n7430), .B(n7429), .Z(n7432) );
  XOR U8513 ( .A(n7431), .B(n7432), .Z(n7445) );
  XNOR U8514 ( .A(n7445), .B(sreg[1266]), .Z(n7447) );
  NANDN U8515 ( .A(n7424), .B(sreg[1265]), .Z(n7428) );
  NAND U8516 ( .A(n7426), .B(n7425), .Z(n7427) );
  NAND U8517 ( .A(n7428), .B(n7427), .Z(n7446) );
  XOR U8518 ( .A(n7447), .B(n7446), .Z(c[1266]) );
  NANDN U8519 ( .A(n7430), .B(n7429), .Z(n7434) );
  OR U8520 ( .A(n7432), .B(n7431), .Z(n7433) );
  AND U8521 ( .A(n7434), .B(n7433), .Z(n7452) );
  XOR U8522 ( .A(a[245]), .B(n2211), .Z(n7456) );
  AND U8523 ( .A(a[247]), .B(b[0]), .Z(n7436) );
  XNOR U8524 ( .A(n7436), .B(n2175), .Z(n7438) );
  NANDN U8525 ( .A(b[0]), .B(a[246]), .Z(n7437) );
  NAND U8526 ( .A(n7438), .B(n7437), .Z(n7461) );
  AND U8527 ( .A(a[243]), .B(b[3]), .Z(n7460) );
  XOR U8528 ( .A(n7461), .B(n7460), .Z(n7463) );
  XOR U8529 ( .A(n7462), .B(n7463), .Z(n7451) );
  NANDN U8530 ( .A(n7440), .B(n7439), .Z(n7444) );
  OR U8531 ( .A(n7442), .B(n7441), .Z(n7443) );
  AND U8532 ( .A(n7444), .B(n7443), .Z(n7450) );
  XOR U8533 ( .A(n7451), .B(n7450), .Z(n7453) );
  XOR U8534 ( .A(n7452), .B(n7453), .Z(n7466) );
  XNOR U8535 ( .A(n7466), .B(sreg[1267]), .Z(n7468) );
  NANDN U8536 ( .A(n7445), .B(sreg[1266]), .Z(n7449) );
  NAND U8537 ( .A(n7447), .B(n7446), .Z(n7448) );
  NAND U8538 ( .A(n7449), .B(n7448), .Z(n7467) );
  XOR U8539 ( .A(n7468), .B(n7467), .Z(c[1267]) );
  NANDN U8540 ( .A(n7451), .B(n7450), .Z(n7455) );
  OR U8541 ( .A(n7453), .B(n7452), .Z(n7454) );
  AND U8542 ( .A(n7455), .B(n7454), .Z(n7473) );
  XOR U8543 ( .A(a[246]), .B(n2211), .Z(n7477) );
  AND U8544 ( .A(a[248]), .B(b[0]), .Z(n7457) );
  XNOR U8545 ( .A(n7457), .B(n2175), .Z(n7459) );
  NANDN U8546 ( .A(b[0]), .B(a[247]), .Z(n7458) );
  NAND U8547 ( .A(n7459), .B(n7458), .Z(n7482) );
  AND U8548 ( .A(a[244]), .B(b[3]), .Z(n7481) );
  XOR U8549 ( .A(n7482), .B(n7481), .Z(n7484) );
  XOR U8550 ( .A(n7483), .B(n7484), .Z(n7472) );
  NANDN U8551 ( .A(n7461), .B(n7460), .Z(n7465) );
  OR U8552 ( .A(n7463), .B(n7462), .Z(n7464) );
  AND U8553 ( .A(n7465), .B(n7464), .Z(n7471) );
  XOR U8554 ( .A(n7472), .B(n7471), .Z(n7474) );
  XOR U8555 ( .A(n7473), .B(n7474), .Z(n7487) );
  XNOR U8556 ( .A(n7487), .B(sreg[1268]), .Z(n7489) );
  NANDN U8557 ( .A(n7466), .B(sreg[1267]), .Z(n7470) );
  NAND U8558 ( .A(n7468), .B(n7467), .Z(n7469) );
  NAND U8559 ( .A(n7470), .B(n7469), .Z(n7488) );
  XOR U8560 ( .A(n7489), .B(n7488), .Z(c[1268]) );
  NANDN U8561 ( .A(n7472), .B(n7471), .Z(n7476) );
  OR U8562 ( .A(n7474), .B(n7473), .Z(n7475) );
  AND U8563 ( .A(n7476), .B(n7475), .Z(n7494) );
  XOR U8564 ( .A(a[247]), .B(n2211), .Z(n7498) );
  AND U8565 ( .A(a[249]), .B(b[0]), .Z(n7478) );
  XNOR U8566 ( .A(n7478), .B(n2175), .Z(n7480) );
  NANDN U8567 ( .A(b[0]), .B(a[248]), .Z(n7479) );
  NAND U8568 ( .A(n7480), .B(n7479), .Z(n7503) );
  AND U8569 ( .A(a[245]), .B(b[3]), .Z(n7502) );
  XOR U8570 ( .A(n7503), .B(n7502), .Z(n7505) );
  XOR U8571 ( .A(n7504), .B(n7505), .Z(n7493) );
  NANDN U8572 ( .A(n7482), .B(n7481), .Z(n7486) );
  OR U8573 ( .A(n7484), .B(n7483), .Z(n7485) );
  AND U8574 ( .A(n7486), .B(n7485), .Z(n7492) );
  XOR U8575 ( .A(n7493), .B(n7492), .Z(n7495) );
  XOR U8576 ( .A(n7494), .B(n7495), .Z(n7508) );
  XNOR U8577 ( .A(n7508), .B(sreg[1269]), .Z(n7510) );
  NANDN U8578 ( .A(n7487), .B(sreg[1268]), .Z(n7491) );
  NAND U8579 ( .A(n7489), .B(n7488), .Z(n7490) );
  NAND U8580 ( .A(n7491), .B(n7490), .Z(n7509) );
  XOR U8581 ( .A(n7510), .B(n7509), .Z(c[1269]) );
  NANDN U8582 ( .A(n7493), .B(n7492), .Z(n7497) );
  OR U8583 ( .A(n7495), .B(n7494), .Z(n7496) );
  AND U8584 ( .A(n7497), .B(n7496), .Z(n7515) );
  XOR U8585 ( .A(a[248]), .B(n2211), .Z(n7519) );
  AND U8586 ( .A(a[246]), .B(b[3]), .Z(n7523) );
  AND U8587 ( .A(a[250]), .B(b[0]), .Z(n7499) );
  XNOR U8588 ( .A(n7499), .B(n2175), .Z(n7501) );
  NANDN U8589 ( .A(b[0]), .B(a[249]), .Z(n7500) );
  NAND U8590 ( .A(n7501), .B(n7500), .Z(n7524) );
  XOR U8591 ( .A(n7523), .B(n7524), .Z(n7526) );
  XOR U8592 ( .A(n7525), .B(n7526), .Z(n7514) );
  NANDN U8593 ( .A(n7503), .B(n7502), .Z(n7507) );
  OR U8594 ( .A(n7505), .B(n7504), .Z(n7506) );
  AND U8595 ( .A(n7507), .B(n7506), .Z(n7513) );
  XOR U8596 ( .A(n7514), .B(n7513), .Z(n7516) );
  XOR U8597 ( .A(n7515), .B(n7516), .Z(n7529) );
  XNOR U8598 ( .A(n7529), .B(sreg[1270]), .Z(n7531) );
  NANDN U8599 ( .A(n7508), .B(sreg[1269]), .Z(n7512) );
  NAND U8600 ( .A(n7510), .B(n7509), .Z(n7511) );
  NAND U8601 ( .A(n7512), .B(n7511), .Z(n7530) );
  XOR U8602 ( .A(n7531), .B(n7530), .Z(c[1270]) );
  NANDN U8603 ( .A(n7514), .B(n7513), .Z(n7518) );
  OR U8604 ( .A(n7516), .B(n7515), .Z(n7517) );
  AND U8605 ( .A(n7518), .B(n7517), .Z(n7537) );
  XOR U8606 ( .A(a[249]), .B(n2211), .Z(n7538) );
  AND U8607 ( .A(b[0]), .B(a[251]), .Z(n7520) );
  XOR U8608 ( .A(b[1]), .B(n7520), .Z(n7522) );
  NANDN U8609 ( .A(b[0]), .B(a[250]), .Z(n7521) );
  AND U8610 ( .A(n7522), .B(n7521), .Z(n7542) );
  AND U8611 ( .A(a[247]), .B(b[3]), .Z(n7543) );
  XOR U8612 ( .A(n7542), .B(n7543), .Z(n7544) );
  XNOR U8613 ( .A(n7545), .B(n7544), .Z(n7534) );
  NANDN U8614 ( .A(n7524), .B(n7523), .Z(n7528) );
  OR U8615 ( .A(n7526), .B(n7525), .Z(n7527) );
  AND U8616 ( .A(n7528), .B(n7527), .Z(n7535) );
  XNOR U8617 ( .A(n7534), .B(n7535), .Z(n7536) );
  XNOR U8618 ( .A(n7537), .B(n7536), .Z(n7548) );
  XNOR U8619 ( .A(n7548), .B(sreg[1271]), .Z(n7550) );
  NANDN U8620 ( .A(n7529), .B(sreg[1270]), .Z(n7533) );
  NAND U8621 ( .A(n7531), .B(n7530), .Z(n7532) );
  NAND U8622 ( .A(n7533), .B(n7532), .Z(n7549) );
  XOR U8623 ( .A(n7550), .B(n7549), .Z(c[1271]) );
  XOR U8624 ( .A(a[250]), .B(n2211), .Z(n7557) );
  AND U8625 ( .A(a[252]), .B(b[0]), .Z(n7539) );
  XNOR U8626 ( .A(n7539), .B(n2175), .Z(n7541) );
  NANDN U8627 ( .A(b[0]), .B(a[251]), .Z(n7540) );
  NAND U8628 ( .A(n7541), .B(n7540), .Z(n7562) );
  AND U8629 ( .A(a[248]), .B(b[3]), .Z(n7561) );
  XOR U8630 ( .A(n7562), .B(n7561), .Z(n7564) );
  XOR U8631 ( .A(n7563), .B(n7564), .Z(n7552) );
  NAND U8632 ( .A(n7543), .B(n7542), .Z(n7547) );
  NANDN U8633 ( .A(n7545), .B(n7544), .Z(n7546) );
  AND U8634 ( .A(n7547), .B(n7546), .Z(n7551) );
  XOR U8635 ( .A(n7552), .B(n7551), .Z(n7554) );
  XOR U8636 ( .A(n7553), .B(n7554), .Z(n7567) );
  XNOR U8637 ( .A(n7567), .B(sreg[1272]), .Z(n7569) );
  XOR U8638 ( .A(n7569), .B(n7568), .Z(c[1272]) );
  NANDN U8639 ( .A(n7552), .B(n7551), .Z(n7556) );
  OR U8640 ( .A(n7554), .B(n7553), .Z(n7555) );
  AND U8641 ( .A(n7556), .B(n7555), .Z(n7574) );
  XOR U8642 ( .A(a[251]), .B(n2212), .Z(n7578) );
  AND U8643 ( .A(a[253]), .B(b[0]), .Z(n7558) );
  XNOR U8644 ( .A(n7558), .B(n2175), .Z(n7560) );
  NANDN U8645 ( .A(b[0]), .B(a[252]), .Z(n7559) );
  NAND U8646 ( .A(n7560), .B(n7559), .Z(n7583) );
  AND U8647 ( .A(a[249]), .B(b[3]), .Z(n7582) );
  XOR U8648 ( .A(n7583), .B(n7582), .Z(n7585) );
  XOR U8649 ( .A(n7584), .B(n7585), .Z(n7573) );
  NANDN U8650 ( .A(n7562), .B(n7561), .Z(n7566) );
  OR U8651 ( .A(n7564), .B(n7563), .Z(n7565) );
  AND U8652 ( .A(n7566), .B(n7565), .Z(n7572) );
  XOR U8653 ( .A(n7573), .B(n7572), .Z(n7575) );
  XOR U8654 ( .A(n7574), .B(n7575), .Z(n7588) );
  XNOR U8655 ( .A(n7588), .B(sreg[1273]), .Z(n7590) );
  NANDN U8656 ( .A(n7567), .B(sreg[1272]), .Z(n7571) );
  NAND U8657 ( .A(n7569), .B(n7568), .Z(n7570) );
  NAND U8658 ( .A(n7571), .B(n7570), .Z(n7589) );
  XOR U8659 ( .A(n7590), .B(n7589), .Z(c[1273]) );
  NANDN U8660 ( .A(n7573), .B(n7572), .Z(n7577) );
  OR U8661 ( .A(n7575), .B(n7574), .Z(n7576) );
  AND U8662 ( .A(n7577), .B(n7576), .Z(n7595) );
  XOR U8663 ( .A(a[252]), .B(n2212), .Z(n7599) );
  AND U8664 ( .A(a[254]), .B(b[0]), .Z(n7579) );
  XNOR U8665 ( .A(n7579), .B(n2175), .Z(n7581) );
  NANDN U8666 ( .A(b[0]), .B(a[253]), .Z(n7580) );
  NAND U8667 ( .A(n7581), .B(n7580), .Z(n7604) );
  AND U8668 ( .A(a[250]), .B(b[3]), .Z(n7603) );
  XOR U8669 ( .A(n7604), .B(n7603), .Z(n7606) );
  XOR U8670 ( .A(n7605), .B(n7606), .Z(n7594) );
  NANDN U8671 ( .A(n7583), .B(n7582), .Z(n7587) );
  OR U8672 ( .A(n7585), .B(n7584), .Z(n7586) );
  AND U8673 ( .A(n7587), .B(n7586), .Z(n7593) );
  XOR U8674 ( .A(n7594), .B(n7593), .Z(n7596) );
  XOR U8675 ( .A(n7595), .B(n7596), .Z(n7609) );
  XNOR U8676 ( .A(n7609), .B(sreg[1274]), .Z(n7611) );
  NANDN U8677 ( .A(n7588), .B(sreg[1273]), .Z(n7592) );
  NAND U8678 ( .A(n7590), .B(n7589), .Z(n7591) );
  NAND U8679 ( .A(n7592), .B(n7591), .Z(n7610) );
  XOR U8680 ( .A(n7611), .B(n7610), .Z(c[1274]) );
  NANDN U8681 ( .A(n7594), .B(n7593), .Z(n7598) );
  OR U8682 ( .A(n7596), .B(n7595), .Z(n7597) );
  AND U8683 ( .A(n7598), .B(n7597), .Z(n7616) );
  XOR U8684 ( .A(a[253]), .B(n2212), .Z(n7620) );
  AND U8685 ( .A(a[255]), .B(b[0]), .Z(n7600) );
  XNOR U8686 ( .A(n7600), .B(n2175), .Z(n7602) );
  NANDN U8687 ( .A(b[0]), .B(a[254]), .Z(n7601) );
  NAND U8688 ( .A(n7602), .B(n7601), .Z(n7625) );
  AND U8689 ( .A(a[251]), .B(b[3]), .Z(n7624) );
  XOR U8690 ( .A(n7625), .B(n7624), .Z(n7627) );
  XOR U8691 ( .A(n7626), .B(n7627), .Z(n7615) );
  NANDN U8692 ( .A(n7604), .B(n7603), .Z(n7608) );
  OR U8693 ( .A(n7606), .B(n7605), .Z(n7607) );
  AND U8694 ( .A(n7608), .B(n7607), .Z(n7614) );
  XOR U8695 ( .A(n7615), .B(n7614), .Z(n7617) );
  XOR U8696 ( .A(n7616), .B(n7617), .Z(n7630) );
  XNOR U8697 ( .A(n7630), .B(sreg[1275]), .Z(n7632) );
  NANDN U8698 ( .A(n7609), .B(sreg[1274]), .Z(n7613) );
  NAND U8699 ( .A(n7611), .B(n7610), .Z(n7612) );
  NAND U8700 ( .A(n7613), .B(n7612), .Z(n7631) );
  XOR U8701 ( .A(n7632), .B(n7631), .Z(c[1275]) );
  NANDN U8702 ( .A(n7615), .B(n7614), .Z(n7619) );
  OR U8703 ( .A(n7617), .B(n7616), .Z(n7618) );
  AND U8704 ( .A(n7619), .B(n7618), .Z(n7637) );
  XOR U8705 ( .A(a[254]), .B(n2212), .Z(n7641) );
  AND U8706 ( .A(a[252]), .B(b[3]), .Z(n7645) );
  AND U8707 ( .A(a[256]), .B(b[0]), .Z(n7621) );
  XNOR U8708 ( .A(n7621), .B(n2175), .Z(n7623) );
  NANDN U8709 ( .A(b[0]), .B(a[255]), .Z(n7622) );
  NAND U8710 ( .A(n7623), .B(n7622), .Z(n7646) );
  XOR U8711 ( .A(n7645), .B(n7646), .Z(n7648) );
  XOR U8712 ( .A(n7647), .B(n7648), .Z(n7636) );
  NANDN U8713 ( .A(n7625), .B(n7624), .Z(n7629) );
  OR U8714 ( .A(n7627), .B(n7626), .Z(n7628) );
  AND U8715 ( .A(n7629), .B(n7628), .Z(n7635) );
  XOR U8716 ( .A(n7636), .B(n7635), .Z(n7638) );
  XOR U8717 ( .A(n7637), .B(n7638), .Z(n7651) );
  XNOR U8718 ( .A(n7651), .B(sreg[1276]), .Z(n7653) );
  NANDN U8719 ( .A(n7630), .B(sreg[1275]), .Z(n7634) );
  NAND U8720 ( .A(n7632), .B(n7631), .Z(n7633) );
  NAND U8721 ( .A(n7634), .B(n7633), .Z(n7652) );
  XOR U8722 ( .A(n7653), .B(n7652), .Z(c[1276]) );
  NANDN U8723 ( .A(n7636), .B(n7635), .Z(n7640) );
  OR U8724 ( .A(n7638), .B(n7637), .Z(n7639) );
  AND U8725 ( .A(n7640), .B(n7639), .Z(n7658) );
  XOR U8726 ( .A(a[255]), .B(n2212), .Z(n7662) );
  AND U8727 ( .A(a[257]), .B(b[0]), .Z(n7642) );
  XNOR U8728 ( .A(n7642), .B(n2175), .Z(n7644) );
  NANDN U8729 ( .A(b[0]), .B(a[256]), .Z(n7643) );
  NAND U8730 ( .A(n7644), .B(n7643), .Z(n7667) );
  AND U8731 ( .A(a[253]), .B(b[3]), .Z(n7666) );
  XOR U8732 ( .A(n7667), .B(n7666), .Z(n7669) );
  XOR U8733 ( .A(n7668), .B(n7669), .Z(n7657) );
  NANDN U8734 ( .A(n7646), .B(n7645), .Z(n7650) );
  OR U8735 ( .A(n7648), .B(n7647), .Z(n7649) );
  AND U8736 ( .A(n7650), .B(n7649), .Z(n7656) );
  XOR U8737 ( .A(n7657), .B(n7656), .Z(n7659) );
  XOR U8738 ( .A(n7658), .B(n7659), .Z(n7672) );
  XNOR U8739 ( .A(n7672), .B(sreg[1277]), .Z(n7674) );
  NANDN U8740 ( .A(n7651), .B(sreg[1276]), .Z(n7655) );
  NAND U8741 ( .A(n7653), .B(n7652), .Z(n7654) );
  NAND U8742 ( .A(n7655), .B(n7654), .Z(n7673) );
  XOR U8743 ( .A(n7674), .B(n7673), .Z(c[1277]) );
  NANDN U8744 ( .A(n7657), .B(n7656), .Z(n7661) );
  OR U8745 ( .A(n7659), .B(n7658), .Z(n7660) );
  AND U8746 ( .A(n7661), .B(n7660), .Z(n7679) );
  XOR U8747 ( .A(a[256]), .B(n2212), .Z(n7683) );
  AND U8748 ( .A(a[258]), .B(b[0]), .Z(n7663) );
  XNOR U8749 ( .A(n7663), .B(n2175), .Z(n7665) );
  NANDN U8750 ( .A(b[0]), .B(a[257]), .Z(n7664) );
  NAND U8751 ( .A(n7665), .B(n7664), .Z(n7688) );
  AND U8752 ( .A(a[254]), .B(b[3]), .Z(n7687) );
  XOR U8753 ( .A(n7688), .B(n7687), .Z(n7690) );
  XOR U8754 ( .A(n7689), .B(n7690), .Z(n7678) );
  NANDN U8755 ( .A(n7667), .B(n7666), .Z(n7671) );
  OR U8756 ( .A(n7669), .B(n7668), .Z(n7670) );
  AND U8757 ( .A(n7671), .B(n7670), .Z(n7677) );
  XOR U8758 ( .A(n7678), .B(n7677), .Z(n7680) );
  XOR U8759 ( .A(n7679), .B(n7680), .Z(n7693) );
  XNOR U8760 ( .A(n7693), .B(sreg[1278]), .Z(n7695) );
  NANDN U8761 ( .A(n7672), .B(sreg[1277]), .Z(n7676) );
  NAND U8762 ( .A(n7674), .B(n7673), .Z(n7675) );
  NAND U8763 ( .A(n7676), .B(n7675), .Z(n7694) );
  XOR U8764 ( .A(n7695), .B(n7694), .Z(c[1278]) );
  NANDN U8765 ( .A(n7678), .B(n7677), .Z(n7682) );
  OR U8766 ( .A(n7680), .B(n7679), .Z(n7681) );
  AND U8767 ( .A(n7682), .B(n7681), .Z(n7700) );
  XOR U8768 ( .A(a[257]), .B(n2212), .Z(n7704) );
  AND U8769 ( .A(a[255]), .B(b[3]), .Z(n7708) );
  AND U8770 ( .A(a[259]), .B(b[0]), .Z(n7684) );
  XNOR U8771 ( .A(n7684), .B(n2175), .Z(n7686) );
  NANDN U8772 ( .A(b[0]), .B(a[258]), .Z(n7685) );
  NAND U8773 ( .A(n7686), .B(n7685), .Z(n7709) );
  XOR U8774 ( .A(n7708), .B(n7709), .Z(n7711) );
  XOR U8775 ( .A(n7710), .B(n7711), .Z(n7699) );
  NANDN U8776 ( .A(n7688), .B(n7687), .Z(n7692) );
  OR U8777 ( .A(n7690), .B(n7689), .Z(n7691) );
  AND U8778 ( .A(n7692), .B(n7691), .Z(n7698) );
  XOR U8779 ( .A(n7699), .B(n7698), .Z(n7701) );
  XOR U8780 ( .A(n7700), .B(n7701), .Z(n7714) );
  XNOR U8781 ( .A(n7714), .B(sreg[1279]), .Z(n7716) );
  NANDN U8782 ( .A(n7693), .B(sreg[1278]), .Z(n7697) );
  NAND U8783 ( .A(n7695), .B(n7694), .Z(n7696) );
  NAND U8784 ( .A(n7697), .B(n7696), .Z(n7715) );
  XOR U8785 ( .A(n7716), .B(n7715), .Z(c[1279]) );
  NANDN U8786 ( .A(n7699), .B(n7698), .Z(n7703) );
  OR U8787 ( .A(n7701), .B(n7700), .Z(n7702) );
  AND U8788 ( .A(n7703), .B(n7702), .Z(n7721) );
  XOR U8789 ( .A(a[258]), .B(n2213), .Z(n7725) );
  AND U8790 ( .A(a[260]), .B(b[0]), .Z(n7705) );
  XNOR U8791 ( .A(n7705), .B(n2175), .Z(n7707) );
  NANDN U8792 ( .A(b[0]), .B(a[259]), .Z(n7706) );
  NAND U8793 ( .A(n7707), .B(n7706), .Z(n7730) );
  AND U8794 ( .A(a[256]), .B(b[3]), .Z(n7729) );
  XOR U8795 ( .A(n7730), .B(n7729), .Z(n7732) );
  XOR U8796 ( .A(n7731), .B(n7732), .Z(n7720) );
  NANDN U8797 ( .A(n7709), .B(n7708), .Z(n7713) );
  OR U8798 ( .A(n7711), .B(n7710), .Z(n7712) );
  AND U8799 ( .A(n7713), .B(n7712), .Z(n7719) );
  XOR U8800 ( .A(n7720), .B(n7719), .Z(n7722) );
  XOR U8801 ( .A(n7721), .B(n7722), .Z(n7735) );
  XNOR U8802 ( .A(n7735), .B(sreg[1280]), .Z(n7737) );
  NANDN U8803 ( .A(n7714), .B(sreg[1279]), .Z(n7718) );
  NAND U8804 ( .A(n7716), .B(n7715), .Z(n7717) );
  NAND U8805 ( .A(n7718), .B(n7717), .Z(n7736) );
  XOR U8806 ( .A(n7737), .B(n7736), .Z(c[1280]) );
  NANDN U8807 ( .A(n7720), .B(n7719), .Z(n7724) );
  OR U8808 ( .A(n7722), .B(n7721), .Z(n7723) );
  AND U8809 ( .A(n7724), .B(n7723), .Z(n7742) );
  XOR U8810 ( .A(a[259]), .B(n2213), .Z(n7746) );
  AND U8811 ( .A(a[261]), .B(b[0]), .Z(n7726) );
  XNOR U8812 ( .A(n7726), .B(n2175), .Z(n7728) );
  NANDN U8813 ( .A(b[0]), .B(a[260]), .Z(n7727) );
  NAND U8814 ( .A(n7728), .B(n7727), .Z(n7751) );
  AND U8815 ( .A(a[257]), .B(b[3]), .Z(n7750) );
  XOR U8816 ( .A(n7751), .B(n7750), .Z(n7753) );
  XOR U8817 ( .A(n7752), .B(n7753), .Z(n7741) );
  NANDN U8818 ( .A(n7730), .B(n7729), .Z(n7734) );
  OR U8819 ( .A(n7732), .B(n7731), .Z(n7733) );
  AND U8820 ( .A(n7734), .B(n7733), .Z(n7740) );
  XOR U8821 ( .A(n7741), .B(n7740), .Z(n7743) );
  XOR U8822 ( .A(n7742), .B(n7743), .Z(n7756) );
  XNOR U8823 ( .A(n7756), .B(sreg[1281]), .Z(n7758) );
  NANDN U8824 ( .A(n7735), .B(sreg[1280]), .Z(n7739) );
  NAND U8825 ( .A(n7737), .B(n7736), .Z(n7738) );
  NAND U8826 ( .A(n7739), .B(n7738), .Z(n7757) );
  XOR U8827 ( .A(n7758), .B(n7757), .Z(c[1281]) );
  NANDN U8828 ( .A(n7741), .B(n7740), .Z(n7745) );
  OR U8829 ( .A(n7743), .B(n7742), .Z(n7744) );
  AND U8830 ( .A(n7745), .B(n7744), .Z(n7763) );
  XOR U8831 ( .A(a[260]), .B(n2213), .Z(n7767) );
  AND U8832 ( .A(a[258]), .B(b[3]), .Z(n7771) );
  AND U8833 ( .A(a[262]), .B(b[0]), .Z(n7747) );
  XNOR U8834 ( .A(n7747), .B(n2175), .Z(n7749) );
  NANDN U8835 ( .A(b[0]), .B(a[261]), .Z(n7748) );
  NAND U8836 ( .A(n7749), .B(n7748), .Z(n7772) );
  XOR U8837 ( .A(n7771), .B(n7772), .Z(n7774) );
  XOR U8838 ( .A(n7773), .B(n7774), .Z(n7762) );
  NANDN U8839 ( .A(n7751), .B(n7750), .Z(n7755) );
  OR U8840 ( .A(n7753), .B(n7752), .Z(n7754) );
  AND U8841 ( .A(n7755), .B(n7754), .Z(n7761) );
  XOR U8842 ( .A(n7762), .B(n7761), .Z(n7764) );
  XOR U8843 ( .A(n7763), .B(n7764), .Z(n7777) );
  XNOR U8844 ( .A(n7777), .B(sreg[1282]), .Z(n7779) );
  NANDN U8845 ( .A(n7756), .B(sreg[1281]), .Z(n7760) );
  NAND U8846 ( .A(n7758), .B(n7757), .Z(n7759) );
  NAND U8847 ( .A(n7760), .B(n7759), .Z(n7778) );
  XOR U8848 ( .A(n7779), .B(n7778), .Z(c[1282]) );
  NANDN U8849 ( .A(n7762), .B(n7761), .Z(n7766) );
  OR U8850 ( .A(n7764), .B(n7763), .Z(n7765) );
  AND U8851 ( .A(n7766), .B(n7765), .Z(n7784) );
  XOR U8852 ( .A(a[261]), .B(n2213), .Z(n7788) );
  AND U8853 ( .A(a[263]), .B(b[0]), .Z(n7768) );
  XNOR U8854 ( .A(n7768), .B(n2175), .Z(n7770) );
  NANDN U8855 ( .A(b[0]), .B(a[262]), .Z(n7769) );
  NAND U8856 ( .A(n7770), .B(n7769), .Z(n7793) );
  AND U8857 ( .A(a[259]), .B(b[3]), .Z(n7792) );
  XOR U8858 ( .A(n7793), .B(n7792), .Z(n7795) );
  XOR U8859 ( .A(n7794), .B(n7795), .Z(n7783) );
  NANDN U8860 ( .A(n7772), .B(n7771), .Z(n7776) );
  OR U8861 ( .A(n7774), .B(n7773), .Z(n7775) );
  AND U8862 ( .A(n7776), .B(n7775), .Z(n7782) );
  XOR U8863 ( .A(n7783), .B(n7782), .Z(n7785) );
  XOR U8864 ( .A(n7784), .B(n7785), .Z(n7798) );
  XNOR U8865 ( .A(n7798), .B(sreg[1283]), .Z(n7800) );
  NANDN U8866 ( .A(n7777), .B(sreg[1282]), .Z(n7781) );
  NAND U8867 ( .A(n7779), .B(n7778), .Z(n7780) );
  NAND U8868 ( .A(n7781), .B(n7780), .Z(n7799) );
  XOR U8869 ( .A(n7800), .B(n7799), .Z(c[1283]) );
  NANDN U8870 ( .A(n7783), .B(n7782), .Z(n7787) );
  OR U8871 ( .A(n7785), .B(n7784), .Z(n7786) );
  AND U8872 ( .A(n7787), .B(n7786), .Z(n7806) );
  XOR U8873 ( .A(a[262]), .B(n2213), .Z(n7807) );
  AND U8874 ( .A(b[0]), .B(a[264]), .Z(n7789) );
  XOR U8875 ( .A(b[1]), .B(n7789), .Z(n7791) );
  NANDN U8876 ( .A(b[0]), .B(a[263]), .Z(n7790) );
  AND U8877 ( .A(n7791), .B(n7790), .Z(n7811) );
  AND U8878 ( .A(a[260]), .B(b[3]), .Z(n7812) );
  XOR U8879 ( .A(n7811), .B(n7812), .Z(n7813) );
  XNOR U8880 ( .A(n7814), .B(n7813), .Z(n7803) );
  NANDN U8881 ( .A(n7793), .B(n7792), .Z(n7797) );
  OR U8882 ( .A(n7795), .B(n7794), .Z(n7796) );
  AND U8883 ( .A(n7797), .B(n7796), .Z(n7804) );
  XNOR U8884 ( .A(n7803), .B(n7804), .Z(n7805) );
  XNOR U8885 ( .A(n7806), .B(n7805), .Z(n7817) );
  XNOR U8886 ( .A(n7817), .B(sreg[1284]), .Z(n7819) );
  NANDN U8887 ( .A(n7798), .B(sreg[1283]), .Z(n7802) );
  NAND U8888 ( .A(n7800), .B(n7799), .Z(n7801) );
  NAND U8889 ( .A(n7802), .B(n7801), .Z(n7818) );
  XOR U8890 ( .A(n7819), .B(n7818), .Z(c[1284]) );
  XOR U8891 ( .A(a[263]), .B(n2213), .Z(n7826) );
  AND U8892 ( .A(a[265]), .B(b[0]), .Z(n7808) );
  XNOR U8893 ( .A(n7808), .B(n2175), .Z(n7810) );
  NANDN U8894 ( .A(b[0]), .B(a[264]), .Z(n7809) );
  NAND U8895 ( .A(n7810), .B(n7809), .Z(n7831) );
  AND U8896 ( .A(a[261]), .B(b[3]), .Z(n7830) );
  XOR U8897 ( .A(n7831), .B(n7830), .Z(n7833) );
  XOR U8898 ( .A(n7832), .B(n7833), .Z(n7821) );
  NAND U8899 ( .A(n7812), .B(n7811), .Z(n7816) );
  NANDN U8900 ( .A(n7814), .B(n7813), .Z(n7815) );
  AND U8901 ( .A(n7816), .B(n7815), .Z(n7820) );
  XOR U8902 ( .A(n7821), .B(n7820), .Z(n7823) );
  XOR U8903 ( .A(n7822), .B(n7823), .Z(n7836) );
  XNOR U8904 ( .A(n7836), .B(sreg[1285]), .Z(n7838) );
  XOR U8905 ( .A(n7838), .B(n7837), .Z(c[1285]) );
  NANDN U8906 ( .A(n7821), .B(n7820), .Z(n7825) );
  OR U8907 ( .A(n7823), .B(n7822), .Z(n7824) );
  AND U8908 ( .A(n7825), .B(n7824), .Z(n7843) );
  XOR U8909 ( .A(a[264]), .B(n2213), .Z(n7847) );
  AND U8910 ( .A(a[266]), .B(b[0]), .Z(n7827) );
  XNOR U8911 ( .A(n7827), .B(n2175), .Z(n7829) );
  NANDN U8912 ( .A(b[0]), .B(a[265]), .Z(n7828) );
  NAND U8913 ( .A(n7829), .B(n7828), .Z(n7852) );
  AND U8914 ( .A(a[262]), .B(b[3]), .Z(n7851) );
  XOR U8915 ( .A(n7852), .B(n7851), .Z(n7854) );
  XOR U8916 ( .A(n7853), .B(n7854), .Z(n7842) );
  NANDN U8917 ( .A(n7831), .B(n7830), .Z(n7835) );
  OR U8918 ( .A(n7833), .B(n7832), .Z(n7834) );
  AND U8919 ( .A(n7835), .B(n7834), .Z(n7841) );
  XOR U8920 ( .A(n7842), .B(n7841), .Z(n7844) );
  XOR U8921 ( .A(n7843), .B(n7844), .Z(n7857) );
  XNOR U8922 ( .A(n7857), .B(sreg[1286]), .Z(n7859) );
  NANDN U8923 ( .A(n7836), .B(sreg[1285]), .Z(n7840) );
  NAND U8924 ( .A(n7838), .B(n7837), .Z(n7839) );
  NAND U8925 ( .A(n7840), .B(n7839), .Z(n7858) );
  XOR U8926 ( .A(n7859), .B(n7858), .Z(c[1286]) );
  NANDN U8927 ( .A(n7842), .B(n7841), .Z(n7846) );
  OR U8928 ( .A(n7844), .B(n7843), .Z(n7845) );
  AND U8929 ( .A(n7846), .B(n7845), .Z(n7864) );
  XOR U8930 ( .A(a[265]), .B(n2214), .Z(n7868) );
  AND U8931 ( .A(a[263]), .B(b[3]), .Z(n7872) );
  AND U8932 ( .A(a[267]), .B(b[0]), .Z(n7848) );
  XNOR U8933 ( .A(n7848), .B(n2175), .Z(n7850) );
  NANDN U8934 ( .A(b[0]), .B(a[266]), .Z(n7849) );
  NAND U8935 ( .A(n7850), .B(n7849), .Z(n7873) );
  XOR U8936 ( .A(n7872), .B(n7873), .Z(n7875) );
  XOR U8937 ( .A(n7874), .B(n7875), .Z(n7863) );
  NANDN U8938 ( .A(n7852), .B(n7851), .Z(n7856) );
  OR U8939 ( .A(n7854), .B(n7853), .Z(n7855) );
  AND U8940 ( .A(n7856), .B(n7855), .Z(n7862) );
  XOR U8941 ( .A(n7863), .B(n7862), .Z(n7865) );
  XOR U8942 ( .A(n7864), .B(n7865), .Z(n7878) );
  XNOR U8943 ( .A(n7878), .B(sreg[1287]), .Z(n7880) );
  NANDN U8944 ( .A(n7857), .B(sreg[1286]), .Z(n7861) );
  NAND U8945 ( .A(n7859), .B(n7858), .Z(n7860) );
  NAND U8946 ( .A(n7861), .B(n7860), .Z(n7879) );
  XOR U8947 ( .A(n7880), .B(n7879), .Z(c[1287]) );
  NANDN U8948 ( .A(n7863), .B(n7862), .Z(n7867) );
  OR U8949 ( .A(n7865), .B(n7864), .Z(n7866) );
  AND U8950 ( .A(n7867), .B(n7866), .Z(n7885) );
  XOR U8951 ( .A(a[266]), .B(n2214), .Z(n7889) );
  AND U8952 ( .A(a[268]), .B(b[0]), .Z(n7869) );
  XNOR U8953 ( .A(n7869), .B(n2175), .Z(n7871) );
  NANDN U8954 ( .A(b[0]), .B(a[267]), .Z(n7870) );
  NAND U8955 ( .A(n7871), .B(n7870), .Z(n7894) );
  AND U8956 ( .A(a[264]), .B(b[3]), .Z(n7893) );
  XOR U8957 ( .A(n7894), .B(n7893), .Z(n7896) );
  XOR U8958 ( .A(n7895), .B(n7896), .Z(n7884) );
  NANDN U8959 ( .A(n7873), .B(n7872), .Z(n7877) );
  OR U8960 ( .A(n7875), .B(n7874), .Z(n7876) );
  AND U8961 ( .A(n7877), .B(n7876), .Z(n7883) );
  XOR U8962 ( .A(n7884), .B(n7883), .Z(n7886) );
  XOR U8963 ( .A(n7885), .B(n7886), .Z(n7899) );
  XNOR U8964 ( .A(n7899), .B(sreg[1288]), .Z(n7901) );
  NANDN U8965 ( .A(n7878), .B(sreg[1287]), .Z(n7882) );
  NAND U8966 ( .A(n7880), .B(n7879), .Z(n7881) );
  NAND U8967 ( .A(n7882), .B(n7881), .Z(n7900) );
  XOR U8968 ( .A(n7901), .B(n7900), .Z(c[1288]) );
  NANDN U8969 ( .A(n7884), .B(n7883), .Z(n7888) );
  OR U8970 ( .A(n7886), .B(n7885), .Z(n7887) );
  AND U8971 ( .A(n7888), .B(n7887), .Z(n7906) );
  XOR U8972 ( .A(a[267]), .B(n2214), .Z(n7910) );
  AND U8973 ( .A(a[269]), .B(b[0]), .Z(n7890) );
  XNOR U8974 ( .A(n7890), .B(n2175), .Z(n7892) );
  NANDN U8975 ( .A(b[0]), .B(a[268]), .Z(n7891) );
  NAND U8976 ( .A(n7892), .B(n7891), .Z(n7915) );
  AND U8977 ( .A(a[265]), .B(b[3]), .Z(n7914) );
  XOR U8978 ( .A(n7915), .B(n7914), .Z(n7917) );
  XOR U8979 ( .A(n7916), .B(n7917), .Z(n7905) );
  NANDN U8980 ( .A(n7894), .B(n7893), .Z(n7898) );
  OR U8981 ( .A(n7896), .B(n7895), .Z(n7897) );
  AND U8982 ( .A(n7898), .B(n7897), .Z(n7904) );
  XOR U8983 ( .A(n7905), .B(n7904), .Z(n7907) );
  XOR U8984 ( .A(n7906), .B(n7907), .Z(n7920) );
  XNOR U8985 ( .A(n7920), .B(sreg[1289]), .Z(n7922) );
  NANDN U8986 ( .A(n7899), .B(sreg[1288]), .Z(n7903) );
  NAND U8987 ( .A(n7901), .B(n7900), .Z(n7902) );
  NAND U8988 ( .A(n7903), .B(n7902), .Z(n7921) );
  XOR U8989 ( .A(n7922), .B(n7921), .Z(c[1289]) );
  NANDN U8990 ( .A(n7905), .B(n7904), .Z(n7909) );
  OR U8991 ( .A(n7907), .B(n7906), .Z(n7908) );
  AND U8992 ( .A(n7909), .B(n7908), .Z(n7928) );
  XOR U8993 ( .A(a[268]), .B(n2214), .Z(n7929) );
  AND U8994 ( .A(b[0]), .B(a[270]), .Z(n7911) );
  XOR U8995 ( .A(b[1]), .B(n7911), .Z(n7913) );
  NANDN U8996 ( .A(b[0]), .B(a[269]), .Z(n7912) );
  AND U8997 ( .A(n7913), .B(n7912), .Z(n7933) );
  AND U8998 ( .A(a[266]), .B(b[3]), .Z(n7934) );
  XOR U8999 ( .A(n7933), .B(n7934), .Z(n7935) );
  XNOR U9000 ( .A(n7936), .B(n7935), .Z(n7925) );
  NANDN U9001 ( .A(n7915), .B(n7914), .Z(n7919) );
  OR U9002 ( .A(n7917), .B(n7916), .Z(n7918) );
  AND U9003 ( .A(n7919), .B(n7918), .Z(n7926) );
  XNOR U9004 ( .A(n7925), .B(n7926), .Z(n7927) );
  XNOR U9005 ( .A(n7928), .B(n7927), .Z(n7939) );
  XNOR U9006 ( .A(n7939), .B(sreg[1290]), .Z(n7941) );
  NANDN U9007 ( .A(n7920), .B(sreg[1289]), .Z(n7924) );
  NAND U9008 ( .A(n7922), .B(n7921), .Z(n7923) );
  NAND U9009 ( .A(n7924), .B(n7923), .Z(n7940) );
  XOR U9010 ( .A(n7941), .B(n7940), .Z(c[1290]) );
  XOR U9011 ( .A(a[269]), .B(n2214), .Z(n7948) );
  AND U9012 ( .A(a[271]), .B(b[0]), .Z(n7930) );
  XNOR U9013 ( .A(n7930), .B(n2175), .Z(n7932) );
  NANDN U9014 ( .A(b[0]), .B(a[270]), .Z(n7931) );
  NAND U9015 ( .A(n7932), .B(n7931), .Z(n7953) );
  AND U9016 ( .A(a[267]), .B(b[3]), .Z(n7952) );
  XOR U9017 ( .A(n7953), .B(n7952), .Z(n7955) );
  XOR U9018 ( .A(n7954), .B(n7955), .Z(n7943) );
  NAND U9019 ( .A(n7934), .B(n7933), .Z(n7938) );
  NANDN U9020 ( .A(n7936), .B(n7935), .Z(n7937) );
  AND U9021 ( .A(n7938), .B(n7937), .Z(n7942) );
  XOR U9022 ( .A(n7943), .B(n7942), .Z(n7945) );
  XOR U9023 ( .A(n7944), .B(n7945), .Z(n7958) );
  XNOR U9024 ( .A(n7958), .B(sreg[1291]), .Z(n7960) );
  XOR U9025 ( .A(n7960), .B(n7959), .Z(c[1291]) );
  NANDN U9026 ( .A(n7943), .B(n7942), .Z(n7947) );
  OR U9027 ( .A(n7945), .B(n7944), .Z(n7946) );
  AND U9028 ( .A(n7947), .B(n7946), .Z(n7965) );
  XOR U9029 ( .A(a[270]), .B(n2214), .Z(n7969) );
  AND U9030 ( .A(a[272]), .B(b[0]), .Z(n7949) );
  XNOR U9031 ( .A(n7949), .B(n2175), .Z(n7951) );
  NANDN U9032 ( .A(b[0]), .B(a[271]), .Z(n7950) );
  NAND U9033 ( .A(n7951), .B(n7950), .Z(n7974) );
  AND U9034 ( .A(a[268]), .B(b[3]), .Z(n7973) );
  XOR U9035 ( .A(n7974), .B(n7973), .Z(n7976) );
  XOR U9036 ( .A(n7975), .B(n7976), .Z(n7964) );
  NANDN U9037 ( .A(n7953), .B(n7952), .Z(n7957) );
  OR U9038 ( .A(n7955), .B(n7954), .Z(n7956) );
  AND U9039 ( .A(n7957), .B(n7956), .Z(n7963) );
  XOR U9040 ( .A(n7964), .B(n7963), .Z(n7966) );
  XOR U9041 ( .A(n7965), .B(n7966), .Z(n7979) );
  XNOR U9042 ( .A(n7979), .B(sreg[1292]), .Z(n7981) );
  NANDN U9043 ( .A(n7958), .B(sreg[1291]), .Z(n7962) );
  NAND U9044 ( .A(n7960), .B(n7959), .Z(n7961) );
  NAND U9045 ( .A(n7962), .B(n7961), .Z(n7980) );
  XOR U9046 ( .A(n7981), .B(n7980), .Z(c[1292]) );
  NANDN U9047 ( .A(n7964), .B(n7963), .Z(n7968) );
  OR U9048 ( .A(n7966), .B(n7965), .Z(n7967) );
  AND U9049 ( .A(n7968), .B(n7967), .Z(n7986) );
  XOR U9050 ( .A(a[271]), .B(n2214), .Z(n7990) );
  AND U9051 ( .A(a[273]), .B(b[0]), .Z(n7970) );
  XNOR U9052 ( .A(n7970), .B(n2175), .Z(n7972) );
  NANDN U9053 ( .A(b[0]), .B(a[272]), .Z(n7971) );
  NAND U9054 ( .A(n7972), .B(n7971), .Z(n7995) );
  AND U9055 ( .A(a[269]), .B(b[3]), .Z(n7994) );
  XOR U9056 ( .A(n7995), .B(n7994), .Z(n7997) );
  XOR U9057 ( .A(n7996), .B(n7997), .Z(n7985) );
  NANDN U9058 ( .A(n7974), .B(n7973), .Z(n7978) );
  OR U9059 ( .A(n7976), .B(n7975), .Z(n7977) );
  AND U9060 ( .A(n7978), .B(n7977), .Z(n7984) );
  XOR U9061 ( .A(n7985), .B(n7984), .Z(n7987) );
  XOR U9062 ( .A(n7986), .B(n7987), .Z(n8000) );
  XNOR U9063 ( .A(n8000), .B(sreg[1293]), .Z(n8002) );
  NANDN U9064 ( .A(n7979), .B(sreg[1292]), .Z(n7983) );
  NAND U9065 ( .A(n7981), .B(n7980), .Z(n7982) );
  NAND U9066 ( .A(n7983), .B(n7982), .Z(n8001) );
  XOR U9067 ( .A(n8002), .B(n8001), .Z(c[1293]) );
  NANDN U9068 ( .A(n7985), .B(n7984), .Z(n7989) );
  OR U9069 ( .A(n7987), .B(n7986), .Z(n7988) );
  AND U9070 ( .A(n7989), .B(n7988), .Z(n8007) );
  XOR U9071 ( .A(a[272]), .B(n2215), .Z(n8011) );
  AND U9072 ( .A(a[274]), .B(b[0]), .Z(n7991) );
  XNOR U9073 ( .A(n7991), .B(n2175), .Z(n7993) );
  NANDN U9074 ( .A(b[0]), .B(a[273]), .Z(n7992) );
  NAND U9075 ( .A(n7993), .B(n7992), .Z(n8016) );
  AND U9076 ( .A(a[270]), .B(b[3]), .Z(n8015) );
  XOR U9077 ( .A(n8016), .B(n8015), .Z(n8018) );
  XOR U9078 ( .A(n8017), .B(n8018), .Z(n8006) );
  NANDN U9079 ( .A(n7995), .B(n7994), .Z(n7999) );
  OR U9080 ( .A(n7997), .B(n7996), .Z(n7998) );
  AND U9081 ( .A(n7999), .B(n7998), .Z(n8005) );
  XOR U9082 ( .A(n8006), .B(n8005), .Z(n8008) );
  XOR U9083 ( .A(n8007), .B(n8008), .Z(n8021) );
  XNOR U9084 ( .A(n8021), .B(sreg[1294]), .Z(n8023) );
  NANDN U9085 ( .A(n8000), .B(sreg[1293]), .Z(n8004) );
  NAND U9086 ( .A(n8002), .B(n8001), .Z(n8003) );
  NAND U9087 ( .A(n8004), .B(n8003), .Z(n8022) );
  XOR U9088 ( .A(n8023), .B(n8022), .Z(c[1294]) );
  NANDN U9089 ( .A(n8006), .B(n8005), .Z(n8010) );
  OR U9090 ( .A(n8008), .B(n8007), .Z(n8009) );
  AND U9091 ( .A(n8010), .B(n8009), .Z(n8028) );
  XOR U9092 ( .A(a[273]), .B(n2215), .Z(n8032) );
  AND U9093 ( .A(a[275]), .B(b[0]), .Z(n8012) );
  XNOR U9094 ( .A(n8012), .B(n2175), .Z(n8014) );
  NANDN U9095 ( .A(b[0]), .B(a[274]), .Z(n8013) );
  NAND U9096 ( .A(n8014), .B(n8013), .Z(n8037) );
  AND U9097 ( .A(a[271]), .B(b[3]), .Z(n8036) );
  XOR U9098 ( .A(n8037), .B(n8036), .Z(n8039) );
  XOR U9099 ( .A(n8038), .B(n8039), .Z(n8027) );
  NANDN U9100 ( .A(n8016), .B(n8015), .Z(n8020) );
  OR U9101 ( .A(n8018), .B(n8017), .Z(n8019) );
  AND U9102 ( .A(n8020), .B(n8019), .Z(n8026) );
  XOR U9103 ( .A(n8027), .B(n8026), .Z(n8029) );
  XOR U9104 ( .A(n8028), .B(n8029), .Z(n8042) );
  XNOR U9105 ( .A(n8042), .B(sreg[1295]), .Z(n8044) );
  NANDN U9106 ( .A(n8021), .B(sreg[1294]), .Z(n8025) );
  NAND U9107 ( .A(n8023), .B(n8022), .Z(n8024) );
  NAND U9108 ( .A(n8025), .B(n8024), .Z(n8043) );
  XOR U9109 ( .A(n8044), .B(n8043), .Z(c[1295]) );
  NANDN U9110 ( .A(n8027), .B(n8026), .Z(n8031) );
  OR U9111 ( .A(n8029), .B(n8028), .Z(n8030) );
  AND U9112 ( .A(n8031), .B(n8030), .Z(n8049) );
  XOR U9113 ( .A(a[274]), .B(n2215), .Z(n8053) );
  AND U9114 ( .A(a[272]), .B(b[3]), .Z(n8057) );
  AND U9115 ( .A(a[276]), .B(b[0]), .Z(n8033) );
  XNOR U9116 ( .A(n8033), .B(n2175), .Z(n8035) );
  NANDN U9117 ( .A(b[0]), .B(a[275]), .Z(n8034) );
  NAND U9118 ( .A(n8035), .B(n8034), .Z(n8058) );
  XOR U9119 ( .A(n8057), .B(n8058), .Z(n8060) );
  XOR U9120 ( .A(n8059), .B(n8060), .Z(n8048) );
  NANDN U9121 ( .A(n8037), .B(n8036), .Z(n8041) );
  OR U9122 ( .A(n8039), .B(n8038), .Z(n8040) );
  AND U9123 ( .A(n8041), .B(n8040), .Z(n8047) );
  XOR U9124 ( .A(n8048), .B(n8047), .Z(n8050) );
  XOR U9125 ( .A(n8049), .B(n8050), .Z(n8063) );
  XNOR U9126 ( .A(n8063), .B(sreg[1296]), .Z(n8065) );
  NANDN U9127 ( .A(n8042), .B(sreg[1295]), .Z(n8046) );
  NAND U9128 ( .A(n8044), .B(n8043), .Z(n8045) );
  NAND U9129 ( .A(n8046), .B(n8045), .Z(n8064) );
  XOR U9130 ( .A(n8065), .B(n8064), .Z(c[1296]) );
  NANDN U9131 ( .A(n8048), .B(n8047), .Z(n8052) );
  OR U9132 ( .A(n8050), .B(n8049), .Z(n8051) );
  AND U9133 ( .A(n8052), .B(n8051), .Z(n8070) );
  XOR U9134 ( .A(a[275]), .B(n2215), .Z(n8074) );
  AND U9135 ( .A(a[273]), .B(b[3]), .Z(n8078) );
  AND U9136 ( .A(a[277]), .B(b[0]), .Z(n8054) );
  XNOR U9137 ( .A(n8054), .B(n2175), .Z(n8056) );
  NANDN U9138 ( .A(b[0]), .B(a[276]), .Z(n8055) );
  NAND U9139 ( .A(n8056), .B(n8055), .Z(n8079) );
  XOR U9140 ( .A(n8078), .B(n8079), .Z(n8081) );
  XOR U9141 ( .A(n8080), .B(n8081), .Z(n8069) );
  NANDN U9142 ( .A(n8058), .B(n8057), .Z(n8062) );
  OR U9143 ( .A(n8060), .B(n8059), .Z(n8061) );
  AND U9144 ( .A(n8062), .B(n8061), .Z(n8068) );
  XOR U9145 ( .A(n8069), .B(n8068), .Z(n8071) );
  XOR U9146 ( .A(n8070), .B(n8071), .Z(n8084) );
  XNOR U9147 ( .A(n8084), .B(sreg[1297]), .Z(n8086) );
  NANDN U9148 ( .A(n8063), .B(sreg[1296]), .Z(n8067) );
  NAND U9149 ( .A(n8065), .B(n8064), .Z(n8066) );
  NAND U9150 ( .A(n8067), .B(n8066), .Z(n8085) );
  XOR U9151 ( .A(n8086), .B(n8085), .Z(c[1297]) );
  NANDN U9152 ( .A(n8069), .B(n8068), .Z(n8073) );
  OR U9153 ( .A(n8071), .B(n8070), .Z(n8072) );
  AND U9154 ( .A(n8073), .B(n8072), .Z(n8091) );
  XOR U9155 ( .A(a[276]), .B(n2215), .Z(n8095) );
  AND U9156 ( .A(a[278]), .B(b[0]), .Z(n8075) );
  XNOR U9157 ( .A(n8075), .B(n2175), .Z(n8077) );
  NANDN U9158 ( .A(b[0]), .B(a[277]), .Z(n8076) );
  NAND U9159 ( .A(n8077), .B(n8076), .Z(n8100) );
  AND U9160 ( .A(a[274]), .B(b[3]), .Z(n8099) );
  XOR U9161 ( .A(n8100), .B(n8099), .Z(n8102) );
  XOR U9162 ( .A(n8101), .B(n8102), .Z(n8090) );
  NANDN U9163 ( .A(n8079), .B(n8078), .Z(n8083) );
  OR U9164 ( .A(n8081), .B(n8080), .Z(n8082) );
  AND U9165 ( .A(n8083), .B(n8082), .Z(n8089) );
  XOR U9166 ( .A(n8090), .B(n8089), .Z(n8092) );
  XOR U9167 ( .A(n8091), .B(n8092), .Z(n8105) );
  XNOR U9168 ( .A(n8105), .B(sreg[1298]), .Z(n8107) );
  NANDN U9169 ( .A(n8084), .B(sreg[1297]), .Z(n8088) );
  NAND U9170 ( .A(n8086), .B(n8085), .Z(n8087) );
  NAND U9171 ( .A(n8088), .B(n8087), .Z(n8106) );
  XOR U9172 ( .A(n8107), .B(n8106), .Z(c[1298]) );
  NANDN U9173 ( .A(n8090), .B(n8089), .Z(n8094) );
  OR U9174 ( .A(n8092), .B(n8091), .Z(n8093) );
  AND U9175 ( .A(n8094), .B(n8093), .Z(n8112) );
  XOR U9176 ( .A(a[277]), .B(n2215), .Z(n8116) );
  AND U9177 ( .A(a[275]), .B(b[3]), .Z(n8120) );
  AND U9178 ( .A(a[279]), .B(b[0]), .Z(n8096) );
  XNOR U9179 ( .A(n8096), .B(n2175), .Z(n8098) );
  NANDN U9180 ( .A(b[0]), .B(a[278]), .Z(n8097) );
  NAND U9181 ( .A(n8098), .B(n8097), .Z(n8121) );
  XOR U9182 ( .A(n8120), .B(n8121), .Z(n8123) );
  XOR U9183 ( .A(n8122), .B(n8123), .Z(n8111) );
  NANDN U9184 ( .A(n8100), .B(n8099), .Z(n8104) );
  OR U9185 ( .A(n8102), .B(n8101), .Z(n8103) );
  AND U9186 ( .A(n8104), .B(n8103), .Z(n8110) );
  XOR U9187 ( .A(n8111), .B(n8110), .Z(n8113) );
  XOR U9188 ( .A(n8112), .B(n8113), .Z(n8126) );
  XNOR U9189 ( .A(n8126), .B(sreg[1299]), .Z(n8128) );
  NANDN U9190 ( .A(n8105), .B(sreg[1298]), .Z(n8109) );
  NAND U9191 ( .A(n8107), .B(n8106), .Z(n8108) );
  NAND U9192 ( .A(n8109), .B(n8108), .Z(n8127) );
  XOR U9193 ( .A(n8128), .B(n8127), .Z(c[1299]) );
  NANDN U9194 ( .A(n8111), .B(n8110), .Z(n8115) );
  OR U9195 ( .A(n8113), .B(n8112), .Z(n8114) );
  AND U9196 ( .A(n8115), .B(n8114), .Z(n8133) );
  XOR U9197 ( .A(a[278]), .B(n2215), .Z(n8137) );
  AND U9198 ( .A(a[280]), .B(b[0]), .Z(n8117) );
  XNOR U9199 ( .A(n8117), .B(n2175), .Z(n8119) );
  NANDN U9200 ( .A(b[0]), .B(a[279]), .Z(n8118) );
  NAND U9201 ( .A(n8119), .B(n8118), .Z(n8142) );
  AND U9202 ( .A(a[276]), .B(b[3]), .Z(n8141) );
  XOR U9203 ( .A(n8142), .B(n8141), .Z(n8144) );
  XOR U9204 ( .A(n8143), .B(n8144), .Z(n8132) );
  NANDN U9205 ( .A(n8121), .B(n8120), .Z(n8125) );
  OR U9206 ( .A(n8123), .B(n8122), .Z(n8124) );
  AND U9207 ( .A(n8125), .B(n8124), .Z(n8131) );
  XOR U9208 ( .A(n8132), .B(n8131), .Z(n8134) );
  XOR U9209 ( .A(n8133), .B(n8134), .Z(n8147) );
  XNOR U9210 ( .A(n8147), .B(sreg[1300]), .Z(n8149) );
  NANDN U9211 ( .A(n8126), .B(sreg[1299]), .Z(n8130) );
  NAND U9212 ( .A(n8128), .B(n8127), .Z(n8129) );
  NAND U9213 ( .A(n8130), .B(n8129), .Z(n8148) );
  XOR U9214 ( .A(n8149), .B(n8148), .Z(c[1300]) );
  NANDN U9215 ( .A(n8132), .B(n8131), .Z(n8136) );
  OR U9216 ( .A(n8134), .B(n8133), .Z(n8135) );
  AND U9217 ( .A(n8136), .B(n8135), .Z(n8154) );
  XOR U9218 ( .A(a[279]), .B(n2216), .Z(n8158) );
  AND U9219 ( .A(a[281]), .B(b[0]), .Z(n8138) );
  XNOR U9220 ( .A(n8138), .B(n2175), .Z(n8140) );
  NANDN U9221 ( .A(b[0]), .B(a[280]), .Z(n8139) );
  NAND U9222 ( .A(n8140), .B(n8139), .Z(n8163) );
  AND U9223 ( .A(a[277]), .B(b[3]), .Z(n8162) );
  XOR U9224 ( .A(n8163), .B(n8162), .Z(n8165) );
  XOR U9225 ( .A(n8164), .B(n8165), .Z(n8153) );
  NANDN U9226 ( .A(n8142), .B(n8141), .Z(n8146) );
  OR U9227 ( .A(n8144), .B(n8143), .Z(n8145) );
  AND U9228 ( .A(n8146), .B(n8145), .Z(n8152) );
  XOR U9229 ( .A(n8153), .B(n8152), .Z(n8155) );
  XOR U9230 ( .A(n8154), .B(n8155), .Z(n8168) );
  XNOR U9231 ( .A(n8168), .B(sreg[1301]), .Z(n8170) );
  NANDN U9232 ( .A(n8147), .B(sreg[1300]), .Z(n8151) );
  NAND U9233 ( .A(n8149), .B(n8148), .Z(n8150) );
  NAND U9234 ( .A(n8151), .B(n8150), .Z(n8169) );
  XOR U9235 ( .A(n8170), .B(n8169), .Z(c[1301]) );
  NANDN U9236 ( .A(n8153), .B(n8152), .Z(n8157) );
  OR U9237 ( .A(n8155), .B(n8154), .Z(n8156) );
  AND U9238 ( .A(n8157), .B(n8156), .Z(n8175) );
  XOR U9239 ( .A(a[280]), .B(n2216), .Z(n8179) );
  AND U9240 ( .A(a[282]), .B(b[0]), .Z(n8159) );
  XNOR U9241 ( .A(n8159), .B(n2175), .Z(n8161) );
  NANDN U9242 ( .A(b[0]), .B(a[281]), .Z(n8160) );
  NAND U9243 ( .A(n8161), .B(n8160), .Z(n8184) );
  AND U9244 ( .A(a[278]), .B(b[3]), .Z(n8183) );
  XOR U9245 ( .A(n8184), .B(n8183), .Z(n8186) );
  XOR U9246 ( .A(n8185), .B(n8186), .Z(n8174) );
  NANDN U9247 ( .A(n8163), .B(n8162), .Z(n8167) );
  OR U9248 ( .A(n8165), .B(n8164), .Z(n8166) );
  AND U9249 ( .A(n8167), .B(n8166), .Z(n8173) );
  XOR U9250 ( .A(n8174), .B(n8173), .Z(n8176) );
  XOR U9251 ( .A(n8175), .B(n8176), .Z(n8189) );
  XNOR U9252 ( .A(n8189), .B(sreg[1302]), .Z(n8191) );
  NANDN U9253 ( .A(n8168), .B(sreg[1301]), .Z(n8172) );
  NAND U9254 ( .A(n8170), .B(n8169), .Z(n8171) );
  NAND U9255 ( .A(n8172), .B(n8171), .Z(n8190) );
  XOR U9256 ( .A(n8191), .B(n8190), .Z(c[1302]) );
  NANDN U9257 ( .A(n8174), .B(n8173), .Z(n8178) );
  OR U9258 ( .A(n8176), .B(n8175), .Z(n8177) );
  AND U9259 ( .A(n8178), .B(n8177), .Z(n8197) );
  XOR U9260 ( .A(a[281]), .B(n2216), .Z(n8198) );
  AND U9261 ( .A(b[0]), .B(a[283]), .Z(n8180) );
  XOR U9262 ( .A(b[1]), .B(n8180), .Z(n8182) );
  NANDN U9263 ( .A(b[0]), .B(a[282]), .Z(n8181) );
  AND U9264 ( .A(n8182), .B(n8181), .Z(n8202) );
  AND U9265 ( .A(a[279]), .B(b[3]), .Z(n8203) );
  XOR U9266 ( .A(n8202), .B(n8203), .Z(n8204) );
  XNOR U9267 ( .A(n8205), .B(n8204), .Z(n8194) );
  NANDN U9268 ( .A(n8184), .B(n8183), .Z(n8188) );
  OR U9269 ( .A(n8186), .B(n8185), .Z(n8187) );
  AND U9270 ( .A(n8188), .B(n8187), .Z(n8195) );
  XNOR U9271 ( .A(n8194), .B(n8195), .Z(n8196) );
  XNOR U9272 ( .A(n8197), .B(n8196), .Z(n8208) );
  XNOR U9273 ( .A(n8208), .B(sreg[1303]), .Z(n8210) );
  NANDN U9274 ( .A(n8189), .B(sreg[1302]), .Z(n8193) );
  NAND U9275 ( .A(n8191), .B(n8190), .Z(n8192) );
  NAND U9276 ( .A(n8193), .B(n8192), .Z(n8209) );
  XOR U9277 ( .A(n8210), .B(n8209), .Z(c[1303]) );
  XOR U9278 ( .A(a[282]), .B(n2216), .Z(n8217) );
  AND U9279 ( .A(a[284]), .B(b[0]), .Z(n8199) );
  XNOR U9280 ( .A(n8199), .B(n2175), .Z(n8201) );
  NANDN U9281 ( .A(b[0]), .B(a[283]), .Z(n8200) );
  NAND U9282 ( .A(n8201), .B(n8200), .Z(n8222) );
  AND U9283 ( .A(a[280]), .B(b[3]), .Z(n8221) );
  XOR U9284 ( .A(n8222), .B(n8221), .Z(n8224) );
  XOR U9285 ( .A(n8223), .B(n8224), .Z(n8212) );
  NAND U9286 ( .A(n8203), .B(n8202), .Z(n8207) );
  NANDN U9287 ( .A(n8205), .B(n8204), .Z(n8206) );
  AND U9288 ( .A(n8207), .B(n8206), .Z(n8211) );
  XOR U9289 ( .A(n8212), .B(n8211), .Z(n8214) );
  XOR U9290 ( .A(n8213), .B(n8214), .Z(n8227) );
  XNOR U9291 ( .A(n8227), .B(sreg[1304]), .Z(n8229) );
  XOR U9292 ( .A(n8229), .B(n8228), .Z(c[1304]) );
  NANDN U9293 ( .A(n8212), .B(n8211), .Z(n8216) );
  OR U9294 ( .A(n8214), .B(n8213), .Z(n8215) );
  AND U9295 ( .A(n8216), .B(n8215), .Z(n8234) );
  XOR U9296 ( .A(a[283]), .B(n2216), .Z(n8238) );
  AND U9297 ( .A(a[285]), .B(b[0]), .Z(n8218) );
  XNOR U9298 ( .A(n8218), .B(n2175), .Z(n8220) );
  NANDN U9299 ( .A(b[0]), .B(a[284]), .Z(n8219) );
  NAND U9300 ( .A(n8220), .B(n8219), .Z(n8243) );
  AND U9301 ( .A(a[281]), .B(b[3]), .Z(n8242) );
  XOR U9302 ( .A(n8243), .B(n8242), .Z(n8245) );
  XOR U9303 ( .A(n8244), .B(n8245), .Z(n8233) );
  NANDN U9304 ( .A(n8222), .B(n8221), .Z(n8226) );
  OR U9305 ( .A(n8224), .B(n8223), .Z(n8225) );
  AND U9306 ( .A(n8226), .B(n8225), .Z(n8232) );
  XOR U9307 ( .A(n8233), .B(n8232), .Z(n8235) );
  XOR U9308 ( .A(n8234), .B(n8235), .Z(n8248) );
  XNOR U9309 ( .A(n8248), .B(sreg[1305]), .Z(n8250) );
  NANDN U9310 ( .A(n8227), .B(sreg[1304]), .Z(n8231) );
  NAND U9311 ( .A(n8229), .B(n8228), .Z(n8230) );
  NAND U9312 ( .A(n8231), .B(n8230), .Z(n8249) );
  XOR U9313 ( .A(n8250), .B(n8249), .Z(c[1305]) );
  NANDN U9314 ( .A(n8233), .B(n8232), .Z(n8237) );
  OR U9315 ( .A(n8235), .B(n8234), .Z(n8236) );
  AND U9316 ( .A(n8237), .B(n8236), .Z(n8255) );
  XOR U9317 ( .A(a[284]), .B(n2216), .Z(n8259) );
  AND U9318 ( .A(a[286]), .B(b[0]), .Z(n8239) );
  XNOR U9319 ( .A(n8239), .B(n2175), .Z(n8241) );
  NANDN U9320 ( .A(b[0]), .B(a[285]), .Z(n8240) );
  NAND U9321 ( .A(n8241), .B(n8240), .Z(n8264) );
  AND U9322 ( .A(a[282]), .B(b[3]), .Z(n8263) );
  XOR U9323 ( .A(n8264), .B(n8263), .Z(n8266) );
  XOR U9324 ( .A(n8265), .B(n8266), .Z(n8254) );
  NANDN U9325 ( .A(n8243), .B(n8242), .Z(n8247) );
  OR U9326 ( .A(n8245), .B(n8244), .Z(n8246) );
  AND U9327 ( .A(n8247), .B(n8246), .Z(n8253) );
  XOR U9328 ( .A(n8254), .B(n8253), .Z(n8256) );
  XOR U9329 ( .A(n8255), .B(n8256), .Z(n8269) );
  XNOR U9330 ( .A(n8269), .B(sreg[1306]), .Z(n8271) );
  NANDN U9331 ( .A(n8248), .B(sreg[1305]), .Z(n8252) );
  NAND U9332 ( .A(n8250), .B(n8249), .Z(n8251) );
  NAND U9333 ( .A(n8252), .B(n8251), .Z(n8270) );
  XOR U9334 ( .A(n8271), .B(n8270), .Z(c[1306]) );
  NANDN U9335 ( .A(n8254), .B(n8253), .Z(n8258) );
  OR U9336 ( .A(n8256), .B(n8255), .Z(n8257) );
  AND U9337 ( .A(n8258), .B(n8257), .Z(n8276) );
  XOR U9338 ( .A(a[285]), .B(n2216), .Z(n8280) );
  AND U9339 ( .A(a[287]), .B(b[0]), .Z(n8260) );
  XNOR U9340 ( .A(n8260), .B(n2175), .Z(n8262) );
  NANDN U9341 ( .A(b[0]), .B(a[286]), .Z(n8261) );
  NAND U9342 ( .A(n8262), .B(n8261), .Z(n8285) );
  AND U9343 ( .A(a[283]), .B(b[3]), .Z(n8284) );
  XOR U9344 ( .A(n8285), .B(n8284), .Z(n8287) );
  XOR U9345 ( .A(n8286), .B(n8287), .Z(n8275) );
  NANDN U9346 ( .A(n8264), .B(n8263), .Z(n8268) );
  OR U9347 ( .A(n8266), .B(n8265), .Z(n8267) );
  AND U9348 ( .A(n8268), .B(n8267), .Z(n8274) );
  XOR U9349 ( .A(n8275), .B(n8274), .Z(n8277) );
  XOR U9350 ( .A(n8276), .B(n8277), .Z(n8290) );
  XNOR U9351 ( .A(n8290), .B(sreg[1307]), .Z(n8292) );
  NANDN U9352 ( .A(n8269), .B(sreg[1306]), .Z(n8273) );
  NAND U9353 ( .A(n8271), .B(n8270), .Z(n8272) );
  NAND U9354 ( .A(n8273), .B(n8272), .Z(n8291) );
  XOR U9355 ( .A(n8292), .B(n8291), .Z(c[1307]) );
  NANDN U9356 ( .A(n8275), .B(n8274), .Z(n8279) );
  OR U9357 ( .A(n8277), .B(n8276), .Z(n8278) );
  AND U9358 ( .A(n8279), .B(n8278), .Z(n8297) );
  XOR U9359 ( .A(a[286]), .B(n2217), .Z(n8301) );
  AND U9360 ( .A(a[284]), .B(b[3]), .Z(n8305) );
  AND U9361 ( .A(a[288]), .B(b[0]), .Z(n8281) );
  XNOR U9362 ( .A(n8281), .B(n2175), .Z(n8283) );
  NANDN U9363 ( .A(b[0]), .B(a[287]), .Z(n8282) );
  NAND U9364 ( .A(n8283), .B(n8282), .Z(n8306) );
  XOR U9365 ( .A(n8305), .B(n8306), .Z(n8308) );
  XOR U9366 ( .A(n8307), .B(n8308), .Z(n8296) );
  NANDN U9367 ( .A(n8285), .B(n8284), .Z(n8289) );
  OR U9368 ( .A(n8287), .B(n8286), .Z(n8288) );
  AND U9369 ( .A(n8289), .B(n8288), .Z(n8295) );
  XOR U9370 ( .A(n8296), .B(n8295), .Z(n8298) );
  XOR U9371 ( .A(n8297), .B(n8298), .Z(n8311) );
  XNOR U9372 ( .A(n8311), .B(sreg[1308]), .Z(n8313) );
  NANDN U9373 ( .A(n8290), .B(sreg[1307]), .Z(n8294) );
  NAND U9374 ( .A(n8292), .B(n8291), .Z(n8293) );
  NAND U9375 ( .A(n8294), .B(n8293), .Z(n8312) );
  XOR U9376 ( .A(n8313), .B(n8312), .Z(c[1308]) );
  NANDN U9377 ( .A(n8296), .B(n8295), .Z(n8300) );
  OR U9378 ( .A(n8298), .B(n8297), .Z(n8299) );
  AND U9379 ( .A(n8300), .B(n8299), .Z(n8318) );
  XOR U9380 ( .A(a[287]), .B(n2217), .Z(n8322) );
  AND U9381 ( .A(a[285]), .B(b[3]), .Z(n8326) );
  AND U9382 ( .A(a[289]), .B(b[0]), .Z(n8302) );
  XNOR U9383 ( .A(n8302), .B(n2175), .Z(n8304) );
  NANDN U9384 ( .A(b[0]), .B(a[288]), .Z(n8303) );
  NAND U9385 ( .A(n8304), .B(n8303), .Z(n8327) );
  XOR U9386 ( .A(n8326), .B(n8327), .Z(n8329) );
  XOR U9387 ( .A(n8328), .B(n8329), .Z(n8317) );
  NANDN U9388 ( .A(n8306), .B(n8305), .Z(n8310) );
  OR U9389 ( .A(n8308), .B(n8307), .Z(n8309) );
  AND U9390 ( .A(n8310), .B(n8309), .Z(n8316) );
  XOR U9391 ( .A(n8317), .B(n8316), .Z(n8319) );
  XOR U9392 ( .A(n8318), .B(n8319), .Z(n8332) );
  XNOR U9393 ( .A(n8332), .B(sreg[1309]), .Z(n8334) );
  NANDN U9394 ( .A(n8311), .B(sreg[1308]), .Z(n8315) );
  NAND U9395 ( .A(n8313), .B(n8312), .Z(n8314) );
  NAND U9396 ( .A(n8315), .B(n8314), .Z(n8333) );
  XOR U9397 ( .A(n8334), .B(n8333), .Z(c[1309]) );
  NANDN U9398 ( .A(n8317), .B(n8316), .Z(n8321) );
  OR U9399 ( .A(n8319), .B(n8318), .Z(n8320) );
  AND U9400 ( .A(n8321), .B(n8320), .Z(n8339) );
  XOR U9401 ( .A(a[288]), .B(n2217), .Z(n8343) );
  AND U9402 ( .A(a[290]), .B(b[0]), .Z(n8323) );
  XNOR U9403 ( .A(n8323), .B(n2175), .Z(n8325) );
  NANDN U9404 ( .A(b[0]), .B(a[289]), .Z(n8324) );
  NAND U9405 ( .A(n8325), .B(n8324), .Z(n8348) );
  AND U9406 ( .A(a[286]), .B(b[3]), .Z(n8347) );
  XOR U9407 ( .A(n8348), .B(n8347), .Z(n8350) );
  XOR U9408 ( .A(n8349), .B(n8350), .Z(n8338) );
  NANDN U9409 ( .A(n8327), .B(n8326), .Z(n8331) );
  OR U9410 ( .A(n8329), .B(n8328), .Z(n8330) );
  AND U9411 ( .A(n8331), .B(n8330), .Z(n8337) );
  XOR U9412 ( .A(n8338), .B(n8337), .Z(n8340) );
  XOR U9413 ( .A(n8339), .B(n8340), .Z(n8353) );
  XNOR U9414 ( .A(n8353), .B(sreg[1310]), .Z(n8355) );
  NANDN U9415 ( .A(n8332), .B(sreg[1309]), .Z(n8336) );
  NAND U9416 ( .A(n8334), .B(n8333), .Z(n8335) );
  NAND U9417 ( .A(n8336), .B(n8335), .Z(n8354) );
  XOR U9418 ( .A(n8355), .B(n8354), .Z(c[1310]) );
  NANDN U9419 ( .A(n8338), .B(n8337), .Z(n8342) );
  OR U9420 ( .A(n8340), .B(n8339), .Z(n8341) );
  AND U9421 ( .A(n8342), .B(n8341), .Z(n8360) );
  XOR U9422 ( .A(a[289]), .B(n2217), .Z(n8364) );
  AND U9423 ( .A(a[291]), .B(b[0]), .Z(n8344) );
  XNOR U9424 ( .A(n8344), .B(n2175), .Z(n8346) );
  NANDN U9425 ( .A(b[0]), .B(a[290]), .Z(n8345) );
  NAND U9426 ( .A(n8346), .B(n8345), .Z(n8369) );
  AND U9427 ( .A(a[287]), .B(b[3]), .Z(n8368) );
  XOR U9428 ( .A(n8369), .B(n8368), .Z(n8371) );
  XOR U9429 ( .A(n8370), .B(n8371), .Z(n8359) );
  NANDN U9430 ( .A(n8348), .B(n8347), .Z(n8352) );
  OR U9431 ( .A(n8350), .B(n8349), .Z(n8351) );
  AND U9432 ( .A(n8352), .B(n8351), .Z(n8358) );
  XOR U9433 ( .A(n8359), .B(n8358), .Z(n8361) );
  XOR U9434 ( .A(n8360), .B(n8361), .Z(n8374) );
  XNOR U9435 ( .A(n8374), .B(sreg[1311]), .Z(n8376) );
  NANDN U9436 ( .A(n8353), .B(sreg[1310]), .Z(n8357) );
  NAND U9437 ( .A(n8355), .B(n8354), .Z(n8356) );
  NAND U9438 ( .A(n8357), .B(n8356), .Z(n8375) );
  XOR U9439 ( .A(n8376), .B(n8375), .Z(c[1311]) );
  NANDN U9440 ( .A(n8359), .B(n8358), .Z(n8363) );
  OR U9441 ( .A(n8361), .B(n8360), .Z(n8362) );
  AND U9442 ( .A(n8363), .B(n8362), .Z(n8381) );
  XOR U9443 ( .A(a[290]), .B(n2217), .Z(n8385) );
  AND U9444 ( .A(a[292]), .B(b[0]), .Z(n8365) );
  XNOR U9445 ( .A(n8365), .B(n2175), .Z(n8367) );
  NANDN U9446 ( .A(b[0]), .B(a[291]), .Z(n8366) );
  NAND U9447 ( .A(n8367), .B(n8366), .Z(n8390) );
  AND U9448 ( .A(a[288]), .B(b[3]), .Z(n8389) );
  XOR U9449 ( .A(n8390), .B(n8389), .Z(n8392) );
  XOR U9450 ( .A(n8391), .B(n8392), .Z(n8380) );
  NANDN U9451 ( .A(n8369), .B(n8368), .Z(n8373) );
  OR U9452 ( .A(n8371), .B(n8370), .Z(n8372) );
  AND U9453 ( .A(n8373), .B(n8372), .Z(n8379) );
  XOR U9454 ( .A(n8380), .B(n8379), .Z(n8382) );
  XOR U9455 ( .A(n8381), .B(n8382), .Z(n8395) );
  XNOR U9456 ( .A(n8395), .B(sreg[1312]), .Z(n8397) );
  NANDN U9457 ( .A(n8374), .B(sreg[1311]), .Z(n8378) );
  NAND U9458 ( .A(n8376), .B(n8375), .Z(n8377) );
  NAND U9459 ( .A(n8378), .B(n8377), .Z(n8396) );
  XOR U9460 ( .A(n8397), .B(n8396), .Z(c[1312]) );
  NANDN U9461 ( .A(n8380), .B(n8379), .Z(n8384) );
  OR U9462 ( .A(n8382), .B(n8381), .Z(n8383) );
  AND U9463 ( .A(n8384), .B(n8383), .Z(n8402) );
  XOR U9464 ( .A(a[291]), .B(n2217), .Z(n8406) );
  AND U9465 ( .A(a[293]), .B(b[0]), .Z(n8386) );
  XNOR U9466 ( .A(n8386), .B(n2175), .Z(n8388) );
  NANDN U9467 ( .A(b[0]), .B(a[292]), .Z(n8387) );
  NAND U9468 ( .A(n8388), .B(n8387), .Z(n8411) );
  AND U9469 ( .A(a[289]), .B(b[3]), .Z(n8410) );
  XOR U9470 ( .A(n8411), .B(n8410), .Z(n8413) );
  XOR U9471 ( .A(n8412), .B(n8413), .Z(n8401) );
  NANDN U9472 ( .A(n8390), .B(n8389), .Z(n8394) );
  OR U9473 ( .A(n8392), .B(n8391), .Z(n8393) );
  AND U9474 ( .A(n8394), .B(n8393), .Z(n8400) );
  XOR U9475 ( .A(n8401), .B(n8400), .Z(n8403) );
  XOR U9476 ( .A(n8402), .B(n8403), .Z(n8416) );
  XNOR U9477 ( .A(n8416), .B(sreg[1313]), .Z(n8418) );
  NANDN U9478 ( .A(n8395), .B(sreg[1312]), .Z(n8399) );
  NAND U9479 ( .A(n8397), .B(n8396), .Z(n8398) );
  NAND U9480 ( .A(n8399), .B(n8398), .Z(n8417) );
  XOR U9481 ( .A(n8418), .B(n8417), .Z(c[1313]) );
  NANDN U9482 ( .A(n8401), .B(n8400), .Z(n8405) );
  OR U9483 ( .A(n8403), .B(n8402), .Z(n8404) );
  AND U9484 ( .A(n8405), .B(n8404), .Z(n8423) );
  XOR U9485 ( .A(a[292]), .B(n2217), .Z(n8427) );
  AND U9486 ( .A(a[294]), .B(b[0]), .Z(n8407) );
  XNOR U9487 ( .A(n8407), .B(n2175), .Z(n8409) );
  NANDN U9488 ( .A(b[0]), .B(a[293]), .Z(n8408) );
  NAND U9489 ( .A(n8409), .B(n8408), .Z(n8432) );
  AND U9490 ( .A(a[290]), .B(b[3]), .Z(n8431) );
  XOR U9491 ( .A(n8432), .B(n8431), .Z(n8434) );
  XOR U9492 ( .A(n8433), .B(n8434), .Z(n8422) );
  NANDN U9493 ( .A(n8411), .B(n8410), .Z(n8415) );
  OR U9494 ( .A(n8413), .B(n8412), .Z(n8414) );
  AND U9495 ( .A(n8415), .B(n8414), .Z(n8421) );
  XOR U9496 ( .A(n8422), .B(n8421), .Z(n8424) );
  XOR U9497 ( .A(n8423), .B(n8424), .Z(n8437) );
  XNOR U9498 ( .A(n8437), .B(sreg[1314]), .Z(n8439) );
  NANDN U9499 ( .A(n8416), .B(sreg[1313]), .Z(n8420) );
  NAND U9500 ( .A(n8418), .B(n8417), .Z(n8419) );
  NAND U9501 ( .A(n8420), .B(n8419), .Z(n8438) );
  XOR U9502 ( .A(n8439), .B(n8438), .Z(c[1314]) );
  NANDN U9503 ( .A(n8422), .B(n8421), .Z(n8426) );
  OR U9504 ( .A(n8424), .B(n8423), .Z(n8425) );
  AND U9505 ( .A(n8426), .B(n8425), .Z(n8444) );
  XOR U9506 ( .A(a[293]), .B(n2218), .Z(n8448) );
  AND U9507 ( .A(a[295]), .B(b[0]), .Z(n8428) );
  XNOR U9508 ( .A(n8428), .B(n2175), .Z(n8430) );
  NANDN U9509 ( .A(b[0]), .B(a[294]), .Z(n8429) );
  NAND U9510 ( .A(n8430), .B(n8429), .Z(n8453) );
  AND U9511 ( .A(a[291]), .B(b[3]), .Z(n8452) );
  XOR U9512 ( .A(n8453), .B(n8452), .Z(n8455) );
  XOR U9513 ( .A(n8454), .B(n8455), .Z(n8443) );
  NANDN U9514 ( .A(n8432), .B(n8431), .Z(n8436) );
  OR U9515 ( .A(n8434), .B(n8433), .Z(n8435) );
  AND U9516 ( .A(n8436), .B(n8435), .Z(n8442) );
  XOR U9517 ( .A(n8443), .B(n8442), .Z(n8445) );
  XOR U9518 ( .A(n8444), .B(n8445), .Z(n8458) );
  XNOR U9519 ( .A(n8458), .B(sreg[1315]), .Z(n8460) );
  NANDN U9520 ( .A(n8437), .B(sreg[1314]), .Z(n8441) );
  NAND U9521 ( .A(n8439), .B(n8438), .Z(n8440) );
  NAND U9522 ( .A(n8441), .B(n8440), .Z(n8459) );
  XOR U9523 ( .A(n8460), .B(n8459), .Z(c[1315]) );
  NANDN U9524 ( .A(n8443), .B(n8442), .Z(n8447) );
  OR U9525 ( .A(n8445), .B(n8444), .Z(n8446) );
  AND U9526 ( .A(n8447), .B(n8446), .Z(n8465) );
  XOR U9527 ( .A(a[294]), .B(n2218), .Z(n8469) );
  AND U9528 ( .A(a[292]), .B(b[3]), .Z(n8473) );
  AND U9529 ( .A(a[296]), .B(b[0]), .Z(n8449) );
  XNOR U9530 ( .A(n8449), .B(n2175), .Z(n8451) );
  NANDN U9531 ( .A(b[0]), .B(a[295]), .Z(n8450) );
  NAND U9532 ( .A(n8451), .B(n8450), .Z(n8474) );
  XOR U9533 ( .A(n8473), .B(n8474), .Z(n8476) );
  XOR U9534 ( .A(n8475), .B(n8476), .Z(n8464) );
  NANDN U9535 ( .A(n8453), .B(n8452), .Z(n8457) );
  OR U9536 ( .A(n8455), .B(n8454), .Z(n8456) );
  AND U9537 ( .A(n8457), .B(n8456), .Z(n8463) );
  XOR U9538 ( .A(n8464), .B(n8463), .Z(n8466) );
  XOR U9539 ( .A(n8465), .B(n8466), .Z(n8479) );
  XNOR U9540 ( .A(n8479), .B(sreg[1316]), .Z(n8481) );
  NANDN U9541 ( .A(n8458), .B(sreg[1315]), .Z(n8462) );
  NAND U9542 ( .A(n8460), .B(n8459), .Z(n8461) );
  NAND U9543 ( .A(n8462), .B(n8461), .Z(n8480) );
  XOR U9544 ( .A(n8481), .B(n8480), .Z(c[1316]) );
  NANDN U9545 ( .A(n8464), .B(n8463), .Z(n8468) );
  OR U9546 ( .A(n8466), .B(n8465), .Z(n8467) );
  AND U9547 ( .A(n8468), .B(n8467), .Z(n8486) );
  XOR U9548 ( .A(a[295]), .B(n2218), .Z(n8490) );
  AND U9549 ( .A(a[297]), .B(b[0]), .Z(n8470) );
  XNOR U9550 ( .A(n8470), .B(n2175), .Z(n8472) );
  NANDN U9551 ( .A(b[0]), .B(a[296]), .Z(n8471) );
  NAND U9552 ( .A(n8472), .B(n8471), .Z(n8495) );
  AND U9553 ( .A(a[293]), .B(b[3]), .Z(n8494) );
  XOR U9554 ( .A(n8495), .B(n8494), .Z(n8497) );
  XOR U9555 ( .A(n8496), .B(n8497), .Z(n8485) );
  NANDN U9556 ( .A(n8474), .B(n8473), .Z(n8478) );
  OR U9557 ( .A(n8476), .B(n8475), .Z(n8477) );
  AND U9558 ( .A(n8478), .B(n8477), .Z(n8484) );
  XOR U9559 ( .A(n8485), .B(n8484), .Z(n8487) );
  XOR U9560 ( .A(n8486), .B(n8487), .Z(n8500) );
  XNOR U9561 ( .A(n8500), .B(sreg[1317]), .Z(n8502) );
  NANDN U9562 ( .A(n8479), .B(sreg[1316]), .Z(n8483) );
  NAND U9563 ( .A(n8481), .B(n8480), .Z(n8482) );
  NAND U9564 ( .A(n8483), .B(n8482), .Z(n8501) );
  XOR U9565 ( .A(n8502), .B(n8501), .Z(c[1317]) );
  NANDN U9566 ( .A(n8485), .B(n8484), .Z(n8489) );
  OR U9567 ( .A(n8487), .B(n8486), .Z(n8488) );
  AND U9568 ( .A(n8489), .B(n8488), .Z(n8507) );
  XOR U9569 ( .A(a[296]), .B(n2218), .Z(n8511) );
  AND U9570 ( .A(a[298]), .B(b[0]), .Z(n8491) );
  XNOR U9571 ( .A(n8491), .B(n2175), .Z(n8493) );
  NANDN U9572 ( .A(b[0]), .B(a[297]), .Z(n8492) );
  NAND U9573 ( .A(n8493), .B(n8492), .Z(n8516) );
  AND U9574 ( .A(a[294]), .B(b[3]), .Z(n8515) );
  XOR U9575 ( .A(n8516), .B(n8515), .Z(n8518) );
  XOR U9576 ( .A(n8517), .B(n8518), .Z(n8506) );
  NANDN U9577 ( .A(n8495), .B(n8494), .Z(n8499) );
  OR U9578 ( .A(n8497), .B(n8496), .Z(n8498) );
  AND U9579 ( .A(n8499), .B(n8498), .Z(n8505) );
  XOR U9580 ( .A(n8506), .B(n8505), .Z(n8508) );
  XOR U9581 ( .A(n8507), .B(n8508), .Z(n8521) );
  XNOR U9582 ( .A(n8521), .B(sreg[1318]), .Z(n8523) );
  NANDN U9583 ( .A(n8500), .B(sreg[1317]), .Z(n8504) );
  NAND U9584 ( .A(n8502), .B(n8501), .Z(n8503) );
  NAND U9585 ( .A(n8504), .B(n8503), .Z(n8522) );
  XOR U9586 ( .A(n8523), .B(n8522), .Z(c[1318]) );
  NANDN U9587 ( .A(n8506), .B(n8505), .Z(n8510) );
  OR U9588 ( .A(n8508), .B(n8507), .Z(n8509) );
  AND U9589 ( .A(n8510), .B(n8509), .Z(n8528) );
  XOR U9590 ( .A(a[297]), .B(n2218), .Z(n8532) );
  AND U9591 ( .A(a[299]), .B(b[0]), .Z(n8512) );
  XNOR U9592 ( .A(n8512), .B(n2175), .Z(n8514) );
  NANDN U9593 ( .A(b[0]), .B(a[298]), .Z(n8513) );
  NAND U9594 ( .A(n8514), .B(n8513), .Z(n8537) );
  AND U9595 ( .A(a[295]), .B(b[3]), .Z(n8536) );
  XOR U9596 ( .A(n8537), .B(n8536), .Z(n8539) );
  XOR U9597 ( .A(n8538), .B(n8539), .Z(n8527) );
  NANDN U9598 ( .A(n8516), .B(n8515), .Z(n8520) );
  OR U9599 ( .A(n8518), .B(n8517), .Z(n8519) );
  AND U9600 ( .A(n8520), .B(n8519), .Z(n8526) );
  XOR U9601 ( .A(n8527), .B(n8526), .Z(n8529) );
  XOR U9602 ( .A(n8528), .B(n8529), .Z(n8542) );
  XNOR U9603 ( .A(n8542), .B(sreg[1319]), .Z(n8544) );
  NANDN U9604 ( .A(n8521), .B(sreg[1318]), .Z(n8525) );
  NAND U9605 ( .A(n8523), .B(n8522), .Z(n8524) );
  NAND U9606 ( .A(n8525), .B(n8524), .Z(n8543) );
  XOR U9607 ( .A(n8544), .B(n8543), .Z(c[1319]) );
  NANDN U9608 ( .A(n8527), .B(n8526), .Z(n8531) );
  OR U9609 ( .A(n8529), .B(n8528), .Z(n8530) );
  AND U9610 ( .A(n8531), .B(n8530), .Z(n8549) );
  XOR U9611 ( .A(a[298]), .B(n2218), .Z(n8553) );
  AND U9612 ( .A(a[300]), .B(b[0]), .Z(n8533) );
  XNOR U9613 ( .A(n8533), .B(n2175), .Z(n8535) );
  NANDN U9614 ( .A(b[0]), .B(a[299]), .Z(n8534) );
  NAND U9615 ( .A(n8535), .B(n8534), .Z(n8558) );
  AND U9616 ( .A(a[296]), .B(b[3]), .Z(n8557) );
  XOR U9617 ( .A(n8558), .B(n8557), .Z(n8560) );
  XOR U9618 ( .A(n8559), .B(n8560), .Z(n8548) );
  NANDN U9619 ( .A(n8537), .B(n8536), .Z(n8541) );
  OR U9620 ( .A(n8539), .B(n8538), .Z(n8540) );
  AND U9621 ( .A(n8541), .B(n8540), .Z(n8547) );
  XOR U9622 ( .A(n8548), .B(n8547), .Z(n8550) );
  XOR U9623 ( .A(n8549), .B(n8550), .Z(n8563) );
  XNOR U9624 ( .A(n8563), .B(sreg[1320]), .Z(n8565) );
  NANDN U9625 ( .A(n8542), .B(sreg[1319]), .Z(n8546) );
  NAND U9626 ( .A(n8544), .B(n8543), .Z(n8545) );
  NAND U9627 ( .A(n8546), .B(n8545), .Z(n8564) );
  XOR U9628 ( .A(n8565), .B(n8564), .Z(c[1320]) );
  NANDN U9629 ( .A(n8548), .B(n8547), .Z(n8552) );
  OR U9630 ( .A(n8550), .B(n8549), .Z(n8551) );
  AND U9631 ( .A(n8552), .B(n8551), .Z(n8570) );
  XOR U9632 ( .A(a[299]), .B(n2218), .Z(n8574) );
  AND U9633 ( .A(a[301]), .B(b[0]), .Z(n8554) );
  XNOR U9634 ( .A(n8554), .B(n2175), .Z(n8556) );
  NANDN U9635 ( .A(b[0]), .B(a[300]), .Z(n8555) );
  NAND U9636 ( .A(n8556), .B(n8555), .Z(n8579) );
  AND U9637 ( .A(a[297]), .B(b[3]), .Z(n8578) );
  XOR U9638 ( .A(n8579), .B(n8578), .Z(n8581) );
  XOR U9639 ( .A(n8580), .B(n8581), .Z(n8569) );
  NANDN U9640 ( .A(n8558), .B(n8557), .Z(n8562) );
  OR U9641 ( .A(n8560), .B(n8559), .Z(n8561) );
  AND U9642 ( .A(n8562), .B(n8561), .Z(n8568) );
  XOR U9643 ( .A(n8569), .B(n8568), .Z(n8571) );
  XOR U9644 ( .A(n8570), .B(n8571), .Z(n8584) );
  XNOR U9645 ( .A(n8584), .B(sreg[1321]), .Z(n8586) );
  NANDN U9646 ( .A(n8563), .B(sreg[1320]), .Z(n8567) );
  NAND U9647 ( .A(n8565), .B(n8564), .Z(n8566) );
  NAND U9648 ( .A(n8567), .B(n8566), .Z(n8585) );
  XOR U9649 ( .A(n8586), .B(n8585), .Z(c[1321]) );
  NANDN U9650 ( .A(n8569), .B(n8568), .Z(n8573) );
  OR U9651 ( .A(n8571), .B(n8570), .Z(n8572) );
  AND U9652 ( .A(n8573), .B(n8572), .Z(n8591) );
  XOR U9653 ( .A(a[300]), .B(n2219), .Z(n8595) );
  AND U9654 ( .A(a[302]), .B(b[0]), .Z(n8575) );
  XNOR U9655 ( .A(n8575), .B(n2175), .Z(n8577) );
  NANDN U9656 ( .A(b[0]), .B(a[301]), .Z(n8576) );
  NAND U9657 ( .A(n8577), .B(n8576), .Z(n8600) );
  AND U9658 ( .A(a[298]), .B(b[3]), .Z(n8599) );
  XOR U9659 ( .A(n8600), .B(n8599), .Z(n8602) );
  XOR U9660 ( .A(n8601), .B(n8602), .Z(n8590) );
  NANDN U9661 ( .A(n8579), .B(n8578), .Z(n8583) );
  OR U9662 ( .A(n8581), .B(n8580), .Z(n8582) );
  AND U9663 ( .A(n8583), .B(n8582), .Z(n8589) );
  XOR U9664 ( .A(n8590), .B(n8589), .Z(n8592) );
  XOR U9665 ( .A(n8591), .B(n8592), .Z(n8605) );
  XNOR U9666 ( .A(n8605), .B(sreg[1322]), .Z(n8607) );
  NANDN U9667 ( .A(n8584), .B(sreg[1321]), .Z(n8588) );
  NAND U9668 ( .A(n8586), .B(n8585), .Z(n8587) );
  NAND U9669 ( .A(n8588), .B(n8587), .Z(n8606) );
  XOR U9670 ( .A(n8607), .B(n8606), .Z(c[1322]) );
  NANDN U9671 ( .A(n8590), .B(n8589), .Z(n8594) );
  OR U9672 ( .A(n8592), .B(n8591), .Z(n8593) );
  AND U9673 ( .A(n8594), .B(n8593), .Z(n8612) );
  XOR U9674 ( .A(a[301]), .B(n2219), .Z(n8616) );
  AND U9675 ( .A(a[303]), .B(b[0]), .Z(n8596) );
  XNOR U9676 ( .A(n8596), .B(n2175), .Z(n8598) );
  NANDN U9677 ( .A(b[0]), .B(a[302]), .Z(n8597) );
  NAND U9678 ( .A(n8598), .B(n8597), .Z(n8621) );
  AND U9679 ( .A(a[299]), .B(b[3]), .Z(n8620) );
  XOR U9680 ( .A(n8621), .B(n8620), .Z(n8623) );
  XOR U9681 ( .A(n8622), .B(n8623), .Z(n8611) );
  NANDN U9682 ( .A(n8600), .B(n8599), .Z(n8604) );
  OR U9683 ( .A(n8602), .B(n8601), .Z(n8603) );
  AND U9684 ( .A(n8604), .B(n8603), .Z(n8610) );
  XOR U9685 ( .A(n8611), .B(n8610), .Z(n8613) );
  XOR U9686 ( .A(n8612), .B(n8613), .Z(n8626) );
  XNOR U9687 ( .A(n8626), .B(sreg[1323]), .Z(n8628) );
  NANDN U9688 ( .A(n8605), .B(sreg[1322]), .Z(n8609) );
  NAND U9689 ( .A(n8607), .B(n8606), .Z(n8608) );
  NAND U9690 ( .A(n8609), .B(n8608), .Z(n8627) );
  XOR U9691 ( .A(n8628), .B(n8627), .Z(c[1323]) );
  NANDN U9692 ( .A(n8611), .B(n8610), .Z(n8615) );
  OR U9693 ( .A(n8613), .B(n8612), .Z(n8614) );
  AND U9694 ( .A(n8615), .B(n8614), .Z(n8633) );
  XOR U9695 ( .A(a[302]), .B(n2219), .Z(n8637) );
  AND U9696 ( .A(a[304]), .B(b[0]), .Z(n8617) );
  XNOR U9697 ( .A(n8617), .B(n2175), .Z(n8619) );
  NANDN U9698 ( .A(b[0]), .B(a[303]), .Z(n8618) );
  NAND U9699 ( .A(n8619), .B(n8618), .Z(n8642) );
  AND U9700 ( .A(a[300]), .B(b[3]), .Z(n8641) );
  XOR U9701 ( .A(n8642), .B(n8641), .Z(n8644) );
  XOR U9702 ( .A(n8643), .B(n8644), .Z(n8632) );
  NANDN U9703 ( .A(n8621), .B(n8620), .Z(n8625) );
  OR U9704 ( .A(n8623), .B(n8622), .Z(n8624) );
  AND U9705 ( .A(n8625), .B(n8624), .Z(n8631) );
  XOR U9706 ( .A(n8632), .B(n8631), .Z(n8634) );
  XOR U9707 ( .A(n8633), .B(n8634), .Z(n8647) );
  XNOR U9708 ( .A(n8647), .B(sreg[1324]), .Z(n8649) );
  NANDN U9709 ( .A(n8626), .B(sreg[1323]), .Z(n8630) );
  NAND U9710 ( .A(n8628), .B(n8627), .Z(n8629) );
  NAND U9711 ( .A(n8630), .B(n8629), .Z(n8648) );
  XOR U9712 ( .A(n8649), .B(n8648), .Z(c[1324]) );
  NANDN U9713 ( .A(n8632), .B(n8631), .Z(n8636) );
  OR U9714 ( .A(n8634), .B(n8633), .Z(n8635) );
  AND U9715 ( .A(n8636), .B(n8635), .Z(n8654) );
  XOR U9716 ( .A(a[303]), .B(n2219), .Z(n8658) );
  AND U9717 ( .A(a[301]), .B(b[3]), .Z(n8662) );
  AND U9718 ( .A(a[305]), .B(b[0]), .Z(n8638) );
  XNOR U9719 ( .A(n8638), .B(n2175), .Z(n8640) );
  NANDN U9720 ( .A(b[0]), .B(a[304]), .Z(n8639) );
  NAND U9721 ( .A(n8640), .B(n8639), .Z(n8663) );
  XOR U9722 ( .A(n8662), .B(n8663), .Z(n8665) );
  XOR U9723 ( .A(n8664), .B(n8665), .Z(n8653) );
  NANDN U9724 ( .A(n8642), .B(n8641), .Z(n8646) );
  OR U9725 ( .A(n8644), .B(n8643), .Z(n8645) );
  AND U9726 ( .A(n8646), .B(n8645), .Z(n8652) );
  XOR U9727 ( .A(n8653), .B(n8652), .Z(n8655) );
  XOR U9728 ( .A(n8654), .B(n8655), .Z(n8668) );
  XNOR U9729 ( .A(n8668), .B(sreg[1325]), .Z(n8670) );
  NANDN U9730 ( .A(n8647), .B(sreg[1324]), .Z(n8651) );
  NAND U9731 ( .A(n8649), .B(n8648), .Z(n8650) );
  NAND U9732 ( .A(n8651), .B(n8650), .Z(n8669) );
  XOR U9733 ( .A(n8670), .B(n8669), .Z(c[1325]) );
  NANDN U9734 ( .A(n8653), .B(n8652), .Z(n8657) );
  OR U9735 ( .A(n8655), .B(n8654), .Z(n8656) );
  AND U9736 ( .A(n8657), .B(n8656), .Z(n8675) );
  XOR U9737 ( .A(a[304]), .B(n2219), .Z(n8679) );
  AND U9738 ( .A(a[306]), .B(b[0]), .Z(n8659) );
  XNOR U9739 ( .A(n8659), .B(n2175), .Z(n8661) );
  NANDN U9740 ( .A(b[0]), .B(a[305]), .Z(n8660) );
  NAND U9741 ( .A(n8661), .B(n8660), .Z(n8684) );
  AND U9742 ( .A(a[302]), .B(b[3]), .Z(n8683) );
  XOR U9743 ( .A(n8684), .B(n8683), .Z(n8686) );
  XOR U9744 ( .A(n8685), .B(n8686), .Z(n8674) );
  NANDN U9745 ( .A(n8663), .B(n8662), .Z(n8667) );
  OR U9746 ( .A(n8665), .B(n8664), .Z(n8666) );
  AND U9747 ( .A(n8667), .B(n8666), .Z(n8673) );
  XOR U9748 ( .A(n8674), .B(n8673), .Z(n8676) );
  XOR U9749 ( .A(n8675), .B(n8676), .Z(n8689) );
  XNOR U9750 ( .A(n8689), .B(sreg[1326]), .Z(n8691) );
  NANDN U9751 ( .A(n8668), .B(sreg[1325]), .Z(n8672) );
  NAND U9752 ( .A(n8670), .B(n8669), .Z(n8671) );
  NAND U9753 ( .A(n8672), .B(n8671), .Z(n8690) );
  XOR U9754 ( .A(n8691), .B(n8690), .Z(c[1326]) );
  NANDN U9755 ( .A(n8674), .B(n8673), .Z(n8678) );
  OR U9756 ( .A(n8676), .B(n8675), .Z(n8677) );
  AND U9757 ( .A(n8678), .B(n8677), .Z(n8696) );
  XOR U9758 ( .A(a[305]), .B(n2219), .Z(n8700) );
  AND U9759 ( .A(a[303]), .B(b[3]), .Z(n8704) );
  AND U9760 ( .A(a[307]), .B(b[0]), .Z(n8680) );
  XNOR U9761 ( .A(n8680), .B(n2175), .Z(n8682) );
  NANDN U9762 ( .A(b[0]), .B(a[306]), .Z(n8681) );
  NAND U9763 ( .A(n8682), .B(n8681), .Z(n8705) );
  XOR U9764 ( .A(n8704), .B(n8705), .Z(n8707) );
  XOR U9765 ( .A(n8706), .B(n8707), .Z(n8695) );
  NANDN U9766 ( .A(n8684), .B(n8683), .Z(n8688) );
  OR U9767 ( .A(n8686), .B(n8685), .Z(n8687) );
  AND U9768 ( .A(n8688), .B(n8687), .Z(n8694) );
  XOR U9769 ( .A(n8695), .B(n8694), .Z(n8697) );
  XOR U9770 ( .A(n8696), .B(n8697), .Z(n8710) );
  XNOR U9771 ( .A(n8710), .B(sreg[1327]), .Z(n8712) );
  NANDN U9772 ( .A(n8689), .B(sreg[1326]), .Z(n8693) );
  NAND U9773 ( .A(n8691), .B(n8690), .Z(n8692) );
  NAND U9774 ( .A(n8693), .B(n8692), .Z(n8711) );
  XOR U9775 ( .A(n8712), .B(n8711), .Z(c[1327]) );
  NANDN U9776 ( .A(n8695), .B(n8694), .Z(n8699) );
  OR U9777 ( .A(n8697), .B(n8696), .Z(n8698) );
  AND U9778 ( .A(n8699), .B(n8698), .Z(n8717) );
  XOR U9779 ( .A(a[306]), .B(n2219), .Z(n8721) );
  AND U9780 ( .A(a[308]), .B(b[0]), .Z(n8701) );
  XNOR U9781 ( .A(n8701), .B(n2175), .Z(n8703) );
  NANDN U9782 ( .A(b[0]), .B(a[307]), .Z(n8702) );
  NAND U9783 ( .A(n8703), .B(n8702), .Z(n8726) );
  AND U9784 ( .A(a[304]), .B(b[3]), .Z(n8725) );
  XOR U9785 ( .A(n8726), .B(n8725), .Z(n8728) );
  XOR U9786 ( .A(n8727), .B(n8728), .Z(n8716) );
  NANDN U9787 ( .A(n8705), .B(n8704), .Z(n8709) );
  OR U9788 ( .A(n8707), .B(n8706), .Z(n8708) );
  AND U9789 ( .A(n8709), .B(n8708), .Z(n8715) );
  XOR U9790 ( .A(n8716), .B(n8715), .Z(n8718) );
  XOR U9791 ( .A(n8717), .B(n8718), .Z(n8731) );
  XNOR U9792 ( .A(n8731), .B(sreg[1328]), .Z(n8733) );
  NANDN U9793 ( .A(n8710), .B(sreg[1327]), .Z(n8714) );
  NAND U9794 ( .A(n8712), .B(n8711), .Z(n8713) );
  NAND U9795 ( .A(n8714), .B(n8713), .Z(n8732) );
  XOR U9796 ( .A(n8733), .B(n8732), .Z(c[1328]) );
  NANDN U9797 ( .A(n8716), .B(n8715), .Z(n8720) );
  OR U9798 ( .A(n8718), .B(n8717), .Z(n8719) );
  AND U9799 ( .A(n8720), .B(n8719), .Z(n8738) );
  XOR U9800 ( .A(a[307]), .B(n2220), .Z(n8742) );
  AND U9801 ( .A(a[309]), .B(b[0]), .Z(n8722) );
  XNOR U9802 ( .A(n8722), .B(n2175), .Z(n8724) );
  NANDN U9803 ( .A(b[0]), .B(a[308]), .Z(n8723) );
  NAND U9804 ( .A(n8724), .B(n8723), .Z(n8747) );
  AND U9805 ( .A(a[305]), .B(b[3]), .Z(n8746) );
  XOR U9806 ( .A(n8747), .B(n8746), .Z(n8749) );
  XOR U9807 ( .A(n8748), .B(n8749), .Z(n8737) );
  NANDN U9808 ( .A(n8726), .B(n8725), .Z(n8730) );
  OR U9809 ( .A(n8728), .B(n8727), .Z(n8729) );
  AND U9810 ( .A(n8730), .B(n8729), .Z(n8736) );
  XOR U9811 ( .A(n8737), .B(n8736), .Z(n8739) );
  XOR U9812 ( .A(n8738), .B(n8739), .Z(n8752) );
  XNOR U9813 ( .A(n8752), .B(sreg[1329]), .Z(n8754) );
  NANDN U9814 ( .A(n8731), .B(sreg[1328]), .Z(n8735) );
  NAND U9815 ( .A(n8733), .B(n8732), .Z(n8734) );
  NAND U9816 ( .A(n8735), .B(n8734), .Z(n8753) );
  XOR U9817 ( .A(n8754), .B(n8753), .Z(c[1329]) );
  NANDN U9818 ( .A(n8737), .B(n8736), .Z(n8741) );
  OR U9819 ( .A(n8739), .B(n8738), .Z(n8740) );
  AND U9820 ( .A(n8741), .B(n8740), .Z(n8759) );
  XOR U9821 ( .A(a[308]), .B(n2220), .Z(n8763) );
  AND U9822 ( .A(a[310]), .B(b[0]), .Z(n8743) );
  XNOR U9823 ( .A(n8743), .B(n2175), .Z(n8745) );
  NANDN U9824 ( .A(b[0]), .B(a[309]), .Z(n8744) );
  NAND U9825 ( .A(n8745), .B(n8744), .Z(n8768) );
  AND U9826 ( .A(a[306]), .B(b[3]), .Z(n8767) );
  XOR U9827 ( .A(n8768), .B(n8767), .Z(n8770) );
  XOR U9828 ( .A(n8769), .B(n8770), .Z(n8758) );
  NANDN U9829 ( .A(n8747), .B(n8746), .Z(n8751) );
  OR U9830 ( .A(n8749), .B(n8748), .Z(n8750) );
  AND U9831 ( .A(n8751), .B(n8750), .Z(n8757) );
  XOR U9832 ( .A(n8758), .B(n8757), .Z(n8760) );
  XOR U9833 ( .A(n8759), .B(n8760), .Z(n8773) );
  XNOR U9834 ( .A(n8773), .B(sreg[1330]), .Z(n8775) );
  NANDN U9835 ( .A(n8752), .B(sreg[1329]), .Z(n8756) );
  NAND U9836 ( .A(n8754), .B(n8753), .Z(n8755) );
  NAND U9837 ( .A(n8756), .B(n8755), .Z(n8774) );
  XOR U9838 ( .A(n8775), .B(n8774), .Z(c[1330]) );
  NANDN U9839 ( .A(n8758), .B(n8757), .Z(n8762) );
  OR U9840 ( .A(n8760), .B(n8759), .Z(n8761) );
  AND U9841 ( .A(n8762), .B(n8761), .Z(n8780) );
  XOR U9842 ( .A(a[309]), .B(n2220), .Z(n8784) );
  AND U9843 ( .A(a[307]), .B(b[3]), .Z(n8788) );
  AND U9844 ( .A(a[311]), .B(b[0]), .Z(n8764) );
  XNOR U9845 ( .A(n8764), .B(n2175), .Z(n8766) );
  NANDN U9846 ( .A(b[0]), .B(a[310]), .Z(n8765) );
  NAND U9847 ( .A(n8766), .B(n8765), .Z(n8789) );
  XOR U9848 ( .A(n8788), .B(n8789), .Z(n8791) );
  XOR U9849 ( .A(n8790), .B(n8791), .Z(n8779) );
  NANDN U9850 ( .A(n8768), .B(n8767), .Z(n8772) );
  OR U9851 ( .A(n8770), .B(n8769), .Z(n8771) );
  AND U9852 ( .A(n8772), .B(n8771), .Z(n8778) );
  XOR U9853 ( .A(n8779), .B(n8778), .Z(n8781) );
  XOR U9854 ( .A(n8780), .B(n8781), .Z(n8794) );
  XNOR U9855 ( .A(n8794), .B(sreg[1331]), .Z(n8796) );
  NANDN U9856 ( .A(n8773), .B(sreg[1330]), .Z(n8777) );
  NAND U9857 ( .A(n8775), .B(n8774), .Z(n8776) );
  NAND U9858 ( .A(n8777), .B(n8776), .Z(n8795) );
  XOR U9859 ( .A(n8796), .B(n8795), .Z(c[1331]) );
  NANDN U9860 ( .A(n8779), .B(n8778), .Z(n8783) );
  OR U9861 ( .A(n8781), .B(n8780), .Z(n8782) );
  AND U9862 ( .A(n8783), .B(n8782), .Z(n8801) );
  XOR U9863 ( .A(a[310]), .B(n2220), .Z(n8805) );
  AND U9864 ( .A(a[312]), .B(b[0]), .Z(n8785) );
  XNOR U9865 ( .A(n8785), .B(n2175), .Z(n8787) );
  NANDN U9866 ( .A(b[0]), .B(a[311]), .Z(n8786) );
  NAND U9867 ( .A(n8787), .B(n8786), .Z(n8810) );
  AND U9868 ( .A(a[308]), .B(b[3]), .Z(n8809) );
  XOR U9869 ( .A(n8810), .B(n8809), .Z(n8812) );
  XOR U9870 ( .A(n8811), .B(n8812), .Z(n8800) );
  NANDN U9871 ( .A(n8789), .B(n8788), .Z(n8793) );
  OR U9872 ( .A(n8791), .B(n8790), .Z(n8792) );
  AND U9873 ( .A(n8793), .B(n8792), .Z(n8799) );
  XOR U9874 ( .A(n8800), .B(n8799), .Z(n8802) );
  XOR U9875 ( .A(n8801), .B(n8802), .Z(n8815) );
  XNOR U9876 ( .A(n8815), .B(sreg[1332]), .Z(n8817) );
  NANDN U9877 ( .A(n8794), .B(sreg[1331]), .Z(n8798) );
  NAND U9878 ( .A(n8796), .B(n8795), .Z(n8797) );
  NAND U9879 ( .A(n8798), .B(n8797), .Z(n8816) );
  XOR U9880 ( .A(n8817), .B(n8816), .Z(c[1332]) );
  NANDN U9881 ( .A(n8800), .B(n8799), .Z(n8804) );
  OR U9882 ( .A(n8802), .B(n8801), .Z(n8803) );
  AND U9883 ( .A(n8804), .B(n8803), .Z(n8822) );
  XOR U9884 ( .A(a[311]), .B(n2220), .Z(n8826) );
  AND U9885 ( .A(a[309]), .B(b[3]), .Z(n8830) );
  AND U9886 ( .A(a[313]), .B(b[0]), .Z(n8806) );
  XNOR U9887 ( .A(n8806), .B(n2175), .Z(n8808) );
  NANDN U9888 ( .A(b[0]), .B(a[312]), .Z(n8807) );
  NAND U9889 ( .A(n8808), .B(n8807), .Z(n8831) );
  XOR U9890 ( .A(n8830), .B(n8831), .Z(n8833) );
  XOR U9891 ( .A(n8832), .B(n8833), .Z(n8821) );
  NANDN U9892 ( .A(n8810), .B(n8809), .Z(n8814) );
  OR U9893 ( .A(n8812), .B(n8811), .Z(n8813) );
  AND U9894 ( .A(n8814), .B(n8813), .Z(n8820) );
  XOR U9895 ( .A(n8821), .B(n8820), .Z(n8823) );
  XOR U9896 ( .A(n8822), .B(n8823), .Z(n8836) );
  XNOR U9897 ( .A(n8836), .B(sreg[1333]), .Z(n8838) );
  NANDN U9898 ( .A(n8815), .B(sreg[1332]), .Z(n8819) );
  NAND U9899 ( .A(n8817), .B(n8816), .Z(n8818) );
  NAND U9900 ( .A(n8819), .B(n8818), .Z(n8837) );
  XOR U9901 ( .A(n8838), .B(n8837), .Z(c[1333]) );
  NANDN U9902 ( .A(n8821), .B(n8820), .Z(n8825) );
  OR U9903 ( .A(n8823), .B(n8822), .Z(n8824) );
  AND U9904 ( .A(n8825), .B(n8824), .Z(n8843) );
  XOR U9905 ( .A(a[312]), .B(n2220), .Z(n8847) );
  AND U9906 ( .A(a[314]), .B(b[0]), .Z(n8827) );
  XNOR U9907 ( .A(n8827), .B(n2175), .Z(n8829) );
  NANDN U9908 ( .A(b[0]), .B(a[313]), .Z(n8828) );
  NAND U9909 ( .A(n8829), .B(n8828), .Z(n8852) );
  AND U9910 ( .A(a[310]), .B(b[3]), .Z(n8851) );
  XOR U9911 ( .A(n8852), .B(n8851), .Z(n8854) );
  XOR U9912 ( .A(n8853), .B(n8854), .Z(n8842) );
  NANDN U9913 ( .A(n8831), .B(n8830), .Z(n8835) );
  OR U9914 ( .A(n8833), .B(n8832), .Z(n8834) );
  AND U9915 ( .A(n8835), .B(n8834), .Z(n8841) );
  XOR U9916 ( .A(n8842), .B(n8841), .Z(n8844) );
  XOR U9917 ( .A(n8843), .B(n8844), .Z(n8857) );
  XNOR U9918 ( .A(n8857), .B(sreg[1334]), .Z(n8859) );
  NANDN U9919 ( .A(n8836), .B(sreg[1333]), .Z(n8840) );
  NAND U9920 ( .A(n8838), .B(n8837), .Z(n8839) );
  NAND U9921 ( .A(n8840), .B(n8839), .Z(n8858) );
  XOR U9922 ( .A(n8859), .B(n8858), .Z(c[1334]) );
  NANDN U9923 ( .A(n8842), .B(n8841), .Z(n8846) );
  OR U9924 ( .A(n8844), .B(n8843), .Z(n8845) );
  AND U9925 ( .A(n8846), .B(n8845), .Z(n8864) );
  XOR U9926 ( .A(a[313]), .B(n2220), .Z(n8868) );
  AND U9927 ( .A(a[311]), .B(b[3]), .Z(n8872) );
  AND U9928 ( .A(a[315]), .B(b[0]), .Z(n8848) );
  XNOR U9929 ( .A(n8848), .B(n2175), .Z(n8850) );
  NANDN U9930 ( .A(b[0]), .B(a[314]), .Z(n8849) );
  NAND U9931 ( .A(n8850), .B(n8849), .Z(n8873) );
  XOR U9932 ( .A(n8872), .B(n8873), .Z(n8875) );
  XOR U9933 ( .A(n8874), .B(n8875), .Z(n8863) );
  NANDN U9934 ( .A(n8852), .B(n8851), .Z(n8856) );
  OR U9935 ( .A(n8854), .B(n8853), .Z(n8855) );
  AND U9936 ( .A(n8856), .B(n8855), .Z(n8862) );
  XOR U9937 ( .A(n8863), .B(n8862), .Z(n8865) );
  XOR U9938 ( .A(n8864), .B(n8865), .Z(n8878) );
  XNOR U9939 ( .A(n8878), .B(sreg[1335]), .Z(n8880) );
  NANDN U9940 ( .A(n8857), .B(sreg[1334]), .Z(n8861) );
  NAND U9941 ( .A(n8859), .B(n8858), .Z(n8860) );
  NAND U9942 ( .A(n8861), .B(n8860), .Z(n8879) );
  XOR U9943 ( .A(n8880), .B(n8879), .Z(c[1335]) );
  NANDN U9944 ( .A(n8863), .B(n8862), .Z(n8867) );
  OR U9945 ( .A(n8865), .B(n8864), .Z(n8866) );
  AND U9946 ( .A(n8867), .B(n8866), .Z(n8885) );
  XOR U9947 ( .A(a[314]), .B(n2221), .Z(n8889) );
  AND U9948 ( .A(a[312]), .B(b[3]), .Z(n8893) );
  AND U9949 ( .A(a[316]), .B(b[0]), .Z(n8869) );
  XNOR U9950 ( .A(n8869), .B(n2175), .Z(n8871) );
  NANDN U9951 ( .A(b[0]), .B(a[315]), .Z(n8870) );
  NAND U9952 ( .A(n8871), .B(n8870), .Z(n8894) );
  XOR U9953 ( .A(n8893), .B(n8894), .Z(n8896) );
  XOR U9954 ( .A(n8895), .B(n8896), .Z(n8884) );
  NANDN U9955 ( .A(n8873), .B(n8872), .Z(n8877) );
  OR U9956 ( .A(n8875), .B(n8874), .Z(n8876) );
  AND U9957 ( .A(n8877), .B(n8876), .Z(n8883) );
  XOR U9958 ( .A(n8884), .B(n8883), .Z(n8886) );
  XOR U9959 ( .A(n8885), .B(n8886), .Z(n8899) );
  XNOR U9960 ( .A(n8899), .B(sreg[1336]), .Z(n8901) );
  NANDN U9961 ( .A(n8878), .B(sreg[1335]), .Z(n8882) );
  NAND U9962 ( .A(n8880), .B(n8879), .Z(n8881) );
  NAND U9963 ( .A(n8882), .B(n8881), .Z(n8900) );
  XOR U9964 ( .A(n8901), .B(n8900), .Z(c[1336]) );
  NANDN U9965 ( .A(n8884), .B(n8883), .Z(n8888) );
  OR U9966 ( .A(n8886), .B(n8885), .Z(n8887) );
  AND U9967 ( .A(n8888), .B(n8887), .Z(n8906) );
  XOR U9968 ( .A(a[315]), .B(n2221), .Z(n8910) );
  AND U9969 ( .A(a[317]), .B(b[0]), .Z(n8890) );
  XNOR U9970 ( .A(n8890), .B(n2175), .Z(n8892) );
  NANDN U9971 ( .A(b[0]), .B(a[316]), .Z(n8891) );
  NAND U9972 ( .A(n8892), .B(n8891), .Z(n8915) );
  AND U9973 ( .A(a[313]), .B(b[3]), .Z(n8914) );
  XOR U9974 ( .A(n8915), .B(n8914), .Z(n8917) );
  XOR U9975 ( .A(n8916), .B(n8917), .Z(n8905) );
  NANDN U9976 ( .A(n8894), .B(n8893), .Z(n8898) );
  OR U9977 ( .A(n8896), .B(n8895), .Z(n8897) );
  AND U9978 ( .A(n8898), .B(n8897), .Z(n8904) );
  XOR U9979 ( .A(n8905), .B(n8904), .Z(n8907) );
  XOR U9980 ( .A(n8906), .B(n8907), .Z(n8920) );
  XNOR U9981 ( .A(n8920), .B(sreg[1337]), .Z(n8922) );
  NANDN U9982 ( .A(n8899), .B(sreg[1336]), .Z(n8903) );
  NAND U9983 ( .A(n8901), .B(n8900), .Z(n8902) );
  NAND U9984 ( .A(n8903), .B(n8902), .Z(n8921) );
  XOR U9985 ( .A(n8922), .B(n8921), .Z(c[1337]) );
  NANDN U9986 ( .A(n8905), .B(n8904), .Z(n8909) );
  OR U9987 ( .A(n8907), .B(n8906), .Z(n8908) );
  AND U9988 ( .A(n8909), .B(n8908), .Z(n8927) );
  XOR U9989 ( .A(a[316]), .B(n2221), .Z(n8931) );
  AND U9990 ( .A(a[318]), .B(b[0]), .Z(n8911) );
  XNOR U9991 ( .A(n8911), .B(n2175), .Z(n8913) );
  NANDN U9992 ( .A(b[0]), .B(a[317]), .Z(n8912) );
  NAND U9993 ( .A(n8913), .B(n8912), .Z(n8936) );
  AND U9994 ( .A(a[314]), .B(b[3]), .Z(n8935) );
  XOR U9995 ( .A(n8936), .B(n8935), .Z(n8938) );
  XOR U9996 ( .A(n8937), .B(n8938), .Z(n8926) );
  NANDN U9997 ( .A(n8915), .B(n8914), .Z(n8919) );
  OR U9998 ( .A(n8917), .B(n8916), .Z(n8918) );
  AND U9999 ( .A(n8919), .B(n8918), .Z(n8925) );
  XOR U10000 ( .A(n8926), .B(n8925), .Z(n8928) );
  XOR U10001 ( .A(n8927), .B(n8928), .Z(n8941) );
  XNOR U10002 ( .A(n8941), .B(sreg[1338]), .Z(n8943) );
  NANDN U10003 ( .A(n8920), .B(sreg[1337]), .Z(n8924) );
  NAND U10004 ( .A(n8922), .B(n8921), .Z(n8923) );
  NAND U10005 ( .A(n8924), .B(n8923), .Z(n8942) );
  XOR U10006 ( .A(n8943), .B(n8942), .Z(c[1338]) );
  NANDN U10007 ( .A(n8926), .B(n8925), .Z(n8930) );
  OR U10008 ( .A(n8928), .B(n8927), .Z(n8929) );
  AND U10009 ( .A(n8930), .B(n8929), .Z(n8948) );
  XOR U10010 ( .A(a[317]), .B(n2221), .Z(n8952) );
  AND U10011 ( .A(a[315]), .B(b[3]), .Z(n8956) );
  AND U10012 ( .A(a[319]), .B(b[0]), .Z(n8932) );
  XNOR U10013 ( .A(n8932), .B(n2175), .Z(n8934) );
  NANDN U10014 ( .A(b[0]), .B(a[318]), .Z(n8933) );
  NAND U10015 ( .A(n8934), .B(n8933), .Z(n8957) );
  XOR U10016 ( .A(n8956), .B(n8957), .Z(n8959) );
  XOR U10017 ( .A(n8958), .B(n8959), .Z(n8947) );
  NANDN U10018 ( .A(n8936), .B(n8935), .Z(n8940) );
  OR U10019 ( .A(n8938), .B(n8937), .Z(n8939) );
  AND U10020 ( .A(n8940), .B(n8939), .Z(n8946) );
  XOR U10021 ( .A(n8947), .B(n8946), .Z(n8949) );
  XOR U10022 ( .A(n8948), .B(n8949), .Z(n8962) );
  XNOR U10023 ( .A(n8962), .B(sreg[1339]), .Z(n8964) );
  NANDN U10024 ( .A(n8941), .B(sreg[1338]), .Z(n8945) );
  NAND U10025 ( .A(n8943), .B(n8942), .Z(n8944) );
  NAND U10026 ( .A(n8945), .B(n8944), .Z(n8963) );
  XOR U10027 ( .A(n8964), .B(n8963), .Z(c[1339]) );
  NANDN U10028 ( .A(n8947), .B(n8946), .Z(n8951) );
  OR U10029 ( .A(n8949), .B(n8948), .Z(n8950) );
  AND U10030 ( .A(n8951), .B(n8950), .Z(n8969) );
  XOR U10031 ( .A(a[318]), .B(n2221), .Z(n8973) );
  AND U10032 ( .A(a[320]), .B(b[0]), .Z(n8953) );
  XNOR U10033 ( .A(n8953), .B(n2175), .Z(n8955) );
  NANDN U10034 ( .A(b[0]), .B(a[319]), .Z(n8954) );
  NAND U10035 ( .A(n8955), .B(n8954), .Z(n8978) );
  AND U10036 ( .A(a[316]), .B(b[3]), .Z(n8977) );
  XOR U10037 ( .A(n8978), .B(n8977), .Z(n8980) );
  XOR U10038 ( .A(n8979), .B(n8980), .Z(n8968) );
  NANDN U10039 ( .A(n8957), .B(n8956), .Z(n8961) );
  OR U10040 ( .A(n8959), .B(n8958), .Z(n8960) );
  AND U10041 ( .A(n8961), .B(n8960), .Z(n8967) );
  XOR U10042 ( .A(n8968), .B(n8967), .Z(n8970) );
  XOR U10043 ( .A(n8969), .B(n8970), .Z(n8983) );
  XNOR U10044 ( .A(n8983), .B(sreg[1340]), .Z(n8985) );
  NANDN U10045 ( .A(n8962), .B(sreg[1339]), .Z(n8966) );
  NAND U10046 ( .A(n8964), .B(n8963), .Z(n8965) );
  NAND U10047 ( .A(n8966), .B(n8965), .Z(n8984) );
  XOR U10048 ( .A(n8985), .B(n8984), .Z(c[1340]) );
  NANDN U10049 ( .A(n8968), .B(n8967), .Z(n8972) );
  OR U10050 ( .A(n8970), .B(n8969), .Z(n8971) );
  AND U10051 ( .A(n8972), .B(n8971), .Z(n8990) );
  XOR U10052 ( .A(a[319]), .B(n2221), .Z(n8994) );
  AND U10053 ( .A(a[321]), .B(b[0]), .Z(n8974) );
  XNOR U10054 ( .A(n8974), .B(n2175), .Z(n8976) );
  NANDN U10055 ( .A(b[0]), .B(a[320]), .Z(n8975) );
  NAND U10056 ( .A(n8976), .B(n8975), .Z(n8999) );
  AND U10057 ( .A(a[317]), .B(b[3]), .Z(n8998) );
  XOR U10058 ( .A(n8999), .B(n8998), .Z(n9001) );
  XOR U10059 ( .A(n9000), .B(n9001), .Z(n8989) );
  NANDN U10060 ( .A(n8978), .B(n8977), .Z(n8982) );
  OR U10061 ( .A(n8980), .B(n8979), .Z(n8981) );
  AND U10062 ( .A(n8982), .B(n8981), .Z(n8988) );
  XOR U10063 ( .A(n8989), .B(n8988), .Z(n8991) );
  XOR U10064 ( .A(n8990), .B(n8991), .Z(n9004) );
  XNOR U10065 ( .A(n9004), .B(sreg[1341]), .Z(n9006) );
  NANDN U10066 ( .A(n8983), .B(sreg[1340]), .Z(n8987) );
  NAND U10067 ( .A(n8985), .B(n8984), .Z(n8986) );
  NAND U10068 ( .A(n8987), .B(n8986), .Z(n9005) );
  XOR U10069 ( .A(n9006), .B(n9005), .Z(c[1341]) );
  NANDN U10070 ( .A(n8989), .B(n8988), .Z(n8993) );
  OR U10071 ( .A(n8991), .B(n8990), .Z(n8992) );
  AND U10072 ( .A(n8993), .B(n8992), .Z(n9011) );
  XOR U10073 ( .A(a[320]), .B(n2221), .Z(n9015) );
  AND U10074 ( .A(a[322]), .B(b[0]), .Z(n8995) );
  XNOR U10075 ( .A(n8995), .B(n2175), .Z(n8997) );
  NANDN U10076 ( .A(b[0]), .B(a[321]), .Z(n8996) );
  NAND U10077 ( .A(n8997), .B(n8996), .Z(n9020) );
  AND U10078 ( .A(a[318]), .B(b[3]), .Z(n9019) );
  XOR U10079 ( .A(n9020), .B(n9019), .Z(n9022) );
  XOR U10080 ( .A(n9021), .B(n9022), .Z(n9010) );
  NANDN U10081 ( .A(n8999), .B(n8998), .Z(n9003) );
  OR U10082 ( .A(n9001), .B(n9000), .Z(n9002) );
  AND U10083 ( .A(n9003), .B(n9002), .Z(n9009) );
  XOR U10084 ( .A(n9010), .B(n9009), .Z(n9012) );
  XOR U10085 ( .A(n9011), .B(n9012), .Z(n9025) );
  XNOR U10086 ( .A(n9025), .B(sreg[1342]), .Z(n9027) );
  NANDN U10087 ( .A(n9004), .B(sreg[1341]), .Z(n9008) );
  NAND U10088 ( .A(n9006), .B(n9005), .Z(n9007) );
  NAND U10089 ( .A(n9008), .B(n9007), .Z(n9026) );
  XOR U10090 ( .A(n9027), .B(n9026), .Z(c[1342]) );
  NANDN U10091 ( .A(n9010), .B(n9009), .Z(n9014) );
  OR U10092 ( .A(n9012), .B(n9011), .Z(n9013) );
  AND U10093 ( .A(n9014), .B(n9013), .Z(n9032) );
  XOR U10094 ( .A(a[321]), .B(n2222), .Z(n9036) );
  AND U10095 ( .A(a[323]), .B(b[0]), .Z(n9016) );
  XNOR U10096 ( .A(n9016), .B(n2175), .Z(n9018) );
  NANDN U10097 ( .A(b[0]), .B(a[322]), .Z(n9017) );
  NAND U10098 ( .A(n9018), .B(n9017), .Z(n9041) );
  AND U10099 ( .A(a[319]), .B(b[3]), .Z(n9040) );
  XOR U10100 ( .A(n9041), .B(n9040), .Z(n9043) );
  XOR U10101 ( .A(n9042), .B(n9043), .Z(n9031) );
  NANDN U10102 ( .A(n9020), .B(n9019), .Z(n9024) );
  OR U10103 ( .A(n9022), .B(n9021), .Z(n9023) );
  AND U10104 ( .A(n9024), .B(n9023), .Z(n9030) );
  XOR U10105 ( .A(n9031), .B(n9030), .Z(n9033) );
  XOR U10106 ( .A(n9032), .B(n9033), .Z(n9046) );
  XNOR U10107 ( .A(n9046), .B(sreg[1343]), .Z(n9048) );
  NANDN U10108 ( .A(n9025), .B(sreg[1342]), .Z(n9029) );
  NAND U10109 ( .A(n9027), .B(n9026), .Z(n9028) );
  NAND U10110 ( .A(n9029), .B(n9028), .Z(n9047) );
  XOR U10111 ( .A(n9048), .B(n9047), .Z(c[1343]) );
  NANDN U10112 ( .A(n9031), .B(n9030), .Z(n9035) );
  OR U10113 ( .A(n9033), .B(n9032), .Z(n9034) );
  AND U10114 ( .A(n9035), .B(n9034), .Z(n9054) );
  XOR U10115 ( .A(a[322]), .B(n2222), .Z(n9055) );
  AND U10116 ( .A(b[0]), .B(a[324]), .Z(n9037) );
  XOR U10117 ( .A(b[1]), .B(n9037), .Z(n9039) );
  NANDN U10118 ( .A(b[0]), .B(a[323]), .Z(n9038) );
  AND U10119 ( .A(n9039), .B(n9038), .Z(n9059) );
  AND U10120 ( .A(a[320]), .B(b[3]), .Z(n9060) );
  XOR U10121 ( .A(n9059), .B(n9060), .Z(n9061) );
  XNOR U10122 ( .A(n9062), .B(n9061), .Z(n9051) );
  NANDN U10123 ( .A(n9041), .B(n9040), .Z(n9045) );
  OR U10124 ( .A(n9043), .B(n9042), .Z(n9044) );
  AND U10125 ( .A(n9045), .B(n9044), .Z(n9052) );
  XNOR U10126 ( .A(n9051), .B(n9052), .Z(n9053) );
  XNOR U10127 ( .A(n9054), .B(n9053), .Z(n9065) );
  XNOR U10128 ( .A(n9065), .B(sreg[1344]), .Z(n9067) );
  NANDN U10129 ( .A(n9046), .B(sreg[1343]), .Z(n9050) );
  NAND U10130 ( .A(n9048), .B(n9047), .Z(n9049) );
  NAND U10131 ( .A(n9050), .B(n9049), .Z(n9066) );
  XOR U10132 ( .A(n9067), .B(n9066), .Z(c[1344]) );
  XOR U10133 ( .A(a[323]), .B(n2222), .Z(n9074) );
  AND U10134 ( .A(a[325]), .B(b[0]), .Z(n9056) );
  XNOR U10135 ( .A(n9056), .B(n2175), .Z(n9058) );
  NANDN U10136 ( .A(b[0]), .B(a[324]), .Z(n9057) );
  NAND U10137 ( .A(n9058), .B(n9057), .Z(n9079) );
  AND U10138 ( .A(a[321]), .B(b[3]), .Z(n9078) );
  XOR U10139 ( .A(n9079), .B(n9078), .Z(n9081) );
  XOR U10140 ( .A(n9080), .B(n9081), .Z(n9069) );
  NAND U10141 ( .A(n9060), .B(n9059), .Z(n9064) );
  NANDN U10142 ( .A(n9062), .B(n9061), .Z(n9063) );
  AND U10143 ( .A(n9064), .B(n9063), .Z(n9068) );
  XOR U10144 ( .A(n9069), .B(n9068), .Z(n9071) );
  XOR U10145 ( .A(n9070), .B(n9071), .Z(n9084) );
  XNOR U10146 ( .A(n9084), .B(sreg[1345]), .Z(n9086) );
  XOR U10147 ( .A(n9086), .B(n9085), .Z(c[1345]) );
  NANDN U10148 ( .A(n9069), .B(n9068), .Z(n9073) );
  OR U10149 ( .A(n9071), .B(n9070), .Z(n9072) );
  AND U10150 ( .A(n9073), .B(n9072), .Z(n9091) );
  XOR U10151 ( .A(a[324]), .B(n2222), .Z(n9095) );
  AND U10152 ( .A(a[326]), .B(b[0]), .Z(n9075) );
  XNOR U10153 ( .A(n9075), .B(n2175), .Z(n9077) );
  NANDN U10154 ( .A(b[0]), .B(a[325]), .Z(n9076) );
  NAND U10155 ( .A(n9077), .B(n9076), .Z(n9100) );
  AND U10156 ( .A(a[322]), .B(b[3]), .Z(n9099) );
  XOR U10157 ( .A(n9100), .B(n9099), .Z(n9102) );
  XOR U10158 ( .A(n9101), .B(n9102), .Z(n9090) );
  NANDN U10159 ( .A(n9079), .B(n9078), .Z(n9083) );
  OR U10160 ( .A(n9081), .B(n9080), .Z(n9082) );
  AND U10161 ( .A(n9083), .B(n9082), .Z(n9089) );
  XOR U10162 ( .A(n9090), .B(n9089), .Z(n9092) );
  XOR U10163 ( .A(n9091), .B(n9092), .Z(n9105) );
  XNOR U10164 ( .A(n9105), .B(sreg[1346]), .Z(n9107) );
  NANDN U10165 ( .A(n9084), .B(sreg[1345]), .Z(n9088) );
  NAND U10166 ( .A(n9086), .B(n9085), .Z(n9087) );
  NAND U10167 ( .A(n9088), .B(n9087), .Z(n9106) );
  XOR U10168 ( .A(n9107), .B(n9106), .Z(c[1346]) );
  NANDN U10169 ( .A(n9090), .B(n9089), .Z(n9094) );
  OR U10170 ( .A(n9092), .B(n9091), .Z(n9093) );
  AND U10171 ( .A(n9094), .B(n9093), .Z(n9112) );
  XOR U10172 ( .A(a[325]), .B(n2222), .Z(n9116) );
  AND U10173 ( .A(a[327]), .B(b[0]), .Z(n9096) );
  XNOR U10174 ( .A(n9096), .B(n2175), .Z(n9098) );
  NANDN U10175 ( .A(b[0]), .B(a[326]), .Z(n9097) );
  NAND U10176 ( .A(n9098), .B(n9097), .Z(n9121) );
  AND U10177 ( .A(a[323]), .B(b[3]), .Z(n9120) );
  XOR U10178 ( .A(n9121), .B(n9120), .Z(n9123) );
  XOR U10179 ( .A(n9122), .B(n9123), .Z(n9111) );
  NANDN U10180 ( .A(n9100), .B(n9099), .Z(n9104) );
  OR U10181 ( .A(n9102), .B(n9101), .Z(n9103) );
  AND U10182 ( .A(n9104), .B(n9103), .Z(n9110) );
  XOR U10183 ( .A(n9111), .B(n9110), .Z(n9113) );
  XOR U10184 ( .A(n9112), .B(n9113), .Z(n9126) );
  XNOR U10185 ( .A(n9126), .B(sreg[1347]), .Z(n9128) );
  NANDN U10186 ( .A(n9105), .B(sreg[1346]), .Z(n9109) );
  NAND U10187 ( .A(n9107), .B(n9106), .Z(n9108) );
  NAND U10188 ( .A(n9109), .B(n9108), .Z(n9127) );
  XOR U10189 ( .A(n9128), .B(n9127), .Z(c[1347]) );
  NANDN U10190 ( .A(n9111), .B(n9110), .Z(n9115) );
  OR U10191 ( .A(n9113), .B(n9112), .Z(n9114) );
  AND U10192 ( .A(n9115), .B(n9114), .Z(n9133) );
  XOR U10193 ( .A(a[326]), .B(n2222), .Z(n9137) );
  AND U10194 ( .A(a[328]), .B(b[0]), .Z(n9117) );
  XNOR U10195 ( .A(n9117), .B(n2175), .Z(n9119) );
  NANDN U10196 ( .A(b[0]), .B(a[327]), .Z(n9118) );
  NAND U10197 ( .A(n9119), .B(n9118), .Z(n9142) );
  AND U10198 ( .A(a[324]), .B(b[3]), .Z(n9141) );
  XOR U10199 ( .A(n9142), .B(n9141), .Z(n9144) );
  XOR U10200 ( .A(n9143), .B(n9144), .Z(n9132) );
  NANDN U10201 ( .A(n9121), .B(n9120), .Z(n9125) );
  OR U10202 ( .A(n9123), .B(n9122), .Z(n9124) );
  AND U10203 ( .A(n9125), .B(n9124), .Z(n9131) );
  XOR U10204 ( .A(n9132), .B(n9131), .Z(n9134) );
  XOR U10205 ( .A(n9133), .B(n9134), .Z(n9147) );
  XNOR U10206 ( .A(n9147), .B(sreg[1348]), .Z(n9149) );
  NANDN U10207 ( .A(n9126), .B(sreg[1347]), .Z(n9130) );
  NAND U10208 ( .A(n9128), .B(n9127), .Z(n9129) );
  NAND U10209 ( .A(n9130), .B(n9129), .Z(n9148) );
  XOR U10210 ( .A(n9149), .B(n9148), .Z(c[1348]) );
  NANDN U10211 ( .A(n9132), .B(n9131), .Z(n9136) );
  OR U10212 ( .A(n9134), .B(n9133), .Z(n9135) );
  AND U10213 ( .A(n9136), .B(n9135), .Z(n9154) );
  XOR U10214 ( .A(a[327]), .B(n2222), .Z(n9158) );
  AND U10215 ( .A(a[329]), .B(b[0]), .Z(n9138) );
  XNOR U10216 ( .A(n9138), .B(n2175), .Z(n9140) );
  NANDN U10217 ( .A(b[0]), .B(a[328]), .Z(n9139) );
  NAND U10218 ( .A(n9140), .B(n9139), .Z(n9163) );
  AND U10219 ( .A(a[325]), .B(b[3]), .Z(n9162) );
  XOR U10220 ( .A(n9163), .B(n9162), .Z(n9165) );
  XOR U10221 ( .A(n9164), .B(n9165), .Z(n9153) );
  NANDN U10222 ( .A(n9142), .B(n9141), .Z(n9146) );
  OR U10223 ( .A(n9144), .B(n9143), .Z(n9145) );
  AND U10224 ( .A(n9146), .B(n9145), .Z(n9152) );
  XOR U10225 ( .A(n9153), .B(n9152), .Z(n9155) );
  XOR U10226 ( .A(n9154), .B(n9155), .Z(n9168) );
  XNOR U10227 ( .A(n9168), .B(sreg[1349]), .Z(n9170) );
  NANDN U10228 ( .A(n9147), .B(sreg[1348]), .Z(n9151) );
  NAND U10229 ( .A(n9149), .B(n9148), .Z(n9150) );
  NAND U10230 ( .A(n9151), .B(n9150), .Z(n9169) );
  XOR U10231 ( .A(n9170), .B(n9169), .Z(c[1349]) );
  NANDN U10232 ( .A(n9153), .B(n9152), .Z(n9157) );
  OR U10233 ( .A(n9155), .B(n9154), .Z(n9156) );
  AND U10234 ( .A(n9157), .B(n9156), .Z(n9175) );
  XOR U10235 ( .A(a[328]), .B(n2223), .Z(n9179) );
  AND U10236 ( .A(a[326]), .B(b[3]), .Z(n9183) );
  AND U10237 ( .A(a[330]), .B(b[0]), .Z(n9159) );
  XNOR U10238 ( .A(n9159), .B(n2175), .Z(n9161) );
  NANDN U10239 ( .A(b[0]), .B(a[329]), .Z(n9160) );
  NAND U10240 ( .A(n9161), .B(n9160), .Z(n9184) );
  XOR U10241 ( .A(n9183), .B(n9184), .Z(n9186) );
  XOR U10242 ( .A(n9185), .B(n9186), .Z(n9174) );
  NANDN U10243 ( .A(n9163), .B(n9162), .Z(n9167) );
  OR U10244 ( .A(n9165), .B(n9164), .Z(n9166) );
  AND U10245 ( .A(n9167), .B(n9166), .Z(n9173) );
  XOR U10246 ( .A(n9174), .B(n9173), .Z(n9176) );
  XOR U10247 ( .A(n9175), .B(n9176), .Z(n9189) );
  XNOR U10248 ( .A(n9189), .B(sreg[1350]), .Z(n9191) );
  NANDN U10249 ( .A(n9168), .B(sreg[1349]), .Z(n9172) );
  NAND U10250 ( .A(n9170), .B(n9169), .Z(n9171) );
  NAND U10251 ( .A(n9172), .B(n9171), .Z(n9190) );
  XOR U10252 ( .A(n9191), .B(n9190), .Z(c[1350]) );
  NANDN U10253 ( .A(n9174), .B(n9173), .Z(n9178) );
  OR U10254 ( .A(n9176), .B(n9175), .Z(n9177) );
  AND U10255 ( .A(n9178), .B(n9177), .Z(n9197) );
  XOR U10256 ( .A(a[329]), .B(n2223), .Z(n9198) );
  NAND U10257 ( .A(a[331]), .B(b[0]), .Z(n9180) );
  XNOR U10258 ( .A(b[1]), .B(n9180), .Z(n9182) );
  NANDN U10259 ( .A(b[0]), .B(a[330]), .Z(n9181) );
  AND U10260 ( .A(n9182), .B(n9181), .Z(n9202) );
  AND U10261 ( .A(a[327]), .B(b[3]), .Z(n9203) );
  XOR U10262 ( .A(n9202), .B(n9203), .Z(n9204) );
  XNOR U10263 ( .A(n9205), .B(n9204), .Z(n9194) );
  NANDN U10264 ( .A(n9184), .B(n9183), .Z(n9188) );
  OR U10265 ( .A(n9186), .B(n9185), .Z(n9187) );
  AND U10266 ( .A(n9188), .B(n9187), .Z(n9195) );
  XNOR U10267 ( .A(n9194), .B(n9195), .Z(n9196) );
  XNOR U10268 ( .A(n9197), .B(n9196), .Z(n9208) );
  XNOR U10269 ( .A(n9208), .B(sreg[1351]), .Z(n9210) );
  NANDN U10270 ( .A(n9189), .B(sreg[1350]), .Z(n9193) );
  NAND U10271 ( .A(n9191), .B(n9190), .Z(n9192) );
  NAND U10272 ( .A(n9193), .B(n9192), .Z(n9209) );
  XOR U10273 ( .A(n9210), .B(n9209), .Z(c[1351]) );
  XOR U10274 ( .A(a[330]), .B(n2223), .Z(n9217) );
  AND U10275 ( .A(a[332]), .B(b[0]), .Z(n9199) );
  XNOR U10276 ( .A(n9199), .B(n2175), .Z(n9201) );
  NANDN U10277 ( .A(b[0]), .B(a[331]), .Z(n9200) );
  NAND U10278 ( .A(n9201), .B(n9200), .Z(n9222) );
  AND U10279 ( .A(a[328]), .B(b[3]), .Z(n9221) );
  XOR U10280 ( .A(n9222), .B(n9221), .Z(n9224) );
  XOR U10281 ( .A(n9223), .B(n9224), .Z(n9212) );
  NAND U10282 ( .A(n9203), .B(n9202), .Z(n9207) );
  NANDN U10283 ( .A(n9205), .B(n9204), .Z(n9206) );
  AND U10284 ( .A(n9207), .B(n9206), .Z(n9211) );
  XOR U10285 ( .A(n9212), .B(n9211), .Z(n9214) );
  XOR U10286 ( .A(n9213), .B(n9214), .Z(n9227) );
  XNOR U10287 ( .A(n9227), .B(sreg[1352]), .Z(n9229) );
  XOR U10288 ( .A(n9229), .B(n9228), .Z(c[1352]) );
  NANDN U10289 ( .A(n9212), .B(n9211), .Z(n9216) );
  OR U10290 ( .A(n9214), .B(n9213), .Z(n9215) );
  AND U10291 ( .A(n9216), .B(n9215), .Z(n9234) );
  XOR U10292 ( .A(a[331]), .B(n2223), .Z(n9238) );
  AND U10293 ( .A(a[329]), .B(b[3]), .Z(n9242) );
  AND U10294 ( .A(a[333]), .B(b[0]), .Z(n9218) );
  XNOR U10295 ( .A(n9218), .B(n2175), .Z(n9220) );
  NANDN U10296 ( .A(b[0]), .B(a[332]), .Z(n9219) );
  NAND U10297 ( .A(n9220), .B(n9219), .Z(n9243) );
  XOR U10298 ( .A(n9242), .B(n9243), .Z(n9245) );
  XOR U10299 ( .A(n9244), .B(n9245), .Z(n9233) );
  NANDN U10300 ( .A(n9222), .B(n9221), .Z(n9226) );
  OR U10301 ( .A(n9224), .B(n9223), .Z(n9225) );
  AND U10302 ( .A(n9226), .B(n9225), .Z(n9232) );
  XOR U10303 ( .A(n9233), .B(n9232), .Z(n9235) );
  XOR U10304 ( .A(n9234), .B(n9235), .Z(n9248) );
  XNOR U10305 ( .A(n9248), .B(sreg[1353]), .Z(n9250) );
  NANDN U10306 ( .A(n9227), .B(sreg[1352]), .Z(n9231) );
  NAND U10307 ( .A(n9229), .B(n9228), .Z(n9230) );
  NAND U10308 ( .A(n9231), .B(n9230), .Z(n9249) );
  XOR U10309 ( .A(n9250), .B(n9249), .Z(c[1353]) );
  NANDN U10310 ( .A(n9233), .B(n9232), .Z(n9237) );
  OR U10311 ( .A(n9235), .B(n9234), .Z(n9236) );
  AND U10312 ( .A(n9237), .B(n9236), .Z(n9255) );
  XOR U10313 ( .A(a[332]), .B(n2223), .Z(n9259) );
  AND U10314 ( .A(a[334]), .B(b[0]), .Z(n9239) );
  XNOR U10315 ( .A(n9239), .B(n2175), .Z(n9241) );
  NANDN U10316 ( .A(b[0]), .B(a[333]), .Z(n9240) );
  NAND U10317 ( .A(n9241), .B(n9240), .Z(n9264) );
  AND U10318 ( .A(a[330]), .B(b[3]), .Z(n9263) );
  XOR U10319 ( .A(n9264), .B(n9263), .Z(n9266) );
  XOR U10320 ( .A(n9265), .B(n9266), .Z(n9254) );
  NANDN U10321 ( .A(n9243), .B(n9242), .Z(n9247) );
  OR U10322 ( .A(n9245), .B(n9244), .Z(n9246) );
  AND U10323 ( .A(n9247), .B(n9246), .Z(n9253) );
  XOR U10324 ( .A(n9254), .B(n9253), .Z(n9256) );
  XOR U10325 ( .A(n9255), .B(n9256), .Z(n9269) );
  XNOR U10326 ( .A(n9269), .B(sreg[1354]), .Z(n9271) );
  NANDN U10327 ( .A(n9248), .B(sreg[1353]), .Z(n9252) );
  NAND U10328 ( .A(n9250), .B(n9249), .Z(n9251) );
  NAND U10329 ( .A(n9252), .B(n9251), .Z(n9270) );
  XOR U10330 ( .A(n9271), .B(n9270), .Z(c[1354]) );
  NANDN U10331 ( .A(n9254), .B(n9253), .Z(n9258) );
  OR U10332 ( .A(n9256), .B(n9255), .Z(n9257) );
  AND U10333 ( .A(n9258), .B(n9257), .Z(n9276) );
  XOR U10334 ( .A(a[333]), .B(n2223), .Z(n9280) );
  AND U10335 ( .A(a[335]), .B(b[0]), .Z(n9260) );
  XNOR U10336 ( .A(n9260), .B(n2175), .Z(n9262) );
  NANDN U10337 ( .A(b[0]), .B(a[334]), .Z(n9261) );
  NAND U10338 ( .A(n9262), .B(n9261), .Z(n9285) );
  AND U10339 ( .A(a[331]), .B(b[3]), .Z(n9284) );
  XOR U10340 ( .A(n9285), .B(n9284), .Z(n9287) );
  XOR U10341 ( .A(n9286), .B(n9287), .Z(n9275) );
  NANDN U10342 ( .A(n9264), .B(n9263), .Z(n9268) );
  OR U10343 ( .A(n9266), .B(n9265), .Z(n9267) );
  AND U10344 ( .A(n9268), .B(n9267), .Z(n9274) );
  XOR U10345 ( .A(n9275), .B(n9274), .Z(n9277) );
  XOR U10346 ( .A(n9276), .B(n9277), .Z(n9290) );
  XNOR U10347 ( .A(n9290), .B(sreg[1355]), .Z(n9292) );
  NANDN U10348 ( .A(n9269), .B(sreg[1354]), .Z(n9273) );
  NAND U10349 ( .A(n9271), .B(n9270), .Z(n9272) );
  NAND U10350 ( .A(n9273), .B(n9272), .Z(n9291) );
  XOR U10351 ( .A(n9292), .B(n9291), .Z(c[1355]) );
  NANDN U10352 ( .A(n9275), .B(n9274), .Z(n9279) );
  OR U10353 ( .A(n9277), .B(n9276), .Z(n9278) );
  AND U10354 ( .A(n9279), .B(n9278), .Z(n9297) );
  XOR U10355 ( .A(a[334]), .B(n2223), .Z(n9301) );
  AND U10356 ( .A(a[336]), .B(b[0]), .Z(n9281) );
  XNOR U10357 ( .A(n9281), .B(n2175), .Z(n9283) );
  NANDN U10358 ( .A(b[0]), .B(a[335]), .Z(n9282) );
  NAND U10359 ( .A(n9283), .B(n9282), .Z(n9306) );
  AND U10360 ( .A(a[332]), .B(b[3]), .Z(n9305) );
  XOR U10361 ( .A(n9306), .B(n9305), .Z(n9308) );
  XOR U10362 ( .A(n9307), .B(n9308), .Z(n9296) );
  NANDN U10363 ( .A(n9285), .B(n9284), .Z(n9289) );
  OR U10364 ( .A(n9287), .B(n9286), .Z(n9288) );
  AND U10365 ( .A(n9289), .B(n9288), .Z(n9295) );
  XOR U10366 ( .A(n9296), .B(n9295), .Z(n9298) );
  XOR U10367 ( .A(n9297), .B(n9298), .Z(n9311) );
  XNOR U10368 ( .A(n9311), .B(sreg[1356]), .Z(n9313) );
  NANDN U10369 ( .A(n9290), .B(sreg[1355]), .Z(n9294) );
  NAND U10370 ( .A(n9292), .B(n9291), .Z(n9293) );
  NAND U10371 ( .A(n9294), .B(n9293), .Z(n9312) );
  XOR U10372 ( .A(n9313), .B(n9312), .Z(c[1356]) );
  NANDN U10373 ( .A(n9296), .B(n9295), .Z(n9300) );
  OR U10374 ( .A(n9298), .B(n9297), .Z(n9299) );
  AND U10375 ( .A(n9300), .B(n9299), .Z(n9318) );
  XOR U10376 ( .A(a[335]), .B(n2224), .Z(n9322) );
  AND U10377 ( .A(a[337]), .B(b[0]), .Z(n9302) );
  XNOR U10378 ( .A(n9302), .B(n2175), .Z(n9304) );
  NANDN U10379 ( .A(b[0]), .B(a[336]), .Z(n9303) );
  NAND U10380 ( .A(n9304), .B(n9303), .Z(n9327) );
  AND U10381 ( .A(a[333]), .B(b[3]), .Z(n9326) );
  XOR U10382 ( .A(n9327), .B(n9326), .Z(n9329) );
  XOR U10383 ( .A(n9328), .B(n9329), .Z(n9317) );
  NANDN U10384 ( .A(n9306), .B(n9305), .Z(n9310) );
  OR U10385 ( .A(n9308), .B(n9307), .Z(n9309) );
  AND U10386 ( .A(n9310), .B(n9309), .Z(n9316) );
  XOR U10387 ( .A(n9317), .B(n9316), .Z(n9319) );
  XOR U10388 ( .A(n9318), .B(n9319), .Z(n9332) );
  XNOR U10389 ( .A(n9332), .B(sreg[1357]), .Z(n9334) );
  NANDN U10390 ( .A(n9311), .B(sreg[1356]), .Z(n9315) );
  NAND U10391 ( .A(n9313), .B(n9312), .Z(n9314) );
  NAND U10392 ( .A(n9315), .B(n9314), .Z(n9333) );
  XOR U10393 ( .A(n9334), .B(n9333), .Z(c[1357]) );
  NANDN U10394 ( .A(n9317), .B(n9316), .Z(n9321) );
  OR U10395 ( .A(n9319), .B(n9318), .Z(n9320) );
  AND U10396 ( .A(n9321), .B(n9320), .Z(n9339) );
  XOR U10397 ( .A(a[336]), .B(n2224), .Z(n9343) );
  AND U10398 ( .A(a[334]), .B(b[3]), .Z(n9347) );
  AND U10399 ( .A(a[338]), .B(b[0]), .Z(n9323) );
  XNOR U10400 ( .A(n9323), .B(n2175), .Z(n9325) );
  NANDN U10401 ( .A(b[0]), .B(a[337]), .Z(n9324) );
  NAND U10402 ( .A(n9325), .B(n9324), .Z(n9348) );
  XOR U10403 ( .A(n9347), .B(n9348), .Z(n9350) );
  XOR U10404 ( .A(n9349), .B(n9350), .Z(n9338) );
  NANDN U10405 ( .A(n9327), .B(n9326), .Z(n9331) );
  OR U10406 ( .A(n9329), .B(n9328), .Z(n9330) );
  AND U10407 ( .A(n9331), .B(n9330), .Z(n9337) );
  XOR U10408 ( .A(n9338), .B(n9337), .Z(n9340) );
  XOR U10409 ( .A(n9339), .B(n9340), .Z(n9353) );
  XNOR U10410 ( .A(n9353), .B(sreg[1358]), .Z(n9355) );
  NANDN U10411 ( .A(n9332), .B(sreg[1357]), .Z(n9336) );
  NAND U10412 ( .A(n9334), .B(n9333), .Z(n9335) );
  NAND U10413 ( .A(n9336), .B(n9335), .Z(n9354) );
  XOR U10414 ( .A(n9355), .B(n9354), .Z(c[1358]) );
  NANDN U10415 ( .A(n9338), .B(n9337), .Z(n9342) );
  OR U10416 ( .A(n9340), .B(n9339), .Z(n9341) );
  AND U10417 ( .A(n9342), .B(n9341), .Z(n9360) );
  XOR U10418 ( .A(a[337]), .B(n2224), .Z(n9364) );
  AND U10419 ( .A(a[335]), .B(b[3]), .Z(n9368) );
  AND U10420 ( .A(a[339]), .B(b[0]), .Z(n9344) );
  XNOR U10421 ( .A(n9344), .B(n2175), .Z(n9346) );
  NANDN U10422 ( .A(b[0]), .B(a[338]), .Z(n9345) );
  NAND U10423 ( .A(n9346), .B(n9345), .Z(n9369) );
  XOR U10424 ( .A(n9368), .B(n9369), .Z(n9371) );
  XOR U10425 ( .A(n9370), .B(n9371), .Z(n9359) );
  NANDN U10426 ( .A(n9348), .B(n9347), .Z(n9352) );
  OR U10427 ( .A(n9350), .B(n9349), .Z(n9351) );
  AND U10428 ( .A(n9352), .B(n9351), .Z(n9358) );
  XOR U10429 ( .A(n9359), .B(n9358), .Z(n9361) );
  XOR U10430 ( .A(n9360), .B(n9361), .Z(n9374) );
  XNOR U10431 ( .A(n9374), .B(sreg[1359]), .Z(n9376) );
  NANDN U10432 ( .A(n9353), .B(sreg[1358]), .Z(n9357) );
  NAND U10433 ( .A(n9355), .B(n9354), .Z(n9356) );
  NAND U10434 ( .A(n9357), .B(n9356), .Z(n9375) );
  XOR U10435 ( .A(n9376), .B(n9375), .Z(c[1359]) );
  NANDN U10436 ( .A(n9359), .B(n9358), .Z(n9363) );
  OR U10437 ( .A(n9361), .B(n9360), .Z(n9362) );
  AND U10438 ( .A(n9363), .B(n9362), .Z(n9381) );
  XOR U10439 ( .A(a[338]), .B(n2224), .Z(n9385) );
  AND U10440 ( .A(a[340]), .B(b[0]), .Z(n9365) );
  XNOR U10441 ( .A(n9365), .B(n2175), .Z(n9367) );
  NANDN U10442 ( .A(b[0]), .B(a[339]), .Z(n9366) );
  NAND U10443 ( .A(n9367), .B(n9366), .Z(n9390) );
  AND U10444 ( .A(a[336]), .B(b[3]), .Z(n9389) );
  XOR U10445 ( .A(n9390), .B(n9389), .Z(n9392) );
  XOR U10446 ( .A(n9391), .B(n9392), .Z(n9380) );
  NANDN U10447 ( .A(n9369), .B(n9368), .Z(n9373) );
  OR U10448 ( .A(n9371), .B(n9370), .Z(n9372) );
  AND U10449 ( .A(n9373), .B(n9372), .Z(n9379) );
  XOR U10450 ( .A(n9380), .B(n9379), .Z(n9382) );
  XOR U10451 ( .A(n9381), .B(n9382), .Z(n9395) );
  XNOR U10452 ( .A(n9395), .B(sreg[1360]), .Z(n9397) );
  NANDN U10453 ( .A(n9374), .B(sreg[1359]), .Z(n9378) );
  NAND U10454 ( .A(n9376), .B(n9375), .Z(n9377) );
  NAND U10455 ( .A(n9378), .B(n9377), .Z(n9396) );
  XOR U10456 ( .A(n9397), .B(n9396), .Z(c[1360]) );
  NANDN U10457 ( .A(n9380), .B(n9379), .Z(n9384) );
  OR U10458 ( .A(n9382), .B(n9381), .Z(n9383) );
  AND U10459 ( .A(n9384), .B(n9383), .Z(n9402) );
  XOR U10460 ( .A(a[339]), .B(n2224), .Z(n9406) );
  AND U10461 ( .A(a[341]), .B(b[0]), .Z(n9386) );
  XNOR U10462 ( .A(n9386), .B(n2175), .Z(n9388) );
  NANDN U10463 ( .A(b[0]), .B(a[340]), .Z(n9387) );
  NAND U10464 ( .A(n9388), .B(n9387), .Z(n9411) );
  AND U10465 ( .A(a[337]), .B(b[3]), .Z(n9410) );
  XOR U10466 ( .A(n9411), .B(n9410), .Z(n9413) );
  XOR U10467 ( .A(n9412), .B(n9413), .Z(n9401) );
  NANDN U10468 ( .A(n9390), .B(n9389), .Z(n9394) );
  OR U10469 ( .A(n9392), .B(n9391), .Z(n9393) );
  AND U10470 ( .A(n9394), .B(n9393), .Z(n9400) );
  XOR U10471 ( .A(n9401), .B(n9400), .Z(n9403) );
  XOR U10472 ( .A(n9402), .B(n9403), .Z(n9416) );
  XNOR U10473 ( .A(n9416), .B(sreg[1361]), .Z(n9418) );
  NANDN U10474 ( .A(n9395), .B(sreg[1360]), .Z(n9399) );
  NAND U10475 ( .A(n9397), .B(n9396), .Z(n9398) );
  NAND U10476 ( .A(n9399), .B(n9398), .Z(n9417) );
  XOR U10477 ( .A(n9418), .B(n9417), .Z(c[1361]) );
  NANDN U10478 ( .A(n9401), .B(n9400), .Z(n9405) );
  OR U10479 ( .A(n9403), .B(n9402), .Z(n9404) );
  AND U10480 ( .A(n9405), .B(n9404), .Z(n9423) );
  XOR U10481 ( .A(a[340]), .B(n2224), .Z(n9427) );
  AND U10482 ( .A(a[338]), .B(b[3]), .Z(n9431) );
  AND U10483 ( .A(a[342]), .B(b[0]), .Z(n9407) );
  XNOR U10484 ( .A(n9407), .B(n2175), .Z(n9409) );
  NANDN U10485 ( .A(b[0]), .B(a[341]), .Z(n9408) );
  NAND U10486 ( .A(n9409), .B(n9408), .Z(n9432) );
  XOR U10487 ( .A(n9431), .B(n9432), .Z(n9434) );
  XOR U10488 ( .A(n9433), .B(n9434), .Z(n9422) );
  NANDN U10489 ( .A(n9411), .B(n9410), .Z(n9415) );
  OR U10490 ( .A(n9413), .B(n9412), .Z(n9414) );
  AND U10491 ( .A(n9415), .B(n9414), .Z(n9421) );
  XOR U10492 ( .A(n9422), .B(n9421), .Z(n9424) );
  XOR U10493 ( .A(n9423), .B(n9424), .Z(n9437) );
  XNOR U10494 ( .A(n9437), .B(sreg[1362]), .Z(n9439) );
  NANDN U10495 ( .A(n9416), .B(sreg[1361]), .Z(n9420) );
  NAND U10496 ( .A(n9418), .B(n9417), .Z(n9419) );
  NAND U10497 ( .A(n9420), .B(n9419), .Z(n9438) );
  XOR U10498 ( .A(n9439), .B(n9438), .Z(c[1362]) );
  NANDN U10499 ( .A(n9422), .B(n9421), .Z(n9426) );
  OR U10500 ( .A(n9424), .B(n9423), .Z(n9425) );
  AND U10501 ( .A(n9426), .B(n9425), .Z(n9444) );
  XOR U10502 ( .A(a[341]), .B(n2224), .Z(n9448) );
  AND U10503 ( .A(a[343]), .B(b[0]), .Z(n9428) );
  XNOR U10504 ( .A(n9428), .B(n2175), .Z(n9430) );
  NANDN U10505 ( .A(b[0]), .B(a[342]), .Z(n9429) );
  NAND U10506 ( .A(n9430), .B(n9429), .Z(n9453) );
  AND U10507 ( .A(a[339]), .B(b[3]), .Z(n9452) );
  XOR U10508 ( .A(n9453), .B(n9452), .Z(n9455) );
  XOR U10509 ( .A(n9454), .B(n9455), .Z(n9443) );
  NANDN U10510 ( .A(n9432), .B(n9431), .Z(n9436) );
  OR U10511 ( .A(n9434), .B(n9433), .Z(n9435) );
  AND U10512 ( .A(n9436), .B(n9435), .Z(n9442) );
  XOR U10513 ( .A(n9443), .B(n9442), .Z(n9445) );
  XOR U10514 ( .A(n9444), .B(n9445), .Z(n9458) );
  XNOR U10515 ( .A(n9458), .B(sreg[1363]), .Z(n9460) );
  NANDN U10516 ( .A(n9437), .B(sreg[1362]), .Z(n9441) );
  NAND U10517 ( .A(n9439), .B(n9438), .Z(n9440) );
  NAND U10518 ( .A(n9441), .B(n9440), .Z(n9459) );
  XOR U10519 ( .A(n9460), .B(n9459), .Z(c[1363]) );
  NANDN U10520 ( .A(n9443), .B(n9442), .Z(n9447) );
  OR U10521 ( .A(n9445), .B(n9444), .Z(n9446) );
  AND U10522 ( .A(n9447), .B(n9446), .Z(n9465) );
  XOR U10523 ( .A(a[342]), .B(n2225), .Z(n9469) );
  AND U10524 ( .A(a[344]), .B(b[0]), .Z(n9449) );
  XNOR U10525 ( .A(n9449), .B(n2175), .Z(n9451) );
  NANDN U10526 ( .A(b[0]), .B(a[343]), .Z(n9450) );
  NAND U10527 ( .A(n9451), .B(n9450), .Z(n9474) );
  AND U10528 ( .A(a[340]), .B(b[3]), .Z(n9473) );
  XOR U10529 ( .A(n9474), .B(n9473), .Z(n9476) );
  XOR U10530 ( .A(n9475), .B(n9476), .Z(n9464) );
  NANDN U10531 ( .A(n9453), .B(n9452), .Z(n9457) );
  OR U10532 ( .A(n9455), .B(n9454), .Z(n9456) );
  AND U10533 ( .A(n9457), .B(n9456), .Z(n9463) );
  XOR U10534 ( .A(n9464), .B(n9463), .Z(n9466) );
  XOR U10535 ( .A(n9465), .B(n9466), .Z(n9479) );
  XNOR U10536 ( .A(n9479), .B(sreg[1364]), .Z(n9481) );
  NANDN U10537 ( .A(n9458), .B(sreg[1363]), .Z(n9462) );
  NAND U10538 ( .A(n9460), .B(n9459), .Z(n9461) );
  NAND U10539 ( .A(n9462), .B(n9461), .Z(n9480) );
  XOR U10540 ( .A(n9481), .B(n9480), .Z(c[1364]) );
  NANDN U10541 ( .A(n9464), .B(n9463), .Z(n9468) );
  OR U10542 ( .A(n9466), .B(n9465), .Z(n9467) );
  AND U10543 ( .A(n9468), .B(n9467), .Z(n9486) );
  XOR U10544 ( .A(a[343]), .B(n2225), .Z(n9490) );
  AND U10545 ( .A(a[345]), .B(b[0]), .Z(n9470) );
  XNOR U10546 ( .A(n9470), .B(n2175), .Z(n9472) );
  NANDN U10547 ( .A(b[0]), .B(a[344]), .Z(n9471) );
  NAND U10548 ( .A(n9472), .B(n9471), .Z(n9495) );
  AND U10549 ( .A(a[341]), .B(b[3]), .Z(n9494) );
  XOR U10550 ( .A(n9495), .B(n9494), .Z(n9497) );
  XOR U10551 ( .A(n9496), .B(n9497), .Z(n9485) );
  NANDN U10552 ( .A(n9474), .B(n9473), .Z(n9478) );
  OR U10553 ( .A(n9476), .B(n9475), .Z(n9477) );
  AND U10554 ( .A(n9478), .B(n9477), .Z(n9484) );
  XOR U10555 ( .A(n9485), .B(n9484), .Z(n9487) );
  XOR U10556 ( .A(n9486), .B(n9487), .Z(n9500) );
  XNOR U10557 ( .A(n9500), .B(sreg[1365]), .Z(n9502) );
  NANDN U10558 ( .A(n9479), .B(sreg[1364]), .Z(n9483) );
  NAND U10559 ( .A(n9481), .B(n9480), .Z(n9482) );
  NAND U10560 ( .A(n9483), .B(n9482), .Z(n9501) );
  XOR U10561 ( .A(n9502), .B(n9501), .Z(c[1365]) );
  NANDN U10562 ( .A(n9485), .B(n9484), .Z(n9489) );
  OR U10563 ( .A(n9487), .B(n9486), .Z(n9488) );
  AND U10564 ( .A(n9489), .B(n9488), .Z(n9507) );
  XOR U10565 ( .A(a[344]), .B(n2225), .Z(n9511) );
  AND U10566 ( .A(a[346]), .B(b[0]), .Z(n9491) );
  XNOR U10567 ( .A(n9491), .B(n2175), .Z(n9493) );
  NANDN U10568 ( .A(b[0]), .B(a[345]), .Z(n9492) );
  NAND U10569 ( .A(n9493), .B(n9492), .Z(n9516) );
  AND U10570 ( .A(a[342]), .B(b[3]), .Z(n9515) );
  XOR U10571 ( .A(n9516), .B(n9515), .Z(n9518) );
  XOR U10572 ( .A(n9517), .B(n9518), .Z(n9506) );
  NANDN U10573 ( .A(n9495), .B(n9494), .Z(n9499) );
  OR U10574 ( .A(n9497), .B(n9496), .Z(n9498) );
  AND U10575 ( .A(n9499), .B(n9498), .Z(n9505) );
  XOR U10576 ( .A(n9506), .B(n9505), .Z(n9508) );
  XOR U10577 ( .A(n9507), .B(n9508), .Z(n9521) );
  XNOR U10578 ( .A(n9521), .B(sreg[1366]), .Z(n9523) );
  NANDN U10579 ( .A(n9500), .B(sreg[1365]), .Z(n9504) );
  NAND U10580 ( .A(n9502), .B(n9501), .Z(n9503) );
  NAND U10581 ( .A(n9504), .B(n9503), .Z(n9522) );
  XOR U10582 ( .A(n9523), .B(n9522), .Z(c[1366]) );
  NANDN U10583 ( .A(n9506), .B(n9505), .Z(n9510) );
  OR U10584 ( .A(n9508), .B(n9507), .Z(n9509) );
  AND U10585 ( .A(n9510), .B(n9509), .Z(n9528) );
  XOR U10586 ( .A(a[345]), .B(n2225), .Z(n9532) );
  AND U10587 ( .A(a[347]), .B(b[0]), .Z(n9512) );
  XNOR U10588 ( .A(n9512), .B(n2175), .Z(n9514) );
  NANDN U10589 ( .A(b[0]), .B(a[346]), .Z(n9513) );
  NAND U10590 ( .A(n9514), .B(n9513), .Z(n9537) );
  AND U10591 ( .A(a[343]), .B(b[3]), .Z(n9536) );
  XOR U10592 ( .A(n9537), .B(n9536), .Z(n9539) );
  XOR U10593 ( .A(n9538), .B(n9539), .Z(n9527) );
  NANDN U10594 ( .A(n9516), .B(n9515), .Z(n9520) );
  OR U10595 ( .A(n9518), .B(n9517), .Z(n9519) );
  AND U10596 ( .A(n9520), .B(n9519), .Z(n9526) );
  XOR U10597 ( .A(n9527), .B(n9526), .Z(n9529) );
  XOR U10598 ( .A(n9528), .B(n9529), .Z(n9542) );
  XNOR U10599 ( .A(n9542), .B(sreg[1367]), .Z(n9544) );
  NANDN U10600 ( .A(n9521), .B(sreg[1366]), .Z(n9525) );
  NAND U10601 ( .A(n9523), .B(n9522), .Z(n9524) );
  NAND U10602 ( .A(n9525), .B(n9524), .Z(n9543) );
  XOR U10603 ( .A(n9544), .B(n9543), .Z(c[1367]) );
  NANDN U10604 ( .A(n9527), .B(n9526), .Z(n9531) );
  OR U10605 ( .A(n9529), .B(n9528), .Z(n9530) );
  AND U10606 ( .A(n9531), .B(n9530), .Z(n9549) );
  XOR U10607 ( .A(a[346]), .B(n2225), .Z(n9553) );
  AND U10608 ( .A(a[348]), .B(b[0]), .Z(n9533) );
  XNOR U10609 ( .A(n9533), .B(n2175), .Z(n9535) );
  NANDN U10610 ( .A(b[0]), .B(a[347]), .Z(n9534) );
  NAND U10611 ( .A(n9535), .B(n9534), .Z(n9558) );
  AND U10612 ( .A(a[344]), .B(b[3]), .Z(n9557) );
  XOR U10613 ( .A(n9558), .B(n9557), .Z(n9560) );
  XOR U10614 ( .A(n9559), .B(n9560), .Z(n9548) );
  NANDN U10615 ( .A(n9537), .B(n9536), .Z(n9541) );
  OR U10616 ( .A(n9539), .B(n9538), .Z(n9540) );
  AND U10617 ( .A(n9541), .B(n9540), .Z(n9547) );
  XOR U10618 ( .A(n9548), .B(n9547), .Z(n9550) );
  XOR U10619 ( .A(n9549), .B(n9550), .Z(n9563) );
  XNOR U10620 ( .A(n9563), .B(sreg[1368]), .Z(n9565) );
  NANDN U10621 ( .A(n9542), .B(sreg[1367]), .Z(n9546) );
  NAND U10622 ( .A(n9544), .B(n9543), .Z(n9545) );
  NAND U10623 ( .A(n9546), .B(n9545), .Z(n9564) );
  XOR U10624 ( .A(n9565), .B(n9564), .Z(c[1368]) );
  NANDN U10625 ( .A(n9548), .B(n9547), .Z(n9552) );
  OR U10626 ( .A(n9550), .B(n9549), .Z(n9551) );
  AND U10627 ( .A(n9552), .B(n9551), .Z(n9570) );
  XOR U10628 ( .A(a[347]), .B(n2225), .Z(n9574) );
  AND U10629 ( .A(a[345]), .B(b[3]), .Z(n9578) );
  AND U10630 ( .A(a[349]), .B(b[0]), .Z(n9554) );
  XNOR U10631 ( .A(n9554), .B(n2175), .Z(n9556) );
  NANDN U10632 ( .A(b[0]), .B(a[348]), .Z(n9555) );
  NAND U10633 ( .A(n9556), .B(n9555), .Z(n9579) );
  XOR U10634 ( .A(n9578), .B(n9579), .Z(n9581) );
  XOR U10635 ( .A(n9580), .B(n9581), .Z(n9569) );
  NANDN U10636 ( .A(n9558), .B(n9557), .Z(n9562) );
  OR U10637 ( .A(n9560), .B(n9559), .Z(n9561) );
  AND U10638 ( .A(n9562), .B(n9561), .Z(n9568) );
  XOR U10639 ( .A(n9569), .B(n9568), .Z(n9571) );
  XOR U10640 ( .A(n9570), .B(n9571), .Z(n9584) );
  XNOR U10641 ( .A(n9584), .B(sreg[1369]), .Z(n9586) );
  NANDN U10642 ( .A(n9563), .B(sreg[1368]), .Z(n9567) );
  NAND U10643 ( .A(n9565), .B(n9564), .Z(n9566) );
  NAND U10644 ( .A(n9567), .B(n9566), .Z(n9585) );
  XOR U10645 ( .A(n9586), .B(n9585), .Z(c[1369]) );
  NANDN U10646 ( .A(n9569), .B(n9568), .Z(n9573) );
  OR U10647 ( .A(n9571), .B(n9570), .Z(n9572) );
  AND U10648 ( .A(n9573), .B(n9572), .Z(n9591) );
  XOR U10649 ( .A(a[348]), .B(n2225), .Z(n9595) );
  AND U10650 ( .A(a[350]), .B(b[0]), .Z(n9575) );
  XNOR U10651 ( .A(n9575), .B(n2175), .Z(n9577) );
  NANDN U10652 ( .A(b[0]), .B(a[349]), .Z(n9576) );
  NAND U10653 ( .A(n9577), .B(n9576), .Z(n9600) );
  AND U10654 ( .A(a[346]), .B(b[3]), .Z(n9599) );
  XOR U10655 ( .A(n9600), .B(n9599), .Z(n9602) );
  XOR U10656 ( .A(n9601), .B(n9602), .Z(n9590) );
  NANDN U10657 ( .A(n9579), .B(n9578), .Z(n9583) );
  OR U10658 ( .A(n9581), .B(n9580), .Z(n9582) );
  AND U10659 ( .A(n9583), .B(n9582), .Z(n9589) );
  XOR U10660 ( .A(n9590), .B(n9589), .Z(n9592) );
  XOR U10661 ( .A(n9591), .B(n9592), .Z(n9605) );
  XNOR U10662 ( .A(n9605), .B(sreg[1370]), .Z(n9607) );
  NANDN U10663 ( .A(n9584), .B(sreg[1369]), .Z(n9588) );
  NAND U10664 ( .A(n9586), .B(n9585), .Z(n9587) );
  NAND U10665 ( .A(n9588), .B(n9587), .Z(n9606) );
  XOR U10666 ( .A(n9607), .B(n9606), .Z(c[1370]) );
  NANDN U10667 ( .A(n9590), .B(n9589), .Z(n9594) );
  OR U10668 ( .A(n9592), .B(n9591), .Z(n9593) );
  AND U10669 ( .A(n9594), .B(n9593), .Z(n9612) );
  XOR U10670 ( .A(a[349]), .B(n2226), .Z(n9616) );
  AND U10671 ( .A(a[351]), .B(b[0]), .Z(n9596) );
  XNOR U10672 ( .A(n9596), .B(n2175), .Z(n9598) );
  NANDN U10673 ( .A(b[0]), .B(a[350]), .Z(n9597) );
  NAND U10674 ( .A(n9598), .B(n9597), .Z(n9621) );
  AND U10675 ( .A(a[347]), .B(b[3]), .Z(n9620) );
  XOR U10676 ( .A(n9621), .B(n9620), .Z(n9623) );
  XOR U10677 ( .A(n9622), .B(n9623), .Z(n9611) );
  NANDN U10678 ( .A(n9600), .B(n9599), .Z(n9604) );
  OR U10679 ( .A(n9602), .B(n9601), .Z(n9603) );
  AND U10680 ( .A(n9604), .B(n9603), .Z(n9610) );
  XOR U10681 ( .A(n9611), .B(n9610), .Z(n9613) );
  XOR U10682 ( .A(n9612), .B(n9613), .Z(n9626) );
  XNOR U10683 ( .A(n9626), .B(sreg[1371]), .Z(n9628) );
  NANDN U10684 ( .A(n9605), .B(sreg[1370]), .Z(n9609) );
  NAND U10685 ( .A(n9607), .B(n9606), .Z(n9608) );
  NAND U10686 ( .A(n9609), .B(n9608), .Z(n9627) );
  XOR U10687 ( .A(n9628), .B(n9627), .Z(c[1371]) );
  NANDN U10688 ( .A(n9611), .B(n9610), .Z(n9615) );
  OR U10689 ( .A(n9613), .B(n9612), .Z(n9614) );
  AND U10690 ( .A(n9615), .B(n9614), .Z(n9633) );
  XOR U10691 ( .A(a[350]), .B(n2226), .Z(n9637) );
  AND U10692 ( .A(a[352]), .B(b[0]), .Z(n9617) );
  XNOR U10693 ( .A(n9617), .B(n2175), .Z(n9619) );
  NANDN U10694 ( .A(b[0]), .B(a[351]), .Z(n9618) );
  NAND U10695 ( .A(n9619), .B(n9618), .Z(n9642) );
  AND U10696 ( .A(a[348]), .B(b[3]), .Z(n9641) );
  XOR U10697 ( .A(n9642), .B(n9641), .Z(n9644) );
  XOR U10698 ( .A(n9643), .B(n9644), .Z(n9632) );
  NANDN U10699 ( .A(n9621), .B(n9620), .Z(n9625) );
  OR U10700 ( .A(n9623), .B(n9622), .Z(n9624) );
  AND U10701 ( .A(n9625), .B(n9624), .Z(n9631) );
  XOR U10702 ( .A(n9632), .B(n9631), .Z(n9634) );
  XOR U10703 ( .A(n9633), .B(n9634), .Z(n9647) );
  XNOR U10704 ( .A(n9647), .B(sreg[1372]), .Z(n9649) );
  NANDN U10705 ( .A(n9626), .B(sreg[1371]), .Z(n9630) );
  NAND U10706 ( .A(n9628), .B(n9627), .Z(n9629) );
  NAND U10707 ( .A(n9630), .B(n9629), .Z(n9648) );
  XOR U10708 ( .A(n9649), .B(n9648), .Z(c[1372]) );
  NANDN U10709 ( .A(n9632), .B(n9631), .Z(n9636) );
  OR U10710 ( .A(n9634), .B(n9633), .Z(n9635) );
  AND U10711 ( .A(n9636), .B(n9635), .Z(n9654) );
  XOR U10712 ( .A(a[351]), .B(n2226), .Z(n9658) );
  AND U10713 ( .A(a[353]), .B(b[0]), .Z(n9638) );
  XNOR U10714 ( .A(n9638), .B(n2175), .Z(n9640) );
  NANDN U10715 ( .A(b[0]), .B(a[352]), .Z(n9639) );
  NAND U10716 ( .A(n9640), .B(n9639), .Z(n9663) );
  AND U10717 ( .A(a[349]), .B(b[3]), .Z(n9662) );
  XOR U10718 ( .A(n9663), .B(n9662), .Z(n9665) );
  XOR U10719 ( .A(n9664), .B(n9665), .Z(n9653) );
  NANDN U10720 ( .A(n9642), .B(n9641), .Z(n9646) );
  OR U10721 ( .A(n9644), .B(n9643), .Z(n9645) );
  AND U10722 ( .A(n9646), .B(n9645), .Z(n9652) );
  XOR U10723 ( .A(n9653), .B(n9652), .Z(n9655) );
  XOR U10724 ( .A(n9654), .B(n9655), .Z(n9668) );
  XNOR U10725 ( .A(n9668), .B(sreg[1373]), .Z(n9670) );
  NANDN U10726 ( .A(n9647), .B(sreg[1372]), .Z(n9651) );
  NAND U10727 ( .A(n9649), .B(n9648), .Z(n9650) );
  NAND U10728 ( .A(n9651), .B(n9650), .Z(n9669) );
  XOR U10729 ( .A(n9670), .B(n9669), .Z(c[1373]) );
  NANDN U10730 ( .A(n9653), .B(n9652), .Z(n9657) );
  OR U10731 ( .A(n9655), .B(n9654), .Z(n9656) );
  AND U10732 ( .A(n9657), .B(n9656), .Z(n9675) );
  XOR U10733 ( .A(a[352]), .B(n2226), .Z(n9679) );
  AND U10734 ( .A(a[354]), .B(b[0]), .Z(n9659) );
  XNOR U10735 ( .A(n9659), .B(n2175), .Z(n9661) );
  NANDN U10736 ( .A(b[0]), .B(a[353]), .Z(n9660) );
  NAND U10737 ( .A(n9661), .B(n9660), .Z(n9684) );
  AND U10738 ( .A(a[350]), .B(b[3]), .Z(n9683) );
  XOR U10739 ( .A(n9684), .B(n9683), .Z(n9686) );
  XOR U10740 ( .A(n9685), .B(n9686), .Z(n9674) );
  NANDN U10741 ( .A(n9663), .B(n9662), .Z(n9667) );
  OR U10742 ( .A(n9665), .B(n9664), .Z(n9666) );
  AND U10743 ( .A(n9667), .B(n9666), .Z(n9673) );
  XOR U10744 ( .A(n9674), .B(n9673), .Z(n9676) );
  XOR U10745 ( .A(n9675), .B(n9676), .Z(n9689) );
  XNOR U10746 ( .A(n9689), .B(sreg[1374]), .Z(n9691) );
  NANDN U10747 ( .A(n9668), .B(sreg[1373]), .Z(n9672) );
  NAND U10748 ( .A(n9670), .B(n9669), .Z(n9671) );
  NAND U10749 ( .A(n9672), .B(n9671), .Z(n9690) );
  XOR U10750 ( .A(n9691), .B(n9690), .Z(c[1374]) );
  NANDN U10751 ( .A(n9674), .B(n9673), .Z(n9678) );
  OR U10752 ( .A(n9676), .B(n9675), .Z(n9677) );
  AND U10753 ( .A(n9678), .B(n9677), .Z(n9696) );
  XOR U10754 ( .A(a[353]), .B(n2226), .Z(n9700) );
  AND U10755 ( .A(a[351]), .B(b[3]), .Z(n9704) );
  AND U10756 ( .A(a[355]), .B(b[0]), .Z(n9680) );
  XNOR U10757 ( .A(n9680), .B(n2175), .Z(n9682) );
  NANDN U10758 ( .A(b[0]), .B(a[354]), .Z(n9681) );
  NAND U10759 ( .A(n9682), .B(n9681), .Z(n9705) );
  XOR U10760 ( .A(n9704), .B(n9705), .Z(n9707) );
  XOR U10761 ( .A(n9706), .B(n9707), .Z(n9695) );
  NANDN U10762 ( .A(n9684), .B(n9683), .Z(n9688) );
  OR U10763 ( .A(n9686), .B(n9685), .Z(n9687) );
  AND U10764 ( .A(n9688), .B(n9687), .Z(n9694) );
  XOR U10765 ( .A(n9695), .B(n9694), .Z(n9697) );
  XOR U10766 ( .A(n9696), .B(n9697), .Z(n9710) );
  XNOR U10767 ( .A(n9710), .B(sreg[1375]), .Z(n9712) );
  NANDN U10768 ( .A(n9689), .B(sreg[1374]), .Z(n9693) );
  NAND U10769 ( .A(n9691), .B(n9690), .Z(n9692) );
  NAND U10770 ( .A(n9693), .B(n9692), .Z(n9711) );
  XOR U10771 ( .A(n9712), .B(n9711), .Z(c[1375]) );
  NANDN U10772 ( .A(n9695), .B(n9694), .Z(n9699) );
  OR U10773 ( .A(n9697), .B(n9696), .Z(n9698) );
  AND U10774 ( .A(n9699), .B(n9698), .Z(n9717) );
  XOR U10775 ( .A(a[354]), .B(n2226), .Z(n9721) );
  AND U10776 ( .A(a[356]), .B(b[0]), .Z(n9701) );
  XNOR U10777 ( .A(n9701), .B(n2175), .Z(n9703) );
  NANDN U10778 ( .A(b[0]), .B(a[355]), .Z(n9702) );
  NAND U10779 ( .A(n9703), .B(n9702), .Z(n9726) );
  AND U10780 ( .A(a[352]), .B(b[3]), .Z(n9725) );
  XOR U10781 ( .A(n9726), .B(n9725), .Z(n9728) );
  XOR U10782 ( .A(n9727), .B(n9728), .Z(n9716) );
  NANDN U10783 ( .A(n9705), .B(n9704), .Z(n9709) );
  OR U10784 ( .A(n9707), .B(n9706), .Z(n9708) );
  AND U10785 ( .A(n9709), .B(n9708), .Z(n9715) );
  XOR U10786 ( .A(n9716), .B(n9715), .Z(n9718) );
  XOR U10787 ( .A(n9717), .B(n9718), .Z(n9731) );
  XNOR U10788 ( .A(n9731), .B(sreg[1376]), .Z(n9733) );
  NANDN U10789 ( .A(n9710), .B(sreg[1375]), .Z(n9714) );
  NAND U10790 ( .A(n9712), .B(n9711), .Z(n9713) );
  NAND U10791 ( .A(n9714), .B(n9713), .Z(n9732) );
  XOR U10792 ( .A(n9733), .B(n9732), .Z(c[1376]) );
  NANDN U10793 ( .A(n9716), .B(n9715), .Z(n9720) );
  OR U10794 ( .A(n9718), .B(n9717), .Z(n9719) );
  AND U10795 ( .A(n9720), .B(n9719), .Z(n9738) );
  XOR U10796 ( .A(a[355]), .B(n2226), .Z(n9742) );
  AND U10797 ( .A(a[357]), .B(b[0]), .Z(n9722) );
  XNOR U10798 ( .A(n9722), .B(n2175), .Z(n9724) );
  NANDN U10799 ( .A(b[0]), .B(a[356]), .Z(n9723) );
  NAND U10800 ( .A(n9724), .B(n9723), .Z(n9747) );
  AND U10801 ( .A(a[353]), .B(b[3]), .Z(n9746) );
  XOR U10802 ( .A(n9747), .B(n9746), .Z(n9749) );
  XOR U10803 ( .A(n9748), .B(n9749), .Z(n9737) );
  NANDN U10804 ( .A(n9726), .B(n9725), .Z(n9730) );
  OR U10805 ( .A(n9728), .B(n9727), .Z(n9729) );
  AND U10806 ( .A(n9730), .B(n9729), .Z(n9736) );
  XOR U10807 ( .A(n9737), .B(n9736), .Z(n9739) );
  XOR U10808 ( .A(n9738), .B(n9739), .Z(n9752) );
  XNOR U10809 ( .A(n9752), .B(sreg[1377]), .Z(n9754) );
  NANDN U10810 ( .A(n9731), .B(sreg[1376]), .Z(n9735) );
  NAND U10811 ( .A(n9733), .B(n9732), .Z(n9734) );
  NAND U10812 ( .A(n9735), .B(n9734), .Z(n9753) );
  XOR U10813 ( .A(n9754), .B(n9753), .Z(c[1377]) );
  NANDN U10814 ( .A(n9737), .B(n9736), .Z(n9741) );
  OR U10815 ( .A(n9739), .B(n9738), .Z(n9740) );
  AND U10816 ( .A(n9741), .B(n9740), .Z(n9759) );
  XOR U10817 ( .A(a[356]), .B(n2227), .Z(n9763) );
  AND U10818 ( .A(a[358]), .B(b[0]), .Z(n9743) );
  XNOR U10819 ( .A(n9743), .B(n2175), .Z(n9745) );
  NANDN U10820 ( .A(b[0]), .B(a[357]), .Z(n9744) );
  NAND U10821 ( .A(n9745), .B(n9744), .Z(n9768) );
  AND U10822 ( .A(a[354]), .B(b[3]), .Z(n9767) );
  XOR U10823 ( .A(n9768), .B(n9767), .Z(n9770) );
  XOR U10824 ( .A(n9769), .B(n9770), .Z(n9758) );
  NANDN U10825 ( .A(n9747), .B(n9746), .Z(n9751) );
  OR U10826 ( .A(n9749), .B(n9748), .Z(n9750) );
  AND U10827 ( .A(n9751), .B(n9750), .Z(n9757) );
  XOR U10828 ( .A(n9758), .B(n9757), .Z(n9760) );
  XOR U10829 ( .A(n9759), .B(n9760), .Z(n9773) );
  XNOR U10830 ( .A(n9773), .B(sreg[1378]), .Z(n9775) );
  NANDN U10831 ( .A(n9752), .B(sreg[1377]), .Z(n9756) );
  NAND U10832 ( .A(n9754), .B(n9753), .Z(n9755) );
  NAND U10833 ( .A(n9756), .B(n9755), .Z(n9774) );
  XOR U10834 ( .A(n9775), .B(n9774), .Z(c[1378]) );
  NANDN U10835 ( .A(n9758), .B(n9757), .Z(n9762) );
  OR U10836 ( .A(n9760), .B(n9759), .Z(n9761) );
  AND U10837 ( .A(n9762), .B(n9761), .Z(n9780) );
  XOR U10838 ( .A(a[357]), .B(n2227), .Z(n9784) );
  AND U10839 ( .A(a[355]), .B(b[3]), .Z(n9788) );
  AND U10840 ( .A(a[359]), .B(b[0]), .Z(n9764) );
  XNOR U10841 ( .A(n9764), .B(n2175), .Z(n9766) );
  NANDN U10842 ( .A(b[0]), .B(a[358]), .Z(n9765) );
  NAND U10843 ( .A(n9766), .B(n9765), .Z(n9789) );
  XOR U10844 ( .A(n9788), .B(n9789), .Z(n9791) );
  XOR U10845 ( .A(n9790), .B(n9791), .Z(n9779) );
  NANDN U10846 ( .A(n9768), .B(n9767), .Z(n9772) );
  OR U10847 ( .A(n9770), .B(n9769), .Z(n9771) );
  AND U10848 ( .A(n9772), .B(n9771), .Z(n9778) );
  XOR U10849 ( .A(n9779), .B(n9778), .Z(n9781) );
  XOR U10850 ( .A(n9780), .B(n9781), .Z(n9794) );
  XNOR U10851 ( .A(n9794), .B(sreg[1379]), .Z(n9796) );
  NANDN U10852 ( .A(n9773), .B(sreg[1378]), .Z(n9777) );
  NAND U10853 ( .A(n9775), .B(n9774), .Z(n9776) );
  NAND U10854 ( .A(n9777), .B(n9776), .Z(n9795) );
  XOR U10855 ( .A(n9796), .B(n9795), .Z(c[1379]) );
  NANDN U10856 ( .A(n9779), .B(n9778), .Z(n9783) );
  OR U10857 ( .A(n9781), .B(n9780), .Z(n9782) );
  AND U10858 ( .A(n9783), .B(n9782), .Z(n9801) );
  XOR U10859 ( .A(a[358]), .B(n2227), .Z(n9805) );
  AND U10860 ( .A(a[356]), .B(b[3]), .Z(n9809) );
  AND U10861 ( .A(a[360]), .B(b[0]), .Z(n9785) );
  XNOR U10862 ( .A(n9785), .B(n2175), .Z(n9787) );
  NANDN U10863 ( .A(b[0]), .B(a[359]), .Z(n9786) );
  NAND U10864 ( .A(n9787), .B(n9786), .Z(n9810) );
  XOR U10865 ( .A(n9809), .B(n9810), .Z(n9812) );
  XOR U10866 ( .A(n9811), .B(n9812), .Z(n9800) );
  NANDN U10867 ( .A(n9789), .B(n9788), .Z(n9793) );
  OR U10868 ( .A(n9791), .B(n9790), .Z(n9792) );
  AND U10869 ( .A(n9793), .B(n9792), .Z(n9799) );
  XOR U10870 ( .A(n9800), .B(n9799), .Z(n9802) );
  XOR U10871 ( .A(n9801), .B(n9802), .Z(n9815) );
  XNOR U10872 ( .A(n9815), .B(sreg[1380]), .Z(n9817) );
  NANDN U10873 ( .A(n9794), .B(sreg[1379]), .Z(n9798) );
  NAND U10874 ( .A(n9796), .B(n9795), .Z(n9797) );
  NAND U10875 ( .A(n9798), .B(n9797), .Z(n9816) );
  XOR U10876 ( .A(n9817), .B(n9816), .Z(c[1380]) );
  NANDN U10877 ( .A(n9800), .B(n9799), .Z(n9804) );
  OR U10878 ( .A(n9802), .B(n9801), .Z(n9803) );
  AND U10879 ( .A(n9804), .B(n9803), .Z(n9822) );
  XOR U10880 ( .A(a[359]), .B(n2227), .Z(n9826) );
  AND U10881 ( .A(a[361]), .B(b[0]), .Z(n9806) );
  XNOR U10882 ( .A(n9806), .B(n2175), .Z(n9808) );
  NANDN U10883 ( .A(b[0]), .B(a[360]), .Z(n9807) );
  NAND U10884 ( .A(n9808), .B(n9807), .Z(n9831) );
  AND U10885 ( .A(a[357]), .B(b[3]), .Z(n9830) );
  XOR U10886 ( .A(n9831), .B(n9830), .Z(n9833) );
  XOR U10887 ( .A(n9832), .B(n9833), .Z(n9821) );
  NANDN U10888 ( .A(n9810), .B(n9809), .Z(n9814) );
  OR U10889 ( .A(n9812), .B(n9811), .Z(n9813) );
  AND U10890 ( .A(n9814), .B(n9813), .Z(n9820) );
  XOR U10891 ( .A(n9821), .B(n9820), .Z(n9823) );
  XOR U10892 ( .A(n9822), .B(n9823), .Z(n9836) );
  XNOR U10893 ( .A(n9836), .B(sreg[1381]), .Z(n9838) );
  NANDN U10894 ( .A(n9815), .B(sreg[1380]), .Z(n9819) );
  NAND U10895 ( .A(n9817), .B(n9816), .Z(n9818) );
  NAND U10896 ( .A(n9819), .B(n9818), .Z(n9837) );
  XOR U10897 ( .A(n9838), .B(n9837), .Z(c[1381]) );
  NANDN U10898 ( .A(n9821), .B(n9820), .Z(n9825) );
  OR U10899 ( .A(n9823), .B(n9822), .Z(n9824) );
  AND U10900 ( .A(n9825), .B(n9824), .Z(n9843) );
  XOR U10901 ( .A(a[360]), .B(n2227), .Z(n9847) );
  AND U10902 ( .A(a[358]), .B(b[3]), .Z(n9851) );
  AND U10903 ( .A(a[362]), .B(b[0]), .Z(n9827) );
  XNOR U10904 ( .A(n9827), .B(n2175), .Z(n9829) );
  NANDN U10905 ( .A(b[0]), .B(a[361]), .Z(n9828) );
  NAND U10906 ( .A(n9829), .B(n9828), .Z(n9852) );
  XOR U10907 ( .A(n9851), .B(n9852), .Z(n9854) );
  XOR U10908 ( .A(n9853), .B(n9854), .Z(n9842) );
  NANDN U10909 ( .A(n9831), .B(n9830), .Z(n9835) );
  OR U10910 ( .A(n9833), .B(n9832), .Z(n9834) );
  AND U10911 ( .A(n9835), .B(n9834), .Z(n9841) );
  XOR U10912 ( .A(n9842), .B(n9841), .Z(n9844) );
  XOR U10913 ( .A(n9843), .B(n9844), .Z(n9857) );
  XNOR U10914 ( .A(n9857), .B(sreg[1382]), .Z(n9859) );
  NANDN U10915 ( .A(n9836), .B(sreg[1381]), .Z(n9840) );
  NAND U10916 ( .A(n9838), .B(n9837), .Z(n9839) );
  NAND U10917 ( .A(n9840), .B(n9839), .Z(n9858) );
  XOR U10918 ( .A(n9859), .B(n9858), .Z(c[1382]) );
  NANDN U10919 ( .A(n9842), .B(n9841), .Z(n9846) );
  OR U10920 ( .A(n9844), .B(n9843), .Z(n9845) );
  AND U10921 ( .A(n9846), .B(n9845), .Z(n9864) );
  XOR U10922 ( .A(a[361]), .B(n2227), .Z(n9868) );
  AND U10923 ( .A(a[363]), .B(b[0]), .Z(n9848) );
  XNOR U10924 ( .A(n9848), .B(n2175), .Z(n9850) );
  NANDN U10925 ( .A(b[0]), .B(a[362]), .Z(n9849) );
  NAND U10926 ( .A(n9850), .B(n9849), .Z(n9873) );
  AND U10927 ( .A(a[359]), .B(b[3]), .Z(n9872) );
  XOR U10928 ( .A(n9873), .B(n9872), .Z(n9875) );
  XOR U10929 ( .A(n9874), .B(n9875), .Z(n9863) );
  NANDN U10930 ( .A(n9852), .B(n9851), .Z(n9856) );
  OR U10931 ( .A(n9854), .B(n9853), .Z(n9855) );
  AND U10932 ( .A(n9856), .B(n9855), .Z(n9862) );
  XOR U10933 ( .A(n9863), .B(n9862), .Z(n9865) );
  XOR U10934 ( .A(n9864), .B(n9865), .Z(n9878) );
  XNOR U10935 ( .A(n9878), .B(sreg[1383]), .Z(n9880) );
  NANDN U10936 ( .A(n9857), .B(sreg[1382]), .Z(n9861) );
  NAND U10937 ( .A(n9859), .B(n9858), .Z(n9860) );
  NAND U10938 ( .A(n9861), .B(n9860), .Z(n9879) );
  XOR U10939 ( .A(n9880), .B(n9879), .Z(c[1383]) );
  NANDN U10940 ( .A(n9863), .B(n9862), .Z(n9867) );
  OR U10941 ( .A(n9865), .B(n9864), .Z(n9866) );
  AND U10942 ( .A(n9867), .B(n9866), .Z(n9885) );
  XOR U10943 ( .A(a[362]), .B(n2227), .Z(n9889) );
  AND U10944 ( .A(a[364]), .B(b[0]), .Z(n9869) );
  XNOR U10945 ( .A(n9869), .B(n2175), .Z(n9871) );
  NANDN U10946 ( .A(b[0]), .B(a[363]), .Z(n9870) );
  NAND U10947 ( .A(n9871), .B(n9870), .Z(n9894) );
  AND U10948 ( .A(a[360]), .B(b[3]), .Z(n9893) );
  XOR U10949 ( .A(n9894), .B(n9893), .Z(n9896) );
  XOR U10950 ( .A(n9895), .B(n9896), .Z(n9884) );
  NANDN U10951 ( .A(n9873), .B(n9872), .Z(n9877) );
  OR U10952 ( .A(n9875), .B(n9874), .Z(n9876) );
  AND U10953 ( .A(n9877), .B(n9876), .Z(n9883) );
  XOR U10954 ( .A(n9884), .B(n9883), .Z(n9886) );
  XOR U10955 ( .A(n9885), .B(n9886), .Z(n9899) );
  XNOR U10956 ( .A(n9899), .B(sreg[1384]), .Z(n9901) );
  NANDN U10957 ( .A(n9878), .B(sreg[1383]), .Z(n9882) );
  NAND U10958 ( .A(n9880), .B(n9879), .Z(n9881) );
  NAND U10959 ( .A(n9882), .B(n9881), .Z(n9900) );
  XOR U10960 ( .A(n9901), .B(n9900), .Z(c[1384]) );
  NANDN U10961 ( .A(n9884), .B(n9883), .Z(n9888) );
  OR U10962 ( .A(n9886), .B(n9885), .Z(n9887) );
  AND U10963 ( .A(n9888), .B(n9887), .Z(n9906) );
  XOR U10964 ( .A(a[363]), .B(n2228), .Z(n9910) );
  AND U10965 ( .A(a[361]), .B(b[3]), .Z(n9914) );
  AND U10966 ( .A(a[365]), .B(b[0]), .Z(n9890) );
  XNOR U10967 ( .A(n9890), .B(n2175), .Z(n9892) );
  NANDN U10968 ( .A(b[0]), .B(a[364]), .Z(n9891) );
  NAND U10969 ( .A(n9892), .B(n9891), .Z(n9915) );
  XOR U10970 ( .A(n9914), .B(n9915), .Z(n9917) );
  XOR U10971 ( .A(n9916), .B(n9917), .Z(n9905) );
  NANDN U10972 ( .A(n9894), .B(n9893), .Z(n9898) );
  OR U10973 ( .A(n9896), .B(n9895), .Z(n9897) );
  AND U10974 ( .A(n9898), .B(n9897), .Z(n9904) );
  XOR U10975 ( .A(n9905), .B(n9904), .Z(n9907) );
  XOR U10976 ( .A(n9906), .B(n9907), .Z(n9920) );
  XNOR U10977 ( .A(n9920), .B(sreg[1385]), .Z(n9922) );
  NANDN U10978 ( .A(n9899), .B(sreg[1384]), .Z(n9903) );
  NAND U10979 ( .A(n9901), .B(n9900), .Z(n9902) );
  NAND U10980 ( .A(n9903), .B(n9902), .Z(n9921) );
  XOR U10981 ( .A(n9922), .B(n9921), .Z(c[1385]) );
  NANDN U10982 ( .A(n9905), .B(n9904), .Z(n9909) );
  OR U10983 ( .A(n9907), .B(n9906), .Z(n9908) );
  AND U10984 ( .A(n9909), .B(n9908), .Z(n9927) );
  XOR U10985 ( .A(a[364]), .B(n2228), .Z(n9931) );
  AND U10986 ( .A(a[366]), .B(b[0]), .Z(n9911) );
  XNOR U10987 ( .A(n9911), .B(n2175), .Z(n9913) );
  NANDN U10988 ( .A(b[0]), .B(a[365]), .Z(n9912) );
  NAND U10989 ( .A(n9913), .B(n9912), .Z(n9936) );
  AND U10990 ( .A(a[362]), .B(b[3]), .Z(n9935) );
  XOR U10991 ( .A(n9936), .B(n9935), .Z(n9938) );
  XOR U10992 ( .A(n9937), .B(n9938), .Z(n9926) );
  NANDN U10993 ( .A(n9915), .B(n9914), .Z(n9919) );
  OR U10994 ( .A(n9917), .B(n9916), .Z(n9918) );
  AND U10995 ( .A(n9919), .B(n9918), .Z(n9925) );
  XOR U10996 ( .A(n9926), .B(n9925), .Z(n9928) );
  XOR U10997 ( .A(n9927), .B(n9928), .Z(n9941) );
  XNOR U10998 ( .A(n9941), .B(sreg[1386]), .Z(n9943) );
  NANDN U10999 ( .A(n9920), .B(sreg[1385]), .Z(n9924) );
  NAND U11000 ( .A(n9922), .B(n9921), .Z(n9923) );
  NAND U11001 ( .A(n9924), .B(n9923), .Z(n9942) );
  XOR U11002 ( .A(n9943), .B(n9942), .Z(c[1386]) );
  NANDN U11003 ( .A(n9926), .B(n9925), .Z(n9930) );
  OR U11004 ( .A(n9928), .B(n9927), .Z(n9929) );
  AND U11005 ( .A(n9930), .B(n9929), .Z(n9948) );
  XOR U11006 ( .A(a[365]), .B(n2228), .Z(n9952) );
  AND U11007 ( .A(a[363]), .B(b[3]), .Z(n9956) );
  AND U11008 ( .A(a[367]), .B(b[0]), .Z(n9932) );
  XNOR U11009 ( .A(n9932), .B(n2175), .Z(n9934) );
  NANDN U11010 ( .A(b[0]), .B(a[366]), .Z(n9933) );
  NAND U11011 ( .A(n9934), .B(n9933), .Z(n9957) );
  XOR U11012 ( .A(n9956), .B(n9957), .Z(n9959) );
  XOR U11013 ( .A(n9958), .B(n9959), .Z(n9947) );
  NANDN U11014 ( .A(n9936), .B(n9935), .Z(n9940) );
  OR U11015 ( .A(n9938), .B(n9937), .Z(n9939) );
  AND U11016 ( .A(n9940), .B(n9939), .Z(n9946) );
  XOR U11017 ( .A(n9947), .B(n9946), .Z(n9949) );
  XOR U11018 ( .A(n9948), .B(n9949), .Z(n9962) );
  XNOR U11019 ( .A(n9962), .B(sreg[1387]), .Z(n9964) );
  NANDN U11020 ( .A(n9941), .B(sreg[1386]), .Z(n9945) );
  NAND U11021 ( .A(n9943), .B(n9942), .Z(n9944) );
  NAND U11022 ( .A(n9945), .B(n9944), .Z(n9963) );
  XOR U11023 ( .A(n9964), .B(n9963), .Z(c[1387]) );
  NANDN U11024 ( .A(n9947), .B(n9946), .Z(n9951) );
  OR U11025 ( .A(n9949), .B(n9948), .Z(n9950) );
  AND U11026 ( .A(n9951), .B(n9950), .Z(n9969) );
  XOR U11027 ( .A(a[366]), .B(n2228), .Z(n9973) );
  AND U11028 ( .A(a[364]), .B(b[3]), .Z(n9977) );
  AND U11029 ( .A(a[368]), .B(b[0]), .Z(n9953) );
  XNOR U11030 ( .A(n9953), .B(n2175), .Z(n9955) );
  NANDN U11031 ( .A(b[0]), .B(a[367]), .Z(n9954) );
  NAND U11032 ( .A(n9955), .B(n9954), .Z(n9978) );
  XOR U11033 ( .A(n9977), .B(n9978), .Z(n9980) );
  XOR U11034 ( .A(n9979), .B(n9980), .Z(n9968) );
  NANDN U11035 ( .A(n9957), .B(n9956), .Z(n9961) );
  OR U11036 ( .A(n9959), .B(n9958), .Z(n9960) );
  AND U11037 ( .A(n9961), .B(n9960), .Z(n9967) );
  XOR U11038 ( .A(n9968), .B(n9967), .Z(n9970) );
  XOR U11039 ( .A(n9969), .B(n9970), .Z(n9983) );
  XNOR U11040 ( .A(n9983), .B(sreg[1388]), .Z(n9985) );
  NANDN U11041 ( .A(n9962), .B(sreg[1387]), .Z(n9966) );
  NAND U11042 ( .A(n9964), .B(n9963), .Z(n9965) );
  NAND U11043 ( .A(n9966), .B(n9965), .Z(n9984) );
  XOR U11044 ( .A(n9985), .B(n9984), .Z(c[1388]) );
  NANDN U11045 ( .A(n9968), .B(n9967), .Z(n9972) );
  OR U11046 ( .A(n9970), .B(n9969), .Z(n9971) );
  AND U11047 ( .A(n9972), .B(n9971), .Z(n9990) );
  XOR U11048 ( .A(a[367]), .B(n2228), .Z(n9994) );
  AND U11049 ( .A(a[369]), .B(b[0]), .Z(n9974) );
  XNOR U11050 ( .A(n9974), .B(n2175), .Z(n9976) );
  NANDN U11051 ( .A(b[0]), .B(a[368]), .Z(n9975) );
  NAND U11052 ( .A(n9976), .B(n9975), .Z(n9999) );
  AND U11053 ( .A(a[365]), .B(b[3]), .Z(n9998) );
  XOR U11054 ( .A(n9999), .B(n9998), .Z(n10001) );
  XOR U11055 ( .A(n10000), .B(n10001), .Z(n9989) );
  NANDN U11056 ( .A(n9978), .B(n9977), .Z(n9982) );
  OR U11057 ( .A(n9980), .B(n9979), .Z(n9981) );
  AND U11058 ( .A(n9982), .B(n9981), .Z(n9988) );
  XOR U11059 ( .A(n9989), .B(n9988), .Z(n9991) );
  XOR U11060 ( .A(n9990), .B(n9991), .Z(n10004) );
  XNOR U11061 ( .A(n10004), .B(sreg[1389]), .Z(n10006) );
  NANDN U11062 ( .A(n9983), .B(sreg[1388]), .Z(n9987) );
  NAND U11063 ( .A(n9985), .B(n9984), .Z(n9986) );
  NAND U11064 ( .A(n9987), .B(n9986), .Z(n10005) );
  XOR U11065 ( .A(n10006), .B(n10005), .Z(c[1389]) );
  NANDN U11066 ( .A(n9989), .B(n9988), .Z(n9993) );
  OR U11067 ( .A(n9991), .B(n9990), .Z(n9992) );
  AND U11068 ( .A(n9993), .B(n9992), .Z(n10011) );
  XOR U11069 ( .A(a[368]), .B(n2228), .Z(n10015) );
  AND U11070 ( .A(a[370]), .B(b[0]), .Z(n9995) );
  XNOR U11071 ( .A(n9995), .B(n2175), .Z(n9997) );
  NANDN U11072 ( .A(b[0]), .B(a[369]), .Z(n9996) );
  NAND U11073 ( .A(n9997), .B(n9996), .Z(n10020) );
  AND U11074 ( .A(a[366]), .B(b[3]), .Z(n10019) );
  XOR U11075 ( .A(n10020), .B(n10019), .Z(n10022) );
  XOR U11076 ( .A(n10021), .B(n10022), .Z(n10010) );
  NANDN U11077 ( .A(n9999), .B(n9998), .Z(n10003) );
  OR U11078 ( .A(n10001), .B(n10000), .Z(n10002) );
  AND U11079 ( .A(n10003), .B(n10002), .Z(n10009) );
  XOR U11080 ( .A(n10010), .B(n10009), .Z(n10012) );
  XOR U11081 ( .A(n10011), .B(n10012), .Z(n10025) );
  XNOR U11082 ( .A(n10025), .B(sreg[1390]), .Z(n10027) );
  NANDN U11083 ( .A(n10004), .B(sreg[1389]), .Z(n10008) );
  NAND U11084 ( .A(n10006), .B(n10005), .Z(n10007) );
  NAND U11085 ( .A(n10008), .B(n10007), .Z(n10026) );
  XOR U11086 ( .A(n10027), .B(n10026), .Z(c[1390]) );
  NANDN U11087 ( .A(n10010), .B(n10009), .Z(n10014) );
  OR U11088 ( .A(n10012), .B(n10011), .Z(n10013) );
  AND U11089 ( .A(n10014), .B(n10013), .Z(n10032) );
  XOR U11090 ( .A(a[369]), .B(n2228), .Z(n10036) );
  AND U11091 ( .A(a[371]), .B(b[0]), .Z(n10016) );
  XNOR U11092 ( .A(n10016), .B(n2175), .Z(n10018) );
  NANDN U11093 ( .A(b[0]), .B(a[370]), .Z(n10017) );
  NAND U11094 ( .A(n10018), .B(n10017), .Z(n10041) );
  AND U11095 ( .A(a[367]), .B(b[3]), .Z(n10040) );
  XOR U11096 ( .A(n10041), .B(n10040), .Z(n10043) );
  XOR U11097 ( .A(n10042), .B(n10043), .Z(n10031) );
  NANDN U11098 ( .A(n10020), .B(n10019), .Z(n10024) );
  OR U11099 ( .A(n10022), .B(n10021), .Z(n10023) );
  AND U11100 ( .A(n10024), .B(n10023), .Z(n10030) );
  XOR U11101 ( .A(n10031), .B(n10030), .Z(n10033) );
  XOR U11102 ( .A(n10032), .B(n10033), .Z(n10046) );
  XNOR U11103 ( .A(n10046), .B(sreg[1391]), .Z(n10048) );
  NANDN U11104 ( .A(n10025), .B(sreg[1390]), .Z(n10029) );
  NAND U11105 ( .A(n10027), .B(n10026), .Z(n10028) );
  NAND U11106 ( .A(n10029), .B(n10028), .Z(n10047) );
  XOR U11107 ( .A(n10048), .B(n10047), .Z(c[1391]) );
  NANDN U11108 ( .A(n10031), .B(n10030), .Z(n10035) );
  OR U11109 ( .A(n10033), .B(n10032), .Z(n10034) );
  AND U11110 ( .A(n10035), .B(n10034), .Z(n10053) );
  XOR U11111 ( .A(a[370]), .B(n2229), .Z(n10057) );
  AND U11112 ( .A(a[368]), .B(b[3]), .Z(n10061) );
  AND U11113 ( .A(a[372]), .B(b[0]), .Z(n10037) );
  XNOR U11114 ( .A(n10037), .B(n2175), .Z(n10039) );
  NANDN U11115 ( .A(b[0]), .B(a[371]), .Z(n10038) );
  NAND U11116 ( .A(n10039), .B(n10038), .Z(n10062) );
  XOR U11117 ( .A(n10061), .B(n10062), .Z(n10064) );
  XOR U11118 ( .A(n10063), .B(n10064), .Z(n10052) );
  NANDN U11119 ( .A(n10041), .B(n10040), .Z(n10045) );
  OR U11120 ( .A(n10043), .B(n10042), .Z(n10044) );
  AND U11121 ( .A(n10045), .B(n10044), .Z(n10051) );
  XOR U11122 ( .A(n10052), .B(n10051), .Z(n10054) );
  XOR U11123 ( .A(n10053), .B(n10054), .Z(n10067) );
  XNOR U11124 ( .A(n10067), .B(sreg[1392]), .Z(n10069) );
  NANDN U11125 ( .A(n10046), .B(sreg[1391]), .Z(n10050) );
  NAND U11126 ( .A(n10048), .B(n10047), .Z(n10049) );
  NAND U11127 ( .A(n10050), .B(n10049), .Z(n10068) );
  XOR U11128 ( .A(n10069), .B(n10068), .Z(c[1392]) );
  NANDN U11129 ( .A(n10052), .B(n10051), .Z(n10056) );
  OR U11130 ( .A(n10054), .B(n10053), .Z(n10055) );
  AND U11131 ( .A(n10056), .B(n10055), .Z(n10074) );
  XOR U11132 ( .A(a[371]), .B(n2229), .Z(n10078) );
  AND U11133 ( .A(a[373]), .B(b[0]), .Z(n10058) );
  XNOR U11134 ( .A(n10058), .B(n2175), .Z(n10060) );
  NANDN U11135 ( .A(b[0]), .B(a[372]), .Z(n10059) );
  NAND U11136 ( .A(n10060), .B(n10059), .Z(n10083) );
  AND U11137 ( .A(a[369]), .B(b[3]), .Z(n10082) );
  XOR U11138 ( .A(n10083), .B(n10082), .Z(n10085) );
  XOR U11139 ( .A(n10084), .B(n10085), .Z(n10073) );
  NANDN U11140 ( .A(n10062), .B(n10061), .Z(n10066) );
  OR U11141 ( .A(n10064), .B(n10063), .Z(n10065) );
  AND U11142 ( .A(n10066), .B(n10065), .Z(n10072) );
  XOR U11143 ( .A(n10073), .B(n10072), .Z(n10075) );
  XOR U11144 ( .A(n10074), .B(n10075), .Z(n10088) );
  XNOR U11145 ( .A(n10088), .B(sreg[1393]), .Z(n10090) );
  NANDN U11146 ( .A(n10067), .B(sreg[1392]), .Z(n10071) );
  NAND U11147 ( .A(n10069), .B(n10068), .Z(n10070) );
  NAND U11148 ( .A(n10071), .B(n10070), .Z(n10089) );
  XOR U11149 ( .A(n10090), .B(n10089), .Z(c[1393]) );
  NANDN U11150 ( .A(n10073), .B(n10072), .Z(n10077) );
  OR U11151 ( .A(n10075), .B(n10074), .Z(n10076) );
  AND U11152 ( .A(n10077), .B(n10076), .Z(n10095) );
  XOR U11153 ( .A(a[372]), .B(n2229), .Z(n10099) );
  AND U11154 ( .A(a[374]), .B(b[0]), .Z(n10079) );
  XNOR U11155 ( .A(n10079), .B(n2175), .Z(n10081) );
  NANDN U11156 ( .A(b[0]), .B(a[373]), .Z(n10080) );
  NAND U11157 ( .A(n10081), .B(n10080), .Z(n10104) );
  AND U11158 ( .A(a[370]), .B(b[3]), .Z(n10103) );
  XOR U11159 ( .A(n10104), .B(n10103), .Z(n10106) );
  XOR U11160 ( .A(n10105), .B(n10106), .Z(n10094) );
  NANDN U11161 ( .A(n10083), .B(n10082), .Z(n10087) );
  OR U11162 ( .A(n10085), .B(n10084), .Z(n10086) );
  AND U11163 ( .A(n10087), .B(n10086), .Z(n10093) );
  XOR U11164 ( .A(n10094), .B(n10093), .Z(n10096) );
  XOR U11165 ( .A(n10095), .B(n10096), .Z(n10109) );
  XNOR U11166 ( .A(n10109), .B(sreg[1394]), .Z(n10111) );
  NANDN U11167 ( .A(n10088), .B(sreg[1393]), .Z(n10092) );
  NAND U11168 ( .A(n10090), .B(n10089), .Z(n10091) );
  NAND U11169 ( .A(n10092), .B(n10091), .Z(n10110) );
  XOR U11170 ( .A(n10111), .B(n10110), .Z(c[1394]) );
  NANDN U11171 ( .A(n10094), .B(n10093), .Z(n10098) );
  OR U11172 ( .A(n10096), .B(n10095), .Z(n10097) );
  AND U11173 ( .A(n10098), .B(n10097), .Z(n10116) );
  XOR U11174 ( .A(a[373]), .B(n2229), .Z(n10120) );
  AND U11175 ( .A(a[375]), .B(b[0]), .Z(n10100) );
  XNOR U11176 ( .A(n10100), .B(n2175), .Z(n10102) );
  NANDN U11177 ( .A(b[0]), .B(a[374]), .Z(n10101) );
  NAND U11178 ( .A(n10102), .B(n10101), .Z(n10125) );
  AND U11179 ( .A(a[371]), .B(b[3]), .Z(n10124) );
  XOR U11180 ( .A(n10125), .B(n10124), .Z(n10127) );
  XOR U11181 ( .A(n10126), .B(n10127), .Z(n10115) );
  NANDN U11182 ( .A(n10104), .B(n10103), .Z(n10108) );
  OR U11183 ( .A(n10106), .B(n10105), .Z(n10107) );
  AND U11184 ( .A(n10108), .B(n10107), .Z(n10114) );
  XOR U11185 ( .A(n10115), .B(n10114), .Z(n10117) );
  XOR U11186 ( .A(n10116), .B(n10117), .Z(n10130) );
  XNOR U11187 ( .A(n10130), .B(sreg[1395]), .Z(n10132) );
  NANDN U11188 ( .A(n10109), .B(sreg[1394]), .Z(n10113) );
  NAND U11189 ( .A(n10111), .B(n10110), .Z(n10112) );
  NAND U11190 ( .A(n10113), .B(n10112), .Z(n10131) );
  XOR U11191 ( .A(n10132), .B(n10131), .Z(c[1395]) );
  NANDN U11192 ( .A(n10115), .B(n10114), .Z(n10119) );
  OR U11193 ( .A(n10117), .B(n10116), .Z(n10118) );
  AND U11194 ( .A(n10119), .B(n10118), .Z(n10137) );
  XOR U11195 ( .A(a[374]), .B(n2229), .Z(n10141) );
  AND U11196 ( .A(a[376]), .B(b[0]), .Z(n10121) );
  XNOR U11197 ( .A(n10121), .B(n2175), .Z(n10123) );
  NANDN U11198 ( .A(b[0]), .B(a[375]), .Z(n10122) );
  NAND U11199 ( .A(n10123), .B(n10122), .Z(n10146) );
  AND U11200 ( .A(a[372]), .B(b[3]), .Z(n10145) );
  XOR U11201 ( .A(n10146), .B(n10145), .Z(n10148) );
  XOR U11202 ( .A(n10147), .B(n10148), .Z(n10136) );
  NANDN U11203 ( .A(n10125), .B(n10124), .Z(n10129) );
  OR U11204 ( .A(n10127), .B(n10126), .Z(n10128) );
  AND U11205 ( .A(n10129), .B(n10128), .Z(n10135) );
  XOR U11206 ( .A(n10136), .B(n10135), .Z(n10138) );
  XOR U11207 ( .A(n10137), .B(n10138), .Z(n10151) );
  XNOR U11208 ( .A(n10151), .B(sreg[1396]), .Z(n10153) );
  NANDN U11209 ( .A(n10130), .B(sreg[1395]), .Z(n10134) );
  NAND U11210 ( .A(n10132), .B(n10131), .Z(n10133) );
  NAND U11211 ( .A(n10134), .B(n10133), .Z(n10152) );
  XOR U11212 ( .A(n10153), .B(n10152), .Z(c[1396]) );
  NANDN U11213 ( .A(n10136), .B(n10135), .Z(n10140) );
  OR U11214 ( .A(n10138), .B(n10137), .Z(n10139) );
  AND U11215 ( .A(n10140), .B(n10139), .Z(n10158) );
  XOR U11216 ( .A(a[375]), .B(n2229), .Z(n10162) );
  AND U11217 ( .A(a[373]), .B(b[3]), .Z(n10166) );
  AND U11218 ( .A(a[377]), .B(b[0]), .Z(n10142) );
  XNOR U11219 ( .A(n10142), .B(n2175), .Z(n10144) );
  NANDN U11220 ( .A(b[0]), .B(a[376]), .Z(n10143) );
  NAND U11221 ( .A(n10144), .B(n10143), .Z(n10167) );
  XOR U11222 ( .A(n10166), .B(n10167), .Z(n10169) );
  XOR U11223 ( .A(n10168), .B(n10169), .Z(n10157) );
  NANDN U11224 ( .A(n10146), .B(n10145), .Z(n10150) );
  OR U11225 ( .A(n10148), .B(n10147), .Z(n10149) );
  AND U11226 ( .A(n10150), .B(n10149), .Z(n10156) );
  XOR U11227 ( .A(n10157), .B(n10156), .Z(n10159) );
  XOR U11228 ( .A(n10158), .B(n10159), .Z(n10172) );
  XNOR U11229 ( .A(n10172), .B(sreg[1397]), .Z(n10174) );
  NANDN U11230 ( .A(n10151), .B(sreg[1396]), .Z(n10155) );
  NAND U11231 ( .A(n10153), .B(n10152), .Z(n10154) );
  NAND U11232 ( .A(n10155), .B(n10154), .Z(n10173) );
  XOR U11233 ( .A(n10174), .B(n10173), .Z(c[1397]) );
  NANDN U11234 ( .A(n10157), .B(n10156), .Z(n10161) );
  OR U11235 ( .A(n10159), .B(n10158), .Z(n10160) );
  AND U11236 ( .A(n10161), .B(n10160), .Z(n10179) );
  XOR U11237 ( .A(a[376]), .B(n2229), .Z(n10183) );
  AND U11238 ( .A(a[378]), .B(b[0]), .Z(n10163) );
  XNOR U11239 ( .A(n10163), .B(n2175), .Z(n10165) );
  NANDN U11240 ( .A(b[0]), .B(a[377]), .Z(n10164) );
  NAND U11241 ( .A(n10165), .B(n10164), .Z(n10188) );
  AND U11242 ( .A(a[374]), .B(b[3]), .Z(n10187) );
  XOR U11243 ( .A(n10188), .B(n10187), .Z(n10190) );
  XOR U11244 ( .A(n10189), .B(n10190), .Z(n10178) );
  NANDN U11245 ( .A(n10167), .B(n10166), .Z(n10171) );
  OR U11246 ( .A(n10169), .B(n10168), .Z(n10170) );
  AND U11247 ( .A(n10171), .B(n10170), .Z(n10177) );
  XOR U11248 ( .A(n10178), .B(n10177), .Z(n10180) );
  XOR U11249 ( .A(n10179), .B(n10180), .Z(n10193) );
  XNOR U11250 ( .A(n10193), .B(sreg[1398]), .Z(n10195) );
  NANDN U11251 ( .A(n10172), .B(sreg[1397]), .Z(n10176) );
  NAND U11252 ( .A(n10174), .B(n10173), .Z(n10175) );
  NAND U11253 ( .A(n10176), .B(n10175), .Z(n10194) );
  XOR U11254 ( .A(n10195), .B(n10194), .Z(c[1398]) );
  NANDN U11255 ( .A(n10178), .B(n10177), .Z(n10182) );
  OR U11256 ( .A(n10180), .B(n10179), .Z(n10181) );
  AND U11257 ( .A(n10182), .B(n10181), .Z(n10200) );
  XOR U11258 ( .A(a[377]), .B(n2230), .Z(n10204) );
  AND U11259 ( .A(a[379]), .B(b[0]), .Z(n10184) );
  XNOR U11260 ( .A(n10184), .B(n2175), .Z(n10186) );
  NANDN U11261 ( .A(b[0]), .B(a[378]), .Z(n10185) );
  NAND U11262 ( .A(n10186), .B(n10185), .Z(n10209) );
  AND U11263 ( .A(a[375]), .B(b[3]), .Z(n10208) );
  XOR U11264 ( .A(n10209), .B(n10208), .Z(n10211) );
  XOR U11265 ( .A(n10210), .B(n10211), .Z(n10199) );
  NANDN U11266 ( .A(n10188), .B(n10187), .Z(n10192) );
  OR U11267 ( .A(n10190), .B(n10189), .Z(n10191) );
  AND U11268 ( .A(n10192), .B(n10191), .Z(n10198) );
  XOR U11269 ( .A(n10199), .B(n10198), .Z(n10201) );
  XOR U11270 ( .A(n10200), .B(n10201), .Z(n10214) );
  XNOR U11271 ( .A(n10214), .B(sreg[1399]), .Z(n10216) );
  NANDN U11272 ( .A(n10193), .B(sreg[1398]), .Z(n10197) );
  NAND U11273 ( .A(n10195), .B(n10194), .Z(n10196) );
  NAND U11274 ( .A(n10197), .B(n10196), .Z(n10215) );
  XOR U11275 ( .A(n10216), .B(n10215), .Z(c[1399]) );
  NANDN U11276 ( .A(n10199), .B(n10198), .Z(n10203) );
  OR U11277 ( .A(n10201), .B(n10200), .Z(n10202) );
  AND U11278 ( .A(n10203), .B(n10202), .Z(n10221) );
  XOR U11279 ( .A(a[378]), .B(n2230), .Z(n10225) );
  AND U11280 ( .A(a[376]), .B(b[3]), .Z(n10229) );
  AND U11281 ( .A(a[380]), .B(b[0]), .Z(n10205) );
  XNOR U11282 ( .A(n10205), .B(n2175), .Z(n10207) );
  NANDN U11283 ( .A(b[0]), .B(a[379]), .Z(n10206) );
  NAND U11284 ( .A(n10207), .B(n10206), .Z(n10230) );
  XOR U11285 ( .A(n10229), .B(n10230), .Z(n10232) );
  XOR U11286 ( .A(n10231), .B(n10232), .Z(n10220) );
  NANDN U11287 ( .A(n10209), .B(n10208), .Z(n10213) );
  OR U11288 ( .A(n10211), .B(n10210), .Z(n10212) );
  AND U11289 ( .A(n10213), .B(n10212), .Z(n10219) );
  XOR U11290 ( .A(n10220), .B(n10219), .Z(n10222) );
  XOR U11291 ( .A(n10221), .B(n10222), .Z(n10235) );
  XNOR U11292 ( .A(n10235), .B(sreg[1400]), .Z(n10237) );
  NANDN U11293 ( .A(n10214), .B(sreg[1399]), .Z(n10218) );
  NAND U11294 ( .A(n10216), .B(n10215), .Z(n10217) );
  NAND U11295 ( .A(n10218), .B(n10217), .Z(n10236) );
  XOR U11296 ( .A(n10237), .B(n10236), .Z(c[1400]) );
  NANDN U11297 ( .A(n10220), .B(n10219), .Z(n10224) );
  OR U11298 ( .A(n10222), .B(n10221), .Z(n10223) );
  AND U11299 ( .A(n10224), .B(n10223), .Z(n10242) );
  XOR U11300 ( .A(a[379]), .B(n2230), .Z(n10246) );
  AND U11301 ( .A(a[381]), .B(b[0]), .Z(n10226) );
  XNOR U11302 ( .A(n10226), .B(n2175), .Z(n10228) );
  NANDN U11303 ( .A(b[0]), .B(a[380]), .Z(n10227) );
  NAND U11304 ( .A(n10228), .B(n10227), .Z(n10251) );
  AND U11305 ( .A(a[377]), .B(b[3]), .Z(n10250) );
  XOR U11306 ( .A(n10251), .B(n10250), .Z(n10253) );
  XOR U11307 ( .A(n10252), .B(n10253), .Z(n10241) );
  NANDN U11308 ( .A(n10230), .B(n10229), .Z(n10234) );
  OR U11309 ( .A(n10232), .B(n10231), .Z(n10233) );
  AND U11310 ( .A(n10234), .B(n10233), .Z(n10240) );
  XOR U11311 ( .A(n10241), .B(n10240), .Z(n10243) );
  XOR U11312 ( .A(n10242), .B(n10243), .Z(n10256) );
  XNOR U11313 ( .A(n10256), .B(sreg[1401]), .Z(n10258) );
  NANDN U11314 ( .A(n10235), .B(sreg[1400]), .Z(n10239) );
  NAND U11315 ( .A(n10237), .B(n10236), .Z(n10238) );
  NAND U11316 ( .A(n10239), .B(n10238), .Z(n10257) );
  XOR U11317 ( .A(n10258), .B(n10257), .Z(c[1401]) );
  NANDN U11318 ( .A(n10241), .B(n10240), .Z(n10245) );
  OR U11319 ( .A(n10243), .B(n10242), .Z(n10244) );
  AND U11320 ( .A(n10245), .B(n10244), .Z(n10263) );
  XOR U11321 ( .A(a[380]), .B(n2230), .Z(n10267) );
  AND U11322 ( .A(a[378]), .B(b[3]), .Z(n10271) );
  AND U11323 ( .A(a[382]), .B(b[0]), .Z(n10247) );
  XNOR U11324 ( .A(n10247), .B(n2175), .Z(n10249) );
  NANDN U11325 ( .A(b[0]), .B(a[381]), .Z(n10248) );
  NAND U11326 ( .A(n10249), .B(n10248), .Z(n10272) );
  XOR U11327 ( .A(n10271), .B(n10272), .Z(n10274) );
  XOR U11328 ( .A(n10273), .B(n10274), .Z(n10262) );
  NANDN U11329 ( .A(n10251), .B(n10250), .Z(n10255) );
  OR U11330 ( .A(n10253), .B(n10252), .Z(n10254) );
  AND U11331 ( .A(n10255), .B(n10254), .Z(n10261) );
  XOR U11332 ( .A(n10262), .B(n10261), .Z(n10264) );
  XOR U11333 ( .A(n10263), .B(n10264), .Z(n10277) );
  XNOR U11334 ( .A(n10277), .B(sreg[1402]), .Z(n10279) );
  NANDN U11335 ( .A(n10256), .B(sreg[1401]), .Z(n10260) );
  NAND U11336 ( .A(n10258), .B(n10257), .Z(n10259) );
  NAND U11337 ( .A(n10260), .B(n10259), .Z(n10278) );
  XOR U11338 ( .A(n10279), .B(n10278), .Z(c[1402]) );
  NANDN U11339 ( .A(n10262), .B(n10261), .Z(n10266) );
  OR U11340 ( .A(n10264), .B(n10263), .Z(n10265) );
  AND U11341 ( .A(n10266), .B(n10265), .Z(n10284) );
  XOR U11342 ( .A(a[381]), .B(n2230), .Z(n10288) );
  AND U11343 ( .A(a[383]), .B(b[0]), .Z(n10268) );
  XNOR U11344 ( .A(n10268), .B(n2175), .Z(n10270) );
  NANDN U11345 ( .A(b[0]), .B(a[382]), .Z(n10269) );
  NAND U11346 ( .A(n10270), .B(n10269), .Z(n10293) );
  AND U11347 ( .A(a[379]), .B(b[3]), .Z(n10292) );
  XOR U11348 ( .A(n10293), .B(n10292), .Z(n10295) );
  XOR U11349 ( .A(n10294), .B(n10295), .Z(n10283) );
  NANDN U11350 ( .A(n10272), .B(n10271), .Z(n10276) );
  OR U11351 ( .A(n10274), .B(n10273), .Z(n10275) );
  AND U11352 ( .A(n10276), .B(n10275), .Z(n10282) );
  XOR U11353 ( .A(n10283), .B(n10282), .Z(n10285) );
  XOR U11354 ( .A(n10284), .B(n10285), .Z(n10298) );
  XNOR U11355 ( .A(n10298), .B(sreg[1403]), .Z(n10300) );
  NANDN U11356 ( .A(n10277), .B(sreg[1402]), .Z(n10281) );
  NAND U11357 ( .A(n10279), .B(n10278), .Z(n10280) );
  NAND U11358 ( .A(n10281), .B(n10280), .Z(n10299) );
  XOR U11359 ( .A(n10300), .B(n10299), .Z(c[1403]) );
  NANDN U11360 ( .A(n10283), .B(n10282), .Z(n10287) );
  OR U11361 ( .A(n10285), .B(n10284), .Z(n10286) );
  AND U11362 ( .A(n10287), .B(n10286), .Z(n10305) );
  XOR U11363 ( .A(a[382]), .B(n2230), .Z(n10309) );
  AND U11364 ( .A(a[380]), .B(b[3]), .Z(n10313) );
  AND U11365 ( .A(a[384]), .B(b[0]), .Z(n10289) );
  XNOR U11366 ( .A(n10289), .B(n2175), .Z(n10291) );
  NANDN U11367 ( .A(b[0]), .B(a[383]), .Z(n10290) );
  NAND U11368 ( .A(n10291), .B(n10290), .Z(n10314) );
  XOR U11369 ( .A(n10313), .B(n10314), .Z(n10316) );
  XOR U11370 ( .A(n10315), .B(n10316), .Z(n10304) );
  NANDN U11371 ( .A(n10293), .B(n10292), .Z(n10297) );
  OR U11372 ( .A(n10295), .B(n10294), .Z(n10296) );
  AND U11373 ( .A(n10297), .B(n10296), .Z(n10303) );
  XOR U11374 ( .A(n10304), .B(n10303), .Z(n10306) );
  XOR U11375 ( .A(n10305), .B(n10306), .Z(n10319) );
  XNOR U11376 ( .A(n10319), .B(sreg[1404]), .Z(n10321) );
  NANDN U11377 ( .A(n10298), .B(sreg[1403]), .Z(n10302) );
  NAND U11378 ( .A(n10300), .B(n10299), .Z(n10301) );
  NAND U11379 ( .A(n10302), .B(n10301), .Z(n10320) );
  XOR U11380 ( .A(n10321), .B(n10320), .Z(c[1404]) );
  NANDN U11381 ( .A(n10304), .B(n10303), .Z(n10308) );
  OR U11382 ( .A(n10306), .B(n10305), .Z(n10307) );
  AND U11383 ( .A(n10308), .B(n10307), .Z(n10326) );
  XOR U11384 ( .A(a[383]), .B(n2230), .Z(n10330) );
  AND U11385 ( .A(a[385]), .B(b[0]), .Z(n10310) );
  XNOR U11386 ( .A(n10310), .B(n2175), .Z(n10312) );
  NANDN U11387 ( .A(b[0]), .B(a[384]), .Z(n10311) );
  NAND U11388 ( .A(n10312), .B(n10311), .Z(n10335) );
  AND U11389 ( .A(a[381]), .B(b[3]), .Z(n10334) );
  XOR U11390 ( .A(n10335), .B(n10334), .Z(n10337) );
  XOR U11391 ( .A(n10336), .B(n10337), .Z(n10325) );
  NANDN U11392 ( .A(n10314), .B(n10313), .Z(n10318) );
  OR U11393 ( .A(n10316), .B(n10315), .Z(n10317) );
  AND U11394 ( .A(n10318), .B(n10317), .Z(n10324) );
  XOR U11395 ( .A(n10325), .B(n10324), .Z(n10327) );
  XOR U11396 ( .A(n10326), .B(n10327), .Z(n10340) );
  XNOR U11397 ( .A(n10340), .B(sreg[1405]), .Z(n10342) );
  NANDN U11398 ( .A(n10319), .B(sreg[1404]), .Z(n10323) );
  NAND U11399 ( .A(n10321), .B(n10320), .Z(n10322) );
  NAND U11400 ( .A(n10323), .B(n10322), .Z(n10341) );
  XOR U11401 ( .A(n10342), .B(n10341), .Z(c[1405]) );
  NANDN U11402 ( .A(n10325), .B(n10324), .Z(n10329) );
  OR U11403 ( .A(n10327), .B(n10326), .Z(n10328) );
  AND U11404 ( .A(n10329), .B(n10328), .Z(n10347) );
  XOR U11405 ( .A(a[384]), .B(n2231), .Z(n10351) );
  AND U11406 ( .A(a[382]), .B(b[3]), .Z(n10355) );
  AND U11407 ( .A(a[386]), .B(b[0]), .Z(n10331) );
  XNOR U11408 ( .A(n10331), .B(n2175), .Z(n10333) );
  NANDN U11409 ( .A(b[0]), .B(a[385]), .Z(n10332) );
  NAND U11410 ( .A(n10333), .B(n10332), .Z(n10356) );
  XOR U11411 ( .A(n10355), .B(n10356), .Z(n10358) );
  XOR U11412 ( .A(n10357), .B(n10358), .Z(n10346) );
  NANDN U11413 ( .A(n10335), .B(n10334), .Z(n10339) );
  OR U11414 ( .A(n10337), .B(n10336), .Z(n10338) );
  AND U11415 ( .A(n10339), .B(n10338), .Z(n10345) );
  XOR U11416 ( .A(n10346), .B(n10345), .Z(n10348) );
  XOR U11417 ( .A(n10347), .B(n10348), .Z(n10361) );
  XNOR U11418 ( .A(n10361), .B(sreg[1406]), .Z(n10363) );
  NANDN U11419 ( .A(n10340), .B(sreg[1405]), .Z(n10344) );
  NAND U11420 ( .A(n10342), .B(n10341), .Z(n10343) );
  NAND U11421 ( .A(n10344), .B(n10343), .Z(n10362) );
  XOR U11422 ( .A(n10363), .B(n10362), .Z(c[1406]) );
  NANDN U11423 ( .A(n10346), .B(n10345), .Z(n10350) );
  OR U11424 ( .A(n10348), .B(n10347), .Z(n10349) );
  AND U11425 ( .A(n10350), .B(n10349), .Z(n10368) );
  XOR U11426 ( .A(a[385]), .B(n2231), .Z(n10372) );
  AND U11427 ( .A(a[387]), .B(b[0]), .Z(n10352) );
  XNOR U11428 ( .A(n10352), .B(n2175), .Z(n10354) );
  NANDN U11429 ( .A(b[0]), .B(a[386]), .Z(n10353) );
  NAND U11430 ( .A(n10354), .B(n10353), .Z(n10377) );
  AND U11431 ( .A(a[383]), .B(b[3]), .Z(n10376) );
  XOR U11432 ( .A(n10377), .B(n10376), .Z(n10379) );
  XOR U11433 ( .A(n10378), .B(n10379), .Z(n10367) );
  NANDN U11434 ( .A(n10356), .B(n10355), .Z(n10360) );
  OR U11435 ( .A(n10358), .B(n10357), .Z(n10359) );
  AND U11436 ( .A(n10360), .B(n10359), .Z(n10366) );
  XOR U11437 ( .A(n10367), .B(n10366), .Z(n10369) );
  XOR U11438 ( .A(n10368), .B(n10369), .Z(n10382) );
  XNOR U11439 ( .A(n10382), .B(sreg[1407]), .Z(n10384) );
  NANDN U11440 ( .A(n10361), .B(sreg[1406]), .Z(n10365) );
  NAND U11441 ( .A(n10363), .B(n10362), .Z(n10364) );
  NAND U11442 ( .A(n10365), .B(n10364), .Z(n10383) );
  XOR U11443 ( .A(n10384), .B(n10383), .Z(c[1407]) );
  NANDN U11444 ( .A(n10367), .B(n10366), .Z(n10371) );
  OR U11445 ( .A(n10369), .B(n10368), .Z(n10370) );
  AND U11446 ( .A(n10371), .B(n10370), .Z(n10389) );
  XOR U11447 ( .A(a[386]), .B(n2231), .Z(n10393) );
  AND U11448 ( .A(a[384]), .B(b[3]), .Z(n10397) );
  AND U11449 ( .A(a[388]), .B(b[0]), .Z(n10373) );
  XNOR U11450 ( .A(n10373), .B(n2175), .Z(n10375) );
  NANDN U11451 ( .A(b[0]), .B(a[387]), .Z(n10374) );
  NAND U11452 ( .A(n10375), .B(n10374), .Z(n10398) );
  XOR U11453 ( .A(n10397), .B(n10398), .Z(n10400) );
  XOR U11454 ( .A(n10399), .B(n10400), .Z(n10388) );
  NANDN U11455 ( .A(n10377), .B(n10376), .Z(n10381) );
  OR U11456 ( .A(n10379), .B(n10378), .Z(n10380) );
  AND U11457 ( .A(n10381), .B(n10380), .Z(n10387) );
  XOR U11458 ( .A(n10388), .B(n10387), .Z(n10390) );
  XOR U11459 ( .A(n10389), .B(n10390), .Z(n10403) );
  XNOR U11460 ( .A(n10403), .B(sreg[1408]), .Z(n10405) );
  NANDN U11461 ( .A(n10382), .B(sreg[1407]), .Z(n10386) );
  NAND U11462 ( .A(n10384), .B(n10383), .Z(n10385) );
  NAND U11463 ( .A(n10386), .B(n10385), .Z(n10404) );
  XOR U11464 ( .A(n10405), .B(n10404), .Z(c[1408]) );
  NANDN U11465 ( .A(n10388), .B(n10387), .Z(n10392) );
  OR U11466 ( .A(n10390), .B(n10389), .Z(n10391) );
  AND U11467 ( .A(n10392), .B(n10391), .Z(n10410) );
  XOR U11468 ( .A(a[387]), .B(n2231), .Z(n10414) );
  AND U11469 ( .A(a[389]), .B(b[0]), .Z(n10394) );
  XNOR U11470 ( .A(n10394), .B(n2175), .Z(n10396) );
  NANDN U11471 ( .A(b[0]), .B(a[388]), .Z(n10395) );
  NAND U11472 ( .A(n10396), .B(n10395), .Z(n10419) );
  AND U11473 ( .A(a[385]), .B(b[3]), .Z(n10418) );
  XOR U11474 ( .A(n10419), .B(n10418), .Z(n10421) );
  XOR U11475 ( .A(n10420), .B(n10421), .Z(n10409) );
  NANDN U11476 ( .A(n10398), .B(n10397), .Z(n10402) );
  OR U11477 ( .A(n10400), .B(n10399), .Z(n10401) );
  AND U11478 ( .A(n10402), .B(n10401), .Z(n10408) );
  XOR U11479 ( .A(n10409), .B(n10408), .Z(n10411) );
  XOR U11480 ( .A(n10410), .B(n10411), .Z(n10424) );
  XNOR U11481 ( .A(n10424), .B(sreg[1409]), .Z(n10426) );
  NANDN U11482 ( .A(n10403), .B(sreg[1408]), .Z(n10407) );
  NAND U11483 ( .A(n10405), .B(n10404), .Z(n10406) );
  NAND U11484 ( .A(n10407), .B(n10406), .Z(n10425) );
  XOR U11485 ( .A(n10426), .B(n10425), .Z(c[1409]) );
  NANDN U11486 ( .A(n10409), .B(n10408), .Z(n10413) );
  OR U11487 ( .A(n10411), .B(n10410), .Z(n10412) );
  AND U11488 ( .A(n10413), .B(n10412), .Z(n10431) );
  XOR U11489 ( .A(a[388]), .B(n2231), .Z(n10435) );
  AND U11490 ( .A(a[390]), .B(b[0]), .Z(n10415) );
  XNOR U11491 ( .A(n10415), .B(n2175), .Z(n10417) );
  NANDN U11492 ( .A(b[0]), .B(a[389]), .Z(n10416) );
  NAND U11493 ( .A(n10417), .B(n10416), .Z(n10440) );
  AND U11494 ( .A(a[386]), .B(b[3]), .Z(n10439) );
  XOR U11495 ( .A(n10440), .B(n10439), .Z(n10442) );
  XOR U11496 ( .A(n10441), .B(n10442), .Z(n10430) );
  NANDN U11497 ( .A(n10419), .B(n10418), .Z(n10423) );
  OR U11498 ( .A(n10421), .B(n10420), .Z(n10422) );
  AND U11499 ( .A(n10423), .B(n10422), .Z(n10429) );
  XOR U11500 ( .A(n10430), .B(n10429), .Z(n10432) );
  XOR U11501 ( .A(n10431), .B(n10432), .Z(n10445) );
  XNOR U11502 ( .A(n10445), .B(sreg[1410]), .Z(n10447) );
  NANDN U11503 ( .A(n10424), .B(sreg[1409]), .Z(n10428) );
  NAND U11504 ( .A(n10426), .B(n10425), .Z(n10427) );
  NAND U11505 ( .A(n10428), .B(n10427), .Z(n10446) );
  XOR U11506 ( .A(n10447), .B(n10446), .Z(c[1410]) );
  NANDN U11507 ( .A(n10430), .B(n10429), .Z(n10434) );
  OR U11508 ( .A(n10432), .B(n10431), .Z(n10433) );
  AND U11509 ( .A(n10434), .B(n10433), .Z(n10452) );
  XOR U11510 ( .A(a[389]), .B(n2231), .Z(n10456) );
  AND U11511 ( .A(a[391]), .B(b[0]), .Z(n10436) );
  XNOR U11512 ( .A(n10436), .B(n2175), .Z(n10438) );
  NANDN U11513 ( .A(b[0]), .B(a[390]), .Z(n10437) );
  NAND U11514 ( .A(n10438), .B(n10437), .Z(n10461) );
  AND U11515 ( .A(a[387]), .B(b[3]), .Z(n10460) );
  XOR U11516 ( .A(n10461), .B(n10460), .Z(n10463) );
  XOR U11517 ( .A(n10462), .B(n10463), .Z(n10451) );
  NANDN U11518 ( .A(n10440), .B(n10439), .Z(n10444) );
  OR U11519 ( .A(n10442), .B(n10441), .Z(n10443) );
  AND U11520 ( .A(n10444), .B(n10443), .Z(n10450) );
  XOR U11521 ( .A(n10451), .B(n10450), .Z(n10453) );
  XOR U11522 ( .A(n10452), .B(n10453), .Z(n10466) );
  XNOR U11523 ( .A(n10466), .B(sreg[1411]), .Z(n10468) );
  NANDN U11524 ( .A(n10445), .B(sreg[1410]), .Z(n10449) );
  NAND U11525 ( .A(n10447), .B(n10446), .Z(n10448) );
  NAND U11526 ( .A(n10449), .B(n10448), .Z(n10467) );
  XOR U11527 ( .A(n10468), .B(n10467), .Z(c[1411]) );
  NANDN U11528 ( .A(n10451), .B(n10450), .Z(n10455) );
  OR U11529 ( .A(n10453), .B(n10452), .Z(n10454) );
  AND U11530 ( .A(n10455), .B(n10454), .Z(n10473) );
  XOR U11531 ( .A(a[390]), .B(n2231), .Z(n10477) );
  AND U11532 ( .A(a[388]), .B(b[3]), .Z(n10481) );
  AND U11533 ( .A(a[392]), .B(b[0]), .Z(n10457) );
  XNOR U11534 ( .A(n10457), .B(n2175), .Z(n10459) );
  NANDN U11535 ( .A(b[0]), .B(a[391]), .Z(n10458) );
  NAND U11536 ( .A(n10459), .B(n10458), .Z(n10482) );
  XOR U11537 ( .A(n10481), .B(n10482), .Z(n10484) );
  XOR U11538 ( .A(n10483), .B(n10484), .Z(n10472) );
  NANDN U11539 ( .A(n10461), .B(n10460), .Z(n10465) );
  OR U11540 ( .A(n10463), .B(n10462), .Z(n10464) );
  AND U11541 ( .A(n10465), .B(n10464), .Z(n10471) );
  XOR U11542 ( .A(n10472), .B(n10471), .Z(n10474) );
  XOR U11543 ( .A(n10473), .B(n10474), .Z(n10487) );
  XNOR U11544 ( .A(n10487), .B(sreg[1412]), .Z(n10489) );
  NANDN U11545 ( .A(n10466), .B(sreg[1411]), .Z(n10470) );
  NAND U11546 ( .A(n10468), .B(n10467), .Z(n10469) );
  NAND U11547 ( .A(n10470), .B(n10469), .Z(n10488) );
  XOR U11548 ( .A(n10489), .B(n10488), .Z(c[1412]) );
  NANDN U11549 ( .A(n10472), .B(n10471), .Z(n10476) );
  OR U11550 ( .A(n10474), .B(n10473), .Z(n10475) );
  AND U11551 ( .A(n10476), .B(n10475), .Z(n10494) );
  XOR U11552 ( .A(a[391]), .B(n2232), .Z(n10498) );
  AND U11553 ( .A(a[393]), .B(b[0]), .Z(n10478) );
  XNOR U11554 ( .A(n10478), .B(n2175), .Z(n10480) );
  NANDN U11555 ( .A(b[0]), .B(a[392]), .Z(n10479) );
  NAND U11556 ( .A(n10480), .B(n10479), .Z(n10503) );
  AND U11557 ( .A(a[389]), .B(b[3]), .Z(n10502) );
  XOR U11558 ( .A(n10503), .B(n10502), .Z(n10505) );
  XOR U11559 ( .A(n10504), .B(n10505), .Z(n10493) );
  NANDN U11560 ( .A(n10482), .B(n10481), .Z(n10486) );
  OR U11561 ( .A(n10484), .B(n10483), .Z(n10485) );
  AND U11562 ( .A(n10486), .B(n10485), .Z(n10492) );
  XOR U11563 ( .A(n10493), .B(n10492), .Z(n10495) );
  XOR U11564 ( .A(n10494), .B(n10495), .Z(n10508) );
  XNOR U11565 ( .A(n10508), .B(sreg[1413]), .Z(n10510) );
  NANDN U11566 ( .A(n10487), .B(sreg[1412]), .Z(n10491) );
  NAND U11567 ( .A(n10489), .B(n10488), .Z(n10490) );
  NAND U11568 ( .A(n10491), .B(n10490), .Z(n10509) );
  XOR U11569 ( .A(n10510), .B(n10509), .Z(c[1413]) );
  NANDN U11570 ( .A(n10493), .B(n10492), .Z(n10497) );
  OR U11571 ( .A(n10495), .B(n10494), .Z(n10496) );
  AND U11572 ( .A(n10497), .B(n10496), .Z(n10515) );
  XOR U11573 ( .A(a[392]), .B(n2232), .Z(n10519) );
  AND U11574 ( .A(a[390]), .B(b[3]), .Z(n10523) );
  AND U11575 ( .A(a[394]), .B(b[0]), .Z(n10499) );
  XNOR U11576 ( .A(n10499), .B(n2175), .Z(n10501) );
  NANDN U11577 ( .A(b[0]), .B(a[393]), .Z(n10500) );
  NAND U11578 ( .A(n10501), .B(n10500), .Z(n10524) );
  XOR U11579 ( .A(n10523), .B(n10524), .Z(n10526) );
  XOR U11580 ( .A(n10525), .B(n10526), .Z(n10514) );
  NANDN U11581 ( .A(n10503), .B(n10502), .Z(n10507) );
  OR U11582 ( .A(n10505), .B(n10504), .Z(n10506) );
  AND U11583 ( .A(n10507), .B(n10506), .Z(n10513) );
  XOR U11584 ( .A(n10514), .B(n10513), .Z(n10516) );
  XOR U11585 ( .A(n10515), .B(n10516), .Z(n10529) );
  XNOR U11586 ( .A(n10529), .B(sreg[1414]), .Z(n10531) );
  NANDN U11587 ( .A(n10508), .B(sreg[1413]), .Z(n10512) );
  NAND U11588 ( .A(n10510), .B(n10509), .Z(n10511) );
  NAND U11589 ( .A(n10512), .B(n10511), .Z(n10530) );
  XOR U11590 ( .A(n10531), .B(n10530), .Z(c[1414]) );
  NANDN U11591 ( .A(n10514), .B(n10513), .Z(n10518) );
  OR U11592 ( .A(n10516), .B(n10515), .Z(n10517) );
  AND U11593 ( .A(n10518), .B(n10517), .Z(n10536) );
  XOR U11594 ( .A(a[393]), .B(n2232), .Z(n10540) );
  AND U11595 ( .A(a[395]), .B(b[0]), .Z(n10520) );
  XNOR U11596 ( .A(n10520), .B(n2175), .Z(n10522) );
  NANDN U11597 ( .A(b[0]), .B(a[394]), .Z(n10521) );
  NAND U11598 ( .A(n10522), .B(n10521), .Z(n10545) );
  AND U11599 ( .A(a[391]), .B(b[3]), .Z(n10544) );
  XOR U11600 ( .A(n10545), .B(n10544), .Z(n10547) );
  XOR U11601 ( .A(n10546), .B(n10547), .Z(n10535) );
  NANDN U11602 ( .A(n10524), .B(n10523), .Z(n10528) );
  OR U11603 ( .A(n10526), .B(n10525), .Z(n10527) );
  AND U11604 ( .A(n10528), .B(n10527), .Z(n10534) );
  XOR U11605 ( .A(n10535), .B(n10534), .Z(n10537) );
  XOR U11606 ( .A(n10536), .B(n10537), .Z(n10550) );
  XNOR U11607 ( .A(n10550), .B(sreg[1415]), .Z(n10552) );
  NANDN U11608 ( .A(n10529), .B(sreg[1414]), .Z(n10533) );
  NAND U11609 ( .A(n10531), .B(n10530), .Z(n10532) );
  NAND U11610 ( .A(n10533), .B(n10532), .Z(n10551) );
  XOR U11611 ( .A(n10552), .B(n10551), .Z(c[1415]) );
  NANDN U11612 ( .A(n10535), .B(n10534), .Z(n10539) );
  OR U11613 ( .A(n10537), .B(n10536), .Z(n10538) );
  AND U11614 ( .A(n10539), .B(n10538), .Z(n10557) );
  XOR U11615 ( .A(a[394]), .B(n2232), .Z(n10561) );
  AND U11616 ( .A(a[396]), .B(b[0]), .Z(n10541) );
  XNOR U11617 ( .A(n10541), .B(n2175), .Z(n10543) );
  NANDN U11618 ( .A(b[0]), .B(a[395]), .Z(n10542) );
  NAND U11619 ( .A(n10543), .B(n10542), .Z(n10566) );
  AND U11620 ( .A(a[392]), .B(b[3]), .Z(n10565) );
  XOR U11621 ( .A(n10566), .B(n10565), .Z(n10568) );
  XOR U11622 ( .A(n10567), .B(n10568), .Z(n10556) );
  NANDN U11623 ( .A(n10545), .B(n10544), .Z(n10549) );
  OR U11624 ( .A(n10547), .B(n10546), .Z(n10548) );
  AND U11625 ( .A(n10549), .B(n10548), .Z(n10555) );
  XOR U11626 ( .A(n10556), .B(n10555), .Z(n10558) );
  XOR U11627 ( .A(n10557), .B(n10558), .Z(n10571) );
  XNOR U11628 ( .A(n10571), .B(sreg[1416]), .Z(n10573) );
  NANDN U11629 ( .A(n10550), .B(sreg[1415]), .Z(n10554) );
  NAND U11630 ( .A(n10552), .B(n10551), .Z(n10553) );
  NAND U11631 ( .A(n10554), .B(n10553), .Z(n10572) );
  XOR U11632 ( .A(n10573), .B(n10572), .Z(c[1416]) );
  NANDN U11633 ( .A(n10556), .B(n10555), .Z(n10560) );
  OR U11634 ( .A(n10558), .B(n10557), .Z(n10559) );
  AND U11635 ( .A(n10560), .B(n10559), .Z(n10578) );
  XOR U11636 ( .A(a[395]), .B(n2232), .Z(n10582) );
  AND U11637 ( .A(a[397]), .B(b[0]), .Z(n10562) );
  XNOR U11638 ( .A(n10562), .B(n2175), .Z(n10564) );
  NANDN U11639 ( .A(b[0]), .B(a[396]), .Z(n10563) );
  NAND U11640 ( .A(n10564), .B(n10563), .Z(n10587) );
  AND U11641 ( .A(a[393]), .B(b[3]), .Z(n10586) );
  XOR U11642 ( .A(n10587), .B(n10586), .Z(n10589) );
  XOR U11643 ( .A(n10588), .B(n10589), .Z(n10577) );
  NANDN U11644 ( .A(n10566), .B(n10565), .Z(n10570) );
  OR U11645 ( .A(n10568), .B(n10567), .Z(n10569) );
  AND U11646 ( .A(n10570), .B(n10569), .Z(n10576) );
  XOR U11647 ( .A(n10577), .B(n10576), .Z(n10579) );
  XOR U11648 ( .A(n10578), .B(n10579), .Z(n10592) );
  XNOR U11649 ( .A(n10592), .B(sreg[1417]), .Z(n10594) );
  NANDN U11650 ( .A(n10571), .B(sreg[1416]), .Z(n10575) );
  NAND U11651 ( .A(n10573), .B(n10572), .Z(n10574) );
  NAND U11652 ( .A(n10575), .B(n10574), .Z(n10593) );
  XOR U11653 ( .A(n10594), .B(n10593), .Z(c[1417]) );
  NANDN U11654 ( .A(n10577), .B(n10576), .Z(n10581) );
  OR U11655 ( .A(n10579), .B(n10578), .Z(n10580) );
  AND U11656 ( .A(n10581), .B(n10580), .Z(n10599) );
  XOR U11657 ( .A(a[396]), .B(n2232), .Z(n10603) );
  AND U11658 ( .A(a[394]), .B(b[3]), .Z(n10607) );
  AND U11659 ( .A(a[398]), .B(b[0]), .Z(n10583) );
  XNOR U11660 ( .A(n10583), .B(n2175), .Z(n10585) );
  NANDN U11661 ( .A(b[0]), .B(a[397]), .Z(n10584) );
  NAND U11662 ( .A(n10585), .B(n10584), .Z(n10608) );
  XOR U11663 ( .A(n10607), .B(n10608), .Z(n10610) );
  XOR U11664 ( .A(n10609), .B(n10610), .Z(n10598) );
  NANDN U11665 ( .A(n10587), .B(n10586), .Z(n10591) );
  OR U11666 ( .A(n10589), .B(n10588), .Z(n10590) );
  AND U11667 ( .A(n10591), .B(n10590), .Z(n10597) );
  XOR U11668 ( .A(n10598), .B(n10597), .Z(n10600) );
  XOR U11669 ( .A(n10599), .B(n10600), .Z(n10613) );
  XNOR U11670 ( .A(n10613), .B(sreg[1418]), .Z(n10615) );
  NANDN U11671 ( .A(n10592), .B(sreg[1417]), .Z(n10596) );
  NAND U11672 ( .A(n10594), .B(n10593), .Z(n10595) );
  NAND U11673 ( .A(n10596), .B(n10595), .Z(n10614) );
  XOR U11674 ( .A(n10615), .B(n10614), .Z(c[1418]) );
  NANDN U11675 ( .A(n10598), .B(n10597), .Z(n10602) );
  OR U11676 ( .A(n10600), .B(n10599), .Z(n10601) );
  AND U11677 ( .A(n10602), .B(n10601), .Z(n10620) );
  XOR U11678 ( .A(a[397]), .B(n2232), .Z(n10624) );
  AND U11679 ( .A(a[395]), .B(b[3]), .Z(n10628) );
  AND U11680 ( .A(a[399]), .B(b[0]), .Z(n10604) );
  XNOR U11681 ( .A(n10604), .B(n2175), .Z(n10606) );
  NANDN U11682 ( .A(b[0]), .B(a[398]), .Z(n10605) );
  NAND U11683 ( .A(n10606), .B(n10605), .Z(n10629) );
  XOR U11684 ( .A(n10628), .B(n10629), .Z(n10631) );
  XOR U11685 ( .A(n10630), .B(n10631), .Z(n10619) );
  NANDN U11686 ( .A(n10608), .B(n10607), .Z(n10612) );
  OR U11687 ( .A(n10610), .B(n10609), .Z(n10611) );
  AND U11688 ( .A(n10612), .B(n10611), .Z(n10618) );
  XOR U11689 ( .A(n10619), .B(n10618), .Z(n10621) );
  XOR U11690 ( .A(n10620), .B(n10621), .Z(n10634) );
  XNOR U11691 ( .A(n10634), .B(sreg[1419]), .Z(n10636) );
  NANDN U11692 ( .A(n10613), .B(sreg[1418]), .Z(n10617) );
  NAND U11693 ( .A(n10615), .B(n10614), .Z(n10616) );
  NAND U11694 ( .A(n10617), .B(n10616), .Z(n10635) );
  XOR U11695 ( .A(n10636), .B(n10635), .Z(c[1419]) );
  NANDN U11696 ( .A(n10619), .B(n10618), .Z(n10623) );
  OR U11697 ( .A(n10621), .B(n10620), .Z(n10622) );
  AND U11698 ( .A(n10623), .B(n10622), .Z(n10641) );
  XOR U11699 ( .A(a[398]), .B(n2233), .Z(n10645) );
  AND U11700 ( .A(a[400]), .B(b[0]), .Z(n10625) );
  XNOR U11701 ( .A(n10625), .B(n2175), .Z(n10627) );
  NANDN U11702 ( .A(b[0]), .B(a[399]), .Z(n10626) );
  NAND U11703 ( .A(n10627), .B(n10626), .Z(n10650) );
  AND U11704 ( .A(a[396]), .B(b[3]), .Z(n10649) );
  XOR U11705 ( .A(n10650), .B(n10649), .Z(n10652) );
  XOR U11706 ( .A(n10651), .B(n10652), .Z(n10640) );
  NANDN U11707 ( .A(n10629), .B(n10628), .Z(n10633) );
  OR U11708 ( .A(n10631), .B(n10630), .Z(n10632) );
  AND U11709 ( .A(n10633), .B(n10632), .Z(n10639) );
  XOR U11710 ( .A(n10640), .B(n10639), .Z(n10642) );
  XOR U11711 ( .A(n10641), .B(n10642), .Z(n10655) );
  XNOR U11712 ( .A(n10655), .B(sreg[1420]), .Z(n10657) );
  NANDN U11713 ( .A(n10634), .B(sreg[1419]), .Z(n10638) );
  NAND U11714 ( .A(n10636), .B(n10635), .Z(n10637) );
  NAND U11715 ( .A(n10638), .B(n10637), .Z(n10656) );
  XOR U11716 ( .A(n10657), .B(n10656), .Z(c[1420]) );
  NANDN U11717 ( .A(n10640), .B(n10639), .Z(n10644) );
  OR U11718 ( .A(n10642), .B(n10641), .Z(n10643) );
  AND U11719 ( .A(n10644), .B(n10643), .Z(n10662) );
  XOR U11720 ( .A(a[399]), .B(n2233), .Z(n10666) );
  AND U11721 ( .A(a[401]), .B(b[0]), .Z(n10646) );
  XNOR U11722 ( .A(n10646), .B(n2175), .Z(n10648) );
  NANDN U11723 ( .A(b[0]), .B(a[400]), .Z(n10647) );
  NAND U11724 ( .A(n10648), .B(n10647), .Z(n10671) );
  AND U11725 ( .A(a[397]), .B(b[3]), .Z(n10670) );
  XOR U11726 ( .A(n10671), .B(n10670), .Z(n10673) );
  XOR U11727 ( .A(n10672), .B(n10673), .Z(n10661) );
  NANDN U11728 ( .A(n10650), .B(n10649), .Z(n10654) );
  OR U11729 ( .A(n10652), .B(n10651), .Z(n10653) );
  AND U11730 ( .A(n10654), .B(n10653), .Z(n10660) );
  XOR U11731 ( .A(n10661), .B(n10660), .Z(n10663) );
  XOR U11732 ( .A(n10662), .B(n10663), .Z(n10676) );
  XNOR U11733 ( .A(n10676), .B(sreg[1421]), .Z(n10678) );
  NANDN U11734 ( .A(n10655), .B(sreg[1420]), .Z(n10659) );
  NAND U11735 ( .A(n10657), .B(n10656), .Z(n10658) );
  NAND U11736 ( .A(n10659), .B(n10658), .Z(n10677) );
  XOR U11737 ( .A(n10678), .B(n10677), .Z(c[1421]) );
  NANDN U11738 ( .A(n10661), .B(n10660), .Z(n10665) );
  OR U11739 ( .A(n10663), .B(n10662), .Z(n10664) );
  AND U11740 ( .A(n10665), .B(n10664), .Z(n10683) );
  XOR U11741 ( .A(a[400]), .B(n2233), .Z(n10687) );
  AND U11742 ( .A(a[402]), .B(b[0]), .Z(n10667) );
  XNOR U11743 ( .A(n10667), .B(n2175), .Z(n10669) );
  NANDN U11744 ( .A(b[0]), .B(a[401]), .Z(n10668) );
  NAND U11745 ( .A(n10669), .B(n10668), .Z(n10692) );
  AND U11746 ( .A(a[398]), .B(b[3]), .Z(n10691) );
  XOR U11747 ( .A(n10692), .B(n10691), .Z(n10694) );
  XOR U11748 ( .A(n10693), .B(n10694), .Z(n10682) );
  NANDN U11749 ( .A(n10671), .B(n10670), .Z(n10675) );
  OR U11750 ( .A(n10673), .B(n10672), .Z(n10674) );
  AND U11751 ( .A(n10675), .B(n10674), .Z(n10681) );
  XOR U11752 ( .A(n10682), .B(n10681), .Z(n10684) );
  XOR U11753 ( .A(n10683), .B(n10684), .Z(n10697) );
  XNOR U11754 ( .A(n10697), .B(sreg[1422]), .Z(n10699) );
  NANDN U11755 ( .A(n10676), .B(sreg[1421]), .Z(n10680) );
  NAND U11756 ( .A(n10678), .B(n10677), .Z(n10679) );
  NAND U11757 ( .A(n10680), .B(n10679), .Z(n10698) );
  XOR U11758 ( .A(n10699), .B(n10698), .Z(c[1422]) );
  NANDN U11759 ( .A(n10682), .B(n10681), .Z(n10686) );
  OR U11760 ( .A(n10684), .B(n10683), .Z(n10685) );
  AND U11761 ( .A(n10686), .B(n10685), .Z(n10704) );
  XOR U11762 ( .A(a[401]), .B(n2233), .Z(n10708) );
  AND U11763 ( .A(a[399]), .B(b[3]), .Z(n10712) );
  AND U11764 ( .A(a[403]), .B(b[0]), .Z(n10688) );
  XNOR U11765 ( .A(n10688), .B(n2175), .Z(n10690) );
  NANDN U11766 ( .A(b[0]), .B(a[402]), .Z(n10689) );
  NAND U11767 ( .A(n10690), .B(n10689), .Z(n10713) );
  XOR U11768 ( .A(n10712), .B(n10713), .Z(n10715) );
  XOR U11769 ( .A(n10714), .B(n10715), .Z(n10703) );
  NANDN U11770 ( .A(n10692), .B(n10691), .Z(n10696) );
  OR U11771 ( .A(n10694), .B(n10693), .Z(n10695) );
  AND U11772 ( .A(n10696), .B(n10695), .Z(n10702) );
  XOR U11773 ( .A(n10703), .B(n10702), .Z(n10705) );
  XOR U11774 ( .A(n10704), .B(n10705), .Z(n10718) );
  XNOR U11775 ( .A(n10718), .B(sreg[1423]), .Z(n10720) );
  NANDN U11776 ( .A(n10697), .B(sreg[1422]), .Z(n10701) );
  NAND U11777 ( .A(n10699), .B(n10698), .Z(n10700) );
  NAND U11778 ( .A(n10701), .B(n10700), .Z(n10719) );
  XOR U11779 ( .A(n10720), .B(n10719), .Z(c[1423]) );
  NANDN U11780 ( .A(n10703), .B(n10702), .Z(n10707) );
  OR U11781 ( .A(n10705), .B(n10704), .Z(n10706) );
  AND U11782 ( .A(n10707), .B(n10706), .Z(n10725) );
  XOR U11783 ( .A(a[402]), .B(n2233), .Z(n10729) );
  AND U11784 ( .A(a[404]), .B(b[0]), .Z(n10709) );
  XNOR U11785 ( .A(n10709), .B(n2175), .Z(n10711) );
  NANDN U11786 ( .A(b[0]), .B(a[403]), .Z(n10710) );
  NAND U11787 ( .A(n10711), .B(n10710), .Z(n10734) );
  AND U11788 ( .A(a[400]), .B(b[3]), .Z(n10733) );
  XOR U11789 ( .A(n10734), .B(n10733), .Z(n10736) );
  XOR U11790 ( .A(n10735), .B(n10736), .Z(n10724) );
  NANDN U11791 ( .A(n10713), .B(n10712), .Z(n10717) );
  OR U11792 ( .A(n10715), .B(n10714), .Z(n10716) );
  AND U11793 ( .A(n10717), .B(n10716), .Z(n10723) );
  XOR U11794 ( .A(n10724), .B(n10723), .Z(n10726) );
  XOR U11795 ( .A(n10725), .B(n10726), .Z(n10739) );
  XNOR U11796 ( .A(n10739), .B(sreg[1424]), .Z(n10741) );
  NANDN U11797 ( .A(n10718), .B(sreg[1423]), .Z(n10722) );
  NAND U11798 ( .A(n10720), .B(n10719), .Z(n10721) );
  NAND U11799 ( .A(n10722), .B(n10721), .Z(n10740) );
  XOR U11800 ( .A(n10741), .B(n10740), .Z(c[1424]) );
  NANDN U11801 ( .A(n10724), .B(n10723), .Z(n10728) );
  OR U11802 ( .A(n10726), .B(n10725), .Z(n10727) );
  AND U11803 ( .A(n10728), .B(n10727), .Z(n10746) );
  XOR U11804 ( .A(a[403]), .B(n2233), .Z(n10750) );
  AND U11805 ( .A(a[401]), .B(b[3]), .Z(n10754) );
  AND U11806 ( .A(a[405]), .B(b[0]), .Z(n10730) );
  XNOR U11807 ( .A(n10730), .B(n2175), .Z(n10732) );
  NANDN U11808 ( .A(b[0]), .B(a[404]), .Z(n10731) );
  NAND U11809 ( .A(n10732), .B(n10731), .Z(n10755) );
  XOR U11810 ( .A(n10754), .B(n10755), .Z(n10757) );
  XOR U11811 ( .A(n10756), .B(n10757), .Z(n10745) );
  NANDN U11812 ( .A(n10734), .B(n10733), .Z(n10738) );
  OR U11813 ( .A(n10736), .B(n10735), .Z(n10737) );
  AND U11814 ( .A(n10738), .B(n10737), .Z(n10744) );
  XOR U11815 ( .A(n10745), .B(n10744), .Z(n10747) );
  XOR U11816 ( .A(n10746), .B(n10747), .Z(n10760) );
  XNOR U11817 ( .A(n10760), .B(sreg[1425]), .Z(n10762) );
  NANDN U11818 ( .A(n10739), .B(sreg[1424]), .Z(n10743) );
  NAND U11819 ( .A(n10741), .B(n10740), .Z(n10742) );
  NAND U11820 ( .A(n10743), .B(n10742), .Z(n10761) );
  XOR U11821 ( .A(n10762), .B(n10761), .Z(c[1425]) );
  NANDN U11822 ( .A(n10745), .B(n10744), .Z(n10749) );
  OR U11823 ( .A(n10747), .B(n10746), .Z(n10748) );
  AND U11824 ( .A(n10749), .B(n10748), .Z(n10767) );
  XOR U11825 ( .A(a[404]), .B(n2233), .Z(n10771) );
  AND U11826 ( .A(a[406]), .B(b[0]), .Z(n10751) );
  XNOR U11827 ( .A(n10751), .B(n2175), .Z(n10753) );
  NANDN U11828 ( .A(b[0]), .B(a[405]), .Z(n10752) );
  NAND U11829 ( .A(n10753), .B(n10752), .Z(n10776) );
  AND U11830 ( .A(a[402]), .B(b[3]), .Z(n10775) );
  XOR U11831 ( .A(n10776), .B(n10775), .Z(n10778) );
  XOR U11832 ( .A(n10777), .B(n10778), .Z(n10766) );
  NANDN U11833 ( .A(n10755), .B(n10754), .Z(n10759) );
  OR U11834 ( .A(n10757), .B(n10756), .Z(n10758) );
  AND U11835 ( .A(n10759), .B(n10758), .Z(n10765) );
  XOR U11836 ( .A(n10766), .B(n10765), .Z(n10768) );
  XOR U11837 ( .A(n10767), .B(n10768), .Z(n10781) );
  XNOR U11838 ( .A(n10781), .B(sreg[1426]), .Z(n10783) );
  NANDN U11839 ( .A(n10760), .B(sreg[1425]), .Z(n10764) );
  NAND U11840 ( .A(n10762), .B(n10761), .Z(n10763) );
  NAND U11841 ( .A(n10764), .B(n10763), .Z(n10782) );
  XOR U11842 ( .A(n10783), .B(n10782), .Z(c[1426]) );
  NANDN U11843 ( .A(n10766), .B(n10765), .Z(n10770) );
  OR U11844 ( .A(n10768), .B(n10767), .Z(n10769) );
  AND U11845 ( .A(n10770), .B(n10769), .Z(n10788) );
  XOR U11846 ( .A(a[405]), .B(n2234), .Z(n10792) );
  AND U11847 ( .A(a[403]), .B(b[3]), .Z(n10796) );
  AND U11848 ( .A(a[407]), .B(b[0]), .Z(n10772) );
  XNOR U11849 ( .A(n10772), .B(n2175), .Z(n10774) );
  NANDN U11850 ( .A(b[0]), .B(a[406]), .Z(n10773) );
  NAND U11851 ( .A(n10774), .B(n10773), .Z(n10797) );
  XOR U11852 ( .A(n10796), .B(n10797), .Z(n10799) );
  XOR U11853 ( .A(n10798), .B(n10799), .Z(n10787) );
  NANDN U11854 ( .A(n10776), .B(n10775), .Z(n10780) );
  OR U11855 ( .A(n10778), .B(n10777), .Z(n10779) );
  AND U11856 ( .A(n10780), .B(n10779), .Z(n10786) );
  XOR U11857 ( .A(n10787), .B(n10786), .Z(n10789) );
  XOR U11858 ( .A(n10788), .B(n10789), .Z(n10802) );
  XNOR U11859 ( .A(n10802), .B(sreg[1427]), .Z(n10804) );
  NANDN U11860 ( .A(n10781), .B(sreg[1426]), .Z(n10785) );
  NAND U11861 ( .A(n10783), .B(n10782), .Z(n10784) );
  NAND U11862 ( .A(n10785), .B(n10784), .Z(n10803) );
  XOR U11863 ( .A(n10804), .B(n10803), .Z(c[1427]) );
  NANDN U11864 ( .A(n10787), .B(n10786), .Z(n10791) );
  OR U11865 ( .A(n10789), .B(n10788), .Z(n10790) );
  AND U11866 ( .A(n10791), .B(n10790), .Z(n10809) );
  XOR U11867 ( .A(a[406]), .B(n2234), .Z(n10813) );
  AND U11868 ( .A(a[408]), .B(b[0]), .Z(n10793) );
  XNOR U11869 ( .A(n10793), .B(n2175), .Z(n10795) );
  NANDN U11870 ( .A(b[0]), .B(a[407]), .Z(n10794) );
  NAND U11871 ( .A(n10795), .B(n10794), .Z(n10818) );
  AND U11872 ( .A(a[404]), .B(b[3]), .Z(n10817) );
  XOR U11873 ( .A(n10818), .B(n10817), .Z(n10820) );
  XOR U11874 ( .A(n10819), .B(n10820), .Z(n10808) );
  NANDN U11875 ( .A(n10797), .B(n10796), .Z(n10801) );
  OR U11876 ( .A(n10799), .B(n10798), .Z(n10800) );
  AND U11877 ( .A(n10801), .B(n10800), .Z(n10807) );
  XOR U11878 ( .A(n10808), .B(n10807), .Z(n10810) );
  XOR U11879 ( .A(n10809), .B(n10810), .Z(n10823) );
  XNOR U11880 ( .A(n10823), .B(sreg[1428]), .Z(n10825) );
  NANDN U11881 ( .A(n10802), .B(sreg[1427]), .Z(n10806) );
  NAND U11882 ( .A(n10804), .B(n10803), .Z(n10805) );
  NAND U11883 ( .A(n10806), .B(n10805), .Z(n10824) );
  XOR U11884 ( .A(n10825), .B(n10824), .Z(c[1428]) );
  NANDN U11885 ( .A(n10808), .B(n10807), .Z(n10812) );
  OR U11886 ( .A(n10810), .B(n10809), .Z(n10811) );
  AND U11887 ( .A(n10812), .B(n10811), .Z(n10830) );
  XOR U11888 ( .A(a[407]), .B(n2234), .Z(n10834) );
  AND U11889 ( .A(a[409]), .B(b[0]), .Z(n10814) );
  XNOR U11890 ( .A(n10814), .B(n2175), .Z(n10816) );
  NANDN U11891 ( .A(b[0]), .B(a[408]), .Z(n10815) );
  NAND U11892 ( .A(n10816), .B(n10815), .Z(n10839) );
  AND U11893 ( .A(a[405]), .B(b[3]), .Z(n10838) );
  XOR U11894 ( .A(n10839), .B(n10838), .Z(n10841) );
  XOR U11895 ( .A(n10840), .B(n10841), .Z(n10829) );
  NANDN U11896 ( .A(n10818), .B(n10817), .Z(n10822) );
  OR U11897 ( .A(n10820), .B(n10819), .Z(n10821) );
  AND U11898 ( .A(n10822), .B(n10821), .Z(n10828) );
  XOR U11899 ( .A(n10829), .B(n10828), .Z(n10831) );
  XOR U11900 ( .A(n10830), .B(n10831), .Z(n10844) );
  XNOR U11901 ( .A(n10844), .B(sreg[1429]), .Z(n10846) );
  NANDN U11902 ( .A(n10823), .B(sreg[1428]), .Z(n10827) );
  NAND U11903 ( .A(n10825), .B(n10824), .Z(n10826) );
  NAND U11904 ( .A(n10827), .B(n10826), .Z(n10845) );
  XOR U11905 ( .A(n10846), .B(n10845), .Z(c[1429]) );
  NANDN U11906 ( .A(n10829), .B(n10828), .Z(n10833) );
  OR U11907 ( .A(n10831), .B(n10830), .Z(n10832) );
  AND U11908 ( .A(n10833), .B(n10832), .Z(n10851) );
  XOR U11909 ( .A(a[408]), .B(n2234), .Z(n10855) );
  AND U11910 ( .A(a[410]), .B(b[0]), .Z(n10835) );
  XNOR U11911 ( .A(n10835), .B(n2175), .Z(n10837) );
  NANDN U11912 ( .A(b[0]), .B(a[409]), .Z(n10836) );
  NAND U11913 ( .A(n10837), .B(n10836), .Z(n10860) );
  AND U11914 ( .A(a[406]), .B(b[3]), .Z(n10859) );
  XOR U11915 ( .A(n10860), .B(n10859), .Z(n10862) );
  XOR U11916 ( .A(n10861), .B(n10862), .Z(n10850) );
  NANDN U11917 ( .A(n10839), .B(n10838), .Z(n10843) );
  OR U11918 ( .A(n10841), .B(n10840), .Z(n10842) );
  AND U11919 ( .A(n10843), .B(n10842), .Z(n10849) );
  XOR U11920 ( .A(n10850), .B(n10849), .Z(n10852) );
  XOR U11921 ( .A(n10851), .B(n10852), .Z(n10865) );
  XNOR U11922 ( .A(n10865), .B(sreg[1430]), .Z(n10867) );
  NANDN U11923 ( .A(n10844), .B(sreg[1429]), .Z(n10848) );
  NAND U11924 ( .A(n10846), .B(n10845), .Z(n10847) );
  NAND U11925 ( .A(n10848), .B(n10847), .Z(n10866) );
  XOR U11926 ( .A(n10867), .B(n10866), .Z(c[1430]) );
  NANDN U11927 ( .A(n10850), .B(n10849), .Z(n10854) );
  OR U11928 ( .A(n10852), .B(n10851), .Z(n10853) );
  AND U11929 ( .A(n10854), .B(n10853), .Z(n10872) );
  XOR U11930 ( .A(a[409]), .B(n2234), .Z(n10876) );
  AND U11931 ( .A(a[411]), .B(b[0]), .Z(n10856) );
  XNOR U11932 ( .A(n10856), .B(n2175), .Z(n10858) );
  NANDN U11933 ( .A(b[0]), .B(a[410]), .Z(n10857) );
  NAND U11934 ( .A(n10858), .B(n10857), .Z(n10881) );
  AND U11935 ( .A(a[407]), .B(b[3]), .Z(n10880) );
  XOR U11936 ( .A(n10881), .B(n10880), .Z(n10883) );
  XOR U11937 ( .A(n10882), .B(n10883), .Z(n10871) );
  NANDN U11938 ( .A(n10860), .B(n10859), .Z(n10864) );
  OR U11939 ( .A(n10862), .B(n10861), .Z(n10863) );
  AND U11940 ( .A(n10864), .B(n10863), .Z(n10870) );
  XOR U11941 ( .A(n10871), .B(n10870), .Z(n10873) );
  XOR U11942 ( .A(n10872), .B(n10873), .Z(n10886) );
  XNOR U11943 ( .A(n10886), .B(sreg[1431]), .Z(n10888) );
  NANDN U11944 ( .A(n10865), .B(sreg[1430]), .Z(n10869) );
  NAND U11945 ( .A(n10867), .B(n10866), .Z(n10868) );
  NAND U11946 ( .A(n10869), .B(n10868), .Z(n10887) );
  XOR U11947 ( .A(n10888), .B(n10887), .Z(c[1431]) );
  NANDN U11948 ( .A(n10871), .B(n10870), .Z(n10875) );
  OR U11949 ( .A(n10873), .B(n10872), .Z(n10874) );
  AND U11950 ( .A(n10875), .B(n10874), .Z(n10893) );
  XOR U11951 ( .A(a[410]), .B(n2234), .Z(n10897) );
  AND U11952 ( .A(a[412]), .B(b[0]), .Z(n10877) );
  XNOR U11953 ( .A(n10877), .B(n2175), .Z(n10879) );
  NANDN U11954 ( .A(b[0]), .B(a[411]), .Z(n10878) );
  NAND U11955 ( .A(n10879), .B(n10878), .Z(n10902) );
  AND U11956 ( .A(a[408]), .B(b[3]), .Z(n10901) );
  XOR U11957 ( .A(n10902), .B(n10901), .Z(n10904) );
  XOR U11958 ( .A(n10903), .B(n10904), .Z(n10892) );
  NANDN U11959 ( .A(n10881), .B(n10880), .Z(n10885) );
  OR U11960 ( .A(n10883), .B(n10882), .Z(n10884) );
  AND U11961 ( .A(n10885), .B(n10884), .Z(n10891) );
  XOR U11962 ( .A(n10892), .B(n10891), .Z(n10894) );
  XOR U11963 ( .A(n10893), .B(n10894), .Z(n10907) );
  XNOR U11964 ( .A(n10907), .B(sreg[1432]), .Z(n10909) );
  NANDN U11965 ( .A(n10886), .B(sreg[1431]), .Z(n10890) );
  NAND U11966 ( .A(n10888), .B(n10887), .Z(n10889) );
  NAND U11967 ( .A(n10890), .B(n10889), .Z(n10908) );
  XOR U11968 ( .A(n10909), .B(n10908), .Z(c[1432]) );
  NANDN U11969 ( .A(n10892), .B(n10891), .Z(n10896) );
  OR U11970 ( .A(n10894), .B(n10893), .Z(n10895) );
  AND U11971 ( .A(n10896), .B(n10895), .Z(n10914) );
  XOR U11972 ( .A(a[411]), .B(n2234), .Z(n10918) );
  AND U11973 ( .A(a[413]), .B(b[0]), .Z(n10898) );
  XNOR U11974 ( .A(n10898), .B(n2175), .Z(n10900) );
  NANDN U11975 ( .A(b[0]), .B(a[412]), .Z(n10899) );
  NAND U11976 ( .A(n10900), .B(n10899), .Z(n10923) );
  AND U11977 ( .A(a[409]), .B(b[3]), .Z(n10922) );
  XOR U11978 ( .A(n10923), .B(n10922), .Z(n10925) );
  XOR U11979 ( .A(n10924), .B(n10925), .Z(n10913) );
  NANDN U11980 ( .A(n10902), .B(n10901), .Z(n10906) );
  OR U11981 ( .A(n10904), .B(n10903), .Z(n10905) );
  AND U11982 ( .A(n10906), .B(n10905), .Z(n10912) );
  XOR U11983 ( .A(n10913), .B(n10912), .Z(n10915) );
  XOR U11984 ( .A(n10914), .B(n10915), .Z(n10928) );
  XNOR U11985 ( .A(n10928), .B(sreg[1433]), .Z(n10930) );
  NANDN U11986 ( .A(n10907), .B(sreg[1432]), .Z(n10911) );
  NAND U11987 ( .A(n10909), .B(n10908), .Z(n10910) );
  NAND U11988 ( .A(n10911), .B(n10910), .Z(n10929) );
  XOR U11989 ( .A(n10930), .B(n10929), .Z(c[1433]) );
  NANDN U11990 ( .A(n10913), .B(n10912), .Z(n10917) );
  OR U11991 ( .A(n10915), .B(n10914), .Z(n10916) );
  AND U11992 ( .A(n10917), .B(n10916), .Z(n10935) );
  XOR U11993 ( .A(a[412]), .B(n2235), .Z(n10939) );
  AND U11994 ( .A(a[414]), .B(b[0]), .Z(n10919) );
  XNOR U11995 ( .A(n10919), .B(n2175), .Z(n10921) );
  NANDN U11996 ( .A(b[0]), .B(a[413]), .Z(n10920) );
  NAND U11997 ( .A(n10921), .B(n10920), .Z(n10944) );
  AND U11998 ( .A(a[410]), .B(b[3]), .Z(n10943) );
  XOR U11999 ( .A(n10944), .B(n10943), .Z(n10946) );
  XOR U12000 ( .A(n10945), .B(n10946), .Z(n10934) );
  NANDN U12001 ( .A(n10923), .B(n10922), .Z(n10927) );
  OR U12002 ( .A(n10925), .B(n10924), .Z(n10926) );
  AND U12003 ( .A(n10927), .B(n10926), .Z(n10933) );
  XOR U12004 ( .A(n10934), .B(n10933), .Z(n10936) );
  XOR U12005 ( .A(n10935), .B(n10936), .Z(n10949) );
  XNOR U12006 ( .A(n10949), .B(sreg[1434]), .Z(n10951) );
  NANDN U12007 ( .A(n10928), .B(sreg[1433]), .Z(n10932) );
  NAND U12008 ( .A(n10930), .B(n10929), .Z(n10931) );
  NAND U12009 ( .A(n10932), .B(n10931), .Z(n10950) );
  XOR U12010 ( .A(n10951), .B(n10950), .Z(c[1434]) );
  NANDN U12011 ( .A(n10934), .B(n10933), .Z(n10938) );
  OR U12012 ( .A(n10936), .B(n10935), .Z(n10937) );
  AND U12013 ( .A(n10938), .B(n10937), .Z(n10956) );
  XOR U12014 ( .A(a[413]), .B(n2235), .Z(n10960) );
  AND U12015 ( .A(a[411]), .B(b[3]), .Z(n10964) );
  AND U12016 ( .A(a[415]), .B(b[0]), .Z(n10940) );
  XNOR U12017 ( .A(n10940), .B(n2175), .Z(n10942) );
  NANDN U12018 ( .A(b[0]), .B(a[414]), .Z(n10941) );
  NAND U12019 ( .A(n10942), .B(n10941), .Z(n10965) );
  XOR U12020 ( .A(n10964), .B(n10965), .Z(n10967) );
  XOR U12021 ( .A(n10966), .B(n10967), .Z(n10955) );
  NANDN U12022 ( .A(n10944), .B(n10943), .Z(n10948) );
  OR U12023 ( .A(n10946), .B(n10945), .Z(n10947) );
  AND U12024 ( .A(n10948), .B(n10947), .Z(n10954) );
  XOR U12025 ( .A(n10955), .B(n10954), .Z(n10957) );
  XOR U12026 ( .A(n10956), .B(n10957), .Z(n10970) );
  XNOR U12027 ( .A(n10970), .B(sreg[1435]), .Z(n10972) );
  NANDN U12028 ( .A(n10949), .B(sreg[1434]), .Z(n10953) );
  NAND U12029 ( .A(n10951), .B(n10950), .Z(n10952) );
  NAND U12030 ( .A(n10953), .B(n10952), .Z(n10971) );
  XOR U12031 ( .A(n10972), .B(n10971), .Z(c[1435]) );
  NANDN U12032 ( .A(n10955), .B(n10954), .Z(n10959) );
  OR U12033 ( .A(n10957), .B(n10956), .Z(n10958) );
  AND U12034 ( .A(n10959), .B(n10958), .Z(n10977) );
  XOR U12035 ( .A(a[414]), .B(n2235), .Z(n10981) );
  AND U12036 ( .A(a[416]), .B(b[0]), .Z(n10961) );
  XNOR U12037 ( .A(n10961), .B(n2175), .Z(n10963) );
  NANDN U12038 ( .A(b[0]), .B(a[415]), .Z(n10962) );
  NAND U12039 ( .A(n10963), .B(n10962), .Z(n10986) );
  AND U12040 ( .A(a[412]), .B(b[3]), .Z(n10985) );
  XOR U12041 ( .A(n10986), .B(n10985), .Z(n10988) );
  XOR U12042 ( .A(n10987), .B(n10988), .Z(n10976) );
  NANDN U12043 ( .A(n10965), .B(n10964), .Z(n10969) );
  OR U12044 ( .A(n10967), .B(n10966), .Z(n10968) );
  AND U12045 ( .A(n10969), .B(n10968), .Z(n10975) );
  XOR U12046 ( .A(n10976), .B(n10975), .Z(n10978) );
  XOR U12047 ( .A(n10977), .B(n10978), .Z(n10991) );
  XNOR U12048 ( .A(n10991), .B(sreg[1436]), .Z(n10993) );
  NANDN U12049 ( .A(n10970), .B(sreg[1435]), .Z(n10974) );
  NAND U12050 ( .A(n10972), .B(n10971), .Z(n10973) );
  NAND U12051 ( .A(n10974), .B(n10973), .Z(n10992) );
  XOR U12052 ( .A(n10993), .B(n10992), .Z(c[1436]) );
  NANDN U12053 ( .A(n10976), .B(n10975), .Z(n10980) );
  OR U12054 ( .A(n10978), .B(n10977), .Z(n10979) );
  AND U12055 ( .A(n10980), .B(n10979), .Z(n10998) );
  XOR U12056 ( .A(a[415]), .B(n2235), .Z(n11002) );
  AND U12057 ( .A(a[413]), .B(b[3]), .Z(n11006) );
  AND U12058 ( .A(a[417]), .B(b[0]), .Z(n10982) );
  XNOR U12059 ( .A(n10982), .B(n2175), .Z(n10984) );
  NANDN U12060 ( .A(b[0]), .B(a[416]), .Z(n10983) );
  NAND U12061 ( .A(n10984), .B(n10983), .Z(n11007) );
  XOR U12062 ( .A(n11006), .B(n11007), .Z(n11009) );
  XOR U12063 ( .A(n11008), .B(n11009), .Z(n10997) );
  NANDN U12064 ( .A(n10986), .B(n10985), .Z(n10990) );
  OR U12065 ( .A(n10988), .B(n10987), .Z(n10989) );
  AND U12066 ( .A(n10990), .B(n10989), .Z(n10996) );
  XOR U12067 ( .A(n10997), .B(n10996), .Z(n10999) );
  XOR U12068 ( .A(n10998), .B(n10999), .Z(n11012) );
  XNOR U12069 ( .A(n11012), .B(sreg[1437]), .Z(n11014) );
  NANDN U12070 ( .A(n10991), .B(sreg[1436]), .Z(n10995) );
  NAND U12071 ( .A(n10993), .B(n10992), .Z(n10994) );
  NAND U12072 ( .A(n10995), .B(n10994), .Z(n11013) );
  XOR U12073 ( .A(n11014), .B(n11013), .Z(c[1437]) );
  NANDN U12074 ( .A(n10997), .B(n10996), .Z(n11001) );
  OR U12075 ( .A(n10999), .B(n10998), .Z(n11000) );
  AND U12076 ( .A(n11001), .B(n11000), .Z(n11019) );
  XOR U12077 ( .A(a[416]), .B(n2235), .Z(n11023) );
  AND U12078 ( .A(a[414]), .B(b[3]), .Z(n11027) );
  AND U12079 ( .A(a[418]), .B(b[0]), .Z(n11003) );
  XNOR U12080 ( .A(n11003), .B(n2175), .Z(n11005) );
  NANDN U12081 ( .A(b[0]), .B(a[417]), .Z(n11004) );
  NAND U12082 ( .A(n11005), .B(n11004), .Z(n11028) );
  XOR U12083 ( .A(n11027), .B(n11028), .Z(n11030) );
  XOR U12084 ( .A(n11029), .B(n11030), .Z(n11018) );
  NANDN U12085 ( .A(n11007), .B(n11006), .Z(n11011) );
  OR U12086 ( .A(n11009), .B(n11008), .Z(n11010) );
  AND U12087 ( .A(n11011), .B(n11010), .Z(n11017) );
  XOR U12088 ( .A(n11018), .B(n11017), .Z(n11020) );
  XOR U12089 ( .A(n11019), .B(n11020), .Z(n11033) );
  XNOR U12090 ( .A(n11033), .B(sreg[1438]), .Z(n11035) );
  NANDN U12091 ( .A(n11012), .B(sreg[1437]), .Z(n11016) );
  NAND U12092 ( .A(n11014), .B(n11013), .Z(n11015) );
  NAND U12093 ( .A(n11016), .B(n11015), .Z(n11034) );
  XOR U12094 ( .A(n11035), .B(n11034), .Z(c[1438]) );
  NANDN U12095 ( .A(n11018), .B(n11017), .Z(n11022) );
  OR U12096 ( .A(n11020), .B(n11019), .Z(n11021) );
  AND U12097 ( .A(n11022), .B(n11021), .Z(n11040) );
  XOR U12098 ( .A(a[417]), .B(n2235), .Z(n11044) );
  AND U12099 ( .A(a[419]), .B(b[0]), .Z(n11024) );
  XNOR U12100 ( .A(n11024), .B(n2175), .Z(n11026) );
  NANDN U12101 ( .A(b[0]), .B(a[418]), .Z(n11025) );
  NAND U12102 ( .A(n11026), .B(n11025), .Z(n11049) );
  AND U12103 ( .A(a[415]), .B(b[3]), .Z(n11048) );
  XOR U12104 ( .A(n11049), .B(n11048), .Z(n11051) );
  XOR U12105 ( .A(n11050), .B(n11051), .Z(n11039) );
  NANDN U12106 ( .A(n11028), .B(n11027), .Z(n11032) );
  OR U12107 ( .A(n11030), .B(n11029), .Z(n11031) );
  AND U12108 ( .A(n11032), .B(n11031), .Z(n11038) );
  XOR U12109 ( .A(n11039), .B(n11038), .Z(n11041) );
  XOR U12110 ( .A(n11040), .B(n11041), .Z(n11054) );
  XNOR U12111 ( .A(n11054), .B(sreg[1439]), .Z(n11056) );
  NANDN U12112 ( .A(n11033), .B(sreg[1438]), .Z(n11037) );
  NAND U12113 ( .A(n11035), .B(n11034), .Z(n11036) );
  NAND U12114 ( .A(n11037), .B(n11036), .Z(n11055) );
  XOR U12115 ( .A(n11056), .B(n11055), .Z(c[1439]) );
  NANDN U12116 ( .A(n11039), .B(n11038), .Z(n11043) );
  OR U12117 ( .A(n11041), .B(n11040), .Z(n11042) );
  AND U12118 ( .A(n11043), .B(n11042), .Z(n11061) );
  XOR U12119 ( .A(a[418]), .B(n2235), .Z(n11065) );
  AND U12120 ( .A(a[420]), .B(b[0]), .Z(n11045) );
  XNOR U12121 ( .A(n11045), .B(n2175), .Z(n11047) );
  NANDN U12122 ( .A(b[0]), .B(a[419]), .Z(n11046) );
  NAND U12123 ( .A(n11047), .B(n11046), .Z(n11070) );
  AND U12124 ( .A(a[416]), .B(b[3]), .Z(n11069) );
  XOR U12125 ( .A(n11070), .B(n11069), .Z(n11072) );
  XOR U12126 ( .A(n11071), .B(n11072), .Z(n11060) );
  NANDN U12127 ( .A(n11049), .B(n11048), .Z(n11053) );
  OR U12128 ( .A(n11051), .B(n11050), .Z(n11052) );
  AND U12129 ( .A(n11053), .B(n11052), .Z(n11059) );
  XOR U12130 ( .A(n11060), .B(n11059), .Z(n11062) );
  XOR U12131 ( .A(n11061), .B(n11062), .Z(n11075) );
  XNOR U12132 ( .A(n11075), .B(sreg[1440]), .Z(n11077) );
  NANDN U12133 ( .A(n11054), .B(sreg[1439]), .Z(n11058) );
  NAND U12134 ( .A(n11056), .B(n11055), .Z(n11057) );
  NAND U12135 ( .A(n11058), .B(n11057), .Z(n11076) );
  XOR U12136 ( .A(n11077), .B(n11076), .Z(c[1440]) );
  NANDN U12137 ( .A(n11060), .B(n11059), .Z(n11064) );
  OR U12138 ( .A(n11062), .B(n11061), .Z(n11063) );
  AND U12139 ( .A(n11064), .B(n11063), .Z(n11082) );
  XOR U12140 ( .A(a[419]), .B(n2236), .Z(n11086) );
  AND U12141 ( .A(a[421]), .B(b[0]), .Z(n11066) );
  XNOR U12142 ( .A(n11066), .B(n2175), .Z(n11068) );
  NANDN U12143 ( .A(b[0]), .B(a[420]), .Z(n11067) );
  NAND U12144 ( .A(n11068), .B(n11067), .Z(n11091) );
  AND U12145 ( .A(a[417]), .B(b[3]), .Z(n11090) );
  XOR U12146 ( .A(n11091), .B(n11090), .Z(n11093) );
  XOR U12147 ( .A(n11092), .B(n11093), .Z(n11081) );
  NANDN U12148 ( .A(n11070), .B(n11069), .Z(n11074) );
  OR U12149 ( .A(n11072), .B(n11071), .Z(n11073) );
  AND U12150 ( .A(n11074), .B(n11073), .Z(n11080) );
  XOR U12151 ( .A(n11081), .B(n11080), .Z(n11083) );
  XOR U12152 ( .A(n11082), .B(n11083), .Z(n11096) );
  XNOR U12153 ( .A(n11096), .B(sreg[1441]), .Z(n11098) );
  NANDN U12154 ( .A(n11075), .B(sreg[1440]), .Z(n11079) );
  NAND U12155 ( .A(n11077), .B(n11076), .Z(n11078) );
  NAND U12156 ( .A(n11079), .B(n11078), .Z(n11097) );
  XOR U12157 ( .A(n11098), .B(n11097), .Z(c[1441]) );
  NANDN U12158 ( .A(n11081), .B(n11080), .Z(n11085) );
  OR U12159 ( .A(n11083), .B(n11082), .Z(n11084) );
  AND U12160 ( .A(n11085), .B(n11084), .Z(n11103) );
  XOR U12161 ( .A(a[420]), .B(n2236), .Z(n11107) );
  AND U12162 ( .A(a[418]), .B(b[3]), .Z(n11111) );
  AND U12163 ( .A(a[422]), .B(b[0]), .Z(n11087) );
  XNOR U12164 ( .A(n11087), .B(n2175), .Z(n11089) );
  NANDN U12165 ( .A(b[0]), .B(a[421]), .Z(n11088) );
  NAND U12166 ( .A(n11089), .B(n11088), .Z(n11112) );
  XOR U12167 ( .A(n11111), .B(n11112), .Z(n11114) );
  XOR U12168 ( .A(n11113), .B(n11114), .Z(n11102) );
  NANDN U12169 ( .A(n11091), .B(n11090), .Z(n11095) );
  OR U12170 ( .A(n11093), .B(n11092), .Z(n11094) );
  AND U12171 ( .A(n11095), .B(n11094), .Z(n11101) );
  XOR U12172 ( .A(n11102), .B(n11101), .Z(n11104) );
  XOR U12173 ( .A(n11103), .B(n11104), .Z(n11117) );
  XNOR U12174 ( .A(n11117), .B(sreg[1442]), .Z(n11119) );
  NANDN U12175 ( .A(n11096), .B(sreg[1441]), .Z(n11100) );
  NAND U12176 ( .A(n11098), .B(n11097), .Z(n11099) );
  NAND U12177 ( .A(n11100), .B(n11099), .Z(n11118) );
  XOR U12178 ( .A(n11119), .B(n11118), .Z(c[1442]) );
  NANDN U12179 ( .A(n11102), .B(n11101), .Z(n11106) );
  OR U12180 ( .A(n11104), .B(n11103), .Z(n11105) );
  AND U12181 ( .A(n11106), .B(n11105), .Z(n11124) );
  XOR U12182 ( .A(a[421]), .B(n2236), .Z(n11128) );
  AND U12183 ( .A(a[419]), .B(b[3]), .Z(n11132) );
  AND U12184 ( .A(a[423]), .B(b[0]), .Z(n11108) );
  XNOR U12185 ( .A(n11108), .B(n2175), .Z(n11110) );
  NANDN U12186 ( .A(b[0]), .B(a[422]), .Z(n11109) );
  NAND U12187 ( .A(n11110), .B(n11109), .Z(n11133) );
  XOR U12188 ( .A(n11132), .B(n11133), .Z(n11135) );
  XOR U12189 ( .A(n11134), .B(n11135), .Z(n11123) );
  NANDN U12190 ( .A(n11112), .B(n11111), .Z(n11116) );
  OR U12191 ( .A(n11114), .B(n11113), .Z(n11115) );
  AND U12192 ( .A(n11116), .B(n11115), .Z(n11122) );
  XOR U12193 ( .A(n11123), .B(n11122), .Z(n11125) );
  XOR U12194 ( .A(n11124), .B(n11125), .Z(n11138) );
  XNOR U12195 ( .A(n11138), .B(sreg[1443]), .Z(n11140) );
  NANDN U12196 ( .A(n11117), .B(sreg[1442]), .Z(n11121) );
  NAND U12197 ( .A(n11119), .B(n11118), .Z(n11120) );
  NAND U12198 ( .A(n11121), .B(n11120), .Z(n11139) );
  XOR U12199 ( .A(n11140), .B(n11139), .Z(c[1443]) );
  NANDN U12200 ( .A(n11123), .B(n11122), .Z(n11127) );
  OR U12201 ( .A(n11125), .B(n11124), .Z(n11126) );
  AND U12202 ( .A(n11127), .B(n11126), .Z(n11145) );
  XOR U12203 ( .A(a[422]), .B(n2236), .Z(n11149) );
  AND U12204 ( .A(a[424]), .B(b[0]), .Z(n11129) );
  XNOR U12205 ( .A(n11129), .B(n2175), .Z(n11131) );
  NANDN U12206 ( .A(b[0]), .B(a[423]), .Z(n11130) );
  NAND U12207 ( .A(n11131), .B(n11130), .Z(n11154) );
  AND U12208 ( .A(a[420]), .B(b[3]), .Z(n11153) );
  XOR U12209 ( .A(n11154), .B(n11153), .Z(n11156) );
  XOR U12210 ( .A(n11155), .B(n11156), .Z(n11144) );
  NANDN U12211 ( .A(n11133), .B(n11132), .Z(n11137) );
  OR U12212 ( .A(n11135), .B(n11134), .Z(n11136) );
  AND U12213 ( .A(n11137), .B(n11136), .Z(n11143) );
  XOR U12214 ( .A(n11144), .B(n11143), .Z(n11146) );
  XOR U12215 ( .A(n11145), .B(n11146), .Z(n11159) );
  XNOR U12216 ( .A(n11159), .B(sreg[1444]), .Z(n11161) );
  NANDN U12217 ( .A(n11138), .B(sreg[1443]), .Z(n11142) );
  NAND U12218 ( .A(n11140), .B(n11139), .Z(n11141) );
  NAND U12219 ( .A(n11142), .B(n11141), .Z(n11160) );
  XOR U12220 ( .A(n11161), .B(n11160), .Z(c[1444]) );
  NANDN U12221 ( .A(n11144), .B(n11143), .Z(n11148) );
  OR U12222 ( .A(n11146), .B(n11145), .Z(n11147) );
  AND U12223 ( .A(n11148), .B(n11147), .Z(n11166) );
  XOR U12224 ( .A(a[423]), .B(n2236), .Z(n11170) );
  AND U12225 ( .A(a[425]), .B(b[0]), .Z(n11150) );
  XNOR U12226 ( .A(n11150), .B(n2175), .Z(n11152) );
  NANDN U12227 ( .A(b[0]), .B(a[424]), .Z(n11151) );
  NAND U12228 ( .A(n11152), .B(n11151), .Z(n11175) );
  AND U12229 ( .A(a[421]), .B(b[3]), .Z(n11174) );
  XOR U12230 ( .A(n11175), .B(n11174), .Z(n11177) );
  XOR U12231 ( .A(n11176), .B(n11177), .Z(n11165) );
  NANDN U12232 ( .A(n11154), .B(n11153), .Z(n11158) );
  OR U12233 ( .A(n11156), .B(n11155), .Z(n11157) );
  AND U12234 ( .A(n11158), .B(n11157), .Z(n11164) );
  XOR U12235 ( .A(n11165), .B(n11164), .Z(n11167) );
  XOR U12236 ( .A(n11166), .B(n11167), .Z(n11180) );
  XNOR U12237 ( .A(n11180), .B(sreg[1445]), .Z(n11182) );
  NANDN U12238 ( .A(n11159), .B(sreg[1444]), .Z(n11163) );
  NAND U12239 ( .A(n11161), .B(n11160), .Z(n11162) );
  NAND U12240 ( .A(n11163), .B(n11162), .Z(n11181) );
  XOR U12241 ( .A(n11182), .B(n11181), .Z(c[1445]) );
  NANDN U12242 ( .A(n11165), .B(n11164), .Z(n11169) );
  OR U12243 ( .A(n11167), .B(n11166), .Z(n11168) );
  AND U12244 ( .A(n11169), .B(n11168), .Z(n11187) );
  XOR U12245 ( .A(a[424]), .B(n2236), .Z(n11191) );
  AND U12246 ( .A(a[422]), .B(b[3]), .Z(n11195) );
  AND U12247 ( .A(a[426]), .B(b[0]), .Z(n11171) );
  XNOR U12248 ( .A(n11171), .B(n2175), .Z(n11173) );
  NANDN U12249 ( .A(b[0]), .B(a[425]), .Z(n11172) );
  NAND U12250 ( .A(n11173), .B(n11172), .Z(n11196) );
  XOR U12251 ( .A(n11195), .B(n11196), .Z(n11198) );
  XOR U12252 ( .A(n11197), .B(n11198), .Z(n11186) );
  NANDN U12253 ( .A(n11175), .B(n11174), .Z(n11179) );
  OR U12254 ( .A(n11177), .B(n11176), .Z(n11178) );
  AND U12255 ( .A(n11179), .B(n11178), .Z(n11185) );
  XOR U12256 ( .A(n11186), .B(n11185), .Z(n11188) );
  XOR U12257 ( .A(n11187), .B(n11188), .Z(n11201) );
  XNOR U12258 ( .A(n11201), .B(sreg[1446]), .Z(n11203) );
  NANDN U12259 ( .A(n11180), .B(sreg[1445]), .Z(n11184) );
  NAND U12260 ( .A(n11182), .B(n11181), .Z(n11183) );
  NAND U12261 ( .A(n11184), .B(n11183), .Z(n11202) );
  XOR U12262 ( .A(n11203), .B(n11202), .Z(c[1446]) );
  NANDN U12263 ( .A(n11186), .B(n11185), .Z(n11190) );
  OR U12264 ( .A(n11188), .B(n11187), .Z(n11189) );
  AND U12265 ( .A(n11190), .B(n11189), .Z(n11208) );
  XOR U12266 ( .A(a[425]), .B(n2236), .Z(n11212) );
  AND U12267 ( .A(a[423]), .B(b[3]), .Z(n11216) );
  AND U12268 ( .A(a[427]), .B(b[0]), .Z(n11192) );
  XNOR U12269 ( .A(n11192), .B(n2175), .Z(n11194) );
  NANDN U12270 ( .A(b[0]), .B(a[426]), .Z(n11193) );
  NAND U12271 ( .A(n11194), .B(n11193), .Z(n11217) );
  XOR U12272 ( .A(n11216), .B(n11217), .Z(n11219) );
  XOR U12273 ( .A(n11218), .B(n11219), .Z(n11207) );
  NANDN U12274 ( .A(n11196), .B(n11195), .Z(n11200) );
  OR U12275 ( .A(n11198), .B(n11197), .Z(n11199) );
  AND U12276 ( .A(n11200), .B(n11199), .Z(n11206) );
  XOR U12277 ( .A(n11207), .B(n11206), .Z(n11209) );
  XOR U12278 ( .A(n11208), .B(n11209), .Z(n11222) );
  XNOR U12279 ( .A(n11222), .B(sreg[1447]), .Z(n11224) );
  NANDN U12280 ( .A(n11201), .B(sreg[1446]), .Z(n11205) );
  NAND U12281 ( .A(n11203), .B(n11202), .Z(n11204) );
  NAND U12282 ( .A(n11205), .B(n11204), .Z(n11223) );
  XOR U12283 ( .A(n11224), .B(n11223), .Z(c[1447]) );
  NANDN U12284 ( .A(n11207), .B(n11206), .Z(n11211) );
  OR U12285 ( .A(n11209), .B(n11208), .Z(n11210) );
  AND U12286 ( .A(n11211), .B(n11210), .Z(n11229) );
  XOR U12287 ( .A(a[426]), .B(n2237), .Z(n11233) );
  AND U12288 ( .A(a[428]), .B(b[0]), .Z(n11213) );
  XNOR U12289 ( .A(n11213), .B(n2175), .Z(n11215) );
  NANDN U12290 ( .A(b[0]), .B(a[427]), .Z(n11214) );
  NAND U12291 ( .A(n11215), .B(n11214), .Z(n11238) );
  AND U12292 ( .A(a[424]), .B(b[3]), .Z(n11237) );
  XOR U12293 ( .A(n11238), .B(n11237), .Z(n11240) );
  XOR U12294 ( .A(n11239), .B(n11240), .Z(n11228) );
  NANDN U12295 ( .A(n11217), .B(n11216), .Z(n11221) );
  OR U12296 ( .A(n11219), .B(n11218), .Z(n11220) );
  AND U12297 ( .A(n11221), .B(n11220), .Z(n11227) );
  XOR U12298 ( .A(n11228), .B(n11227), .Z(n11230) );
  XOR U12299 ( .A(n11229), .B(n11230), .Z(n11243) );
  XNOR U12300 ( .A(n11243), .B(sreg[1448]), .Z(n11245) );
  NANDN U12301 ( .A(n11222), .B(sreg[1447]), .Z(n11226) );
  NAND U12302 ( .A(n11224), .B(n11223), .Z(n11225) );
  NAND U12303 ( .A(n11226), .B(n11225), .Z(n11244) );
  XOR U12304 ( .A(n11245), .B(n11244), .Z(c[1448]) );
  NANDN U12305 ( .A(n11228), .B(n11227), .Z(n11232) );
  OR U12306 ( .A(n11230), .B(n11229), .Z(n11231) );
  AND U12307 ( .A(n11232), .B(n11231), .Z(n11250) );
  XOR U12308 ( .A(a[427]), .B(n2237), .Z(n11254) );
  AND U12309 ( .A(a[429]), .B(b[0]), .Z(n11234) );
  XNOR U12310 ( .A(n11234), .B(n2175), .Z(n11236) );
  NANDN U12311 ( .A(b[0]), .B(a[428]), .Z(n11235) );
  NAND U12312 ( .A(n11236), .B(n11235), .Z(n11259) );
  AND U12313 ( .A(a[425]), .B(b[3]), .Z(n11258) );
  XOR U12314 ( .A(n11259), .B(n11258), .Z(n11261) );
  XOR U12315 ( .A(n11260), .B(n11261), .Z(n11249) );
  NANDN U12316 ( .A(n11238), .B(n11237), .Z(n11242) );
  OR U12317 ( .A(n11240), .B(n11239), .Z(n11241) );
  AND U12318 ( .A(n11242), .B(n11241), .Z(n11248) );
  XOR U12319 ( .A(n11249), .B(n11248), .Z(n11251) );
  XOR U12320 ( .A(n11250), .B(n11251), .Z(n11264) );
  XNOR U12321 ( .A(n11264), .B(sreg[1449]), .Z(n11266) );
  NANDN U12322 ( .A(n11243), .B(sreg[1448]), .Z(n11247) );
  NAND U12323 ( .A(n11245), .B(n11244), .Z(n11246) );
  NAND U12324 ( .A(n11247), .B(n11246), .Z(n11265) );
  XOR U12325 ( .A(n11266), .B(n11265), .Z(c[1449]) );
  NANDN U12326 ( .A(n11249), .B(n11248), .Z(n11253) );
  OR U12327 ( .A(n11251), .B(n11250), .Z(n11252) );
  AND U12328 ( .A(n11253), .B(n11252), .Z(n11271) );
  XOR U12329 ( .A(a[428]), .B(n2237), .Z(n11275) );
  AND U12330 ( .A(a[426]), .B(b[3]), .Z(n11279) );
  AND U12331 ( .A(a[430]), .B(b[0]), .Z(n11255) );
  XNOR U12332 ( .A(n11255), .B(n2175), .Z(n11257) );
  NANDN U12333 ( .A(b[0]), .B(a[429]), .Z(n11256) );
  NAND U12334 ( .A(n11257), .B(n11256), .Z(n11280) );
  XOR U12335 ( .A(n11279), .B(n11280), .Z(n11282) );
  XOR U12336 ( .A(n11281), .B(n11282), .Z(n11270) );
  NANDN U12337 ( .A(n11259), .B(n11258), .Z(n11263) );
  OR U12338 ( .A(n11261), .B(n11260), .Z(n11262) );
  AND U12339 ( .A(n11263), .B(n11262), .Z(n11269) );
  XOR U12340 ( .A(n11270), .B(n11269), .Z(n11272) );
  XOR U12341 ( .A(n11271), .B(n11272), .Z(n11285) );
  XNOR U12342 ( .A(n11285), .B(sreg[1450]), .Z(n11287) );
  NANDN U12343 ( .A(n11264), .B(sreg[1449]), .Z(n11268) );
  NAND U12344 ( .A(n11266), .B(n11265), .Z(n11267) );
  NAND U12345 ( .A(n11268), .B(n11267), .Z(n11286) );
  XOR U12346 ( .A(n11287), .B(n11286), .Z(c[1450]) );
  NANDN U12347 ( .A(n11270), .B(n11269), .Z(n11274) );
  OR U12348 ( .A(n11272), .B(n11271), .Z(n11273) );
  AND U12349 ( .A(n11274), .B(n11273), .Z(n11292) );
  XOR U12350 ( .A(a[429]), .B(n2237), .Z(n11296) );
  AND U12351 ( .A(a[431]), .B(b[0]), .Z(n11276) );
  XNOR U12352 ( .A(n11276), .B(n2175), .Z(n11278) );
  NANDN U12353 ( .A(b[0]), .B(a[430]), .Z(n11277) );
  NAND U12354 ( .A(n11278), .B(n11277), .Z(n11301) );
  AND U12355 ( .A(a[427]), .B(b[3]), .Z(n11300) );
  XOR U12356 ( .A(n11301), .B(n11300), .Z(n11303) );
  XOR U12357 ( .A(n11302), .B(n11303), .Z(n11291) );
  NANDN U12358 ( .A(n11280), .B(n11279), .Z(n11284) );
  OR U12359 ( .A(n11282), .B(n11281), .Z(n11283) );
  AND U12360 ( .A(n11284), .B(n11283), .Z(n11290) );
  XOR U12361 ( .A(n11291), .B(n11290), .Z(n11293) );
  XOR U12362 ( .A(n11292), .B(n11293), .Z(n11306) );
  XNOR U12363 ( .A(n11306), .B(sreg[1451]), .Z(n11308) );
  NANDN U12364 ( .A(n11285), .B(sreg[1450]), .Z(n11289) );
  NAND U12365 ( .A(n11287), .B(n11286), .Z(n11288) );
  NAND U12366 ( .A(n11289), .B(n11288), .Z(n11307) );
  XOR U12367 ( .A(n11308), .B(n11307), .Z(c[1451]) );
  NANDN U12368 ( .A(n11291), .B(n11290), .Z(n11295) );
  OR U12369 ( .A(n11293), .B(n11292), .Z(n11294) );
  AND U12370 ( .A(n11295), .B(n11294), .Z(n11313) );
  XOR U12371 ( .A(a[430]), .B(n2237), .Z(n11317) );
  AND U12372 ( .A(a[432]), .B(b[0]), .Z(n11297) );
  XNOR U12373 ( .A(n11297), .B(n2175), .Z(n11299) );
  NANDN U12374 ( .A(b[0]), .B(a[431]), .Z(n11298) );
  NAND U12375 ( .A(n11299), .B(n11298), .Z(n11322) );
  AND U12376 ( .A(a[428]), .B(b[3]), .Z(n11321) );
  XOR U12377 ( .A(n11322), .B(n11321), .Z(n11324) );
  XOR U12378 ( .A(n11323), .B(n11324), .Z(n11312) );
  NANDN U12379 ( .A(n11301), .B(n11300), .Z(n11305) );
  OR U12380 ( .A(n11303), .B(n11302), .Z(n11304) );
  AND U12381 ( .A(n11305), .B(n11304), .Z(n11311) );
  XOR U12382 ( .A(n11312), .B(n11311), .Z(n11314) );
  XOR U12383 ( .A(n11313), .B(n11314), .Z(n11327) );
  XNOR U12384 ( .A(n11327), .B(sreg[1452]), .Z(n11329) );
  NANDN U12385 ( .A(n11306), .B(sreg[1451]), .Z(n11310) );
  NAND U12386 ( .A(n11308), .B(n11307), .Z(n11309) );
  NAND U12387 ( .A(n11310), .B(n11309), .Z(n11328) );
  XOR U12388 ( .A(n11329), .B(n11328), .Z(c[1452]) );
  NANDN U12389 ( .A(n11312), .B(n11311), .Z(n11316) );
  OR U12390 ( .A(n11314), .B(n11313), .Z(n11315) );
  AND U12391 ( .A(n11316), .B(n11315), .Z(n11334) );
  XOR U12392 ( .A(a[431]), .B(n2237), .Z(n11338) );
  AND U12393 ( .A(a[429]), .B(b[3]), .Z(n11342) );
  AND U12394 ( .A(a[433]), .B(b[0]), .Z(n11318) );
  XNOR U12395 ( .A(n11318), .B(n2175), .Z(n11320) );
  NANDN U12396 ( .A(b[0]), .B(a[432]), .Z(n11319) );
  NAND U12397 ( .A(n11320), .B(n11319), .Z(n11343) );
  XOR U12398 ( .A(n11342), .B(n11343), .Z(n11345) );
  XOR U12399 ( .A(n11344), .B(n11345), .Z(n11333) );
  NANDN U12400 ( .A(n11322), .B(n11321), .Z(n11326) );
  OR U12401 ( .A(n11324), .B(n11323), .Z(n11325) );
  AND U12402 ( .A(n11326), .B(n11325), .Z(n11332) );
  XOR U12403 ( .A(n11333), .B(n11332), .Z(n11335) );
  XOR U12404 ( .A(n11334), .B(n11335), .Z(n11348) );
  XNOR U12405 ( .A(n11348), .B(sreg[1453]), .Z(n11350) );
  NANDN U12406 ( .A(n11327), .B(sreg[1452]), .Z(n11331) );
  NAND U12407 ( .A(n11329), .B(n11328), .Z(n11330) );
  NAND U12408 ( .A(n11331), .B(n11330), .Z(n11349) );
  XOR U12409 ( .A(n11350), .B(n11349), .Z(c[1453]) );
  NANDN U12410 ( .A(n11333), .B(n11332), .Z(n11337) );
  OR U12411 ( .A(n11335), .B(n11334), .Z(n11336) );
  AND U12412 ( .A(n11337), .B(n11336), .Z(n11355) );
  XOR U12413 ( .A(a[432]), .B(n2237), .Z(n11359) );
  AND U12414 ( .A(a[434]), .B(b[0]), .Z(n11339) );
  XNOR U12415 ( .A(n11339), .B(n2175), .Z(n11341) );
  NANDN U12416 ( .A(b[0]), .B(a[433]), .Z(n11340) );
  NAND U12417 ( .A(n11341), .B(n11340), .Z(n11364) );
  AND U12418 ( .A(a[430]), .B(b[3]), .Z(n11363) );
  XOR U12419 ( .A(n11364), .B(n11363), .Z(n11366) );
  XOR U12420 ( .A(n11365), .B(n11366), .Z(n11354) );
  NANDN U12421 ( .A(n11343), .B(n11342), .Z(n11347) );
  OR U12422 ( .A(n11345), .B(n11344), .Z(n11346) );
  AND U12423 ( .A(n11347), .B(n11346), .Z(n11353) );
  XOR U12424 ( .A(n11354), .B(n11353), .Z(n11356) );
  XOR U12425 ( .A(n11355), .B(n11356), .Z(n11369) );
  XNOR U12426 ( .A(n11369), .B(sreg[1454]), .Z(n11371) );
  NANDN U12427 ( .A(n11348), .B(sreg[1453]), .Z(n11352) );
  NAND U12428 ( .A(n11350), .B(n11349), .Z(n11351) );
  NAND U12429 ( .A(n11352), .B(n11351), .Z(n11370) );
  XOR U12430 ( .A(n11371), .B(n11370), .Z(c[1454]) );
  NANDN U12431 ( .A(n11354), .B(n11353), .Z(n11358) );
  OR U12432 ( .A(n11356), .B(n11355), .Z(n11357) );
  AND U12433 ( .A(n11358), .B(n11357), .Z(n11376) );
  XOR U12434 ( .A(a[433]), .B(n2238), .Z(n11380) );
  AND U12435 ( .A(a[435]), .B(b[0]), .Z(n11360) );
  XNOR U12436 ( .A(n11360), .B(n2175), .Z(n11362) );
  NANDN U12437 ( .A(b[0]), .B(a[434]), .Z(n11361) );
  NAND U12438 ( .A(n11362), .B(n11361), .Z(n11385) );
  AND U12439 ( .A(a[431]), .B(b[3]), .Z(n11384) );
  XOR U12440 ( .A(n11385), .B(n11384), .Z(n11387) );
  XOR U12441 ( .A(n11386), .B(n11387), .Z(n11375) );
  NANDN U12442 ( .A(n11364), .B(n11363), .Z(n11368) );
  OR U12443 ( .A(n11366), .B(n11365), .Z(n11367) );
  AND U12444 ( .A(n11368), .B(n11367), .Z(n11374) );
  XOR U12445 ( .A(n11375), .B(n11374), .Z(n11377) );
  XOR U12446 ( .A(n11376), .B(n11377), .Z(n11390) );
  XNOR U12447 ( .A(n11390), .B(sreg[1455]), .Z(n11392) );
  NANDN U12448 ( .A(n11369), .B(sreg[1454]), .Z(n11373) );
  NAND U12449 ( .A(n11371), .B(n11370), .Z(n11372) );
  NAND U12450 ( .A(n11373), .B(n11372), .Z(n11391) );
  XOR U12451 ( .A(n11392), .B(n11391), .Z(c[1455]) );
  NANDN U12452 ( .A(n11375), .B(n11374), .Z(n11379) );
  OR U12453 ( .A(n11377), .B(n11376), .Z(n11378) );
  AND U12454 ( .A(n11379), .B(n11378), .Z(n11397) );
  XOR U12455 ( .A(a[434]), .B(n2238), .Z(n11401) );
  AND U12456 ( .A(a[432]), .B(b[3]), .Z(n11405) );
  AND U12457 ( .A(a[436]), .B(b[0]), .Z(n11381) );
  XNOR U12458 ( .A(n11381), .B(n2175), .Z(n11383) );
  NANDN U12459 ( .A(b[0]), .B(a[435]), .Z(n11382) );
  NAND U12460 ( .A(n11383), .B(n11382), .Z(n11406) );
  XOR U12461 ( .A(n11405), .B(n11406), .Z(n11408) );
  XOR U12462 ( .A(n11407), .B(n11408), .Z(n11396) );
  NANDN U12463 ( .A(n11385), .B(n11384), .Z(n11389) );
  OR U12464 ( .A(n11387), .B(n11386), .Z(n11388) );
  AND U12465 ( .A(n11389), .B(n11388), .Z(n11395) );
  XOR U12466 ( .A(n11396), .B(n11395), .Z(n11398) );
  XOR U12467 ( .A(n11397), .B(n11398), .Z(n11411) );
  XNOR U12468 ( .A(n11411), .B(sreg[1456]), .Z(n11413) );
  NANDN U12469 ( .A(n11390), .B(sreg[1455]), .Z(n11394) );
  NAND U12470 ( .A(n11392), .B(n11391), .Z(n11393) );
  NAND U12471 ( .A(n11394), .B(n11393), .Z(n11412) );
  XOR U12472 ( .A(n11413), .B(n11412), .Z(c[1456]) );
  NANDN U12473 ( .A(n11396), .B(n11395), .Z(n11400) );
  OR U12474 ( .A(n11398), .B(n11397), .Z(n11399) );
  AND U12475 ( .A(n11400), .B(n11399), .Z(n11418) );
  XOR U12476 ( .A(a[435]), .B(n2238), .Z(n11422) );
  AND U12477 ( .A(a[437]), .B(b[0]), .Z(n11402) );
  XNOR U12478 ( .A(n11402), .B(n2175), .Z(n11404) );
  NANDN U12479 ( .A(b[0]), .B(a[436]), .Z(n11403) );
  NAND U12480 ( .A(n11404), .B(n11403), .Z(n11427) );
  AND U12481 ( .A(a[433]), .B(b[3]), .Z(n11426) );
  XOR U12482 ( .A(n11427), .B(n11426), .Z(n11429) );
  XOR U12483 ( .A(n11428), .B(n11429), .Z(n11417) );
  NANDN U12484 ( .A(n11406), .B(n11405), .Z(n11410) );
  OR U12485 ( .A(n11408), .B(n11407), .Z(n11409) );
  AND U12486 ( .A(n11410), .B(n11409), .Z(n11416) );
  XOR U12487 ( .A(n11417), .B(n11416), .Z(n11419) );
  XOR U12488 ( .A(n11418), .B(n11419), .Z(n11432) );
  XNOR U12489 ( .A(n11432), .B(sreg[1457]), .Z(n11434) );
  NANDN U12490 ( .A(n11411), .B(sreg[1456]), .Z(n11415) );
  NAND U12491 ( .A(n11413), .B(n11412), .Z(n11414) );
  NAND U12492 ( .A(n11415), .B(n11414), .Z(n11433) );
  XOR U12493 ( .A(n11434), .B(n11433), .Z(c[1457]) );
  NANDN U12494 ( .A(n11417), .B(n11416), .Z(n11421) );
  OR U12495 ( .A(n11419), .B(n11418), .Z(n11420) );
  AND U12496 ( .A(n11421), .B(n11420), .Z(n11439) );
  XOR U12497 ( .A(a[436]), .B(n2238), .Z(n11443) );
  AND U12498 ( .A(a[434]), .B(b[3]), .Z(n11447) );
  AND U12499 ( .A(a[438]), .B(b[0]), .Z(n11423) );
  XNOR U12500 ( .A(n11423), .B(n2175), .Z(n11425) );
  NANDN U12501 ( .A(b[0]), .B(a[437]), .Z(n11424) );
  NAND U12502 ( .A(n11425), .B(n11424), .Z(n11448) );
  XOR U12503 ( .A(n11447), .B(n11448), .Z(n11450) );
  XOR U12504 ( .A(n11449), .B(n11450), .Z(n11438) );
  NANDN U12505 ( .A(n11427), .B(n11426), .Z(n11431) );
  OR U12506 ( .A(n11429), .B(n11428), .Z(n11430) );
  AND U12507 ( .A(n11431), .B(n11430), .Z(n11437) );
  XOR U12508 ( .A(n11438), .B(n11437), .Z(n11440) );
  XOR U12509 ( .A(n11439), .B(n11440), .Z(n11453) );
  XNOR U12510 ( .A(n11453), .B(sreg[1458]), .Z(n11455) );
  NANDN U12511 ( .A(n11432), .B(sreg[1457]), .Z(n11436) );
  NAND U12512 ( .A(n11434), .B(n11433), .Z(n11435) );
  NAND U12513 ( .A(n11436), .B(n11435), .Z(n11454) );
  XOR U12514 ( .A(n11455), .B(n11454), .Z(c[1458]) );
  NANDN U12515 ( .A(n11438), .B(n11437), .Z(n11442) );
  OR U12516 ( .A(n11440), .B(n11439), .Z(n11441) );
  AND U12517 ( .A(n11442), .B(n11441), .Z(n11460) );
  XOR U12518 ( .A(a[437]), .B(n2238), .Z(n11464) );
  AND U12519 ( .A(a[439]), .B(b[0]), .Z(n11444) );
  XNOR U12520 ( .A(n11444), .B(n2175), .Z(n11446) );
  NANDN U12521 ( .A(b[0]), .B(a[438]), .Z(n11445) );
  NAND U12522 ( .A(n11446), .B(n11445), .Z(n11469) );
  AND U12523 ( .A(a[435]), .B(b[3]), .Z(n11468) );
  XOR U12524 ( .A(n11469), .B(n11468), .Z(n11471) );
  XOR U12525 ( .A(n11470), .B(n11471), .Z(n11459) );
  NANDN U12526 ( .A(n11448), .B(n11447), .Z(n11452) );
  OR U12527 ( .A(n11450), .B(n11449), .Z(n11451) );
  AND U12528 ( .A(n11452), .B(n11451), .Z(n11458) );
  XOR U12529 ( .A(n11459), .B(n11458), .Z(n11461) );
  XOR U12530 ( .A(n11460), .B(n11461), .Z(n11474) );
  XNOR U12531 ( .A(n11474), .B(sreg[1459]), .Z(n11476) );
  NANDN U12532 ( .A(n11453), .B(sreg[1458]), .Z(n11457) );
  NAND U12533 ( .A(n11455), .B(n11454), .Z(n11456) );
  NAND U12534 ( .A(n11457), .B(n11456), .Z(n11475) );
  XOR U12535 ( .A(n11476), .B(n11475), .Z(c[1459]) );
  NANDN U12536 ( .A(n11459), .B(n11458), .Z(n11463) );
  OR U12537 ( .A(n11461), .B(n11460), .Z(n11462) );
  AND U12538 ( .A(n11463), .B(n11462), .Z(n11481) );
  XOR U12539 ( .A(a[438]), .B(n2238), .Z(n11485) );
  AND U12540 ( .A(a[436]), .B(b[3]), .Z(n11489) );
  AND U12541 ( .A(a[440]), .B(b[0]), .Z(n11465) );
  XNOR U12542 ( .A(n11465), .B(n2175), .Z(n11467) );
  NANDN U12543 ( .A(b[0]), .B(a[439]), .Z(n11466) );
  NAND U12544 ( .A(n11467), .B(n11466), .Z(n11490) );
  XOR U12545 ( .A(n11489), .B(n11490), .Z(n11492) );
  XOR U12546 ( .A(n11491), .B(n11492), .Z(n11480) );
  NANDN U12547 ( .A(n11469), .B(n11468), .Z(n11473) );
  OR U12548 ( .A(n11471), .B(n11470), .Z(n11472) );
  AND U12549 ( .A(n11473), .B(n11472), .Z(n11479) );
  XOR U12550 ( .A(n11480), .B(n11479), .Z(n11482) );
  XOR U12551 ( .A(n11481), .B(n11482), .Z(n11495) );
  XNOR U12552 ( .A(n11495), .B(sreg[1460]), .Z(n11497) );
  NANDN U12553 ( .A(n11474), .B(sreg[1459]), .Z(n11478) );
  NAND U12554 ( .A(n11476), .B(n11475), .Z(n11477) );
  NAND U12555 ( .A(n11478), .B(n11477), .Z(n11496) );
  XOR U12556 ( .A(n11497), .B(n11496), .Z(c[1460]) );
  NANDN U12557 ( .A(n11480), .B(n11479), .Z(n11484) );
  OR U12558 ( .A(n11482), .B(n11481), .Z(n11483) );
  AND U12559 ( .A(n11484), .B(n11483), .Z(n11502) );
  XOR U12560 ( .A(a[439]), .B(n2238), .Z(n11506) );
  AND U12561 ( .A(a[437]), .B(b[3]), .Z(n11510) );
  AND U12562 ( .A(a[441]), .B(b[0]), .Z(n11486) );
  XNOR U12563 ( .A(n11486), .B(n2175), .Z(n11488) );
  NANDN U12564 ( .A(b[0]), .B(a[440]), .Z(n11487) );
  NAND U12565 ( .A(n11488), .B(n11487), .Z(n11511) );
  XOR U12566 ( .A(n11510), .B(n11511), .Z(n11513) );
  XOR U12567 ( .A(n11512), .B(n11513), .Z(n11501) );
  NANDN U12568 ( .A(n11490), .B(n11489), .Z(n11494) );
  OR U12569 ( .A(n11492), .B(n11491), .Z(n11493) );
  AND U12570 ( .A(n11494), .B(n11493), .Z(n11500) );
  XOR U12571 ( .A(n11501), .B(n11500), .Z(n11503) );
  XOR U12572 ( .A(n11502), .B(n11503), .Z(n11516) );
  XNOR U12573 ( .A(n11516), .B(sreg[1461]), .Z(n11518) );
  NANDN U12574 ( .A(n11495), .B(sreg[1460]), .Z(n11499) );
  NAND U12575 ( .A(n11497), .B(n11496), .Z(n11498) );
  NAND U12576 ( .A(n11499), .B(n11498), .Z(n11517) );
  XOR U12577 ( .A(n11518), .B(n11517), .Z(c[1461]) );
  NANDN U12578 ( .A(n11501), .B(n11500), .Z(n11505) );
  OR U12579 ( .A(n11503), .B(n11502), .Z(n11504) );
  AND U12580 ( .A(n11505), .B(n11504), .Z(n11523) );
  XOR U12581 ( .A(a[440]), .B(n2239), .Z(n11527) );
  AND U12582 ( .A(a[442]), .B(b[0]), .Z(n11507) );
  XNOR U12583 ( .A(n11507), .B(n2175), .Z(n11509) );
  NANDN U12584 ( .A(b[0]), .B(a[441]), .Z(n11508) );
  NAND U12585 ( .A(n11509), .B(n11508), .Z(n11532) );
  AND U12586 ( .A(a[438]), .B(b[3]), .Z(n11531) );
  XOR U12587 ( .A(n11532), .B(n11531), .Z(n11534) );
  XOR U12588 ( .A(n11533), .B(n11534), .Z(n11522) );
  NANDN U12589 ( .A(n11511), .B(n11510), .Z(n11515) );
  OR U12590 ( .A(n11513), .B(n11512), .Z(n11514) );
  AND U12591 ( .A(n11515), .B(n11514), .Z(n11521) );
  XOR U12592 ( .A(n11522), .B(n11521), .Z(n11524) );
  XOR U12593 ( .A(n11523), .B(n11524), .Z(n11537) );
  XNOR U12594 ( .A(n11537), .B(sreg[1462]), .Z(n11539) );
  NANDN U12595 ( .A(n11516), .B(sreg[1461]), .Z(n11520) );
  NAND U12596 ( .A(n11518), .B(n11517), .Z(n11519) );
  NAND U12597 ( .A(n11520), .B(n11519), .Z(n11538) );
  XOR U12598 ( .A(n11539), .B(n11538), .Z(c[1462]) );
  NANDN U12599 ( .A(n11522), .B(n11521), .Z(n11526) );
  OR U12600 ( .A(n11524), .B(n11523), .Z(n11525) );
  AND U12601 ( .A(n11526), .B(n11525), .Z(n11544) );
  XOR U12602 ( .A(a[441]), .B(n2239), .Z(n11548) );
  AND U12603 ( .A(a[443]), .B(b[0]), .Z(n11528) );
  XNOR U12604 ( .A(n11528), .B(n2175), .Z(n11530) );
  NANDN U12605 ( .A(b[0]), .B(a[442]), .Z(n11529) );
  NAND U12606 ( .A(n11530), .B(n11529), .Z(n11553) );
  AND U12607 ( .A(a[439]), .B(b[3]), .Z(n11552) );
  XOR U12608 ( .A(n11553), .B(n11552), .Z(n11555) );
  XOR U12609 ( .A(n11554), .B(n11555), .Z(n11543) );
  NANDN U12610 ( .A(n11532), .B(n11531), .Z(n11536) );
  OR U12611 ( .A(n11534), .B(n11533), .Z(n11535) );
  AND U12612 ( .A(n11536), .B(n11535), .Z(n11542) );
  XOR U12613 ( .A(n11543), .B(n11542), .Z(n11545) );
  XOR U12614 ( .A(n11544), .B(n11545), .Z(n11558) );
  XNOR U12615 ( .A(n11558), .B(sreg[1463]), .Z(n11560) );
  NANDN U12616 ( .A(n11537), .B(sreg[1462]), .Z(n11541) );
  NAND U12617 ( .A(n11539), .B(n11538), .Z(n11540) );
  NAND U12618 ( .A(n11541), .B(n11540), .Z(n11559) );
  XOR U12619 ( .A(n11560), .B(n11559), .Z(c[1463]) );
  NANDN U12620 ( .A(n11543), .B(n11542), .Z(n11547) );
  OR U12621 ( .A(n11545), .B(n11544), .Z(n11546) );
  AND U12622 ( .A(n11547), .B(n11546), .Z(n11565) );
  XOR U12623 ( .A(a[442]), .B(n2239), .Z(n11569) );
  AND U12624 ( .A(a[440]), .B(b[3]), .Z(n11573) );
  AND U12625 ( .A(a[444]), .B(b[0]), .Z(n11549) );
  XNOR U12626 ( .A(n11549), .B(n2175), .Z(n11551) );
  NANDN U12627 ( .A(b[0]), .B(a[443]), .Z(n11550) );
  NAND U12628 ( .A(n11551), .B(n11550), .Z(n11574) );
  XOR U12629 ( .A(n11573), .B(n11574), .Z(n11576) );
  XOR U12630 ( .A(n11575), .B(n11576), .Z(n11564) );
  NANDN U12631 ( .A(n11553), .B(n11552), .Z(n11557) );
  OR U12632 ( .A(n11555), .B(n11554), .Z(n11556) );
  AND U12633 ( .A(n11557), .B(n11556), .Z(n11563) );
  XOR U12634 ( .A(n11564), .B(n11563), .Z(n11566) );
  XOR U12635 ( .A(n11565), .B(n11566), .Z(n11579) );
  XNOR U12636 ( .A(n11579), .B(sreg[1464]), .Z(n11581) );
  NANDN U12637 ( .A(n11558), .B(sreg[1463]), .Z(n11562) );
  NAND U12638 ( .A(n11560), .B(n11559), .Z(n11561) );
  NAND U12639 ( .A(n11562), .B(n11561), .Z(n11580) );
  XOR U12640 ( .A(n11581), .B(n11580), .Z(c[1464]) );
  NANDN U12641 ( .A(n11564), .B(n11563), .Z(n11568) );
  OR U12642 ( .A(n11566), .B(n11565), .Z(n11567) );
  AND U12643 ( .A(n11568), .B(n11567), .Z(n11586) );
  XOR U12644 ( .A(a[443]), .B(n2239), .Z(n11590) );
  AND U12645 ( .A(a[441]), .B(b[3]), .Z(n11594) );
  AND U12646 ( .A(a[445]), .B(b[0]), .Z(n11570) );
  XNOR U12647 ( .A(n11570), .B(n2175), .Z(n11572) );
  NANDN U12648 ( .A(b[0]), .B(a[444]), .Z(n11571) );
  NAND U12649 ( .A(n11572), .B(n11571), .Z(n11595) );
  XOR U12650 ( .A(n11594), .B(n11595), .Z(n11597) );
  XOR U12651 ( .A(n11596), .B(n11597), .Z(n11585) );
  NANDN U12652 ( .A(n11574), .B(n11573), .Z(n11578) );
  OR U12653 ( .A(n11576), .B(n11575), .Z(n11577) );
  AND U12654 ( .A(n11578), .B(n11577), .Z(n11584) );
  XOR U12655 ( .A(n11585), .B(n11584), .Z(n11587) );
  XOR U12656 ( .A(n11586), .B(n11587), .Z(n11600) );
  XNOR U12657 ( .A(n11600), .B(sreg[1465]), .Z(n11602) );
  NANDN U12658 ( .A(n11579), .B(sreg[1464]), .Z(n11583) );
  NAND U12659 ( .A(n11581), .B(n11580), .Z(n11582) );
  NAND U12660 ( .A(n11583), .B(n11582), .Z(n11601) );
  XOR U12661 ( .A(n11602), .B(n11601), .Z(c[1465]) );
  NANDN U12662 ( .A(n11585), .B(n11584), .Z(n11589) );
  OR U12663 ( .A(n11587), .B(n11586), .Z(n11588) );
  AND U12664 ( .A(n11589), .B(n11588), .Z(n11607) );
  XOR U12665 ( .A(a[444]), .B(n2239), .Z(n11611) );
  AND U12666 ( .A(a[446]), .B(b[0]), .Z(n11591) );
  XNOR U12667 ( .A(n11591), .B(n2175), .Z(n11593) );
  NANDN U12668 ( .A(b[0]), .B(a[445]), .Z(n11592) );
  NAND U12669 ( .A(n11593), .B(n11592), .Z(n11616) );
  AND U12670 ( .A(a[442]), .B(b[3]), .Z(n11615) );
  XOR U12671 ( .A(n11616), .B(n11615), .Z(n11618) );
  XOR U12672 ( .A(n11617), .B(n11618), .Z(n11606) );
  NANDN U12673 ( .A(n11595), .B(n11594), .Z(n11599) );
  OR U12674 ( .A(n11597), .B(n11596), .Z(n11598) );
  AND U12675 ( .A(n11599), .B(n11598), .Z(n11605) );
  XOR U12676 ( .A(n11606), .B(n11605), .Z(n11608) );
  XOR U12677 ( .A(n11607), .B(n11608), .Z(n11621) );
  XNOR U12678 ( .A(n11621), .B(sreg[1466]), .Z(n11623) );
  NANDN U12679 ( .A(n11600), .B(sreg[1465]), .Z(n11604) );
  NAND U12680 ( .A(n11602), .B(n11601), .Z(n11603) );
  NAND U12681 ( .A(n11604), .B(n11603), .Z(n11622) );
  XOR U12682 ( .A(n11623), .B(n11622), .Z(c[1466]) );
  NANDN U12683 ( .A(n11606), .B(n11605), .Z(n11610) );
  OR U12684 ( .A(n11608), .B(n11607), .Z(n11609) );
  AND U12685 ( .A(n11610), .B(n11609), .Z(n11628) );
  XOR U12686 ( .A(a[445]), .B(n2239), .Z(n11632) );
  AND U12687 ( .A(a[443]), .B(b[3]), .Z(n11636) );
  AND U12688 ( .A(a[447]), .B(b[0]), .Z(n11612) );
  XNOR U12689 ( .A(n11612), .B(n2175), .Z(n11614) );
  NANDN U12690 ( .A(b[0]), .B(a[446]), .Z(n11613) );
  NAND U12691 ( .A(n11614), .B(n11613), .Z(n11637) );
  XOR U12692 ( .A(n11636), .B(n11637), .Z(n11639) );
  XOR U12693 ( .A(n11638), .B(n11639), .Z(n11627) );
  NANDN U12694 ( .A(n11616), .B(n11615), .Z(n11620) );
  OR U12695 ( .A(n11618), .B(n11617), .Z(n11619) );
  AND U12696 ( .A(n11620), .B(n11619), .Z(n11626) );
  XOR U12697 ( .A(n11627), .B(n11626), .Z(n11629) );
  XOR U12698 ( .A(n11628), .B(n11629), .Z(n11642) );
  XNOR U12699 ( .A(n11642), .B(sreg[1467]), .Z(n11644) );
  NANDN U12700 ( .A(n11621), .B(sreg[1466]), .Z(n11625) );
  NAND U12701 ( .A(n11623), .B(n11622), .Z(n11624) );
  NAND U12702 ( .A(n11625), .B(n11624), .Z(n11643) );
  XOR U12703 ( .A(n11644), .B(n11643), .Z(c[1467]) );
  NANDN U12704 ( .A(n11627), .B(n11626), .Z(n11631) );
  OR U12705 ( .A(n11629), .B(n11628), .Z(n11630) );
  AND U12706 ( .A(n11631), .B(n11630), .Z(n11649) );
  XOR U12707 ( .A(a[446]), .B(n2239), .Z(n11653) );
  AND U12708 ( .A(a[448]), .B(b[0]), .Z(n11633) );
  XNOR U12709 ( .A(n11633), .B(n2175), .Z(n11635) );
  NANDN U12710 ( .A(b[0]), .B(a[447]), .Z(n11634) );
  NAND U12711 ( .A(n11635), .B(n11634), .Z(n11658) );
  AND U12712 ( .A(a[444]), .B(b[3]), .Z(n11657) );
  XOR U12713 ( .A(n11658), .B(n11657), .Z(n11660) );
  XOR U12714 ( .A(n11659), .B(n11660), .Z(n11648) );
  NANDN U12715 ( .A(n11637), .B(n11636), .Z(n11641) );
  OR U12716 ( .A(n11639), .B(n11638), .Z(n11640) );
  AND U12717 ( .A(n11641), .B(n11640), .Z(n11647) );
  XOR U12718 ( .A(n11648), .B(n11647), .Z(n11650) );
  XOR U12719 ( .A(n11649), .B(n11650), .Z(n11663) );
  XNOR U12720 ( .A(n11663), .B(sreg[1468]), .Z(n11665) );
  NANDN U12721 ( .A(n11642), .B(sreg[1467]), .Z(n11646) );
  NAND U12722 ( .A(n11644), .B(n11643), .Z(n11645) );
  NAND U12723 ( .A(n11646), .B(n11645), .Z(n11664) );
  XOR U12724 ( .A(n11665), .B(n11664), .Z(c[1468]) );
  NANDN U12725 ( .A(n11648), .B(n11647), .Z(n11652) );
  OR U12726 ( .A(n11650), .B(n11649), .Z(n11651) );
  AND U12727 ( .A(n11652), .B(n11651), .Z(n11670) );
  XOR U12728 ( .A(a[447]), .B(n2240), .Z(n11674) );
  AND U12729 ( .A(a[445]), .B(b[3]), .Z(n11678) );
  AND U12730 ( .A(a[449]), .B(b[0]), .Z(n11654) );
  XNOR U12731 ( .A(n11654), .B(n2175), .Z(n11656) );
  NANDN U12732 ( .A(b[0]), .B(a[448]), .Z(n11655) );
  NAND U12733 ( .A(n11656), .B(n11655), .Z(n11679) );
  XOR U12734 ( .A(n11678), .B(n11679), .Z(n11681) );
  XOR U12735 ( .A(n11680), .B(n11681), .Z(n11669) );
  NANDN U12736 ( .A(n11658), .B(n11657), .Z(n11662) );
  OR U12737 ( .A(n11660), .B(n11659), .Z(n11661) );
  AND U12738 ( .A(n11662), .B(n11661), .Z(n11668) );
  XOR U12739 ( .A(n11669), .B(n11668), .Z(n11671) );
  XOR U12740 ( .A(n11670), .B(n11671), .Z(n11684) );
  XNOR U12741 ( .A(n11684), .B(sreg[1469]), .Z(n11686) );
  NANDN U12742 ( .A(n11663), .B(sreg[1468]), .Z(n11667) );
  NAND U12743 ( .A(n11665), .B(n11664), .Z(n11666) );
  NAND U12744 ( .A(n11667), .B(n11666), .Z(n11685) );
  XOR U12745 ( .A(n11686), .B(n11685), .Z(c[1469]) );
  NANDN U12746 ( .A(n11669), .B(n11668), .Z(n11673) );
  OR U12747 ( .A(n11671), .B(n11670), .Z(n11672) );
  AND U12748 ( .A(n11673), .B(n11672), .Z(n11691) );
  XOR U12749 ( .A(a[448]), .B(n2240), .Z(n11695) );
  AND U12750 ( .A(a[450]), .B(b[0]), .Z(n11675) );
  XNOR U12751 ( .A(n11675), .B(n2175), .Z(n11677) );
  NANDN U12752 ( .A(b[0]), .B(a[449]), .Z(n11676) );
  NAND U12753 ( .A(n11677), .B(n11676), .Z(n11700) );
  AND U12754 ( .A(a[446]), .B(b[3]), .Z(n11699) );
  XOR U12755 ( .A(n11700), .B(n11699), .Z(n11702) );
  XOR U12756 ( .A(n11701), .B(n11702), .Z(n11690) );
  NANDN U12757 ( .A(n11679), .B(n11678), .Z(n11683) );
  OR U12758 ( .A(n11681), .B(n11680), .Z(n11682) );
  AND U12759 ( .A(n11683), .B(n11682), .Z(n11689) );
  XOR U12760 ( .A(n11690), .B(n11689), .Z(n11692) );
  XOR U12761 ( .A(n11691), .B(n11692), .Z(n11705) );
  XNOR U12762 ( .A(n11705), .B(sreg[1470]), .Z(n11707) );
  NANDN U12763 ( .A(n11684), .B(sreg[1469]), .Z(n11688) );
  NAND U12764 ( .A(n11686), .B(n11685), .Z(n11687) );
  NAND U12765 ( .A(n11688), .B(n11687), .Z(n11706) );
  XOR U12766 ( .A(n11707), .B(n11706), .Z(c[1470]) );
  NANDN U12767 ( .A(n11690), .B(n11689), .Z(n11694) );
  OR U12768 ( .A(n11692), .B(n11691), .Z(n11693) );
  AND U12769 ( .A(n11694), .B(n11693), .Z(n11712) );
  XOR U12770 ( .A(a[449]), .B(n2240), .Z(n11716) );
  AND U12771 ( .A(a[451]), .B(b[0]), .Z(n11696) );
  XNOR U12772 ( .A(n11696), .B(n2175), .Z(n11698) );
  NANDN U12773 ( .A(b[0]), .B(a[450]), .Z(n11697) );
  NAND U12774 ( .A(n11698), .B(n11697), .Z(n11721) );
  AND U12775 ( .A(a[447]), .B(b[3]), .Z(n11720) );
  XOR U12776 ( .A(n11721), .B(n11720), .Z(n11723) );
  XOR U12777 ( .A(n11722), .B(n11723), .Z(n11711) );
  NANDN U12778 ( .A(n11700), .B(n11699), .Z(n11704) );
  OR U12779 ( .A(n11702), .B(n11701), .Z(n11703) );
  AND U12780 ( .A(n11704), .B(n11703), .Z(n11710) );
  XOR U12781 ( .A(n11711), .B(n11710), .Z(n11713) );
  XOR U12782 ( .A(n11712), .B(n11713), .Z(n11726) );
  XNOR U12783 ( .A(n11726), .B(sreg[1471]), .Z(n11728) );
  NANDN U12784 ( .A(n11705), .B(sreg[1470]), .Z(n11709) );
  NAND U12785 ( .A(n11707), .B(n11706), .Z(n11708) );
  NAND U12786 ( .A(n11709), .B(n11708), .Z(n11727) );
  XOR U12787 ( .A(n11728), .B(n11727), .Z(c[1471]) );
  NANDN U12788 ( .A(n11711), .B(n11710), .Z(n11715) );
  OR U12789 ( .A(n11713), .B(n11712), .Z(n11714) );
  AND U12790 ( .A(n11715), .B(n11714), .Z(n11733) );
  XOR U12791 ( .A(a[450]), .B(n2240), .Z(n11737) );
  AND U12792 ( .A(a[452]), .B(b[0]), .Z(n11717) );
  XNOR U12793 ( .A(n11717), .B(n2175), .Z(n11719) );
  NANDN U12794 ( .A(b[0]), .B(a[451]), .Z(n11718) );
  NAND U12795 ( .A(n11719), .B(n11718), .Z(n11742) );
  AND U12796 ( .A(a[448]), .B(b[3]), .Z(n11741) );
  XOR U12797 ( .A(n11742), .B(n11741), .Z(n11744) );
  XOR U12798 ( .A(n11743), .B(n11744), .Z(n11732) );
  NANDN U12799 ( .A(n11721), .B(n11720), .Z(n11725) );
  OR U12800 ( .A(n11723), .B(n11722), .Z(n11724) );
  AND U12801 ( .A(n11725), .B(n11724), .Z(n11731) );
  XOR U12802 ( .A(n11732), .B(n11731), .Z(n11734) );
  XOR U12803 ( .A(n11733), .B(n11734), .Z(n11747) );
  XNOR U12804 ( .A(n11747), .B(sreg[1472]), .Z(n11749) );
  NANDN U12805 ( .A(n11726), .B(sreg[1471]), .Z(n11730) );
  NAND U12806 ( .A(n11728), .B(n11727), .Z(n11729) );
  NAND U12807 ( .A(n11730), .B(n11729), .Z(n11748) );
  XOR U12808 ( .A(n11749), .B(n11748), .Z(c[1472]) );
  NANDN U12809 ( .A(n11732), .B(n11731), .Z(n11736) );
  OR U12810 ( .A(n11734), .B(n11733), .Z(n11735) );
  AND U12811 ( .A(n11736), .B(n11735), .Z(n11755) );
  XOR U12812 ( .A(a[451]), .B(n2240), .Z(n11756) );
  AND U12813 ( .A(b[0]), .B(a[453]), .Z(n11738) );
  XOR U12814 ( .A(b[1]), .B(n11738), .Z(n11740) );
  NANDN U12815 ( .A(b[0]), .B(a[452]), .Z(n11739) );
  AND U12816 ( .A(n11740), .B(n11739), .Z(n11760) );
  AND U12817 ( .A(a[449]), .B(b[3]), .Z(n11761) );
  XOR U12818 ( .A(n11760), .B(n11761), .Z(n11762) );
  XNOR U12819 ( .A(n11763), .B(n11762), .Z(n11752) );
  NANDN U12820 ( .A(n11742), .B(n11741), .Z(n11746) );
  OR U12821 ( .A(n11744), .B(n11743), .Z(n11745) );
  AND U12822 ( .A(n11746), .B(n11745), .Z(n11753) );
  XNOR U12823 ( .A(n11752), .B(n11753), .Z(n11754) );
  XNOR U12824 ( .A(n11755), .B(n11754), .Z(n11766) );
  XNOR U12825 ( .A(n11766), .B(sreg[1473]), .Z(n11768) );
  NANDN U12826 ( .A(n11747), .B(sreg[1472]), .Z(n11751) );
  NAND U12827 ( .A(n11749), .B(n11748), .Z(n11750) );
  NAND U12828 ( .A(n11751), .B(n11750), .Z(n11767) );
  XOR U12829 ( .A(n11768), .B(n11767), .Z(c[1473]) );
  XOR U12830 ( .A(a[452]), .B(n2240), .Z(n11775) );
  AND U12831 ( .A(a[454]), .B(b[0]), .Z(n11757) );
  XNOR U12832 ( .A(n11757), .B(n2175), .Z(n11759) );
  NANDN U12833 ( .A(b[0]), .B(a[453]), .Z(n11758) );
  NAND U12834 ( .A(n11759), .B(n11758), .Z(n11780) );
  AND U12835 ( .A(a[450]), .B(b[3]), .Z(n11779) );
  XOR U12836 ( .A(n11780), .B(n11779), .Z(n11782) );
  XOR U12837 ( .A(n11781), .B(n11782), .Z(n11770) );
  NAND U12838 ( .A(n11761), .B(n11760), .Z(n11765) );
  NANDN U12839 ( .A(n11763), .B(n11762), .Z(n11764) );
  AND U12840 ( .A(n11765), .B(n11764), .Z(n11769) );
  XOR U12841 ( .A(n11770), .B(n11769), .Z(n11772) );
  XOR U12842 ( .A(n11771), .B(n11772), .Z(n11785) );
  XNOR U12843 ( .A(n11785), .B(sreg[1474]), .Z(n11787) );
  XOR U12844 ( .A(n11787), .B(n11786), .Z(c[1474]) );
  NANDN U12845 ( .A(n11770), .B(n11769), .Z(n11774) );
  OR U12846 ( .A(n11772), .B(n11771), .Z(n11773) );
  AND U12847 ( .A(n11774), .B(n11773), .Z(n11793) );
  XOR U12848 ( .A(a[453]), .B(n2240), .Z(n11794) );
  AND U12849 ( .A(b[0]), .B(a[455]), .Z(n11776) );
  XOR U12850 ( .A(b[1]), .B(n11776), .Z(n11778) );
  ANDN U12851 ( .B(b[1]), .A(b[0]), .Z(n23588) );
  NAND U12852 ( .A(n23588), .B(a[454]), .Z(n11777) );
  AND U12853 ( .A(n11778), .B(n11777), .Z(n11798) );
  AND U12854 ( .A(a[451]), .B(b[3]), .Z(n11799) );
  XOR U12855 ( .A(n11798), .B(n11799), .Z(n11800) );
  XNOR U12856 ( .A(n11801), .B(n11800), .Z(n11790) );
  NANDN U12857 ( .A(n11780), .B(n11779), .Z(n11784) );
  OR U12858 ( .A(n11782), .B(n11781), .Z(n11783) );
  AND U12859 ( .A(n11784), .B(n11783), .Z(n11791) );
  XNOR U12860 ( .A(n11790), .B(n11791), .Z(n11792) );
  XNOR U12861 ( .A(n11793), .B(n11792), .Z(n11804) );
  XNOR U12862 ( .A(n11804), .B(sreg[1475]), .Z(n11806) );
  NANDN U12863 ( .A(n11785), .B(sreg[1474]), .Z(n11789) );
  NAND U12864 ( .A(n11787), .B(n11786), .Z(n11788) );
  NAND U12865 ( .A(n11789), .B(n11788), .Z(n11805) );
  XOR U12866 ( .A(n11806), .B(n11805), .Z(c[1475]) );
  XOR U12867 ( .A(a[454]), .B(n2241), .Z(n11813) );
  AND U12868 ( .A(a[456]), .B(b[0]), .Z(n11795) );
  XNOR U12869 ( .A(n11795), .B(n2175), .Z(n11797) );
  NANDN U12870 ( .A(b[0]), .B(a[455]), .Z(n11796) );
  NAND U12871 ( .A(n11797), .B(n11796), .Z(n11818) );
  AND U12872 ( .A(a[452]), .B(b[3]), .Z(n11817) );
  XOR U12873 ( .A(n11818), .B(n11817), .Z(n11820) );
  XOR U12874 ( .A(n11819), .B(n11820), .Z(n11808) );
  NAND U12875 ( .A(n11799), .B(n11798), .Z(n11803) );
  NANDN U12876 ( .A(n11801), .B(n11800), .Z(n11802) );
  AND U12877 ( .A(n11803), .B(n11802), .Z(n11807) );
  XOR U12878 ( .A(n11808), .B(n11807), .Z(n11810) );
  XOR U12879 ( .A(n11809), .B(n11810), .Z(n11823) );
  XNOR U12880 ( .A(n11823), .B(sreg[1476]), .Z(n11825) );
  XOR U12881 ( .A(n11825), .B(n11824), .Z(c[1476]) );
  NANDN U12882 ( .A(n11808), .B(n11807), .Z(n11812) );
  OR U12883 ( .A(n11810), .B(n11809), .Z(n11811) );
  AND U12884 ( .A(n11812), .B(n11811), .Z(n11830) );
  XOR U12885 ( .A(a[455]), .B(n2241), .Z(n11834) );
  AND U12886 ( .A(a[457]), .B(b[0]), .Z(n11814) );
  XNOR U12887 ( .A(n11814), .B(n2175), .Z(n11816) );
  NANDN U12888 ( .A(b[0]), .B(a[456]), .Z(n11815) );
  NAND U12889 ( .A(n11816), .B(n11815), .Z(n11839) );
  AND U12890 ( .A(a[453]), .B(b[3]), .Z(n11838) );
  XOR U12891 ( .A(n11839), .B(n11838), .Z(n11841) );
  XOR U12892 ( .A(n11840), .B(n11841), .Z(n11829) );
  NANDN U12893 ( .A(n11818), .B(n11817), .Z(n11822) );
  OR U12894 ( .A(n11820), .B(n11819), .Z(n11821) );
  AND U12895 ( .A(n11822), .B(n11821), .Z(n11828) );
  XOR U12896 ( .A(n11829), .B(n11828), .Z(n11831) );
  XOR U12897 ( .A(n11830), .B(n11831), .Z(n11844) );
  XNOR U12898 ( .A(n11844), .B(sreg[1477]), .Z(n11846) );
  NANDN U12899 ( .A(n11823), .B(sreg[1476]), .Z(n11827) );
  NAND U12900 ( .A(n11825), .B(n11824), .Z(n11826) );
  NAND U12901 ( .A(n11827), .B(n11826), .Z(n11845) );
  XOR U12902 ( .A(n11846), .B(n11845), .Z(c[1477]) );
  NANDN U12903 ( .A(n11829), .B(n11828), .Z(n11833) );
  OR U12904 ( .A(n11831), .B(n11830), .Z(n11832) );
  AND U12905 ( .A(n11833), .B(n11832), .Z(n11851) );
  XOR U12906 ( .A(a[456]), .B(n2241), .Z(n11855) );
  AND U12907 ( .A(a[454]), .B(b[3]), .Z(n11859) );
  AND U12908 ( .A(a[458]), .B(b[0]), .Z(n11835) );
  XNOR U12909 ( .A(n11835), .B(n2175), .Z(n11837) );
  NANDN U12910 ( .A(b[0]), .B(a[457]), .Z(n11836) );
  NAND U12911 ( .A(n11837), .B(n11836), .Z(n11860) );
  XOR U12912 ( .A(n11859), .B(n11860), .Z(n11862) );
  XOR U12913 ( .A(n11861), .B(n11862), .Z(n11850) );
  NANDN U12914 ( .A(n11839), .B(n11838), .Z(n11843) );
  OR U12915 ( .A(n11841), .B(n11840), .Z(n11842) );
  AND U12916 ( .A(n11843), .B(n11842), .Z(n11849) );
  XOR U12917 ( .A(n11850), .B(n11849), .Z(n11852) );
  XOR U12918 ( .A(n11851), .B(n11852), .Z(n11865) );
  XNOR U12919 ( .A(n11865), .B(sreg[1478]), .Z(n11867) );
  NANDN U12920 ( .A(n11844), .B(sreg[1477]), .Z(n11848) );
  NAND U12921 ( .A(n11846), .B(n11845), .Z(n11847) );
  NAND U12922 ( .A(n11848), .B(n11847), .Z(n11866) );
  XOR U12923 ( .A(n11867), .B(n11866), .Z(c[1478]) );
  NANDN U12924 ( .A(n11850), .B(n11849), .Z(n11854) );
  OR U12925 ( .A(n11852), .B(n11851), .Z(n11853) );
  AND U12926 ( .A(n11854), .B(n11853), .Z(n11872) );
  XOR U12927 ( .A(a[457]), .B(n2241), .Z(n11876) );
  AND U12928 ( .A(a[459]), .B(b[0]), .Z(n11856) );
  XNOR U12929 ( .A(n11856), .B(n2175), .Z(n11858) );
  NANDN U12930 ( .A(b[0]), .B(a[458]), .Z(n11857) );
  NAND U12931 ( .A(n11858), .B(n11857), .Z(n11881) );
  AND U12932 ( .A(a[455]), .B(b[3]), .Z(n11880) );
  XOR U12933 ( .A(n11881), .B(n11880), .Z(n11883) );
  XOR U12934 ( .A(n11882), .B(n11883), .Z(n11871) );
  NANDN U12935 ( .A(n11860), .B(n11859), .Z(n11864) );
  OR U12936 ( .A(n11862), .B(n11861), .Z(n11863) );
  AND U12937 ( .A(n11864), .B(n11863), .Z(n11870) );
  XOR U12938 ( .A(n11871), .B(n11870), .Z(n11873) );
  XOR U12939 ( .A(n11872), .B(n11873), .Z(n11886) );
  XNOR U12940 ( .A(n11886), .B(sreg[1479]), .Z(n11888) );
  NANDN U12941 ( .A(n11865), .B(sreg[1478]), .Z(n11869) );
  NAND U12942 ( .A(n11867), .B(n11866), .Z(n11868) );
  NAND U12943 ( .A(n11869), .B(n11868), .Z(n11887) );
  XOR U12944 ( .A(n11888), .B(n11887), .Z(c[1479]) );
  NANDN U12945 ( .A(n11871), .B(n11870), .Z(n11875) );
  OR U12946 ( .A(n11873), .B(n11872), .Z(n11874) );
  AND U12947 ( .A(n11875), .B(n11874), .Z(n11893) );
  XOR U12948 ( .A(a[458]), .B(n2241), .Z(n11897) );
  AND U12949 ( .A(a[460]), .B(b[0]), .Z(n11877) );
  XNOR U12950 ( .A(n11877), .B(n2175), .Z(n11879) );
  NANDN U12951 ( .A(b[0]), .B(a[459]), .Z(n11878) );
  NAND U12952 ( .A(n11879), .B(n11878), .Z(n11902) );
  AND U12953 ( .A(a[456]), .B(b[3]), .Z(n11901) );
  XOR U12954 ( .A(n11902), .B(n11901), .Z(n11904) );
  XOR U12955 ( .A(n11903), .B(n11904), .Z(n11892) );
  NANDN U12956 ( .A(n11881), .B(n11880), .Z(n11885) );
  OR U12957 ( .A(n11883), .B(n11882), .Z(n11884) );
  AND U12958 ( .A(n11885), .B(n11884), .Z(n11891) );
  XOR U12959 ( .A(n11892), .B(n11891), .Z(n11894) );
  XOR U12960 ( .A(n11893), .B(n11894), .Z(n11907) );
  XNOR U12961 ( .A(n11907), .B(sreg[1480]), .Z(n11909) );
  NANDN U12962 ( .A(n11886), .B(sreg[1479]), .Z(n11890) );
  NAND U12963 ( .A(n11888), .B(n11887), .Z(n11889) );
  NAND U12964 ( .A(n11890), .B(n11889), .Z(n11908) );
  XOR U12965 ( .A(n11909), .B(n11908), .Z(c[1480]) );
  NANDN U12966 ( .A(n11892), .B(n11891), .Z(n11896) );
  OR U12967 ( .A(n11894), .B(n11893), .Z(n11895) );
  AND U12968 ( .A(n11896), .B(n11895), .Z(n11914) );
  XOR U12969 ( .A(a[459]), .B(n2241), .Z(n11918) );
  AND U12970 ( .A(a[457]), .B(b[3]), .Z(n11922) );
  AND U12971 ( .A(a[461]), .B(b[0]), .Z(n11898) );
  XNOR U12972 ( .A(n11898), .B(n2175), .Z(n11900) );
  NANDN U12973 ( .A(b[0]), .B(a[460]), .Z(n11899) );
  NAND U12974 ( .A(n11900), .B(n11899), .Z(n11923) );
  XOR U12975 ( .A(n11922), .B(n11923), .Z(n11925) );
  XOR U12976 ( .A(n11924), .B(n11925), .Z(n11913) );
  NANDN U12977 ( .A(n11902), .B(n11901), .Z(n11906) );
  OR U12978 ( .A(n11904), .B(n11903), .Z(n11905) );
  AND U12979 ( .A(n11906), .B(n11905), .Z(n11912) );
  XOR U12980 ( .A(n11913), .B(n11912), .Z(n11915) );
  XOR U12981 ( .A(n11914), .B(n11915), .Z(n11928) );
  XNOR U12982 ( .A(n11928), .B(sreg[1481]), .Z(n11930) );
  NANDN U12983 ( .A(n11907), .B(sreg[1480]), .Z(n11911) );
  NAND U12984 ( .A(n11909), .B(n11908), .Z(n11910) );
  NAND U12985 ( .A(n11911), .B(n11910), .Z(n11929) );
  XOR U12986 ( .A(n11930), .B(n11929), .Z(c[1481]) );
  NANDN U12987 ( .A(n11913), .B(n11912), .Z(n11917) );
  OR U12988 ( .A(n11915), .B(n11914), .Z(n11916) );
  AND U12989 ( .A(n11917), .B(n11916), .Z(n11935) );
  XOR U12990 ( .A(a[460]), .B(n2241), .Z(n11939) );
  AND U12991 ( .A(a[462]), .B(b[0]), .Z(n11919) );
  XNOR U12992 ( .A(n11919), .B(n2175), .Z(n11921) );
  NANDN U12993 ( .A(b[0]), .B(a[461]), .Z(n11920) );
  NAND U12994 ( .A(n11921), .B(n11920), .Z(n11944) );
  AND U12995 ( .A(a[458]), .B(b[3]), .Z(n11943) );
  XOR U12996 ( .A(n11944), .B(n11943), .Z(n11946) );
  XOR U12997 ( .A(n11945), .B(n11946), .Z(n11934) );
  NANDN U12998 ( .A(n11923), .B(n11922), .Z(n11927) );
  OR U12999 ( .A(n11925), .B(n11924), .Z(n11926) );
  AND U13000 ( .A(n11927), .B(n11926), .Z(n11933) );
  XOR U13001 ( .A(n11934), .B(n11933), .Z(n11936) );
  XOR U13002 ( .A(n11935), .B(n11936), .Z(n11949) );
  XNOR U13003 ( .A(n11949), .B(sreg[1482]), .Z(n11951) );
  NANDN U13004 ( .A(n11928), .B(sreg[1481]), .Z(n11932) );
  NAND U13005 ( .A(n11930), .B(n11929), .Z(n11931) );
  NAND U13006 ( .A(n11932), .B(n11931), .Z(n11950) );
  XOR U13007 ( .A(n11951), .B(n11950), .Z(c[1482]) );
  NANDN U13008 ( .A(n11934), .B(n11933), .Z(n11938) );
  OR U13009 ( .A(n11936), .B(n11935), .Z(n11937) );
  AND U13010 ( .A(n11938), .B(n11937), .Z(n11956) );
  XOR U13011 ( .A(a[461]), .B(n2242), .Z(n11960) );
  AND U13012 ( .A(a[463]), .B(b[0]), .Z(n11940) );
  XNOR U13013 ( .A(n11940), .B(n2175), .Z(n11942) );
  NANDN U13014 ( .A(b[0]), .B(a[462]), .Z(n11941) );
  NAND U13015 ( .A(n11942), .B(n11941), .Z(n11965) );
  AND U13016 ( .A(a[459]), .B(b[3]), .Z(n11964) );
  XOR U13017 ( .A(n11965), .B(n11964), .Z(n11967) );
  XOR U13018 ( .A(n11966), .B(n11967), .Z(n11955) );
  NANDN U13019 ( .A(n11944), .B(n11943), .Z(n11948) );
  OR U13020 ( .A(n11946), .B(n11945), .Z(n11947) );
  AND U13021 ( .A(n11948), .B(n11947), .Z(n11954) );
  XOR U13022 ( .A(n11955), .B(n11954), .Z(n11957) );
  XOR U13023 ( .A(n11956), .B(n11957), .Z(n11970) );
  XNOR U13024 ( .A(n11970), .B(sreg[1483]), .Z(n11972) );
  NANDN U13025 ( .A(n11949), .B(sreg[1482]), .Z(n11953) );
  NAND U13026 ( .A(n11951), .B(n11950), .Z(n11952) );
  NAND U13027 ( .A(n11953), .B(n11952), .Z(n11971) );
  XOR U13028 ( .A(n11972), .B(n11971), .Z(c[1483]) );
  NANDN U13029 ( .A(n11955), .B(n11954), .Z(n11959) );
  OR U13030 ( .A(n11957), .B(n11956), .Z(n11958) );
  AND U13031 ( .A(n11959), .B(n11958), .Z(n11977) );
  XOR U13032 ( .A(a[462]), .B(n2242), .Z(n11981) );
  AND U13033 ( .A(a[464]), .B(b[0]), .Z(n11961) );
  XNOR U13034 ( .A(n11961), .B(n2175), .Z(n11963) );
  NANDN U13035 ( .A(b[0]), .B(a[463]), .Z(n11962) );
  NAND U13036 ( .A(n11963), .B(n11962), .Z(n11986) );
  AND U13037 ( .A(a[460]), .B(b[3]), .Z(n11985) );
  XOR U13038 ( .A(n11986), .B(n11985), .Z(n11988) );
  XOR U13039 ( .A(n11987), .B(n11988), .Z(n11976) );
  NANDN U13040 ( .A(n11965), .B(n11964), .Z(n11969) );
  OR U13041 ( .A(n11967), .B(n11966), .Z(n11968) );
  AND U13042 ( .A(n11969), .B(n11968), .Z(n11975) );
  XOR U13043 ( .A(n11976), .B(n11975), .Z(n11978) );
  XOR U13044 ( .A(n11977), .B(n11978), .Z(n11991) );
  XNOR U13045 ( .A(n11991), .B(sreg[1484]), .Z(n11993) );
  NANDN U13046 ( .A(n11970), .B(sreg[1483]), .Z(n11974) );
  NAND U13047 ( .A(n11972), .B(n11971), .Z(n11973) );
  NAND U13048 ( .A(n11974), .B(n11973), .Z(n11992) );
  XOR U13049 ( .A(n11993), .B(n11992), .Z(c[1484]) );
  NANDN U13050 ( .A(n11976), .B(n11975), .Z(n11980) );
  OR U13051 ( .A(n11978), .B(n11977), .Z(n11979) );
  AND U13052 ( .A(n11980), .B(n11979), .Z(n11998) );
  XOR U13053 ( .A(a[463]), .B(n2242), .Z(n12002) );
  AND U13054 ( .A(a[465]), .B(b[0]), .Z(n11982) );
  XNOR U13055 ( .A(n11982), .B(n2175), .Z(n11984) );
  NANDN U13056 ( .A(b[0]), .B(a[464]), .Z(n11983) );
  NAND U13057 ( .A(n11984), .B(n11983), .Z(n12007) );
  AND U13058 ( .A(a[461]), .B(b[3]), .Z(n12006) );
  XOR U13059 ( .A(n12007), .B(n12006), .Z(n12009) );
  XOR U13060 ( .A(n12008), .B(n12009), .Z(n11997) );
  NANDN U13061 ( .A(n11986), .B(n11985), .Z(n11990) );
  OR U13062 ( .A(n11988), .B(n11987), .Z(n11989) );
  AND U13063 ( .A(n11990), .B(n11989), .Z(n11996) );
  XOR U13064 ( .A(n11997), .B(n11996), .Z(n11999) );
  XOR U13065 ( .A(n11998), .B(n11999), .Z(n12012) );
  XNOR U13066 ( .A(n12012), .B(sreg[1485]), .Z(n12014) );
  NANDN U13067 ( .A(n11991), .B(sreg[1484]), .Z(n11995) );
  NAND U13068 ( .A(n11993), .B(n11992), .Z(n11994) );
  NAND U13069 ( .A(n11995), .B(n11994), .Z(n12013) );
  XOR U13070 ( .A(n12014), .B(n12013), .Z(c[1485]) );
  NANDN U13071 ( .A(n11997), .B(n11996), .Z(n12001) );
  OR U13072 ( .A(n11999), .B(n11998), .Z(n12000) );
  AND U13073 ( .A(n12001), .B(n12000), .Z(n12019) );
  XOR U13074 ( .A(a[464]), .B(n2242), .Z(n12023) );
  AND U13075 ( .A(a[466]), .B(b[0]), .Z(n12003) );
  XNOR U13076 ( .A(n12003), .B(n2175), .Z(n12005) );
  NANDN U13077 ( .A(b[0]), .B(a[465]), .Z(n12004) );
  NAND U13078 ( .A(n12005), .B(n12004), .Z(n12028) );
  AND U13079 ( .A(a[462]), .B(b[3]), .Z(n12027) );
  XOR U13080 ( .A(n12028), .B(n12027), .Z(n12030) );
  XOR U13081 ( .A(n12029), .B(n12030), .Z(n12018) );
  NANDN U13082 ( .A(n12007), .B(n12006), .Z(n12011) );
  OR U13083 ( .A(n12009), .B(n12008), .Z(n12010) );
  AND U13084 ( .A(n12011), .B(n12010), .Z(n12017) );
  XOR U13085 ( .A(n12018), .B(n12017), .Z(n12020) );
  XOR U13086 ( .A(n12019), .B(n12020), .Z(n12033) );
  XNOR U13087 ( .A(n12033), .B(sreg[1486]), .Z(n12035) );
  NANDN U13088 ( .A(n12012), .B(sreg[1485]), .Z(n12016) );
  NAND U13089 ( .A(n12014), .B(n12013), .Z(n12015) );
  NAND U13090 ( .A(n12016), .B(n12015), .Z(n12034) );
  XOR U13091 ( .A(n12035), .B(n12034), .Z(c[1486]) );
  NANDN U13092 ( .A(n12018), .B(n12017), .Z(n12022) );
  OR U13093 ( .A(n12020), .B(n12019), .Z(n12021) );
  AND U13094 ( .A(n12022), .B(n12021), .Z(n12040) );
  XOR U13095 ( .A(a[465]), .B(n2242), .Z(n12044) );
  AND U13096 ( .A(a[467]), .B(b[0]), .Z(n12024) );
  XNOR U13097 ( .A(n12024), .B(n2175), .Z(n12026) );
  NANDN U13098 ( .A(b[0]), .B(a[466]), .Z(n12025) );
  NAND U13099 ( .A(n12026), .B(n12025), .Z(n12049) );
  AND U13100 ( .A(a[463]), .B(b[3]), .Z(n12048) );
  XOR U13101 ( .A(n12049), .B(n12048), .Z(n12051) );
  XOR U13102 ( .A(n12050), .B(n12051), .Z(n12039) );
  NANDN U13103 ( .A(n12028), .B(n12027), .Z(n12032) );
  OR U13104 ( .A(n12030), .B(n12029), .Z(n12031) );
  AND U13105 ( .A(n12032), .B(n12031), .Z(n12038) );
  XOR U13106 ( .A(n12039), .B(n12038), .Z(n12041) );
  XOR U13107 ( .A(n12040), .B(n12041), .Z(n12054) );
  XNOR U13108 ( .A(n12054), .B(sreg[1487]), .Z(n12056) );
  NANDN U13109 ( .A(n12033), .B(sreg[1486]), .Z(n12037) );
  NAND U13110 ( .A(n12035), .B(n12034), .Z(n12036) );
  NAND U13111 ( .A(n12037), .B(n12036), .Z(n12055) );
  XOR U13112 ( .A(n12056), .B(n12055), .Z(c[1487]) );
  NANDN U13113 ( .A(n12039), .B(n12038), .Z(n12043) );
  OR U13114 ( .A(n12041), .B(n12040), .Z(n12042) );
  AND U13115 ( .A(n12043), .B(n12042), .Z(n12061) );
  XOR U13116 ( .A(a[466]), .B(n2242), .Z(n12065) );
  AND U13117 ( .A(a[468]), .B(b[0]), .Z(n12045) );
  XNOR U13118 ( .A(n12045), .B(n2175), .Z(n12047) );
  NANDN U13119 ( .A(b[0]), .B(a[467]), .Z(n12046) );
  NAND U13120 ( .A(n12047), .B(n12046), .Z(n12070) );
  AND U13121 ( .A(a[464]), .B(b[3]), .Z(n12069) );
  XOR U13122 ( .A(n12070), .B(n12069), .Z(n12072) );
  XOR U13123 ( .A(n12071), .B(n12072), .Z(n12060) );
  NANDN U13124 ( .A(n12049), .B(n12048), .Z(n12053) );
  OR U13125 ( .A(n12051), .B(n12050), .Z(n12052) );
  AND U13126 ( .A(n12053), .B(n12052), .Z(n12059) );
  XOR U13127 ( .A(n12060), .B(n12059), .Z(n12062) );
  XOR U13128 ( .A(n12061), .B(n12062), .Z(n12075) );
  XNOR U13129 ( .A(n12075), .B(sreg[1488]), .Z(n12077) );
  NANDN U13130 ( .A(n12054), .B(sreg[1487]), .Z(n12058) );
  NAND U13131 ( .A(n12056), .B(n12055), .Z(n12057) );
  NAND U13132 ( .A(n12058), .B(n12057), .Z(n12076) );
  XOR U13133 ( .A(n12077), .B(n12076), .Z(c[1488]) );
  NANDN U13134 ( .A(n12060), .B(n12059), .Z(n12064) );
  OR U13135 ( .A(n12062), .B(n12061), .Z(n12063) );
  AND U13136 ( .A(n12064), .B(n12063), .Z(n12082) );
  XOR U13137 ( .A(a[467]), .B(n2242), .Z(n12086) );
  AND U13138 ( .A(a[469]), .B(b[0]), .Z(n12066) );
  XNOR U13139 ( .A(n12066), .B(n2175), .Z(n12068) );
  NANDN U13140 ( .A(b[0]), .B(a[468]), .Z(n12067) );
  NAND U13141 ( .A(n12068), .B(n12067), .Z(n12091) );
  AND U13142 ( .A(a[465]), .B(b[3]), .Z(n12090) );
  XOR U13143 ( .A(n12091), .B(n12090), .Z(n12093) );
  XOR U13144 ( .A(n12092), .B(n12093), .Z(n12081) );
  NANDN U13145 ( .A(n12070), .B(n12069), .Z(n12074) );
  OR U13146 ( .A(n12072), .B(n12071), .Z(n12073) );
  AND U13147 ( .A(n12074), .B(n12073), .Z(n12080) );
  XOR U13148 ( .A(n12081), .B(n12080), .Z(n12083) );
  XOR U13149 ( .A(n12082), .B(n12083), .Z(n12096) );
  XNOR U13150 ( .A(n12096), .B(sreg[1489]), .Z(n12098) );
  NANDN U13151 ( .A(n12075), .B(sreg[1488]), .Z(n12079) );
  NAND U13152 ( .A(n12077), .B(n12076), .Z(n12078) );
  NAND U13153 ( .A(n12079), .B(n12078), .Z(n12097) );
  XOR U13154 ( .A(n12098), .B(n12097), .Z(c[1489]) );
  NANDN U13155 ( .A(n12081), .B(n12080), .Z(n12085) );
  OR U13156 ( .A(n12083), .B(n12082), .Z(n12084) );
  AND U13157 ( .A(n12085), .B(n12084), .Z(n12103) );
  XOR U13158 ( .A(a[468]), .B(n2243), .Z(n12107) );
  AND U13159 ( .A(a[470]), .B(b[0]), .Z(n12087) );
  XNOR U13160 ( .A(n12087), .B(n2175), .Z(n12089) );
  NANDN U13161 ( .A(b[0]), .B(a[469]), .Z(n12088) );
  NAND U13162 ( .A(n12089), .B(n12088), .Z(n12112) );
  AND U13163 ( .A(a[466]), .B(b[3]), .Z(n12111) );
  XOR U13164 ( .A(n12112), .B(n12111), .Z(n12114) );
  XOR U13165 ( .A(n12113), .B(n12114), .Z(n12102) );
  NANDN U13166 ( .A(n12091), .B(n12090), .Z(n12095) );
  OR U13167 ( .A(n12093), .B(n12092), .Z(n12094) );
  AND U13168 ( .A(n12095), .B(n12094), .Z(n12101) );
  XOR U13169 ( .A(n12102), .B(n12101), .Z(n12104) );
  XOR U13170 ( .A(n12103), .B(n12104), .Z(n12117) );
  XNOR U13171 ( .A(n12117), .B(sreg[1490]), .Z(n12119) );
  NANDN U13172 ( .A(n12096), .B(sreg[1489]), .Z(n12100) );
  NAND U13173 ( .A(n12098), .B(n12097), .Z(n12099) );
  NAND U13174 ( .A(n12100), .B(n12099), .Z(n12118) );
  XOR U13175 ( .A(n12119), .B(n12118), .Z(c[1490]) );
  NANDN U13176 ( .A(n12102), .B(n12101), .Z(n12106) );
  OR U13177 ( .A(n12104), .B(n12103), .Z(n12105) );
  AND U13178 ( .A(n12106), .B(n12105), .Z(n12124) );
  XOR U13179 ( .A(a[469]), .B(n2243), .Z(n12128) );
  AND U13180 ( .A(a[471]), .B(b[0]), .Z(n12108) );
  XNOR U13181 ( .A(n12108), .B(n2175), .Z(n12110) );
  NANDN U13182 ( .A(b[0]), .B(a[470]), .Z(n12109) );
  NAND U13183 ( .A(n12110), .B(n12109), .Z(n12133) );
  AND U13184 ( .A(a[467]), .B(b[3]), .Z(n12132) );
  XOR U13185 ( .A(n12133), .B(n12132), .Z(n12135) );
  XOR U13186 ( .A(n12134), .B(n12135), .Z(n12123) );
  NANDN U13187 ( .A(n12112), .B(n12111), .Z(n12116) );
  OR U13188 ( .A(n12114), .B(n12113), .Z(n12115) );
  AND U13189 ( .A(n12116), .B(n12115), .Z(n12122) );
  XOR U13190 ( .A(n12123), .B(n12122), .Z(n12125) );
  XOR U13191 ( .A(n12124), .B(n12125), .Z(n12138) );
  XNOR U13192 ( .A(n12138), .B(sreg[1491]), .Z(n12140) );
  NANDN U13193 ( .A(n12117), .B(sreg[1490]), .Z(n12121) );
  NAND U13194 ( .A(n12119), .B(n12118), .Z(n12120) );
  NAND U13195 ( .A(n12121), .B(n12120), .Z(n12139) );
  XOR U13196 ( .A(n12140), .B(n12139), .Z(c[1491]) );
  NANDN U13197 ( .A(n12123), .B(n12122), .Z(n12127) );
  OR U13198 ( .A(n12125), .B(n12124), .Z(n12126) );
  AND U13199 ( .A(n12127), .B(n12126), .Z(n12145) );
  XOR U13200 ( .A(a[470]), .B(n2243), .Z(n12149) );
  AND U13201 ( .A(a[468]), .B(b[3]), .Z(n12153) );
  AND U13202 ( .A(a[472]), .B(b[0]), .Z(n12129) );
  XNOR U13203 ( .A(n12129), .B(n2175), .Z(n12131) );
  NANDN U13204 ( .A(b[0]), .B(a[471]), .Z(n12130) );
  NAND U13205 ( .A(n12131), .B(n12130), .Z(n12154) );
  XOR U13206 ( .A(n12153), .B(n12154), .Z(n12156) );
  XOR U13207 ( .A(n12155), .B(n12156), .Z(n12144) );
  NANDN U13208 ( .A(n12133), .B(n12132), .Z(n12137) );
  OR U13209 ( .A(n12135), .B(n12134), .Z(n12136) );
  AND U13210 ( .A(n12137), .B(n12136), .Z(n12143) );
  XOR U13211 ( .A(n12144), .B(n12143), .Z(n12146) );
  XOR U13212 ( .A(n12145), .B(n12146), .Z(n12159) );
  XNOR U13213 ( .A(n12159), .B(sreg[1492]), .Z(n12161) );
  NANDN U13214 ( .A(n12138), .B(sreg[1491]), .Z(n12142) );
  NAND U13215 ( .A(n12140), .B(n12139), .Z(n12141) );
  NAND U13216 ( .A(n12142), .B(n12141), .Z(n12160) );
  XOR U13217 ( .A(n12161), .B(n12160), .Z(c[1492]) );
  NANDN U13218 ( .A(n12144), .B(n12143), .Z(n12148) );
  OR U13219 ( .A(n12146), .B(n12145), .Z(n12147) );
  AND U13220 ( .A(n12148), .B(n12147), .Z(n12166) );
  XOR U13221 ( .A(a[471]), .B(n2243), .Z(n12170) );
  AND U13222 ( .A(a[473]), .B(b[0]), .Z(n12150) );
  XNOR U13223 ( .A(n12150), .B(n2175), .Z(n12152) );
  NANDN U13224 ( .A(b[0]), .B(a[472]), .Z(n12151) );
  NAND U13225 ( .A(n12152), .B(n12151), .Z(n12175) );
  AND U13226 ( .A(a[469]), .B(b[3]), .Z(n12174) );
  XOR U13227 ( .A(n12175), .B(n12174), .Z(n12177) );
  XOR U13228 ( .A(n12176), .B(n12177), .Z(n12165) );
  NANDN U13229 ( .A(n12154), .B(n12153), .Z(n12158) );
  OR U13230 ( .A(n12156), .B(n12155), .Z(n12157) );
  AND U13231 ( .A(n12158), .B(n12157), .Z(n12164) );
  XOR U13232 ( .A(n12165), .B(n12164), .Z(n12167) );
  XOR U13233 ( .A(n12166), .B(n12167), .Z(n12180) );
  XNOR U13234 ( .A(n12180), .B(sreg[1493]), .Z(n12182) );
  NANDN U13235 ( .A(n12159), .B(sreg[1492]), .Z(n12163) );
  NAND U13236 ( .A(n12161), .B(n12160), .Z(n12162) );
  NAND U13237 ( .A(n12163), .B(n12162), .Z(n12181) );
  XOR U13238 ( .A(n12182), .B(n12181), .Z(c[1493]) );
  NANDN U13239 ( .A(n12165), .B(n12164), .Z(n12169) );
  OR U13240 ( .A(n12167), .B(n12166), .Z(n12168) );
  AND U13241 ( .A(n12169), .B(n12168), .Z(n12187) );
  XOR U13242 ( .A(a[472]), .B(n2243), .Z(n12191) );
  AND U13243 ( .A(a[474]), .B(b[0]), .Z(n12171) );
  XNOR U13244 ( .A(n12171), .B(n2175), .Z(n12173) );
  NANDN U13245 ( .A(b[0]), .B(a[473]), .Z(n12172) );
  NAND U13246 ( .A(n12173), .B(n12172), .Z(n12196) );
  AND U13247 ( .A(a[470]), .B(b[3]), .Z(n12195) );
  XOR U13248 ( .A(n12196), .B(n12195), .Z(n12198) );
  XOR U13249 ( .A(n12197), .B(n12198), .Z(n12186) );
  NANDN U13250 ( .A(n12175), .B(n12174), .Z(n12179) );
  OR U13251 ( .A(n12177), .B(n12176), .Z(n12178) );
  AND U13252 ( .A(n12179), .B(n12178), .Z(n12185) );
  XOR U13253 ( .A(n12186), .B(n12185), .Z(n12188) );
  XOR U13254 ( .A(n12187), .B(n12188), .Z(n12201) );
  XNOR U13255 ( .A(n12201), .B(sreg[1494]), .Z(n12203) );
  NANDN U13256 ( .A(n12180), .B(sreg[1493]), .Z(n12184) );
  NAND U13257 ( .A(n12182), .B(n12181), .Z(n12183) );
  NAND U13258 ( .A(n12184), .B(n12183), .Z(n12202) );
  XOR U13259 ( .A(n12203), .B(n12202), .Z(c[1494]) );
  NANDN U13260 ( .A(n12186), .B(n12185), .Z(n12190) );
  OR U13261 ( .A(n12188), .B(n12187), .Z(n12189) );
  AND U13262 ( .A(n12190), .B(n12189), .Z(n12208) );
  XOR U13263 ( .A(a[473]), .B(n2243), .Z(n12212) );
  AND U13264 ( .A(a[475]), .B(b[0]), .Z(n12192) );
  XNOR U13265 ( .A(n12192), .B(n2175), .Z(n12194) );
  NANDN U13266 ( .A(b[0]), .B(a[474]), .Z(n12193) );
  NAND U13267 ( .A(n12194), .B(n12193), .Z(n12217) );
  AND U13268 ( .A(a[471]), .B(b[3]), .Z(n12216) );
  XOR U13269 ( .A(n12217), .B(n12216), .Z(n12219) );
  XOR U13270 ( .A(n12218), .B(n12219), .Z(n12207) );
  NANDN U13271 ( .A(n12196), .B(n12195), .Z(n12200) );
  OR U13272 ( .A(n12198), .B(n12197), .Z(n12199) );
  AND U13273 ( .A(n12200), .B(n12199), .Z(n12206) );
  XOR U13274 ( .A(n12207), .B(n12206), .Z(n12209) );
  XOR U13275 ( .A(n12208), .B(n12209), .Z(n12222) );
  XNOR U13276 ( .A(n12222), .B(sreg[1495]), .Z(n12224) );
  NANDN U13277 ( .A(n12201), .B(sreg[1494]), .Z(n12205) );
  NAND U13278 ( .A(n12203), .B(n12202), .Z(n12204) );
  NAND U13279 ( .A(n12205), .B(n12204), .Z(n12223) );
  XOR U13280 ( .A(n12224), .B(n12223), .Z(c[1495]) );
  NANDN U13281 ( .A(n12207), .B(n12206), .Z(n12211) );
  OR U13282 ( .A(n12209), .B(n12208), .Z(n12210) );
  AND U13283 ( .A(n12211), .B(n12210), .Z(n12229) );
  XOR U13284 ( .A(a[474]), .B(n2243), .Z(n12233) );
  AND U13285 ( .A(a[472]), .B(b[3]), .Z(n12237) );
  AND U13286 ( .A(a[476]), .B(b[0]), .Z(n12213) );
  XNOR U13287 ( .A(n12213), .B(n2175), .Z(n12215) );
  NANDN U13288 ( .A(b[0]), .B(a[475]), .Z(n12214) );
  NAND U13289 ( .A(n12215), .B(n12214), .Z(n12238) );
  XOR U13290 ( .A(n12237), .B(n12238), .Z(n12240) );
  XOR U13291 ( .A(n12239), .B(n12240), .Z(n12228) );
  NANDN U13292 ( .A(n12217), .B(n12216), .Z(n12221) );
  OR U13293 ( .A(n12219), .B(n12218), .Z(n12220) );
  AND U13294 ( .A(n12221), .B(n12220), .Z(n12227) );
  XOR U13295 ( .A(n12228), .B(n12227), .Z(n12230) );
  XOR U13296 ( .A(n12229), .B(n12230), .Z(n12243) );
  XNOR U13297 ( .A(n12243), .B(sreg[1496]), .Z(n12245) );
  NANDN U13298 ( .A(n12222), .B(sreg[1495]), .Z(n12226) );
  NAND U13299 ( .A(n12224), .B(n12223), .Z(n12225) );
  NAND U13300 ( .A(n12226), .B(n12225), .Z(n12244) );
  XOR U13301 ( .A(n12245), .B(n12244), .Z(c[1496]) );
  NANDN U13302 ( .A(n12228), .B(n12227), .Z(n12232) );
  OR U13303 ( .A(n12230), .B(n12229), .Z(n12231) );
  AND U13304 ( .A(n12232), .B(n12231), .Z(n12250) );
  XOR U13305 ( .A(a[475]), .B(n2244), .Z(n12254) );
  AND U13306 ( .A(a[477]), .B(b[0]), .Z(n12234) );
  XNOR U13307 ( .A(n12234), .B(n2175), .Z(n12236) );
  NANDN U13308 ( .A(b[0]), .B(a[476]), .Z(n12235) );
  NAND U13309 ( .A(n12236), .B(n12235), .Z(n12259) );
  AND U13310 ( .A(a[473]), .B(b[3]), .Z(n12258) );
  XOR U13311 ( .A(n12259), .B(n12258), .Z(n12261) );
  XOR U13312 ( .A(n12260), .B(n12261), .Z(n12249) );
  NANDN U13313 ( .A(n12238), .B(n12237), .Z(n12242) );
  OR U13314 ( .A(n12240), .B(n12239), .Z(n12241) );
  AND U13315 ( .A(n12242), .B(n12241), .Z(n12248) );
  XOR U13316 ( .A(n12249), .B(n12248), .Z(n12251) );
  XOR U13317 ( .A(n12250), .B(n12251), .Z(n12264) );
  XNOR U13318 ( .A(n12264), .B(sreg[1497]), .Z(n12266) );
  NANDN U13319 ( .A(n12243), .B(sreg[1496]), .Z(n12247) );
  NAND U13320 ( .A(n12245), .B(n12244), .Z(n12246) );
  NAND U13321 ( .A(n12247), .B(n12246), .Z(n12265) );
  XOR U13322 ( .A(n12266), .B(n12265), .Z(c[1497]) );
  NANDN U13323 ( .A(n12249), .B(n12248), .Z(n12253) );
  OR U13324 ( .A(n12251), .B(n12250), .Z(n12252) );
  AND U13325 ( .A(n12253), .B(n12252), .Z(n12271) );
  XOR U13326 ( .A(a[476]), .B(n2244), .Z(n12275) );
  AND U13327 ( .A(a[478]), .B(b[0]), .Z(n12255) );
  XNOR U13328 ( .A(n12255), .B(n2175), .Z(n12257) );
  NANDN U13329 ( .A(b[0]), .B(a[477]), .Z(n12256) );
  NAND U13330 ( .A(n12257), .B(n12256), .Z(n12280) );
  AND U13331 ( .A(a[474]), .B(b[3]), .Z(n12279) );
  XOR U13332 ( .A(n12280), .B(n12279), .Z(n12282) );
  XOR U13333 ( .A(n12281), .B(n12282), .Z(n12270) );
  NANDN U13334 ( .A(n12259), .B(n12258), .Z(n12263) );
  OR U13335 ( .A(n12261), .B(n12260), .Z(n12262) );
  AND U13336 ( .A(n12263), .B(n12262), .Z(n12269) );
  XOR U13337 ( .A(n12270), .B(n12269), .Z(n12272) );
  XOR U13338 ( .A(n12271), .B(n12272), .Z(n12285) );
  XNOR U13339 ( .A(n12285), .B(sreg[1498]), .Z(n12287) );
  NANDN U13340 ( .A(n12264), .B(sreg[1497]), .Z(n12268) );
  NAND U13341 ( .A(n12266), .B(n12265), .Z(n12267) );
  NAND U13342 ( .A(n12268), .B(n12267), .Z(n12286) );
  XOR U13343 ( .A(n12287), .B(n12286), .Z(c[1498]) );
  NANDN U13344 ( .A(n12270), .B(n12269), .Z(n12274) );
  OR U13345 ( .A(n12272), .B(n12271), .Z(n12273) );
  AND U13346 ( .A(n12274), .B(n12273), .Z(n12292) );
  XOR U13347 ( .A(a[477]), .B(n2244), .Z(n12296) );
  AND U13348 ( .A(a[475]), .B(b[3]), .Z(n12300) );
  AND U13349 ( .A(a[479]), .B(b[0]), .Z(n12276) );
  XNOR U13350 ( .A(n12276), .B(n2175), .Z(n12278) );
  NANDN U13351 ( .A(b[0]), .B(a[478]), .Z(n12277) );
  NAND U13352 ( .A(n12278), .B(n12277), .Z(n12301) );
  XOR U13353 ( .A(n12300), .B(n12301), .Z(n12303) );
  XOR U13354 ( .A(n12302), .B(n12303), .Z(n12291) );
  NANDN U13355 ( .A(n12280), .B(n12279), .Z(n12284) );
  OR U13356 ( .A(n12282), .B(n12281), .Z(n12283) );
  AND U13357 ( .A(n12284), .B(n12283), .Z(n12290) );
  XOR U13358 ( .A(n12291), .B(n12290), .Z(n12293) );
  XOR U13359 ( .A(n12292), .B(n12293), .Z(n12306) );
  XNOR U13360 ( .A(n12306), .B(sreg[1499]), .Z(n12308) );
  NANDN U13361 ( .A(n12285), .B(sreg[1498]), .Z(n12289) );
  NAND U13362 ( .A(n12287), .B(n12286), .Z(n12288) );
  NAND U13363 ( .A(n12289), .B(n12288), .Z(n12307) );
  XOR U13364 ( .A(n12308), .B(n12307), .Z(c[1499]) );
  NANDN U13365 ( .A(n12291), .B(n12290), .Z(n12295) );
  OR U13366 ( .A(n12293), .B(n12292), .Z(n12294) );
  AND U13367 ( .A(n12295), .B(n12294), .Z(n12313) );
  XOR U13368 ( .A(a[478]), .B(n2244), .Z(n12317) );
  AND U13369 ( .A(a[476]), .B(b[3]), .Z(n12321) );
  AND U13370 ( .A(a[480]), .B(b[0]), .Z(n12297) );
  XNOR U13371 ( .A(n12297), .B(n2175), .Z(n12299) );
  NANDN U13372 ( .A(b[0]), .B(a[479]), .Z(n12298) );
  NAND U13373 ( .A(n12299), .B(n12298), .Z(n12322) );
  XOR U13374 ( .A(n12321), .B(n12322), .Z(n12324) );
  XOR U13375 ( .A(n12323), .B(n12324), .Z(n12312) );
  NANDN U13376 ( .A(n12301), .B(n12300), .Z(n12305) );
  OR U13377 ( .A(n12303), .B(n12302), .Z(n12304) );
  AND U13378 ( .A(n12305), .B(n12304), .Z(n12311) );
  XOR U13379 ( .A(n12312), .B(n12311), .Z(n12314) );
  XOR U13380 ( .A(n12313), .B(n12314), .Z(n12327) );
  XNOR U13381 ( .A(n12327), .B(sreg[1500]), .Z(n12329) );
  NANDN U13382 ( .A(n12306), .B(sreg[1499]), .Z(n12310) );
  NAND U13383 ( .A(n12308), .B(n12307), .Z(n12309) );
  NAND U13384 ( .A(n12310), .B(n12309), .Z(n12328) );
  XOR U13385 ( .A(n12329), .B(n12328), .Z(c[1500]) );
  NANDN U13386 ( .A(n12312), .B(n12311), .Z(n12316) );
  OR U13387 ( .A(n12314), .B(n12313), .Z(n12315) );
  AND U13388 ( .A(n12316), .B(n12315), .Z(n12334) );
  XOR U13389 ( .A(a[479]), .B(n2244), .Z(n12338) );
  AND U13390 ( .A(a[481]), .B(b[0]), .Z(n12318) );
  XNOR U13391 ( .A(n12318), .B(n2175), .Z(n12320) );
  NANDN U13392 ( .A(b[0]), .B(a[480]), .Z(n12319) );
  NAND U13393 ( .A(n12320), .B(n12319), .Z(n12343) );
  AND U13394 ( .A(a[477]), .B(b[3]), .Z(n12342) );
  XOR U13395 ( .A(n12343), .B(n12342), .Z(n12345) );
  XOR U13396 ( .A(n12344), .B(n12345), .Z(n12333) );
  NANDN U13397 ( .A(n12322), .B(n12321), .Z(n12326) );
  OR U13398 ( .A(n12324), .B(n12323), .Z(n12325) );
  AND U13399 ( .A(n12326), .B(n12325), .Z(n12332) );
  XOR U13400 ( .A(n12333), .B(n12332), .Z(n12335) );
  XOR U13401 ( .A(n12334), .B(n12335), .Z(n12348) );
  XNOR U13402 ( .A(n12348), .B(sreg[1501]), .Z(n12350) );
  NANDN U13403 ( .A(n12327), .B(sreg[1500]), .Z(n12331) );
  NAND U13404 ( .A(n12329), .B(n12328), .Z(n12330) );
  NAND U13405 ( .A(n12331), .B(n12330), .Z(n12349) );
  XOR U13406 ( .A(n12350), .B(n12349), .Z(c[1501]) );
  NANDN U13407 ( .A(n12333), .B(n12332), .Z(n12337) );
  OR U13408 ( .A(n12335), .B(n12334), .Z(n12336) );
  AND U13409 ( .A(n12337), .B(n12336), .Z(n12355) );
  XOR U13410 ( .A(a[480]), .B(n2244), .Z(n12359) );
  AND U13411 ( .A(a[478]), .B(b[3]), .Z(n12363) );
  AND U13412 ( .A(a[482]), .B(b[0]), .Z(n12339) );
  XNOR U13413 ( .A(n12339), .B(n2175), .Z(n12341) );
  NANDN U13414 ( .A(b[0]), .B(a[481]), .Z(n12340) );
  NAND U13415 ( .A(n12341), .B(n12340), .Z(n12364) );
  XOR U13416 ( .A(n12363), .B(n12364), .Z(n12366) );
  XOR U13417 ( .A(n12365), .B(n12366), .Z(n12354) );
  NANDN U13418 ( .A(n12343), .B(n12342), .Z(n12347) );
  OR U13419 ( .A(n12345), .B(n12344), .Z(n12346) );
  AND U13420 ( .A(n12347), .B(n12346), .Z(n12353) );
  XOR U13421 ( .A(n12354), .B(n12353), .Z(n12356) );
  XOR U13422 ( .A(n12355), .B(n12356), .Z(n12369) );
  XNOR U13423 ( .A(n12369), .B(sreg[1502]), .Z(n12371) );
  NANDN U13424 ( .A(n12348), .B(sreg[1501]), .Z(n12352) );
  NAND U13425 ( .A(n12350), .B(n12349), .Z(n12351) );
  NAND U13426 ( .A(n12352), .B(n12351), .Z(n12370) );
  XOR U13427 ( .A(n12371), .B(n12370), .Z(c[1502]) );
  NANDN U13428 ( .A(n12354), .B(n12353), .Z(n12358) );
  OR U13429 ( .A(n12356), .B(n12355), .Z(n12357) );
  AND U13430 ( .A(n12358), .B(n12357), .Z(n12376) );
  XOR U13431 ( .A(a[481]), .B(n2244), .Z(n12380) );
  AND U13432 ( .A(a[483]), .B(b[0]), .Z(n12360) );
  XNOR U13433 ( .A(n12360), .B(n2175), .Z(n12362) );
  NANDN U13434 ( .A(b[0]), .B(a[482]), .Z(n12361) );
  NAND U13435 ( .A(n12362), .B(n12361), .Z(n12385) );
  AND U13436 ( .A(a[479]), .B(b[3]), .Z(n12384) );
  XOR U13437 ( .A(n12385), .B(n12384), .Z(n12387) );
  XOR U13438 ( .A(n12386), .B(n12387), .Z(n12375) );
  NANDN U13439 ( .A(n12364), .B(n12363), .Z(n12368) );
  OR U13440 ( .A(n12366), .B(n12365), .Z(n12367) );
  AND U13441 ( .A(n12368), .B(n12367), .Z(n12374) );
  XOR U13442 ( .A(n12375), .B(n12374), .Z(n12377) );
  XOR U13443 ( .A(n12376), .B(n12377), .Z(n12390) );
  XNOR U13444 ( .A(n12390), .B(sreg[1503]), .Z(n12392) );
  NANDN U13445 ( .A(n12369), .B(sreg[1502]), .Z(n12373) );
  NAND U13446 ( .A(n12371), .B(n12370), .Z(n12372) );
  NAND U13447 ( .A(n12373), .B(n12372), .Z(n12391) );
  XOR U13448 ( .A(n12392), .B(n12391), .Z(c[1503]) );
  NANDN U13449 ( .A(n12375), .B(n12374), .Z(n12379) );
  OR U13450 ( .A(n12377), .B(n12376), .Z(n12378) );
  AND U13451 ( .A(n12379), .B(n12378), .Z(n12397) );
  XOR U13452 ( .A(a[482]), .B(n2245), .Z(n12401) );
  AND U13453 ( .A(a[480]), .B(b[3]), .Z(n12405) );
  AND U13454 ( .A(a[484]), .B(b[0]), .Z(n12381) );
  XNOR U13455 ( .A(n12381), .B(n2175), .Z(n12383) );
  NANDN U13456 ( .A(b[0]), .B(a[483]), .Z(n12382) );
  NAND U13457 ( .A(n12383), .B(n12382), .Z(n12406) );
  XOR U13458 ( .A(n12405), .B(n12406), .Z(n12408) );
  XOR U13459 ( .A(n12407), .B(n12408), .Z(n12396) );
  NANDN U13460 ( .A(n12385), .B(n12384), .Z(n12389) );
  OR U13461 ( .A(n12387), .B(n12386), .Z(n12388) );
  AND U13462 ( .A(n12389), .B(n12388), .Z(n12395) );
  XOR U13463 ( .A(n12396), .B(n12395), .Z(n12398) );
  XOR U13464 ( .A(n12397), .B(n12398), .Z(n12411) );
  XNOR U13465 ( .A(n12411), .B(sreg[1504]), .Z(n12413) );
  NANDN U13466 ( .A(n12390), .B(sreg[1503]), .Z(n12394) );
  NAND U13467 ( .A(n12392), .B(n12391), .Z(n12393) );
  NAND U13468 ( .A(n12394), .B(n12393), .Z(n12412) );
  XOR U13469 ( .A(n12413), .B(n12412), .Z(c[1504]) );
  NANDN U13470 ( .A(n12396), .B(n12395), .Z(n12400) );
  OR U13471 ( .A(n12398), .B(n12397), .Z(n12399) );
  AND U13472 ( .A(n12400), .B(n12399), .Z(n12418) );
  XOR U13473 ( .A(a[483]), .B(n2245), .Z(n12422) );
  AND U13474 ( .A(a[481]), .B(b[3]), .Z(n12426) );
  AND U13475 ( .A(a[485]), .B(b[0]), .Z(n12402) );
  XNOR U13476 ( .A(n12402), .B(n2175), .Z(n12404) );
  NANDN U13477 ( .A(b[0]), .B(a[484]), .Z(n12403) );
  NAND U13478 ( .A(n12404), .B(n12403), .Z(n12427) );
  XOR U13479 ( .A(n12426), .B(n12427), .Z(n12429) );
  XOR U13480 ( .A(n12428), .B(n12429), .Z(n12417) );
  NANDN U13481 ( .A(n12406), .B(n12405), .Z(n12410) );
  OR U13482 ( .A(n12408), .B(n12407), .Z(n12409) );
  AND U13483 ( .A(n12410), .B(n12409), .Z(n12416) );
  XOR U13484 ( .A(n12417), .B(n12416), .Z(n12419) );
  XOR U13485 ( .A(n12418), .B(n12419), .Z(n12432) );
  XNOR U13486 ( .A(n12432), .B(sreg[1505]), .Z(n12434) );
  NANDN U13487 ( .A(n12411), .B(sreg[1504]), .Z(n12415) );
  NAND U13488 ( .A(n12413), .B(n12412), .Z(n12414) );
  NAND U13489 ( .A(n12415), .B(n12414), .Z(n12433) );
  XOR U13490 ( .A(n12434), .B(n12433), .Z(c[1505]) );
  NANDN U13491 ( .A(n12417), .B(n12416), .Z(n12421) );
  OR U13492 ( .A(n12419), .B(n12418), .Z(n12420) );
  AND U13493 ( .A(n12421), .B(n12420), .Z(n12439) );
  XOR U13494 ( .A(a[484]), .B(n2245), .Z(n12443) );
  AND U13495 ( .A(a[486]), .B(b[0]), .Z(n12423) );
  XNOR U13496 ( .A(n12423), .B(n2175), .Z(n12425) );
  NANDN U13497 ( .A(b[0]), .B(a[485]), .Z(n12424) );
  NAND U13498 ( .A(n12425), .B(n12424), .Z(n12448) );
  AND U13499 ( .A(a[482]), .B(b[3]), .Z(n12447) );
  XOR U13500 ( .A(n12448), .B(n12447), .Z(n12450) );
  XOR U13501 ( .A(n12449), .B(n12450), .Z(n12438) );
  NANDN U13502 ( .A(n12427), .B(n12426), .Z(n12431) );
  OR U13503 ( .A(n12429), .B(n12428), .Z(n12430) );
  AND U13504 ( .A(n12431), .B(n12430), .Z(n12437) );
  XOR U13505 ( .A(n12438), .B(n12437), .Z(n12440) );
  XOR U13506 ( .A(n12439), .B(n12440), .Z(n12453) );
  XNOR U13507 ( .A(n12453), .B(sreg[1506]), .Z(n12455) );
  NANDN U13508 ( .A(n12432), .B(sreg[1505]), .Z(n12436) );
  NAND U13509 ( .A(n12434), .B(n12433), .Z(n12435) );
  NAND U13510 ( .A(n12436), .B(n12435), .Z(n12454) );
  XOR U13511 ( .A(n12455), .B(n12454), .Z(c[1506]) );
  NANDN U13512 ( .A(n12438), .B(n12437), .Z(n12442) );
  OR U13513 ( .A(n12440), .B(n12439), .Z(n12441) );
  AND U13514 ( .A(n12442), .B(n12441), .Z(n12460) );
  XOR U13515 ( .A(a[485]), .B(n2245), .Z(n12464) );
  AND U13516 ( .A(a[487]), .B(b[0]), .Z(n12444) );
  XNOR U13517 ( .A(n12444), .B(n2175), .Z(n12446) );
  NANDN U13518 ( .A(b[0]), .B(a[486]), .Z(n12445) );
  NAND U13519 ( .A(n12446), .B(n12445), .Z(n12469) );
  AND U13520 ( .A(a[483]), .B(b[3]), .Z(n12468) );
  XOR U13521 ( .A(n12469), .B(n12468), .Z(n12471) );
  XOR U13522 ( .A(n12470), .B(n12471), .Z(n12459) );
  NANDN U13523 ( .A(n12448), .B(n12447), .Z(n12452) );
  OR U13524 ( .A(n12450), .B(n12449), .Z(n12451) );
  AND U13525 ( .A(n12452), .B(n12451), .Z(n12458) );
  XOR U13526 ( .A(n12459), .B(n12458), .Z(n12461) );
  XOR U13527 ( .A(n12460), .B(n12461), .Z(n12474) );
  XNOR U13528 ( .A(n12474), .B(sreg[1507]), .Z(n12476) );
  NANDN U13529 ( .A(n12453), .B(sreg[1506]), .Z(n12457) );
  NAND U13530 ( .A(n12455), .B(n12454), .Z(n12456) );
  NAND U13531 ( .A(n12457), .B(n12456), .Z(n12475) );
  XOR U13532 ( .A(n12476), .B(n12475), .Z(c[1507]) );
  NANDN U13533 ( .A(n12459), .B(n12458), .Z(n12463) );
  OR U13534 ( .A(n12461), .B(n12460), .Z(n12462) );
  AND U13535 ( .A(n12463), .B(n12462), .Z(n12481) );
  XOR U13536 ( .A(a[486]), .B(n2245), .Z(n12485) );
  AND U13537 ( .A(a[488]), .B(b[0]), .Z(n12465) );
  XNOR U13538 ( .A(n12465), .B(n2175), .Z(n12467) );
  NANDN U13539 ( .A(b[0]), .B(a[487]), .Z(n12466) );
  NAND U13540 ( .A(n12467), .B(n12466), .Z(n12490) );
  AND U13541 ( .A(a[484]), .B(b[3]), .Z(n12489) );
  XOR U13542 ( .A(n12490), .B(n12489), .Z(n12492) );
  XOR U13543 ( .A(n12491), .B(n12492), .Z(n12480) );
  NANDN U13544 ( .A(n12469), .B(n12468), .Z(n12473) );
  OR U13545 ( .A(n12471), .B(n12470), .Z(n12472) );
  AND U13546 ( .A(n12473), .B(n12472), .Z(n12479) );
  XOR U13547 ( .A(n12480), .B(n12479), .Z(n12482) );
  XOR U13548 ( .A(n12481), .B(n12482), .Z(n12495) );
  XNOR U13549 ( .A(n12495), .B(sreg[1508]), .Z(n12497) );
  NANDN U13550 ( .A(n12474), .B(sreg[1507]), .Z(n12478) );
  NAND U13551 ( .A(n12476), .B(n12475), .Z(n12477) );
  NAND U13552 ( .A(n12478), .B(n12477), .Z(n12496) );
  XOR U13553 ( .A(n12497), .B(n12496), .Z(c[1508]) );
  NANDN U13554 ( .A(n12480), .B(n12479), .Z(n12484) );
  OR U13555 ( .A(n12482), .B(n12481), .Z(n12483) );
  AND U13556 ( .A(n12484), .B(n12483), .Z(n12502) );
  XOR U13557 ( .A(a[487]), .B(n2245), .Z(n12506) );
  AND U13558 ( .A(a[489]), .B(b[0]), .Z(n12486) );
  XNOR U13559 ( .A(n12486), .B(n2175), .Z(n12488) );
  NANDN U13560 ( .A(b[0]), .B(a[488]), .Z(n12487) );
  NAND U13561 ( .A(n12488), .B(n12487), .Z(n12511) );
  AND U13562 ( .A(a[485]), .B(b[3]), .Z(n12510) );
  XOR U13563 ( .A(n12511), .B(n12510), .Z(n12513) );
  XOR U13564 ( .A(n12512), .B(n12513), .Z(n12501) );
  NANDN U13565 ( .A(n12490), .B(n12489), .Z(n12494) );
  OR U13566 ( .A(n12492), .B(n12491), .Z(n12493) );
  AND U13567 ( .A(n12494), .B(n12493), .Z(n12500) );
  XOR U13568 ( .A(n12501), .B(n12500), .Z(n12503) );
  XOR U13569 ( .A(n12502), .B(n12503), .Z(n12516) );
  XNOR U13570 ( .A(n12516), .B(sreg[1509]), .Z(n12518) );
  NANDN U13571 ( .A(n12495), .B(sreg[1508]), .Z(n12499) );
  NAND U13572 ( .A(n12497), .B(n12496), .Z(n12498) );
  NAND U13573 ( .A(n12499), .B(n12498), .Z(n12517) );
  XOR U13574 ( .A(n12518), .B(n12517), .Z(c[1509]) );
  NANDN U13575 ( .A(n12501), .B(n12500), .Z(n12505) );
  OR U13576 ( .A(n12503), .B(n12502), .Z(n12504) );
  AND U13577 ( .A(n12505), .B(n12504), .Z(n12523) );
  XOR U13578 ( .A(a[488]), .B(n2245), .Z(n12527) );
  AND U13579 ( .A(a[486]), .B(b[3]), .Z(n12531) );
  AND U13580 ( .A(a[490]), .B(b[0]), .Z(n12507) );
  XNOR U13581 ( .A(n12507), .B(n2175), .Z(n12509) );
  NANDN U13582 ( .A(b[0]), .B(a[489]), .Z(n12508) );
  NAND U13583 ( .A(n12509), .B(n12508), .Z(n12532) );
  XOR U13584 ( .A(n12531), .B(n12532), .Z(n12534) );
  XOR U13585 ( .A(n12533), .B(n12534), .Z(n12522) );
  NANDN U13586 ( .A(n12511), .B(n12510), .Z(n12515) );
  OR U13587 ( .A(n12513), .B(n12512), .Z(n12514) );
  AND U13588 ( .A(n12515), .B(n12514), .Z(n12521) );
  XOR U13589 ( .A(n12522), .B(n12521), .Z(n12524) );
  XOR U13590 ( .A(n12523), .B(n12524), .Z(n12537) );
  XNOR U13591 ( .A(n12537), .B(sreg[1510]), .Z(n12539) );
  NANDN U13592 ( .A(n12516), .B(sreg[1509]), .Z(n12520) );
  NAND U13593 ( .A(n12518), .B(n12517), .Z(n12519) );
  NAND U13594 ( .A(n12520), .B(n12519), .Z(n12538) );
  XOR U13595 ( .A(n12539), .B(n12538), .Z(c[1510]) );
  NANDN U13596 ( .A(n12522), .B(n12521), .Z(n12526) );
  OR U13597 ( .A(n12524), .B(n12523), .Z(n12525) );
  AND U13598 ( .A(n12526), .B(n12525), .Z(n12544) );
  XOR U13599 ( .A(a[489]), .B(n2246), .Z(n12548) );
  AND U13600 ( .A(a[491]), .B(b[0]), .Z(n12528) );
  XNOR U13601 ( .A(n12528), .B(n2175), .Z(n12530) );
  NANDN U13602 ( .A(b[0]), .B(a[490]), .Z(n12529) );
  NAND U13603 ( .A(n12530), .B(n12529), .Z(n12553) );
  AND U13604 ( .A(a[487]), .B(b[3]), .Z(n12552) );
  XOR U13605 ( .A(n12553), .B(n12552), .Z(n12555) );
  XOR U13606 ( .A(n12554), .B(n12555), .Z(n12543) );
  NANDN U13607 ( .A(n12532), .B(n12531), .Z(n12536) );
  OR U13608 ( .A(n12534), .B(n12533), .Z(n12535) );
  AND U13609 ( .A(n12536), .B(n12535), .Z(n12542) );
  XOR U13610 ( .A(n12543), .B(n12542), .Z(n12545) );
  XOR U13611 ( .A(n12544), .B(n12545), .Z(n12558) );
  XNOR U13612 ( .A(n12558), .B(sreg[1511]), .Z(n12560) );
  NANDN U13613 ( .A(n12537), .B(sreg[1510]), .Z(n12541) );
  NAND U13614 ( .A(n12539), .B(n12538), .Z(n12540) );
  NAND U13615 ( .A(n12541), .B(n12540), .Z(n12559) );
  XOR U13616 ( .A(n12560), .B(n12559), .Z(c[1511]) );
  NANDN U13617 ( .A(n12543), .B(n12542), .Z(n12547) );
  OR U13618 ( .A(n12545), .B(n12544), .Z(n12546) );
  AND U13619 ( .A(n12547), .B(n12546), .Z(n12565) );
  XOR U13620 ( .A(a[490]), .B(n2246), .Z(n12569) );
  AND U13621 ( .A(a[492]), .B(b[0]), .Z(n12549) );
  XNOR U13622 ( .A(n12549), .B(n2175), .Z(n12551) );
  NANDN U13623 ( .A(b[0]), .B(a[491]), .Z(n12550) );
  NAND U13624 ( .A(n12551), .B(n12550), .Z(n12574) );
  AND U13625 ( .A(a[488]), .B(b[3]), .Z(n12573) );
  XOR U13626 ( .A(n12574), .B(n12573), .Z(n12576) );
  XOR U13627 ( .A(n12575), .B(n12576), .Z(n12564) );
  NANDN U13628 ( .A(n12553), .B(n12552), .Z(n12557) );
  OR U13629 ( .A(n12555), .B(n12554), .Z(n12556) );
  AND U13630 ( .A(n12557), .B(n12556), .Z(n12563) );
  XOR U13631 ( .A(n12564), .B(n12563), .Z(n12566) );
  XOR U13632 ( .A(n12565), .B(n12566), .Z(n12579) );
  XNOR U13633 ( .A(n12579), .B(sreg[1512]), .Z(n12581) );
  NANDN U13634 ( .A(n12558), .B(sreg[1511]), .Z(n12562) );
  NAND U13635 ( .A(n12560), .B(n12559), .Z(n12561) );
  NAND U13636 ( .A(n12562), .B(n12561), .Z(n12580) );
  XOR U13637 ( .A(n12581), .B(n12580), .Z(c[1512]) );
  NANDN U13638 ( .A(n12564), .B(n12563), .Z(n12568) );
  OR U13639 ( .A(n12566), .B(n12565), .Z(n12567) );
  AND U13640 ( .A(n12568), .B(n12567), .Z(n12586) );
  XOR U13641 ( .A(a[491]), .B(n2246), .Z(n12590) );
  AND U13642 ( .A(a[489]), .B(b[3]), .Z(n12594) );
  AND U13643 ( .A(a[493]), .B(b[0]), .Z(n12570) );
  XNOR U13644 ( .A(n12570), .B(n2175), .Z(n12572) );
  NANDN U13645 ( .A(b[0]), .B(a[492]), .Z(n12571) );
  NAND U13646 ( .A(n12572), .B(n12571), .Z(n12595) );
  XOR U13647 ( .A(n12594), .B(n12595), .Z(n12597) );
  XOR U13648 ( .A(n12596), .B(n12597), .Z(n12585) );
  NANDN U13649 ( .A(n12574), .B(n12573), .Z(n12578) );
  OR U13650 ( .A(n12576), .B(n12575), .Z(n12577) );
  AND U13651 ( .A(n12578), .B(n12577), .Z(n12584) );
  XOR U13652 ( .A(n12585), .B(n12584), .Z(n12587) );
  XOR U13653 ( .A(n12586), .B(n12587), .Z(n12600) );
  XNOR U13654 ( .A(n12600), .B(sreg[1513]), .Z(n12602) );
  NANDN U13655 ( .A(n12579), .B(sreg[1512]), .Z(n12583) );
  NAND U13656 ( .A(n12581), .B(n12580), .Z(n12582) );
  NAND U13657 ( .A(n12583), .B(n12582), .Z(n12601) );
  XOR U13658 ( .A(n12602), .B(n12601), .Z(c[1513]) );
  NANDN U13659 ( .A(n12585), .B(n12584), .Z(n12589) );
  OR U13660 ( .A(n12587), .B(n12586), .Z(n12588) );
  AND U13661 ( .A(n12589), .B(n12588), .Z(n12607) );
  XOR U13662 ( .A(a[492]), .B(n2246), .Z(n12611) );
  AND U13663 ( .A(a[494]), .B(b[0]), .Z(n12591) );
  XNOR U13664 ( .A(n12591), .B(n2175), .Z(n12593) );
  NANDN U13665 ( .A(b[0]), .B(a[493]), .Z(n12592) );
  NAND U13666 ( .A(n12593), .B(n12592), .Z(n12616) );
  AND U13667 ( .A(a[490]), .B(b[3]), .Z(n12615) );
  XOR U13668 ( .A(n12616), .B(n12615), .Z(n12618) );
  XOR U13669 ( .A(n12617), .B(n12618), .Z(n12606) );
  NANDN U13670 ( .A(n12595), .B(n12594), .Z(n12599) );
  OR U13671 ( .A(n12597), .B(n12596), .Z(n12598) );
  AND U13672 ( .A(n12599), .B(n12598), .Z(n12605) );
  XOR U13673 ( .A(n12606), .B(n12605), .Z(n12608) );
  XOR U13674 ( .A(n12607), .B(n12608), .Z(n12621) );
  XNOR U13675 ( .A(n12621), .B(sreg[1514]), .Z(n12623) );
  NANDN U13676 ( .A(n12600), .B(sreg[1513]), .Z(n12604) );
  NAND U13677 ( .A(n12602), .B(n12601), .Z(n12603) );
  NAND U13678 ( .A(n12604), .B(n12603), .Z(n12622) );
  XOR U13679 ( .A(n12623), .B(n12622), .Z(c[1514]) );
  NANDN U13680 ( .A(n12606), .B(n12605), .Z(n12610) );
  OR U13681 ( .A(n12608), .B(n12607), .Z(n12609) );
  AND U13682 ( .A(n12610), .B(n12609), .Z(n12628) );
  XOR U13683 ( .A(a[493]), .B(n2246), .Z(n12632) );
  AND U13684 ( .A(a[491]), .B(b[3]), .Z(n12636) );
  AND U13685 ( .A(a[495]), .B(b[0]), .Z(n12612) );
  XNOR U13686 ( .A(n12612), .B(n2175), .Z(n12614) );
  NANDN U13687 ( .A(b[0]), .B(a[494]), .Z(n12613) );
  NAND U13688 ( .A(n12614), .B(n12613), .Z(n12637) );
  XOR U13689 ( .A(n12636), .B(n12637), .Z(n12639) );
  XOR U13690 ( .A(n12638), .B(n12639), .Z(n12627) );
  NANDN U13691 ( .A(n12616), .B(n12615), .Z(n12620) );
  OR U13692 ( .A(n12618), .B(n12617), .Z(n12619) );
  AND U13693 ( .A(n12620), .B(n12619), .Z(n12626) );
  XOR U13694 ( .A(n12627), .B(n12626), .Z(n12629) );
  XOR U13695 ( .A(n12628), .B(n12629), .Z(n12642) );
  XNOR U13696 ( .A(n12642), .B(sreg[1515]), .Z(n12644) );
  NANDN U13697 ( .A(n12621), .B(sreg[1514]), .Z(n12625) );
  NAND U13698 ( .A(n12623), .B(n12622), .Z(n12624) );
  NAND U13699 ( .A(n12625), .B(n12624), .Z(n12643) );
  XOR U13700 ( .A(n12644), .B(n12643), .Z(c[1515]) );
  NANDN U13701 ( .A(n12627), .B(n12626), .Z(n12631) );
  OR U13702 ( .A(n12629), .B(n12628), .Z(n12630) );
  AND U13703 ( .A(n12631), .B(n12630), .Z(n12650) );
  XOR U13704 ( .A(a[494]), .B(n2246), .Z(n12651) );
  AND U13705 ( .A(b[0]), .B(a[496]), .Z(n12633) );
  XOR U13706 ( .A(b[1]), .B(n12633), .Z(n12635) );
  NANDN U13707 ( .A(b[0]), .B(a[495]), .Z(n12634) );
  AND U13708 ( .A(n12635), .B(n12634), .Z(n12655) );
  AND U13709 ( .A(a[492]), .B(b[3]), .Z(n12656) );
  XOR U13710 ( .A(n12655), .B(n12656), .Z(n12657) );
  XNOR U13711 ( .A(n12658), .B(n12657), .Z(n12647) );
  NANDN U13712 ( .A(n12637), .B(n12636), .Z(n12641) );
  OR U13713 ( .A(n12639), .B(n12638), .Z(n12640) );
  AND U13714 ( .A(n12641), .B(n12640), .Z(n12648) );
  XNOR U13715 ( .A(n12647), .B(n12648), .Z(n12649) );
  XNOR U13716 ( .A(n12650), .B(n12649), .Z(n12661) );
  XNOR U13717 ( .A(n12661), .B(sreg[1516]), .Z(n12663) );
  NANDN U13718 ( .A(n12642), .B(sreg[1515]), .Z(n12646) );
  NAND U13719 ( .A(n12644), .B(n12643), .Z(n12645) );
  NAND U13720 ( .A(n12646), .B(n12645), .Z(n12662) );
  XOR U13721 ( .A(n12663), .B(n12662), .Z(c[1516]) );
  XOR U13722 ( .A(a[495]), .B(n2246), .Z(n12670) );
  AND U13723 ( .A(a[497]), .B(b[0]), .Z(n12652) );
  XNOR U13724 ( .A(n12652), .B(n2175), .Z(n12654) );
  NANDN U13725 ( .A(b[0]), .B(a[496]), .Z(n12653) );
  NAND U13726 ( .A(n12654), .B(n12653), .Z(n12675) );
  AND U13727 ( .A(a[493]), .B(b[3]), .Z(n12674) );
  XOR U13728 ( .A(n12675), .B(n12674), .Z(n12677) );
  XOR U13729 ( .A(n12676), .B(n12677), .Z(n12665) );
  NAND U13730 ( .A(n12656), .B(n12655), .Z(n12660) );
  NANDN U13731 ( .A(n12658), .B(n12657), .Z(n12659) );
  AND U13732 ( .A(n12660), .B(n12659), .Z(n12664) );
  XOR U13733 ( .A(n12665), .B(n12664), .Z(n12667) );
  XOR U13734 ( .A(n12666), .B(n12667), .Z(n12680) );
  XNOR U13735 ( .A(n12680), .B(sreg[1517]), .Z(n12682) );
  XOR U13736 ( .A(n12682), .B(n12681), .Z(c[1517]) );
  NANDN U13737 ( .A(n12665), .B(n12664), .Z(n12669) );
  OR U13738 ( .A(n12667), .B(n12666), .Z(n12668) );
  AND U13739 ( .A(n12669), .B(n12668), .Z(n12687) );
  XOR U13740 ( .A(a[496]), .B(n2247), .Z(n12691) );
  AND U13741 ( .A(a[498]), .B(b[0]), .Z(n12671) );
  XNOR U13742 ( .A(n12671), .B(n2175), .Z(n12673) );
  NANDN U13743 ( .A(b[0]), .B(a[497]), .Z(n12672) );
  NAND U13744 ( .A(n12673), .B(n12672), .Z(n12696) );
  AND U13745 ( .A(a[494]), .B(b[3]), .Z(n12695) );
  XOR U13746 ( .A(n12696), .B(n12695), .Z(n12698) );
  XOR U13747 ( .A(n12697), .B(n12698), .Z(n12686) );
  NANDN U13748 ( .A(n12675), .B(n12674), .Z(n12679) );
  OR U13749 ( .A(n12677), .B(n12676), .Z(n12678) );
  AND U13750 ( .A(n12679), .B(n12678), .Z(n12685) );
  XOR U13751 ( .A(n12686), .B(n12685), .Z(n12688) );
  XOR U13752 ( .A(n12687), .B(n12688), .Z(n12701) );
  XNOR U13753 ( .A(n12701), .B(sreg[1518]), .Z(n12703) );
  NANDN U13754 ( .A(n12680), .B(sreg[1517]), .Z(n12684) );
  NAND U13755 ( .A(n12682), .B(n12681), .Z(n12683) );
  NAND U13756 ( .A(n12684), .B(n12683), .Z(n12702) );
  XOR U13757 ( .A(n12703), .B(n12702), .Z(c[1518]) );
  NANDN U13758 ( .A(n12686), .B(n12685), .Z(n12690) );
  OR U13759 ( .A(n12688), .B(n12687), .Z(n12689) );
  AND U13760 ( .A(n12690), .B(n12689), .Z(n12708) );
  XOR U13761 ( .A(a[497]), .B(n2247), .Z(n12712) );
  AND U13762 ( .A(a[499]), .B(b[0]), .Z(n12692) );
  XNOR U13763 ( .A(n12692), .B(n2175), .Z(n12694) );
  NANDN U13764 ( .A(b[0]), .B(a[498]), .Z(n12693) );
  NAND U13765 ( .A(n12694), .B(n12693), .Z(n12717) );
  AND U13766 ( .A(a[495]), .B(b[3]), .Z(n12716) );
  XOR U13767 ( .A(n12717), .B(n12716), .Z(n12719) );
  XOR U13768 ( .A(n12718), .B(n12719), .Z(n12707) );
  NANDN U13769 ( .A(n12696), .B(n12695), .Z(n12700) );
  OR U13770 ( .A(n12698), .B(n12697), .Z(n12699) );
  AND U13771 ( .A(n12700), .B(n12699), .Z(n12706) );
  XOR U13772 ( .A(n12707), .B(n12706), .Z(n12709) );
  XOR U13773 ( .A(n12708), .B(n12709), .Z(n12722) );
  XNOR U13774 ( .A(n12722), .B(sreg[1519]), .Z(n12724) );
  NANDN U13775 ( .A(n12701), .B(sreg[1518]), .Z(n12705) );
  NAND U13776 ( .A(n12703), .B(n12702), .Z(n12704) );
  NAND U13777 ( .A(n12705), .B(n12704), .Z(n12723) );
  XOR U13778 ( .A(n12724), .B(n12723), .Z(c[1519]) );
  NANDN U13779 ( .A(n12707), .B(n12706), .Z(n12711) );
  OR U13780 ( .A(n12709), .B(n12708), .Z(n12710) );
  AND U13781 ( .A(n12711), .B(n12710), .Z(n12729) );
  XOR U13782 ( .A(a[498]), .B(n2247), .Z(n12733) );
  AND U13783 ( .A(a[500]), .B(b[0]), .Z(n12713) );
  XNOR U13784 ( .A(n12713), .B(n2175), .Z(n12715) );
  NANDN U13785 ( .A(b[0]), .B(a[499]), .Z(n12714) );
  NAND U13786 ( .A(n12715), .B(n12714), .Z(n12738) );
  AND U13787 ( .A(a[496]), .B(b[3]), .Z(n12737) );
  XOR U13788 ( .A(n12738), .B(n12737), .Z(n12740) );
  XOR U13789 ( .A(n12739), .B(n12740), .Z(n12728) );
  NANDN U13790 ( .A(n12717), .B(n12716), .Z(n12721) );
  OR U13791 ( .A(n12719), .B(n12718), .Z(n12720) );
  AND U13792 ( .A(n12721), .B(n12720), .Z(n12727) );
  XOR U13793 ( .A(n12728), .B(n12727), .Z(n12730) );
  XOR U13794 ( .A(n12729), .B(n12730), .Z(n12743) );
  XNOR U13795 ( .A(n12743), .B(sreg[1520]), .Z(n12745) );
  NANDN U13796 ( .A(n12722), .B(sreg[1519]), .Z(n12726) );
  NAND U13797 ( .A(n12724), .B(n12723), .Z(n12725) );
  NAND U13798 ( .A(n12726), .B(n12725), .Z(n12744) );
  XOR U13799 ( .A(n12745), .B(n12744), .Z(c[1520]) );
  NANDN U13800 ( .A(n12728), .B(n12727), .Z(n12732) );
  OR U13801 ( .A(n12730), .B(n12729), .Z(n12731) );
  AND U13802 ( .A(n12732), .B(n12731), .Z(n12750) );
  XOR U13803 ( .A(a[499]), .B(n2247), .Z(n12754) );
  AND U13804 ( .A(a[501]), .B(b[0]), .Z(n12734) );
  XNOR U13805 ( .A(n12734), .B(n2175), .Z(n12736) );
  NANDN U13806 ( .A(b[0]), .B(a[500]), .Z(n12735) );
  NAND U13807 ( .A(n12736), .B(n12735), .Z(n12759) );
  AND U13808 ( .A(a[497]), .B(b[3]), .Z(n12758) );
  XOR U13809 ( .A(n12759), .B(n12758), .Z(n12761) );
  XOR U13810 ( .A(n12760), .B(n12761), .Z(n12749) );
  NANDN U13811 ( .A(n12738), .B(n12737), .Z(n12742) );
  OR U13812 ( .A(n12740), .B(n12739), .Z(n12741) );
  AND U13813 ( .A(n12742), .B(n12741), .Z(n12748) );
  XOR U13814 ( .A(n12749), .B(n12748), .Z(n12751) );
  XOR U13815 ( .A(n12750), .B(n12751), .Z(n12764) );
  XNOR U13816 ( .A(n12764), .B(sreg[1521]), .Z(n12766) );
  NANDN U13817 ( .A(n12743), .B(sreg[1520]), .Z(n12747) );
  NAND U13818 ( .A(n12745), .B(n12744), .Z(n12746) );
  NAND U13819 ( .A(n12747), .B(n12746), .Z(n12765) );
  XOR U13820 ( .A(n12766), .B(n12765), .Z(c[1521]) );
  NANDN U13821 ( .A(n12749), .B(n12748), .Z(n12753) );
  OR U13822 ( .A(n12751), .B(n12750), .Z(n12752) );
  AND U13823 ( .A(n12753), .B(n12752), .Z(n12771) );
  XOR U13824 ( .A(a[500]), .B(n2247), .Z(n12775) );
  AND U13825 ( .A(a[502]), .B(b[0]), .Z(n12755) );
  XNOR U13826 ( .A(n12755), .B(n2175), .Z(n12757) );
  NANDN U13827 ( .A(b[0]), .B(a[501]), .Z(n12756) );
  NAND U13828 ( .A(n12757), .B(n12756), .Z(n12780) );
  AND U13829 ( .A(a[498]), .B(b[3]), .Z(n12779) );
  XOR U13830 ( .A(n12780), .B(n12779), .Z(n12782) );
  XOR U13831 ( .A(n12781), .B(n12782), .Z(n12770) );
  NANDN U13832 ( .A(n12759), .B(n12758), .Z(n12763) );
  OR U13833 ( .A(n12761), .B(n12760), .Z(n12762) );
  AND U13834 ( .A(n12763), .B(n12762), .Z(n12769) );
  XOR U13835 ( .A(n12770), .B(n12769), .Z(n12772) );
  XOR U13836 ( .A(n12771), .B(n12772), .Z(n12785) );
  XNOR U13837 ( .A(n12785), .B(sreg[1522]), .Z(n12787) );
  NANDN U13838 ( .A(n12764), .B(sreg[1521]), .Z(n12768) );
  NAND U13839 ( .A(n12766), .B(n12765), .Z(n12767) );
  NAND U13840 ( .A(n12768), .B(n12767), .Z(n12786) );
  XOR U13841 ( .A(n12787), .B(n12786), .Z(c[1522]) );
  NANDN U13842 ( .A(n12770), .B(n12769), .Z(n12774) );
  OR U13843 ( .A(n12772), .B(n12771), .Z(n12773) );
  AND U13844 ( .A(n12774), .B(n12773), .Z(n12792) );
  XOR U13845 ( .A(a[501]), .B(n2247), .Z(n12796) );
  AND U13846 ( .A(a[499]), .B(b[3]), .Z(n12800) );
  AND U13847 ( .A(a[503]), .B(b[0]), .Z(n12776) );
  XNOR U13848 ( .A(n12776), .B(n2175), .Z(n12778) );
  NANDN U13849 ( .A(b[0]), .B(a[502]), .Z(n12777) );
  NAND U13850 ( .A(n12778), .B(n12777), .Z(n12801) );
  XOR U13851 ( .A(n12800), .B(n12801), .Z(n12803) );
  XOR U13852 ( .A(n12802), .B(n12803), .Z(n12791) );
  NANDN U13853 ( .A(n12780), .B(n12779), .Z(n12784) );
  OR U13854 ( .A(n12782), .B(n12781), .Z(n12783) );
  AND U13855 ( .A(n12784), .B(n12783), .Z(n12790) );
  XOR U13856 ( .A(n12791), .B(n12790), .Z(n12793) );
  XOR U13857 ( .A(n12792), .B(n12793), .Z(n12806) );
  XNOR U13858 ( .A(n12806), .B(sreg[1523]), .Z(n12808) );
  NANDN U13859 ( .A(n12785), .B(sreg[1522]), .Z(n12789) );
  NAND U13860 ( .A(n12787), .B(n12786), .Z(n12788) );
  NAND U13861 ( .A(n12789), .B(n12788), .Z(n12807) );
  XOR U13862 ( .A(n12808), .B(n12807), .Z(c[1523]) );
  NANDN U13863 ( .A(n12791), .B(n12790), .Z(n12795) );
  OR U13864 ( .A(n12793), .B(n12792), .Z(n12794) );
  AND U13865 ( .A(n12795), .B(n12794), .Z(n12813) );
  XOR U13866 ( .A(a[502]), .B(n2247), .Z(n12817) );
  AND U13867 ( .A(a[504]), .B(b[0]), .Z(n12797) );
  XNOR U13868 ( .A(n12797), .B(n2175), .Z(n12799) );
  NANDN U13869 ( .A(b[0]), .B(a[503]), .Z(n12798) );
  NAND U13870 ( .A(n12799), .B(n12798), .Z(n12822) );
  AND U13871 ( .A(a[500]), .B(b[3]), .Z(n12821) );
  XOR U13872 ( .A(n12822), .B(n12821), .Z(n12824) );
  XOR U13873 ( .A(n12823), .B(n12824), .Z(n12812) );
  NANDN U13874 ( .A(n12801), .B(n12800), .Z(n12805) );
  OR U13875 ( .A(n12803), .B(n12802), .Z(n12804) );
  AND U13876 ( .A(n12805), .B(n12804), .Z(n12811) );
  XOR U13877 ( .A(n12812), .B(n12811), .Z(n12814) );
  XOR U13878 ( .A(n12813), .B(n12814), .Z(n12827) );
  XNOR U13879 ( .A(n12827), .B(sreg[1524]), .Z(n12829) );
  NANDN U13880 ( .A(n12806), .B(sreg[1523]), .Z(n12810) );
  NAND U13881 ( .A(n12808), .B(n12807), .Z(n12809) );
  NAND U13882 ( .A(n12810), .B(n12809), .Z(n12828) );
  XOR U13883 ( .A(n12829), .B(n12828), .Z(c[1524]) );
  NANDN U13884 ( .A(n12812), .B(n12811), .Z(n12816) );
  OR U13885 ( .A(n12814), .B(n12813), .Z(n12815) );
  AND U13886 ( .A(n12816), .B(n12815), .Z(n12834) );
  XOR U13887 ( .A(a[503]), .B(n2248), .Z(n12838) );
  AND U13888 ( .A(a[505]), .B(b[0]), .Z(n12818) );
  XNOR U13889 ( .A(n12818), .B(n2175), .Z(n12820) );
  NANDN U13890 ( .A(b[0]), .B(a[504]), .Z(n12819) );
  NAND U13891 ( .A(n12820), .B(n12819), .Z(n12843) );
  AND U13892 ( .A(a[501]), .B(b[3]), .Z(n12842) );
  XOR U13893 ( .A(n12843), .B(n12842), .Z(n12845) );
  XOR U13894 ( .A(n12844), .B(n12845), .Z(n12833) );
  NANDN U13895 ( .A(n12822), .B(n12821), .Z(n12826) );
  OR U13896 ( .A(n12824), .B(n12823), .Z(n12825) );
  AND U13897 ( .A(n12826), .B(n12825), .Z(n12832) );
  XOR U13898 ( .A(n12833), .B(n12832), .Z(n12835) );
  XOR U13899 ( .A(n12834), .B(n12835), .Z(n12848) );
  XNOR U13900 ( .A(n12848), .B(sreg[1525]), .Z(n12850) );
  NANDN U13901 ( .A(n12827), .B(sreg[1524]), .Z(n12831) );
  NAND U13902 ( .A(n12829), .B(n12828), .Z(n12830) );
  NAND U13903 ( .A(n12831), .B(n12830), .Z(n12849) );
  XOR U13904 ( .A(n12850), .B(n12849), .Z(c[1525]) );
  NANDN U13905 ( .A(n12833), .B(n12832), .Z(n12837) );
  OR U13906 ( .A(n12835), .B(n12834), .Z(n12836) );
  AND U13907 ( .A(n12837), .B(n12836), .Z(n12855) );
  XOR U13908 ( .A(a[504]), .B(n2248), .Z(n12859) );
  AND U13909 ( .A(a[502]), .B(b[3]), .Z(n12863) );
  AND U13910 ( .A(a[506]), .B(b[0]), .Z(n12839) );
  XNOR U13911 ( .A(n12839), .B(n2175), .Z(n12841) );
  NANDN U13912 ( .A(b[0]), .B(a[505]), .Z(n12840) );
  NAND U13913 ( .A(n12841), .B(n12840), .Z(n12864) );
  XOR U13914 ( .A(n12863), .B(n12864), .Z(n12866) );
  XOR U13915 ( .A(n12865), .B(n12866), .Z(n12854) );
  NANDN U13916 ( .A(n12843), .B(n12842), .Z(n12847) );
  OR U13917 ( .A(n12845), .B(n12844), .Z(n12846) );
  AND U13918 ( .A(n12847), .B(n12846), .Z(n12853) );
  XOR U13919 ( .A(n12854), .B(n12853), .Z(n12856) );
  XOR U13920 ( .A(n12855), .B(n12856), .Z(n12869) );
  XNOR U13921 ( .A(n12869), .B(sreg[1526]), .Z(n12871) );
  NANDN U13922 ( .A(n12848), .B(sreg[1525]), .Z(n12852) );
  NAND U13923 ( .A(n12850), .B(n12849), .Z(n12851) );
  NAND U13924 ( .A(n12852), .B(n12851), .Z(n12870) );
  XOR U13925 ( .A(n12871), .B(n12870), .Z(c[1526]) );
  NANDN U13926 ( .A(n12854), .B(n12853), .Z(n12858) );
  OR U13927 ( .A(n12856), .B(n12855), .Z(n12857) );
  AND U13928 ( .A(n12858), .B(n12857), .Z(n12876) );
  XOR U13929 ( .A(a[505]), .B(n2248), .Z(n12880) );
  AND U13930 ( .A(a[507]), .B(b[0]), .Z(n12860) );
  XNOR U13931 ( .A(n12860), .B(n2175), .Z(n12862) );
  NANDN U13932 ( .A(b[0]), .B(a[506]), .Z(n12861) );
  NAND U13933 ( .A(n12862), .B(n12861), .Z(n12885) );
  AND U13934 ( .A(a[503]), .B(b[3]), .Z(n12884) );
  XOR U13935 ( .A(n12885), .B(n12884), .Z(n12887) );
  XOR U13936 ( .A(n12886), .B(n12887), .Z(n12875) );
  NANDN U13937 ( .A(n12864), .B(n12863), .Z(n12868) );
  OR U13938 ( .A(n12866), .B(n12865), .Z(n12867) );
  AND U13939 ( .A(n12868), .B(n12867), .Z(n12874) );
  XOR U13940 ( .A(n12875), .B(n12874), .Z(n12877) );
  XOR U13941 ( .A(n12876), .B(n12877), .Z(n12890) );
  XNOR U13942 ( .A(n12890), .B(sreg[1527]), .Z(n12892) );
  NANDN U13943 ( .A(n12869), .B(sreg[1526]), .Z(n12873) );
  NAND U13944 ( .A(n12871), .B(n12870), .Z(n12872) );
  NAND U13945 ( .A(n12873), .B(n12872), .Z(n12891) );
  XOR U13946 ( .A(n12892), .B(n12891), .Z(c[1527]) );
  NANDN U13947 ( .A(n12875), .B(n12874), .Z(n12879) );
  OR U13948 ( .A(n12877), .B(n12876), .Z(n12878) );
  AND U13949 ( .A(n12879), .B(n12878), .Z(n12897) );
  XOR U13950 ( .A(a[506]), .B(n2248), .Z(n12901) );
  AND U13951 ( .A(a[504]), .B(b[3]), .Z(n12905) );
  AND U13952 ( .A(a[508]), .B(b[0]), .Z(n12881) );
  XNOR U13953 ( .A(n12881), .B(n2175), .Z(n12883) );
  NANDN U13954 ( .A(b[0]), .B(a[507]), .Z(n12882) );
  NAND U13955 ( .A(n12883), .B(n12882), .Z(n12906) );
  XOR U13956 ( .A(n12905), .B(n12906), .Z(n12908) );
  XOR U13957 ( .A(n12907), .B(n12908), .Z(n12896) );
  NANDN U13958 ( .A(n12885), .B(n12884), .Z(n12889) );
  OR U13959 ( .A(n12887), .B(n12886), .Z(n12888) );
  AND U13960 ( .A(n12889), .B(n12888), .Z(n12895) );
  XOR U13961 ( .A(n12896), .B(n12895), .Z(n12898) );
  XOR U13962 ( .A(n12897), .B(n12898), .Z(n12911) );
  XNOR U13963 ( .A(n12911), .B(sreg[1528]), .Z(n12913) );
  NANDN U13964 ( .A(n12890), .B(sreg[1527]), .Z(n12894) );
  NAND U13965 ( .A(n12892), .B(n12891), .Z(n12893) );
  NAND U13966 ( .A(n12894), .B(n12893), .Z(n12912) );
  XOR U13967 ( .A(n12913), .B(n12912), .Z(c[1528]) );
  NANDN U13968 ( .A(n12896), .B(n12895), .Z(n12900) );
  OR U13969 ( .A(n12898), .B(n12897), .Z(n12899) );
  AND U13970 ( .A(n12900), .B(n12899), .Z(n12918) );
  XOR U13971 ( .A(a[507]), .B(n2248), .Z(n12922) );
  AND U13972 ( .A(a[509]), .B(b[0]), .Z(n12902) );
  XNOR U13973 ( .A(n12902), .B(n2175), .Z(n12904) );
  NANDN U13974 ( .A(b[0]), .B(a[508]), .Z(n12903) );
  NAND U13975 ( .A(n12904), .B(n12903), .Z(n12927) );
  AND U13976 ( .A(a[505]), .B(b[3]), .Z(n12926) );
  XOR U13977 ( .A(n12927), .B(n12926), .Z(n12929) );
  XOR U13978 ( .A(n12928), .B(n12929), .Z(n12917) );
  NANDN U13979 ( .A(n12906), .B(n12905), .Z(n12910) );
  OR U13980 ( .A(n12908), .B(n12907), .Z(n12909) );
  AND U13981 ( .A(n12910), .B(n12909), .Z(n12916) );
  XOR U13982 ( .A(n12917), .B(n12916), .Z(n12919) );
  XOR U13983 ( .A(n12918), .B(n12919), .Z(n12932) );
  XNOR U13984 ( .A(n12932), .B(sreg[1529]), .Z(n12934) );
  NANDN U13985 ( .A(n12911), .B(sreg[1528]), .Z(n12915) );
  NAND U13986 ( .A(n12913), .B(n12912), .Z(n12914) );
  NAND U13987 ( .A(n12915), .B(n12914), .Z(n12933) );
  XOR U13988 ( .A(n12934), .B(n12933), .Z(c[1529]) );
  NANDN U13989 ( .A(n12917), .B(n12916), .Z(n12921) );
  OR U13990 ( .A(n12919), .B(n12918), .Z(n12920) );
  AND U13991 ( .A(n12921), .B(n12920), .Z(n12939) );
  XOR U13992 ( .A(a[508]), .B(n2248), .Z(n12943) );
  AND U13993 ( .A(a[510]), .B(b[0]), .Z(n12923) );
  XNOR U13994 ( .A(n12923), .B(n2175), .Z(n12925) );
  NANDN U13995 ( .A(b[0]), .B(a[509]), .Z(n12924) );
  NAND U13996 ( .A(n12925), .B(n12924), .Z(n12948) );
  AND U13997 ( .A(a[506]), .B(b[3]), .Z(n12947) );
  XOR U13998 ( .A(n12948), .B(n12947), .Z(n12950) );
  XOR U13999 ( .A(n12949), .B(n12950), .Z(n12938) );
  NANDN U14000 ( .A(n12927), .B(n12926), .Z(n12931) );
  OR U14001 ( .A(n12929), .B(n12928), .Z(n12930) );
  AND U14002 ( .A(n12931), .B(n12930), .Z(n12937) );
  XOR U14003 ( .A(n12938), .B(n12937), .Z(n12940) );
  XOR U14004 ( .A(n12939), .B(n12940), .Z(n12953) );
  XNOR U14005 ( .A(n12953), .B(sreg[1530]), .Z(n12955) );
  NANDN U14006 ( .A(n12932), .B(sreg[1529]), .Z(n12936) );
  NAND U14007 ( .A(n12934), .B(n12933), .Z(n12935) );
  NAND U14008 ( .A(n12936), .B(n12935), .Z(n12954) );
  XOR U14009 ( .A(n12955), .B(n12954), .Z(c[1530]) );
  NANDN U14010 ( .A(n12938), .B(n12937), .Z(n12942) );
  OR U14011 ( .A(n12940), .B(n12939), .Z(n12941) );
  AND U14012 ( .A(n12942), .B(n12941), .Z(n12960) );
  XOR U14013 ( .A(a[509]), .B(n2248), .Z(n12964) );
  AND U14014 ( .A(a[511]), .B(b[0]), .Z(n12944) );
  XNOR U14015 ( .A(n12944), .B(n2175), .Z(n12946) );
  NANDN U14016 ( .A(b[0]), .B(a[510]), .Z(n12945) );
  NAND U14017 ( .A(n12946), .B(n12945), .Z(n12969) );
  AND U14018 ( .A(a[507]), .B(b[3]), .Z(n12968) );
  XOR U14019 ( .A(n12969), .B(n12968), .Z(n12971) );
  XOR U14020 ( .A(n12970), .B(n12971), .Z(n12959) );
  NANDN U14021 ( .A(n12948), .B(n12947), .Z(n12952) );
  OR U14022 ( .A(n12950), .B(n12949), .Z(n12951) );
  AND U14023 ( .A(n12952), .B(n12951), .Z(n12958) );
  XOR U14024 ( .A(n12959), .B(n12958), .Z(n12961) );
  XOR U14025 ( .A(n12960), .B(n12961), .Z(n12974) );
  XNOR U14026 ( .A(n12974), .B(sreg[1531]), .Z(n12976) );
  NANDN U14027 ( .A(n12953), .B(sreg[1530]), .Z(n12957) );
  NAND U14028 ( .A(n12955), .B(n12954), .Z(n12956) );
  NAND U14029 ( .A(n12957), .B(n12956), .Z(n12975) );
  XOR U14030 ( .A(n12976), .B(n12975), .Z(c[1531]) );
  NANDN U14031 ( .A(n12959), .B(n12958), .Z(n12963) );
  OR U14032 ( .A(n12961), .B(n12960), .Z(n12962) );
  AND U14033 ( .A(n12963), .B(n12962), .Z(n12981) );
  XOR U14034 ( .A(a[510]), .B(n2249), .Z(n12985) );
  AND U14035 ( .A(a[512]), .B(b[0]), .Z(n12965) );
  XNOR U14036 ( .A(n12965), .B(n2175), .Z(n12967) );
  NANDN U14037 ( .A(b[0]), .B(a[511]), .Z(n12966) );
  NAND U14038 ( .A(n12967), .B(n12966), .Z(n12990) );
  AND U14039 ( .A(a[508]), .B(b[3]), .Z(n12989) );
  XOR U14040 ( .A(n12990), .B(n12989), .Z(n12992) );
  XOR U14041 ( .A(n12991), .B(n12992), .Z(n12980) );
  NANDN U14042 ( .A(n12969), .B(n12968), .Z(n12973) );
  OR U14043 ( .A(n12971), .B(n12970), .Z(n12972) );
  AND U14044 ( .A(n12973), .B(n12972), .Z(n12979) );
  XOR U14045 ( .A(n12980), .B(n12979), .Z(n12982) );
  XOR U14046 ( .A(n12981), .B(n12982), .Z(n12995) );
  XNOR U14047 ( .A(n12995), .B(sreg[1532]), .Z(n12997) );
  NANDN U14048 ( .A(n12974), .B(sreg[1531]), .Z(n12978) );
  NAND U14049 ( .A(n12976), .B(n12975), .Z(n12977) );
  NAND U14050 ( .A(n12978), .B(n12977), .Z(n12996) );
  XOR U14051 ( .A(n12997), .B(n12996), .Z(c[1532]) );
  NANDN U14052 ( .A(n12980), .B(n12979), .Z(n12984) );
  OR U14053 ( .A(n12982), .B(n12981), .Z(n12983) );
  AND U14054 ( .A(n12984), .B(n12983), .Z(n13002) );
  XOR U14055 ( .A(a[511]), .B(n2249), .Z(n13006) );
  AND U14056 ( .A(a[513]), .B(b[0]), .Z(n12986) );
  XNOR U14057 ( .A(n12986), .B(n2175), .Z(n12988) );
  NANDN U14058 ( .A(b[0]), .B(a[512]), .Z(n12987) );
  NAND U14059 ( .A(n12988), .B(n12987), .Z(n13011) );
  AND U14060 ( .A(a[509]), .B(b[3]), .Z(n13010) );
  XOR U14061 ( .A(n13011), .B(n13010), .Z(n13013) );
  XOR U14062 ( .A(n13012), .B(n13013), .Z(n13001) );
  NANDN U14063 ( .A(n12990), .B(n12989), .Z(n12994) );
  OR U14064 ( .A(n12992), .B(n12991), .Z(n12993) );
  AND U14065 ( .A(n12994), .B(n12993), .Z(n13000) );
  XOR U14066 ( .A(n13001), .B(n13000), .Z(n13003) );
  XOR U14067 ( .A(n13002), .B(n13003), .Z(n13016) );
  XNOR U14068 ( .A(n13016), .B(sreg[1533]), .Z(n13018) );
  NANDN U14069 ( .A(n12995), .B(sreg[1532]), .Z(n12999) );
  NAND U14070 ( .A(n12997), .B(n12996), .Z(n12998) );
  NAND U14071 ( .A(n12999), .B(n12998), .Z(n13017) );
  XOR U14072 ( .A(n13018), .B(n13017), .Z(c[1533]) );
  NANDN U14073 ( .A(n13001), .B(n13000), .Z(n13005) );
  OR U14074 ( .A(n13003), .B(n13002), .Z(n13004) );
  AND U14075 ( .A(n13005), .B(n13004), .Z(n13023) );
  XOR U14076 ( .A(a[512]), .B(n2249), .Z(n13027) );
  AND U14077 ( .A(a[514]), .B(b[0]), .Z(n13007) );
  XNOR U14078 ( .A(n13007), .B(n2175), .Z(n13009) );
  NANDN U14079 ( .A(b[0]), .B(a[513]), .Z(n13008) );
  NAND U14080 ( .A(n13009), .B(n13008), .Z(n13032) );
  AND U14081 ( .A(a[510]), .B(b[3]), .Z(n13031) );
  XOR U14082 ( .A(n13032), .B(n13031), .Z(n13034) );
  XOR U14083 ( .A(n13033), .B(n13034), .Z(n13022) );
  NANDN U14084 ( .A(n13011), .B(n13010), .Z(n13015) );
  OR U14085 ( .A(n13013), .B(n13012), .Z(n13014) );
  AND U14086 ( .A(n13015), .B(n13014), .Z(n13021) );
  XOR U14087 ( .A(n13022), .B(n13021), .Z(n13024) );
  XOR U14088 ( .A(n13023), .B(n13024), .Z(n13037) );
  XNOR U14089 ( .A(n13037), .B(sreg[1534]), .Z(n13039) );
  NANDN U14090 ( .A(n13016), .B(sreg[1533]), .Z(n13020) );
  NAND U14091 ( .A(n13018), .B(n13017), .Z(n13019) );
  NAND U14092 ( .A(n13020), .B(n13019), .Z(n13038) );
  XOR U14093 ( .A(n13039), .B(n13038), .Z(c[1534]) );
  NANDN U14094 ( .A(n13022), .B(n13021), .Z(n13026) );
  OR U14095 ( .A(n13024), .B(n13023), .Z(n13025) );
  AND U14096 ( .A(n13026), .B(n13025), .Z(n13044) );
  XOR U14097 ( .A(a[513]), .B(n2249), .Z(n13048) );
  AND U14098 ( .A(a[515]), .B(b[0]), .Z(n13028) );
  XNOR U14099 ( .A(n13028), .B(n2175), .Z(n13030) );
  NANDN U14100 ( .A(b[0]), .B(a[514]), .Z(n13029) );
  NAND U14101 ( .A(n13030), .B(n13029), .Z(n13053) );
  AND U14102 ( .A(a[511]), .B(b[3]), .Z(n13052) );
  XOR U14103 ( .A(n13053), .B(n13052), .Z(n13055) );
  XOR U14104 ( .A(n13054), .B(n13055), .Z(n13043) );
  NANDN U14105 ( .A(n13032), .B(n13031), .Z(n13036) );
  OR U14106 ( .A(n13034), .B(n13033), .Z(n13035) );
  AND U14107 ( .A(n13036), .B(n13035), .Z(n13042) );
  XOR U14108 ( .A(n13043), .B(n13042), .Z(n13045) );
  XOR U14109 ( .A(n13044), .B(n13045), .Z(n13058) );
  XNOR U14110 ( .A(n13058), .B(sreg[1535]), .Z(n13060) );
  NANDN U14111 ( .A(n13037), .B(sreg[1534]), .Z(n13041) );
  NAND U14112 ( .A(n13039), .B(n13038), .Z(n13040) );
  NAND U14113 ( .A(n13041), .B(n13040), .Z(n13059) );
  XOR U14114 ( .A(n13060), .B(n13059), .Z(c[1535]) );
  NANDN U14115 ( .A(n13043), .B(n13042), .Z(n13047) );
  OR U14116 ( .A(n13045), .B(n13044), .Z(n13046) );
  AND U14117 ( .A(n13047), .B(n13046), .Z(n13065) );
  XOR U14118 ( .A(a[514]), .B(n2249), .Z(n13069) );
  AND U14119 ( .A(a[512]), .B(b[3]), .Z(n13073) );
  AND U14120 ( .A(a[516]), .B(b[0]), .Z(n13049) );
  XNOR U14121 ( .A(n13049), .B(n2175), .Z(n13051) );
  NANDN U14122 ( .A(b[0]), .B(a[515]), .Z(n13050) );
  NAND U14123 ( .A(n13051), .B(n13050), .Z(n13074) );
  XOR U14124 ( .A(n13073), .B(n13074), .Z(n13076) );
  XOR U14125 ( .A(n13075), .B(n13076), .Z(n13064) );
  NANDN U14126 ( .A(n13053), .B(n13052), .Z(n13057) );
  OR U14127 ( .A(n13055), .B(n13054), .Z(n13056) );
  AND U14128 ( .A(n13057), .B(n13056), .Z(n13063) );
  XOR U14129 ( .A(n13064), .B(n13063), .Z(n13066) );
  XOR U14130 ( .A(n13065), .B(n13066), .Z(n13079) );
  XNOR U14131 ( .A(n13079), .B(sreg[1536]), .Z(n13081) );
  NANDN U14132 ( .A(n13058), .B(sreg[1535]), .Z(n13062) );
  NAND U14133 ( .A(n13060), .B(n13059), .Z(n13061) );
  NAND U14134 ( .A(n13062), .B(n13061), .Z(n13080) );
  XOR U14135 ( .A(n13081), .B(n13080), .Z(c[1536]) );
  NANDN U14136 ( .A(n13064), .B(n13063), .Z(n13068) );
  OR U14137 ( .A(n13066), .B(n13065), .Z(n13067) );
  AND U14138 ( .A(n13068), .B(n13067), .Z(n13086) );
  XOR U14139 ( .A(a[515]), .B(n2249), .Z(n13090) );
  AND U14140 ( .A(a[513]), .B(b[3]), .Z(n13094) );
  AND U14141 ( .A(a[517]), .B(b[0]), .Z(n13070) );
  XNOR U14142 ( .A(n13070), .B(n2175), .Z(n13072) );
  NANDN U14143 ( .A(b[0]), .B(a[516]), .Z(n13071) );
  NAND U14144 ( .A(n13072), .B(n13071), .Z(n13095) );
  XOR U14145 ( .A(n13094), .B(n13095), .Z(n13097) );
  XOR U14146 ( .A(n13096), .B(n13097), .Z(n13085) );
  NANDN U14147 ( .A(n13074), .B(n13073), .Z(n13078) );
  OR U14148 ( .A(n13076), .B(n13075), .Z(n13077) );
  AND U14149 ( .A(n13078), .B(n13077), .Z(n13084) );
  XOR U14150 ( .A(n13085), .B(n13084), .Z(n13087) );
  XOR U14151 ( .A(n13086), .B(n13087), .Z(n13100) );
  XNOR U14152 ( .A(n13100), .B(sreg[1537]), .Z(n13102) );
  NANDN U14153 ( .A(n13079), .B(sreg[1536]), .Z(n13083) );
  NAND U14154 ( .A(n13081), .B(n13080), .Z(n13082) );
  NAND U14155 ( .A(n13083), .B(n13082), .Z(n13101) );
  XOR U14156 ( .A(n13102), .B(n13101), .Z(c[1537]) );
  NANDN U14157 ( .A(n13085), .B(n13084), .Z(n13089) );
  OR U14158 ( .A(n13087), .B(n13086), .Z(n13088) );
  AND U14159 ( .A(n13089), .B(n13088), .Z(n13107) );
  XOR U14160 ( .A(a[516]), .B(n2249), .Z(n13111) );
  AND U14161 ( .A(a[518]), .B(b[0]), .Z(n13091) );
  XNOR U14162 ( .A(n13091), .B(n2175), .Z(n13093) );
  NANDN U14163 ( .A(b[0]), .B(a[517]), .Z(n13092) );
  NAND U14164 ( .A(n13093), .B(n13092), .Z(n13116) );
  AND U14165 ( .A(a[514]), .B(b[3]), .Z(n13115) );
  XOR U14166 ( .A(n13116), .B(n13115), .Z(n13118) );
  XOR U14167 ( .A(n13117), .B(n13118), .Z(n13106) );
  NANDN U14168 ( .A(n13095), .B(n13094), .Z(n13099) );
  OR U14169 ( .A(n13097), .B(n13096), .Z(n13098) );
  AND U14170 ( .A(n13099), .B(n13098), .Z(n13105) );
  XOR U14171 ( .A(n13106), .B(n13105), .Z(n13108) );
  XOR U14172 ( .A(n13107), .B(n13108), .Z(n13121) );
  XNOR U14173 ( .A(n13121), .B(sreg[1538]), .Z(n13123) );
  NANDN U14174 ( .A(n13100), .B(sreg[1537]), .Z(n13104) );
  NAND U14175 ( .A(n13102), .B(n13101), .Z(n13103) );
  NAND U14176 ( .A(n13104), .B(n13103), .Z(n13122) );
  XOR U14177 ( .A(n13123), .B(n13122), .Z(c[1538]) );
  NANDN U14178 ( .A(n13106), .B(n13105), .Z(n13110) );
  OR U14179 ( .A(n13108), .B(n13107), .Z(n13109) );
  AND U14180 ( .A(n13110), .B(n13109), .Z(n13128) );
  XOR U14181 ( .A(a[517]), .B(n2250), .Z(n13132) );
  AND U14182 ( .A(a[515]), .B(b[3]), .Z(n13136) );
  AND U14183 ( .A(a[519]), .B(b[0]), .Z(n13112) );
  XNOR U14184 ( .A(n13112), .B(n2175), .Z(n13114) );
  NANDN U14185 ( .A(b[0]), .B(a[518]), .Z(n13113) );
  NAND U14186 ( .A(n13114), .B(n13113), .Z(n13137) );
  XOR U14187 ( .A(n13136), .B(n13137), .Z(n13139) );
  XOR U14188 ( .A(n13138), .B(n13139), .Z(n13127) );
  NANDN U14189 ( .A(n13116), .B(n13115), .Z(n13120) );
  OR U14190 ( .A(n13118), .B(n13117), .Z(n13119) );
  AND U14191 ( .A(n13120), .B(n13119), .Z(n13126) );
  XOR U14192 ( .A(n13127), .B(n13126), .Z(n13129) );
  XOR U14193 ( .A(n13128), .B(n13129), .Z(n13142) );
  XNOR U14194 ( .A(n13142), .B(sreg[1539]), .Z(n13144) );
  NANDN U14195 ( .A(n13121), .B(sreg[1538]), .Z(n13125) );
  NAND U14196 ( .A(n13123), .B(n13122), .Z(n13124) );
  NAND U14197 ( .A(n13125), .B(n13124), .Z(n13143) );
  XOR U14198 ( .A(n13144), .B(n13143), .Z(c[1539]) );
  NANDN U14199 ( .A(n13127), .B(n13126), .Z(n13131) );
  OR U14200 ( .A(n13129), .B(n13128), .Z(n13130) );
  AND U14201 ( .A(n13131), .B(n13130), .Z(n13149) );
  XOR U14202 ( .A(a[518]), .B(n2250), .Z(n13153) );
  AND U14203 ( .A(a[520]), .B(b[0]), .Z(n13133) );
  XNOR U14204 ( .A(n13133), .B(n2175), .Z(n13135) );
  NANDN U14205 ( .A(b[0]), .B(a[519]), .Z(n13134) );
  NAND U14206 ( .A(n13135), .B(n13134), .Z(n13158) );
  AND U14207 ( .A(a[516]), .B(b[3]), .Z(n13157) );
  XOR U14208 ( .A(n13158), .B(n13157), .Z(n13160) );
  XOR U14209 ( .A(n13159), .B(n13160), .Z(n13148) );
  NANDN U14210 ( .A(n13137), .B(n13136), .Z(n13141) );
  OR U14211 ( .A(n13139), .B(n13138), .Z(n13140) );
  AND U14212 ( .A(n13141), .B(n13140), .Z(n13147) );
  XOR U14213 ( .A(n13148), .B(n13147), .Z(n13150) );
  XOR U14214 ( .A(n13149), .B(n13150), .Z(n13163) );
  XNOR U14215 ( .A(n13163), .B(sreg[1540]), .Z(n13165) );
  NANDN U14216 ( .A(n13142), .B(sreg[1539]), .Z(n13146) );
  NAND U14217 ( .A(n13144), .B(n13143), .Z(n13145) );
  NAND U14218 ( .A(n13146), .B(n13145), .Z(n13164) );
  XOR U14219 ( .A(n13165), .B(n13164), .Z(c[1540]) );
  NANDN U14220 ( .A(n13148), .B(n13147), .Z(n13152) );
  OR U14221 ( .A(n13150), .B(n13149), .Z(n13151) );
  AND U14222 ( .A(n13152), .B(n13151), .Z(n13170) );
  XOR U14223 ( .A(a[519]), .B(n2250), .Z(n13174) );
  AND U14224 ( .A(a[517]), .B(b[3]), .Z(n13178) );
  AND U14225 ( .A(a[521]), .B(b[0]), .Z(n13154) );
  XNOR U14226 ( .A(n13154), .B(n2175), .Z(n13156) );
  NANDN U14227 ( .A(b[0]), .B(a[520]), .Z(n13155) );
  NAND U14228 ( .A(n13156), .B(n13155), .Z(n13179) );
  XOR U14229 ( .A(n13178), .B(n13179), .Z(n13181) );
  XOR U14230 ( .A(n13180), .B(n13181), .Z(n13169) );
  NANDN U14231 ( .A(n13158), .B(n13157), .Z(n13162) );
  OR U14232 ( .A(n13160), .B(n13159), .Z(n13161) );
  AND U14233 ( .A(n13162), .B(n13161), .Z(n13168) );
  XOR U14234 ( .A(n13169), .B(n13168), .Z(n13171) );
  XOR U14235 ( .A(n13170), .B(n13171), .Z(n13184) );
  XNOR U14236 ( .A(n13184), .B(sreg[1541]), .Z(n13186) );
  NANDN U14237 ( .A(n13163), .B(sreg[1540]), .Z(n13167) );
  NAND U14238 ( .A(n13165), .B(n13164), .Z(n13166) );
  NAND U14239 ( .A(n13167), .B(n13166), .Z(n13185) );
  XOR U14240 ( .A(n13186), .B(n13185), .Z(c[1541]) );
  NANDN U14241 ( .A(n13169), .B(n13168), .Z(n13173) );
  OR U14242 ( .A(n13171), .B(n13170), .Z(n13172) );
  AND U14243 ( .A(n13173), .B(n13172), .Z(n13191) );
  XOR U14244 ( .A(a[520]), .B(n2250), .Z(n13195) );
  AND U14245 ( .A(a[522]), .B(b[0]), .Z(n13175) );
  XNOR U14246 ( .A(n13175), .B(n2175), .Z(n13177) );
  NANDN U14247 ( .A(b[0]), .B(a[521]), .Z(n13176) );
  NAND U14248 ( .A(n13177), .B(n13176), .Z(n13200) );
  AND U14249 ( .A(a[518]), .B(b[3]), .Z(n13199) );
  XOR U14250 ( .A(n13200), .B(n13199), .Z(n13202) );
  XOR U14251 ( .A(n13201), .B(n13202), .Z(n13190) );
  NANDN U14252 ( .A(n13179), .B(n13178), .Z(n13183) );
  OR U14253 ( .A(n13181), .B(n13180), .Z(n13182) );
  AND U14254 ( .A(n13183), .B(n13182), .Z(n13189) );
  XOR U14255 ( .A(n13190), .B(n13189), .Z(n13192) );
  XOR U14256 ( .A(n13191), .B(n13192), .Z(n13205) );
  XNOR U14257 ( .A(n13205), .B(sreg[1542]), .Z(n13207) );
  NANDN U14258 ( .A(n13184), .B(sreg[1541]), .Z(n13188) );
  NAND U14259 ( .A(n13186), .B(n13185), .Z(n13187) );
  NAND U14260 ( .A(n13188), .B(n13187), .Z(n13206) );
  XOR U14261 ( .A(n13207), .B(n13206), .Z(c[1542]) );
  NANDN U14262 ( .A(n13190), .B(n13189), .Z(n13194) );
  OR U14263 ( .A(n13192), .B(n13191), .Z(n13193) );
  AND U14264 ( .A(n13194), .B(n13193), .Z(n13212) );
  XOR U14265 ( .A(a[521]), .B(n2250), .Z(n13216) );
  AND U14266 ( .A(a[519]), .B(b[3]), .Z(n13220) );
  AND U14267 ( .A(a[523]), .B(b[0]), .Z(n13196) );
  XNOR U14268 ( .A(n13196), .B(n2175), .Z(n13198) );
  NANDN U14269 ( .A(b[0]), .B(a[522]), .Z(n13197) );
  NAND U14270 ( .A(n13198), .B(n13197), .Z(n13221) );
  XOR U14271 ( .A(n13220), .B(n13221), .Z(n13223) );
  XOR U14272 ( .A(n13222), .B(n13223), .Z(n13211) );
  NANDN U14273 ( .A(n13200), .B(n13199), .Z(n13204) );
  OR U14274 ( .A(n13202), .B(n13201), .Z(n13203) );
  AND U14275 ( .A(n13204), .B(n13203), .Z(n13210) );
  XOR U14276 ( .A(n13211), .B(n13210), .Z(n13213) );
  XOR U14277 ( .A(n13212), .B(n13213), .Z(n13226) );
  XNOR U14278 ( .A(n13226), .B(sreg[1543]), .Z(n13228) );
  NANDN U14279 ( .A(n13205), .B(sreg[1542]), .Z(n13209) );
  NAND U14280 ( .A(n13207), .B(n13206), .Z(n13208) );
  NAND U14281 ( .A(n13209), .B(n13208), .Z(n13227) );
  XOR U14282 ( .A(n13228), .B(n13227), .Z(c[1543]) );
  NANDN U14283 ( .A(n13211), .B(n13210), .Z(n13215) );
  OR U14284 ( .A(n13213), .B(n13212), .Z(n13214) );
  AND U14285 ( .A(n13215), .B(n13214), .Z(n13233) );
  XOR U14286 ( .A(a[522]), .B(n2250), .Z(n13237) );
  AND U14287 ( .A(a[524]), .B(b[0]), .Z(n13217) );
  XNOR U14288 ( .A(n13217), .B(n2175), .Z(n13219) );
  NANDN U14289 ( .A(b[0]), .B(a[523]), .Z(n13218) );
  NAND U14290 ( .A(n13219), .B(n13218), .Z(n13242) );
  AND U14291 ( .A(a[520]), .B(b[3]), .Z(n13241) );
  XOR U14292 ( .A(n13242), .B(n13241), .Z(n13244) );
  XOR U14293 ( .A(n13243), .B(n13244), .Z(n13232) );
  NANDN U14294 ( .A(n13221), .B(n13220), .Z(n13225) );
  OR U14295 ( .A(n13223), .B(n13222), .Z(n13224) );
  AND U14296 ( .A(n13225), .B(n13224), .Z(n13231) );
  XOR U14297 ( .A(n13232), .B(n13231), .Z(n13234) );
  XOR U14298 ( .A(n13233), .B(n13234), .Z(n13247) );
  XNOR U14299 ( .A(n13247), .B(sreg[1544]), .Z(n13249) );
  NANDN U14300 ( .A(n13226), .B(sreg[1543]), .Z(n13230) );
  NAND U14301 ( .A(n13228), .B(n13227), .Z(n13229) );
  NAND U14302 ( .A(n13230), .B(n13229), .Z(n13248) );
  XOR U14303 ( .A(n13249), .B(n13248), .Z(c[1544]) );
  NANDN U14304 ( .A(n13232), .B(n13231), .Z(n13236) );
  OR U14305 ( .A(n13234), .B(n13233), .Z(n13235) );
  AND U14306 ( .A(n13236), .B(n13235), .Z(n13254) );
  XOR U14307 ( .A(a[523]), .B(n2250), .Z(n13258) );
  AND U14308 ( .A(a[525]), .B(b[0]), .Z(n13238) );
  XNOR U14309 ( .A(n13238), .B(n2175), .Z(n13240) );
  NANDN U14310 ( .A(b[0]), .B(a[524]), .Z(n13239) );
  NAND U14311 ( .A(n13240), .B(n13239), .Z(n13263) );
  AND U14312 ( .A(a[521]), .B(b[3]), .Z(n13262) );
  XOR U14313 ( .A(n13263), .B(n13262), .Z(n13265) );
  XOR U14314 ( .A(n13264), .B(n13265), .Z(n13253) );
  NANDN U14315 ( .A(n13242), .B(n13241), .Z(n13246) );
  OR U14316 ( .A(n13244), .B(n13243), .Z(n13245) );
  AND U14317 ( .A(n13246), .B(n13245), .Z(n13252) );
  XOR U14318 ( .A(n13253), .B(n13252), .Z(n13255) );
  XOR U14319 ( .A(n13254), .B(n13255), .Z(n13268) );
  XNOR U14320 ( .A(n13268), .B(sreg[1545]), .Z(n13270) );
  NANDN U14321 ( .A(n13247), .B(sreg[1544]), .Z(n13251) );
  NAND U14322 ( .A(n13249), .B(n13248), .Z(n13250) );
  NAND U14323 ( .A(n13251), .B(n13250), .Z(n13269) );
  XOR U14324 ( .A(n13270), .B(n13269), .Z(c[1545]) );
  NANDN U14325 ( .A(n13253), .B(n13252), .Z(n13257) );
  OR U14326 ( .A(n13255), .B(n13254), .Z(n13256) );
  AND U14327 ( .A(n13257), .B(n13256), .Z(n13275) );
  XOR U14328 ( .A(a[524]), .B(n2251), .Z(n13279) );
  AND U14329 ( .A(a[522]), .B(b[3]), .Z(n13283) );
  AND U14330 ( .A(a[526]), .B(b[0]), .Z(n13259) );
  XNOR U14331 ( .A(n13259), .B(n2175), .Z(n13261) );
  NANDN U14332 ( .A(b[0]), .B(a[525]), .Z(n13260) );
  NAND U14333 ( .A(n13261), .B(n13260), .Z(n13284) );
  XOR U14334 ( .A(n13283), .B(n13284), .Z(n13286) );
  XOR U14335 ( .A(n13285), .B(n13286), .Z(n13274) );
  NANDN U14336 ( .A(n13263), .B(n13262), .Z(n13267) );
  OR U14337 ( .A(n13265), .B(n13264), .Z(n13266) );
  AND U14338 ( .A(n13267), .B(n13266), .Z(n13273) );
  XOR U14339 ( .A(n13274), .B(n13273), .Z(n13276) );
  XOR U14340 ( .A(n13275), .B(n13276), .Z(n13289) );
  XNOR U14341 ( .A(n13289), .B(sreg[1546]), .Z(n13291) );
  NANDN U14342 ( .A(n13268), .B(sreg[1545]), .Z(n13272) );
  NAND U14343 ( .A(n13270), .B(n13269), .Z(n13271) );
  NAND U14344 ( .A(n13272), .B(n13271), .Z(n13290) );
  XOR U14345 ( .A(n13291), .B(n13290), .Z(c[1546]) );
  NANDN U14346 ( .A(n13274), .B(n13273), .Z(n13278) );
  OR U14347 ( .A(n13276), .B(n13275), .Z(n13277) );
  AND U14348 ( .A(n13278), .B(n13277), .Z(n13296) );
  XOR U14349 ( .A(a[525]), .B(n2251), .Z(n13300) );
  AND U14350 ( .A(a[527]), .B(b[0]), .Z(n13280) );
  XNOR U14351 ( .A(n13280), .B(n2175), .Z(n13282) );
  NANDN U14352 ( .A(b[0]), .B(a[526]), .Z(n13281) );
  NAND U14353 ( .A(n13282), .B(n13281), .Z(n13305) );
  AND U14354 ( .A(a[523]), .B(b[3]), .Z(n13304) );
  XOR U14355 ( .A(n13305), .B(n13304), .Z(n13307) );
  XOR U14356 ( .A(n13306), .B(n13307), .Z(n13295) );
  NANDN U14357 ( .A(n13284), .B(n13283), .Z(n13288) );
  OR U14358 ( .A(n13286), .B(n13285), .Z(n13287) );
  AND U14359 ( .A(n13288), .B(n13287), .Z(n13294) );
  XOR U14360 ( .A(n13295), .B(n13294), .Z(n13297) );
  XOR U14361 ( .A(n13296), .B(n13297), .Z(n13310) );
  XNOR U14362 ( .A(n13310), .B(sreg[1547]), .Z(n13312) );
  NANDN U14363 ( .A(n13289), .B(sreg[1546]), .Z(n13293) );
  NAND U14364 ( .A(n13291), .B(n13290), .Z(n13292) );
  NAND U14365 ( .A(n13293), .B(n13292), .Z(n13311) );
  XOR U14366 ( .A(n13312), .B(n13311), .Z(c[1547]) );
  NANDN U14367 ( .A(n13295), .B(n13294), .Z(n13299) );
  OR U14368 ( .A(n13297), .B(n13296), .Z(n13298) );
  AND U14369 ( .A(n13299), .B(n13298), .Z(n13317) );
  XOR U14370 ( .A(a[526]), .B(n2251), .Z(n13321) );
  AND U14371 ( .A(a[528]), .B(b[0]), .Z(n13301) );
  XNOR U14372 ( .A(n13301), .B(n2175), .Z(n13303) );
  NANDN U14373 ( .A(b[0]), .B(a[527]), .Z(n13302) );
  NAND U14374 ( .A(n13303), .B(n13302), .Z(n13326) );
  AND U14375 ( .A(a[524]), .B(b[3]), .Z(n13325) );
  XOR U14376 ( .A(n13326), .B(n13325), .Z(n13328) );
  XOR U14377 ( .A(n13327), .B(n13328), .Z(n13316) );
  NANDN U14378 ( .A(n13305), .B(n13304), .Z(n13309) );
  OR U14379 ( .A(n13307), .B(n13306), .Z(n13308) );
  AND U14380 ( .A(n13309), .B(n13308), .Z(n13315) );
  XOR U14381 ( .A(n13316), .B(n13315), .Z(n13318) );
  XOR U14382 ( .A(n13317), .B(n13318), .Z(n13331) );
  XNOR U14383 ( .A(n13331), .B(sreg[1548]), .Z(n13333) );
  NANDN U14384 ( .A(n13310), .B(sreg[1547]), .Z(n13314) );
  NAND U14385 ( .A(n13312), .B(n13311), .Z(n13313) );
  NAND U14386 ( .A(n13314), .B(n13313), .Z(n13332) );
  XOR U14387 ( .A(n13333), .B(n13332), .Z(c[1548]) );
  NANDN U14388 ( .A(n13316), .B(n13315), .Z(n13320) );
  OR U14389 ( .A(n13318), .B(n13317), .Z(n13319) );
  AND U14390 ( .A(n13320), .B(n13319), .Z(n13338) );
  XOR U14391 ( .A(a[527]), .B(n2251), .Z(n13342) );
  AND U14392 ( .A(a[529]), .B(b[0]), .Z(n13322) );
  XNOR U14393 ( .A(n13322), .B(n2175), .Z(n13324) );
  NANDN U14394 ( .A(b[0]), .B(a[528]), .Z(n13323) );
  NAND U14395 ( .A(n13324), .B(n13323), .Z(n13347) );
  AND U14396 ( .A(a[525]), .B(b[3]), .Z(n13346) );
  XOR U14397 ( .A(n13347), .B(n13346), .Z(n13349) );
  XOR U14398 ( .A(n13348), .B(n13349), .Z(n13337) );
  NANDN U14399 ( .A(n13326), .B(n13325), .Z(n13330) );
  OR U14400 ( .A(n13328), .B(n13327), .Z(n13329) );
  AND U14401 ( .A(n13330), .B(n13329), .Z(n13336) );
  XOR U14402 ( .A(n13337), .B(n13336), .Z(n13339) );
  XOR U14403 ( .A(n13338), .B(n13339), .Z(n13352) );
  XNOR U14404 ( .A(n13352), .B(sreg[1549]), .Z(n13354) );
  NANDN U14405 ( .A(n13331), .B(sreg[1548]), .Z(n13335) );
  NAND U14406 ( .A(n13333), .B(n13332), .Z(n13334) );
  NAND U14407 ( .A(n13335), .B(n13334), .Z(n13353) );
  XOR U14408 ( .A(n13354), .B(n13353), .Z(c[1549]) );
  NANDN U14409 ( .A(n13337), .B(n13336), .Z(n13341) );
  OR U14410 ( .A(n13339), .B(n13338), .Z(n13340) );
  AND U14411 ( .A(n13341), .B(n13340), .Z(n13359) );
  XOR U14412 ( .A(a[528]), .B(n2251), .Z(n13363) );
  AND U14413 ( .A(a[530]), .B(b[0]), .Z(n13343) );
  XNOR U14414 ( .A(n13343), .B(n2175), .Z(n13345) );
  NANDN U14415 ( .A(b[0]), .B(a[529]), .Z(n13344) );
  NAND U14416 ( .A(n13345), .B(n13344), .Z(n13368) );
  AND U14417 ( .A(a[526]), .B(b[3]), .Z(n13367) );
  XOR U14418 ( .A(n13368), .B(n13367), .Z(n13370) );
  XOR U14419 ( .A(n13369), .B(n13370), .Z(n13358) );
  NANDN U14420 ( .A(n13347), .B(n13346), .Z(n13351) );
  OR U14421 ( .A(n13349), .B(n13348), .Z(n13350) );
  AND U14422 ( .A(n13351), .B(n13350), .Z(n13357) );
  XOR U14423 ( .A(n13358), .B(n13357), .Z(n13360) );
  XOR U14424 ( .A(n13359), .B(n13360), .Z(n13373) );
  XNOR U14425 ( .A(n13373), .B(sreg[1550]), .Z(n13375) );
  NANDN U14426 ( .A(n13352), .B(sreg[1549]), .Z(n13356) );
  NAND U14427 ( .A(n13354), .B(n13353), .Z(n13355) );
  NAND U14428 ( .A(n13356), .B(n13355), .Z(n13374) );
  XOR U14429 ( .A(n13375), .B(n13374), .Z(c[1550]) );
  NANDN U14430 ( .A(n13358), .B(n13357), .Z(n13362) );
  OR U14431 ( .A(n13360), .B(n13359), .Z(n13361) );
  AND U14432 ( .A(n13362), .B(n13361), .Z(n13380) );
  XOR U14433 ( .A(a[529]), .B(n2251), .Z(n13384) );
  AND U14434 ( .A(a[531]), .B(b[0]), .Z(n13364) );
  XNOR U14435 ( .A(n13364), .B(n2175), .Z(n13366) );
  NANDN U14436 ( .A(b[0]), .B(a[530]), .Z(n13365) );
  NAND U14437 ( .A(n13366), .B(n13365), .Z(n13389) );
  AND U14438 ( .A(a[527]), .B(b[3]), .Z(n13388) );
  XOR U14439 ( .A(n13389), .B(n13388), .Z(n13391) );
  XOR U14440 ( .A(n13390), .B(n13391), .Z(n13379) );
  NANDN U14441 ( .A(n13368), .B(n13367), .Z(n13372) );
  OR U14442 ( .A(n13370), .B(n13369), .Z(n13371) );
  AND U14443 ( .A(n13372), .B(n13371), .Z(n13378) );
  XOR U14444 ( .A(n13379), .B(n13378), .Z(n13381) );
  XOR U14445 ( .A(n13380), .B(n13381), .Z(n13394) );
  XNOR U14446 ( .A(n13394), .B(sreg[1551]), .Z(n13396) );
  NANDN U14447 ( .A(n13373), .B(sreg[1550]), .Z(n13377) );
  NAND U14448 ( .A(n13375), .B(n13374), .Z(n13376) );
  NAND U14449 ( .A(n13377), .B(n13376), .Z(n13395) );
  XOR U14450 ( .A(n13396), .B(n13395), .Z(c[1551]) );
  NANDN U14451 ( .A(n13379), .B(n13378), .Z(n13383) );
  OR U14452 ( .A(n13381), .B(n13380), .Z(n13382) );
  AND U14453 ( .A(n13383), .B(n13382), .Z(n13401) );
  XOR U14454 ( .A(a[530]), .B(n2251), .Z(n13405) );
  AND U14455 ( .A(a[532]), .B(b[0]), .Z(n13385) );
  XNOR U14456 ( .A(n13385), .B(n2175), .Z(n13387) );
  NANDN U14457 ( .A(b[0]), .B(a[531]), .Z(n13386) );
  NAND U14458 ( .A(n13387), .B(n13386), .Z(n13410) );
  AND U14459 ( .A(a[528]), .B(b[3]), .Z(n13409) );
  XOR U14460 ( .A(n13410), .B(n13409), .Z(n13412) );
  XOR U14461 ( .A(n13411), .B(n13412), .Z(n13400) );
  NANDN U14462 ( .A(n13389), .B(n13388), .Z(n13393) );
  OR U14463 ( .A(n13391), .B(n13390), .Z(n13392) );
  AND U14464 ( .A(n13393), .B(n13392), .Z(n13399) );
  XOR U14465 ( .A(n13400), .B(n13399), .Z(n13402) );
  XOR U14466 ( .A(n13401), .B(n13402), .Z(n13415) );
  XNOR U14467 ( .A(n13415), .B(sreg[1552]), .Z(n13417) );
  NANDN U14468 ( .A(n13394), .B(sreg[1551]), .Z(n13398) );
  NAND U14469 ( .A(n13396), .B(n13395), .Z(n13397) );
  NAND U14470 ( .A(n13398), .B(n13397), .Z(n13416) );
  XOR U14471 ( .A(n13417), .B(n13416), .Z(c[1552]) );
  NANDN U14472 ( .A(n13400), .B(n13399), .Z(n13404) );
  OR U14473 ( .A(n13402), .B(n13401), .Z(n13403) );
  AND U14474 ( .A(n13404), .B(n13403), .Z(n13422) );
  XOR U14475 ( .A(a[531]), .B(n2252), .Z(n13426) );
  AND U14476 ( .A(a[533]), .B(b[0]), .Z(n13406) );
  XNOR U14477 ( .A(n13406), .B(n2175), .Z(n13408) );
  NANDN U14478 ( .A(b[0]), .B(a[532]), .Z(n13407) );
  NAND U14479 ( .A(n13408), .B(n13407), .Z(n13431) );
  AND U14480 ( .A(a[529]), .B(b[3]), .Z(n13430) );
  XOR U14481 ( .A(n13431), .B(n13430), .Z(n13433) );
  XOR U14482 ( .A(n13432), .B(n13433), .Z(n13421) );
  NANDN U14483 ( .A(n13410), .B(n13409), .Z(n13414) );
  OR U14484 ( .A(n13412), .B(n13411), .Z(n13413) );
  AND U14485 ( .A(n13414), .B(n13413), .Z(n13420) );
  XOR U14486 ( .A(n13421), .B(n13420), .Z(n13423) );
  XOR U14487 ( .A(n13422), .B(n13423), .Z(n13436) );
  XNOR U14488 ( .A(n13436), .B(sreg[1553]), .Z(n13438) );
  NANDN U14489 ( .A(n13415), .B(sreg[1552]), .Z(n13419) );
  NAND U14490 ( .A(n13417), .B(n13416), .Z(n13418) );
  NAND U14491 ( .A(n13419), .B(n13418), .Z(n13437) );
  XOR U14492 ( .A(n13438), .B(n13437), .Z(c[1553]) );
  NANDN U14493 ( .A(n13421), .B(n13420), .Z(n13425) );
  OR U14494 ( .A(n13423), .B(n13422), .Z(n13424) );
  AND U14495 ( .A(n13425), .B(n13424), .Z(n13443) );
  XOR U14496 ( .A(a[532]), .B(n2252), .Z(n13447) );
  AND U14497 ( .A(a[534]), .B(b[0]), .Z(n13427) );
  XNOR U14498 ( .A(n13427), .B(n2175), .Z(n13429) );
  NANDN U14499 ( .A(b[0]), .B(a[533]), .Z(n13428) );
  NAND U14500 ( .A(n13429), .B(n13428), .Z(n13452) );
  AND U14501 ( .A(a[530]), .B(b[3]), .Z(n13451) );
  XOR U14502 ( .A(n13452), .B(n13451), .Z(n13454) );
  XOR U14503 ( .A(n13453), .B(n13454), .Z(n13442) );
  NANDN U14504 ( .A(n13431), .B(n13430), .Z(n13435) );
  OR U14505 ( .A(n13433), .B(n13432), .Z(n13434) );
  AND U14506 ( .A(n13435), .B(n13434), .Z(n13441) );
  XOR U14507 ( .A(n13442), .B(n13441), .Z(n13444) );
  XOR U14508 ( .A(n13443), .B(n13444), .Z(n13457) );
  XNOR U14509 ( .A(n13457), .B(sreg[1554]), .Z(n13459) );
  NANDN U14510 ( .A(n13436), .B(sreg[1553]), .Z(n13440) );
  NAND U14511 ( .A(n13438), .B(n13437), .Z(n13439) );
  NAND U14512 ( .A(n13440), .B(n13439), .Z(n13458) );
  XOR U14513 ( .A(n13459), .B(n13458), .Z(c[1554]) );
  NANDN U14514 ( .A(n13442), .B(n13441), .Z(n13446) );
  OR U14515 ( .A(n13444), .B(n13443), .Z(n13445) );
  AND U14516 ( .A(n13446), .B(n13445), .Z(n13464) );
  XOR U14517 ( .A(a[533]), .B(n2252), .Z(n13468) );
  AND U14518 ( .A(a[535]), .B(b[0]), .Z(n13448) );
  XNOR U14519 ( .A(n13448), .B(n2175), .Z(n13450) );
  NANDN U14520 ( .A(b[0]), .B(a[534]), .Z(n13449) );
  NAND U14521 ( .A(n13450), .B(n13449), .Z(n13473) );
  AND U14522 ( .A(a[531]), .B(b[3]), .Z(n13472) );
  XOR U14523 ( .A(n13473), .B(n13472), .Z(n13475) );
  XOR U14524 ( .A(n13474), .B(n13475), .Z(n13463) );
  NANDN U14525 ( .A(n13452), .B(n13451), .Z(n13456) );
  OR U14526 ( .A(n13454), .B(n13453), .Z(n13455) );
  AND U14527 ( .A(n13456), .B(n13455), .Z(n13462) );
  XOR U14528 ( .A(n13463), .B(n13462), .Z(n13465) );
  XOR U14529 ( .A(n13464), .B(n13465), .Z(n13478) );
  XNOR U14530 ( .A(n13478), .B(sreg[1555]), .Z(n13480) );
  NANDN U14531 ( .A(n13457), .B(sreg[1554]), .Z(n13461) );
  NAND U14532 ( .A(n13459), .B(n13458), .Z(n13460) );
  NAND U14533 ( .A(n13461), .B(n13460), .Z(n13479) );
  XOR U14534 ( .A(n13480), .B(n13479), .Z(c[1555]) );
  NANDN U14535 ( .A(n13463), .B(n13462), .Z(n13467) );
  OR U14536 ( .A(n13465), .B(n13464), .Z(n13466) );
  AND U14537 ( .A(n13467), .B(n13466), .Z(n13485) );
  XOR U14538 ( .A(a[534]), .B(n2252), .Z(n13489) );
  AND U14539 ( .A(a[532]), .B(b[3]), .Z(n13493) );
  AND U14540 ( .A(a[536]), .B(b[0]), .Z(n13469) );
  XNOR U14541 ( .A(n13469), .B(n2175), .Z(n13471) );
  NANDN U14542 ( .A(b[0]), .B(a[535]), .Z(n13470) );
  NAND U14543 ( .A(n13471), .B(n13470), .Z(n13494) );
  XOR U14544 ( .A(n13493), .B(n13494), .Z(n13496) );
  XOR U14545 ( .A(n13495), .B(n13496), .Z(n13484) );
  NANDN U14546 ( .A(n13473), .B(n13472), .Z(n13477) );
  OR U14547 ( .A(n13475), .B(n13474), .Z(n13476) );
  AND U14548 ( .A(n13477), .B(n13476), .Z(n13483) );
  XOR U14549 ( .A(n13484), .B(n13483), .Z(n13486) );
  XOR U14550 ( .A(n13485), .B(n13486), .Z(n13499) );
  XNOR U14551 ( .A(n13499), .B(sreg[1556]), .Z(n13501) );
  NANDN U14552 ( .A(n13478), .B(sreg[1555]), .Z(n13482) );
  NAND U14553 ( .A(n13480), .B(n13479), .Z(n13481) );
  NAND U14554 ( .A(n13482), .B(n13481), .Z(n13500) );
  XOR U14555 ( .A(n13501), .B(n13500), .Z(c[1556]) );
  NANDN U14556 ( .A(n13484), .B(n13483), .Z(n13488) );
  OR U14557 ( .A(n13486), .B(n13485), .Z(n13487) );
  AND U14558 ( .A(n13488), .B(n13487), .Z(n13506) );
  XOR U14559 ( .A(a[535]), .B(n2252), .Z(n13510) );
  AND U14560 ( .A(a[537]), .B(b[0]), .Z(n13490) );
  XNOR U14561 ( .A(n13490), .B(n2175), .Z(n13492) );
  NANDN U14562 ( .A(b[0]), .B(a[536]), .Z(n13491) );
  NAND U14563 ( .A(n13492), .B(n13491), .Z(n13515) );
  AND U14564 ( .A(a[533]), .B(b[3]), .Z(n13514) );
  XOR U14565 ( .A(n13515), .B(n13514), .Z(n13517) );
  XOR U14566 ( .A(n13516), .B(n13517), .Z(n13505) );
  NANDN U14567 ( .A(n13494), .B(n13493), .Z(n13498) );
  OR U14568 ( .A(n13496), .B(n13495), .Z(n13497) );
  AND U14569 ( .A(n13498), .B(n13497), .Z(n13504) );
  XOR U14570 ( .A(n13505), .B(n13504), .Z(n13507) );
  XOR U14571 ( .A(n13506), .B(n13507), .Z(n13520) );
  XNOR U14572 ( .A(n13520), .B(sreg[1557]), .Z(n13522) );
  NANDN U14573 ( .A(n13499), .B(sreg[1556]), .Z(n13503) );
  NAND U14574 ( .A(n13501), .B(n13500), .Z(n13502) );
  NAND U14575 ( .A(n13503), .B(n13502), .Z(n13521) );
  XOR U14576 ( .A(n13522), .B(n13521), .Z(c[1557]) );
  NANDN U14577 ( .A(n13505), .B(n13504), .Z(n13509) );
  OR U14578 ( .A(n13507), .B(n13506), .Z(n13508) );
  AND U14579 ( .A(n13509), .B(n13508), .Z(n13527) );
  XOR U14580 ( .A(a[536]), .B(n2252), .Z(n13531) );
  AND U14581 ( .A(a[534]), .B(b[3]), .Z(n13535) );
  AND U14582 ( .A(a[538]), .B(b[0]), .Z(n13511) );
  XNOR U14583 ( .A(n13511), .B(n2175), .Z(n13513) );
  NANDN U14584 ( .A(b[0]), .B(a[537]), .Z(n13512) );
  NAND U14585 ( .A(n13513), .B(n13512), .Z(n13536) );
  XOR U14586 ( .A(n13535), .B(n13536), .Z(n13538) );
  XOR U14587 ( .A(n13537), .B(n13538), .Z(n13526) );
  NANDN U14588 ( .A(n13515), .B(n13514), .Z(n13519) );
  OR U14589 ( .A(n13517), .B(n13516), .Z(n13518) );
  AND U14590 ( .A(n13519), .B(n13518), .Z(n13525) );
  XOR U14591 ( .A(n13526), .B(n13525), .Z(n13528) );
  XOR U14592 ( .A(n13527), .B(n13528), .Z(n13541) );
  XNOR U14593 ( .A(n13541), .B(sreg[1558]), .Z(n13543) );
  NANDN U14594 ( .A(n13520), .B(sreg[1557]), .Z(n13524) );
  NAND U14595 ( .A(n13522), .B(n13521), .Z(n13523) );
  NAND U14596 ( .A(n13524), .B(n13523), .Z(n13542) );
  XOR U14597 ( .A(n13543), .B(n13542), .Z(c[1558]) );
  NANDN U14598 ( .A(n13526), .B(n13525), .Z(n13530) );
  OR U14599 ( .A(n13528), .B(n13527), .Z(n13529) );
  AND U14600 ( .A(n13530), .B(n13529), .Z(n13548) );
  XOR U14601 ( .A(a[537]), .B(n2252), .Z(n13552) );
  AND U14602 ( .A(a[539]), .B(b[0]), .Z(n13532) );
  XNOR U14603 ( .A(n13532), .B(n2175), .Z(n13534) );
  NANDN U14604 ( .A(b[0]), .B(a[538]), .Z(n13533) );
  NAND U14605 ( .A(n13534), .B(n13533), .Z(n13557) );
  AND U14606 ( .A(a[535]), .B(b[3]), .Z(n13556) );
  XOR U14607 ( .A(n13557), .B(n13556), .Z(n13559) );
  XOR U14608 ( .A(n13558), .B(n13559), .Z(n13547) );
  NANDN U14609 ( .A(n13536), .B(n13535), .Z(n13540) );
  OR U14610 ( .A(n13538), .B(n13537), .Z(n13539) );
  AND U14611 ( .A(n13540), .B(n13539), .Z(n13546) );
  XOR U14612 ( .A(n13547), .B(n13546), .Z(n13549) );
  XOR U14613 ( .A(n13548), .B(n13549), .Z(n13562) );
  XNOR U14614 ( .A(n13562), .B(sreg[1559]), .Z(n13564) );
  NANDN U14615 ( .A(n13541), .B(sreg[1558]), .Z(n13545) );
  NAND U14616 ( .A(n13543), .B(n13542), .Z(n13544) );
  NAND U14617 ( .A(n13545), .B(n13544), .Z(n13563) );
  XOR U14618 ( .A(n13564), .B(n13563), .Z(c[1559]) );
  NANDN U14619 ( .A(n13547), .B(n13546), .Z(n13551) );
  OR U14620 ( .A(n13549), .B(n13548), .Z(n13550) );
  AND U14621 ( .A(n13551), .B(n13550), .Z(n13569) );
  XOR U14622 ( .A(a[538]), .B(n2253), .Z(n13573) );
  AND U14623 ( .A(a[540]), .B(b[0]), .Z(n13553) );
  XNOR U14624 ( .A(n13553), .B(n2175), .Z(n13555) );
  NANDN U14625 ( .A(b[0]), .B(a[539]), .Z(n13554) );
  NAND U14626 ( .A(n13555), .B(n13554), .Z(n13578) );
  AND U14627 ( .A(a[536]), .B(b[3]), .Z(n13577) );
  XOR U14628 ( .A(n13578), .B(n13577), .Z(n13580) );
  XOR U14629 ( .A(n13579), .B(n13580), .Z(n13568) );
  NANDN U14630 ( .A(n13557), .B(n13556), .Z(n13561) );
  OR U14631 ( .A(n13559), .B(n13558), .Z(n13560) );
  AND U14632 ( .A(n13561), .B(n13560), .Z(n13567) );
  XOR U14633 ( .A(n13568), .B(n13567), .Z(n13570) );
  XOR U14634 ( .A(n13569), .B(n13570), .Z(n13583) );
  XNOR U14635 ( .A(n13583), .B(sreg[1560]), .Z(n13585) );
  NANDN U14636 ( .A(n13562), .B(sreg[1559]), .Z(n13566) );
  NAND U14637 ( .A(n13564), .B(n13563), .Z(n13565) );
  NAND U14638 ( .A(n13566), .B(n13565), .Z(n13584) );
  XOR U14639 ( .A(n13585), .B(n13584), .Z(c[1560]) );
  NANDN U14640 ( .A(n13568), .B(n13567), .Z(n13572) );
  OR U14641 ( .A(n13570), .B(n13569), .Z(n13571) );
  AND U14642 ( .A(n13572), .B(n13571), .Z(n13590) );
  XOR U14643 ( .A(a[539]), .B(n2253), .Z(n13594) );
  AND U14644 ( .A(a[541]), .B(b[0]), .Z(n13574) );
  XNOR U14645 ( .A(n13574), .B(n2175), .Z(n13576) );
  NANDN U14646 ( .A(b[0]), .B(a[540]), .Z(n13575) );
  NAND U14647 ( .A(n13576), .B(n13575), .Z(n13599) );
  AND U14648 ( .A(a[537]), .B(b[3]), .Z(n13598) );
  XOR U14649 ( .A(n13599), .B(n13598), .Z(n13601) );
  XOR U14650 ( .A(n13600), .B(n13601), .Z(n13589) );
  NANDN U14651 ( .A(n13578), .B(n13577), .Z(n13582) );
  OR U14652 ( .A(n13580), .B(n13579), .Z(n13581) );
  AND U14653 ( .A(n13582), .B(n13581), .Z(n13588) );
  XOR U14654 ( .A(n13589), .B(n13588), .Z(n13591) );
  XOR U14655 ( .A(n13590), .B(n13591), .Z(n13604) );
  XNOR U14656 ( .A(n13604), .B(sreg[1561]), .Z(n13606) );
  NANDN U14657 ( .A(n13583), .B(sreg[1560]), .Z(n13587) );
  NAND U14658 ( .A(n13585), .B(n13584), .Z(n13586) );
  NAND U14659 ( .A(n13587), .B(n13586), .Z(n13605) );
  XOR U14660 ( .A(n13606), .B(n13605), .Z(c[1561]) );
  NANDN U14661 ( .A(n13589), .B(n13588), .Z(n13593) );
  OR U14662 ( .A(n13591), .B(n13590), .Z(n13592) );
  AND U14663 ( .A(n13593), .B(n13592), .Z(n13611) );
  XOR U14664 ( .A(a[540]), .B(n2253), .Z(n13615) );
  AND U14665 ( .A(a[542]), .B(b[0]), .Z(n13595) );
  XNOR U14666 ( .A(n13595), .B(n2175), .Z(n13597) );
  NANDN U14667 ( .A(b[0]), .B(a[541]), .Z(n13596) );
  NAND U14668 ( .A(n13597), .B(n13596), .Z(n13620) );
  AND U14669 ( .A(a[538]), .B(b[3]), .Z(n13619) );
  XOR U14670 ( .A(n13620), .B(n13619), .Z(n13622) );
  XOR U14671 ( .A(n13621), .B(n13622), .Z(n13610) );
  NANDN U14672 ( .A(n13599), .B(n13598), .Z(n13603) );
  OR U14673 ( .A(n13601), .B(n13600), .Z(n13602) );
  AND U14674 ( .A(n13603), .B(n13602), .Z(n13609) );
  XOR U14675 ( .A(n13610), .B(n13609), .Z(n13612) );
  XOR U14676 ( .A(n13611), .B(n13612), .Z(n13625) );
  XNOR U14677 ( .A(n13625), .B(sreg[1562]), .Z(n13627) );
  NANDN U14678 ( .A(n13604), .B(sreg[1561]), .Z(n13608) );
  NAND U14679 ( .A(n13606), .B(n13605), .Z(n13607) );
  NAND U14680 ( .A(n13608), .B(n13607), .Z(n13626) );
  XOR U14681 ( .A(n13627), .B(n13626), .Z(c[1562]) );
  NANDN U14682 ( .A(n13610), .B(n13609), .Z(n13614) );
  OR U14683 ( .A(n13612), .B(n13611), .Z(n13613) );
  AND U14684 ( .A(n13614), .B(n13613), .Z(n13632) );
  XOR U14685 ( .A(a[541]), .B(n2253), .Z(n13636) );
  AND U14686 ( .A(a[543]), .B(b[0]), .Z(n13616) );
  XNOR U14687 ( .A(n13616), .B(n2175), .Z(n13618) );
  NANDN U14688 ( .A(b[0]), .B(a[542]), .Z(n13617) );
  NAND U14689 ( .A(n13618), .B(n13617), .Z(n13641) );
  AND U14690 ( .A(a[539]), .B(b[3]), .Z(n13640) );
  XOR U14691 ( .A(n13641), .B(n13640), .Z(n13643) );
  XOR U14692 ( .A(n13642), .B(n13643), .Z(n13631) );
  NANDN U14693 ( .A(n13620), .B(n13619), .Z(n13624) );
  OR U14694 ( .A(n13622), .B(n13621), .Z(n13623) );
  AND U14695 ( .A(n13624), .B(n13623), .Z(n13630) );
  XOR U14696 ( .A(n13631), .B(n13630), .Z(n13633) );
  XOR U14697 ( .A(n13632), .B(n13633), .Z(n13646) );
  XNOR U14698 ( .A(n13646), .B(sreg[1563]), .Z(n13648) );
  NANDN U14699 ( .A(n13625), .B(sreg[1562]), .Z(n13629) );
  NAND U14700 ( .A(n13627), .B(n13626), .Z(n13628) );
  NAND U14701 ( .A(n13629), .B(n13628), .Z(n13647) );
  XOR U14702 ( .A(n13648), .B(n13647), .Z(c[1563]) );
  NANDN U14703 ( .A(n13631), .B(n13630), .Z(n13635) );
  OR U14704 ( .A(n13633), .B(n13632), .Z(n13634) );
  AND U14705 ( .A(n13635), .B(n13634), .Z(n13653) );
  XOR U14706 ( .A(a[542]), .B(n2253), .Z(n13657) );
  AND U14707 ( .A(a[544]), .B(b[0]), .Z(n13637) );
  XNOR U14708 ( .A(n13637), .B(n2175), .Z(n13639) );
  NANDN U14709 ( .A(b[0]), .B(a[543]), .Z(n13638) );
  NAND U14710 ( .A(n13639), .B(n13638), .Z(n13662) );
  AND U14711 ( .A(a[540]), .B(b[3]), .Z(n13661) );
  XOR U14712 ( .A(n13662), .B(n13661), .Z(n13664) );
  XOR U14713 ( .A(n13663), .B(n13664), .Z(n13652) );
  NANDN U14714 ( .A(n13641), .B(n13640), .Z(n13645) );
  OR U14715 ( .A(n13643), .B(n13642), .Z(n13644) );
  AND U14716 ( .A(n13645), .B(n13644), .Z(n13651) );
  XOR U14717 ( .A(n13652), .B(n13651), .Z(n13654) );
  XOR U14718 ( .A(n13653), .B(n13654), .Z(n13667) );
  XNOR U14719 ( .A(n13667), .B(sreg[1564]), .Z(n13669) );
  NANDN U14720 ( .A(n13646), .B(sreg[1563]), .Z(n13650) );
  NAND U14721 ( .A(n13648), .B(n13647), .Z(n13649) );
  NAND U14722 ( .A(n13650), .B(n13649), .Z(n13668) );
  XOR U14723 ( .A(n13669), .B(n13668), .Z(c[1564]) );
  NANDN U14724 ( .A(n13652), .B(n13651), .Z(n13656) );
  OR U14725 ( .A(n13654), .B(n13653), .Z(n13655) );
  AND U14726 ( .A(n13656), .B(n13655), .Z(n13674) );
  XOR U14727 ( .A(a[543]), .B(n2253), .Z(n13678) );
  AND U14728 ( .A(a[541]), .B(b[3]), .Z(n13682) );
  AND U14729 ( .A(a[545]), .B(b[0]), .Z(n13658) );
  XNOR U14730 ( .A(n13658), .B(n2175), .Z(n13660) );
  NANDN U14731 ( .A(b[0]), .B(a[544]), .Z(n13659) );
  NAND U14732 ( .A(n13660), .B(n13659), .Z(n13683) );
  XOR U14733 ( .A(n13682), .B(n13683), .Z(n13685) );
  XOR U14734 ( .A(n13684), .B(n13685), .Z(n13673) );
  NANDN U14735 ( .A(n13662), .B(n13661), .Z(n13666) );
  OR U14736 ( .A(n13664), .B(n13663), .Z(n13665) );
  AND U14737 ( .A(n13666), .B(n13665), .Z(n13672) );
  XOR U14738 ( .A(n13673), .B(n13672), .Z(n13675) );
  XOR U14739 ( .A(n13674), .B(n13675), .Z(n13688) );
  XNOR U14740 ( .A(n13688), .B(sreg[1565]), .Z(n13690) );
  NANDN U14741 ( .A(n13667), .B(sreg[1564]), .Z(n13671) );
  NAND U14742 ( .A(n13669), .B(n13668), .Z(n13670) );
  NAND U14743 ( .A(n13671), .B(n13670), .Z(n13689) );
  XOR U14744 ( .A(n13690), .B(n13689), .Z(c[1565]) );
  NANDN U14745 ( .A(n13673), .B(n13672), .Z(n13677) );
  OR U14746 ( .A(n13675), .B(n13674), .Z(n13676) );
  AND U14747 ( .A(n13677), .B(n13676), .Z(n13695) );
  XOR U14748 ( .A(a[544]), .B(n2253), .Z(n13699) );
  AND U14749 ( .A(a[546]), .B(b[0]), .Z(n13679) );
  XNOR U14750 ( .A(n13679), .B(n2175), .Z(n13681) );
  NANDN U14751 ( .A(b[0]), .B(a[545]), .Z(n13680) );
  NAND U14752 ( .A(n13681), .B(n13680), .Z(n13704) );
  AND U14753 ( .A(a[542]), .B(b[3]), .Z(n13703) );
  XOR U14754 ( .A(n13704), .B(n13703), .Z(n13706) );
  XOR U14755 ( .A(n13705), .B(n13706), .Z(n13694) );
  NANDN U14756 ( .A(n13683), .B(n13682), .Z(n13687) );
  OR U14757 ( .A(n13685), .B(n13684), .Z(n13686) );
  AND U14758 ( .A(n13687), .B(n13686), .Z(n13693) );
  XOR U14759 ( .A(n13694), .B(n13693), .Z(n13696) );
  XOR U14760 ( .A(n13695), .B(n13696), .Z(n13709) );
  XNOR U14761 ( .A(n13709), .B(sreg[1566]), .Z(n13711) );
  NANDN U14762 ( .A(n13688), .B(sreg[1565]), .Z(n13692) );
  NAND U14763 ( .A(n13690), .B(n13689), .Z(n13691) );
  NAND U14764 ( .A(n13692), .B(n13691), .Z(n13710) );
  XOR U14765 ( .A(n13711), .B(n13710), .Z(c[1566]) );
  NANDN U14766 ( .A(n13694), .B(n13693), .Z(n13698) );
  OR U14767 ( .A(n13696), .B(n13695), .Z(n13697) );
  AND U14768 ( .A(n13698), .B(n13697), .Z(n13716) );
  XOR U14769 ( .A(a[545]), .B(n2254), .Z(n13720) );
  AND U14770 ( .A(a[543]), .B(b[3]), .Z(n13724) );
  AND U14771 ( .A(a[547]), .B(b[0]), .Z(n13700) );
  XNOR U14772 ( .A(n13700), .B(n2175), .Z(n13702) );
  NANDN U14773 ( .A(b[0]), .B(a[546]), .Z(n13701) );
  NAND U14774 ( .A(n13702), .B(n13701), .Z(n13725) );
  XOR U14775 ( .A(n13724), .B(n13725), .Z(n13727) );
  XOR U14776 ( .A(n13726), .B(n13727), .Z(n13715) );
  NANDN U14777 ( .A(n13704), .B(n13703), .Z(n13708) );
  OR U14778 ( .A(n13706), .B(n13705), .Z(n13707) );
  AND U14779 ( .A(n13708), .B(n13707), .Z(n13714) );
  XOR U14780 ( .A(n13715), .B(n13714), .Z(n13717) );
  XOR U14781 ( .A(n13716), .B(n13717), .Z(n13730) );
  XNOR U14782 ( .A(n13730), .B(sreg[1567]), .Z(n13732) );
  NANDN U14783 ( .A(n13709), .B(sreg[1566]), .Z(n13713) );
  NAND U14784 ( .A(n13711), .B(n13710), .Z(n13712) );
  NAND U14785 ( .A(n13713), .B(n13712), .Z(n13731) );
  XOR U14786 ( .A(n13732), .B(n13731), .Z(c[1567]) );
  NANDN U14787 ( .A(n13715), .B(n13714), .Z(n13719) );
  OR U14788 ( .A(n13717), .B(n13716), .Z(n13718) );
  AND U14789 ( .A(n13719), .B(n13718), .Z(n13737) );
  XOR U14790 ( .A(a[546]), .B(n2254), .Z(n13741) );
  AND U14791 ( .A(a[548]), .B(b[0]), .Z(n13721) );
  XNOR U14792 ( .A(n13721), .B(n2175), .Z(n13723) );
  NANDN U14793 ( .A(b[0]), .B(a[547]), .Z(n13722) );
  NAND U14794 ( .A(n13723), .B(n13722), .Z(n13746) );
  AND U14795 ( .A(a[544]), .B(b[3]), .Z(n13745) );
  XOR U14796 ( .A(n13746), .B(n13745), .Z(n13748) );
  XOR U14797 ( .A(n13747), .B(n13748), .Z(n13736) );
  NANDN U14798 ( .A(n13725), .B(n13724), .Z(n13729) );
  OR U14799 ( .A(n13727), .B(n13726), .Z(n13728) );
  AND U14800 ( .A(n13729), .B(n13728), .Z(n13735) );
  XOR U14801 ( .A(n13736), .B(n13735), .Z(n13738) );
  XOR U14802 ( .A(n13737), .B(n13738), .Z(n13751) );
  XNOR U14803 ( .A(n13751), .B(sreg[1568]), .Z(n13753) );
  NANDN U14804 ( .A(n13730), .B(sreg[1567]), .Z(n13734) );
  NAND U14805 ( .A(n13732), .B(n13731), .Z(n13733) );
  NAND U14806 ( .A(n13734), .B(n13733), .Z(n13752) );
  XOR U14807 ( .A(n13753), .B(n13752), .Z(c[1568]) );
  NANDN U14808 ( .A(n13736), .B(n13735), .Z(n13740) );
  OR U14809 ( .A(n13738), .B(n13737), .Z(n13739) );
  AND U14810 ( .A(n13740), .B(n13739), .Z(n13758) );
  XOR U14811 ( .A(a[547]), .B(n2254), .Z(n13762) );
  AND U14812 ( .A(a[545]), .B(b[3]), .Z(n13766) );
  AND U14813 ( .A(a[549]), .B(b[0]), .Z(n13742) );
  XNOR U14814 ( .A(n13742), .B(n2175), .Z(n13744) );
  NANDN U14815 ( .A(b[0]), .B(a[548]), .Z(n13743) );
  NAND U14816 ( .A(n13744), .B(n13743), .Z(n13767) );
  XOR U14817 ( .A(n13766), .B(n13767), .Z(n13769) );
  XOR U14818 ( .A(n13768), .B(n13769), .Z(n13757) );
  NANDN U14819 ( .A(n13746), .B(n13745), .Z(n13750) );
  OR U14820 ( .A(n13748), .B(n13747), .Z(n13749) );
  AND U14821 ( .A(n13750), .B(n13749), .Z(n13756) );
  XOR U14822 ( .A(n13757), .B(n13756), .Z(n13759) );
  XOR U14823 ( .A(n13758), .B(n13759), .Z(n13772) );
  XNOR U14824 ( .A(n13772), .B(sreg[1569]), .Z(n13774) );
  NANDN U14825 ( .A(n13751), .B(sreg[1568]), .Z(n13755) );
  NAND U14826 ( .A(n13753), .B(n13752), .Z(n13754) );
  NAND U14827 ( .A(n13755), .B(n13754), .Z(n13773) );
  XOR U14828 ( .A(n13774), .B(n13773), .Z(c[1569]) );
  NANDN U14829 ( .A(n13757), .B(n13756), .Z(n13761) );
  OR U14830 ( .A(n13759), .B(n13758), .Z(n13760) );
  AND U14831 ( .A(n13761), .B(n13760), .Z(n13779) );
  XOR U14832 ( .A(a[548]), .B(n2254), .Z(n13783) );
  AND U14833 ( .A(a[550]), .B(b[0]), .Z(n13763) );
  XNOR U14834 ( .A(n13763), .B(n2175), .Z(n13765) );
  NANDN U14835 ( .A(b[0]), .B(a[549]), .Z(n13764) );
  NAND U14836 ( .A(n13765), .B(n13764), .Z(n13788) );
  AND U14837 ( .A(a[546]), .B(b[3]), .Z(n13787) );
  XOR U14838 ( .A(n13788), .B(n13787), .Z(n13790) );
  XOR U14839 ( .A(n13789), .B(n13790), .Z(n13778) );
  NANDN U14840 ( .A(n13767), .B(n13766), .Z(n13771) );
  OR U14841 ( .A(n13769), .B(n13768), .Z(n13770) );
  AND U14842 ( .A(n13771), .B(n13770), .Z(n13777) );
  XOR U14843 ( .A(n13778), .B(n13777), .Z(n13780) );
  XOR U14844 ( .A(n13779), .B(n13780), .Z(n13793) );
  XNOR U14845 ( .A(n13793), .B(sreg[1570]), .Z(n13795) );
  NANDN U14846 ( .A(n13772), .B(sreg[1569]), .Z(n13776) );
  NAND U14847 ( .A(n13774), .B(n13773), .Z(n13775) );
  NAND U14848 ( .A(n13776), .B(n13775), .Z(n13794) );
  XOR U14849 ( .A(n13795), .B(n13794), .Z(c[1570]) );
  NANDN U14850 ( .A(n13778), .B(n13777), .Z(n13782) );
  OR U14851 ( .A(n13780), .B(n13779), .Z(n13781) );
  AND U14852 ( .A(n13782), .B(n13781), .Z(n13800) );
  XOR U14853 ( .A(a[549]), .B(n2254), .Z(n13804) );
  AND U14854 ( .A(a[547]), .B(b[3]), .Z(n13808) );
  AND U14855 ( .A(a[551]), .B(b[0]), .Z(n13784) );
  XNOR U14856 ( .A(n13784), .B(n2175), .Z(n13786) );
  NANDN U14857 ( .A(b[0]), .B(a[550]), .Z(n13785) );
  NAND U14858 ( .A(n13786), .B(n13785), .Z(n13809) );
  XOR U14859 ( .A(n13808), .B(n13809), .Z(n13811) );
  XOR U14860 ( .A(n13810), .B(n13811), .Z(n13799) );
  NANDN U14861 ( .A(n13788), .B(n13787), .Z(n13792) );
  OR U14862 ( .A(n13790), .B(n13789), .Z(n13791) );
  AND U14863 ( .A(n13792), .B(n13791), .Z(n13798) );
  XOR U14864 ( .A(n13799), .B(n13798), .Z(n13801) );
  XOR U14865 ( .A(n13800), .B(n13801), .Z(n13814) );
  XNOR U14866 ( .A(n13814), .B(sreg[1571]), .Z(n13816) );
  NANDN U14867 ( .A(n13793), .B(sreg[1570]), .Z(n13797) );
  NAND U14868 ( .A(n13795), .B(n13794), .Z(n13796) );
  NAND U14869 ( .A(n13797), .B(n13796), .Z(n13815) );
  XOR U14870 ( .A(n13816), .B(n13815), .Z(c[1571]) );
  NANDN U14871 ( .A(n13799), .B(n13798), .Z(n13803) );
  OR U14872 ( .A(n13801), .B(n13800), .Z(n13802) );
  AND U14873 ( .A(n13803), .B(n13802), .Z(n13822) );
  XOR U14874 ( .A(a[550]), .B(n2254), .Z(n13823) );
  NAND U14875 ( .A(a[552]), .B(b[0]), .Z(n13805) );
  XNOR U14876 ( .A(b[1]), .B(n13805), .Z(n13807) );
  NANDN U14877 ( .A(b[0]), .B(a[551]), .Z(n13806) );
  AND U14878 ( .A(n13807), .B(n13806), .Z(n13827) );
  AND U14879 ( .A(a[548]), .B(b[3]), .Z(n13828) );
  XOR U14880 ( .A(n13827), .B(n13828), .Z(n13829) );
  XNOR U14881 ( .A(n13830), .B(n13829), .Z(n13819) );
  NANDN U14882 ( .A(n13809), .B(n13808), .Z(n13813) );
  OR U14883 ( .A(n13811), .B(n13810), .Z(n13812) );
  AND U14884 ( .A(n13813), .B(n13812), .Z(n13820) );
  XNOR U14885 ( .A(n13819), .B(n13820), .Z(n13821) );
  XNOR U14886 ( .A(n13822), .B(n13821), .Z(n13833) );
  XNOR U14887 ( .A(n13833), .B(sreg[1572]), .Z(n13835) );
  NANDN U14888 ( .A(n13814), .B(sreg[1571]), .Z(n13818) );
  NAND U14889 ( .A(n13816), .B(n13815), .Z(n13817) );
  NAND U14890 ( .A(n13818), .B(n13817), .Z(n13834) );
  XOR U14891 ( .A(n13835), .B(n13834), .Z(c[1572]) );
  XOR U14892 ( .A(a[551]), .B(n2254), .Z(n13842) );
  AND U14893 ( .A(a[553]), .B(b[0]), .Z(n13824) );
  XNOR U14894 ( .A(n13824), .B(n2175), .Z(n13826) );
  NANDN U14895 ( .A(b[0]), .B(a[552]), .Z(n13825) );
  NAND U14896 ( .A(n13826), .B(n13825), .Z(n13847) );
  AND U14897 ( .A(a[549]), .B(b[3]), .Z(n13846) );
  XOR U14898 ( .A(n13847), .B(n13846), .Z(n13849) );
  XOR U14899 ( .A(n13848), .B(n13849), .Z(n13837) );
  NAND U14900 ( .A(n13828), .B(n13827), .Z(n13832) );
  NANDN U14901 ( .A(n13830), .B(n13829), .Z(n13831) );
  AND U14902 ( .A(n13832), .B(n13831), .Z(n13836) );
  XOR U14903 ( .A(n13837), .B(n13836), .Z(n13839) );
  XOR U14904 ( .A(n13838), .B(n13839), .Z(n13852) );
  XNOR U14905 ( .A(n13852), .B(sreg[1573]), .Z(n13854) );
  XOR U14906 ( .A(n13854), .B(n13853), .Z(c[1573]) );
  NANDN U14907 ( .A(n13837), .B(n13836), .Z(n13841) );
  OR U14908 ( .A(n13839), .B(n13838), .Z(n13840) );
  AND U14909 ( .A(n13841), .B(n13840), .Z(n13859) );
  XOR U14910 ( .A(a[552]), .B(n2255), .Z(n13863) );
  AND U14911 ( .A(a[550]), .B(b[3]), .Z(n13867) );
  AND U14912 ( .A(a[554]), .B(b[0]), .Z(n13843) );
  XNOR U14913 ( .A(n13843), .B(n2175), .Z(n13845) );
  NANDN U14914 ( .A(b[0]), .B(a[553]), .Z(n13844) );
  NAND U14915 ( .A(n13845), .B(n13844), .Z(n13868) );
  XOR U14916 ( .A(n13867), .B(n13868), .Z(n13870) );
  XOR U14917 ( .A(n13869), .B(n13870), .Z(n13858) );
  NANDN U14918 ( .A(n13847), .B(n13846), .Z(n13851) );
  OR U14919 ( .A(n13849), .B(n13848), .Z(n13850) );
  AND U14920 ( .A(n13851), .B(n13850), .Z(n13857) );
  XOR U14921 ( .A(n13858), .B(n13857), .Z(n13860) );
  XOR U14922 ( .A(n13859), .B(n13860), .Z(n13873) );
  XNOR U14923 ( .A(n13873), .B(sreg[1574]), .Z(n13875) );
  NANDN U14924 ( .A(n13852), .B(sreg[1573]), .Z(n13856) );
  NAND U14925 ( .A(n13854), .B(n13853), .Z(n13855) );
  NAND U14926 ( .A(n13856), .B(n13855), .Z(n13874) );
  XOR U14927 ( .A(n13875), .B(n13874), .Z(c[1574]) );
  NANDN U14928 ( .A(n13858), .B(n13857), .Z(n13862) );
  OR U14929 ( .A(n13860), .B(n13859), .Z(n13861) );
  AND U14930 ( .A(n13862), .B(n13861), .Z(n13880) );
  XOR U14931 ( .A(a[553]), .B(n2255), .Z(n13884) );
  AND U14932 ( .A(a[555]), .B(b[0]), .Z(n13864) );
  XNOR U14933 ( .A(n13864), .B(n2175), .Z(n13866) );
  NANDN U14934 ( .A(b[0]), .B(a[554]), .Z(n13865) );
  NAND U14935 ( .A(n13866), .B(n13865), .Z(n13889) );
  AND U14936 ( .A(a[551]), .B(b[3]), .Z(n13888) );
  XOR U14937 ( .A(n13889), .B(n13888), .Z(n13891) );
  XOR U14938 ( .A(n13890), .B(n13891), .Z(n13879) );
  NANDN U14939 ( .A(n13868), .B(n13867), .Z(n13872) );
  OR U14940 ( .A(n13870), .B(n13869), .Z(n13871) );
  AND U14941 ( .A(n13872), .B(n13871), .Z(n13878) );
  XOR U14942 ( .A(n13879), .B(n13878), .Z(n13881) );
  XOR U14943 ( .A(n13880), .B(n13881), .Z(n13894) );
  XNOR U14944 ( .A(n13894), .B(sreg[1575]), .Z(n13896) );
  NANDN U14945 ( .A(n13873), .B(sreg[1574]), .Z(n13877) );
  NAND U14946 ( .A(n13875), .B(n13874), .Z(n13876) );
  NAND U14947 ( .A(n13877), .B(n13876), .Z(n13895) );
  XOR U14948 ( .A(n13896), .B(n13895), .Z(c[1575]) );
  NANDN U14949 ( .A(n13879), .B(n13878), .Z(n13883) );
  OR U14950 ( .A(n13881), .B(n13880), .Z(n13882) );
  AND U14951 ( .A(n13883), .B(n13882), .Z(n13901) );
  XOR U14952 ( .A(a[554]), .B(n2255), .Z(n13905) );
  AND U14953 ( .A(a[556]), .B(b[0]), .Z(n13885) );
  XNOR U14954 ( .A(n13885), .B(n2175), .Z(n13887) );
  NANDN U14955 ( .A(b[0]), .B(a[555]), .Z(n13886) );
  NAND U14956 ( .A(n13887), .B(n13886), .Z(n13910) );
  AND U14957 ( .A(a[552]), .B(b[3]), .Z(n13909) );
  XOR U14958 ( .A(n13910), .B(n13909), .Z(n13912) );
  XOR U14959 ( .A(n13911), .B(n13912), .Z(n13900) );
  NANDN U14960 ( .A(n13889), .B(n13888), .Z(n13893) );
  OR U14961 ( .A(n13891), .B(n13890), .Z(n13892) );
  AND U14962 ( .A(n13893), .B(n13892), .Z(n13899) );
  XOR U14963 ( .A(n13900), .B(n13899), .Z(n13902) );
  XOR U14964 ( .A(n13901), .B(n13902), .Z(n13915) );
  XNOR U14965 ( .A(n13915), .B(sreg[1576]), .Z(n13917) );
  NANDN U14966 ( .A(n13894), .B(sreg[1575]), .Z(n13898) );
  NAND U14967 ( .A(n13896), .B(n13895), .Z(n13897) );
  NAND U14968 ( .A(n13898), .B(n13897), .Z(n13916) );
  XOR U14969 ( .A(n13917), .B(n13916), .Z(c[1576]) );
  NANDN U14970 ( .A(n13900), .B(n13899), .Z(n13904) );
  OR U14971 ( .A(n13902), .B(n13901), .Z(n13903) );
  AND U14972 ( .A(n13904), .B(n13903), .Z(n13922) );
  XOR U14973 ( .A(a[555]), .B(n2255), .Z(n13926) );
  AND U14974 ( .A(a[553]), .B(b[3]), .Z(n13930) );
  AND U14975 ( .A(a[557]), .B(b[0]), .Z(n13906) );
  XNOR U14976 ( .A(n13906), .B(n2175), .Z(n13908) );
  NANDN U14977 ( .A(b[0]), .B(a[556]), .Z(n13907) );
  NAND U14978 ( .A(n13908), .B(n13907), .Z(n13931) );
  XOR U14979 ( .A(n13930), .B(n13931), .Z(n13933) );
  XOR U14980 ( .A(n13932), .B(n13933), .Z(n13921) );
  NANDN U14981 ( .A(n13910), .B(n13909), .Z(n13914) );
  OR U14982 ( .A(n13912), .B(n13911), .Z(n13913) );
  AND U14983 ( .A(n13914), .B(n13913), .Z(n13920) );
  XOR U14984 ( .A(n13921), .B(n13920), .Z(n13923) );
  XOR U14985 ( .A(n13922), .B(n13923), .Z(n13936) );
  XNOR U14986 ( .A(n13936), .B(sreg[1577]), .Z(n13938) );
  NANDN U14987 ( .A(n13915), .B(sreg[1576]), .Z(n13919) );
  NAND U14988 ( .A(n13917), .B(n13916), .Z(n13918) );
  NAND U14989 ( .A(n13919), .B(n13918), .Z(n13937) );
  XOR U14990 ( .A(n13938), .B(n13937), .Z(c[1577]) );
  NANDN U14991 ( .A(n13921), .B(n13920), .Z(n13925) );
  OR U14992 ( .A(n13923), .B(n13922), .Z(n13924) );
  AND U14993 ( .A(n13925), .B(n13924), .Z(n13943) );
  XOR U14994 ( .A(a[556]), .B(n2255), .Z(n13947) );
  AND U14995 ( .A(a[554]), .B(b[3]), .Z(n13951) );
  AND U14996 ( .A(a[558]), .B(b[0]), .Z(n13927) );
  XNOR U14997 ( .A(n13927), .B(n2175), .Z(n13929) );
  NANDN U14998 ( .A(b[0]), .B(a[557]), .Z(n13928) );
  NAND U14999 ( .A(n13929), .B(n13928), .Z(n13952) );
  XOR U15000 ( .A(n13951), .B(n13952), .Z(n13954) );
  XOR U15001 ( .A(n13953), .B(n13954), .Z(n13942) );
  NANDN U15002 ( .A(n13931), .B(n13930), .Z(n13935) );
  OR U15003 ( .A(n13933), .B(n13932), .Z(n13934) );
  AND U15004 ( .A(n13935), .B(n13934), .Z(n13941) );
  XOR U15005 ( .A(n13942), .B(n13941), .Z(n13944) );
  XOR U15006 ( .A(n13943), .B(n13944), .Z(n13957) );
  XNOR U15007 ( .A(n13957), .B(sreg[1578]), .Z(n13959) );
  NANDN U15008 ( .A(n13936), .B(sreg[1577]), .Z(n13940) );
  NAND U15009 ( .A(n13938), .B(n13937), .Z(n13939) );
  NAND U15010 ( .A(n13940), .B(n13939), .Z(n13958) );
  XOR U15011 ( .A(n13959), .B(n13958), .Z(c[1578]) );
  NANDN U15012 ( .A(n13942), .B(n13941), .Z(n13946) );
  OR U15013 ( .A(n13944), .B(n13943), .Z(n13945) );
  AND U15014 ( .A(n13946), .B(n13945), .Z(n13964) );
  XOR U15015 ( .A(a[557]), .B(n2255), .Z(n13968) );
  AND U15016 ( .A(a[555]), .B(b[3]), .Z(n13972) );
  AND U15017 ( .A(a[559]), .B(b[0]), .Z(n13948) );
  XNOR U15018 ( .A(n13948), .B(n2175), .Z(n13950) );
  NANDN U15019 ( .A(b[0]), .B(a[558]), .Z(n13949) );
  NAND U15020 ( .A(n13950), .B(n13949), .Z(n13973) );
  XOR U15021 ( .A(n13972), .B(n13973), .Z(n13975) );
  XOR U15022 ( .A(n13974), .B(n13975), .Z(n13963) );
  NANDN U15023 ( .A(n13952), .B(n13951), .Z(n13956) );
  OR U15024 ( .A(n13954), .B(n13953), .Z(n13955) );
  AND U15025 ( .A(n13956), .B(n13955), .Z(n13962) );
  XOR U15026 ( .A(n13963), .B(n13962), .Z(n13965) );
  XOR U15027 ( .A(n13964), .B(n13965), .Z(n13978) );
  XNOR U15028 ( .A(n13978), .B(sreg[1579]), .Z(n13980) );
  NANDN U15029 ( .A(n13957), .B(sreg[1578]), .Z(n13961) );
  NAND U15030 ( .A(n13959), .B(n13958), .Z(n13960) );
  NAND U15031 ( .A(n13961), .B(n13960), .Z(n13979) );
  XOR U15032 ( .A(n13980), .B(n13979), .Z(c[1579]) );
  NANDN U15033 ( .A(n13963), .B(n13962), .Z(n13967) );
  OR U15034 ( .A(n13965), .B(n13964), .Z(n13966) );
  AND U15035 ( .A(n13967), .B(n13966), .Z(n13985) );
  XOR U15036 ( .A(a[558]), .B(n2255), .Z(n13989) );
  AND U15037 ( .A(a[560]), .B(b[0]), .Z(n13969) );
  XNOR U15038 ( .A(n13969), .B(n2175), .Z(n13971) );
  NANDN U15039 ( .A(b[0]), .B(a[559]), .Z(n13970) );
  NAND U15040 ( .A(n13971), .B(n13970), .Z(n13994) );
  AND U15041 ( .A(a[556]), .B(b[3]), .Z(n13993) );
  XOR U15042 ( .A(n13994), .B(n13993), .Z(n13996) );
  XOR U15043 ( .A(n13995), .B(n13996), .Z(n13984) );
  NANDN U15044 ( .A(n13973), .B(n13972), .Z(n13977) );
  OR U15045 ( .A(n13975), .B(n13974), .Z(n13976) );
  AND U15046 ( .A(n13977), .B(n13976), .Z(n13983) );
  XOR U15047 ( .A(n13984), .B(n13983), .Z(n13986) );
  XOR U15048 ( .A(n13985), .B(n13986), .Z(n13999) );
  XNOR U15049 ( .A(n13999), .B(sreg[1580]), .Z(n14001) );
  NANDN U15050 ( .A(n13978), .B(sreg[1579]), .Z(n13982) );
  NAND U15051 ( .A(n13980), .B(n13979), .Z(n13981) );
  NAND U15052 ( .A(n13982), .B(n13981), .Z(n14000) );
  XOR U15053 ( .A(n14001), .B(n14000), .Z(c[1580]) );
  NANDN U15054 ( .A(n13984), .B(n13983), .Z(n13988) );
  OR U15055 ( .A(n13986), .B(n13985), .Z(n13987) );
  AND U15056 ( .A(n13988), .B(n13987), .Z(n14006) );
  XOR U15057 ( .A(a[559]), .B(n2256), .Z(n14010) );
  AND U15058 ( .A(a[557]), .B(b[3]), .Z(n14014) );
  AND U15059 ( .A(a[561]), .B(b[0]), .Z(n13990) );
  XNOR U15060 ( .A(n13990), .B(n2175), .Z(n13992) );
  NANDN U15061 ( .A(b[0]), .B(a[560]), .Z(n13991) );
  NAND U15062 ( .A(n13992), .B(n13991), .Z(n14015) );
  XOR U15063 ( .A(n14014), .B(n14015), .Z(n14017) );
  XOR U15064 ( .A(n14016), .B(n14017), .Z(n14005) );
  NANDN U15065 ( .A(n13994), .B(n13993), .Z(n13998) );
  OR U15066 ( .A(n13996), .B(n13995), .Z(n13997) );
  AND U15067 ( .A(n13998), .B(n13997), .Z(n14004) );
  XOR U15068 ( .A(n14005), .B(n14004), .Z(n14007) );
  XOR U15069 ( .A(n14006), .B(n14007), .Z(n14020) );
  XNOR U15070 ( .A(n14020), .B(sreg[1581]), .Z(n14022) );
  NANDN U15071 ( .A(n13999), .B(sreg[1580]), .Z(n14003) );
  NAND U15072 ( .A(n14001), .B(n14000), .Z(n14002) );
  NAND U15073 ( .A(n14003), .B(n14002), .Z(n14021) );
  XOR U15074 ( .A(n14022), .B(n14021), .Z(c[1581]) );
  NANDN U15075 ( .A(n14005), .B(n14004), .Z(n14009) );
  OR U15076 ( .A(n14007), .B(n14006), .Z(n14008) );
  AND U15077 ( .A(n14009), .B(n14008), .Z(n14027) );
  XOR U15078 ( .A(a[560]), .B(n2256), .Z(n14031) );
  AND U15079 ( .A(a[562]), .B(b[0]), .Z(n14011) );
  XNOR U15080 ( .A(n14011), .B(n2175), .Z(n14013) );
  NANDN U15081 ( .A(b[0]), .B(a[561]), .Z(n14012) );
  NAND U15082 ( .A(n14013), .B(n14012), .Z(n14036) );
  AND U15083 ( .A(a[558]), .B(b[3]), .Z(n14035) );
  XOR U15084 ( .A(n14036), .B(n14035), .Z(n14038) );
  XOR U15085 ( .A(n14037), .B(n14038), .Z(n14026) );
  NANDN U15086 ( .A(n14015), .B(n14014), .Z(n14019) );
  OR U15087 ( .A(n14017), .B(n14016), .Z(n14018) );
  AND U15088 ( .A(n14019), .B(n14018), .Z(n14025) );
  XOR U15089 ( .A(n14026), .B(n14025), .Z(n14028) );
  XOR U15090 ( .A(n14027), .B(n14028), .Z(n14041) );
  XNOR U15091 ( .A(n14041), .B(sreg[1582]), .Z(n14043) );
  NANDN U15092 ( .A(n14020), .B(sreg[1581]), .Z(n14024) );
  NAND U15093 ( .A(n14022), .B(n14021), .Z(n14023) );
  NAND U15094 ( .A(n14024), .B(n14023), .Z(n14042) );
  XOR U15095 ( .A(n14043), .B(n14042), .Z(c[1582]) );
  NANDN U15096 ( .A(n14026), .B(n14025), .Z(n14030) );
  OR U15097 ( .A(n14028), .B(n14027), .Z(n14029) );
  AND U15098 ( .A(n14030), .B(n14029), .Z(n14048) );
  XOR U15099 ( .A(a[561]), .B(n2256), .Z(n14052) );
  AND U15100 ( .A(a[563]), .B(b[0]), .Z(n14032) );
  XNOR U15101 ( .A(n14032), .B(n2175), .Z(n14034) );
  NANDN U15102 ( .A(b[0]), .B(a[562]), .Z(n14033) );
  NAND U15103 ( .A(n14034), .B(n14033), .Z(n14057) );
  AND U15104 ( .A(a[559]), .B(b[3]), .Z(n14056) );
  XOR U15105 ( .A(n14057), .B(n14056), .Z(n14059) );
  XOR U15106 ( .A(n14058), .B(n14059), .Z(n14047) );
  NANDN U15107 ( .A(n14036), .B(n14035), .Z(n14040) );
  OR U15108 ( .A(n14038), .B(n14037), .Z(n14039) );
  AND U15109 ( .A(n14040), .B(n14039), .Z(n14046) );
  XOR U15110 ( .A(n14047), .B(n14046), .Z(n14049) );
  XOR U15111 ( .A(n14048), .B(n14049), .Z(n14062) );
  XNOR U15112 ( .A(n14062), .B(sreg[1583]), .Z(n14064) );
  NANDN U15113 ( .A(n14041), .B(sreg[1582]), .Z(n14045) );
  NAND U15114 ( .A(n14043), .B(n14042), .Z(n14044) );
  NAND U15115 ( .A(n14045), .B(n14044), .Z(n14063) );
  XOR U15116 ( .A(n14064), .B(n14063), .Z(c[1583]) );
  NANDN U15117 ( .A(n14047), .B(n14046), .Z(n14051) );
  OR U15118 ( .A(n14049), .B(n14048), .Z(n14050) );
  AND U15119 ( .A(n14051), .B(n14050), .Z(n14069) );
  XOR U15120 ( .A(a[562]), .B(n2256), .Z(n14073) );
  AND U15121 ( .A(a[560]), .B(b[3]), .Z(n14077) );
  AND U15122 ( .A(a[564]), .B(b[0]), .Z(n14053) );
  XNOR U15123 ( .A(n14053), .B(n2175), .Z(n14055) );
  NANDN U15124 ( .A(b[0]), .B(a[563]), .Z(n14054) );
  NAND U15125 ( .A(n14055), .B(n14054), .Z(n14078) );
  XOR U15126 ( .A(n14077), .B(n14078), .Z(n14080) );
  XOR U15127 ( .A(n14079), .B(n14080), .Z(n14068) );
  NANDN U15128 ( .A(n14057), .B(n14056), .Z(n14061) );
  OR U15129 ( .A(n14059), .B(n14058), .Z(n14060) );
  AND U15130 ( .A(n14061), .B(n14060), .Z(n14067) );
  XOR U15131 ( .A(n14068), .B(n14067), .Z(n14070) );
  XOR U15132 ( .A(n14069), .B(n14070), .Z(n14083) );
  XNOR U15133 ( .A(n14083), .B(sreg[1584]), .Z(n14085) );
  NANDN U15134 ( .A(n14062), .B(sreg[1583]), .Z(n14066) );
  NAND U15135 ( .A(n14064), .B(n14063), .Z(n14065) );
  NAND U15136 ( .A(n14066), .B(n14065), .Z(n14084) );
  XOR U15137 ( .A(n14085), .B(n14084), .Z(c[1584]) );
  NANDN U15138 ( .A(n14068), .B(n14067), .Z(n14072) );
  OR U15139 ( .A(n14070), .B(n14069), .Z(n14071) );
  AND U15140 ( .A(n14072), .B(n14071), .Z(n14090) );
  XOR U15141 ( .A(a[563]), .B(n2256), .Z(n14094) );
  AND U15142 ( .A(a[565]), .B(b[0]), .Z(n14074) );
  XNOR U15143 ( .A(n14074), .B(n2175), .Z(n14076) );
  NANDN U15144 ( .A(b[0]), .B(a[564]), .Z(n14075) );
  NAND U15145 ( .A(n14076), .B(n14075), .Z(n14099) );
  AND U15146 ( .A(a[561]), .B(b[3]), .Z(n14098) );
  XOR U15147 ( .A(n14099), .B(n14098), .Z(n14101) );
  XOR U15148 ( .A(n14100), .B(n14101), .Z(n14089) );
  NANDN U15149 ( .A(n14078), .B(n14077), .Z(n14082) );
  OR U15150 ( .A(n14080), .B(n14079), .Z(n14081) );
  AND U15151 ( .A(n14082), .B(n14081), .Z(n14088) );
  XOR U15152 ( .A(n14089), .B(n14088), .Z(n14091) );
  XOR U15153 ( .A(n14090), .B(n14091), .Z(n14104) );
  XNOR U15154 ( .A(n14104), .B(sreg[1585]), .Z(n14106) );
  NANDN U15155 ( .A(n14083), .B(sreg[1584]), .Z(n14087) );
  NAND U15156 ( .A(n14085), .B(n14084), .Z(n14086) );
  NAND U15157 ( .A(n14087), .B(n14086), .Z(n14105) );
  XOR U15158 ( .A(n14106), .B(n14105), .Z(c[1585]) );
  NANDN U15159 ( .A(n14089), .B(n14088), .Z(n14093) );
  OR U15160 ( .A(n14091), .B(n14090), .Z(n14092) );
  AND U15161 ( .A(n14093), .B(n14092), .Z(n14111) );
  XOR U15162 ( .A(a[564]), .B(n2256), .Z(n14115) );
  AND U15163 ( .A(a[566]), .B(b[0]), .Z(n14095) );
  XNOR U15164 ( .A(n14095), .B(n2175), .Z(n14097) );
  NANDN U15165 ( .A(b[0]), .B(a[565]), .Z(n14096) );
  NAND U15166 ( .A(n14097), .B(n14096), .Z(n14120) );
  AND U15167 ( .A(a[562]), .B(b[3]), .Z(n14119) );
  XOR U15168 ( .A(n14120), .B(n14119), .Z(n14122) );
  XOR U15169 ( .A(n14121), .B(n14122), .Z(n14110) );
  NANDN U15170 ( .A(n14099), .B(n14098), .Z(n14103) );
  OR U15171 ( .A(n14101), .B(n14100), .Z(n14102) );
  AND U15172 ( .A(n14103), .B(n14102), .Z(n14109) );
  XOR U15173 ( .A(n14110), .B(n14109), .Z(n14112) );
  XOR U15174 ( .A(n14111), .B(n14112), .Z(n14125) );
  XNOR U15175 ( .A(n14125), .B(sreg[1586]), .Z(n14127) );
  NANDN U15176 ( .A(n14104), .B(sreg[1585]), .Z(n14108) );
  NAND U15177 ( .A(n14106), .B(n14105), .Z(n14107) );
  NAND U15178 ( .A(n14108), .B(n14107), .Z(n14126) );
  XOR U15179 ( .A(n14127), .B(n14126), .Z(c[1586]) );
  NANDN U15180 ( .A(n14110), .B(n14109), .Z(n14114) );
  OR U15181 ( .A(n14112), .B(n14111), .Z(n14113) );
  AND U15182 ( .A(n14114), .B(n14113), .Z(n14132) );
  XOR U15183 ( .A(a[565]), .B(n2256), .Z(n14136) );
  AND U15184 ( .A(a[567]), .B(b[0]), .Z(n14116) );
  XNOR U15185 ( .A(n14116), .B(n2175), .Z(n14118) );
  NANDN U15186 ( .A(b[0]), .B(a[566]), .Z(n14117) );
  NAND U15187 ( .A(n14118), .B(n14117), .Z(n14141) );
  AND U15188 ( .A(a[563]), .B(b[3]), .Z(n14140) );
  XOR U15189 ( .A(n14141), .B(n14140), .Z(n14143) );
  XOR U15190 ( .A(n14142), .B(n14143), .Z(n14131) );
  NANDN U15191 ( .A(n14120), .B(n14119), .Z(n14124) );
  OR U15192 ( .A(n14122), .B(n14121), .Z(n14123) );
  AND U15193 ( .A(n14124), .B(n14123), .Z(n14130) );
  XOR U15194 ( .A(n14131), .B(n14130), .Z(n14133) );
  XOR U15195 ( .A(n14132), .B(n14133), .Z(n14146) );
  XNOR U15196 ( .A(n14146), .B(sreg[1587]), .Z(n14148) );
  NANDN U15197 ( .A(n14125), .B(sreg[1586]), .Z(n14129) );
  NAND U15198 ( .A(n14127), .B(n14126), .Z(n14128) );
  NAND U15199 ( .A(n14129), .B(n14128), .Z(n14147) );
  XOR U15200 ( .A(n14148), .B(n14147), .Z(c[1587]) );
  NANDN U15201 ( .A(n14131), .B(n14130), .Z(n14135) );
  OR U15202 ( .A(n14133), .B(n14132), .Z(n14134) );
  AND U15203 ( .A(n14135), .B(n14134), .Z(n14153) );
  XOR U15204 ( .A(a[566]), .B(n2257), .Z(n14157) );
  AND U15205 ( .A(a[568]), .B(b[0]), .Z(n14137) );
  XNOR U15206 ( .A(n14137), .B(n2175), .Z(n14139) );
  NANDN U15207 ( .A(b[0]), .B(a[567]), .Z(n14138) );
  NAND U15208 ( .A(n14139), .B(n14138), .Z(n14162) );
  AND U15209 ( .A(a[564]), .B(b[3]), .Z(n14161) );
  XOR U15210 ( .A(n14162), .B(n14161), .Z(n14164) );
  XOR U15211 ( .A(n14163), .B(n14164), .Z(n14152) );
  NANDN U15212 ( .A(n14141), .B(n14140), .Z(n14145) );
  OR U15213 ( .A(n14143), .B(n14142), .Z(n14144) );
  AND U15214 ( .A(n14145), .B(n14144), .Z(n14151) );
  XOR U15215 ( .A(n14152), .B(n14151), .Z(n14154) );
  XOR U15216 ( .A(n14153), .B(n14154), .Z(n14167) );
  XNOR U15217 ( .A(n14167), .B(sreg[1588]), .Z(n14169) );
  NANDN U15218 ( .A(n14146), .B(sreg[1587]), .Z(n14150) );
  NAND U15219 ( .A(n14148), .B(n14147), .Z(n14149) );
  NAND U15220 ( .A(n14150), .B(n14149), .Z(n14168) );
  XOR U15221 ( .A(n14169), .B(n14168), .Z(c[1588]) );
  NANDN U15222 ( .A(n14152), .B(n14151), .Z(n14156) );
  OR U15223 ( .A(n14154), .B(n14153), .Z(n14155) );
  AND U15224 ( .A(n14156), .B(n14155), .Z(n14174) );
  XOR U15225 ( .A(a[567]), .B(n2257), .Z(n14178) );
  AND U15226 ( .A(a[565]), .B(b[3]), .Z(n14182) );
  AND U15227 ( .A(a[569]), .B(b[0]), .Z(n14158) );
  XNOR U15228 ( .A(n14158), .B(n2175), .Z(n14160) );
  NANDN U15229 ( .A(b[0]), .B(a[568]), .Z(n14159) );
  NAND U15230 ( .A(n14160), .B(n14159), .Z(n14183) );
  XOR U15231 ( .A(n14182), .B(n14183), .Z(n14185) );
  XOR U15232 ( .A(n14184), .B(n14185), .Z(n14173) );
  NANDN U15233 ( .A(n14162), .B(n14161), .Z(n14166) );
  OR U15234 ( .A(n14164), .B(n14163), .Z(n14165) );
  AND U15235 ( .A(n14166), .B(n14165), .Z(n14172) );
  XOR U15236 ( .A(n14173), .B(n14172), .Z(n14175) );
  XOR U15237 ( .A(n14174), .B(n14175), .Z(n14188) );
  XNOR U15238 ( .A(n14188), .B(sreg[1589]), .Z(n14190) );
  NANDN U15239 ( .A(n14167), .B(sreg[1588]), .Z(n14171) );
  NAND U15240 ( .A(n14169), .B(n14168), .Z(n14170) );
  NAND U15241 ( .A(n14171), .B(n14170), .Z(n14189) );
  XOR U15242 ( .A(n14190), .B(n14189), .Z(c[1589]) );
  NANDN U15243 ( .A(n14173), .B(n14172), .Z(n14177) );
  OR U15244 ( .A(n14175), .B(n14174), .Z(n14176) );
  AND U15245 ( .A(n14177), .B(n14176), .Z(n14195) );
  XOR U15246 ( .A(a[568]), .B(n2257), .Z(n14199) );
  AND U15247 ( .A(a[570]), .B(b[0]), .Z(n14179) );
  XNOR U15248 ( .A(n14179), .B(n2175), .Z(n14181) );
  NANDN U15249 ( .A(b[0]), .B(a[569]), .Z(n14180) );
  NAND U15250 ( .A(n14181), .B(n14180), .Z(n14204) );
  AND U15251 ( .A(a[566]), .B(b[3]), .Z(n14203) );
  XOR U15252 ( .A(n14204), .B(n14203), .Z(n14206) );
  XOR U15253 ( .A(n14205), .B(n14206), .Z(n14194) );
  NANDN U15254 ( .A(n14183), .B(n14182), .Z(n14187) );
  OR U15255 ( .A(n14185), .B(n14184), .Z(n14186) );
  AND U15256 ( .A(n14187), .B(n14186), .Z(n14193) );
  XOR U15257 ( .A(n14194), .B(n14193), .Z(n14196) );
  XOR U15258 ( .A(n14195), .B(n14196), .Z(n14209) );
  XNOR U15259 ( .A(n14209), .B(sreg[1590]), .Z(n14211) );
  NANDN U15260 ( .A(n14188), .B(sreg[1589]), .Z(n14192) );
  NAND U15261 ( .A(n14190), .B(n14189), .Z(n14191) );
  NAND U15262 ( .A(n14192), .B(n14191), .Z(n14210) );
  XOR U15263 ( .A(n14211), .B(n14210), .Z(c[1590]) );
  NANDN U15264 ( .A(n14194), .B(n14193), .Z(n14198) );
  OR U15265 ( .A(n14196), .B(n14195), .Z(n14197) );
  AND U15266 ( .A(n14198), .B(n14197), .Z(n14216) );
  XOR U15267 ( .A(a[569]), .B(n2257), .Z(n14220) );
  AND U15268 ( .A(a[567]), .B(b[3]), .Z(n14224) );
  AND U15269 ( .A(a[571]), .B(b[0]), .Z(n14200) );
  XNOR U15270 ( .A(n14200), .B(n2175), .Z(n14202) );
  NANDN U15271 ( .A(b[0]), .B(a[570]), .Z(n14201) );
  NAND U15272 ( .A(n14202), .B(n14201), .Z(n14225) );
  XOR U15273 ( .A(n14224), .B(n14225), .Z(n14227) );
  XOR U15274 ( .A(n14226), .B(n14227), .Z(n14215) );
  NANDN U15275 ( .A(n14204), .B(n14203), .Z(n14208) );
  OR U15276 ( .A(n14206), .B(n14205), .Z(n14207) );
  AND U15277 ( .A(n14208), .B(n14207), .Z(n14214) );
  XOR U15278 ( .A(n14215), .B(n14214), .Z(n14217) );
  XOR U15279 ( .A(n14216), .B(n14217), .Z(n14230) );
  XNOR U15280 ( .A(n14230), .B(sreg[1591]), .Z(n14232) );
  NANDN U15281 ( .A(n14209), .B(sreg[1590]), .Z(n14213) );
  NAND U15282 ( .A(n14211), .B(n14210), .Z(n14212) );
  NAND U15283 ( .A(n14213), .B(n14212), .Z(n14231) );
  XOR U15284 ( .A(n14232), .B(n14231), .Z(c[1591]) );
  NANDN U15285 ( .A(n14215), .B(n14214), .Z(n14219) );
  OR U15286 ( .A(n14217), .B(n14216), .Z(n14218) );
  AND U15287 ( .A(n14219), .B(n14218), .Z(n14237) );
  XOR U15288 ( .A(a[570]), .B(n2257), .Z(n14241) );
  AND U15289 ( .A(a[572]), .B(b[0]), .Z(n14221) );
  XNOR U15290 ( .A(n14221), .B(n2175), .Z(n14223) );
  NANDN U15291 ( .A(b[0]), .B(a[571]), .Z(n14222) );
  NAND U15292 ( .A(n14223), .B(n14222), .Z(n14246) );
  AND U15293 ( .A(a[568]), .B(b[3]), .Z(n14245) );
  XOR U15294 ( .A(n14246), .B(n14245), .Z(n14248) );
  XOR U15295 ( .A(n14247), .B(n14248), .Z(n14236) );
  NANDN U15296 ( .A(n14225), .B(n14224), .Z(n14229) );
  OR U15297 ( .A(n14227), .B(n14226), .Z(n14228) );
  AND U15298 ( .A(n14229), .B(n14228), .Z(n14235) );
  XOR U15299 ( .A(n14236), .B(n14235), .Z(n14238) );
  XOR U15300 ( .A(n14237), .B(n14238), .Z(n14251) );
  XNOR U15301 ( .A(n14251), .B(sreg[1592]), .Z(n14253) );
  NANDN U15302 ( .A(n14230), .B(sreg[1591]), .Z(n14234) );
  NAND U15303 ( .A(n14232), .B(n14231), .Z(n14233) );
  NAND U15304 ( .A(n14234), .B(n14233), .Z(n14252) );
  XOR U15305 ( .A(n14253), .B(n14252), .Z(c[1592]) );
  NANDN U15306 ( .A(n14236), .B(n14235), .Z(n14240) );
  OR U15307 ( .A(n14238), .B(n14237), .Z(n14239) );
  AND U15308 ( .A(n14240), .B(n14239), .Z(n14258) );
  XOR U15309 ( .A(a[571]), .B(n2257), .Z(n14262) );
  AND U15310 ( .A(a[569]), .B(b[3]), .Z(n14266) );
  AND U15311 ( .A(a[573]), .B(b[0]), .Z(n14242) );
  XNOR U15312 ( .A(n14242), .B(n2175), .Z(n14244) );
  NANDN U15313 ( .A(b[0]), .B(a[572]), .Z(n14243) );
  NAND U15314 ( .A(n14244), .B(n14243), .Z(n14267) );
  XOR U15315 ( .A(n14266), .B(n14267), .Z(n14269) );
  XOR U15316 ( .A(n14268), .B(n14269), .Z(n14257) );
  NANDN U15317 ( .A(n14246), .B(n14245), .Z(n14250) );
  OR U15318 ( .A(n14248), .B(n14247), .Z(n14249) );
  AND U15319 ( .A(n14250), .B(n14249), .Z(n14256) );
  XOR U15320 ( .A(n14257), .B(n14256), .Z(n14259) );
  XOR U15321 ( .A(n14258), .B(n14259), .Z(n14272) );
  XNOR U15322 ( .A(n14272), .B(sreg[1593]), .Z(n14274) );
  NANDN U15323 ( .A(n14251), .B(sreg[1592]), .Z(n14255) );
  NAND U15324 ( .A(n14253), .B(n14252), .Z(n14254) );
  NAND U15325 ( .A(n14255), .B(n14254), .Z(n14273) );
  XOR U15326 ( .A(n14274), .B(n14273), .Z(c[1593]) );
  NANDN U15327 ( .A(n14257), .B(n14256), .Z(n14261) );
  OR U15328 ( .A(n14259), .B(n14258), .Z(n14260) );
  AND U15329 ( .A(n14261), .B(n14260), .Z(n14279) );
  XOR U15330 ( .A(a[572]), .B(n2257), .Z(n14283) );
  AND U15331 ( .A(a[574]), .B(b[0]), .Z(n14263) );
  XNOR U15332 ( .A(n14263), .B(n2175), .Z(n14265) );
  NANDN U15333 ( .A(b[0]), .B(a[573]), .Z(n14264) );
  NAND U15334 ( .A(n14265), .B(n14264), .Z(n14288) );
  AND U15335 ( .A(a[570]), .B(b[3]), .Z(n14287) );
  XOR U15336 ( .A(n14288), .B(n14287), .Z(n14290) );
  XOR U15337 ( .A(n14289), .B(n14290), .Z(n14278) );
  NANDN U15338 ( .A(n14267), .B(n14266), .Z(n14271) );
  OR U15339 ( .A(n14269), .B(n14268), .Z(n14270) );
  AND U15340 ( .A(n14271), .B(n14270), .Z(n14277) );
  XOR U15341 ( .A(n14278), .B(n14277), .Z(n14280) );
  XOR U15342 ( .A(n14279), .B(n14280), .Z(n14293) );
  XNOR U15343 ( .A(n14293), .B(sreg[1594]), .Z(n14295) );
  NANDN U15344 ( .A(n14272), .B(sreg[1593]), .Z(n14276) );
  NAND U15345 ( .A(n14274), .B(n14273), .Z(n14275) );
  NAND U15346 ( .A(n14276), .B(n14275), .Z(n14294) );
  XOR U15347 ( .A(n14295), .B(n14294), .Z(c[1594]) );
  NANDN U15348 ( .A(n14278), .B(n14277), .Z(n14282) );
  OR U15349 ( .A(n14280), .B(n14279), .Z(n14281) );
  AND U15350 ( .A(n14282), .B(n14281), .Z(n14300) );
  XOR U15351 ( .A(a[573]), .B(n2258), .Z(n14304) );
  AND U15352 ( .A(a[575]), .B(b[0]), .Z(n14284) );
  XNOR U15353 ( .A(n14284), .B(n2175), .Z(n14286) );
  NANDN U15354 ( .A(b[0]), .B(a[574]), .Z(n14285) );
  NAND U15355 ( .A(n14286), .B(n14285), .Z(n14309) );
  AND U15356 ( .A(a[571]), .B(b[3]), .Z(n14308) );
  XOR U15357 ( .A(n14309), .B(n14308), .Z(n14311) );
  XOR U15358 ( .A(n14310), .B(n14311), .Z(n14299) );
  NANDN U15359 ( .A(n14288), .B(n14287), .Z(n14292) );
  OR U15360 ( .A(n14290), .B(n14289), .Z(n14291) );
  AND U15361 ( .A(n14292), .B(n14291), .Z(n14298) );
  XOR U15362 ( .A(n14299), .B(n14298), .Z(n14301) );
  XOR U15363 ( .A(n14300), .B(n14301), .Z(n14314) );
  XNOR U15364 ( .A(n14314), .B(sreg[1595]), .Z(n14316) );
  NANDN U15365 ( .A(n14293), .B(sreg[1594]), .Z(n14297) );
  NAND U15366 ( .A(n14295), .B(n14294), .Z(n14296) );
  NAND U15367 ( .A(n14297), .B(n14296), .Z(n14315) );
  XOR U15368 ( .A(n14316), .B(n14315), .Z(c[1595]) );
  NANDN U15369 ( .A(n14299), .B(n14298), .Z(n14303) );
  OR U15370 ( .A(n14301), .B(n14300), .Z(n14302) );
  AND U15371 ( .A(n14303), .B(n14302), .Z(n14321) );
  XOR U15372 ( .A(a[574]), .B(n2258), .Z(n14325) );
  AND U15373 ( .A(a[572]), .B(b[3]), .Z(n14329) );
  AND U15374 ( .A(a[576]), .B(b[0]), .Z(n14305) );
  XNOR U15375 ( .A(n14305), .B(n2175), .Z(n14307) );
  NANDN U15376 ( .A(b[0]), .B(a[575]), .Z(n14306) );
  NAND U15377 ( .A(n14307), .B(n14306), .Z(n14330) );
  XOR U15378 ( .A(n14329), .B(n14330), .Z(n14332) );
  XOR U15379 ( .A(n14331), .B(n14332), .Z(n14320) );
  NANDN U15380 ( .A(n14309), .B(n14308), .Z(n14313) );
  OR U15381 ( .A(n14311), .B(n14310), .Z(n14312) );
  AND U15382 ( .A(n14313), .B(n14312), .Z(n14319) );
  XOR U15383 ( .A(n14320), .B(n14319), .Z(n14322) );
  XOR U15384 ( .A(n14321), .B(n14322), .Z(n14335) );
  XNOR U15385 ( .A(n14335), .B(sreg[1596]), .Z(n14337) );
  NANDN U15386 ( .A(n14314), .B(sreg[1595]), .Z(n14318) );
  NAND U15387 ( .A(n14316), .B(n14315), .Z(n14317) );
  NAND U15388 ( .A(n14318), .B(n14317), .Z(n14336) );
  XOR U15389 ( .A(n14337), .B(n14336), .Z(c[1596]) );
  NANDN U15390 ( .A(n14320), .B(n14319), .Z(n14324) );
  OR U15391 ( .A(n14322), .B(n14321), .Z(n14323) );
  AND U15392 ( .A(n14324), .B(n14323), .Z(n14342) );
  XOR U15393 ( .A(a[575]), .B(n2258), .Z(n14346) );
  AND U15394 ( .A(a[577]), .B(b[0]), .Z(n14326) );
  XNOR U15395 ( .A(n14326), .B(n2175), .Z(n14328) );
  NANDN U15396 ( .A(b[0]), .B(a[576]), .Z(n14327) );
  NAND U15397 ( .A(n14328), .B(n14327), .Z(n14351) );
  AND U15398 ( .A(a[573]), .B(b[3]), .Z(n14350) );
  XOR U15399 ( .A(n14351), .B(n14350), .Z(n14353) );
  XOR U15400 ( .A(n14352), .B(n14353), .Z(n14341) );
  NANDN U15401 ( .A(n14330), .B(n14329), .Z(n14334) );
  OR U15402 ( .A(n14332), .B(n14331), .Z(n14333) );
  AND U15403 ( .A(n14334), .B(n14333), .Z(n14340) );
  XOR U15404 ( .A(n14341), .B(n14340), .Z(n14343) );
  XOR U15405 ( .A(n14342), .B(n14343), .Z(n14356) );
  XNOR U15406 ( .A(n14356), .B(sreg[1597]), .Z(n14358) );
  NANDN U15407 ( .A(n14335), .B(sreg[1596]), .Z(n14339) );
  NAND U15408 ( .A(n14337), .B(n14336), .Z(n14338) );
  NAND U15409 ( .A(n14339), .B(n14338), .Z(n14357) );
  XOR U15410 ( .A(n14358), .B(n14357), .Z(c[1597]) );
  NANDN U15411 ( .A(n14341), .B(n14340), .Z(n14345) );
  OR U15412 ( .A(n14343), .B(n14342), .Z(n14344) );
  AND U15413 ( .A(n14345), .B(n14344), .Z(n14363) );
  XOR U15414 ( .A(a[576]), .B(n2258), .Z(n14367) );
  AND U15415 ( .A(a[578]), .B(b[0]), .Z(n14347) );
  XNOR U15416 ( .A(n14347), .B(n2175), .Z(n14349) );
  NANDN U15417 ( .A(b[0]), .B(a[577]), .Z(n14348) );
  NAND U15418 ( .A(n14349), .B(n14348), .Z(n14372) );
  AND U15419 ( .A(a[574]), .B(b[3]), .Z(n14371) );
  XOR U15420 ( .A(n14372), .B(n14371), .Z(n14374) );
  XOR U15421 ( .A(n14373), .B(n14374), .Z(n14362) );
  NANDN U15422 ( .A(n14351), .B(n14350), .Z(n14355) );
  OR U15423 ( .A(n14353), .B(n14352), .Z(n14354) );
  AND U15424 ( .A(n14355), .B(n14354), .Z(n14361) );
  XOR U15425 ( .A(n14362), .B(n14361), .Z(n14364) );
  XOR U15426 ( .A(n14363), .B(n14364), .Z(n14377) );
  XNOR U15427 ( .A(n14377), .B(sreg[1598]), .Z(n14379) );
  NANDN U15428 ( .A(n14356), .B(sreg[1597]), .Z(n14360) );
  NAND U15429 ( .A(n14358), .B(n14357), .Z(n14359) );
  NAND U15430 ( .A(n14360), .B(n14359), .Z(n14378) );
  XOR U15431 ( .A(n14379), .B(n14378), .Z(c[1598]) );
  NANDN U15432 ( .A(n14362), .B(n14361), .Z(n14366) );
  OR U15433 ( .A(n14364), .B(n14363), .Z(n14365) );
  AND U15434 ( .A(n14366), .B(n14365), .Z(n14384) );
  XOR U15435 ( .A(a[577]), .B(n2258), .Z(n14388) );
  AND U15436 ( .A(a[579]), .B(b[0]), .Z(n14368) );
  XNOR U15437 ( .A(n14368), .B(n2175), .Z(n14370) );
  NANDN U15438 ( .A(b[0]), .B(a[578]), .Z(n14369) );
  NAND U15439 ( .A(n14370), .B(n14369), .Z(n14393) );
  AND U15440 ( .A(a[575]), .B(b[3]), .Z(n14392) );
  XOR U15441 ( .A(n14393), .B(n14392), .Z(n14395) );
  XOR U15442 ( .A(n14394), .B(n14395), .Z(n14383) );
  NANDN U15443 ( .A(n14372), .B(n14371), .Z(n14376) );
  OR U15444 ( .A(n14374), .B(n14373), .Z(n14375) );
  AND U15445 ( .A(n14376), .B(n14375), .Z(n14382) );
  XOR U15446 ( .A(n14383), .B(n14382), .Z(n14385) );
  XOR U15447 ( .A(n14384), .B(n14385), .Z(n14398) );
  XNOR U15448 ( .A(n14398), .B(sreg[1599]), .Z(n14400) );
  NANDN U15449 ( .A(n14377), .B(sreg[1598]), .Z(n14381) );
  NAND U15450 ( .A(n14379), .B(n14378), .Z(n14380) );
  NAND U15451 ( .A(n14381), .B(n14380), .Z(n14399) );
  XOR U15452 ( .A(n14400), .B(n14399), .Z(c[1599]) );
  NANDN U15453 ( .A(n14383), .B(n14382), .Z(n14387) );
  OR U15454 ( .A(n14385), .B(n14384), .Z(n14386) );
  AND U15455 ( .A(n14387), .B(n14386), .Z(n14405) );
  XOR U15456 ( .A(a[578]), .B(n2258), .Z(n14409) );
  AND U15457 ( .A(a[580]), .B(b[0]), .Z(n14389) );
  XNOR U15458 ( .A(n14389), .B(n2175), .Z(n14391) );
  NANDN U15459 ( .A(b[0]), .B(a[579]), .Z(n14390) );
  NAND U15460 ( .A(n14391), .B(n14390), .Z(n14414) );
  AND U15461 ( .A(a[576]), .B(b[3]), .Z(n14413) );
  XOR U15462 ( .A(n14414), .B(n14413), .Z(n14416) );
  XOR U15463 ( .A(n14415), .B(n14416), .Z(n14404) );
  NANDN U15464 ( .A(n14393), .B(n14392), .Z(n14397) );
  OR U15465 ( .A(n14395), .B(n14394), .Z(n14396) );
  AND U15466 ( .A(n14397), .B(n14396), .Z(n14403) );
  XOR U15467 ( .A(n14404), .B(n14403), .Z(n14406) );
  XOR U15468 ( .A(n14405), .B(n14406), .Z(n14419) );
  XNOR U15469 ( .A(n14419), .B(sreg[1600]), .Z(n14421) );
  NANDN U15470 ( .A(n14398), .B(sreg[1599]), .Z(n14402) );
  NAND U15471 ( .A(n14400), .B(n14399), .Z(n14401) );
  NAND U15472 ( .A(n14402), .B(n14401), .Z(n14420) );
  XOR U15473 ( .A(n14421), .B(n14420), .Z(c[1600]) );
  NANDN U15474 ( .A(n14404), .B(n14403), .Z(n14408) );
  OR U15475 ( .A(n14406), .B(n14405), .Z(n14407) );
  AND U15476 ( .A(n14408), .B(n14407), .Z(n14426) );
  XOR U15477 ( .A(a[579]), .B(n2258), .Z(n14430) );
  AND U15478 ( .A(a[581]), .B(b[0]), .Z(n14410) );
  XNOR U15479 ( .A(n14410), .B(n2175), .Z(n14412) );
  NANDN U15480 ( .A(b[0]), .B(a[580]), .Z(n14411) );
  NAND U15481 ( .A(n14412), .B(n14411), .Z(n14435) );
  AND U15482 ( .A(a[577]), .B(b[3]), .Z(n14434) );
  XOR U15483 ( .A(n14435), .B(n14434), .Z(n14437) );
  XOR U15484 ( .A(n14436), .B(n14437), .Z(n14425) );
  NANDN U15485 ( .A(n14414), .B(n14413), .Z(n14418) );
  OR U15486 ( .A(n14416), .B(n14415), .Z(n14417) );
  AND U15487 ( .A(n14418), .B(n14417), .Z(n14424) );
  XOR U15488 ( .A(n14425), .B(n14424), .Z(n14427) );
  XOR U15489 ( .A(n14426), .B(n14427), .Z(n14440) );
  XNOR U15490 ( .A(n14440), .B(sreg[1601]), .Z(n14442) );
  NANDN U15491 ( .A(n14419), .B(sreg[1600]), .Z(n14423) );
  NAND U15492 ( .A(n14421), .B(n14420), .Z(n14422) );
  NAND U15493 ( .A(n14423), .B(n14422), .Z(n14441) );
  XOR U15494 ( .A(n14442), .B(n14441), .Z(c[1601]) );
  NANDN U15495 ( .A(n14425), .B(n14424), .Z(n14429) );
  OR U15496 ( .A(n14427), .B(n14426), .Z(n14428) );
  AND U15497 ( .A(n14429), .B(n14428), .Z(n14447) );
  XOR U15498 ( .A(a[580]), .B(n2259), .Z(n14451) );
  AND U15499 ( .A(a[582]), .B(b[0]), .Z(n14431) );
  XNOR U15500 ( .A(n14431), .B(n2175), .Z(n14433) );
  NANDN U15501 ( .A(b[0]), .B(a[581]), .Z(n14432) );
  NAND U15502 ( .A(n14433), .B(n14432), .Z(n14456) );
  AND U15503 ( .A(a[578]), .B(b[3]), .Z(n14455) );
  XOR U15504 ( .A(n14456), .B(n14455), .Z(n14458) );
  XOR U15505 ( .A(n14457), .B(n14458), .Z(n14446) );
  NANDN U15506 ( .A(n14435), .B(n14434), .Z(n14439) );
  OR U15507 ( .A(n14437), .B(n14436), .Z(n14438) );
  AND U15508 ( .A(n14439), .B(n14438), .Z(n14445) );
  XOR U15509 ( .A(n14446), .B(n14445), .Z(n14448) );
  XOR U15510 ( .A(n14447), .B(n14448), .Z(n14461) );
  XNOR U15511 ( .A(n14461), .B(sreg[1602]), .Z(n14463) );
  NANDN U15512 ( .A(n14440), .B(sreg[1601]), .Z(n14444) );
  NAND U15513 ( .A(n14442), .B(n14441), .Z(n14443) );
  NAND U15514 ( .A(n14444), .B(n14443), .Z(n14462) );
  XOR U15515 ( .A(n14463), .B(n14462), .Z(c[1602]) );
  NANDN U15516 ( .A(n14446), .B(n14445), .Z(n14450) );
  OR U15517 ( .A(n14448), .B(n14447), .Z(n14449) );
  AND U15518 ( .A(n14450), .B(n14449), .Z(n14468) );
  XOR U15519 ( .A(a[581]), .B(n2259), .Z(n14472) );
  AND U15520 ( .A(a[579]), .B(b[3]), .Z(n14476) );
  AND U15521 ( .A(a[583]), .B(b[0]), .Z(n14452) );
  XNOR U15522 ( .A(n14452), .B(n2175), .Z(n14454) );
  NANDN U15523 ( .A(b[0]), .B(a[582]), .Z(n14453) );
  NAND U15524 ( .A(n14454), .B(n14453), .Z(n14477) );
  XOR U15525 ( .A(n14476), .B(n14477), .Z(n14479) );
  XOR U15526 ( .A(n14478), .B(n14479), .Z(n14467) );
  NANDN U15527 ( .A(n14456), .B(n14455), .Z(n14460) );
  OR U15528 ( .A(n14458), .B(n14457), .Z(n14459) );
  AND U15529 ( .A(n14460), .B(n14459), .Z(n14466) );
  XOR U15530 ( .A(n14467), .B(n14466), .Z(n14469) );
  XOR U15531 ( .A(n14468), .B(n14469), .Z(n14482) );
  XNOR U15532 ( .A(n14482), .B(sreg[1603]), .Z(n14484) );
  NANDN U15533 ( .A(n14461), .B(sreg[1602]), .Z(n14465) );
  NAND U15534 ( .A(n14463), .B(n14462), .Z(n14464) );
  NAND U15535 ( .A(n14465), .B(n14464), .Z(n14483) );
  XOR U15536 ( .A(n14484), .B(n14483), .Z(c[1603]) );
  NANDN U15537 ( .A(n14467), .B(n14466), .Z(n14471) );
  OR U15538 ( .A(n14469), .B(n14468), .Z(n14470) );
  AND U15539 ( .A(n14471), .B(n14470), .Z(n14489) );
  XOR U15540 ( .A(a[582]), .B(n2259), .Z(n14493) );
  AND U15541 ( .A(a[584]), .B(b[0]), .Z(n14473) );
  XNOR U15542 ( .A(n14473), .B(n2175), .Z(n14475) );
  NANDN U15543 ( .A(b[0]), .B(a[583]), .Z(n14474) );
  NAND U15544 ( .A(n14475), .B(n14474), .Z(n14498) );
  AND U15545 ( .A(a[580]), .B(b[3]), .Z(n14497) );
  XOR U15546 ( .A(n14498), .B(n14497), .Z(n14500) );
  XOR U15547 ( .A(n14499), .B(n14500), .Z(n14488) );
  NANDN U15548 ( .A(n14477), .B(n14476), .Z(n14481) );
  OR U15549 ( .A(n14479), .B(n14478), .Z(n14480) );
  AND U15550 ( .A(n14481), .B(n14480), .Z(n14487) );
  XOR U15551 ( .A(n14488), .B(n14487), .Z(n14490) );
  XOR U15552 ( .A(n14489), .B(n14490), .Z(n14503) );
  XNOR U15553 ( .A(n14503), .B(sreg[1604]), .Z(n14505) );
  NANDN U15554 ( .A(n14482), .B(sreg[1603]), .Z(n14486) );
  NAND U15555 ( .A(n14484), .B(n14483), .Z(n14485) );
  NAND U15556 ( .A(n14486), .B(n14485), .Z(n14504) );
  XOR U15557 ( .A(n14505), .B(n14504), .Z(c[1604]) );
  NANDN U15558 ( .A(n14488), .B(n14487), .Z(n14492) );
  OR U15559 ( .A(n14490), .B(n14489), .Z(n14491) );
  AND U15560 ( .A(n14492), .B(n14491), .Z(n14510) );
  XOR U15561 ( .A(a[583]), .B(n2259), .Z(n14514) );
  AND U15562 ( .A(a[581]), .B(b[3]), .Z(n14518) );
  AND U15563 ( .A(a[585]), .B(b[0]), .Z(n14494) );
  XNOR U15564 ( .A(n14494), .B(n2175), .Z(n14496) );
  NANDN U15565 ( .A(b[0]), .B(a[584]), .Z(n14495) );
  NAND U15566 ( .A(n14496), .B(n14495), .Z(n14519) );
  XOR U15567 ( .A(n14518), .B(n14519), .Z(n14521) );
  XOR U15568 ( .A(n14520), .B(n14521), .Z(n14509) );
  NANDN U15569 ( .A(n14498), .B(n14497), .Z(n14502) );
  OR U15570 ( .A(n14500), .B(n14499), .Z(n14501) );
  AND U15571 ( .A(n14502), .B(n14501), .Z(n14508) );
  XOR U15572 ( .A(n14509), .B(n14508), .Z(n14511) );
  XOR U15573 ( .A(n14510), .B(n14511), .Z(n14524) );
  XNOR U15574 ( .A(n14524), .B(sreg[1605]), .Z(n14526) );
  NANDN U15575 ( .A(n14503), .B(sreg[1604]), .Z(n14507) );
  NAND U15576 ( .A(n14505), .B(n14504), .Z(n14506) );
  NAND U15577 ( .A(n14507), .B(n14506), .Z(n14525) );
  XOR U15578 ( .A(n14526), .B(n14525), .Z(c[1605]) );
  NANDN U15579 ( .A(n14509), .B(n14508), .Z(n14513) );
  OR U15580 ( .A(n14511), .B(n14510), .Z(n14512) );
  AND U15581 ( .A(n14513), .B(n14512), .Z(n14531) );
  XOR U15582 ( .A(a[584]), .B(n2259), .Z(n14535) );
  AND U15583 ( .A(a[582]), .B(b[3]), .Z(n14539) );
  AND U15584 ( .A(a[586]), .B(b[0]), .Z(n14515) );
  XNOR U15585 ( .A(n14515), .B(n2175), .Z(n14517) );
  NANDN U15586 ( .A(b[0]), .B(a[585]), .Z(n14516) );
  NAND U15587 ( .A(n14517), .B(n14516), .Z(n14540) );
  XOR U15588 ( .A(n14539), .B(n14540), .Z(n14542) );
  XOR U15589 ( .A(n14541), .B(n14542), .Z(n14530) );
  NANDN U15590 ( .A(n14519), .B(n14518), .Z(n14523) );
  OR U15591 ( .A(n14521), .B(n14520), .Z(n14522) );
  AND U15592 ( .A(n14523), .B(n14522), .Z(n14529) );
  XOR U15593 ( .A(n14530), .B(n14529), .Z(n14532) );
  XOR U15594 ( .A(n14531), .B(n14532), .Z(n14545) );
  XNOR U15595 ( .A(n14545), .B(sreg[1606]), .Z(n14547) );
  NANDN U15596 ( .A(n14524), .B(sreg[1605]), .Z(n14528) );
  NAND U15597 ( .A(n14526), .B(n14525), .Z(n14527) );
  NAND U15598 ( .A(n14528), .B(n14527), .Z(n14546) );
  XOR U15599 ( .A(n14547), .B(n14546), .Z(c[1606]) );
  NANDN U15600 ( .A(n14530), .B(n14529), .Z(n14534) );
  OR U15601 ( .A(n14532), .B(n14531), .Z(n14533) );
  AND U15602 ( .A(n14534), .B(n14533), .Z(n14552) );
  XOR U15603 ( .A(a[585]), .B(n2259), .Z(n14556) );
  AND U15604 ( .A(a[587]), .B(b[0]), .Z(n14536) );
  XNOR U15605 ( .A(n14536), .B(n2175), .Z(n14538) );
  NANDN U15606 ( .A(b[0]), .B(a[586]), .Z(n14537) );
  NAND U15607 ( .A(n14538), .B(n14537), .Z(n14561) );
  AND U15608 ( .A(a[583]), .B(b[3]), .Z(n14560) );
  XOR U15609 ( .A(n14561), .B(n14560), .Z(n14563) );
  XOR U15610 ( .A(n14562), .B(n14563), .Z(n14551) );
  NANDN U15611 ( .A(n14540), .B(n14539), .Z(n14544) );
  OR U15612 ( .A(n14542), .B(n14541), .Z(n14543) );
  AND U15613 ( .A(n14544), .B(n14543), .Z(n14550) );
  XOR U15614 ( .A(n14551), .B(n14550), .Z(n14553) );
  XOR U15615 ( .A(n14552), .B(n14553), .Z(n14566) );
  XNOR U15616 ( .A(n14566), .B(sreg[1607]), .Z(n14568) );
  NANDN U15617 ( .A(n14545), .B(sreg[1606]), .Z(n14549) );
  NAND U15618 ( .A(n14547), .B(n14546), .Z(n14548) );
  NAND U15619 ( .A(n14549), .B(n14548), .Z(n14567) );
  XOR U15620 ( .A(n14568), .B(n14567), .Z(c[1607]) );
  NANDN U15621 ( .A(n14551), .B(n14550), .Z(n14555) );
  OR U15622 ( .A(n14553), .B(n14552), .Z(n14554) );
  AND U15623 ( .A(n14555), .B(n14554), .Z(n14573) );
  XOR U15624 ( .A(a[586]), .B(n2259), .Z(n14577) );
  AND U15625 ( .A(a[588]), .B(b[0]), .Z(n14557) );
  XNOR U15626 ( .A(n14557), .B(n2175), .Z(n14559) );
  NANDN U15627 ( .A(b[0]), .B(a[587]), .Z(n14558) );
  NAND U15628 ( .A(n14559), .B(n14558), .Z(n14582) );
  AND U15629 ( .A(a[584]), .B(b[3]), .Z(n14581) );
  XOR U15630 ( .A(n14582), .B(n14581), .Z(n14584) );
  XOR U15631 ( .A(n14583), .B(n14584), .Z(n14572) );
  NANDN U15632 ( .A(n14561), .B(n14560), .Z(n14565) );
  OR U15633 ( .A(n14563), .B(n14562), .Z(n14564) );
  AND U15634 ( .A(n14565), .B(n14564), .Z(n14571) );
  XOR U15635 ( .A(n14572), .B(n14571), .Z(n14574) );
  XOR U15636 ( .A(n14573), .B(n14574), .Z(n14587) );
  XNOR U15637 ( .A(n14587), .B(sreg[1608]), .Z(n14589) );
  NANDN U15638 ( .A(n14566), .B(sreg[1607]), .Z(n14570) );
  NAND U15639 ( .A(n14568), .B(n14567), .Z(n14569) );
  NAND U15640 ( .A(n14570), .B(n14569), .Z(n14588) );
  XOR U15641 ( .A(n14589), .B(n14588), .Z(c[1608]) );
  NANDN U15642 ( .A(n14572), .B(n14571), .Z(n14576) );
  OR U15643 ( .A(n14574), .B(n14573), .Z(n14575) );
  AND U15644 ( .A(n14576), .B(n14575), .Z(n14594) );
  XOR U15645 ( .A(a[587]), .B(n2260), .Z(n14598) );
  AND U15646 ( .A(a[589]), .B(b[0]), .Z(n14578) );
  XNOR U15647 ( .A(n14578), .B(n2175), .Z(n14580) );
  NANDN U15648 ( .A(b[0]), .B(a[588]), .Z(n14579) );
  NAND U15649 ( .A(n14580), .B(n14579), .Z(n14603) );
  AND U15650 ( .A(a[585]), .B(b[3]), .Z(n14602) );
  XOR U15651 ( .A(n14603), .B(n14602), .Z(n14605) );
  XOR U15652 ( .A(n14604), .B(n14605), .Z(n14593) );
  NANDN U15653 ( .A(n14582), .B(n14581), .Z(n14586) );
  OR U15654 ( .A(n14584), .B(n14583), .Z(n14585) );
  AND U15655 ( .A(n14586), .B(n14585), .Z(n14592) );
  XOR U15656 ( .A(n14593), .B(n14592), .Z(n14595) );
  XOR U15657 ( .A(n14594), .B(n14595), .Z(n14608) );
  XNOR U15658 ( .A(n14608), .B(sreg[1609]), .Z(n14610) );
  NANDN U15659 ( .A(n14587), .B(sreg[1608]), .Z(n14591) );
  NAND U15660 ( .A(n14589), .B(n14588), .Z(n14590) );
  NAND U15661 ( .A(n14591), .B(n14590), .Z(n14609) );
  XOR U15662 ( .A(n14610), .B(n14609), .Z(c[1609]) );
  NANDN U15663 ( .A(n14593), .B(n14592), .Z(n14597) );
  OR U15664 ( .A(n14595), .B(n14594), .Z(n14596) );
  AND U15665 ( .A(n14597), .B(n14596), .Z(n14615) );
  XOR U15666 ( .A(a[588]), .B(n2260), .Z(n14619) );
  AND U15667 ( .A(a[586]), .B(b[3]), .Z(n14623) );
  AND U15668 ( .A(a[590]), .B(b[0]), .Z(n14599) );
  XNOR U15669 ( .A(n14599), .B(n2175), .Z(n14601) );
  NANDN U15670 ( .A(b[0]), .B(a[589]), .Z(n14600) );
  NAND U15671 ( .A(n14601), .B(n14600), .Z(n14624) );
  XOR U15672 ( .A(n14623), .B(n14624), .Z(n14626) );
  XOR U15673 ( .A(n14625), .B(n14626), .Z(n14614) );
  NANDN U15674 ( .A(n14603), .B(n14602), .Z(n14607) );
  OR U15675 ( .A(n14605), .B(n14604), .Z(n14606) );
  AND U15676 ( .A(n14607), .B(n14606), .Z(n14613) );
  XOR U15677 ( .A(n14614), .B(n14613), .Z(n14616) );
  XOR U15678 ( .A(n14615), .B(n14616), .Z(n14629) );
  XNOR U15679 ( .A(n14629), .B(sreg[1610]), .Z(n14631) );
  NANDN U15680 ( .A(n14608), .B(sreg[1609]), .Z(n14612) );
  NAND U15681 ( .A(n14610), .B(n14609), .Z(n14611) );
  NAND U15682 ( .A(n14612), .B(n14611), .Z(n14630) );
  XOR U15683 ( .A(n14631), .B(n14630), .Z(c[1610]) );
  NANDN U15684 ( .A(n14614), .B(n14613), .Z(n14618) );
  OR U15685 ( .A(n14616), .B(n14615), .Z(n14617) );
  AND U15686 ( .A(n14618), .B(n14617), .Z(n14636) );
  XOR U15687 ( .A(a[589]), .B(n2260), .Z(n14640) );
  AND U15688 ( .A(a[591]), .B(b[0]), .Z(n14620) );
  XNOR U15689 ( .A(n14620), .B(n2175), .Z(n14622) );
  NANDN U15690 ( .A(b[0]), .B(a[590]), .Z(n14621) );
  NAND U15691 ( .A(n14622), .B(n14621), .Z(n14645) );
  AND U15692 ( .A(a[587]), .B(b[3]), .Z(n14644) );
  XOR U15693 ( .A(n14645), .B(n14644), .Z(n14647) );
  XOR U15694 ( .A(n14646), .B(n14647), .Z(n14635) );
  NANDN U15695 ( .A(n14624), .B(n14623), .Z(n14628) );
  OR U15696 ( .A(n14626), .B(n14625), .Z(n14627) );
  AND U15697 ( .A(n14628), .B(n14627), .Z(n14634) );
  XOR U15698 ( .A(n14635), .B(n14634), .Z(n14637) );
  XOR U15699 ( .A(n14636), .B(n14637), .Z(n14650) );
  XNOR U15700 ( .A(n14650), .B(sreg[1611]), .Z(n14652) );
  NANDN U15701 ( .A(n14629), .B(sreg[1610]), .Z(n14633) );
  NAND U15702 ( .A(n14631), .B(n14630), .Z(n14632) );
  NAND U15703 ( .A(n14633), .B(n14632), .Z(n14651) );
  XOR U15704 ( .A(n14652), .B(n14651), .Z(c[1611]) );
  NANDN U15705 ( .A(n14635), .B(n14634), .Z(n14639) );
  OR U15706 ( .A(n14637), .B(n14636), .Z(n14638) );
  AND U15707 ( .A(n14639), .B(n14638), .Z(n14657) );
  XOR U15708 ( .A(a[590]), .B(n2260), .Z(n14661) );
  AND U15709 ( .A(a[592]), .B(b[0]), .Z(n14641) );
  XNOR U15710 ( .A(n14641), .B(n2175), .Z(n14643) );
  NANDN U15711 ( .A(b[0]), .B(a[591]), .Z(n14642) );
  NAND U15712 ( .A(n14643), .B(n14642), .Z(n14666) );
  AND U15713 ( .A(a[588]), .B(b[3]), .Z(n14665) );
  XOR U15714 ( .A(n14666), .B(n14665), .Z(n14668) );
  XOR U15715 ( .A(n14667), .B(n14668), .Z(n14656) );
  NANDN U15716 ( .A(n14645), .B(n14644), .Z(n14649) );
  OR U15717 ( .A(n14647), .B(n14646), .Z(n14648) );
  AND U15718 ( .A(n14649), .B(n14648), .Z(n14655) );
  XOR U15719 ( .A(n14656), .B(n14655), .Z(n14658) );
  XOR U15720 ( .A(n14657), .B(n14658), .Z(n14671) );
  XNOR U15721 ( .A(n14671), .B(sreg[1612]), .Z(n14673) );
  NANDN U15722 ( .A(n14650), .B(sreg[1611]), .Z(n14654) );
  NAND U15723 ( .A(n14652), .B(n14651), .Z(n14653) );
  NAND U15724 ( .A(n14654), .B(n14653), .Z(n14672) );
  XOR U15725 ( .A(n14673), .B(n14672), .Z(c[1612]) );
  NANDN U15726 ( .A(n14656), .B(n14655), .Z(n14660) );
  OR U15727 ( .A(n14658), .B(n14657), .Z(n14659) );
  AND U15728 ( .A(n14660), .B(n14659), .Z(n14678) );
  XOR U15729 ( .A(a[591]), .B(n2260), .Z(n14682) );
  AND U15730 ( .A(a[589]), .B(b[3]), .Z(n14686) );
  AND U15731 ( .A(a[593]), .B(b[0]), .Z(n14662) );
  XNOR U15732 ( .A(n14662), .B(n2175), .Z(n14664) );
  NANDN U15733 ( .A(b[0]), .B(a[592]), .Z(n14663) );
  NAND U15734 ( .A(n14664), .B(n14663), .Z(n14687) );
  XOR U15735 ( .A(n14686), .B(n14687), .Z(n14689) );
  XOR U15736 ( .A(n14688), .B(n14689), .Z(n14677) );
  NANDN U15737 ( .A(n14666), .B(n14665), .Z(n14670) );
  OR U15738 ( .A(n14668), .B(n14667), .Z(n14669) );
  AND U15739 ( .A(n14670), .B(n14669), .Z(n14676) );
  XOR U15740 ( .A(n14677), .B(n14676), .Z(n14679) );
  XOR U15741 ( .A(n14678), .B(n14679), .Z(n14692) );
  XNOR U15742 ( .A(n14692), .B(sreg[1613]), .Z(n14694) );
  NANDN U15743 ( .A(n14671), .B(sreg[1612]), .Z(n14675) );
  NAND U15744 ( .A(n14673), .B(n14672), .Z(n14674) );
  NAND U15745 ( .A(n14675), .B(n14674), .Z(n14693) );
  XOR U15746 ( .A(n14694), .B(n14693), .Z(c[1613]) );
  NANDN U15747 ( .A(n14677), .B(n14676), .Z(n14681) );
  OR U15748 ( .A(n14679), .B(n14678), .Z(n14680) );
  AND U15749 ( .A(n14681), .B(n14680), .Z(n14699) );
  XOR U15750 ( .A(a[592]), .B(n2260), .Z(n14703) );
  AND U15751 ( .A(a[590]), .B(b[3]), .Z(n14707) );
  AND U15752 ( .A(a[594]), .B(b[0]), .Z(n14683) );
  XNOR U15753 ( .A(n14683), .B(n2175), .Z(n14685) );
  NANDN U15754 ( .A(b[0]), .B(a[593]), .Z(n14684) );
  NAND U15755 ( .A(n14685), .B(n14684), .Z(n14708) );
  XOR U15756 ( .A(n14707), .B(n14708), .Z(n14710) );
  XOR U15757 ( .A(n14709), .B(n14710), .Z(n14698) );
  NANDN U15758 ( .A(n14687), .B(n14686), .Z(n14691) );
  OR U15759 ( .A(n14689), .B(n14688), .Z(n14690) );
  AND U15760 ( .A(n14691), .B(n14690), .Z(n14697) );
  XOR U15761 ( .A(n14698), .B(n14697), .Z(n14700) );
  XOR U15762 ( .A(n14699), .B(n14700), .Z(n14713) );
  XNOR U15763 ( .A(n14713), .B(sreg[1614]), .Z(n14715) );
  NANDN U15764 ( .A(n14692), .B(sreg[1613]), .Z(n14696) );
  NAND U15765 ( .A(n14694), .B(n14693), .Z(n14695) );
  NAND U15766 ( .A(n14696), .B(n14695), .Z(n14714) );
  XOR U15767 ( .A(n14715), .B(n14714), .Z(c[1614]) );
  NANDN U15768 ( .A(n14698), .B(n14697), .Z(n14702) );
  OR U15769 ( .A(n14700), .B(n14699), .Z(n14701) );
  AND U15770 ( .A(n14702), .B(n14701), .Z(n14720) );
  XOR U15771 ( .A(a[593]), .B(n2260), .Z(n14724) );
  AND U15772 ( .A(a[595]), .B(b[0]), .Z(n14704) );
  XNOR U15773 ( .A(n14704), .B(n2175), .Z(n14706) );
  NANDN U15774 ( .A(b[0]), .B(a[594]), .Z(n14705) );
  NAND U15775 ( .A(n14706), .B(n14705), .Z(n14729) );
  AND U15776 ( .A(a[591]), .B(b[3]), .Z(n14728) );
  XOR U15777 ( .A(n14729), .B(n14728), .Z(n14731) );
  XOR U15778 ( .A(n14730), .B(n14731), .Z(n14719) );
  NANDN U15779 ( .A(n14708), .B(n14707), .Z(n14712) );
  OR U15780 ( .A(n14710), .B(n14709), .Z(n14711) );
  AND U15781 ( .A(n14712), .B(n14711), .Z(n14718) );
  XOR U15782 ( .A(n14719), .B(n14718), .Z(n14721) );
  XOR U15783 ( .A(n14720), .B(n14721), .Z(n14734) );
  XNOR U15784 ( .A(n14734), .B(sreg[1615]), .Z(n14736) );
  NANDN U15785 ( .A(n14713), .B(sreg[1614]), .Z(n14717) );
  NAND U15786 ( .A(n14715), .B(n14714), .Z(n14716) );
  NAND U15787 ( .A(n14717), .B(n14716), .Z(n14735) );
  XOR U15788 ( .A(n14736), .B(n14735), .Z(c[1615]) );
  NANDN U15789 ( .A(n14719), .B(n14718), .Z(n14723) );
  OR U15790 ( .A(n14721), .B(n14720), .Z(n14722) );
  AND U15791 ( .A(n14723), .B(n14722), .Z(n14741) );
  XOR U15792 ( .A(a[594]), .B(n2261), .Z(n14745) );
  AND U15793 ( .A(a[596]), .B(b[0]), .Z(n14725) );
  XNOR U15794 ( .A(n14725), .B(n2175), .Z(n14727) );
  NANDN U15795 ( .A(b[0]), .B(a[595]), .Z(n14726) );
  NAND U15796 ( .A(n14727), .B(n14726), .Z(n14750) );
  AND U15797 ( .A(a[592]), .B(b[3]), .Z(n14749) );
  XOR U15798 ( .A(n14750), .B(n14749), .Z(n14752) );
  XOR U15799 ( .A(n14751), .B(n14752), .Z(n14740) );
  NANDN U15800 ( .A(n14729), .B(n14728), .Z(n14733) );
  OR U15801 ( .A(n14731), .B(n14730), .Z(n14732) );
  AND U15802 ( .A(n14733), .B(n14732), .Z(n14739) );
  XOR U15803 ( .A(n14740), .B(n14739), .Z(n14742) );
  XOR U15804 ( .A(n14741), .B(n14742), .Z(n14755) );
  XNOR U15805 ( .A(n14755), .B(sreg[1616]), .Z(n14757) );
  NANDN U15806 ( .A(n14734), .B(sreg[1615]), .Z(n14738) );
  NAND U15807 ( .A(n14736), .B(n14735), .Z(n14737) );
  NAND U15808 ( .A(n14738), .B(n14737), .Z(n14756) );
  XOR U15809 ( .A(n14757), .B(n14756), .Z(c[1616]) );
  NANDN U15810 ( .A(n14740), .B(n14739), .Z(n14744) );
  OR U15811 ( .A(n14742), .B(n14741), .Z(n14743) );
  AND U15812 ( .A(n14744), .B(n14743), .Z(n14763) );
  XOR U15813 ( .A(a[595]), .B(n2261), .Z(n14764) );
  AND U15814 ( .A(b[0]), .B(a[597]), .Z(n14746) );
  XOR U15815 ( .A(b[1]), .B(n14746), .Z(n14748) );
  NANDN U15816 ( .A(b[0]), .B(a[596]), .Z(n14747) );
  AND U15817 ( .A(n14748), .B(n14747), .Z(n14768) );
  AND U15818 ( .A(a[593]), .B(b[3]), .Z(n14769) );
  XOR U15819 ( .A(n14768), .B(n14769), .Z(n14770) );
  XNOR U15820 ( .A(n14771), .B(n14770), .Z(n14760) );
  NANDN U15821 ( .A(n14750), .B(n14749), .Z(n14754) );
  OR U15822 ( .A(n14752), .B(n14751), .Z(n14753) );
  AND U15823 ( .A(n14754), .B(n14753), .Z(n14761) );
  XNOR U15824 ( .A(n14760), .B(n14761), .Z(n14762) );
  XNOR U15825 ( .A(n14763), .B(n14762), .Z(n14774) );
  XNOR U15826 ( .A(n14774), .B(sreg[1617]), .Z(n14776) );
  NANDN U15827 ( .A(n14755), .B(sreg[1616]), .Z(n14759) );
  NAND U15828 ( .A(n14757), .B(n14756), .Z(n14758) );
  NAND U15829 ( .A(n14759), .B(n14758), .Z(n14775) );
  XOR U15830 ( .A(n14776), .B(n14775), .Z(c[1617]) );
  XOR U15831 ( .A(a[596]), .B(n2261), .Z(n14783) );
  AND U15832 ( .A(a[598]), .B(b[0]), .Z(n14765) );
  XNOR U15833 ( .A(n14765), .B(n2175), .Z(n14767) );
  NANDN U15834 ( .A(b[0]), .B(a[597]), .Z(n14766) );
  NAND U15835 ( .A(n14767), .B(n14766), .Z(n14788) );
  AND U15836 ( .A(a[594]), .B(b[3]), .Z(n14787) );
  XOR U15837 ( .A(n14788), .B(n14787), .Z(n14790) );
  XOR U15838 ( .A(n14789), .B(n14790), .Z(n14778) );
  NAND U15839 ( .A(n14769), .B(n14768), .Z(n14773) );
  NANDN U15840 ( .A(n14771), .B(n14770), .Z(n14772) );
  AND U15841 ( .A(n14773), .B(n14772), .Z(n14777) );
  XOR U15842 ( .A(n14778), .B(n14777), .Z(n14780) );
  XOR U15843 ( .A(n14779), .B(n14780), .Z(n14793) );
  XNOR U15844 ( .A(n14793), .B(sreg[1618]), .Z(n14795) );
  XOR U15845 ( .A(n14795), .B(n14794), .Z(c[1618]) );
  NANDN U15846 ( .A(n14778), .B(n14777), .Z(n14782) );
  OR U15847 ( .A(n14780), .B(n14779), .Z(n14781) );
  AND U15848 ( .A(n14782), .B(n14781), .Z(n14800) );
  XOR U15849 ( .A(a[597]), .B(n2261), .Z(n14804) );
  AND U15850 ( .A(a[599]), .B(b[0]), .Z(n14784) );
  XNOR U15851 ( .A(n14784), .B(n2175), .Z(n14786) );
  NANDN U15852 ( .A(b[0]), .B(a[598]), .Z(n14785) );
  NAND U15853 ( .A(n14786), .B(n14785), .Z(n14809) );
  AND U15854 ( .A(a[595]), .B(b[3]), .Z(n14808) );
  XOR U15855 ( .A(n14809), .B(n14808), .Z(n14811) );
  XOR U15856 ( .A(n14810), .B(n14811), .Z(n14799) );
  NANDN U15857 ( .A(n14788), .B(n14787), .Z(n14792) );
  OR U15858 ( .A(n14790), .B(n14789), .Z(n14791) );
  AND U15859 ( .A(n14792), .B(n14791), .Z(n14798) );
  XOR U15860 ( .A(n14799), .B(n14798), .Z(n14801) );
  XOR U15861 ( .A(n14800), .B(n14801), .Z(n14814) );
  XNOR U15862 ( .A(n14814), .B(sreg[1619]), .Z(n14816) );
  NANDN U15863 ( .A(n14793), .B(sreg[1618]), .Z(n14797) );
  NAND U15864 ( .A(n14795), .B(n14794), .Z(n14796) );
  NAND U15865 ( .A(n14797), .B(n14796), .Z(n14815) );
  XOR U15866 ( .A(n14816), .B(n14815), .Z(c[1619]) );
  NANDN U15867 ( .A(n14799), .B(n14798), .Z(n14803) );
  OR U15868 ( .A(n14801), .B(n14800), .Z(n14802) );
  AND U15869 ( .A(n14803), .B(n14802), .Z(n14821) );
  XOR U15870 ( .A(a[598]), .B(n2261), .Z(n14825) );
  AND U15871 ( .A(a[600]), .B(b[0]), .Z(n14805) );
  XNOR U15872 ( .A(n14805), .B(n2175), .Z(n14807) );
  NANDN U15873 ( .A(b[0]), .B(a[599]), .Z(n14806) );
  NAND U15874 ( .A(n14807), .B(n14806), .Z(n14830) );
  AND U15875 ( .A(a[596]), .B(b[3]), .Z(n14829) );
  XOR U15876 ( .A(n14830), .B(n14829), .Z(n14832) );
  XOR U15877 ( .A(n14831), .B(n14832), .Z(n14820) );
  NANDN U15878 ( .A(n14809), .B(n14808), .Z(n14813) );
  OR U15879 ( .A(n14811), .B(n14810), .Z(n14812) );
  AND U15880 ( .A(n14813), .B(n14812), .Z(n14819) );
  XOR U15881 ( .A(n14820), .B(n14819), .Z(n14822) );
  XOR U15882 ( .A(n14821), .B(n14822), .Z(n14835) );
  XNOR U15883 ( .A(n14835), .B(sreg[1620]), .Z(n14837) );
  NANDN U15884 ( .A(n14814), .B(sreg[1619]), .Z(n14818) );
  NAND U15885 ( .A(n14816), .B(n14815), .Z(n14817) );
  NAND U15886 ( .A(n14818), .B(n14817), .Z(n14836) );
  XOR U15887 ( .A(n14837), .B(n14836), .Z(c[1620]) );
  NANDN U15888 ( .A(n14820), .B(n14819), .Z(n14824) );
  OR U15889 ( .A(n14822), .B(n14821), .Z(n14823) );
  AND U15890 ( .A(n14824), .B(n14823), .Z(n14842) );
  XOR U15891 ( .A(a[599]), .B(n2261), .Z(n14846) );
  AND U15892 ( .A(a[601]), .B(b[0]), .Z(n14826) );
  XNOR U15893 ( .A(n14826), .B(n2175), .Z(n14828) );
  NANDN U15894 ( .A(b[0]), .B(a[600]), .Z(n14827) );
  NAND U15895 ( .A(n14828), .B(n14827), .Z(n14851) );
  AND U15896 ( .A(a[597]), .B(b[3]), .Z(n14850) );
  XOR U15897 ( .A(n14851), .B(n14850), .Z(n14853) );
  XOR U15898 ( .A(n14852), .B(n14853), .Z(n14841) );
  NANDN U15899 ( .A(n14830), .B(n14829), .Z(n14834) );
  OR U15900 ( .A(n14832), .B(n14831), .Z(n14833) );
  AND U15901 ( .A(n14834), .B(n14833), .Z(n14840) );
  XOR U15902 ( .A(n14841), .B(n14840), .Z(n14843) );
  XOR U15903 ( .A(n14842), .B(n14843), .Z(n14856) );
  XNOR U15904 ( .A(n14856), .B(sreg[1621]), .Z(n14858) );
  NANDN U15905 ( .A(n14835), .B(sreg[1620]), .Z(n14839) );
  NAND U15906 ( .A(n14837), .B(n14836), .Z(n14838) );
  NAND U15907 ( .A(n14839), .B(n14838), .Z(n14857) );
  XOR U15908 ( .A(n14858), .B(n14857), .Z(c[1621]) );
  NANDN U15909 ( .A(n14841), .B(n14840), .Z(n14845) );
  OR U15910 ( .A(n14843), .B(n14842), .Z(n14844) );
  AND U15911 ( .A(n14845), .B(n14844), .Z(n14863) );
  XOR U15912 ( .A(a[600]), .B(n2261), .Z(n14867) );
  AND U15913 ( .A(a[602]), .B(b[0]), .Z(n14847) );
  XNOR U15914 ( .A(n14847), .B(n2175), .Z(n14849) );
  NANDN U15915 ( .A(b[0]), .B(a[601]), .Z(n14848) );
  NAND U15916 ( .A(n14849), .B(n14848), .Z(n14872) );
  AND U15917 ( .A(a[598]), .B(b[3]), .Z(n14871) );
  XOR U15918 ( .A(n14872), .B(n14871), .Z(n14874) );
  XOR U15919 ( .A(n14873), .B(n14874), .Z(n14862) );
  NANDN U15920 ( .A(n14851), .B(n14850), .Z(n14855) );
  OR U15921 ( .A(n14853), .B(n14852), .Z(n14854) );
  AND U15922 ( .A(n14855), .B(n14854), .Z(n14861) );
  XOR U15923 ( .A(n14862), .B(n14861), .Z(n14864) );
  XOR U15924 ( .A(n14863), .B(n14864), .Z(n14877) );
  XNOR U15925 ( .A(n14877), .B(sreg[1622]), .Z(n14879) );
  NANDN U15926 ( .A(n14856), .B(sreg[1621]), .Z(n14860) );
  NAND U15927 ( .A(n14858), .B(n14857), .Z(n14859) );
  NAND U15928 ( .A(n14860), .B(n14859), .Z(n14878) );
  XOR U15929 ( .A(n14879), .B(n14878), .Z(c[1622]) );
  NANDN U15930 ( .A(n14862), .B(n14861), .Z(n14866) );
  OR U15931 ( .A(n14864), .B(n14863), .Z(n14865) );
  AND U15932 ( .A(n14866), .B(n14865), .Z(n14884) );
  XOR U15933 ( .A(a[601]), .B(n2262), .Z(n14888) );
  AND U15934 ( .A(a[603]), .B(b[0]), .Z(n14868) );
  XNOR U15935 ( .A(n14868), .B(n2175), .Z(n14870) );
  NANDN U15936 ( .A(b[0]), .B(a[602]), .Z(n14869) );
  NAND U15937 ( .A(n14870), .B(n14869), .Z(n14893) );
  AND U15938 ( .A(a[599]), .B(b[3]), .Z(n14892) );
  XOR U15939 ( .A(n14893), .B(n14892), .Z(n14895) );
  XOR U15940 ( .A(n14894), .B(n14895), .Z(n14883) );
  NANDN U15941 ( .A(n14872), .B(n14871), .Z(n14876) );
  OR U15942 ( .A(n14874), .B(n14873), .Z(n14875) );
  AND U15943 ( .A(n14876), .B(n14875), .Z(n14882) );
  XOR U15944 ( .A(n14883), .B(n14882), .Z(n14885) );
  XOR U15945 ( .A(n14884), .B(n14885), .Z(n14898) );
  XNOR U15946 ( .A(n14898), .B(sreg[1623]), .Z(n14900) );
  NANDN U15947 ( .A(n14877), .B(sreg[1622]), .Z(n14881) );
  NAND U15948 ( .A(n14879), .B(n14878), .Z(n14880) );
  NAND U15949 ( .A(n14881), .B(n14880), .Z(n14899) );
  XOR U15950 ( .A(n14900), .B(n14899), .Z(c[1623]) );
  NANDN U15951 ( .A(n14883), .B(n14882), .Z(n14887) );
  OR U15952 ( .A(n14885), .B(n14884), .Z(n14886) );
  AND U15953 ( .A(n14887), .B(n14886), .Z(n14905) );
  XOR U15954 ( .A(a[602]), .B(n2262), .Z(n14909) );
  AND U15955 ( .A(a[600]), .B(b[3]), .Z(n14913) );
  AND U15956 ( .A(a[604]), .B(b[0]), .Z(n14889) );
  XNOR U15957 ( .A(n14889), .B(n2175), .Z(n14891) );
  NANDN U15958 ( .A(b[0]), .B(a[603]), .Z(n14890) );
  NAND U15959 ( .A(n14891), .B(n14890), .Z(n14914) );
  XOR U15960 ( .A(n14913), .B(n14914), .Z(n14916) );
  XOR U15961 ( .A(n14915), .B(n14916), .Z(n14904) );
  NANDN U15962 ( .A(n14893), .B(n14892), .Z(n14897) );
  OR U15963 ( .A(n14895), .B(n14894), .Z(n14896) );
  AND U15964 ( .A(n14897), .B(n14896), .Z(n14903) );
  XOR U15965 ( .A(n14904), .B(n14903), .Z(n14906) );
  XOR U15966 ( .A(n14905), .B(n14906), .Z(n14919) );
  XNOR U15967 ( .A(n14919), .B(sreg[1624]), .Z(n14921) );
  NANDN U15968 ( .A(n14898), .B(sreg[1623]), .Z(n14902) );
  NAND U15969 ( .A(n14900), .B(n14899), .Z(n14901) );
  NAND U15970 ( .A(n14902), .B(n14901), .Z(n14920) );
  XOR U15971 ( .A(n14921), .B(n14920), .Z(c[1624]) );
  NANDN U15972 ( .A(n14904), .B(n14903), .Z(n14908) );
  OR U15973 ( .A(n14906), .B(n14905), .Z(n14907) );
  AND U15974 ( .A(n14908), .B(n14907), .Z(n14926) );
  XOR U15975 ( .A(a[603]), .B(n2262), .Z(n14930) );
  AND U15976 ( .A(a[605]), .B(b[0]), .Z(n14910) );
  XNOR U15977 ( .A(n14910), .B(n2175), .Z(n14912) );
  NANDN U15978 ( .A(b[0]), .B(a[604]), .Z(n14911) );
  NAND U15979 ( .A(n14912), .B(n14911), .Z(n14935) );
  AND U15980 ( .A(a[601]), .B(b[3]), .Z(n14934) );
  XOR U15981 ( .A(n14935), .B(n14934), .Z(n14937) );
  XOR U15982 ( .A(n14936), .B(n14937), .Z(n14925) );
  NANDN U15983 ( .A(n14914), .B(n14913), .Z(n14918) );
  OR U15984 ( .A(n14916), .B(n14915), .Z(n14917) );
  AND U15985 ( .A(n14918), .B(n14917), .Z(n14924) );
  XOR U15986 ( .A(n14925), .B(n14924), .Z(n14927) );
  XOR U15987 ( .A(n14926), .B(n14927), .Z(n14940) );
  XNOR U15988 ( .A(n14940), .B(sreg[1625]), .Z(n14942) );
  NANDN U15989 ( .A(n14919), .B(sreg[1624]), .Z(n14923) );
  NAND U15990 ( .A(n14921), .B(n14920), .Z(n14922) );
  NAND U15991 ( .A(n14923), .B(n14922), .Z(n14941) );
  XOR U15992 ( .A(n14942), .B(n14941), .Z(c[1625]) );
  NANDN U15993 ( .A(n14925), .B(n14924), .Z(n14929) );
  OR U15994 ( .A(n14927), .B(n14926), .Z(n14928) );
  AND U15995 ( .A(n14929), .B(n14928), .Z(n14947) );
  XOR U15996 ( .A(a[604]), .B(n2262), .Z(n14951) );
  AND U15997 ( .A(a[606]), .B(b[0]), .Z(n14931) );
  XNOR U15998 ( .A(n14931), .B(n2175), .Z(n14933) );
  NANDN U15999 ( .A(b[0]), .B(a[605]), .Z(n14932) );
  NAND U16000 ( .A(n14933), .B(n14932), .Z(n14956) );
  AND U16001 ( .A(a[602]), .B(b[3]), .Z(n14955) );
  XOR U16002 ( .A(n14956), .B(n14955), .Z(n14958) );
  XOR U16003 ( .A(n14957), .B(n14958), .Z(n14946) );
  NANDN U16004 ( .A(n14935), .B(n14934), .Z(n14939) );
  OR U16005 ( .A(n14937), .B(n14936), .Z(n14938) );
  AND U16006 ( .A(n14939), .B(n14938), .Z(n14945) );
  XOR U16007 ( .A(n14946), .B(n14945), .Z(n14948) );
  XOR U16008 ( .A(n14947), .B(n14948), .Z(n14961) );
  XNOR U16009 ( .A(n14961), .B(sreg[1626]), .Z(n14963) );
  NANDN U16010 ( .A(n14940), .B(sreg[1625]), .Z(n14944) );
  NAND U16011 ( .A(n14942), .B(n14941), .Z(n14943) );
  NAND U16012 ( .A(n14944), .B(n14943), .Z(n14962) );
  XOR U16013 ( .A(n14963), .B(n14962), .Z(c[1626]) );
  NANDN U16014 ( .A(n14946), .B(n14945), .Z(n14950) );
  OR U16015 ( .A(n14948), .B(n14947), .Z(n14949) );
  AND U16016 ( .A(n14950), .B(n14949), .Z(n14968) );
  XOR U16017 ( .A(a[605]), .B(n2262), .Z(n14972) );
  AND U16018 ( .A(a[607]), .B(b[0]), .Z(n14952) );
  XNOR U16019 ( .A(n14952), .B(n2175), .Z(n14954) );
  NANDN U16020 ( .A(b[0]), .B(a[606]), .Z(n14953) );
  NAND U16021 ( .A(n14954), .B(n14953), .Z(n14977) );
  AND U16022 ( .A(a[603]), .B(b[3]), .Z(n14976) );
  XOR U16023 ( .A(n14977), .B(n14976), .Z(n14979) );
  XOR U16024 ( .A(n14978), .B(n14979), .Z(n14967) );
  NANDN U16025 ( .A(n14956), .B(n14955), .Z(n14960) );
  OR U16026 ( .A(n14958), .B(n14957), .Z(n14959) );
  AND U16027 ( .A(n14960), .B(n14959), .Z(n14966) );
  XOR U16028 ( .A(n14967), .B(n14966), .Z(n14969) );
  XOR U16029 ( .A(n14968), .B(n14969), .Z(n14982) );
  XNOR U16030 ( .A(n14982), .B(sreg[1627]), .Z(n14984) );
  NANDN U16031 ( .A(n14961), .B(sreg[1626]), .Z(n14965) );
  NAND U16032 ( .A(n14963), .B(n14962), .Z(n14964) );
  NAND U16033 ( .A(n14965), .B(n14964), .Z(n14983) );
  XOR U16034 ( .A(n14984), .B(n14983), .Z(c[1627]) );
  NANDN U16035 ( .A(n14967), .B(n14966), .Z(n14971) );
  OR U16036 ( .A(n14969), .B(n14968), .Z(n14970) );
  AND U16037 ( .A(n14971), .B(n14970), .Z(n14989) );
  XOR U16038 ( .A(a[606]), .B(n2262), .Z(n14993) );
  AND U16039 ( .A(a[604]), .B(b[3]), .Z(n14997) );
  AND U16040 ( .A(a[608]), .B(b[0]), .Z(n14973) );
  XNOR U16041 ( .A(n14973), .B(n2175), .Z(n14975) );
  NANDN U16042 ( .A(b[0]), .B(a[607]), .Z(n14974) );
  NAND U16043 ( .A(n14975), .B(n14974), .Z(n14998) );
  XOR U16044 ( .A(n14997), .B(n14998), .Z(n15000) );
  XOR U16045 ( .A(n14999), .B(n15000), .Z(n14988) );
  NANDN U16046 ( .A(n14977), .B(n14976), .Z(n14981) );
  OR U16047 ( .A(n14979), .B(n14978), .Z(n14980) );
  AND U16048 ( .A(n14981), .B(n14980), .Z(n14987) );
  XOR U16049 ( .A(n14988), .B(n14987), .Z(n14990) );
  XOR U16050 ( .A(n14989), .B(n14990), .Z(n15003) );
  XNOR U16051 ( .A(n15003), .B(sreg[1628]), .Z(n15005) );
  NANDN U16052 ( .A(n14982), .B(sreg[1627]), .Z(n14986) );
  NAND U16053 ( .A(n14984), .B(n14983), .Z(n14985) );
  NAND U16054 ( .A(n14986), .B(n14985), .Z(n15004) );
  XOR U16055 ( .A(n15005), .B(n15004), .Z(c[1628]) );
  NANDN U16056 ( .A(n14988), .B(n14987), .Z(n14992) );
  OR U16057 ( .A(n14990), .B(n14989), .Z(n14991) );
  AND U16058 ( .A(n14992), .B(n14991), .Z(n15010) );
  XOR U16059 ( .A(a[607]), .B(n2262), .Z(n15014) );
  AND U16060 ( .A(a[609]), .B(b[0]), .Z(n14994) );
  XNOR U16061 ( .A(n14994), .B(n2175), .Z(n14996) );
  NANDN U16062 ( .A(b[0]), .B(a[608]), .Z(n14995) );
  NAND U16063 ( .A(n14996), .B(n14995), .Z(n15019) );
  AND U16064 ( .A(a[605]), .B(b[3]), .Z(n15018) );
  XOR U16065 ( .A(n15019), .B(n15018), .Z(n15021) );
  XOR U16066 ( .A(n15020), .B(n15021), .Z(n15009) );
  NANDN U16067 ( .A(n14998), .B(n14997), .Z(n15002) );
  OR U16068 ( .A(n15000), .B(n14999), .Z(n15001) );
  AND U16069 ( .A(n15002), .B(n15001), .Z(n15008) );
  XOR U16070 ( .A(n15009), .B(n15008), .Z(n15011) );
  XOR U16071 ( .A(n15010), .B(n15011), .Z(n15024) );
  XNOR U16072 ( .A(n15024), .B(sreg[1629]), .Z(n15026) );
  NANDN U16073 ( .A(n15003), .B(sreg[1628]), .Z(n15007) );
  NAND U16074 ( .A(n15005), .B(n15004), .Z(n15006) );
  NAND U16075 ( .A(n15007), .B(n15006), .Z(n15025) );
  XOR U16076 ( .A(n15026), .B(n15025), .Z(c[1629]) );
  NANDN U16077 ( .A(n15009), .B(n15008), .Z(n15013) );
  OR U16078 ( .A(n15011), .B(n15010), .Z(n15012) );
  AND U16079 ( .A(n15013), .B(n15012), .Z(n15031) );
  XOR U16080 ( .A(a[608]), .B(n2263), .Z(n15035) );
  AND U16081 ( .A(a[606]), .B(b[3]), .Z(n15039) );
  AND U16082 ( .A(a[610]), .B(b[0]), .Z(n15015) );
  XNOR U16083 ( .A(n15015), .B(n2175), .Z(n15017) );
  NANDN U16084 ( .A(b[0]), .B(a[609]), .Z(n15016) );
  NAND U16085 ( .A(n15017), .B(n15016), .Z(n15040) );
  XOR U16086 ( .A(n15039), .B(n15040), .Z(n15042) );
  XOR U16087 ( .A(n15041), .B(n15042), .Z(n15030) );
  NANDN U16088 ( .A(n15019), .B(n15018), .Z(n15023) );
  OR U16089 ( .A(n15021), .B(n15020), .Z(n15022) );
  AND U16090 ( .A(n15023), .B(n15022), .Z(n15029) );
  XOR U16091 ( .A(n15030), .B(n15029), .Z(n15032) );
  XOR U16092 ( .A(n15031), .B(n15032), .Z(n15045) );
  XNOR U16093 ( .A(n15045), .B(sreg[1630]), .Z(n15047) );
  NANDN U16094 ( .A(n15024), .B(sreg[1629]), .Z(n15028) );
  NAND U16095 ( .A(n15026), .B(n15025), .Z(n15027) );
  NAND U16096 ( .A(n15028), .B(n15027), .Z(n15046) );
  XOR U16097 ( .A(n15047), .B(n15046), .Z(c[1630]) );
  NANDN U16098 ( .A(n15030), .B(n15029), .Z(n15034) );
  OR U16099 ( .A(n15032), .B(n15031), .Z(n15033) );
  AND U16100 ( .A(n15034), .B(n15033), .Z(n15052) );
  XOR U16101 ( .A(a[609]), .B(n2263), .Z(n15056) );
  AND U16102 ( .A(a[611]), .B(b[0]), .Z(n15036) );
  XNOR U16103 ( .A(n15036), .B(n2175), .Z(n15038) );
  NANDN U16104 ( .A(b[0]), .B(a[610]), .Z(n15037) );
  NAND U16105 ( .A(n15038), .B(n15037), .Z(n15061) );
  AND U16106 ( .A(a[607]), .B(b[3]), .Z(n15060) );
  XOR U16107 ( .A(n15061), .B(n15060), .Z(n15063) );
  XOR U16108 ( .A(n15062), .B(n15063), .Z(n15051) );
  NANDN U16109 ( .A(n15040), .B(n15039), .Z(n15044) );
  OR U16110 ( .A(n15042), .B(n15041), .Z(n15043) );
  AND U16111 ( .A(n15044), .B(n15043), .Z(n15050) );
  XOR U16112 ( .A(n15051), .B(n15050), .Z(n15053) );
  XOR U16113 ( .A(n15052), .B(n15053), .Z(n15066) );
  XNOR U16114 ( .A(n15066), .B(sreg[1631]), .Z(n15068) );
  NANDN U16115 ( .A(n15045), .B(sreg[1630]), .Z(n15049) );
  NAND U16116 ( .A(n15047), .B(n15046), .Z(n15048) );
  NAND U16117 ( .A(n15049), .B(n15048), .Z(n15067) );
  XOR U16118 ( .A(n15068), .B(n15067), .Z(c[1631]) );
  NANDN U16119 ( .A(n15051), .B(n15050), .Z(n15055) );
  OR U16120 ( .A(n15053), .B(n15052), .Z(n15054) );
  AND U16121 ( .A(n15055), .B(n15054), .Z(n15073) );
  XOR U16122 ( .A(a[610]), .B(n2263), .Z(n15077) );
  AND U16123 ( .A(a[608]), .B(b[3]), .Z(n15081) );
  AND U16124 ( .A(a[612]), .B(b[0]), .Z(n15057) );
  XNOR U16125 ( .A(n15057), .B(n2175), .Z(n15059) );
  NANDN U16126 ( .A(b[0]), .B(a[611]), .Z(n15058) );
  NAND U16127 ( .A(n15059), .B(n15058), .Z(n15082) );
  XOR U16128 ( .A(n15081), .B(n15082), .Z(n15084) );
  XOR U16129 ( .A(n15083), .B(n15084), .Z(n15072) );
  NANDN U16130 ( .A(n15061), .B(n15060), .Z(n15065) );
  OR U16131 ( .A(n15063), .B(n15062), .Z(n15064) );
  AND U16132 ( .A(n15065), .B(n15064), .Z(n15071) );
  XOR U16133 ( .A(n15072), .B(n15071), .Z(n15074) );
  XOR U16134 ( .A(n15073), .B(n15074), .Z(n15087) );
  XNOR U16135 ( .A(n15087), .B(sreg[1632]), .Z(n15089) );
  NANDN U16136 ( .A(n15066), .B(sreg[1631]), .Z(n15070) );
  NAND U16137 ( .A(n15068), .B(n15067), .Z(n15069) );
  NAND U16138 ( .A(n15070), .B(n15069), .Z(n15088) );
  XOR U16139 ( .A(n15089), .B(n15088), .Z(c[1632]) );
  NANDN U16140 ( .A(n15072), .B(n15071), .Z(n15076) );
  OR U16141 ( .A(n15074), .B(n15073), .Z(n15075) );
  AND U16142 ( .A(n15076), .B(n15075), .Z(n15094) );
  XOR U16143 ( .A(a[611]), .B(n2263), .Z(n15098) );
  AND U16144 ( .A(a[613]), .B(b[0]), .Z(n15078) );
  XNOR U16145 ( .A(n15078), .B(n2175), .Z(n15080) );
  NANDN U16146 ( .A(b[0]), .B(a[612]), .Z(n15079) );
  NAND U16147 ( .A(n15080), .B(n15079), .Z(n15103) );
  AND U16148 ( .A(a[609]), .B(b[3]), .Z(n15102) );
  XOR U16149 ( .A(n15103), .B(n15102), .Z(n15105) );
  XOR U16150 ( .A(n15104), .B(n15105), .Z(n15093) );
  NANDN U16151 ( .A(n15082), .B(n15081), .Z(n15086) );
  OR U16152 ( .A(n15084), .B(n15083), .Z(n15085) );
  AND U16153 ( .A(n15086), .B(n15085), .Z(n15092) );
  XOR U16154 ( .A(n15093), .B(n15092), .Z(n15095) );
  XOR U16155 ( .A(n15094), .B(n15095), .Z(n15108) );
  XNOR U16156 ( .A(n15108), .B(sreg[1633]), .Z(n15110) );
  NANDN U16157 ( .A(n15087), .B(sreg[1632]), .Z(n15091) );
  NAND U16158 ( .A(n15089), .B(n15088), .Z(n15090) );
  NAND U16159 ( .A(n15091), .B(n15090), .Z(n15109) );
  XOR U16160 ( .A(n15110), .B(n15109), .Z(c[1633]) );
  NANDN U16161 ( .A(n15093), .B(n15092), .Z(n15097) );
  OR U16162 ( .A(n15095), .B(n15094), .Z(n15096) );
  AND U16163 ( .A(n15097), .B(n15096), .Z(n15115) );
  XOR U16164 ( .A(a[612]), .B(n2263), .Z(n15119) );
  AND U16165 ( .A(a[614]), .B(b[0]), .Z(n15099) );
  XNOR U16166 ( .A(n15099), .B(n2175), .Z(n15101) );
  NANDN U16167 ( .A(b[0]), .B(a[613]), .Z(n15100) );
  NAND U16168 ( .A(n15101), .B(n15100), .Z(n15124) );
  AND U16169 ( .A(a[610]), .B(b[3]), .Z(n15123) );
  XOR U16170 ( .A(n15124), .B(n15123), .Z(n15126) );
  XOR U16171 ( .A(n15125), .B(n15126), .Z(n15114) );
  NANDN U16172 ( .A(n15103), .B(n15102), .Z(n15107) );
  OR U16173 ( .A(n15105), .B(n15104), .Z(n15106) );
  AND U16174 ( .A(n15107), .B(n15106), .Z(n15113) );
  XOR U16175 ( .A(n15114), .B(n15113), .Z(n15116) );
  XOR U16176 ( .A(n15115), .B(n15116), .Z(n15129) );
  XNOR U16177 ( .A(n15129), .B(sreg[1634]), .Z(n15131) );
  NANDN U16178 ( .A(n15108), .B(sreg[1633]), .Z(n15112) );
  NAND U16179 ( .A(n15110), .B(n15109), .Z(n15111) );
  NAND U16180 ( .A(n15112), .B(n15111), .Z(n15130) );
  XOR U16181 ( .A(n15131), .B(n15130), .Z(c[1634]) );
  NANDN U16182 ( .A(n15114), .B(n15113), .Z(n15118) );
  OR U16183 ( .A(n15116), .B(n15115), .Z(n15117) );
  AND U16184 ( .A(n15118), .B(n15117), .Z(n15136) );
  XOR U16185 ( .A(a[613]), .B(n2263), .Z(n15140) );
  AND U16186 ( .A(a[611]), .B(b[3]), .Z(n15144) );
  AND U16187 ( .A(a[615]), .B(b[0]), .Z(n15120) );
  XNOR U16188 ( .A(n15120), .B(n2175), .Z(n15122) );
  NANDN U16189 ( .A(b[0]), .B(a[614]), .Z(n15121) );
  NAND U16190 ( .A(n15122), .B(n15121), .Z(n15145) );
  XOR U16191 ( .A(n15144), .B(n15145), .Z(n15147) );
  XOR U16192 ( .A(n15146), .B(n15147), .Z(n15135) );
  NANDN U16193 ( .A(n15124), .B(n15123), .Z(n15128) );
  OR U16194 ( .A(n15126), .B(n15125), .Z(n15127) );
  AND U16195 ( .A(n15128), .B(n15127), .Z(n15134) );
  XOR U16196 ( .A(n15135), .B(n15134), .Z(n15137) );
  XOR U16197 ( .A(n15136), .B(n15137), .Z(n15150) );
  XNOR U16198 ( .A(n15150), .B(sreg[1635]), .Z(n15152) );
  NANDN U16199 ( .A(n15129), .B(sreg[1634]), .Z(n15133) );
  NAND U16200 ( .A(n15131), .B(n15130), .Z(n15132) );
  NAND U16201 ( .A(n15133), .B(n15132), .Z(n15151) );
  XOR U16202 ( .A(n15152), .B(n15151), .Z(c[1635]) );
  NANDN U16203 ( .A(n15135), .B(n15134), .Z(n15139) );
  OR U16204 ( .A(n15137), .B(n15136), .Z(n15138) );
  AND U16205 ( .A(n15139), .B(n15138), .Z(n15157) );
  XOR U16206 ( .A(a[614]), .B(n2263), .Z(n15161) );
  AND U16207 ( .A(a[616]), .B(b[0]), .Z(n15141) );
  XNOR U16208 ( .A(n15141), .B(n2175), .Z(n15143) );
  NANDN U16209 ( .A(b[0]), .B(a[615]), .Z(n15142) );
  NAND U16210 ( .A(n15143), .B(n15142), .Z(n15166) );
  AND U16211 ( .A(a[612]), .B(b[3]), .Z(n15165) );
  XOR U16212 ( .A(n15166), .B(n15165), .Z(n15168) );
  XOR U16213 ( .A(n15167), .B(n15168), .Z(n15156) );
  NANDN U16214 ( .A(n15145), .B(n15144), .Z(n15149) );
  OR U16215 ( .A(n15147), .B(n15146), .Z(n15148) );
  AND U16216 ( .A(n15149), .B(n15148), .Z(n15155) );
  XOR U16217 ( .A(n15156), .B(n15155), .Z(n15158) );
  XOR U16218 ( .A(n15157), .B(n15158), .Z(n15171) );
  XNOR U16219 ( .A(n15171), .B(sreg[1636]), .Z(n15173) );
  NANDN U16220 ( .A(n15150), .B(sreg[1635]), .Z(n15154) );
  NAND U16221 ( .A(n15152), .B(n15151), .Z(n15153) );
  NAND U16222 ( .A(n15154), .B(n15153), .Z(n15172) );
  XOR U16223 ( .A(n15173), .B(n15172), .Z(c[1636]) );
  NANDN U16224 ( .A(n15156), .B(n15155), .Z(n15160) );
  OR U16225 ( .A(n15158), .B(n15157), .Z(n15159) );
  AND U16226 ( .A(n15160), .B(n15159), .Z(n15178) );
  XOR U16227 ( .A(a[615]), .B(n2264), .Z(n15182) );
  AND U16228 ( .A(a[617]), .B(b[0]), .Z(n15162) );
  XNOR U16229 ( .A(n15162), .B(n2175), .Z(n15164) );
  NANDN U16230 ( .A(b[0]), .B(a[616]), .Z(n15163) );
  NAND U16231 ( .A(n15164), .B(n15163), .Z(n15187) );
  AND U16232 ( .A(a[613]), .B(b[3]), .Z(n15186) );
  XOR U16233 ( .A(n15187), .B(n15186), .Z(n15189) );
  XOR U16234 ( .A(n15188), .B(n15189), .Z(n15177) );
  NANDN U16235 ( .A(n15166), .B(n15165), .Z(n15170) );
  OR U16236 ( .A(n15168), .B(n15167), .Z(n15169) );
  AND U16237 ( .A(n15170), .B(n15169), .Z(n15176) );
  XOR U16238 ( .A(n15177), .B(n15176), .Z(n15179) );
  XOR U16239 ( .A(n15178), .B(n15179), .Z(n15192) );
  XNOR U16240 ( .A(n15192), .B(sreg[1637]), .Z(n15194) );
  NANDN U16241 ( .A(n15171), .B(sreg[1636]), .Z(n15175) );
  NAND U16242 ( .A(n15173), .B(n15172), .Z(n15174) );
  NAND U16243 ( .A(n15175), .B(n15174), .Z(n15193) );
  XOR U16244 ( .A(n15194), .B(n15193), .Z(c[1637]) );
  NANDN U16245 ( .A(n15177), .B(n15176), .Z(n15181) );
  OR U16246 ( .A(n15179), .B(n15178), .Z(n15180) );
  AND U16247 ( .A(n15181), .B(n15180), .Z(n15199) );
  XOR U16248 ( .A(a[616]), .B(n2264), .Z(n15203) );
  AND U16249 ( .A(a[618]), .B(b[0]), .Z(n15183) );
  XNOR U16250 ( .A(n15183), .B(n2175), .Z(n15185) );
  NANDN U16251 ( .A(b[0]), .B(a[617]), .Z(n15184) );
  NAND U16252 ( .A(n15185), .B(n15184), .Z(n15208) );
  AND U16253 ( .A(a[614]), .B(b[3]), .Z(n15207) );
  XOR U16254 ( .A(n15208), .B(n15207), .Z(n15210) );
  XOR U16255 ( .A(n15209), .B(n15210), .Z(n15198) );
  NANDN U16256 ( .A(n15187), .B(n15186), .Z(n15191) );
  OR U16257 ( .A(n15189), .B(n15188), .Z(n15190) );
  AND U16258 ( .A(n15191), .B(n15190), .Z(n15197) );
  XOR U16259 ( .A(n15198), .B(n15197), .Z(n15200) );
  XOR U16260 ( .A(n15199), .B(n15200), .Z(n15213) );
  XNOR U16261 ( .A(n15213), .B(sreg[1638]), .Z(n15215) );
  NANDN U16262 ( .A(n15192), .B(sreg[1637]), .Z(n15196) );
  NAND U16263 ( .A(n15194), .B(n15193), .Z(n15195) );
  NAND U16264 ( .A(n15196), .B(n15195), .Z(n15214) );
  XOR U16265 ( .A(n15215), .B(n15214), .Z(c[1638]) );
  NANDN U16266 ( .A(n15198), .B(n15197), .Z(n15202) );
  OR U16267 ( .A(n15200), .B(n15199), .Z(n15201) );
  AND U16268 ( .A(n15202), .B(n15201), .Z(n15220) );
  XOR U16269 ( .A(a[617]), .B(n2264), .Z(n15224) );
  AND U16270 ( .A(a[615]), .B(b[3]), .Z(n15228) );
  AND U16271 ( .A(a[619]), .B(b[0]), .Z(n15204) );
  XNOR U16272 ( .A(n15204), .B(n2175), .Z(n15206) );
  NANDN U16273 ( .A(b[0]), .B(a[618]), .Z(n15205) );
  NAND U16274 ( .A(n15206), .B(n15205), .Z(n15229) );
  XOR U16275 ( .A(n15228), .B(n15229), .Z(n15231) );
  XOR U16276 ( .A(n15230), .B(n15231), .Z(n15219) );
  NANDN U16277 ( .A(n15208), .B(n15207), .Z(n15212) );
  OR U16278 ( .A(n15210), .B(n15209), .Z(n15211) );
  AND U16279 ( .A(n15212), .B(n15211), .Z(n15218) );
  XOR U16280 ( .A(n15219), .B(n15218), .Z(n15221) );
  XOR U16281 ( .A(n15220), .B(n15221), .Z(n15234) );
  XNOR U16282 ( .A(n15234), .B(sreg[1639]), .Z(n15236) );
  NANDN U16283 ( .A(n15213), .B(sreg[1638]), .Z(n15217) );
  NAND U16284 ( .A(n15215), .B(n15214), .Z(n15216) );
  NAND U16285 ( .A(n15217), .B(n15216), .Z(n15235) );
  XOR U16286 ( .A(n15236), .B(n15235), .Z(c[1639]) );
  NANDN U16287 ( .A(n15219), .B(n15218), .Z(n15223) );
  OR U16288 ( .A(n15221), .B(n15220), .Z(n15222) );
  AND U16289 ( .A(n15223), .B(n15222), .Z(n15241) );
  XOR U16290 ( .A(a[618]), .B(n2264), .Z(n15245) );
  AND U16291 ( .A(a[620]), .B(b[0]), .Z(n15225) );
  XNOR U16292 ( .A(n15225), .B(n2175), .Z(n15227) );
  NANDN U16293 ( .A(b[0]), .B(a[619]), .Z(n15226) );
  NAND U16294 ( .A(n15227), .B(n15226), .Z(n15250) );
  AND U16295 ( .A(a[616]), .B(b[3]), .Z(n15249) );
  XOR U16296 ( .A(n15250), .B(n15249), .Z(n15252) );
  XOR U16297 ( .A(n15251), .B(n15252), .Z(n15240) );
  NANDN U16298 ( .A(n15229), .B(n15228), .Z(n15233) );
  OR U16299 ( .A(n15231), .B(n15230), .Z(n15232) );
  AND U16300 ( .A(n15233), .B(n15232), .Z(n15239) );
  XOR U16301 ( .A(n15240), .B(n15239), .Z(n15242) );
  XOR U16302 ( .A(n15241), .B(n15242), .Z(n15255) );
  XNOR U16303 ( .A(n15255), .B(sreg[1640]), .Z(n15257) );
  NANDN U16304 ( .A(n15234), .B(sreg[1639]), .Z(n15238) );
  NAND U16305 ( .A(n15236), .B(n15235), .Z(n15237) );
  NAND U16306 ( .A(n15238), .B(n15237), .Z(n15256) );
  XOR U16307 ( .A(n15257), .B(n15256), .Z(c[1640]) );
  NANDN U16308 ( .A(n15240), .B(n15239), .Z(n15244) );
  OR U16309 ( .A(n15242), .B(n15241), .Z(n15243) );
  AND U16310 ( .A(n15244), .B(n15243), .Z(n15262) );
  XOR U16311 ( .A(a[619]), .B(n2264), .Z(n15266) );
  AND U16312 ( .A(a[617]), .B(b[3]), .Z(n15270) );
  AND U16313 ( .A(a[621]), .B(b[0]), .Z(n15246) );
  XNOR U16314 ( .A(n15246), .B(n2175), .Z(n15248) );
  NANDN U16315 ( .A(b[0]), .B(a[620]), .Z(n15247) );
  NAND U16316 ( .A(n15248), .B(n15247), .Z(n15271) );
  XOR U16317 ( .A(n15270), .B(n15271), .Z(n15273) );
  XOR U16318 ( .A(n15272), .B(n15273), .Z(n15261) );
  NANDN U16319 ( .A(n15250), .B(n15249), .Z(n15254) );
  OR U16320 ( .A(n15252), .B(n15251), .Z(n15253) );
  AND U16321 ( .A(n15254), .B(n15253), .Z(n15260) );
  XOR U16322 ( .A(n15261), .B(n15260), .Z(n15263) );
  XOR U16323 ( .A(n15262), .B(n15263), .Z(n15276) );
  XNOR U16324 ( .A(n15276), .B(sreg[1641]), .Z(n15278) );
  NANDN U16325 ( .A(n15255), .B(sreg[1640]), .Z(n15259) );
  NAND U16326 ( .A(n15257), .B(n15256), .Z(n15258) );
  NAND U16327 ( .A(n15259), .B(n15258), .Z(n15277) );
  XOR U16328 ( .A(n15278), .B(n15277), .Z(c[1641]) );
  NANDN U16329 ( .A(n15261), .B(n15260), .Z(n15265) );
  OR U16330 ( .A(n15263), .B(n15262), .Z(n15264) );
  AND U16331 ( .A(n15265), .B(n15264), .Z(n15283) );
  XOR U16332 ( .A(a[620]), .B(n2264), .Z(n15287) );
  AND U16333 ( .A(a[622]), .B(b[0]), .Z(n15267) );
  XNOR U16334 ( .A(n15267), .B(n2175), .Z(n15269) );
  NANDN U16335 ( .A(b[0]), .B(a[621]), .Z(n15268) );
  NAND U16336 ( .A(n15269), .B(n15268), .Z(n15292) );
  AND U16337 ( .A(a[618]), .B(b[3]), .Z(n15291) );
  XOR U16338 ( .A(n15292), .B(n15291), .Z(n15294) );
  XOR U16339 ( .A(n15293), .B(n15294), .Z(n15282) );
  NANDN U16340 ( .A(n15271), .B(n15270), .Z(n15275) );
  OR U16341 ( .A(n15273), .B(n15272), .Z(n15274) );
  AND U16342 ( .A(n15275), .B(n15274), .Z(n15281) );
  XOR U16343 ( .A(n15282), .B(n15281), .Z(n15284) );
  XOR U16344 ( .A(n15283), .B(n15284), .Z(n15297) );
  XNOR U16345 ( .A(n15297), .B(sreg[1642]), .Z(n15299) );
  NANDN U16346 ( .A(n15276), .B(sreg[1641]), .Z(n15280) );
  NAND U16347 ( .A(n15278), .B(n15277), .Z(n15279) );
  NAND U16348 ( .A(n15280), .B(n15279), .Z(n15298) );
  XOR U16349 ( .A(n15299), .B(n15298), .Z(c[1642]) );
  NANDN U16350 ( .A(n15282), .B(n15281), .Z(n15286) );
  OR U16351 ( .A(n15284), .B(n15283), .Z(n15285) );
  AND U16352 ( .A(n15286), .B(n15285), .Z(n15304) );
  XOR U16353 ( .A(a[621]), .B(n2264), .Z(n15308) );
  AND U16354 ( .A(a[619]), .B(b[3]), .Z(n15312) );
  AND U16355 ( .A(a[623]), .B(b[0]), .Z(n15288) );
  XNOR U16356 ( .A(n15288), .B(n2175), .Z(n15290) );
  NANDN U16357 ( .A(b[0]), .B(a[622]), .Z(n15289) );
  NAND U16358 ( .A(n15290), .B(n15289), .Z(n15313) );
  XOR U16359 ( .A(n15312), .B(n15313), .Z(n15315) );
  XOR U16360 ( .A(n15314), .B(n15315), .Z(n15303) );
  NANDN U16361 ( .A(n15292), .B(n15291), .Z(n15296) );
  OR U16362 ( .A(n15294), .B(n15293), .Z(n15295) );
  AND U16363 ( .A(n15296), .B(n15295), .Z(n15302) );
  XOR U16364 ( .A(n15303), .B(n15302), .Z(n15305) );
  XOR U16365 ( .A(n15304), .B(n15305), .Z(n15318) );
  XNOR U16366 ( .A(n15318), .B(sreg[1643]), .Z(n15320) );
  NANDN U16367 ( .A(n15297), .B(sreg[1642]), .Z(n15301) );
  NAND U16368 ( .A(n15299), .B(n15298), .Z(n15300) );
  NAND U16369 ( .A(n15301), .B(n15300), .Z(n15319) );
  XOR U16370 ( .A(n15320), .B(n15319), .Z(c[1643]) );
  NANDN U16371 ( .A(n15303), .B(n15302), .Z(n15307) );
  OR U16372 ( .A(n15305), .B(n15304), .Z(n15306) );
  AND U16373 ( .A(n15307), .B(n15306), .Z(n15325) );
  XOR U16374 ( .A(a[622]), .B(n2265), .Z(n15329) );
  AND U16375 ( .A(a[624]), .B(b[0]), .Z(n15309) );
  XNOR U16376 ( .A(n15309), .B(n2175), .Z(n15311) );
  NANDN U16377 ( .A(b[0]), .B(a[623]), .Z(n15310) );
  NAND U16378 ( .A(n15311), .B(n15310), .Z(n15334) );
  AND U16379 ( .A(a[620]), .B(b[3]), .Z(n15333) );
  XOR U16380 ( .A(n15334), .B(n15333), .Z(n15336) );
  XOR U16381 ( .A(n15335), .B(n15336), .Z(n15324) );
  NANDN U16382 ( .A(n15313), .B(n15312), .Z(n15317) );
  OR U16383 ( .A(n15315), .B(n15314), .Z(n15316) );
  AND U16384 ( .A(n15317), .B(n15316), .Z(n15323) );
  XOR U16385 ( .A(n15324), .B(n15323), .Z(n15326) );
  XOR U16386 ( .A(n15325), .B(n15326), .Z(n15339) );
  XNOR U16387 ( .A(n15339), .B(sreg[1644]), .Z(n15341) );
  NANDN U16388 ( .A(n15318), .B(sreg[1643]), .Z(n15322) );
  NAND U16389 ( .A(n15320), .B(n15319), .Z(n15321) );
  NAND U16390 ( .A(n15322), .B(n15321), .Z(n15340) );
  XOR U16391 ( .A(n15341), .B(n15340), .Z(c[1644]) );
  NANDN U16392 ( .A(n15324), .B(n15323), .Z(n15328) );
  OR U16393 ( .A(n15326), .B(n15325), .Z(n15327) );
  AND U16394 ( .A(n15328), .B(n15327), .Z(n15346) );
  XOR U16395 ( .A(a[623]), .B(n2265), .Z(n15350) );
  AND U16396 ( .A(a[621]), .B(b[3]), .Z(n15354) );
  AND U16397 ( .A(a[625]), .B(b[0]), .Z(n15330) );
  XNOR U16398 ( .A(n15330), .B(n2175), .Z(n15332) );
  NANDN U16399 ( .A(b[0]), .B(a[624]), .Z(n15331) );
  NAND U16400 ( .A(n15332), .B(n15331), .Z(n15355) );
  XOR U16401 ( .A(n15354), .B(n15355), .Z(n15357) );
  XOR U16402 ( .A(n15356), .B(n15357), .Z(n15345) );
  NANDN U16403 ( .A(n15334), .B(n15333), .Z(n15338) );
  OR U16404 ( .A(n15336), .B(n15335), .Z(n15337) );
  AND U16405 ( .A(n15338), .B(n15337), .Z(n15344) );
  XOR U16406 ( .A(n15345), .B(n15344), .Z(n15347) );
  XOR U16407 ( .A(n15346), .B(n15347), .Z(n15360) );
  XNOR U16408 ( .A(n15360), .B(sreg[1645]), .Z(n15362) );
  NANDN U16409 ( .A(n15339), .B(sreg[1644]), .Z(n15343) );
  NAND U16410 ( .A(n15341), .B(n15340), .Z(n15342) );
  NAND U16411 ( .A(n15343), .B(n15342), .Z(n15361) );
  XOR U16412 ( .A(n15362), .B(n15361), .Z(c[1645]) );
  NANDN U16413 ( .A(n15345), .B(n15344), .Z(n15349) );
  OR U16414 ( .A(n15347), .B(n15346), .Z(n15348) );
  AND U16415 ( .A(n15349), .B(n15348), .Z(n15367) );
  XOR U16416 ( .A(a[624]), .B(n2265), .Z(n15371) );
  AND U16417 ( .A(a[626]), .B(b[0]), .Z(n15351) );
  XNOR U16418 ( .A(n15351), .B(n2175), .Z(n15353) );
  NANDN U16419 ( .A(b[0]), .B(a[625]), .Z(n15352) );
  NAND U16420 ( .A(n15353), .B(n15352), .Z(n15376) );
  AND U16421 ( .A(a[622]), .B(b[3]), .Z(n15375) );
  XOR U16422 ( .A(n15376), .B(n15375), .Z(n15378) );
  XOR U16423 ( .A(n15377), .B(n15378), .Z(n15366) );
  NANDN U16424 ( .A(n15355), .B(n15354), .Z(n15359) );
  OR U16425 ( .A(n15357), .B(n15356), .Z(n15358) );
  AND U16426 ( .A(n15359), .B(n15358), .Z(n15365) );
  XOR U16427 ( .A(n15366), .B(n15365), .Z(n15368) );
  XOR U16428 ( .A(n15367), .B(n15368), .Z(n15381) );
  XNOR U16429 ( .A(n15381), .B(sreg[1646]), .Z(n15383) );
  NANDN U16430 ( .A(n15360), .B(sreg[1645]), .Z(n15364) );
  NAND U16431 ( .A(n15362), .B(n15361), .Z(n15363) );
  NAND U16432 ( .A(n15364), .B(n15363), .Z(n15382) );
  XOR U16433 ( .A(n15383), .B(n15382), .Z(c[1646]) );
  NANDN U16434 ( .A(n15366), .B(n15365), .Z(n15370) );
  OR U16435 ( .A(n15368), .B(n15367), .Z(n15369) );
  AND U16436 ( .A(n15370), .B(n15369), .Z(n15388) );
  XOR U16437 ( .A(a[625]), .B(n2265), .Z(n15392) );
  AND U16438 ( .A(a[623]), .B(b[3]), .Z(n15396) );
  AND U16439 ( .A(a[627]), .B(b[0]), .Z(n15372) );
  XNOR U16440 ( .A(n15372), .B(n2175), .Z(n15374) );
  NANDN U16441 ( .A(b[0]), .B(a[626]), .Z(n15373) );
  NAND U16442 ( .A(n15374), .B(n15373), .Z(n15397) );
  XOR U16443 ( .A(n15396), .B(n15397), .Z(n15399) );
  XOR U16444 ( .A(n15398), .B(n15399), .Z(n15387) );
  NANDN U16445 ( .A(n15376), .B(n15375), .Z(n15380) );
  OR U16446 ( .A(n15378), .B(n15377), .Z(n15379) );
  AND U16447 ( .A(n15380), .B(n15379), .Z(n15386) );
  XOR U16448 ( .A(n15387), .B(n15386), .Z(n15389) );
  XOR U16449 ( .A(n15388), .B(n15389), .Z(n15402) );
  XNOR U16450 ( .A(n15402), .B(sreg[1647]), .Z(n15404) );
  NANDN U16451 ( .A(n15381), .B(sreg[1646]), .Z(n15385) );
  NAND U16452 ( .A(n15383), .B(n15382), .Z(n15384) );
  NAND U16453 ( .A(n15385), .B(n15384), .Z(n15403) );
  XOR U16454 ( .A(n15404), .B(n15403), .Z(c[1647]) );
  NANDN U16455 ( .A(n15387), .B(n15386), .Z(n15391) );
  OR U16456 ( .A(n15389), .B(n15388), .Z(n15390) );
  AND U16457 ( .A(n15391), .B(n15390), .Z(n15409) );
  XOR U16458 ( .A(a[626]), .B(n2265), .Z(n15413) );
  AND U16459 ( .A(a[628]), .B(b[0]), .Z(n15393) );
  XNOR U16460 ( .A(n15393), .B(n2175), .Z(n15395) );
  NANDN U16461 ( .A(b[0]), .B(a[627]), .Z(n15394) );
  NAND U16462 ( .A(n15395), .B(n15394), .Z(n15418) );
  AND U16463 ( .A(a[624]), .B(b[3]), .Z(n15417) );
  XOR U16464 ( .A(n15418), .B(n15417), .Z(n15420) );
  XOR U16465 ( .A(n15419), .B(n15420), .Z(n15408) );
  NANDN U16466 ( .A(n15397), .B(n15396), .Z(n15401) );
  OR U16467 ( .A(n15399), .B(n15398), .Z(n15400) );
  AND U16468 ( .A(n15401), .B(n15400), .Z(n15407) );
  XOR U16469 ( .A(n15408), .B(n15407), .Z(n15410) );
  XOR U16470 ( .A(n15409), .B(n15410), .Z(n15423) );
  XNOR U16471 ( .A(n15423), .B(sreg[1648]), .Z(n15425) );
  NANDN U16472 ( .A(n15402), .B(sreg[1647]), .Z(n15406) );
  NAND U16473 ( .A(n15404), .B(n15403), .Z(n15405) );
  NAND U16474 ( .A(n15406), .B(n15405), .Z(n15424) );
  XOR U16475 ( .A(n15425), .B(n15424), .Z(c[1648]) );
  NANDN U16476 ( .A(n15408), .B(n15407), .Z(n15412) );
  OR U16477 ( .A(n15410), .B(n15409), .Z(n15411) );
  AND U16478 ( .A(n15412), .B(n15411), .Z(n15430) );
  XOR U16479 ( .A(a[627]), .B(n2265), .Z(n15434) );
  AND U16480 ( .A(a[625]), .B(b[3]), .Z(n15438) );
  AND U16481 ( .A(a[629]), .B(b[0]), .Z(n15414) );
  XNOR U16482 ( .A(n15414), .B(n2175), .Z(n15416) );
  NANDN U16483 ( .A(b[0]), .B(a[628]), .Z(n15415) );
  NAND U16484 ( .A(n15416), .B(n15415), .Z(n15439) );
  XOR U16485 ( .A(n15438), .B(n15439), .Z(n15441) );
  XOR U16486 ( .A(n15440), .B(n15441), .Z(n15429) );
  NANDN U16487 ( .A(n15418), .B(n15417), .Z(n15422) );
  OR U16488 ( .A(n15420), .B(n15419), .Z(n15421) );
  AND U16489 ( .A(n15422), .B(n15421), .Z(n15428) );
  XOR U16490 ( .A(n15429), .B(n15428), .Z(n15431) );
  XOR U16491 ( .A(n15430), .B(n15431), .Z(n15444) );
  XNOR U16492 ( .A(n15444), .B(sreg[1649]), .Z(n15446) );
  NANDN U16493 ( .A(n15423), .B(sreg[1648]), .Z(n15427) );
  NAND U16494 ( .A(n15425), .B(n15424), .Z(n15426) );
  NAND U16495 ( .A(n15427), .B(n15426), .Z(n15445) );
  XOR U16496 ( .A(n15446), .B(n15445), .Z(c[1649]) );
  NANDN U16497 ( .A(n15429), .B(n15428), .Z(n15433) );
  OR U16498 ( .A(n15431), .B(n15430), .Z(n15432) );
  AND U16499 ( .A(n15433), .B(n15432), .Z(n15451) );
  XOR U16500 ( .A(a[628]), .B(n2265), .Z(n15455) );
  AND U16501 ( .A(a[626]), .B(b[3]), .Z(n15459) );
  AND U16502 ( .A(a[630]), .B(b[0]), .Z(n15435) );
  XNOR U16503 ( .A(n15435), .B(n2175), .Z(n15437) );
  NANDN U16504 ( .A(b[0]), .B(a[629]), .Z(n15436) );
  NAND U16505 ( .A(n15437), .B(n15436), .Z(n15460) );
  XOR U16506 ( .A(n15459), .B(n15460), .Z(n15462) );
  XOR U16507 ( .A(n15461), .B(n15462), .Z(n15450) );
  NANDN U16508 ( .A(n15439), .B(n15438), .Z(n15443) );
  OR U16509 ( .A(n15441), .B(n15440), .Z(n15442) );
  AND U16510 ( .A(n15443), .B(n15442), .Z(n15449) );
  XOR U16511 ( .A(n15450), .B(n15449), .Z(n15452) );
  XOR U16512 ( .A(n15451), .B(n15452), .Z(n15465) );
  XNOR U16513 ( .A(n15465), .B(sreg[1650]), .Z(n15467) );
  NANDN U16514 ( .A(n15444), .B(sreg[1649]), .Z(n15448) );
  NAND U16515 ( .A(n15446), .B(n15445), .Z(n15447) );
  NAND U16516 ( .A(n15448), .B(n15447), .Z(n15466) );
  XOR U16517 ( .A(n15467), .B(n15466), .Z(c[1650]) );
  NANDN U16518 ( .A(n15450), .B(n15449), .Z(n15454) );
  OR U16519 ( .A(n15452), .B(n15451), .Z(n15453) );
  AND U16520 ( .A(n15454), .B(n15453), .Z(n15472) );
  XOR U16521 ( .A(a[629]), .B(n2266), .Z(n15476) );
  AND U16522 ( .A(a[631]), .B(b[0]), .Z(n15456) );
  XNOR U16523 ( .A(n15456), .B(n2175), .Z(n15458) );
  NANDN U16524 ( .A(b[0]), .B(a[630]), .Z(n15457) );
  NAND U16525 ( .A(n15458), .B(n15457), .Z(n15481) );
  AND U16526 ( .A(a[627]), .B(b[3]), .Z(n15480) );
  XOR U16527 ( .A(n15481), .B(n15480), .Z(n15483) );
  XOR U16528 ( .A(n15482), .B(n15483), .Z(n15471) );
  NANDN U16529 ( .A(n15460), .B(n15459), .Z(n15464) );
  OR U16530 ( .A(n15462), .B(n15461), .Z(n15463) );
  AND U16531 ( .A(n15464), .B(n15463), .Z(n15470) );
  XOR U16532 ( .A(n15471), .B(n15470), .Z(n15473) );
  XOR U16533 ( .A(n15472), .B(n15473), .Z(n15486) );
  XNOR U16534 ( .A(n15486), .B(sreg[1651]), .Z(n15488) );
  NANDN U16535 ( .A(n15465), .B(sreg[1650]), .Z(n15469) );
  NAND U16536 ( .A(n15467), .B(n15466), .Z(n15468) );
  NAND U16537 ( .A(n15469), .B(n15468), .Z(n15487) );
  XOR U16538 ( .A(n15488), .B(n15487), .Z(c[1651]) );
  NANDN U16539 ( .A(n15471), .B(n15470), .Z(n15475) );
  OR U16540 ( .A(n15473), .B(n15472), .Z(n15474) );
  AND U16541 ( .A(n15475), .B(n15474), .Z(n15493) );
  XOR U16542 ( .A(a[630]), .B(n2266), .Z(n15497) );
  AND U16543 ( .A(a[632]), .B(b[0]), .Z(n15477) );
  XNOR U16544 ( .A(n15477), .B(n2175), .Z(n15479) );
  NANDN U16545 ( .A(b[0]), .B(a[631]), .Z(n15478) );
  NAND U16546 ( .A(n15479), .B(n15478), .Z(n15502) );
  AND U16547 ( .A(a[628]), .B(b[3]), .Z(n15501) );
  XOR U16548 ( .A(n15502), .B(n15501), .Z(n15504) );
  XOR U16549 ( .A(n15503), .B(n15504), .Z(n15492) );
  NANDN U16550 ( .A(n15481), .B(n15480), .Z(n15485) );
  OR U16551 ( .A(n15483), .B(n15482), .Z(n15484) );
  AND U16552 ( .A(n15485), .B(n15484), .Z(n15491) );
  XOR U16553 ( .A(n15492), .B(n15491), .Z(n15494) );
  XOR U16554 ( .A(n15493), .B(n15494), .Z(n15507) );
  XNOR U16555 ( .A(n15507), .B(sreg[1652]), .Z(n15509) );
  NANDN U16556 ( .A(n15486), .B(sreg[1651]), .Z(n15490) );
  NAND U16557 ( .A(n15488), .B(n15487), .Z(n15489) );
  NAND U16558 ( .A(n15490), .B(n15489), .Z(n15508) );
  XOR U16559 ( .A(n15509), .B(n15508), .Z(c[1652]) );
  NANDN U16560 ( .A(n15492), .B(n15491), .Z(n15496) );
  OR U16561 ( .A(n15494), .B(n15493), .Z(n15495) );
  AND U16562 ( .A(n15496), .B(n15495), .Z(n15514) );
  XOR U16563 ( .A(a[631]), .B(n2266), .Z(n15518) );
  AND U16564 ( .A(a[633]), .B(b[0]), .Z(n15498) );
  XNOR U16565 ( .A(n15498), .B(n2175), .Z(n15500) );
  NANDN U16566 ( .A(b[0]), .B(a[632]), .Z(n15499) );
  NAND U16567 ( .A(n15500), .B(n15499), .Z(n15523) );
  AND U16568 ( .A(a[629]), .B(b[3]), .Z(n15522) );
  XOR U16569 ( .A(n15523), .B(n15522), .Z(n15525) );
  XOR U16570 ( .A(n15524), .B(n15525), .Z(n15513) );
  NANDN U16571 ( .A(n15502), .B(n15501), .Z(n15506) );
  OR U16572 ( .A(n15504), .B(n15503), .Z(n15505) );
  AND U16573 ( .A(n15506), .B(n15505), .Z(n15512) );
  XOR U16574 ( .A(n15513), .B(n15512), .Z(n15515) );
  XOR U16575 ( .A(n15514), .B(n15515), .Z(n15528) );
  XNOR U16576 ( .A(n15528), .B(sreg[1653]), .Z(n15530) );
  NANDN U16577 ( .A(n15507), .B(sreg[1652]), .Z(n15511) );
  NAND U16578 ( .A(n15509), .B(n15508), .Z(n15510) );
  NAND U16579 ( .A(n15511), .B(n15510), .Z(n15529) );
  XOR U16580 ( .A(n15530), .B(n15529), .Z(c[1653]) );
  NANDN U16581 ( .A(n15513), .B(n15512), .Z(n15517) );
  OR U16582 ( .A(n15515), .B(n15514), .Z(n15516) );
  AND U16583 ( .A(n15517), .B(n15516), .Z(n15535) );
  XOR U16584 ( .A(a[632]), .B(n2266), .Z(n15539) );
  AND U16585 ( .A(a[634]), .B(b[0]), .Z(n15519) );
  XNOR U16586 ( .A(n15519), .B(n2175), .Z(n15521) );
  NANDN U16587 ( .A(b[0]), .B(a[633]), .Z(n15520) );
  NAND U16588 ( .A(n15521), .B(n15520), .Z(n15544) );
  AND U16589 ( .A(a[630]), .B(b[3]), .Z(n15543) );
  XOR U16590 ( .A(n15544), .B(n15543), .Z(n15546) );
  XOR U16591 ( .A(n15545), .B(n15546), .Z(n15534) );
  NANDN U16592 ( .A(n15523), .B(n15522), .Z(n15527) );
  OR U16593 ( .A(n15525), .B(n15524), .Z(n15526) );
  AND U16594 ( .A(n15527), .B(n15526), .Z(n15533) );
  XOR U16595 ( .A(n15534), .B(n15533), .Z(n15536) );
  XOR U16596 ( .A(n15535), .B(n15536), .Z(n15549) );
  XNOR U16597 ( .A(n15549), .B(sreg[1654]), .Z(n15551) );
  NANDN U16598 ( .A(n15528), .B(sreg[1653]), .Z(n15532) );
  NAND U16599 ( .A(n15530), .B(n15529), .Z(n15531) );
  NAND U16600 ( .A(n15532), .B(n15531), .Z(n15550) );
  XOR U16601 ( .A(n15551), .B(n15550), .Z(c[1654]) );
  NANDN U16602 ( .A(n15534), .B(n15533), .Z(n15538) );
  OR U16603 ( .A(n15536), .B(n15535), .Z(n15537) );
  AND U16604 ( .A(n15538), .B(n15537), .Z(n15556) );
  XOR U16605 ( .A(a[633]), .B(n2266), .Z(n15560) );
  AND U16606 ( .A(a[631]), .B(b[3]), .Z(n15564) );
  AND U16607 ( .A(a[635]), .B(b[0]), .Z(n15540) );
  XNOR U16608 ( .A(n15540), .B(n2175), .Z(n15542) );
  NANDN U16609 ( .A(b[0]), .B(a[634]), .Z(n15541) );
  NAND U16610 ( .A(n15542), .B(n15541), .Z(n15565) );
  XOR U16611 ( .A(n15564), .B(n15565), .Z(n15567) );
  XOR U16612 ( .A(n15566), .B(n15567), .Z(n15555) );
  NANDN U16613 ( .A(n15544), .B(n15543), .Z(n15548) );
  OR U16614 ( .A(n15546), .B(n15545), .Z(n15547) );
  AND U16615 ( .A(n15548), .B(n15547), .Z(n15554) );
  XOR U16616 ( .A(n15555), .B(n15554), .Z(n15557) );
  XOR U16617 ( .A(n15556), .B(n15557), .Z(n15570) );
  XNOR U16618 ( .A(n15570), .B(sreg[1655]), .Z(n15572) );
  NANDN U16619 ( .A(n15549), .B(sreg[1654]), .Z(n15553) );
  NAND U16620 ( .A(n15551), .B(n15550), .Z(n15552) );
  NAND U16621 ( .A(n15553), .B(n15552), .Z(n15571) );
  XOR U16622 ( .A(n15572), .B(n15571), .Z(c[1655]) );
  NANDN U16623 ( .A(n15555), .B(n15554), .Z(n15559) );
  OR U16624 ( .A(n15557), .B(n15556), .Z(n15558) );
  AND U16625 ( .A(n15559), .B(n15558), .Z(n15577) );
  XOR U16626 ( .A(a[634]), .B(n2266), .Z(n15581) );
  AND U16627 ( .A(a[636]), .B(b[0]), .Z(n15561) );
  XNOR U16628 ( .A(n15561), .B(n2175), .Z(n15563) );
  NANDN U16629 ( .A(b[0]), .B(a[635]), .Z(n15562) );
  NAND U16630 ( .A(n15563), .B(n15562), .Z(n15586) );
  AND U16631 ( .A(a[632]), .B(b[3]), .Z(n15585) );
  XOR U16632 ( .A(n15586), .B(n15585), .Z(n15588) );
  XOR U16633 ( .A(n15587), .B(n15588), .Z(n15576) );
  NANDN U16634 ( .A(n15565), .B(n15564), .Z(n15569) );
  OR U16635 ( .A(n15567), .B(n15566), .Z(n15568) );
  AND U16636 ( .A(n15569), .B(n15568), .Z(n15575) );
  XOR U16637 ( .A(n15576), .B(n15575), .Z(n15578) );
  XOR U16638 ( .A(n15577), .B(n15578), .Z(n15591) );
  XNOR U16639 ( .A(n15591), .B(sreg[1656]), .Z(n15593) );
  NANDN U16640 ( .A(n15570), .B(sreg[1655]), .Z(n15574) );
  NAND U16641 ( .A(n15572), .B(n15571), .Z(n15573) );
  NAND U16642 ( .A(n15574), .B(n15573), .Z(n15592) );
  XOR U16643 ( .A(n15593), .B(n15592), .Z(c[1656]) );
  NANDN U16644 ( .A(n15576), .B(n15575), .Z(n15580) );
  OR U16645 ( .A(n15578), .B(n15577), .Z(n15579) );
  AND U16646 ( .A(n15580), .B(n15579), .Z(n15598) );
  XOR U16647 ( .A(a[635]), .B(n2266), .Z(n15602) );
  AND U16648 ( .A(a[637]), .B(b[0]), .Z(n15582) );
  XNOR U16649 ( .A(n15582), .B(n2175), .Z(n15584) );
  NANDN U16650 ( .A(b[0]), .B(a[636]), .Z(n15583) );
  NAND U16651 ( .A(n15584), .B(n15583), .Z(n15607) );
  AND U16652 ( .A(a[633]), .B(b[3]), .Z(n15606) );
  XOR U16653 ( .A(n15607), .B(n15606), .Z(n15609) );
  XOR U16654 ( .A(n15608), .B(n15609), .Z(n15597) );
  NANDN U16655 ( .A(n15586), .B(n15585), .Z(n15590) );
  OR U16656 ( .A(n15588), .B(n15587), .Z(n15589) );
  AND U16657 ( .A(n15590), .B(n15589), .Z(n15596) );
  XOR U16658 ( .A(n15597), .B(n15596), .Z(n15599) );
  XOR U16659 ( .A(n15598), .B(n15599), .Z(n15612) );
  XNOR U16660 ( .A(n15612), .B(sreg[1657]), .Z(n15614) );
  NANDN U16661 ( .A(n15591), .B(sreg[1656]), .Z(n15595) );
  NAND U16662 ( .A(n15593), .B(n15592), .Z(n15594) );
  NAND U16663 ( .A(n15595), .B(n15594), .Z(n15613) );
  XOR U16664 ( .A(n15614), .B(n15613), .Z(c[1657]) );
  NANDN U16665 ( .A(n15597), .B(n15596), .Z(n15601) );
  OR U16666 ( .A(n15599), .B(n15598), .Z(n15600) );
  AND U16667 ( .A(n15601), .B(n15600), .Z(n15620) );
  XOR U16668 ( .A(a[636]), .B(n2267), .Z(n15621) );
  AND U16669 ( .A(b[0]), .B(a[638]), .Z(n15603) );
  XOR U16670 ( .A(b[1]), .B(n15603), .Z(n15605) );
  NAND U16671 ( .A(n23588), .B(a[637]), .Z(n15604) );
  AND U16672 ( .A(n15605), .B(n15604), .Z(n15625) );
  AND U16673 ( .A(a[634]), .B(b[3]), .Z(n15626) );
  XOR U16674 ( .A(n15625), .B(n15626), .Z(n15627) );
  XNOR U16675 ( .A(n15628), .B(n15627), .Z(n15617) );
  NANDN U16676 ( .A(n15607), .B(n15606), .Z(n15611) );
  OR U16677 ( .A(n15609), .B(n15608), .Z(n15610) );
  AND U16678 ( .A(n15611), .B(n15610), .Z(n15618) );
  XNOR U16679 ( .A(n15617), .B(n15618), .Z(n15619) );
  XNOR U16680 ( .A(n15620), .B(n15619), .Z(n15631) );
  XNOR U16681 ( .A(n15631), .B(sreg[1658]), .Z(n15633) );
  NANDN U16682 ( .A(n15612), .B(sreg[1657]), .Z(n15616) );
  NAND U16683 ( .A(n15614), .B(n15613), .Z(n15615) );
  NAND U16684 ( .A(n15616), .B(n15615), .Z(n15632) );
  XOR U16685 ( .A(n15633), .B(n15632), .Z(c[1658]) );
  XOR U16686 ( .A(a[637]), .B(n2267), .Z(n15640) );
  AND U16687 ( .A(a[639]), .B(b[0]), .Z(n15622) );
  XNOR U16688 ( .A(n15622), .B(n2175), .Z(n15624) );
  NANDN U16689 ( .A(b[0]), .B(a[638]), .Z(n15623) );
  NAND U16690 ( .A(n15624), .B(n15623), .Z(n15645) );
  AND U16691 ( .A(a[635]), .B(b[3]), .Z(n15644) );
  XOR U16692 ( .A(n15645), .B(n15644), .Z(n15647) );
  XOR U16693 ( .A(n15646), .B(n15647), .Z(n15635) );
  NAND U16694 ( .A(n15626), .B(n15625), .Z(n15630) );
  NANDN U16695 ( .A(n15628), .B(n15627), .Z(n15629) );
  AND U16696 ( .A(n15630), .B(n15629), .Z(n15634) );
  XOR U16697 ( .A(n15635), .B(n15634), .Z(n15637) );
  XOR U16698 ( .A(n15636), .B(n15637), .Z(n15650) );
  XNOR U16699 ( .A(n15650), .B(sreg[1659]), .Z(n15652) );
  XOR U16700 ( .A(n15652), .B(n15651), .Z(c[1659]) );
  NANDN U16701 ( .A(n15635), .B(n15634), .Z(n15639) );
  OR U16702 ( .A(n15637), .B(n15636), .Z(n15638) );
  AND U16703 ( .A(n15639), .B(n15638), .Z(n15657) );
  XOR U16704 ( .A(a[638]), .B(n2267), .Z(n15661) );
  AND U16705 ( .A(a[636]), .B(b[3]), .Z(n15665) );
  AND U16706 ( .A(a[640]), .B(b[0]), .Z(n15641) );
  XNOR U16707 ( .A(n15641), .B(n2175), .Z(n15643) );
  NANDN U16708 ( .A(b[0]), .B(a[639]), .Z(n15642) );
  NAND U16709 ( .A(n15643), .B(n15642), .Z(n15666) );
  XOR U16710 ( .A(n15665), .B(n15666), .Z(n15668) );
  XOR U16711 ( .A(n15667), .B(n15668), .Z(n15656) );
  NANDN U16712 ( .A(n15645), .B(n15644), .Z(n15649) );
  OR U16713 ( .A(n15647), .B(n15646), .Z(n15648) );
  AND U16714 ( .A(n15649), .B(n15648), .Z(n15655) );
  XOR U16715 ( .A(n15656), .B(n15655), .Z(n15658) );
  XOR U16716 ( .A(n15657), .B(n15658), .Z(n15671) );
  XNOR U16717 ( .A(n15671), .B(sreg[1660]), .Z(n15673) );
  NANDN U16718 ( .A(n15650), .B(sreg[1659]), .Z(n15654) );
  NAND U16719 ( .A(n15652), .B(n15651), .Z(n15653) );
  NAND U16720 ( .A(n15654), .B(n15653), .Z(n15672) );
  XOR U16721 ( .A(n15673), .B(n15672), .Z(c[1660]) );
  NANDN U16722 ( .A(n15656), .B(n15655), .Z(n15660) );
  OR U16723 ( .A(n15658), .B(n15657), .Z(n15659) );
  AND U16724 ( .A(n15660), .B(n15659), .Z(n15678) );
  XOR U16725 ( .A(a[639]), .B(n2267), .Z(n15682) );
  AND U16726 ( .A(a[641]), .B(b[0]), .Z(n15662) );
  XNOR U16727 ( .A(n15662), .B(n2175), .Z(n15664) );
  NANDN U16728 ( .A(b[0]), .B(a[640]), .Z(n15663) );
  NAND U16729 ( .A(n15664), .B(n15663), .Z(n15687) );
  AND U16730 ( .A(a[637]), .B(b[3]), .Z(n15686) );
  XOR U16731 ( .A(n15687), .B(n15686), .Z(n15689) );
  XOR U16732 ( .A(n15688), .B(n15689), .Z(n15677) );
  NANDN U16733 ( .A(n15666), .B(n15665), .Z(n15670) );
  OR U16734 ( .A(n15668), .B(n15667), .Z(n15669) );
  AND U16735 ( .A(n15670), .B(n15669), .Z(n15676) );
  XOR U16736 ( .A(n15677), .B(n15676), .Z(n15679) );
  XOR U16737 ( .A(n15678), .B(n15679), .Z(n15692) );
  XNOR U16738 ( .A(n15692), .B(sreg[1661]), .Z(n15694) );
  NANDN U16739 ( .A(n15671), .B(sreg[1660]), .Z(n15675) );
  NAND U16740 ( .A(n15673), .B(n15672), .Z(n15674) );
  NAND U16741 ( .A(n15675), .B(n15674), .Z(n15693) );
  XOR U16742 ( .A(n15694), .B(n15693), .Z(c[1661]) );
  NANDN U16743 ( .A(n15677), .B(n15676), .Z(n15681) );
  OR U16744 ( .A(n15679), .B(n15678), .Z(n15680) );
  AND U16745 ( .A(n15681), .B(n15680), .Z(n15699) );
  XOR U16746 ( .A(a[640]), .B(n2267), .Z(n15703) );
  AND U16747 ( .A(a[638]), .B(b[3]), .Z(n15707) );
  AND U16748 ( .A(a[642]), .B(b[0]), .Z(n15683) );
  XNOR U16749 ( .A(n15683), .B(n2175), .Z(n15685) );
  NANDN U16750 ( .A(b[0]), .B(a[641]), .Z(n15684) );
  NAND U16751 ( .A(n15685), .B(n15684), .Z(n15708) );
  XOR U16752 ( .A(n15707), .B(n15708), .Z(n15710) );
  XOR U16753 ( .A(n15709), .B(n15710), .Z(n15698) );
  NANDN U16754 ( .A(n15687), .B(n15686), .Z(n15691) );
  OR U16755 ( .A(n15689), .B(n15688), .Z(n15690) );
  AND U16756 ( .A(n15691), .B(n15690), .Z(n15697) );
  XOR U16757 ( .A(n15698), .B(n15697), .Z(n15700) );
  XOR U16758 ( .A(n15699), .B(n15700), .Z(n15713) );
  XNOR U16759 ( .A(n15713), .B(sreg[1662]), .Z(n15715) );
  NANDN U16760 ( .A(n15692), .B(sreg[1661]), .Z(n15696) );
  NAND U16761 ( .A(n15694), .B(n15693), .Z(n15695) );
  NAND U16762 ( .A(n15696), .B(n15695), .Z(n15714) );
  XOR U16763 ( .A(n15715), .B(n15714), .Z(c[1662]) );
  NANDN U16764 ( .A(n15698), .B(n15697), .Z(n15702) );
  OR U16765 ( .A(n15700), .B(n15699), .Z(n15701) );
  AND U16766 ( .A(n15702), .B(n15701), .Z(n15720) );
  XOR U16767 ( .A(a[641]), .B(n2267), .Z(n15724) );
  AND U16768 ( .A(a[643]), .B(b[0]), .Z(n15704) );
  XNOR U16769 ( .A(n15704), .B(n2175), .Z(n15706) );
  NANDN U16770 ( .A(b[0]), .B(a[642]), .Z(n15705) );
  NAND U16771 ( .A(n15706), .B(n15705), .Z(n15729) );
  AND U16772 ( .A(a[639]), .B(b[3]), .Z(n15728) );
  XOR U16773 ( .A(n15729), .B(n15728), .Z(n15731) );
  XOR U16774 ( .A(n15730), .B(n15731), .Z(n15719) );
  NANDN U16775 ( .A(n15708), .B(n15707), .Z(n15712) );
  OR U16776 ( .A(n15710), .B(n15709), .Z(n15711) );
  AND U16777 ( .A(n15712), .B(n15711), .Z(n15718) );
  XOR U16778 ( .A(n15719), .B(n15718), .Z(n15721) );
  XOR U16779 ( .A(n15720), .B(n15721), .Z(n15734) );
  XNOR U16780 ( .A(n15734), .B(sreg[1663]), .Z(n15736) );
  NANDN U16781 ( .A(n15713), .B(sreg[1662]), .Z(n15717) );
  NAND U16782 ( .A(n15715), .B(n15714), .Z(n15716) );
  NAND U16783 ( .A(n15717), .B(n15716), .Z(n15735) );
  XOR U16784 ( .A(n15736), .B(n15735), .Z(c[1663]) );
  NANDN U16785 ( .A(n15719), .B(n15718), .Z(n15723) );
  OR U16786 ( .A(n15721), .B(n15720), .Z(n15722) );
  AND U16787 ( .A(n15723), .B(n15722), .Z(n15741) );
  XOR U16788 ( .A(a[642]), .B(n2267), .Z(n15745) );
  AND U16789 ( .A(a[640]), .B(b[3]), .Z(n15749) );
  AND U16790 ( .A(a[644]), .B(b[0]), .Z(n15725) );
  XNOR U16791 ( .A(n15725), .B(n2175), .Z(n15727) );
  NANDN U16792 ( .A(b[0]), .B(a[643]), .Z(n15726) );
  NAND U16793 ( .A(n15727), .B(n15726), .Z(n15750) );
  XOR U16794 ( .A(n15749), .B(n15750), .Z(n15752) );
  XOR U16795 ( .A(n15751), .B(n15752), .Z(n15740) );
  NANDN U16796 ( .A(n15729), .B(n15728), .Z(n15733) );
  OR U16797 ( .A(n15731), .B(n15730), .Z(n15732) );
  AND U16798 ( .A(n15733), .B(n15732), .Z(n15739) );
  XOR U16799 ( .A(n15740), .B(n15739), .Z(n15742) );
  XOR U16800 ( .A(n15741), .B(n15742), .Z(n15755) );
  XNOR U16801 ( .A(n15755), .B(sreg[1664]), .Z(n15757) );
  NANDN U16802 ( .A(n15734), .B(sreg[1663]), .Z(n15738) );
  NAND U16803 ( .A(n15736), .B(n15735), .Z(n15737) );
  NAND U16804 ( .A(n15738), .B(n15737), .Z(n15756) );
  XOR U16805 ( .A(n15757), .B(n15756), .Z(c[1664]) );
  NANDN U16806 ( .A(n15740), .B(n15739), .Z(n15744) );
  OR U16807 ( .A(n15742), .B(n15741), .Z(n15743) );
  AND U16808 ( .A(n15744), .B(n15743), .Z(n15762) );
  XOR U16809 ( .A(a[643]), .B(n2268), .Z(n15766) );
  AND U16810 ( .A(a[645]), .B(b[0]), .Z(n15746) );
  XNOR U16811 ( .A(n15746), .B(n2175), .Z(n15748) );
  NANDN U16812 ( .A(b[0]), .B(a[644]), .Z(n15747) );
  NAND U16813 ( .A(n15748), .B(n15747), .Z(n15771) );
  AND U16814 ( .A(a[641]), .B(b[3]), .Z(n15770) );
  XOR U16815 ( .A(n15771), .B(n15770), .Z(n15773) );
  XOR U16816 ( .A(n15772), .B(n15773), .Z(n15761) );
  NANDN U16817 ( .A(n15750), .B(n15749), .Z(n15754) );
  OR U16818 ( .A(n15752), .B(n15751), .Z(n15753) );
  AND U16819 ( .A(n15754), .B(n15753), .Z(n15760) );
  XOR U16820 ( .A(n15761), .B(n15760), .Z(n15763) );
  XOR U16821 ( .A(n15762), .B(n15763), .Z(n15776) );
  XNOR U16822 ( .A(n15776), .B(sreg[1665]), .Z(n15778) );
  NANDN U16823 ( .A(n15755), .B(sreg[1664]), .Z(n15759) );
  NAND U16824 ( .A(n15757), .B(n15756), .Z(n15758) );
  NAND U16825 ( .A(n15759), .B(n15758), .Z(n15777) );
  XOR U16826 ( .A(n15778), .B(n15777), .Z(c[1665]) );
  NANDN U16827 ( .A(n15761), .B(n15760), .Z(n15765) );
  OR U16828 ( .A(n15763), .B(n15762), .Z(n15764) );
  AND U16829 ( .A(n15765), .B(n15764), .Z(n15783) );
  XOR U16830 ( .A(a[644]), .B(n2268), .Z(n15787) );
  AND U16831 ( .A(a[646]), .B(b[0]), .Z(n15767) );
  XNOR U16832 ( .A(n15767), .B(n2175), .Z(n15769) );
  NANDN U16833 ( .A(b[0]), .B(a[645]), .Z(n15768) );
  NAND U16834 ( .A(n15769), .B(n15768), .Z(n15792) );
  AND U16835 ( .A(a[642]), .B(b[3]), .Z(n15791) );
  XOR U16836 ( .A(n15792), .B(n15791), .Z(n15794) );
  XOR U16837 ( .A(n15793), .B(n15794), .Z(n15782) );
  NANDN U16838 ( .A(n15771), .B(n15770), .Z(n15775) );
  OR U16839 ( .A(n15773), .B(n15772), .Z(n15774) );
  AND U16840 ( .A(n15775), .B(n15774), .Z(n15781) );
  XOR U16841 ( .A(n15782), .B(n15781), .Z(n15784) );
  XOR U16842 ( .A(n15783), .B(n15784), .Z(n15797) );
  XNOR U16843 ( .A(n15797), .B(sreg[1666]), .Z(n15799) );
  NANDN U16844 ( .A(n15776), .B(sreg[1665]), .Z(n15780) );
  NAND U16845 ( .A(n15778), .B(n15777), .Z(n15779) );
  NAND U16846 ( .A(n15780), .B(n15779), .Z(n15798) );
  XOR U16847 ( .A(n15799), .B(n15798), .Z(c[1666]) );
  NANDN U16848 ( .A(n15782), .B(n15781), .Z(n15786) );
  OR U16849 ( .A(n15784), .B(n15783), .Z(n15785) );
  AND U16850 ( .A(n15786), .B(n15785), .Z(n15804) );
  XOR U16851 ( .A(a[645]), .B(n2268), .Z(n15808) );
  AND U16852 ( .A(a[647]), .B(b[0]), .Z(n15788) );
  XNOR U16853 ( .A(n15788), .B(n2175), .Z(n15790) );
  NANDN U16854 ( .A(b[0]), .B(a[646]), .Z(n15789) );
  NAND U16855 ( .A(n15790), .B(n15789), .Z(n15813) );
  AND U16856 ( .A(a[643]), .B(b[3]), .Z(n15812) );
  XOR U16857 ( .A(n15813), .B(n15812), .Z(n15815) );
  XOR U16858 ( .A(n15814), .B(n15815), .Z(n15803) );
  NANDN U16859 ( .A(n15792), .B(n15791), .Z(n15796) );
  OR U16860 ( .A(n15794), .B(n15793), .Z(n15795) );
  AND U16861 ( .A(n15796), .B(n15795), .Z(n15802) );
  XOR U16862 ( .A(n15803), .B(n15802), .Z(n15805) );
  XOR U16863 ( .A(n15804), .B(n15805), .Z(n15818) );
  XNOR U16864 ( .A(n15818), .B(sreg[1667]), .Z(n15820) );
  NANDN U16865 ( .A(n15797), .B(sreg[1666]), .Z(n15801) );
  NAND U16866 ( .A(n15799), .B(n15798), .Z(n15800) );
  NAND U16867 ( .A(n15801), .B(n15800), .Z(n15819) );
  XOR U16868 ( .A(n15820), .B(n15819), .Z(c[1667]) );
  NANDN U16869 ( .A(n15803), .B(n15802), .Z(n15807) );
  OR U16870 ( .A(n15805), .B(n15804), .Z(n15806) );
  AND U16871 ( .A(n15807), .B(n15806), .Z(n15825) );
  XOR U16872 ( .A(a[646]), .B(n2268), .Z(n15829) );
  AND U16873 ( .A(a[648]), .B(b[0]), .Z(n15809) );
  XNOR U16874 ( .A(n15809), .B(n2175), .Z(n15811) );
  NANDN U16875 ( .A(b[0]), .B(a[647]), .Z(n15810) );
  NAND U16876 ( .A(n15811), .B(n15810), .Z(n15834) );
  AND U16877 ( .A(a[644]), .B(b[3]), .Z(n15833) );
  XOR U16878 ( .A(n15834), .B(n15833), .Z(n15836) );
  XOR U16879 ( .A(n15835), .B(n15836), .Z(n15824) );
  NANDN U16880 ( .A(n15813), .B(n15812), .Z(n15817) );
  OR U16881 ( .A(n15815), .B(n15814), .Z(n15816) );
  AND U16882 ( .A(n15817), .B(n15816), .Z(n15823) );
  XOR U16883 ( .A(n15824), .B(n15823), .Z(n15826) );
  XOR U16884 ( .A(n15825), .B(n15826), .Z(n15839) );
  XNOR U16885 ( .A(n15839), .B(sreg[1668]), .Z(n15841) );
  NANDN U16886 ( .A(n15818), .B(sreg[1667]), .Z(n15822) );
  NAND U16887 ( .A(n15820), .B(n15819), .Z(n15821) );
  NAND U16888 ( .A(n15822), .B(n15821), .Z(n15840) );
  XOR U16889 ( .A(n15841), .B(n15840), .Z(c[1668]) );
  NANDN U16890 ( .A(n15824), .B(n15823), .Z(n15828) );
  OR U16891 ( .A(n15826), .B(n15825), .Z(n15827) );
  AND U16892 ( .A(n15828), .B(n15827), .Z(n15846) );
  XOR U16893 ( .A(a[647]), .B(n2268), .Z(n15850) );
  AND U16894 ( .A(a[649]), .B(b[0]), .Z(n15830) );
  XNOR U16895 ( .A(n15830), .B(n2175), .Z(n15832) );
  NANDN U16896 ( .A(b[0]), .B(a[648]), .Z(n15831) );
  NAND U16897 ( .A(n15832), .B(n15831), .Z(n15855) );
  AND U16898 ( .A(a[645]), .B(b[3]), .Z(n15854) );
  XOR U16899 ( .A(n15855), .B(n15854), .Z(n15857) );
  XOR U16900 ( .A(n15856), .B(n15857), .Z(n15845) );
  NANDN U16901 ( .A(n15834), .B(n15833), .Z(n15838) );
  OR U16902 ( .A(n15836), .B(n15835), .Z(n15837) );
  AND U16903 ( .A(n15838), .B(n15837), .Z(n15844) );
  XOR U16904 ( .A(n15845), .B(n15844), .Z(n15847) );
  XOR U16905 ( .A(n15846), .B(n15847), .Z(n15860) );
  XNOR U16906 ( .A(n15860), .B(sreg[1669]), .Z(n15862) );
  NANDN U16907 ( .A(n15839), .B(sreg[1668]), .Z(n15843) );
  NAND U16908 ( .A(n15841), .B(n15840), .Z(n15842) );
  NAND U16909 ( .A(n15843), .B(n15842), .Z(n15861) );
  XOR U16910 ( .A(n15862), .B(n15861), .Z(c[1669]) );
  NANDN U16911 ( .A(n15845), .B(n15844), .Z(n15849) );
  OR U16912 ( .A(n15847), .B(n15846), .Z(n15848) );
  AND U16913 ( .A(n15849), .B(n15848), .Z(n15867) );
  XOR U16914 ( .A(a[648]), .B(n2268), .Z(n15871) );
  AND U16915 ( .A(a[650]), .B(b[0]), .Z(n15851) );
  XNOR U16916 ( .A(n15851), .B(n2175), .Z(n15853) );
  NANDN U16917 ( .A(b[0]), .B(a[649]), .Z(n15852) );
  NAND U16918 ( .A(n15853), .B(n15852), .Z(n15876) );
  AND U16919 ( .A(a[646]), .B(b[3]), .Z(n15875) );
  XOR U16920 ( .A(n15876), .B(n15875), .Z(n15878) );
  XOR U16921 ( .A(n15877), .B(n15878), .Z(n15866) );
  NANDN U16922 ( .A(n15855), .B(n15854), .Z(n15859) );
  OR U16923 ( .A(n15857), .B(n15856), .Z(n15858) );
  AND U16924 ( .A(n15859), .B(n15858), .Z(n15865) );
  XOR U16925 ( .A(n15866), .B(n15865), .Z(n15868) );
  XOR U16926 ( .A(n15867), .B(n15868), .Z(n15881) );
  XNOR U16927 ( .A(n15881), .B(sreg[1670]), .Z(n15883) );
  NANDN U16928 ( .A(n15860), .B(sreg[1669]), .Z(n15864) );
  NAND U16929 ( .A(n15862), .B(n15861), .Z(n15863) );
  NAND U16930 ( .A(n15864), .B(n15863), .Z(n15882) );
  XOR U16931 ( .A(n15883), .B(n15882), .Z(c[1670]) );
  NANDN U16932 ( .A(n15866), .B(n15865), .Z(n15870) );
  OR U16933 ( .A(n15868), .B(n15867), .Z(n15869) );
  AND U16934 ( .A(n15870), .B(n15869), .Z(n15888) );
  XOR U16935 ( .A(a[649]), .B(n2268), .Z(n15892) );
  AND U16936 ( .A(a[647]), .B(b[3]), .Z(n15896) );
  AND U16937 ( .A(a[651]), .B(b[0]), .Z(n15872) );
  XNOR U16938 ( .A(n15872), .B(n2175), .Z(n15874) );
  NANDN U16939 ( .A(b[0]), .B(a[650]), .Z(n15873) );
  NAND U16940 ( .A(n15874), .B(n15873), .Z(n15897) );
  XOR U16941 ( .A(n15896), .B(n15897), .Z(n15899) );
  XOR U16942 ( .A(n15898), .B(n15899), .Z(n15887) );
  NANDN U16943 ( .A(n15876), .B(n15875), .Z(n15880) );
  OR U16944 ( .A(n15878), .B(n15877), .Z(n15879) );
  AND U16945 ( .A(n15880), .B(n15879), .Z(n15886) );
  XOR U16946 ( .A(n15887), .B(n15886), .Z(n15889) );
  XOR U16947 ( .A(n15888), .B(n15889), .Z(n15902) );
  XNOR U16948 ( .A(n15902), .B(sreg[1671]), .Z(n15904) );
  NANDN U16949 ( .A(n15881), .B(sreg[1670]), .Z(n15885) );
  NAND U16950 ( .A(n15883), .B(n15882), .Z(n15884) );
  NAND U16951 ( .A(n15885), .B(n15884), .Z(n15903) );
  XOR U16952 ( .A(n15904), .B(n15903), .Z(c[1671]) );
  NANDN U16953 ( .A(n15887), .B(n15886), .Z(n15891) );
  OR U16954 ( .A(n15889), .B(n15888), .Z(n15890) );
  AND U16955 ( .A(n15891), .B(n15890), .Z(n15909) );
  XOR U16956 ( .A(a[650]), .B(n2269), .Z(n15913) );
  AND U16957 ( .A(a[652]), .B(b[0]), .Z(n15893) );
  XNOR U16958 ( .A(n15893), .B(n2175), .Z(n15895) );
  NANDN U16959 ( .A(b[0]), .B(a[651]), .Z(n15894) );
  NAND U16960 ( .A(n15895), .B(n15894), .Z(n15918) );
  AND U16961 ( .A(a[648]), .B(b[3]), .Z(n15917) );
  XOR U16962 ( .A(n15918), .B(n15917), .Z(n15920) );
  XOR U16963 ( .A(n15919), .B(n15920), .Z(n15908) );
  NANDN U16964 ( .A(n15897), .B(n15896), .Z(n15901) );
  OR U16965 ( .A(n15899), .B(n15898), .Z(n15900) );
  AND U16966 ( .A(n15901), .B(n15900), .Z(n15907) );
  XOR U16967 ( .A(n15908), .B(n15907), .Z(n15910) );
  XOR U16968 ( .A(n15909), .B(n15910), .Z(n15923) );
  XNOR U16969 ( .A(n15923), .B(sreg[1672]), .Z(n15925) );
  NANDN U16970 ( .A(n15902), .B(sreg[1671]), .Z(n15906) );
  NAND U16971 ( .A(n15904), .B(n15903), .Z(n15905) );
  NAND U16972 ( .A(n15906), .B(n15905), .Z(n15924) );
  XOR U16973 ( .A(n15925), .B(n15924), .Z(c[1672]) );
  NANDN U16974 ( .A(n15908), .B(n15907), .Z(n15912) );
  OR U16975 ( .A(n15910), .B(n15909), .Z(n15911) );
  AND U16976 ( .A(n15912), .B(n15911), .Z(n15930) );
  XOR U16977 ( .A(a[651]), .B(n2269), .Z(n15934) );
  AND U16978 ( .A(a[653]), .B(b[0]), .Z(n15914) );
  XNOR U16979 ( .A(n15914), .B(n2175), .Z(n15916) );
  NANDN U16980 ( .A(b[0]), .B(a[652]), .Z(n15915) );
  NAND U16981 ( .A(n15916), .B(n15915), .Z(n15939) );
  AND U16982 ( .A(a[649]), .B(b[3]), .Z(n15938) );
  XOR U16983 ( .A(n15939), .B(n15938), .Z(n15941) );
  XOR U16984 ( .A(n15940), .B(n15941), .Z(n15929) );
  NANDN U16985 ( .A(n15918), .B(n15917), .Z(n15922) );
  OR U16986 ( .A(n15920), .B(n15919), .Z(n15921) );
  AND U16987 ( .A(n15922), .B(n15921), .Z(n15928) );
  XOR U16988 ( .A(n15929), .B(n15928), .Z(n15931) );
  XOR U16989 ( .A(n15930), .B(n15931), .Z(n15944) );
  XNOR U16990 ( .A(n15944), .B(sreg[1673]), .Z(n15946) );
  NANDN U16991 ( .A(n15923), .B(sreg[1672]), .Z(n15927) );
  NAND U16992 ( .A(n15925), .B(n15924), .Z(n15926) );
  NAND U16993 ( .A(n15927), .B(n15926), .Z(n15945) );
  XOR U16994 ( .A(n15946), .B(n15945), .Z(c[1673]) );
  NANDN U16995 ( .A(n15929), .B(n15928), .Z(n15933) );
  OR U16996 ( .A(n15931), .B(n15930), .Z(n15932) );
  AND U16997 ( .A(n15933), .B(n15932), .Z(n15951) );
  XOR U16998 ( .A(a[652]), .B(n2269), .Z(n15955) );
  AND U16999 ( .A(a[650]), .B(b[3]), .Z(n15959) );
  AND U17000 ( .A(a[654]), .B(b[0]), .Z(n15935) );
  XNOR U17001 ( .A(n15935), .B(n2175), .Z(n15937) );
  NANDN U17002 ( .A(b[0]), .B(a[653]), .Z(n15936) );
  NAND U17003 ( .A(n15937), .B(n15936), .Z(n15960) );
  XOR U17004 ( .A(n15959), .B(n15960), .Z(n15962) );
  XOR U17005 ( .A(n15961), .B(n15962), .Z(n15950) );
  NANDN U17006 ( .A(n15939), .B(n15938), .Z(n15943) );
  OR U17007 ( .A(n15941), .B(n15940), .Z(n15942) );
  AND U17008 ( .A(n15943), .B(n15942), .Z(n15949) );
  XOR U17009 ( .A(n15950), .B(n15949), .Z(n15952) );
  XOR U17010 ( .A(n15951), .B(n15952), .Z(n15965) );
  XNOR U17011 ( .A(n15965), .B(sreg[1674]), .Z(n15967) );
  NANDN U17012 ( .A(n15944), .B(sreg[1673]), .Z(n15948) );
  NAND U17013 ( .A(n15946), .B(n15945), .Z(n15947) );
  NAND U17014 ( .A(n15948), .B(n15947), .Z(n15966) );
  XOR U17015 ( .A(n15967), .B(n15966), .Z(c[1674]) );
  NANDN U17016 ( .A(n15950), .B(n15949), .Z(n15954) );
  OR U17017 ( .A(n15952), .B(n15951), .Z(n15953) );
  AND U17018 ( .A(n15954), .B(n15953), .Z(n15972) );
  XOR U17019 ( .A(a[653]), .B(n2269), .Z(n15976) );
  AND U17020 ( .A(a[655]), .B(b[0]), .Z(n15956) );
  XNOR U17021 ( .A(n15956), .B(n2175), .Z(n15958) );
  NANDN U17022 ( .A(b[0]), .B(a[654]), .Z(n15957) );
  NAND U17023 ( .A(n15958), .B(n15957), .Z(n15981) );
  AND U17024 ( .A(a[651]), .B(b[3]), .Z(n15980) );
  XOR U17025 ( .A(n15981), .B(n15980), .Z(n15983) );
  XOR U17026 ( .A(n15982), .B(n15983), .Z(n15971) );
  NANDN U17027 ( .A(n15960), .B(n15959), .Z(n15964) );
  OR U17028 ( .A(n15962), .B(n15961), .Z(n15963) );
  AND U17029 ( .A(n15964), .B(n15963), .Z(n15970) );
  XOR U17030 ( .A(n15971), .B(n15970), .Z(n15973) );
  XOR U17031 ( .A(n15972), .B(n15973), .Z(n15986) );
  XNOR U17032 ( .A(n15986), .B(sreg[1675]), .Z(n15988) );
  NANDN U17033 ( .A(n15965), .B(sreg[1674]), .Z(n15969) );
  NAND U17034 ( .A(n15967), .B(n15966), .Z(n15968) );
  NAND U17035 ( .A(n15969), .B(n15968), .Z(n15987) );
  XOR U17036 ( .A(n15988), .B(n15987), .Z(c[1675]) );
  NANDN U17037 ( .A(n15971), .B(n15970), .Z(n15975) );
  OR U17038 ( .A(n15973), .B(n15972), .Z(n15974) );
  AND U17039 ( .A(n15975), .B(n15974), .Z(n15993) );
  XOR U17040 ( .A(a[654]), .B(n2269), .Z(n15997) );
  AND U17041 ( .A(a[656]), .B(b[0]), .Z(n15977) );
  XNOR U17042 ( .A(n15977), .B(n2175), .Z(n15979) );
  NANDN U17043 ( .A(b[0]), .B(a[655]), .Z(n15978) );
  NAND U17044 ( .A(n15979), .B(n15978), .Z(n16002) );
  AND U17045 ( .A(a[652]), .B(b[3]), .Z(n16001) );
  XOR U17046 ( .A(n16002), .B(n16001), .Z(n16004) );
  XOR U17047 ( .A(n16003), .B(n16004), .Z(n15992) );
  NANDN U17048 ( .A(n15981), .B(n15980), .Z(n15985) );
  OR U17049 ( .A(n15983), .B(n15982), .Z(n15984) );
  AND U17050 ( .A(n15985), .B(n15984), .Z(n15991) );
  XOR U17051 ( .A(n15992), .B(n15991), .Z(n15994) );
  XOR U17052 ( .A(n15993), .B(n15994), .Z(n16007) );
  XNOR U17053 ( .A(n16007), .B(sreg[1676]), .Z(n16009) );
  NANDN U17054 ( .A(n15986), .B(sreg[1675]), .Z(n15990) );
  NAND U17055 ( .A(n15988), .B(n15987), .Z(n15989) );
  NAND U17056 ( .A(n15990), .B(n15989), .Z(n16008) );
  XOR U17057 ( .A(n16009), .B(n16008), .Z(c[1676]) );
  NANDN U17058 ( .A(n15992), .B(n15991), .Z(n15996) );
  OR U17059 ( .A(n15994), .B(n15993), .Z(n15995) );
  AND U17060 ( .A(n15996), .B(n15995), .Z(n16014) );
  XOR U17061 ( .A(a[655]), .B(n2269), .Z(n16018) );
  AND U17062 ( .A(a[657]), .B(b[0]), .Z(n15998) );
  XNOR U17063 ( .A(n15998), .B(n2175), .Z(n16000) );
  NANDN U17064 ( .A(b[0]), .B(a[656]), .Z(n15999) );
  NAND U17065 ( .A(n16000), .B(n15999), .Z(n16023) );
  AND U17066 ( .A(a[653]), .B(b[3]), .Z(n16022) );
  XOR U17067 ( .A(n16023), .B(n16022), .Z(n16025) );
  XOR U17068 ( .A(n16024), .B(n16025), .Z(n16013) );
  NANDN U17069 ( .A(n16002), .B(n16001), .Z(n16006) );
  OR U17070 ( .A(n16004), .B(n16003), .Z(n16005) );
  AND U17071 ( .A(n16006), .B(n16005), .Z(n16012) );
  XOR U17072 ( .A(n16013), .B(n16012), .Z(n16015) );
  XOR U17073 ( .A(n16014), .B(n16015), .Z(n16028) );
  XNOR U17074 ( .A(n16028), .B(sreg[1677]), .Z(n16030) );
  NANDN U17075 ( .A(n16007), .B(sreg[1676]), .Z(n16011) );
  NAND U17076 ( .A(n16009), .B(n16008), .Z(n16010) );
  NAND U17077 ( .A(n16011), .B(n16010), .Z(n16029) );
  XOR U17078 ( .A(n16030), .B(n16029), .Z(c[1677]) );
  NANDN U17079 ( .A(n16013), .B(n16012), .Z(n16017) );
  OR U17080 ( .A(n16015), .B(n16014), .Z(n16016) );
  AND U17081 ( .A(n16017), .B(n16016), .Z(n16035) );
  XOR U17082 ( .A(a[656]), .B(n2269), .Z(n16039) );
  AND U17083 ( .A(a[654]), .B(b[3]), .Z(n16043) );
  AND U17084 ( .A(a[658]), .B(b[0]), .Z(n16019) );
  XNOR U17085 ( .A(n16019), .B(n2175), .Z(n16021) );
  NANDN U17086 ( .A(b[0]), .B(a[657]), .Z(n16020) );
  NAND U17087 ( .A(n16021), .B(n16020), .Z(n16044) );
  XOR U17088 ( .A(n16043), .B(n16044), .Z(n16046) );
  XOR U17089 ( .A(n16045), .B(n16046), .Z(n16034) );
  NANDN U17090 ( .A(n16023), .B(n16022), .Z(n16027) );
  OR U17091 ( .A(n16025), .B(n16024), .Z(n16026) );
  AND U17092 ( .A(n16027), .B(n16026), .Z(n16033) );
  XOR U17093 ( .A(n16034), .B(n16033), .Z(n16036) );
  XOR U17094 ( .A(n16035), .B(n16036), .Z(n16049) );
  XNOR U17095 ( .A(n16049), .B(sreg[1678]), .Z(n16051) );
  NANDN U17096 ( .A(n16028), .B(sreg[1677]), .Z(n16032) );
  NAND U17097 ( .A(n16030), .B(n16029), .Z(n16031) );
  NAND U17098 ( .A(n16032), .B(n16031), .Z(n16050) );
  XOR U17099 ( .A(n16051), .B(n16050), .Z(c[1678]) );
  NANDN U17100 ( .A(n16034), .B(n16033), .Z(n16038) );
  OR U17101 ( .A(n16036), .B(n16035), .Z(n16037) );
  AND U17102 ( .A(n16038), .B(n16037), .Z(n16056) );
  XOR U17103 ( .A(a[657]), .B(n2270), .Z(n16060) );
  AND U17104 ( .A(a[659]), .B(b[0]), .Z(n16040) );
  XNOR U17105 ( .A(n16040), .B(n2175), .Z(n16042) );
  NANDN U17106 ( .A(b[0]), .B(a[658]), .Z(n16041) );
  NAND U17107 ( .A(n16042), .B(n16041), .Z(n16065) );
  AND U17108 ( .A(a[655]), .B(b[3]), .Z(n16064) );
  XOR U17109 ( .A(n16065), .B(n16064), .Z(n16067) );
  XOR U17110 ( .A(n16066), .B(n16067), .Z(n16055) );
  NANDN U17111 ( .A(n16044), .B(n16043), .Z(n16048) );
  OR U17112 ( .A(n16046), .B(n16045), .Z(n16047) );
  AND U17113 ( .A(n16048), .B(n16047), .Z(n16054) );
  XOR U17114 ( .A(n16055), .B(n16054), .Z(n16057) );
  XOR U17115 ( .A(n16056), .B(n16057), .Z(n16070) );
  XNOR U17116 ( .A(n16070), .B(sreg[1679]), .Z(n16072) );
  NANDN U17117 ( .A(n16049), .B(sreg[1678]), .Z(n16053) );
  NAND U17118 ( .A(n16051), .B(n16050), .Z(n16052) );
  NAND U17119 ( .A(n16053), .B(n16052), .Z(n16071) );
  XOR U17120 ( .A(n16072), .B(n16071), .Z(c[1679]) );
  NANDN U17121 ( .A(n16055), .B(n16054), .Z(n16059) );
  OR U17122 ( .A(n16057), .B(n16056), .Z(n16058) );
  AND U17123 ( .A(n16059), .B(n16058), .Z(n16077) );
  XOR U17124 ( .A(a[658]), .B(n2270), .Z(n16081) );
  AND U17125 ( .A(a[660]), .B(b[0]), .Z(n16061) );
  XNOR U17126 ( .A(n16061), .B(n2175), .Z(n16063) );
  NANDN U17127 ( .A(b[0]), .B(a[659]), .Z(n16062) );
  NAND U17128 ( .A(n16063), .B(n16062), .Z(n16086) );
  AND U17129 ( .A(a[656]), .B(b[3]), .Z(n16085) );
  XOR U17130 ( .A(n16086), .B(n16085), .Z(n16088) );
  XOR U17131 ( .A(n16087), .B(n16088), .Z(n16076) );
  NANDN U17132 ( .A(n16065), .B(n16064), .Z(n16069) );
  OR U17133 ( .A(n16067), .B(n16066), .Z(n16068) );
  AND U17134 ( .A(n16069), .B(n16068), .Z(n16075) );
  XOR U17135 ( .A(n16076), .B(n16075), .Z(n16078) );
  XOR U17136 ( .A(n16077), .B(n16078), .Z(n16091) );
  XNOR U17137 ( .A(n16091), .B(sreg[1680]), .Z(n16093) );
  NANDN U17138 ( .A(n16070), .B(sreg[1679]), .Z(n16074) );
  NAND U17139 ( .A(n16072), .B(n16071), .Z(n16073) );
  NAND U17140 ( .A(n16074), .B(n16073), .Z(n16092) );
  XOR U17141 ( .A(n16093), .B(n16092), .Z(c[1680]) );
  NANDN U17142 ( .A(n16076), .B(n16075), .Z(n16080) );
  OR U17143 ( .A(n16078), .B(n16077), .Z(n16079) );
  AND U17144 ( .A(n16080), .B(n16079), .Z(n16098) );
  XOR U17145 ( .A(a[659]), .B(n2270), .Z(n16102) );
  AND U17146 ( .A(a[657]), .B(b[3]), .Z(n16106) );
  AND U17147 ( .A(a[661]), .B(b[0]), .Z(n16082) );
  XNOR U17148 ( .A(n16082), .B(n2175), .Z(n16084) );
  NANDN U17149 ( .A(b[0]), .B(a[660]), .Z(n16083) );
  NAND U17150 ( .A(n16084), .B(n16083), .Z(n16107) );
  XOR U17151 ( .A(n16106), .B(n16107), .Z(n16109) );
  XOR U17152 ( .A(n16108), .B(n16109), .Z(n16097) );
  NANDN U17153 ( .A(n16086), .B(n16085), .Z(n16090) );
  OR U17154 ( .A(n16088), .B(n16087), .Z(n16089) );
  AND U17155 ( .A(n16090), .B(n16089), .Z(n16096) );
  XOR U17156 ( .A(n16097), .B(n16096), .Z(n16099) );
  XOR U17157 ( .A(n16098), .B(n16099), .Z(n16112) );
  XNOR U17158 ( .A(n16112), .B(sreg[1681]), .Z(n16114) );
  NANDN U17159 ( .A(n16091), .B(sreg[1680]), .Z(n16095) );
  NAND U17160 ( .A(n16093), .B(n16092), .Z(n16094) );
  NAND U17161 ( .A(n16095), .B(n16094), .Z(n16113) );
  XOR U17162 ( .A(n16114), .B(n16113), .Z(c[1681]) );
  NANDN U17163 ( .A(n16097), .B(n16096), .Z(n16101) );
  OR U17164 ( .A(n16099), .B(n16098), .Z(n16100) );
  AND U17165 ( .A(n16101), .B(n16100), .Z(n16119) );
  XOR U17166 ( .A(a[660]), .B(n2270), .Z(n16123) );
  AND U17167 ( .A(a[662]), .B(b[0]), .Z(n16103) );
  XNOR U17168 ( .A(n16103), .B(n2175), .Z(n16105) );
  NANDN U17169 ( .A(b[0]), .B(a[661]), .Z(n16104) );
  NAND U17170 ( .A(n16105), .B(n16104), .Z(n16128) );
  AND U17171 ( .A(a[658]), .B(b[3]), .Z(n16127) );
  XOR U17172 ( .A(n16128), .B(n16127), .Z(n16130) );
  XOR U17173 ( .A(n16129), .B(n16130), .Z(n16118) );
  NANDN U17174 ( .A(n16107), .B(n16106), .Z(n16111) );
  OR U17175 ( .A(n16109), .B(n16108), .Z(n16110) );
  AND U17176 ( .A(n16111), .B(n16110), .Z(n16117) );
  XOR U17177 ( .A(n16118), .B(n16117), .Z(n16120) );
  XOR U17178 ( .A(n16119), .B(n16120), .Z(n16133) );
  XNOR U17179 ( .A(n16133), .B(sreg[1682]), .Z(n16135) );
  NANDN U17180 ( .A(n16112), .B(sreg[1681]), .Z(n16116) );
  NAND U17181 ( .A(n16114), .B(n16113), .Z(n16115) );
  NAND U17182 ( .A(n16116), .B(n16115), .Z(n16134) );
  XOR U17183 ( .A(n16135), .B(n16134), .Z(c[1682]) );
  NANDN U17184 ( .A(n16118), .B(n16117), .Z(n16122) );
  OR U17185 ( .A(n16120), .B(n16119), .Z(n16121) );
  AND U17186 ( .A(n16122), .B(n16121), .Z(n16140) );
  XOR U17187 ( .A(a[661]), .B(n2270), .Z(n16144) );
  AND U17188 ( .A(a[659]), .B(b[3]), .Z(n16148) );
  AND U17189 ( .A(a[663]), .B(b[0]), .Z(n16124) );
  XNOR U17190 ( .A(n16124), .B(n2175), .Z(n16126) );
  NANDN U17191 ( .A(b[0]), .B(a[662]), .Z(n16125) );
  NAND U17192 ( .A(n16126), .B(n16125), .Z(n16149) );
  XOR U17193 ( .A(n16148), .B(n16149), .Z(n16151) );
  XOR U17194 ( .A(n16150), .B(n16151), .Z(n16139) );
  NANDN U17195 ( .A(n16128), .B(n16127), .Z(n16132) );
  OR U17196 ( .A(n16130), .B(n16129), .Z(n16131) );
  AND U17197 ( .A(n16132), .B(n16131), .Z(n16138) );
  XOR U17198 ( .A(n16139), .B(n16138), .Z(n16141) );
  XOR U17199 ( .A(n16140), .B(n16141), .Z(n16154) );
  XNOR U17200 ( .A(n16154), .B(sreg[1683]), .Z(n16156) );
  NANDN U17201 ( .A(n16133), .B(sreg[1682]), .Z(n16137) );
  NAND U17202 ( .A(n16135), .B(n16134), .Z(n16136) );
  NAND U17203 ( .A(n16137), .B(n16136), .Z(n16155) );
  XOR U17204 ( .A(n16156), .B(n16155), .Z(c[1683]) );
  NANDN U17205 ( .A(n16139), .B(n16138), .Z(n16143) );
  OR U17206 ( .A(n16141), .B(n16140), .Z(n16142) );
  AND U17207 ( .A(n16143), .B(n16142), .Z(n16161) );
  XOR U17208 ( .A(a[662]), .B(n2270), .Z(n16165) );
  AND U17209 ( .A(a[664]), .B(b[0]), .Z(n16145) );
  XNOR U17210 ( .A(n16145), .B(n2175), .Z(n16147) );
  NANDN U17211 ( .A(b[0]), .B(a[663]), .Z(n16146) );
  NAND U17212 ( .A(n16147), .B(n16146), .Z(n16170) );
  AND U17213 ( .A(a[660]), .B(b[3]), .Z(n16169) );
  XOR U17214 ( .A(n16170), .B(n16169), .Z(n16172) );
  XOR U17215 ( .A(n16171), .B(n16172), .Z(n16160) );
  NANDN U17216 ( .A(n16149), .B(n16148), .Z(n16153) );
  OR U17217 ( .A(n16151), .B(n16150), .Z(n16152) );
  AND U17218 ( .A(n16153), .B(n16152), .Z(n16159) );
  XOR U17219 ( .A(n16160), .B(n16159), .Z(n16162) );
  XOR U17220 ( .A(n16161), .B(n16162), .Z(n16175) );
  XNOR U17221 ( .A(n16175), .B(sreg[1684]), .Z(n16177) );
  NANDN U17222 ( .A(n16154), .B(sreg[1683]), .Z(n16158) );
  NAND U17223 ( .A(n16156), .B(n16155), .Z(n16157) );
  NAND U17224 ( .A(n16158), .B(n16157), .Z(n16176) );
  XOR U17225 ( .A(n16177), .B(n16176), .Z(c[1684]) );
  NANDN U17226 ( .A(n16160), .B(n16159), .Z(n16164) );
  OR U17227 ( .A(n16162), .B(n16161), .Z(n16163) );
  AND U17228 ( .A(n16164), .B(n16163), .Z(n16182) );
  XOR U17229 ( .A(a[663]), .B(n2270), .Z(n16186) );
  AND U17230 ( .A(a[661]), .B(b[3]), .Z(n16190) );
  AND U17231 ( .A(a[665]), .B(b[0]), .Z(n16166) );
  XNOR U17232 ( .A(n16166), .B(n2175), .Z(n16168) );
  NANDN U17233 ( .A(b[0]), .B(a[664]), .Z(n16167) );
  NAND U17234 ( .A(n16168), .B(n16167), .Z(n16191) );
  XOR U17235 ( .A(n16190), .B(n16191), .Z(n16193) );
  XOR U17236 ( .A(n16192), .B(n16193), .Z(n16181) );
  NANDN U17237 ( .A(n16170), .B(n16169), .Z(n16174) );
  OR U17238 ( .A(n16172), .B(n16171), .Z(n16173) );
  AND U17239 ( .A(n16174), .B(n16173), .Z(n16180) );
  XOR U17240 ( .A(n16181), .B(n16180), .Z(n16183) );
  XOR U17241 ( .A(n16182), .B(n16183), .Z(n16196) );
  XNOR U17242 ( .A(n16196), .B(sreg[1685]), .Z(n16198) );
  NANDN U17243 ( .A(n16175), .B(sreg[1684]), .Z(n16179) );
  NAND U17244 ( .A(n16177), .B(n16176), .Z(n16178) );
  NAND U17245 ( .A(n16179), .B(n16178), .Z(n16197) );
  XOR U17246 ( .A(n16198), .B(n16197), .Z(c[1685]) );
  NANDN U17247 ( .A(n16181), .B(n16180), .Z(n16185) );
  OR U17248 ( .A(n16183), .B(n16182), .Z(n16184) );
  AND U17249 ( .A(n16185), .B(n16184), .Z(n16203) );
  XOR U17250 ( .A(a[664]), .B(n2271), .Z(n16207) );
  AND U17251 ( .A(a[666]), .B(b[0]), .Z(n16187) );
  XNOR U17252 ( .A(n16187), .B(n2175), .Z(n16189) );
  NANDN U17253 ( .A(b[0]), .B(a[665]), .Z(n16188) );
  NAND U17254 ( .A(n16189), .B(n16188), .Z(n16212) );
  AND U17255 ( .A(a[662]), .B(b[3]), .Z(n16211) );
  XOR U17256 ( .A(n16212), .B(n16211), .Z(n16214) );
  XOR U17257 ( .A(n16213), .B(n16214), .Z(n16202) );
  NANDN U17258 ( .A(n16191), .B(n16190), .Z(n16195) );
  OR U17259 ( .A(n16193), .B(n16192), .Z(n16194) );
  AND U17260 ( .A(n16195), .B(n16194), .Z(n16201) );
  XOR U17261 ( .A(n16202), .B(n16201), .Z(n16204) );
  XOR U17262 ( .A(n16203), .B(n16204), .Z(n16217) );
  XNOR U17263 ( .A(n16217), .B(sreg[1686]), .Z(n16219) );
  NANDN U17264 ( .A(n16196), .B(sreg[1685]), .Z(n16200) );
  NAND U17265 ( .A(n16198), .B(n16197), .Z(n16199) );
  NAND U17266 ( .A(n16200), .B(n16199), .Z(n16218) );
  XOR U17267 ( .A(n16219), .B(n16218), .Z(c[1686]) );
  NANDN U17268 ( .A(n16202), .B(n16201), .Z(n16206) );
  OR U17269 ( .A(n16204), .B(n16203), .Z(n16205) );
  AND U17270 ( .A(n16206), .B(n16205), .Z(n16224) );
  XOR U17271 ( .A(a[665]), .B(n2271), .Z(n16228) );
  AND U17272 ( .A(a[663]), .B(b[3]), .Z(n16232) );
  AND U17273 ( .A(a[667]), .B(b[0]), .Z(n16208) );
  XNOR U17274 ( .A(n16208), .B(n2175), .Z(n16210) );
  NANDN U17275 ( .A(b[0]), .B(a[666]), .Z(n16209) );
  NAND U17276 ( .A(n16210), .B(n16209), .Z(n16233) );
  XOR U17277 ( .A(n16232), .B(n16233), .Z(n16235) );
  XOR U17278 ( .A(n16234), .B(n16235), .Z(n16223) );
  NANDN U17279 ( .A(n16212), .B(n16211), .Z(n16216) );
  OR U17280 ( .A(n16214), .B(n16213), .Z(n16215) );
  AND U17281 ( .A(n16216), .B(n16215), .Z(n16222) );
  XOR U17282 ( .A(n16223), .B(n16222), .Z(n16225) );
  XOR U17283 ( .A(n16224), .B(n16225), .Z(n16238) );
  XNOR U17284 ( .A(n16238), .B(sreg[1687]), .Z(n16240) );
  NANDN U17285 ( .A(n16217), .B(sreg[1686]), .Z(n16221) );
  NAND U17286 ( .A(n16219), .B(n16218), .Z(n16220) );
  NAND U17287 ( .A(n16221), .B(n16220), .Z(n16239) );
  XOR U17288 ( .A(n16240), .B(n16239), .Z(c[1687]) );
  NANDN U17289 ( .A(n16223), .B(n16222), .Z(n16227) );
  OR U17290 ( .A(n16225), .B(n16224), .Z(n16226) );
  AND U17291 ( .A(n16227), .B(n16226), .Z(n16245) );
  XOR U17292 ( .A(a[666]), .B(n2271), .Z(n16249) );
  AND U17293 ( .A(a[664]), .B(b[3]), .Z(n16253) );
  AND U17294 ( .A(a[668]), .B(b[0]), .Z(n16229) );
  XNOR U17295 ( .A(n16229), .B(n2175), .Z(n16231) );
  NANDN U17296 ( .A(b[0]), .B(a[667]), .Z(n16230) );
  NAND U17297 ( .A(n16231), .B(n16230), .Z(n16254) );
  XOR U17298 ( .A(n16253), .B(n16254), .Z(n16256) );
  XOR U17299 ( .A(n16255), .B(n16256), .Z(n16244) );
  NANDN U17300 ( .A(n16233), .B(n16232), .Z(n16237) );
  OR U17301 ( .A(n16235), .B(n16234), .Z(n16236) );
  AND U17302 ( .A(n16237), .B(n16236), .Z(n16243) );
  XOR U17303 ( .A(n16244), .B(n16243), .Z(n16246) );
  XOR U17304 ( .A(n16245), .B(n16246), .Z(n16259) );
  XNOR U17305 ( .A(n16259), .B(sreg[1688]), .Z(n16261) );
  NANDN U17306 ( .A(n16238), .B(sreg[1687]), .Z(n16242) );
  NAND U17307 ( .A(n16240), .B(n16239), .Z(n16241) );
  NAND U17308 ( .A(n16242), .B(n16241), .Z(n16260) );
  XOR U17309 ( .A(n16261), .B(n16260), .Z(c[1688]) );
  NANDN U17310 ( .A(n16244), .B(n16243), .Z(n16248) );
  OR U17311 ( .A(n16246), .B(n16245), .Z(n16247) );
  AND U17312 ( .A(n16248), .B(n16247), .Z(n16266) );
  XOR U17313 ( .A(a[667]), .B(n2271), .Z(n16270) );
  AND U17314 ( .A(a[669]), .B(b[0]), .Z(n16250) );
  XNOR U17315 ( .A(n16250), .B(n2175), .Z(n16252) );
  NANDN U17316 ( .A(b[0]), .B(a[668]), .Z(n16251) );
  NAND U17317 ( .A(n16252), .B(n16251), .Z(n16275) );
  AND U17318 ( .A(a[665]), .B(b[3]), .Z(n16274) );
  XOR U17319 ( .A(n16275), .B(n16274), .Z(n16277) );
  XOR U17320 ( .A(n16276), .B(n16277), .Z(n16265) );
  NANDN U17321 ( .A(n16254), .B(n16253), .Z(n16258) );
  OR U17322 ( .A(n16256), .B(n16255), .Z(n16257) );
  AND U17323 ( .A(n16258), .B(n16257), .Z(n16264) );
  XOR U17324 ( .A(n16265), .B(n16264), .Z(n16267) );
  XOR U17325 ( .A(n16266), .B(n16267), .Z(n16280) );
  XNOR U17326 ( .A(n16280), .B(sreg[1689]), .Z(n16282) );
  NANDN U17327 ( .A(n16259), .B(sreg[1688]), .Z(n16263) );
  NAND U17328 ( .A(n16261), .B(n16260), .Z(n16262) );
  NAND U17329 ( .A(n16263), .B(n16262), .Z(n16281) );
  XOR U17330 ( .A(n16282), .B(n16281), .Z(c[1689]) );
  NANDN U17331 ( .A(n16265), .B(n16264), .Z(n16269) );
  OR U17332 ( .A(n16267), .B(n16266), .Z(n16268) );
  AND U17333 ( .A(n16269), .B(n16268), .Z(n16287) );
  XOR U17334 ( .A(a[668]), .B(n2271), .Z(n16291) );
  AND U17335 ( .A(a[670]), .B(b[0]), .Z(n16271) );
  XNOR U17336 ( .A(n16271), .B(n2175), .Z(n16273) );
  NANDN U17337 ( .A(b[0]), .B(a[669]), .Z(n16272) );
  NAND U17338 ( .A(n16273), .B(n16272), .Z(n16296) );
  AND U17339 ( .A(a[666]), .B(b[3]), .Z(n16295) );
  XOR U17340 ( .A(n16296), .B(n16295), .Z(n16298) );
  XOR U17341 ( .A(n16297), .B(n16298), .Z(n16286) );
  NANDN U17342 ( .A(n16275), .B(n16274), .Z(n16279) );
  OR U17343 ( .A(n16277), .B(n16276), .Z(n16278) );
  AND U17344 ( .A(n16279), .B(n16278), .Z(n16285) );
  XOR U17345 ( .A(n16286), .B(n16285), .Z(n16288) );
  XOR U17346 ( .A(n16287), .B(n16288), .Z(n16301) );
  XNOR U17347 ( .A(n16301), .B(sreg[1690]), .Z(n16303) );
  NANDN U17348 ( .A(n16280), .B(sreg[1689]), .Z(n16284) );
  NAND U17349 ( .A(n16282), .B(n16281), .Z(n16283) );
  NAND U17350 ( .A(n16284), .B(n16283), .Z(n16302) );
  XOR U17351 ( .A(n16303), .B(n16302), .Z(c[1690]) );
  NANDN U17352 ( .A(n16286), .B(n16285), .Z(n16290) );
  OR U17353 ( .A(n16288), .B(n16287), .Z(n16289) );
  AND U17354 ( .A(n16290), .B(n16289), .Z(n16308) );
  XOR U17355 ( .A(a[669]), .B(n2271), .Z(n16312) );
  AND U17356 ( .A(a[671]), .B(b[0]), .Z(n16292) );
  XNOR U17357 ( .A(n16292), .B(n2175), .Z(n16294) );
  NANDN U17358 ( .A(b[0]), .B(a[670]), .Z(n16293) );
  NAND U17359 ( .A(n16294), .B(n16293), .Z(n16317) );
  AND U17360 ( .A(a[667]), .B(b[3]), .Z(n16316) );
  XOR U17361 ( .A(n16317), .B(n16316), .Z(n16319) );
  XOR U17362 ( .A(n16318), .B(n16319), .Z(n16307) );
  NANDN U17363 ( .A(n16296), .B(n16295), .Z(n16300) );
  OR U17364 ( .A(n16298), .B(n16297), .Z(n16299) );
  AND U17365 ( .A(n16300), .B(n16299), .Z(n16306) );
  XOR U17366 ( .A(n16307), .B(n16306), .Z(n16309) );
  XOR U17367 ( .A(n16308), .B(n16309), .Z(n16322) );
  XNOR U17368 ( .A(n16322), .B(sreg[1691]), .Z(n16324) );
  NANDN U17369 ( .A(n16301), .B(sreg[1690]), .Z(n16305) );
  NAND U17370 ( .A(n16303), .B(n16302), .Z(n16304) );
  NAND U17371 ( .A(n16305), .B(n16304), .Z(n16323) );
  XOR U17372 ( .A(n16324), .B(n16323), .Z(c[1691]) );
  NANDN U17373 ( .A(n16307), .B(n16306), .Z(n16311) );
  OR U17374 ( .A(n16309), .B(n16308), .Z(n16310) );
  AND U17375 ( .A(n16311), .B(n16310), .Z(n16329) );
  XOR U17376 ( .A(a[670]), .B(n2271), .Z(n16333) );
  AND U17377 ( .A(a[672]), .B(b[0]), .Z(n16313) );
  XNOR U17378 ( .A(n16313), .B(n2175), .Z(n16315) );
  NANDN U17379 ( .A(b[0]), .B(a[671]), .Z(n16314) );
  NAND U17380 ( .A(n16315), .B(n16314), .Z(n16338) );
  AND U17381 ( .A(a[668]), .B(b[3]), .Z(n16337) );
  XOR U17382 ( .A(n16338), .B(n16337), .Z(n16340) );
  XOR U17383 ( .A(n16339), .B(n16340), .Z(n16328) );
  NANDN U17384 ( .A(n16317), .B(n16316), .Z(n16321) );
  OR U17385 ( .A(n16319), .B(n16318), .Z(n16320) );
  AND U17386 ( .A(n16321), .B(n16320), .Z(n16327) );
  XOR U17387 ( .A(n16328), .B(n16327), .Z(n16330) );
  XOR U17388 ( .A(n16329), .B(n16330), .Z(n16343) );
  XNOR U17389 ( .A(n16343), .B(sreg[1692]), .Z(n16345) );
  NANDN U17390 ( .A(n16322), .B(sreg[1691]), .Z(n16326) );
  NAND U17391 ( .A(n16324), .B(n16323), .Z(n16325) );
  NAND U17392 ( .A(n16326), .B(n16325), .Z(n16344) );
  XOR U17393 ( .A(n16345), .B(n16344), .Z(c[1692]) );
  NANDN U17394 ( .A(n16328), .B(n16327), .Z(n16332) );
  OR U17395 ( .A(n16330), .B(n16329), .Z(n16331) );
  AND U17396 ( .A(n16332), .B(n16331), .Z(n16350) );
  XOR U17397 ( .A(a[671]), .B(n2272), .Z(n16354) );
  AND U17398 ( .A(a[673]), .B(b[0]), .Z(n16334) );
  XNOR U17399 ( .A(n16334), .B(n2175), .Z(n16336) );
  NANDN U17400 ( .A(b[0]), .B(a[672]), .Z(n16335) );
  NAND U17401 ( .A(n16336), .B(n16335), .Z(n16359) );
  AND U17402 ( .A(a[669]), .B(b[3]), .Z(n16358) );
  XOR U17403 ( .A(n16359), .B(n16358), .Z(n16361) );
  XOR U17404 ( .A(n16360), .B(n16361), .Z(n16349) );
  NANDN U17405 ( .A(n16338), .B(n16337), .Z(n16342) );
  OR U17406 ( .A(n16340), .B(n16339), .Z(n16341) );
  AND U17407 ( .A(n16342), .B(n16341), .Z(n16348) );
  XOR U17408 ( .A(n16349), .B(n16348), .Z(n16351) );
  XOR U17409 ( .A(n16350), .B(n16351), .Z(n16364) );
  XNOR U17410 ( .A(n16364), .B(sreg[1693]), .Z(n16366) );
  NANDN U17411 ( .A(n16343), .B(sreg[1692]), .Z(n16347) );
  NAND U17412 ( .A(n16345), .B(n16344), .Z(n16346) );
  NAND U17413 ( .A(n16347), .B(n16346), .Z(n16365) );
  XOR U17414 ( .A(n16366), .B(n16365), .Z(c[1693]) );
  NANDN U17415 ( .A(n16349), .B(n16348), .Z(n16353) );
  OR U17416 ( .A(n16351), .B(n16350), .Z(n16352) );
  AND U17417 ( .A(n16353), .B(n16352), .Z(n16371) );
  XOR U17418 ( .A(a[672]), .B(n2272), .Z(n16375) );
  AND U17419 ( .A(a[670]), .B(b[3]), .Z(n16379) );
  AND U17420 ( .A(a[674]), .B(b[0]), .Z(n16355) );
  XNOR U17421 ( .A(n16355), .B(n2175), .Z(n16357) );
  NANDN U17422 ( .A(b[0]), .B(a[673]), .Z(n16356) );
  NAND U17423 ( .A(n16357), .B(n16356), .Z(n16380) );
  XOR U17424 ( .A(n16379), .B(n16380), .Z(n16382) );
  XOR U17425 ( .A(n16381), .B(n16382), .Z(n16370) );
  NANDN U17426 ( .A(n16359), .B(n16358), .Z(n16363) );
  OR U17427 ( .A(n16361), .B(n16360), .Z(n16362) );
  AND U17428 ( .A(n16363), .B(n16362), .Z(n16369) );
  XOR U17429 ( .A(n16370), .B(n16369), .Z(n16372) );
  XOR U17430 ( .A(n16371), .B(n16372), .Z(n16385) );
  XNOR U17431 ( .A(n16385), .B(sreg[1694]), .Z(n16387) );
  NANDN U17432 ( .A(n16364), .B(sreg[1693]), .Z(n16368) );
  NAND U17433 ( .A(n16366), .B(n16365), .Z(n16367) );
  NAND U17434 ( .A(n16368), .B(n16367), .Z(n16386) );
  XOR U17435 ( .A(n16387), .B(n16386), .Z(c[1694]) );
  NANDN U17436 ( .A(n16370), .B(n16369), .Z(n16374) );
  OR U17437 ( .A(n16372), .B(n16371), .Z(n16373) );
  AND U17438 ( .A(n16374), .B(n16373), .Z(n16392) );
  XOR U17439 ( .A(a[673]), .B(n2272), .Z(n16396) );
  AND U17440 ( .A(a[675]), .B(b[0]), .Z(n16376) );
  XNOR U17441 ( .A(n16376), .B(n2175), .Z(n16378) );
  NANDN U17442 ( .A(b[0]), .B(a[674]), .Z(n16377) );
  NAND U17443 ( .A(n16378), .B(n16377), .Z(n16401) );
  AND U17444 ( .A(a[671]), .B(b[3]), .Z(n16400) );
  XOR U17445 ( .A(n16401), .B(n16400), .Z(n16403) );
  XOR U17446 ( .A(n16402), .B(n16403), .Z(n16391) );
  NANDN U17447 ( .A(n16380), .B(n16379), .Z(n16384) );
  OR U17448 ( .A(n16382), .B(n16381), .Z(n16383) );
  AND U17449 ( .A(n16384), .B(n16383), .Z(n16390) );
  XOR U17450 ( .A(n16391), .B(n16390), .Z(n16393) );
  XOR U17451 ( .A(n16392), .B(n16393), .Z(n16406) );
  XNOR U17452 ( .A(n16406), .B(sreg[1695]), .Z(n16408) );
  NANDN U17453 ( .A(n16385), .B(sreg[1694]), .Z(n16389) );
  NAND U17454 ( .A(n16387), .B(n16386), .Z(n16388) );
  NAND U17455 ( .A(n16389), .B(n16388), .Z(n16407) );
  XOR U17456 ( .A(n16408), .B(n16407), .Z(c[1695]) );
  NANDN U17457 ( .A(n16391), .B(n16390), .Z(n16395) );
  OR U17458 ( .A(n16393), .B(n16392), .Z(n16394) );
  AND U17459 ( .A(n16395), .B(n16394), .Z(n16413) );
  XOR U17460 ( .A(a[674]), .B(n2272), .Z(n16417) );
  AND U17461 ( .A(a[672]), .B(b[3]), .Z(n16421) );
  AND U17462 ( .A(a[676]), .B(b[0]), .Z(n16397) );
  XNOR U17463 ( .A(n16397), .B(n2175), .Z(n16399) );
  NANDN U17464 ( .A(b[0]), .B(a[675]), .Z(n16398) );
  NAND U17465 ( .A(n16399), .B(n16398), .Z(n16422) );
  XOR U17466 ( .A(n16421), .B(n16422), .Z(n16424) );
  XOR U17467 ( .A(n16423), .B(n16424), .Z(n16412) );
  NANDN U17468 ( .A(n16401), .B(n16400), .Z(n16405) );
  OR U17469 ( .A(n16403), .B(n16402), .Z(n16404) );
  AND U17470 ( .A(n16405), .B(n16404), .Z(n16411) );
  XOR U17471 ( .A(n16412), .B(n16411), .Z(n16414) );
  XOR U17472 ( .A(n16413), .B(n16414), .Z(n16427) );
  XNOR U17473 ( .A(n16427), .B(sreg[1696]), .Z(n16429) );
  NANDN U17474 ( .A(n16406), .B(sreg[1695]), .Z(n16410) );
  NAND U17475 ( .A(n16408), .B(n16407), .Z(n16409) );
  NAND U17476 ( .A(n16410), .B(n16409), .Z(n16428) );
  XOR U17477 ( .A(n16429), .B(n16428), .Z(c[1696]) );
  NANDN U17478 ( .A(n16412), .B(n16411), .Z(n16416) );
  OR U17479 ( .A(n16414), .B(n16413), .Z(n16415) );
  AND U17480 ( .A(n16416), .B(n16415), .Z(n16434) );
  XOR U17481 ( .A(a[675]), .B(n2272), .Z(n16438) );
  AND U17482 ( .A(a[673]), .B(b[3]), .Z(n16442) );
  AND U17483 ( .A(a[677]), .B(b[0]), .Z(n16418) );
  XNOR U17484 ( .A(n16418), .B(n2175), .Z(n16420) );
  NANDN U17485 ( .A(b[0]), .B(a[676]), .Z(n16419) );
  NAND U17486 ( .A(n16420), .B(n16419), .Z(n16443) );
  XOR U17487 ( .A(n16442), .B(n16443), .Z(n16445) );
  XOR U17488 ( .A(n16444), .B(n16445), .Z(n16433) );
  NANDN U17489 ( .A(n16422), .B(n16421), .Z(n16426) );
  OR U17490 ( .A(n16424), .B(n16423), .Z(n16425) );
  AND U17491 ( .A(n16426), .B(n16425), .Z(n16432) );
  XOR U17492 ( .A(n16433), .B(n16432), .Z(n16435) );
  XOR U17493 ( .A(n16434), .B(n16435), .Z(n16448) );
  XNOR U17494 ( .A(n16448), .B(sreg[1697]), .Z(n16450) );
  NANDN U17495 ( .A(n16427), .B(sreg[1696]), .Z(n16431) );
  NAND U17496 ( .A(n16429), .B(n16428), .Z(n16430) );
  NAND U17497 ( .A(n16431), .B(n16430), .Z(n16449) );
  XOR U17498 ( .A(n16450), .B(n16449), .Z(c[1697]) );
  NANDN U17499 ( .A(n16433), .B(n16432), .Z(n16437) );
  OR U17500 ( .A(n16435), .B(n16434), .Z(n16436) );
  AND U17501 ( .A(n16437), .B(n16436), .Z(n16455) );
  XOR U17502 ( .A(a[676]), .B(n2272), .Z(n16459) );
  AND U17503 ( .A(a[678]), .B(b[0]), .Z(n16439) );
  XNOR U17504 ( .A(n16439), .B(n2175), .Z(n16441) );
  NANDN U17505 ( .A(b[0]), .B(a[677]), .Z(n16440) );
  NAND U17506 ( .A(n16441), .B(n16440), .Z(n16464) );
  AND U17507 ( .A(a[674]), .B(b[3]), .Z(n16463) );
  XOR U17508 ( .A(n16464), .B(n16463), .Z(n16466) );
  XOR U17509 ( .A(n16465), .B(n16466), .Z(n16454) );
  NANDN U17510 ( .A(n16443), .B(n16442), .Z(n16447) );
  OR U17511 ( .A(n16445), .B(n16444), .Z(n16446) );
  AND U17512 ( .A(n16447), .B(n16446), .Z(n16453) );
  XOR U17513 ( .A(n16454), .B(n16453), .Z(n16456) );
  XOR U17514 ( .A(n16455), .B(n16456), .Z(n16469) );
  XNOR U17515 ( .A(n16469), .B(sreg[1698]), .Z(n16471) );
  NANDN U17516 ( .A(n16448), .B(sreg[1697]), .Z(n16452) );
  NAND U17517 ( .A(n16450), .B(n16449), .Z(n16451) );
  NAND U17518 ( .A(n16452), .B(n16451), .Z(n16470) );
  XOR U17519 ( .A(n16471), .B(n16470), .Z(c[1698]) );
  NANDN U17520 ( .A(n16454), .B(n16453), .Z(n16458) );
  OR U17521 ( .A(n16456), .B(n16455), .Z(n16457) );
  AND U17522 ( .A(n16458), .B(n16457), .Z(n16476) );
  XOR U17523 ( .A(a[677]), .B(n2272), .Z(n16480) );
  AND U17524 ( .A(a[675]), .B(b[3]), .Z(n16484) );
  AND U17525 ( .A(a[679]), .B(b[0]), .Z(n16460) );
  XNOR U17526 ( .A(n16460), .B(n2175), .Z(n16462) );
  NANDN U17527 ( .A(b[0]), .B(a[678]), .Z(n16461) );
  NAND U17528 ( .A(n16462), .B(n16461), .Z(n16485) );
  XOR U17529 ( .A(n16484), .B(n16485), .Z(n16487) );
  XOR U17530 ( .A(n16486), .B(n16487), .Z(n16475) );
  NANDN U17531 ( .A(n16464), .B(n16463), .Z(n16468) );
  OR U17532 ( .A(n16466), .B(n16465), .Z(n16467) );
  AND U17533 ( .A(n16468), .B(n16467), .Z(n16474) );
  XOR U17534 ( .A(n16475), .B(n16474), .Z(n16477) );
  XOR U17535 ( .A(n16476), .B(n16477), .Z(n16490) );
  XNOR U17536 ( .A(n16490), .B(sreg[1699]), .Z(n16492) );
  NANDN U17537 ( .A(n16469), .B(sreg[1698]), .Z(n16473) );
  NAND U17538 ( .A(n16471), .B(n16470), .Z(n16472) );
  NAND U17539 ( .A(n16473), .B(n16472), .Z(n16491) );
  XOR U17540 ( .A(n16492), .B(n16491), .Z(c[1699]) );
  NANDN U17541 ( .A(n16475), .B(n16474), .Z(n16479) );
  OR U17542 ( .A(n16477), .B(n16476), .Z(n16478) );
  AND U17543 ( .A(n16479), .B(n16478), .Z(n16497) );
  XOR U17544 ( .A(a[678]), .B(n2273), .Z(n16501) );
  AND U17545 ( .A(a[680]), .B(b[0]), .Z(n16481) );
  XNOR U17546 ( .A(n16481), .B(n2175), .Z(n16483) );
  NANDN U17547 ( .A(b[0]), .B(a[679]), .Z(n16482) );
  NAND U17548 ( .A(n16483), .B(n16482), .Z(n16506) );
  AND U17549 ( .A(a[676]), .B(b[3]), .Z(n16505) );
  XOR U17550 ( .A(n16506), .B(n16505), .Z(n16508) );
  XOR U17551 ( .A(n16507), .B(n16508), .Z(n16496) );
  NANDN U17552 ( .A(n16485), .B(n16484), .Z(n16489) );
  OR U17553 ( .A(n16487), .B(n16486), .Z(n16488) );
  AND U17554 ( .A(n16489), .B(n16488), .Z(n16495) );
  XOR U17555 ( .A(n16496), .B(n16495), .Z(n16498) );
  XOR U17556 ( .A(n16497), .B(n16498), .Z(n16511) );
  XNOR U17557 ( .A(n16511), .B(sreg[1700]), .Z(n16513) );
  NANDN U17558 ( .A(n16490), .B(sreg[1699]), .Z(n16494) );
  NAND U17559 ( .A(n16492), .B(n16491), .Z(n16493) );
  NAND U17560 ( .A(n16494), .B(n16493), .Z(n16512) );
  XOR U17561 ( .A(n16513), .B(n16512), .Z(c[1700]) );
  NANDN U17562 ( .A(n16496), .B(n16495), .Z(n16500) );
  OR U17563 ( .A(n16498), .B(n16497), .Z(n16499) );
  AND U17564 ( .A(n16500), .B(n16499), .Z(n16518) );
  XOR U17565 ( .A(a[679]), .B(n2273), .Z(n16522) );
  AND U17566 ( .A(a[677]), .B(b[3]), .Z(n16526) );
  AND U17567 ( .A(a[681]), .B(b[0]), .Z(n16502) );
  XNOR U17568 ( .A(n16502), .B(n2175), .Z(n16504) );
  NANDN U17569 ( .A(b[0]), .B(a[680]), .Z(n16503) );
  NAND U17570 ( .A(n16504), .B(n16503), .Z(n16527) );
  XOR U17571 ( .A(n16526), .B(n16527), .Z(n16529) );
  XOR U17572 ( .A(n16528), .B(n16529), .Z(n16517) );
  NANDN U17573 ( .A(n16506), .B(n16505), .Z(n16510) );
  OR U17574 ( .A(n16508), .B(n16507), .Z(n16509) );
  AND U17575 ( .A(n16510), .B(n16509), .Z(n16516) );
  XOR U17576 ( .A(n16517), .B(n16516), .Z(n16519) );
  XOR U17577 ( .A(n16518), .B(n16519), .Z(n16532) );
  XNOR U17578 ( .A(n16532), .B(sreg[1701]), .Z(n16534) );
  NANDN U17579 ( .A(n16511), .B(sreg[1700]), .Z(n16515) );
  NAND U17580 ( .A(n16513), .B(n16512), .Z(n16514) );
  NAND U17581 ( .A(n16515), .B(n16514), .Z(n16533) );
  XOR U17582 ( .A(n16534), .B(n16533), .Z(c[1701]) );
  NANDN U17583 ( .A(n16517), .B(n16516), .Z(n16521) );
  OR U17584 ( .A(n16519), .B(n16518), .Z(n16520) );
  AND U17585 ( .A(n16521), .B(n16520), .Z(n16539) );
  XOR U17586 ( .A(a[680]), .B(n2273), .Z(n16543) );
  AND U17587 ( .A(a[682]), .B(b[0]), .Z(n16523) );
  XNOR U17588 ( .A(n16523), .B(n2175), .Z(n16525) );
  NANDN U17589 ( .A(b[0]), .B(a[681]), .Z(n16524) );
  NAND U17590 ( .A(n16525), .B(n16524), .Z(n16548) );
  AND U17591 ( .A(a[678]), .B(b[3]), .Z(n16547) );
  XOR U17592 ( .A(n16548), .B(n16547), .Z(n16550) );
  XOR U17593 ( .A(n16549), .B(n16550), .Z(n16538) );
  NANDN U17594 ( .A(n16527), .B(n16526), .Z(n16531) );
  OR U17595 ( .A(n16529), .B(n16528), .Z(n16530) );
  AND U17596 ( .A(n16531), .B(n16530), .Z(n16537) );
  XOR U17597 ( .A(n16538), .B(n16537), .Z(n16540) );
  XOR U17598 ( .A(n16539), .B(n16540), .Z(n16553) );
  XNOR U17599 ( .A(n16553), .B(sreg[1702]), .Z(n16555) );
  NANDN U17600 ( .A(n16532), .B(sreg[1701]), .Z(n16536) );
  NAND U17601 ( .A(n16534), .B(n16533), .Z(n16535) );
  NAND U17602 ( .A(n16536), .B(n16535), .Z(n16554) );
  XOR U17603 ( .A(n16555), .B(n16554), .Z(c[1702]) );
  NANDN U17604 ( .A(n16538), .B(n16537), .Z(n16542) );
  OR U17605 ( .A(n16540), .B(n16539), .Z(n16541) );
  AND U17606 ( .A(n16542), .B(n16541), .Z(n16560) );
  XOR U17607 ( .A(a[681]), .B(n2273), .Z(n16564) );
  AND U17608 ( .A(a[679]), .B(b[3]), .Z(n16568) );
  AND U17609 ( .A(a[683]), .B(b[0]), .Z(n16544) );
  XNOR U17610 ( .A(n16544), .B(n2175), .Z(n16546) );
  NANDN U17611 ( .A(b[0]), .B(a[682]), .Z(n16545) );
  NAND U17612 ( .A(n16546), .B(n16545), .Z(n16569) );
  XOR U17613 ( .A(n16568), .B(n16569), .Z(n16571) );
  XOR U17614 ( .A(n16570), .B(n16571), .Z(n16559) );
  NANDN U17615 ( .A(n16548), .B(n16547), .Z(n16552) );
  OR U17616 ( .A(n16550), .B(n16549), .Z(n16551) );
  AND U17617 ( .A(n16552), .B(n16551), .Z(n16558) );
  XOR U17618 ( .A(n16559), .B(n16558), .Z(n16561) );
  XOR U17619 ( .A(n16560), .B(n16561), .Z(n16574) );
  XNOR U17620 ( .A(n16574), .B(sreg[1703]), .Z(n16576) );
  NANDN U17621 ( .A(n16553), .B(sreg[1702]), .Z(n16557) );
  NAND U17622 ( .A(n16555), .B(n16554), .Z(n16556) );
  NAND U17623 ( .A(n16557), .B(n16556), .Z(n16575) );
  XOR U17624 ( .A(n16576), .B(n16575), .Z(c[1703]) );
  NANDN U17625 ( .A(n16559), .B(n16558), .Z(n16563) );
  OR U17626 ( .A(n16561), .B(n16560), .Z(n16562) );
  AND U17627 ( .A(n16563), .B(n16562), .Z(n16581) );
  XOR U17628 ( .A(a[682]), .B(n2273), .Z(n16585) );
  AND U17629 ( .A(a[684]), .B(b[0]), .Z(n16565) );
  XNOR U17630 ( .A(n16565), .B(n2175), .Z(n16567) );
  NANDN U17631 ( .A(b[0]), .B(a[683]), .Z(n16566) );
  NAND U17632 ( .A(n16567), .B(n16566), .Z(n16590) );
  AND U17633 ( .A(a[680]), .B(b[3]), .Z(n16589) );
  XOR U17634 ( .A(n16590), .B(n16589), .Z(n16592) );
  XOR U17635 ( .A(n16591), .B(n16592), .Z(n16580) );
  NANDN U17636 ( .A(n16569), .B(n16568), .Z(n16573) );
  OR U17637 ( .A(n16571), .B(n16570), .Z(n16572) );
  AND U17638 ( .A(n16573), .B(n16572), .Z(n16579) );
  XOR U17639 ( .A(n16580), .B(n16579), .Z(n16582) );
  XOR U17640 ( .A(n16581), .B(n16582), .Z(n16595) );
  XNOR U17641 ( .A(n16595), .B(sreg[1704]), .Z(n16597) );
  NANDN U17642 ( .A(n16574), .B(sreg[1703]), .Z(n16578) );
  NAND U17643 ( .A(n16576), .B(n16575), .Z(n16577) );
  NAND U17644 ( .A(n16578), .B(n16577), .Z(n16596) );
  XOR U17645 ( .A(n16597), .B(n16596), .Z(c[1704]) );
  NANDN U17646 ( .A(n16580), .B(n16579), .Z(n16584) );
  OR U17647 ( .A(n16582), .B(n16581), .Z(n16583) );
  AND U17648 ( .A(n16584), .B(n16583), .Z(n16602) );
  XOR U17649 ( .A(a[683]), .B(n2273), .Z(n16606) );
  AND U17650 ( .A(a[685]), .B(b[0]), .Z(n16586) );
  XNOR U17651 ( .A(n16586), .B(n2175), .Z(n16588) );
  NANDN U17652 ( .A(b[0]), .B(a[684]), .Z(n16587) );
  NAND U17653 ( .A(n16588), .B(n16587), .Z(n16611) );
  AND U17654 ( .A(a[681]), .B(b[3]), .Z(n16610) );
  XOR U17655 ( .A(n16611), .B(n16610), .Z(n16613) );
  XOR U17656 ( .A(n16612), .B(n16613), .Z(n16601) );
  NANDN U17657 ( .A(n16590), .B(n16589), .Z(n16594) );
  OR U17658 ( .A(n16592), .B(n16591), .Z(n16593) );
  AND U17659 ( .A(n16594), .B(n16593), .Z(n16600) );
  XOR U17660 ( .A(n16601), .B(n16600), .Z(n16603) );
  XOR U17661 ( .A(n16602), .B(n16603), .Z(n16616) );
  XNOR U17662 ( .A(n16616), .B(sreg[1705]), .Z(n16618) );
  NANDN U17663 ( .A(n16595), .B(sreg[1704]), .Z(n16599) );
  NAND U17664 ( .A(n16597), .B(n16596), .Z(n16598) );
  NAND U17665 ( .A(n16599), .B(n16598), .Z(n16617) );
  XOR U17666 ( .A(n16618), .B(n16617), .Z(c[1705]) );
  NANDN U17667 ( .A(n16601), .B(n16600), .Z(n16605) );
  OR U17668 ( .A(n16603), .B(n16602), .Z(n16604) );
  AND U17669 ( .A(n16605), .B(n16604), .Z(n16623) );
  XOR U17670 ( .A(a[684]), .B(n2273), .Z(n16627) );
  AND U17671 ( .A(a[682]), .B(b[3]), .Z(n16631) );
  AND U17672 ( .A(a[686]), .B(b[0]), .Z(n16607) );
  XNOR U17673 ( .A(n16607), .B(n2175), .Z(n16609) );
  NANDN U17674 ( .A(b[0]), .B(a[685]), .Z(n16608) );
  NAND U17675 ( .A(n16609), .B(n16608), .Z(n16632) );
  XOR U17676 ( .A(n16631), .B(n16632), .Z(n16634) );
  XOR U17677 ( .A(n16633), .B(n16634), .Z(n16622) );
  NANDN U17678 ( .A(n16611), .B(n16610), .Z(n16615) );
  OR U17679 ( .A(n16613), .B(n16612), .Z(n16614) );
  AND U17680 ( .A(n16615), .B(n16614), .Z(n16621) );
  XOR U17681 ( .A(n16622), .B(n16621), .Z(n16624) );
  XOR U17682 ( .A(n16623), .B(n16624), .Z(n16637) );
  XNOR U17683 ( .A(n16637), .B(sreg[1706]), .Z(n16639) );
  NANDN U17684 ( .A(n16616), .B(sreg[1705]), .Z(n16620) );
  NAND U17685 ( .A(n16618), .B(n16617), .Z(n16619) );
  NAND U17686 ( .A(n16620), .B(n16619), .Z(n16638) );
  XOR U17687 ( .A(n16639), .B(n16638), .Z(c[1706]) );
  NANDN U17688 ( .A(n16622), .B(n16621), .Z(n16626) );
  OR U17689 ( .A(n16624), .B(n16623), .Z(n16625) );
  AND U17690 ( .A(n16626), .B(n16625), .Z(n16644) );
  XOR U17691 ( .A(a[685]), .B(n2274), .Z(n16648) );
  AND U17692 ( .A(a[687]), .B(b[0]), .Z(n16628) );
  XNOR U17693 ( .A(n16628), .B(n2175), .Z(n16630) );
  NANDN U17694 ( .A(b[0]), .B(a[686]), .Z(n16629) );
  NAND U17695 ( .A(n16630), .B(n16629), .Z(n16653) );
  AND U17696 ( .A(a[683]), .B(b[3]), .Z(n16652) );
  XOR U17697 ( .A(n16653), .B(n16652), .Z(n16655) );
  XOR U17698 ( .A(n16654), .B(n16655), .Z(n16643) );
  NANDN U17699 ( .A(n16632), .B(n16631), .Z(n16636) );
  OR U17700 ( .A(n16634), .B(n16633), .Z(n16635) );
  AND U17701 ( .A(n16636), .B(n16635), .Z(n16642) );
  XOR U17702 ( .A(n16643), .B(n16642), .Z(n16645) );
  XOR U17703 ( .A(n16644), .B(n16645), .Z(n16658) );
  XNOR U17704 ( .A(n16658), .B(sreg[1707]), .Z(n16660) );
  NANDN U17705 ( .A(n16637), .B(sreg[1706]), .Z(n16641) );
  NAND U17706 ( .A(n16639), .B(n16638), .Z(n16640) );
  NAND U17707 ( .A(n16641), .B(n16640), .Z(n16659) );
  XOR U17708 ( .A(n16660), .B(n16659), .Z(c[1707]) );
  NANDN U17709 ( .A(n16643), .B(n16642), .Z(n16647) );
  OR U17710 ( .A(n16645), .B(n16644), .Z(n16646) );
  AND U17711 ( .A(n16647), .B(n16646), .Z(n16665) );
  XOR U17712 ( .A(a[686]), .B(n2274), .Z(n16669) );
  AND U17713 ( .A(a[688]), .B(b[0]), .Z(n16649) );
  XNOR U17714 ( .A(n16649), .B(n2175), .Z(n16651) );
  NANDN U17715 ( .A(b[0]), .B(a[687]), .Z(n16650) );
  NAND U17716 ( .A(n16651), .B(n16650), .Z(n16674) );
  AND U17717 ( .A(a[684]), .B(b[3]), .Z(n16673) );
  XOR U17718 ( .A(n16674), .B(n16673), .Z(n16676) );
  XOR U17719 ( .A(n16675), .B(n16676), .Z(n16664) );
  NANDN U17720 ( .A(n16653), .B(n16652), .Z(n16657) );
  OR U17721 ( .A(n16655), .B(n16654), .Z(n16656) );
  AND U17722 ( .A(n16657), .B(n16656), .Z(n16663) );
  XOR U17723 ( .A(n16664), .B(n16663), .Z(n16666) );
  XOR U17724 ( .A(n16665), .B(n16666), .Z(n16679) );
  XNOR U17725 ( .A(n16679), .B(sreg[1708]), .Z(n16681) );
  NANDN U17726 ( .A(n16658), .B(sreg[1707]), .Z(n16662) );
  NAND U17727 ( .A(n16660), .B(n16659), .Z(n16661) );
  NAND U17728 ( .A(n16662), .B(n16661), .Z(n16680) );
  XOR U17729 ( .A(n16681), .B(n16680), .Z(c[1708]) );
  NANDN U17730 ( .A(n16664), .B(n16663), .Z(n16668) );
  OR U17731 ( .A(n16666), .B(n16665), .Z(n16667) );
  AND U17732 ( .A(n16668), .B(n16667), .Z(n16686) );
  XOR U17733 ( .A(a[687]), .B(n2274), .Z(n16690) );
  AND U17734 ( .A(a[689]), .B(b[0]), .Z(n16670) );
  XNOR U17735 ( .A(n16670), .B(n2175), .Z(n16672) );
  NANDN U17736 ( .A(b[0]), .B(a[688]), .Z(n16671) );
  NAND U17737 ( .A(n16672), .B(n16671), .Z(n16695) );
  AND U17738 ( .A(a[685]), .B(b[3]), .Z(n16694) );
  XOR U17739 ( .A(n16695), .B(n16694), .Z(n16697) );
  XOR U17740 ( .A(n16696), .B(n16697), .Z(n16685) );
  NANDN U17741 ( .A(n16674), .B(n16673), .Z(n16678) );
  OR U17742 ( .A(n16676), .B(n16675), .Z(n16677) );
  AND U17743 ( .A(n16678), .B(n16677), .Z(n16684) );
  XOR U17744 ( .A(n16685), .B(n16684), .Z(n16687) );
  XOR U17745 ( .A(n16686), .B(n16687), .Z(n16700) );
  XNOR U17746 ( .A(n16700), .B(sreg[1709]), .Z(n16702) );
  NANDN U17747 ( .A(n16679), .B(sreg[1708]), .Z(n16683) );
  NAND U17748 ( .A(n16681), .B(n16680), .Z(n16682) );
  NAND U17749 ( .A(n16683), .B(n16682), .Z(n16701) );
  XOR U17750 ( .A(n16702), .B(n16701), .Z(c[1709]) );
  NANDN U17751 ( .A(n16685), .B(n16684), .Z(n16689) );
  OR U17752 ( .A(n16687), .B(n16686), .Z(n16688) );
  AND U17753 ( .A(n16689), .B(n16688), .Z(n16707) );
  XOR U17754 ( .A(a[688]), .B(n2274), .Z(n16711) );
  AND U17755 ( .A(a[690]), .B(b[0]), .Z(n16691) );
  XNOR U17756 ( .A(n16691), .B(n2175), .Z(n16693) );
  NANDN U17757 ( .A(b[0]), .B(a[689]), .Z(n16692) );
  NAND U17758 ( .A(n16693), .B(n16692), .Z(n16716) );
  AND U17759 ( .A(a[686]), .B(b[3]), .Z(n16715) );
  XOR U17760 ( .A(n16716), .B(n16715), .Z(n16718) );
  XOR U17761 ( .A(n16717), .B(n16718), .Z(n16706) );
  NANDN U17762 ( .A(n16695), .B(n16694), .Z(n16699) );
  OR U17763 ( .A(n16697), .B(n16696), .Z(n16698) );
  AND U17764 ( .A(n16699), .B(n16698), .Z(n16705) );
  XOR U17765 ( .A(n16706), .B(n16705), .Z(n16708) );
  XOR U17766 ( .A(n16707), .B(n16708), .Z(n16721) );
  XNOR U17767 ( .A(n16721), .B(sreg[1710]), .Z(n16723) );
  NANDN U17768 ( .A(n16700), .B(sreg[1709]), .Z(n16704) );
  NAND U17769 ( .A(n16702), .B(n16701), .Z(n16703) );
  NAND U17770 ( .A(n16704), .B(n16703), .Z(n16722) );
  XOR U17771 ( .A(n16723), .B(n16722), .Z(c[1710]) );
  NANDN U17772 ( .A(n16706), .B(n16705), .Z(n16710) );
  OR U17773 ( .A(n16708), .B(n16707), .Z(n16709) );
  AND U17774 ( .A(n16710), .B(n16709), .Z(n16728) );
  XOR U17775 ( .A(a[689]), .B(n2274), .Z(n16732) );
  AND U17776 ( .A(a[687]), .B(b[3]), .Z(n16736) );
  AND U17777 ( .A(a[691]), .B(b[0]), .Z(n16712) );
  XNOR U17778 ( .A(n16712), .B(n2175), .Z(n16714) );
  NANDN U17779 ( .A(b[0]), .B(a[690]), .Z(n16713) );
  NAND U17780 ( .A(n16714), .B(n16713), .Z(n16737) );
  XOR U17781 ( .A(n16736), .B(n16737), .Z(n16739) );
  XOR U17782 ( .A(n16738), .B(n16739), .Z(n16727) );
  NANDN U17783 ( .A(n16716), .B(n16715), .Z(n16720) );
  OR U17784 ( .A(n16718), .B(n16717), .Z(n16719) );
  AND U17785 ( .A(n16720), .B(n16719), .Z(n16726) );
  XOR U17786 ( .A(n16727), .B(n16726), .Z(n16729) );
  XOR U17787 ( .A(n16728), .B(n16729), .Z(n16742) );
  XNOR U17788 ( .A(n16742), .B(sreg[1711]), .Z(n16744) );
  NANDN U17789 ( .A(n16721), .B(sreg[1710]), .Z(n16725) );
  NAND U17790 ( .A(n16723), .B(n16722), .Z(n16724) );
  NAND U17791 ( .A(n16725), .B(n16724), .Z(n16743) );
  XOR U17792 ( .A(n16744), .B(n16743), .Z(c[1711]) );
  NANDN U17793 ( .A(n16727), .B(n16726), .Z(n16731) );
  OR U17794 ( .A(n16729), .B(n16728), .Z(n16730) );
  AND U17795 ( .A(n16731), .B(n16730), .Z(n16749) );
  XOR U17796 ( .A(a[690]), .B(n2274), .Z(n16753) );
  AND U17797 ( .A(a[692]), .B(b[0]), .Z(n16733) );
  XNOR U17798 ( .A(n16733), .B(n2175), .Z(n16735) );
  NANDN U17799 ( .A(b[0]), .B(a[691]), .Z(n16734) );
  NAND U17800 ( .A(n16735), .B(n16734), .Z(n16758) );
  AND U17801 ( .A(a[688]), .B(b[3]), .Z(n16757) );
  XOR U17802 ( .A(n16758), .B(n16757), .Z(n16760) );
  XOR U17803 ( .A(n16759), .B(n16760), .Z(n16748) );
  NANDN U17804 ( .A(n16737), .B(n16736), .Z(n16741) );
  OR U17805 ( .A(n16739), .B(n16738), .Z(n16740) );
  AND U17806 ( .A(n16741), .B(n16740), .Z(n16747) );
  XOR U17807 ( .A(n16748), .B(n16747), .Z(n16750) );
  XOR U17808 ( .A(n16749), .B(n16750), .Z(n16763) );
  XNOR U17809 ( .A(n16763), .B(sreg[1712]), .Z(n16765) );
  NANDN U17810 ( .A(n16742), .B(sreg[1711]), .Z(n16746) );
  NAND U17811 ( .A(n16744), .B(n16743), .Z(n16745) );
  NAND U17812 ( .A(n16746), .B(n16745), .Z(n16764) );
  XOR U17813 ( .A(n16765), .B(n16764), .Z(c[1712]) );
  NANDN U17814 ( .A(n16748), .B(n16747), .Z(n16752) );
  OR U17815 ( .A(n16750), .B(n16749), .Z(n16751) );
  AND U17816 ( .A(n16752), .B(n16751), .Z(n16770) );
  XOR U17817 ( .A(a[691]), .B(n2274), .Z(n16774) );
  AND U17818 ( .A(a[689]), .B(b[3]), .Z(n16778) );
  AND U17819 ( .A(a[693]), .B(b[0]), .Z(n16754) );
  XNOR U17820 ( .A(n16754), .B(n2175), .Z(n16756) );
  NANDN U17821 ( .A(b[0]), .B(a[692]), .Z(n16755) );
  NAND U17822 ( .A(n16756), .B(n16755), .Z(n16779) );
  XOR U17823 ( .A(n16778), .B(n16779), .Z(n16781) );
  XOR U17824 ( .A(n16780), .B(n16781), .Z(n16769) );
  NANDN U17825 ( .A(n16758), .B(n16757), .Z(n16762) );
  OR U17826 ( .A(n16760), .B(n16759), .Z(n16761) );
  AND U17827 ( .A(n16762), .B(n16761), .Z(n16768) );
  XOR U17828 ( .A(n16769), .B(n16768), .Z(n16771) );
  XOR U17829 ( .A(n16770), .B(n16771), .Z(n16784) );
  XNOR U17830 ( .A(n16784), .B(sreg[1713]), .Z(n16786) );
  NANDN U17831 ( .A(n16763), .B(sreg[1712]), .Z(n16767) );
  NAND U17832 ( .A(n16765), .B(n16764), .Z(n16766) );
  NAND U17833 ( .A(n16767), .B(n16766), .Z(n16785) );
  XOR U17834 ( .A(n16786), .B(n16785), .Z(c[1713]) );
  NANDN U17835 ( .A(n16769), .B(n16768), .Z(n16773) );
  OR U17836 ( .A(n16771), .B(n16770), .Z(n16772) );
  AND U17837 ( .A(n16773), .B(n16772), .Z(n16791) );
  XOR U17838 ( .A(a[692]), .B(n2275), .Z(n16795) );
  AND U17839 ( .A(a[694]), .B(b[0]), .Z(n16775) );
  XNOR U17840 ( .A(n16775), .B(n2175), .Z(n16777) );
  NANDN U17841 ( .A(b[0]), .B(a[693]), .Z(n16776) );
  NAND U17842 ( .A(n16777), .B(n16776), .Z(n16800) );
  AND U17843 ( .A(a[690]), .B(b[3]), .Z(n16799) );
  XOR U17844 ( .A(n16800), .B(n16799), .Z(n16802) );
  XOR U17845 ( .A(n16801), .B(n16802), .Z(n16790) );
  NANDN U17846 ( .A(n16779), .B(n16778), .Z(n16783) );
  OR U17847 ( .A(n16781), .B(n16780), .Z(n16782) );
  AND U17848 ( .A(n16783), .B(n16782), .Z(n16789) );
  XOR U17849 ( .A(n16790), .B(n16789), .Z(n16792) );
  XOR U17850 ( .A(n16791), .B(n16792), .Z(n16805) );
  XNOR U17851 ( .A(n16805), .B(sreg[1714]), .Z(n16807) );
  NANDN U17852 ( .A(n16784), .B(sreg[1713]), .Z(n16788) );
  NAND U17853 ( .A(n16786), .B(n16785), .Z(n16787) );
  NAND U17854 ( .A(n16788), .B(n16787), .Z(n16806) );
  XOR U17855 ( .A(n16807), .B(n16806), .Z(c[1714]) );
  NANDN U17856 ( .A(n16790), .B(n16789), .Z(n16794) );
  OR U17857 ( .A(n16792), .B(n16791), .Z(n16793) );
  AND U17858 ( .A(n16794), .B(n16793), .Z(n16812) );
  XOR U17859 ( .A(a[693]), .B(n2275), .Z(n16816) );
  AND U17860 ( .A(a[695]), .B(b[0]), .Z(n16796) );
  XNOR U17861 ( .A(n16796), .B(n2175), .Z(n16798) );
  NANDN U17862 ( .A(b[0]), .B(a[694]), .Z(n16797) );
  NAND U17863 ( .A(n16798), .B(n16797), .Z(n16821) );
  AND U17864 ( .A(a[691]), .B(b[3]), .Z(n16820) );
  XOR U17865 ( .A(n16821), .B(n16820), .Z(n16823) );
  XOR U17866 ( .A(n16822), .B(n16823), .Z(n16811) );
  NANDN U17867 ( .A(n16800), .B(n16799), .Z(n16804) );
  OR U17868 ( .A(n16802), .B(n16801), .Z(n16803) );
  AND U17869 ( .A(n16804), .B(n16803), .Z(n16810) );
  XOR U17870 ( .A(n16811), .B(n16810), .Z(n16813) );
  XOR U17871 ( .A(n16812), .B(n16813), .Z(n16826) );
  XNOR U17872 ( .A(n16826), .B(sreg[1715]), .Z(n16828) );
  NANDN U17873 ( .A(n16805), .B(sreg[1714]), .Z(n16809) );
  NAND U17874 ( .A(n16807), .B(n16806), .Z(n16808) );
  NAND U17875 ( .A(n16809), .B(n16808), .Z(n16827) );
  XOR U17876 ( .A(n16828), .B(n16827), .Z(c[1715]) );
  NANDN U17877 ( .A(n16811), .B(n16810), .Z(n16815) );
  OR U17878 ( .A(n16813), .B(n16812), .Z(n16814) );
  AND U17879 ( .A(n16815), .B(n16814), .Z(n16833) );
  XOR U17880 ( .A(a[694]), .B(n2275), .Z(n16837) );
  AND U17881 ( .A(a[692]), .B(b[3]), .Z(n16841) );
  AND U17882 ( .A(a[696]), .B(b[0]), .Z(n16817) );
  XNOR U17883 ( .A(n16817), .B(n2175), .Z(n16819) );
  NANDN U17884 ( .A(b[0]), .B(a[695]), .Z(n16818) );
  NAND U17885 ( .A(n16819), .B(n16818), .Z(n16842) );
  XOR U17886 ( .A(n16841), .B(n16842), .Z(n16844) );
  XOR U17887 ( .A(n16843), .B(n16844), .Z(n16832) );
  NANDN U17888 ( .A(n16821), .B(n16820), .Z(n16825) );
  OR U17889 ( .A(n16823), .B(n16822), .Z(n16824) );
  AND U17890 ( .A(n16825), .B(n16824), .Z(n16831) );
  XOR U17891 ( .A(n16832), .B(n16831), .Z(n16834) );
  XOR U17892 ( .A(n16833), .B(n16834), .Z(n16847) );
  XNOR U17893 ( .A(n16847), .B(sreg[1716]), .Z(n16849) );
  NANDN U17894 ( .A(n16826), .B(sreg[1715]), .Z(n16830) );
  NAND U17895 ( .A(n16828), .B(n16827), .Z(n16829) );
  NAND U17896 ( .A(n16830), .B(n16829), .Z(n16848) );
  XOR U17897 ( .A(n16849), .B(n16848), .Z(c[1716]) );
  NANDN U17898 ( .A(n16832), .B(n16831), .Z(n16836) );
  OR U17899 ( .A(n16834), .B(n16833), .Z(n16835) );
  AND U17900 ( .A(n16836), .B(n16835), .Z(n16854) );
  XOR U17901 ( .A(a[695]), .B(n2275), .Z(n16858) );
  AND U17902 ( .A(a[697]), .B(b[0]), .Z(n16838) );
  XNOR U17903 ( .A(n16838), .B(n2175), .Z(n16840) );
  NANDN U17904 ( .A(b[0]), .B(a[696]), .Z(n16839) );
  NAND U17905 ( .A(n16840), .B(n16839), .Z(n16863) );
  AND U17906 ( .A(a[693]), .B(b[3]), .Z(n16862) );
  XOR U17907 ( .A(n16863), .B(n16862), .Z(n16865) );
  XOR U17908 ( .A(n16864), .B(n16865), .Z(n16853) );
  NANDN U17909 ( .A(n16842), .B(n16841), .Z(n16846) );
  OR U17910 ( .A(n16844), .B(n16843), .Z(n16845) );
  AND U17911 ( .A(n16846), .B(n16845), .Z(n16852) );
  XOR U17912 ( .A(n16853), .B(n16852), .Z(n16855) );
  XOR U17913 ( .A(n16854), .B(n16855), .Z(n16868) );
  XNOR U17914 ( .A(n16868), .B(sreg[1717]), .Z(n16870) );
  NANDN U17915 ( .A(n16847), .B(sreg[1716]), .Z(n16851) );
  NAND U17916 ( .A(n16849), .B(n16848), .Z(n16850) );
  NAND U17917 ( .A(n16851), .B(n16850), .Z(n16869) );
  XOR U17918 ( .A(n16870), .B(n16869), .Z(c[1717]) );
  NANDN U17919 ( .A(n16853), .B(n16852), .Z(n16857) );
  OR U17920 ( .A(n16855), .B(n16854), .Z(n16856) );
  AND U17921 ( .A(n16857), .B(n16856), .Z(n16875) );
  XOR U17922 ( .A(a[696]), .B(n2275), .Z(n16879) );
  AND U17923 ( .A(a[694]), .B(b[3]), .Z(n16883) );
  AND U17924 ( .A(a[698]), .B(b[0]), .Z(n16859) );
  XNOR U17925 ( .A(n16859), .B(n2175), .Z(n16861) );
  NANDN U17926 ( .A(b[0]), .B(a[697]), .Z(n16860) );
  NAND U17927 ( .A(n16861), .B(n16860), .Z(n16884) );
  XOR U17928 ( .A(n16883), .B(n16884), .Z(n16886) );
  XOR U17929 ( .A(n16885), .B(n16886), .Z(n16874) );
  NANDN U17930 ( .A(n16863), .B(n16862), .Z(n16867) );
  OR U17931 ( .A(n16865), .B(n16864), .Z(n16866) );
  AND U17932 ( .A(n16867), .B(n16866), .Z(n16873) );
  XOR U17933 ( .A(n16874), .B(n16873), .Z(n16876) );
  XOR U17934 ( .A(n16875), .B(n16876), .Z(n16889) );
  XNOR U17935 ( .A(n16889), .B(sreg[1718]), .Z(n16891) );
  NANDN U17936 ( .A(n16868), .B(sreg[1717]), .Z(n16872) );
  NAND U17937 ( .A(n16870), .B(n16869), .Z(n16871) );
  NAND U17938 ( .A(n16872), .B(n16871), .Z(n16890) );
  XOR U17939 ( .A(n16891), .B(n16890), .Z(c[1718]) );
  NANDN U17940 ( .A(n16874), .B(n16873), .Z(n16878) );
  OR U17941 ( .A(n16876), .B(n16875), .Z(n16877) );
  AND U17942 ( .A(n16878), .B(n16877), .Z(n16896) );
  XOR U17943 ( .A(a[697]), .B(n2275), .Z(n16900) );
  AND U17944 ( .A(a[695]), .B(b[3]), .Z(n16904) );
  AND U17945 ( .A(a[699]), .B(b[0]), .Z(n16880) );
  XNOR U17946 ( .A(n16880), .B(n2175), .Z(n16882) );
  NANDN U17947 ( .A(b[0]), .B(a[698]), .Z(n16881) );
  NAND U17948 ( .A(n16882), .B(n16881), .Z(n16905) );
  XOR U17949 ( .A(n16904), .B(n16905), .Z(n16907) );
  XOR U17950 ( .A(n16906), .B(n16907), .Z(n16895) );
  NANDN U17951 ( .A(n16884), .B(n16883), .Z(n16888) );
  OR U17952 ( .A(n16886), .B(n16885), .Z(n16887) );
  AND U17953 ( .A(n16888), .B(n16887), .Z(n16894) );
  XOR U17954 ( .A(n16895), .B(n16894), .Z(n16897) );
  XOR U17955 ( .A(n16896), .B(n16897), .Z(n16910) );
  XNOR U17956 ( .A(n16910), .B(sreg[1719]), .Z(n16912) );
  NANDN U17957 ( .A(n16889), .B(sreg[1718]), .Z(n16893) );
  NAND U17958 ( .A(n16891), .B(n16890), .Z(n16892) );
  NAND U17959 ( .A(n16893), .B(n16892), .Z(n16911) );
  XOR U17960 ( .A(n16912), .B(n16911), .Z(c[1719]) );
  NANDN U17961 ( .A(n16895), .B(n16894), .Z(n16899) );
  OR U17962 ( .A(n16897), .B(n16896), .Z(n16898) );
  AND U17963 ( .A(n16899), .B(n16898), .Z(n16917) );
  XOR U17964 ( .A(a[698]), .B(n2275), .Z(n16921) );
  AND U17965 ( .A(a[700]), .B(b[0]), .Z(n16901) );
  XNOR U17966 ( .A(n16901), .B(n2175), .Z(n16903) );
  NANDN U17967 ( .A(b[0]), .B(a[699]), .Z(n16902) );
  NAND U17968 ( .A(n16903), .B(n16902), .Z(n16926) );
  AND U17969 ( .A(a[696]), .B(b[3]), .Z(n16925) );
  XOR U17970 ( .A(n16926), .B(n16925), .Z(n16928) );
  XOR U17971 ( .A(n16927), .B(n16928), .Z(n16916) );
  NANDN U17972 ( .A(n16905), .B(n16904), .Z(n16909) );
  OR U17973 ( .A(n16907), .B(n16906), .Z(n16908) );
  AND U17974 ( .A(n16909), .B(n16908), .Z(n16915) );
  XOR U17975 ( .A(n16916), .B(n16915), .Z(n16918) );
  XOR U17976 ( .A(n16917), .B(n16918), .Z(n16931) );
  XNOR U17977 ( .A(n16931), .B(sreg[1720]), .Z(n16933) );
  NANDN U17978 ( .A(n16910), .B(sreg[1719]), .Z(n16914) );
  NAND U17979 ( .A(n16912), .B(n16911), .Z(n16913) );
  NAND U17980 ( .A(n16914), .B(n16913), .Z(n16932) );
  XOR U17981 ( .A(n16933), .B(n16932), .Z(c[1720]) );
  NANDN U17982 ( .A(n16916), .B(n16915), .Z(n16920) );
  OR U17983 ( .A(n16918), .B(n16917), .Z(n16919) );
  AND U17984 ( .A(n16920), .B(n16919), .Z(n16938) );
  XOR U17985 ( .A(a[699]), .B(n2276), .Z(n16942) );
  AND U17986 ( .A(a[701]), .B(b[0]), .Z(n16922) );
  XNOR U17987 ( .A(n16922), .B(n2175), .Z(n16924) );
  NANDN U17988 ( .A(b[0]), .B(a[700]), .Z(n16923) );
  NAND U17989 ( .A(n16924), .B(n16923), .Z(n16947) );
  AND U17990 ( .A(a[697]), .B(b[3]), .Z(n16946) );
  XOR U17991 ( .A(n16947), .B(n16946), .Z(n16949) );
  XOR U17992 ( .A(n16948), .B(n16949), .Z(n16937) );
  NANDN U17993 ( .A(n16926), .B(n16925), .Z(n16930) );
  OR U17994 ( .A(n16928), .B(n16927), .Z(n16929) );
  AND U17995 ( .A(n16930), .B(n16929), .Z(n16936) );
  XOR U17996 ( .A(n16937), .B(n16936), .Z(n16939) );
  XOR U17997 ( .A(n16938), .B(n16939), .Z(n16952) );
  XNOR U17998 ( .A(n16952), .B(sreg[1721]), .Z(n16954) );
  NANDN U17999 ( .A(n16931), .B(sreg[1720]), .Z(n16935) );
  NAND U18000 ( .A(n16933), .B(n16932), .Z(n16934) );
  NAND U18001 ( .A(n16935), .B(n16934), .Z(n16953) );
  XOR U18002 ( .A(n16954), .B(n16953), .Z(c[1721]) );
  NANDN U18003 ( .A(n16937), .B(n16936), .Z(n16941) );
  OR U18004 ( .A(n16939), .B(n16938), .Z(n16940) );
  AND U18005 ( .A(n16941), .B(n16940), .Z(n16959) );
  XOR U18006 ( .A(a[700]), .B(n2276), .Z(n16963) );
  AND U18007 ( .A(a[702]), .B(b[0]), .Z(n16943) );
  XNOR U18008 ( .A(n16943), .B(n2175), .Z(n16945) );
  NANDN U18009 ( .A(b[0]), .B(a[701]), .Z(n16944) );
  NAND U18010 ( .A(n16945), .B(n16944), .Z(n16968) );
  AND U18011 ( .A(a[698]), .B(b[3]), .Z(n16967) );
  XOR U18012 ( .A(n16968), .B(n16967), .Z(n16970) );
  XOR U18013 ( .A(n16969), .B(n16970), .Z(n16958) );
  NANDN U18014 ( .A(n16947), .B(n16946), .Z(n16951) );
  OR U18015 ( .A(n16949), .B(n16948), .Z(n16950) );
  AND U18016 ( .A(n16951), .B(n16950), .Z(n16957) );
  XOR U18017 ( .A(n16958), .B(n16957), .Z(n16960) );
  XOR U18018 ( .A(n16959), .B(n16960), .Z(n16973) );
  XNOR U18019 ( .A(n16973), .B(sreg[1722]), .Z(n16975) );
  NANDN U18020 ( .A(n16952), .B(sreg[1721]), .Z(n16956) );
  NAND U18021 ( .A(n16954), .B(n16953), .Z(n16955) );
  NAND U18022 ( .A(n16956), .B(n16955), .Z(n16974) );
  XOR U18023 ( .A(n16975), .B(n16974), .Z(c[1722]) );
  NANDN U18024 ( .A(n16958), .B(n16957), .Z(n16962) );
  OR U18025 ( .A(n16960), .B(n16959), .Z(n16961) );
  AND U18026 ( .A(n16962), .B(n16961), .Z(n16980) );
  XOR U18027 ( .A(a[701]), .B(n2276), .Z(n16984) );
  AND U18028 ( .A(a[699]), .B(b[3]), .Z(n16988) );
  AND U18029 ( .A(a[703]), .B(b[0]), .Z(n16964) );
  XNOR U18030 ( .A(n16964), .B(n2175), .Z(n16966) );
  NANDN U18031 ( .A(b[0]), .B(a[702]), .Z(n16965) );
  NAND U18032 ( .A(n16966), .B(n16965), .Z(n16989) );
  XOR U18033 ( .A(n16988), .B(n16989), .Z(n16991) );
  XOR U18034 ( .A(n16990), .B(n16991), .Z(n16979) );
  NANDN U18035 ( .A(n16968), .B(n16967), .Z(n16972) );
  OR U18036 ( .A(n16970), .B(n16969), .Z(n16971) );
  AND U18037 ( .A(n16972), .B(n16971), .Z(n16978) );
  XOR U18038 ( .A(n16979), .B(n16978), .Z(n16981) );
  XOR U18039 ( .A(n16980), .B(n16981), .Z(n16994) );
  XNOR U18040 ( .A(n16994), .B(sreg[1723]), .Z(n16996) );
  NANDN U18041 ( .A(n16973), .B(sreg[1722]), .Z(n16977) );
  NAND U18042 ( .A(n16975), .B(n16974), .Z(n16976) );
  NAND U18043 ( .A(n16977), .B(n16976), .Z(n16995) );
  XOR U18044 ( .A(n16996), .B(n16995), .Z(c[1723]) );
  NANDN U18045 ( .A(n16979), .B(n16978), .Z(n16983) );
  OR U18046 ( .A(n16981), .B(n16980), .Z(n16982) );
  AND U18047 ( .A(n16983), .B(n16982), .Z(n17001) );
  XOR U18048 ( .A(a[702]), .B(n2276), .Z(n17005) );
  AND U18049 ( .A(a[704]), .B(b[0]), .Z(n16985) );
  XNOR U18050 ( .A(n16985), .B(n2175), .Z(n16987) );
  NANDN U18051 ( .A(b[0]), .B(a[703]), .Z(n16986) );
  NAND U18052 ( .A(n16987), .B(n16986), .Z(n17010) );
  AND U18053 ( .A(a[700]), .B(b[3]), .Z(n17009) );
  XOR U18054 ( .A(n17010), .B(n17009), .Z(n17012) );
  XOR U18055 ( .A(n17011), .B(n17012), .Z(n17000) );
  NANDN U18056 ( .A(n16989), .B(n16988), .Z(n16993) );
  OR U18057 ( .A(n16991), .B(n16990), .Z(n16992) );
  AND U18058 ( .A(n16993), .B(n16992), .Z(n16999) );
  XOR U18059 ( .A(n17000), .B(n16999), .Z(n17002) );
  XOR U18060 ( .A(n17001), .B(n17002), .Z(n17015) );
  XNOR U18061 ( .A(n17015), .B(sreg[1724]), .Z(n17017) );
  NANDN U18062 ( .A(n16994), .B(sreg[1723]), .Z(n16998) );
  NAND U18063 ( .A(n16996), .B(n16995), .Z(n16997) );
  NAND U18064 ( .A(n16998), .B(n16997), .Z(n17016) );
  XOR U18065 ( .A(n17017), .B(n17016), .Z(c[1724]) );
  NANDN U18066 ( .A(n17000), .B(n16999), .Z(n17004) );
  OR U18067 ( .A(n17002), .B(n17001), .Z(n17003) );
  AND U18068 ( .A(n17004), .B(n17003), .Z(n17022) );
  XOR U18069 ( .A(a[703]), .B(n2276), .Z(n17026) );
  AND U18070 ( .A(a[701]), .B(b[3]), .Z(n17030) );
  AND U18071 ( .A(a[705]), .B(b[0]), .Z(n17006) );
  XNOR U18072 ( .A(n17006), .B(n2175), .Z(n17008) );
  NANDN U18073 ( .A(b[0]), .B(a[704]), .Z(n17007) );
  NAND U18074 ( .A(n17008), .B(n17007), .Z(n17031) );
  XOR U18075 ( .A(n17030), .B(n17031), .Z(n17033) );
  XOR U18076 ( .A(n17032), .B(n17033), .Z(n17021) );
  NANDN U18077 ( .A(n17010), .B(n17009), .Z(n17014) );
  OR U18078 ( .A(n17012), .B(n17011), .Z(n17013) );
  AND U18079 ( .A(n17014), .B(n17013), .Z(n17020) );
  XOR U18080 ( .A(n17021), .B(n17020), .Z(n17023) );
  XOR U18081 ( .A(n17022), .B(n17023), .Z(n17036) );
  XNOR U18082 ( .A(n17036), .B(sreg[1725]), .Z(n17038) );
  NANDN U18083 ( .A(n17015), .B(sreg[1724]), .Z(n17019) );
  NAND U18084 ( .A(n17017), .B(n17016), .Z(n17018) );
  NAND U18085 ( .A(n17019), .B(n17018), .Z(n17037) );
  XOR U18086 ( .A(n17038), .B(n17037), .Z(c[1725]) );
  NANDN U18087 ( .A(n17021), .B(n17020), .Z(n17025) );
  OR U18088 ( .A(n17023), .B(n17022), .Z(n17024) );
  AND U18089 ( .A(n17025), .B(n17024), .Z(n17043) );
  XOR U18090 ( .A(a[704]), .B(n2276), .Z(n17047) );
  AND U18091 ( .A(a[706]), .B(b[0]), .Z(n17027) );
  XNOR U18092 ( .A(n17027), .B(n2175), .Z(n17029) );
  NANDN U18093 ( .A(b[0]), .B(a[705]), .Z(n17028) );
  NAND U18094 ( .A(n17029), .B(n17028), .Z(n17052) );
  AND U18095 ( .A(a[702]), .B(b[3]), .Z(n17051) );
  XOR U18096 ( .A(n17052), .B(n17051), .Z(n17054) );
  XOR U18097 ( .A(n17053), .B(n17054), .Z(n17042) );
  NANDN U18098 ( .A(n17031), .B(n17030), .Z(n17035) );
  OR U18099 ( .A(n17033), .B(n17032), .Z(n17034) );
  AND U18100 ( .A(n17035), .B(n17034), .Z(n17041) );
  XOR U18101 ( .A(n17042), .B(n17041), .Z(n17044) );
  XOR U18102 ( .A(n17043), .B(n17044), .Z(n17057) );
  XNOR U18103 ( .A(n17057), .B(sreg[1726]), .Z(n17059) );
  NANDN U18104 ( .A(n17036), .B(sreg[1725]), .Z(n17040) );
  NAND U18105 ( .A(n17038), .B(n17037), .Z(n17039) );
  NAND U18106 ( .A(n17040), .B(n17039), .Z(n17058) );
  XOR U18107 ( .A(n17059), .B(n17058), .Z(c[1726]) );
  NANDN U18108 ( .A(n17042), .B(n17041), .Z(n17046) );
  OR U18109 ( .A(n17044), .B(n17043), .Z(n17045) );
  AND U18110 ( .A(n17046), .B(n17045), .Z(n17064) );
  XOR U18111 ( .A(a[705]), .B(n2276), .Z(n17068) );
  AND U18112 ( .A(a[703]), .B(b[3]), .Z(n17072) );
  AND U18113 ( .A(a[707]), .B(b[0]), .Z(n17048) );
  XNOR U18114 ( .A(n17048), .B(n2175), .Z(n17050) );
  NANDN U18115 ( .A(b[0]), .B(a[706]), .Z(n17049) );
  NAND U18116 ( .A(n17050), .B(n17049), .Z(n17073) );
  XOR U18117 ( .A(n17072), .B(n17073), .Z(n17075) );
  XOR U18118 ( .A(n17074), .B(n17075), .Z(n17063) );
  NANDN U18119 ( .A(n17052), .B(n17051), .Z(n17056) );
  OR U18120 ( .A(n17054), .B(n17053), .Z(n17055) );
  AND U18121 ( .A(n17056), .B(n17055), .Z(n17062) );
  XOR U18122 ( .A(n17063), .B(n17062), .Z(n17065) );
  XOR U18123 ( .A(n17064), .B(n17065), .Z(n17078) );
  XNOR U18124 ( .A(n17078), .B(sreg[1727]), .Z(n17080) );
  NANDN U18125 ( .A(n17057), .B(sreg[1726]), .Z(n17061) );
  NAND U18126 ( .A(n17059), .B(n17058), .Z(n17060) );
  NAND U18127 ( .A(n17061), .B(n17060), .Z(n17079) );
  XOR U18128 ( .A(n17080), .B(n17079), .Z(c[1727]) );
  NANDN U18129 ( .A(n17063), .B(n17062), .Z(n17067) );
  OR U18130 ( .A(n17065), .B(n17064), .Z(n17066) );
  AND U18131 ( .A(n17067), .B(n17066), .Z(n17085) );
  XOR U18132 ( .A(a[706]), .B(n2277), .Z(n17089) );
  AND U18133 ( .A(a[708]), .B(b[0]), .Z(n17069) );
  XNOR U18134 ( .A(n17069), .B(n2175), .Z(n17071) );
  NANDN U18135 ( .A(b[0]), .B(a[707]), .Z(n17070) );
  NAND U18136 ( .A(n17071), .B(n17070), .Z(n17094) );
  AND U18137 ( .A(a[704]), .B(b[3]), .Z(n17093) );
  XOR U18138 ( .A(n17094), .B(n17093), .Z(n17096) );
  XOR U18139 ( .A(n17095), .B(n17096), .Z(n17084) );
  NANDN U18140 ( .A(n17073), .B(n17072), .Z(n17077) );
  OR U18141 ( .A(n17075), .B(n17074), .Z(n17076) );
  AND U18142 ( .A(n17077), .B(n17076), .Z(n17083) );
  XOR U18143 ( .A(n17084), .B(n17083), .Z(n17086) );
  XOR U18144 ( .A(n17085), .B(n17086), .Z(n17099) );
  XNOR U18145 ( .A(n17099), .B(sreg[1728]), .Z(n17101) );
  NANDN U18146 ( .A(n17078), .B(sreg[1727]), .Z(n17082) );
  NAND U18147 ( .A(n17080), .B(n17079), .Z(n17081) );
  NAND U18148 ( .A(n17082), .B(n17081), .Z(n17100) );
  XOR U18149 ( .A(n17101), .B(n17100), .Z(c[1728]) );
  NANDN U18150 ( .A(n17084), .B(n17083), .Z(n17088) );
  OR U18151 ( .A(n17086), .B(n17085), .Z(n17087) );
  AND U18152 ( .A(n17088), .B(n17087), .Z(n17106) );
  XOR U18153 ( .A(a[707]), .B(n2277), .Z(n17110) );
  AND U18154 ( .A(a[705]), .B(b[3]), .Z(n17114) );
  AND U18155 ( .A(a[709]), .B(b[0]), .Z(n17090) );
  XNOR U18156 ( .A(n17090), .B(n2175), .Z(n17092) );
  NANDN U18157 ( .A(b[0]), .B(a[708]), .Z(n17091) );
  NAND U18158 ( .A(n17092), .B(n17091), .Z(n17115) );
  XOR U18159 ( .A(n17114), .B(n17115), .Z(n17117) );
  XOR U18160 ( .A(n17116), .B(n17117), .Z(n17105) );
  NANDN U18161 ( .A(n17094), .B(n17093), .Z(n17098) );
  OR U18162 ( .A(n17096), .B(n17095), .Z(n17097) );
  AND U18163 ( .A(n17098), .B(n17097), .Z(n17104) );
  XOR U18164 ( .A(n17105), .B(n17104), .Z(n17107) );
  XOR U18165 ( .A(n17106), .B(n17107), .Z(n17120) );
  XNOR U18166 ( .A(n17120), .B(sreg[1729]), .Z(n17122) );
  NANDN U18167 ( .A(n17099), .B(sreg[1728]), .Z(n17103) );
  NAND U18168 ( .A(n17101), .B(n17100), .Z(n17102) );
  NAND U18169 ( .A(n17103), .B(n17102), .Z(n17121) );
  XOR U18170 ( .A(n17122), .B(n17121), .Z(c[1729]) );
  NANDN U18171 ( .A(n17105), .B(n17104), .Z(n17109) );
  OR U18172 ( .A(n17107), .B(n17106), .Z(n17108) );
  AND U18173 ( .A(n17109), .B(n17108), .Z(n17127) );
  XOR U18174 ( .A(a[708]), .B(n2277), .Z(n17131) );
  AND U18175 ( .A(a[710]), .B(b[0]), .Z(n17111) );
  XNOR U18176 ( .A(n17111), .B(n2175), .Z(n17113) );
  NANDN U18177 ( .A(b[0]), .B(a[709]), .Z(n17112) );
  NAND U18178 ( .A(n17113), .B(n17112), .Z(n17136) );
  AND U18179 ( .A(a[706]), .B(b[3]), .Z(n17135) );
  XOR U18180 ( .A(n17136), .B(n17135), .Z(n17138) );
  XOR U18181 ( .A(n17137), .B(n17138), .Z(n17126) );
  NANDN U18182 ( .A(n17115), .B(n17114), .Z(n17119) );
  OR U18183 ( .A(n17117), .B(n17116), .Z(n17118) );
  AND U18184 ( .A(n17119), .B(n17118), .Z(n17125) );
  XOR U18185 ( .A(n17126), .B(n17125), .Z(n17128) );
  XOR U18186 ( .A(n17127), .B(n17128), .Z(n17141) );
  XNOR U18187 ( .A(n17141), .B(sreg[1730]), .Z(n17143) );
  NANDN U18188 ( .A(n17120), .B(sreg[1729]), .Z(n17124) );
  NAND U18189 ( .A(n17122), .B(n17121), .Z(n17123) );
  NAND U18190 ( .A(n17124), .B(n17123), .Z(n17142) );
  XOR U18191 ( .A(n17143), .B(n17142), .Z(c[1730]) );
  NANDN U18192 ( .A(n17126), .B(n17125), .Z(n17130) );
  OR U18193 ( .A(n17128), .B(n17127), .Z(n17129) );
  AND U18194 ( .A(n17130), .B(n17129), .Z(n17148) );
  XOR U18195 ( .A(a[709]), .B(n2277), .Z(n17152) );
  AND U18196 ( .A(a[711]), .B(b[0]), .Z(n17132) );
  XNOR U18197 ( .A(n17132), .B(n2175), .Z(n17134) );
  NANDN U18198 ( .A(b[0]), .B(a[710]), .Z(n17133) );
  NAND U18199 ( .A(n17134), .B(n17133), .Z(n17157) );
  AND U18200 ( .A(a[707]), .B(b[3]), .Z(n17156) );
  XOR U18201 ( .A(n17157), .B(n17156), .Z(n17159) );
  XOR U18202 ( .A(n17158), .B(n17159), .Z(n17147) );
  NANDN U18203 ( .A(n17136), .B(n17135), .Z(n17140) );
  OR U18204 ( .A(n17138), .B(n17137), .Z(n17139) );
  AND U18205 ( .A(n17140), .B(n17139), .Z(n17146) );
  XOR U18206 ( .A(n17147), .B(n17146), .Z(n17149) );
  XOR U18207 ( .A(n17148), .B(n17149), .Z(n17162) );
  XNOR U18208 ( .A(n17162), .B(sreg[1731]), .Z(n17164) );
  NANDN U18209 ( .A(n17141), .B(sreg[1730]), .Z(n17145) );
  NAND U18210 ( .A(n17143), .B(n17142), .Z(n17144) );
  NAND U18211 ( .A(n17145), .B(n17144), .Z(n17163) );
  XOR U18212 ( .A(n17164), .B(n17163), .Z(c[1731]) );
  NANDN U18213 ( .A(n17147), .B(n17146), .Z(n17151) );
  OR U18214 ( .A(n17149), .B(n17148), .Z(n17150) );
  AND U18215 ( .A(n17151), .B(n17150), .Z(n17169) );
  XOR U18216 ( .A(a[710]), .B(n2277), .Z(n17173) );
  AND U18217 ( .A(a[708]), .B(b[3]), .Z(n17177) );
  AND U18218 ( .A(a[712]), .B(b[0]), .Z(n17153) );
  XNOR U18219 ( .A(n17153), .B(n2175), .Z(n17155) );
  NANDN U18220 ( .A(b[0]), .B(a[711]), .Z(n17154) );
  NAND U18221 ( .A(n17155), .B(n17154), .Z(n17178) );
  XOR U18222 ( .A(n17177), .B(n17178), .Z(n17180) );
  XOR U18223 ( .A(n17179), .B(n17180), .Z(n17168) );
  NANDN U18224 ( .A(n17157), .B(n17156), .Z(n17161) );
  OR U18225 ( .A(n17159), .B(n17158), .Z(n17160) );
  AND U18226 ( .A(n17161), .B(n17160), .Z(n17167) );
  XOR U18227 ( .A(n17168), .B(n17167), .Z(n17170) );
  XOR U18228 ( .A(n17169), .B(n17170), .Z(n17183) );
  XNOR U18229 ( .A(n17183), .B(sreg[1732]), .Z(n17185) );
  NANDN U18230 ( .A(n17162), .B(sreg[1731]), .Z(n17166) );
  NAND U18231 ( .A(n17164), .B(n17163), .Z(n17165) );
  NAND U18232 ( .A(n17166), .B(n17165), .Z(n17184) );
  XOR U18233 ( .A(n17185), .B(n17184), .Z(c[1732]) );
  NANDN U18234 ( .A(n17168), .B(n17167), .Z(n17172) );
  OR U18235 ( .A(n17170), .B(n17169), .Z(n17171) );
  AND U18236 ( .A(n17172), .B(n17171), .Z(n17190) );
  XOR U18237 ( .A(a[711]), .B(n2277), .Z(n17194) );
  AND U18238 ( .A(a[713]), .B(b[0]), .Z(n17174) );
  XNOR U18239 ( .A(n17174), .B(n2175), .Z(n17176) );
  NANDN U18240 ( .A(b[0]), .B(a[712]), .Z(n17175) );
  NAND U18241 ( .A(n17176), .B(n17175), .Z(n17199) );
  AND U18242 ( .A(a[709]), .B(b[3]), .Z(n17198) );
  XOR U18243 ( .A(n17199), .B(n17198), .Z(n17201) );
  XOR U18244 ( .A(n17200), .B(n17201), .Z(n17189) );
  NANDN U18245 ( .A(n17178), .B(n17177), .Z(n17182) );
  OR U18246 ( .A(n17180), .B(n17179), .Z(n17181) );
  AND U18247 ( .A(n17182), .B(n17181), .Z(n17188) );
  XOR U18248 ( .A(n17189), .B(n17188), .Z(n17191) );
  XOR U18249 ( .A(n17190), .B(n17191), .Z(n17204) );
  XNOR U18250 ( .A(n17204), .B(sreg[1733]), .Z(n17206) );
  NANDN U18251 ( .A(n17183), .B(sreg[1732]), .Z(n17187) );
  NAND U18252 ( .A(n17185), .B(n17184), .Z(n17186) );
  NAND U18253 ( .A(n17187), .B(n17186), .Z(n17205) );
  XOR U18254 ( .A(n17206), .B(n17205), .Z(c[1733]) );
  NANDN U18255 ( .A(n17189), .B(n17188), .Z(n17193) );
  OR U18256 ( .A(n17191), .B(n17190), .Z(n17192) );
  AND U18257 ( .A(n17193), .B(n17192), .Z(n17211) );
  XOR U18258 ( .A(a[712]), .B(n2277), .Z(n17215) );
  AND U18259 ( .A(a[710]), .B(b[3]), .Z(n17219) );
  AND U18260 ( .A(a[714]), .B(b[0]), .Z(n17195) );
  XNOR U18261 ( .A(n17195), .B(n2175), .Z(n17197) );
  NANDN U18262 ( .A(b[0]), .B(a[713]), .Z(n17196) );
  NAND U18263 ( .A(n17197), .B(n17196), .Z(n17220) );
  XOR U18264 ( .A(n17219), .B(n17220), .Z(n17222) );
  XOR U18265 ( .A(n17221), .B(n17222), .Z(n17210) );
  NANDN U18266 ( .A(n17199), .B(n17198), .Z(n17203) );
  OR U18267 ( .A(n17201), .B(n17200), .Z(n17202) );
  AND U18268 ( .A(n17203), .B(n17202), .Z(n17209) );
  XOR U18269 ( .A(n17210), .B(n17209), .Z(n17212) );
  XOR U18270 ( .A(n17211), .B(n17212), .Z(n17225) );
  XNOR U18271 ( .A(n17225), .B(sreg[1734]), .Z(n17227) );
  NANDN U18272 ( .A(n17204), .B(sreg[1733]), .Z(n17208) );
  NAND U18273 ( .A(n17206), .B(n17205), .Z(n17207) );
  NAND U18274 ( .A(n17208), .B(n17207), .Z(n17226) );
  XOR U18275 ( .A(n17227), .B(n17226), .Z(c[1734]) );
  NANDN U18276 ( .A(n17210), .B(n17209), .Z(n17214) );
  OR U18277 ( .A(n17212), .B(n17211), .Z(n17213) );
  AND U18278 ( .A(n17214), .B(n17213), .Z(n17232) );
  XOR U18279 ( .A(a[713]), .B(n2278), .Z(n17236) );
  AND U18280 ( .A(a[711]), .B(b[3]), .Z(n17240) );
  AND U18281 ( .A(a[715]), .B(b[0]), .Z(n17216) );
  XNOR U18282 ( .A(n17216), .B(n2175), .Z(n17218) );
  NANDN U18283 ( .A(b[0]), .B(a[714]), .Z(n17217) );
  NAND U18284 ( .A(n17218), .B(n17217), .Z(n17241) );
  XOR U18285 ( .A(n17240), .B(n17241), .Z(n17243) );
  XOR U18286 ( .A(n17242), .B(n17243), .Z(n17231) );
  NANDN U18287 ( .A(n17220), .B(n17219), .Z(n17224) );
  OR U18288 ( .A(n17222), .B(n17221), .Z(n17223) );
  AND U18289 ( .A(n17224), .B(n17223), .Z(n17230) );
  XOR U18290 ( .A(n17231), .B(n17230), .Z(n17233) );
  XOR U18291 ( .A(n17232), .B(n17233), .Z(n17246) );
  XNOR U18292 ( .A(n17246), .B(sreg[1735]), .Z(n17248) );
  NANDN U18293 ( .A(n17225), .B(sreg[1734]), .Z(n17229) );
  NAND U18294 ( .A(n17227), .B(n17226), .Z(n17228) );
  NAND U18295 ( .A(n17229), .B(n17228), .Z(n17247) );
  XOR U18296 ( .A(n17248), .B(n17247), .Z(c[1735]) );
  NANDN U18297 ( .A(n17231), .B(n17230), .Z(n17235) );
  OR U18298 ( .A(n17233), .B(n17232), .Z(n17234) );
  AND U18299 ( .A(n17235), .B(n17234), .Z(n17253) );
  XOR U18300 ( .A(a[714]), .B(n2278), .Z(n17257) );
  AND U18301 ( .A(a[716]), .B(b[0]), .Z(n17237) );
  XNOR U18302 ( .A(n17237), .B(n2175), .Z(n17239) );
  NANDN U18303 ( .A(b[0]), .B(a[715]), .Z(n17238) );
  NAND U18304 ( .A(n17239), .B(n17238), .Z(n17262) );
  AND U18305 ( .A(a[712]), .B(b[3]), .Z(n17261) );
  XOR U18306 ( .A(n17262), .B(n17261), .Z(n17264) );
  XOR U18307 ( .A(n17263), .B(n17264), .Z(n17252) );
  NANDN U18308 ( .A(n17241), .B(n17240), .Z(n17245) );
  OR U18309 ( .A(n17243), .B(n17242), .Z(n17244) );
  AND U18310 ( .A(n17245), .B(n17244), .Z(n17251) );
  XOR U18311 ( .A(n17252), .B(n17251), .Z(n17254) );
  XOR U18312 ( .A(n17253), .B(n17254), .Z(n17267) );
  XNOR U18313 ( .A(n17267), .B(sreg[1736]), .Z(n17269) );
  NANDN U18314 ( .A(n17246), .B(sreg[1735]), .Z(n17250) );
  NAND U18315 ( .A(n17248), .B(n17247), .Z(n17249) );
  NAND U18316 ( .A(n17250), .B(n17249), .Z(n17268) );
  XOR U18317 ( .A(n17269), .B(n17268), .Z(c[1736]) );
  NANDN U18318 ( .A(n17252), .B(n17251), .Z(n17256) );
  OR U18319 ( .A(n17254), .B(n17253), .Z(n17255) );
  AND U18320 ( .A(n17256), .B(n17255), .Z(n17274) );
  XOR U18321 ( .A(a[715]), .B(n2278), .Z(n17278) );
  AND U18322 ( .A(a[717]), .B(b[0]), .Z(n17258) );
  XNOR U18323 ( .A(n17258), .B(n2175), .Z(n17260) );
  NANDN U18324 ( .A(b[0]), .B(a[716]), .Z(n17259) );
  NAND U18325 ( .A(n17260), .B(n17259), .Z(n17283) );
  AND U18326 ( .A(a[713]), .B(b[3]), .Z(n17282) );
  XOR U18327 ( .A(n17283), .B(n17282), .Z(n17285) );
  XOR U18328 ( .A(n17284), .B(n17285), .Z(n17273) );
  NANDN U18329 ( .A(n17262), .B(n17261), .Z(n17266) );
  OR U18330 ( .A(n17264), .B(n17263), .Z(n17265) );
  AND U18331 ( .A(n17266), .B(n17265), .Z(n17272) );
  XOR U18332 ( .A(n17273), .B(n17272), .Z(n17275) );
  XOR U18333 ( .A(n17274), .B(n17275), .Z(n17288) );
  XNOR U18334 ( .A(n17288), .B(sreg[1737]), .Z(n17290) );
  NANDN U18335 ( .A(n17267), .B(sreg[1736]), .Z(n17271) );
  NAND U18336 ( .A(n17269), .B(n17268), .Z(n17270) );
  NAND U18337 ( .A(n17271), .B(n17270), .Z(n17289) );
  XOR U18338 ( .A(n17290), .B(n17289), .Z(c[1737]) );
  NANDN U18339 ( .A(n17273), .B(n17272), .Z(n17277) );
  OR U18340 ( .A(n17275), .B(n17274), .Z(n17276) );
  AND U18341 ( .A(n17277), .B(n17276), .Z(n17295) );
  XOR U18342 ( .A(a[716]), .B(n2278), .Z(n17299) );
  AND U18343 ( .A(a[714]), .B(b[3]), .Z(n17303) );
  AND U18344 ( .A(a[718]), .B(b[0]), .Z(n17279) );
  XNOR U18345 ( .A(n17279), .B(n2175), .Z(n17281) );
  NANDN U18346 ( .A(b[0]), .B(a[717]), .Z(n17280) );
  NAND U18347 ( .A(n17281), .B(n17280), .Z(n17304) );
  XOR U18348 ( .A(n17303), .B(n17304), .Z(n17306) );
  XOR U18349 ( .A(n17305), .B(n17306), .Z(n17294) );
  NANDN U18350 ( .A(n17283), .B(n17282), .Z(n17287) );
  OR U18351 ( .A(n17285), .B(n17284), .Z(n17286) );
  AND U18352 ( .A(n17287), .B(n17286), .Z(n17293) );
  XOR U18353 ( .A(n17294), .B(n17293), .Z(n17296) );
  XOR U18354 ( .A(n17295), .B(n17296), .Z(n17309) );
  XNOR U18355 ( .A(n17309), .B(sreg[1738]), .Z(n17311) );
  NANDN U18356 ( .A(n17288), .B(sreg[1737]), .Z(n17292) );
  NAND U18357 ( .A(n17290), .B(n17289), .Z(n17291) );
  NAND U18358 ( .A(n17292), .B(n17291), .Z(n17310) );
  XOR U18359 ( .A(n17311), .B(n17310), .Z(c[1738]) );
  NANDN U18360 ( .A(n17294), .B(n17293), .Z(n17298) );
  OR U18361 ( .A(n17296), .B(n17295), .Z(n17297) );
  AND U18362 ( .A(n17298), .B(n17297), .Z(n17316) );
  XOR U18363 ( .A(a[717]), .B(n2278), .Z(n17320) );
  AND U18364 ( .A(a[719]), .B(b[0]), .Z(n17300) );
  XNOR U18365 ( .A(n17300), .B(n2175), .Z(n17302) );
  NANDN U18366 ( .A(b[0]), .B(a[718]), .Z(n17301) );
  NAND U18367 ( .A(n17302), .B(n17301), .Z(n17325) );
  AND U18368 ( .A(a[715]), .B(b[3]), .Z(n17324) );
  XOR U18369 ( .A(n17325), .B(n17324), .Z(n17327) );
  XOR U18370 ( .A(n17326), .B(n17327), .Z(n17315) );
  NANDN U18371 ( .A(n17304), .B(n17303), .Z(n17308) );
  OR U18372 ( .A(n17306), .B(n17305), .Z(n17307) );
  AND U18373 ( .A(n17308), .B(n17307), .Z(n17314) );
  XOR U18374 ( .A(n17315), .B(n17314), .Z(n17317) );
  XOR U18375 ( .A(n17316), .B(n17317), .Z(n17330) );
  XNOR U18376 ( .A(n17330), .B(sreg[1739]), .Z(n17332) );
  NANDN U18377 ( .A(n17309), .B(sreg[1738]), .Z(n17313) );
  NAND U18378 ( .A(n17311), .B(n17310), .Z(n17312) );
  NAND U18379 ( .A(n17313), .B(n17312), .Z(n17331) );
  XOR U18380 ( .A(n17332), .B(n17331), .Z(c[1739]) );
  NANDN U18381 ( .A(n17315), .B(n17314), .Z(n17319) );
  OR U18382 ( .A(n17317), .B(n17316), .Z(n17318) );
  AND U18383 ( .A(n17319), .B(n17318), .Z(n17337) );
  XOR U18384 ( .A(a[718]), .B(n2278), .Z(n17341) );
  AND U18385 ( .A(a[720]), .B(b[0]), .Z(n17321) );
  XNOR U18386 ( .A(n17321), .B(n2175), .Z(n17323) );
  NANDN U18387 ( .A(b[0]), .B(a[719]), .Z(n17322) );
  NAND U18388 ( .A(n17323), .B(n17322), .Z(n17346) );
  AND U18389 ( .A(a[716]), .B(b[3]), .Z(n17345) );
  XOR U18390 ( .A(n17346), .B(n17345), .Z(n17348) );
  XOR U18391 ( .A(n17347), .B(n17348), .Z(n17336) );
  NANDN U18392 ( .A(n17325), .B(n17324), .Z(n17329) );
  OR U18393 ( .A(n17327), .B(n17326), .Z(n17328) );
  AND U18394 ( .A(n17329), .B(n17328), .Z(n17335) );
  XOR U18395 ( .A(n17336), .B(n17335), .Z(n17338) );
  XOR U18396 ( .A(n17337), .B(n17338), .Z(n17351) );
  XNOR U18397 ( .A(n17351), .B(sreg[1740]), .Z(n17353) );
  NANDN U18398 ( .A(n17330), .B(sreg[1739]), .Z(n17334) );
  NAND U18399 ( .A(n17332), .B(n17331), .Z(n17333) );
  NAND U18400 ( .A(n17334), .B(n17333), .Z(n17352) );
  XOR U18401 ( .A(n17353), .B(n17352), .Z(c[1740]) );
  NANDN U18402 ( .A(n17336), .B(n17335), .Z(n17340) );
  OR U18403 ( .A(n17338), .B(n17337), .Z(n17339) );
  AND U18404 ( .A(n17340), .B(n17339), .Z(n17358) );
  XOR U18405 ( .A(a[719]), .B(n2278), .Z(n17362) );
  AND U18406 ( .A(a[721]), .B(b[0]), .Z(n17342) );
  XNOR U18407 ( .A(n17342), .B(n2175), .Z(n17344) );
  NANDN U18408 ( .A(b[0]), .B(a[720]), .Z(n17343) );
  NAND U18409 ( .A(n17344), .B(n17343), .Z(n17367) );
  AND U18410 ( .A(a[717]), .B(b[3]), .Z(n17366) );
  XOR U18411 ( .A(n17367), .B(n17366), .Z(n17369) );
  XOR U18412 ( .A(n17368), .B(n17369), .Z(n17357) );
  NANDN U18413 ( .A(n17346), .B(n17345), .Z(n17350) );
  OR U18414 ( .A(n17348), .B(n17347), .Z(n17349) );
  AND U18415 ( .A(n17350), .B(n17349), .Z(n17356) );
  XOR U18416 ( .A(n17357), .B(n17356), .Z(n17359) );
  XOR U18417 ( .A(n17358), .B(n17359), .Z(n17372) );
  XNOR U18418 ( .A(n17372), .B(sreg[1741]), .Z(n17374) );
  NANDN U18419 ( .A(n17351), .B(sreg[1740]), .Z(n17355) );
  NAND U18420 ( .A(n17353), .B(n17352), .Z(n17354) );
  NAND U18421 ( .A(n17355), .B(n17354), .Z(n17373) );
  XOR U18422 ( .A(n17374), .B(n17373), .Z(c[1741]) );
  NANDN U18423 ( .A(n17357), .B(n17356), .Z(n17361) );
  OR U18424 ( .A(n17359), .B(n17358), .Z(n17360) );
  AND U18425 ( .A(n17361), .B(n17360), .Z(n17379) );
  XOR U18426 ( .A(a[720]), .B(n2279), .Z(n17383) );
  AND U18427 ( .A(a[722]), .B(b[0]), .Z(n17363) );
  XNOR U18428 ( .A(n17363), .B(n2175), .Z(n17365) );
  NANDN U18429 ( .A(b[0]), .B(a[721]), .Z(n17364) );
  NAND U18430 ( .A(n17365), .B(n17364), .Z(n17388) );
  AND U18431 ( .A(a[718]), .B(b[3]), .Z(n17387) );
  XOR U18432 ( .A(n17388), .B(n17387), .Z(n17390) );
  XOR U18433 ( .A(n17389), .B(n17390), .Z(n17378) );
  NANDN U18434 ( .A(n17367), .B(n17366), .Z(n17371) );
  OR U18435 ( .A(n17369), .B(n17368), .Z(n17370) );
  AND U18436 ( .A(n17371), .B(n17370), .Z(n17377) );
  XOR U18437 ( .A(n17378), .B(n17377), .Z(n17380) );
  XOR U18438 ( .A(n17379), .B(n17380), .Z(n17393) );
  XNOR U18439 ( .A(n17393), .B(sreg[1742]), .Z(n17395) );
  NANDN U18440 ( .A(n17372), .B(sreg[1741]), .Z(n17376) );
  NAND U18441 ( .A(n17374), .B(n17373), .Z(n17375) );
  NAND U18442 ( .A(n17376), .B(n17375), .Z(n17394) );
  XOR U18443 ( .A(n17395), .B(n17394), .Z(c[1742]) );
  NANDN U18444 ( .A(n17378), .B(n17377), .Z(n17382) );
  OR U18445 ( .A(n17380), .B(n17379), .Z(n17381) );
  AND U18446 ( .A(n17382), .B(n17381), .Z(n17400) );
  XOR U18447 ( .A(a[721]), .B(n2279), .Z(n17404) );
  AND U18448 ( .A(a[719]), .B(b[3]), .Z(n17408) );
  AND U18449 ( .A(a[723]), .B(b[0]), .Z(n17384) );
  XNOR U18450 ( .A(n17384), .B(n2175), .Z(n17386) );
  NANDN U18451 ( .A(b[0]), .B(a[722]), .Z(n17385) );
  NAND U18452 ( .A(n17386), .B(n17385), .Z(n17409) );
  XOR U18453 ( .A(n17408), .B(n17409), .Z(n17411) );
  XOR U18454 ( .A(n17410), .B(n17411), .Z(n17399) );
  NANDN U18455 ( .A(n17388), .B(n17387), .Z(n17392) );
  OR U18456 ( .A(n17390), .B(n17389), .Z(n17391) );
  AND U18457 ( .A(n17392), .B(n17391), .Z(n17398) );
  XOR U18458 ( .A(n17399), .B(n17398), .Z(n17401) );
  XOR U18459 ( .A(n17400), .B(n17401), .Z(n17414) );
  XNOR U18460 ( .A(n17414), .B(sreg[1743]), .Z(n17416) );
  NANDN U18461 ( .A(n17393), .B(sreg[1742]), .Z(n17397) );
  NAND U18462 ( .A(n17395), .B(n17394), .Z(n17396) );
  NAND U18463 ( .A(n17397), .B(n17396), .Z(n17415) );
  XOR U18464 ( .A(n17416), .B(n17415), .Z(c[1743]) );
  NANDN U18465 ( .A(n17399), .B(n17398), .Z(n17403) );
  OR U18466 ( .A(n17401), .B(n17400), .Z(n17402) );
  AND U18467 ( .A(n17403), .B(n17402), .Z(n17421) );
  XOR U18468 ( .A(a[722]), .B(n2279), .Z(n17425) );
  AND U18469 ( .A(a[720]), .B(b[3]), .Z(n17429) );
  AND U18470 ( .A(a[724]), .B(b[0]), .Z(n17405) );
  XNOR U18471 ( .A(n17405), .B(n2175), .Z(n17407) );
  NANDN U18472 ( .A(b[0]), .B(a[723]), .Z(n17406) );
  NAND U18473 ( .A(n17407), .B(n17406), .Z(n17430) );
  XOR U18474 ( .A(n17429), .B(n17430), .Z(n17432) );
  XOR U18475 ( .A(n17431), .B(n17432), .Z(n17420) );
  NANDN U18476 ( .A(n17409), .B(n17408), .Z(n17413) );
  OR U18477 ( .A(n17411), .B(n17410), .Z(n17412) );
  AND U18478 ( .A(n17413), .B(n17412), .Z(n17419) );
  XOR U18479 ( .A(n17420), .B(n17419), .Z(n17422) );
  XOR U18480 ( .A(n17421), .B(n17422), .Z(n17435) );
  XNOR U18481 ( .A(n17435), .B(sreg[1744]), .Z(n17437) );
  NANDN U18482 ( .A(n17414), .B(sreg[1743]), .Z(n17418) );
  NAND U18483 ( .A(n17416), .B(n17415), .Z(n17417) );
  NAND U18484 ( .A(n17418), .B(n17417), .Z(n17436) );
  XOR U18485 ( .A(n17437), .B(n17436), .Z(c[1744]) );
  NANDN U18486 ( .A(n17420), .B(n17419), .Z(n17424) );
  OR U18487 ( .A(n17422), .B(n17421), .Z(n17423) );
  AND U18488 ( .A(n17424), .B(n17423), .Z(n17442) );
  XOR U18489 ( .A(a[723]), .B(n2279), .Z(n17446) );
  AND U18490 ( .A(a[725]), .B(b[0]), .Z(n17426) );
  XNOR U18491 ( .A(n17426), .B(n2175), .Z(n17428) );
  NANDN U18492 ( .A(b[0]), .B(a[724]), .Z(n17427) );
  NAND U18493 ( .A(n17428), .B(n17427), .Z(n17451) );
  AND U18494 ( .A(a[721]), .B(b[3]), .Z(n17450) );
  XOR U18495 ( .A(n17451), .B(n17450), .Z(n17453) );
  XOR U18496 ( .A(n17452), .B(n17453), .Z(n17441) );
  NANDN U18497 ( .A(n17430), .B(n17429), .Z(n17434) );
  OR U18498 ( .A(n17432), .B(n17431), .Z(n17433) );
  AND U18499 ( .A(n17434), .B(n17433), .Z(n17440) );
  XOR U18500 ( .A(n17441), .B(n17440), .Z(n17443) );
  XOR U18501 ( .A(n17442), .B(n17443), .Z(n17456) );
  XNOR U18502 ( .A(n17456), .B(sreg[1745]), .Z(n17458) );
  NANDN U18503 ( .A(n17435), .B(sreg[1744]), .Z(n17439) );
  NAND U18504 ( .A(n17437), .B(n17436), .Z(n17438) );
  NAND U18505 ( .A(n17439), .B(n17438), .Z(n17457) );
  XOR U18506 ( .A(n17458), .B(n17457), .Z(c[1745]) );
  NANDN U18507 ( .A(n17441), .B(n17440), .Z(n17445) );
  OR U18508 ( .A(n17443), .B(n17442), .Z(n17444) );
  AND U18509 ( .A(n17445), .B(n17444), .Z(n17463) );
  XOR U18510 ( .A(a[724]), .B(n2279), .Z(n17467) );
  AND U18511 ( .A(a[722]), .B(b[3]), .Z(n17471) );
  AND U18512 ( .A(a[726]), .B(b[0]), .Z(n17447) );
  XNOR U18513 ( .A(n17447), .B(n2175), .Z(n17449) );
  NANDN U18514 ( .A(b[0]), .B(a[725]), .Z(n17448) );
  NAND U18515 ( .A(n17449), .B(n17448), .Z(n17472) );
  XOR U18516 ( .A(n17471), .B(n17472), .Z(n17474) );
  XOR U18517 ( .A(n17473), .B(n17474), .Z(n17462) );
  NANDN U18518 ( .A(n17451), .B(n17450), .Z(n17455) );
  OR U18519 ( .A(n17453), .B(n17452), .Z(n17454) );
  AND U18520 ( .A(n17455), .B(n17454), .Z(n17461) );
  XOR U18521 ( .A(n17462), .B(n17461), .Z(n17464) );
  XOR U18522 ( .A(n17463), .B(n17464), .Z(n17477) );
  XNOR U18523 ( .A(n17477), .B(sreg[1746]), .Z(n17479) );
  NANDN U18524 ( .A(n17456), .B(sreg[1745]), .Z(n17460) );
  NAND U18525 ( .A(n17458), .B(n17457), .Z(n17459) );
  NAND U18526 ( .A(n17460), .B(n17459), .Z(n17478) );
  XOR U18527 ( .A(n17479), .B(n17478), .Z(c[1746]) );
  NANDN U18528 ( .A(n17462), .B(n17461), .Z(n17466) );
  OR U18529 ( .A(n17464), .B(n17463), .Z(n17465) );
  AND U18530 ( .A(n17466), .B(n17465), .Z(n17484) );
  XOR U18531 ( .A(a[725]), .B(n2279), .Z(n17488) );
  AND U18532 ( .A(a[727]), .B(b[0]), .Z(n17468) );
  XNOR U18533 ( .A(n17468), .B(n2175), .Z(n17470) );
  NANDN U18534 ( .A(b[0]), .B(a[726]), .Z(n17469) );
  NAND U18535 ( .A(n17470), .B(n17469), .Z(n17493) );
  AND U18536 ( .A(a[723]), .B(b[3]), .Z(n17492) );
  XOR U18537 ( .A(n17493), .B(n17492), .Z(n17495) );
  XOR U18538 ( .A(n17494), .B(n17495), .Z(n17483) );
  NANDN U18539 ( .A(n17472), .B(n17471), .Z(n17476) );
  OR U18540 ( .A(n17474), .B(n17473), .Z(n17475) );
  AND U18541 ( .A(n17476), .B(n17475), .Z(n17482) );
  XOR U18542 ( .A(n17483), .B(n17482), .Z(n17485) );
  XOR U18543 ( .A(n17484), .B(n17485), .Z(n17498) );
  XNOR U18544 ( .A(n17498), .B(sreg[1747]), .Z(n17500) );
  NANDN U18545 ( .A(n17477), .B(sreg[1746]), .Z(n17481) );
  NAND U18546 ( .A(n17479), .B(n17478), .Z(n17480) );
  NAND U18547 ( .A(n17481), .B(n17480), .Z(n17499) );
  XOR U18548 ( .A(n17500), .B(n17499), .Z(c[1747]) );
  NANDN U18549 ( .A(n17483), .B(n17482), .Z(n17487) );
  OR U18550 ( .A(n17485), .B(n17484), .Z(n17486) );
  AND U18551 ( .A(n17487), .B(n17486), .Z(n17505) );
  XOR U18552 ( .A(a[726]), .B(n2279), .Z(n17509) );
  AND U18553 ( .A(a[728]), .B(b[0]), .Z(n17489) );
  XNOR U18554 ( .A(n17489), .B(n2175), .Z(n17491) );
  NANDN U18555 ( .A(b[0]), .B(a[727]), .Z(n17490) );
  NAND U18556 ( .A(n17491), .B(n17490), .Z(n17514) );
  AND U18557 ( .A(a[724]), .B(b[3]), .Z(n17513) );
  XOR U18558 ( .A(n17514), .B(n17513), .Z(n17516) );
  XOR U18559 ( .A(n17515), .B(n17516), .Z(n17504) );
  NANDN U18560 ( .A(n17493), .B(n17492), .Z(n17497) );
  OR U18561 ( .A(n17495), .B(n17494), .Z(n17496) );
  AND U18562 ( .A(n17497), .B(n17496), .Z(n17503) );
  XOR U18563 ( .A(n17504), .B(n17503), .Z(n17506) );
  XOR U18564 ( .A(n17505), .B(n17506), .Z(n17519) );
  XNOR U18565 ( .A(n17519), .B(sreg[1748]), .Z(n17521) );
  NANDN U18566 ( .A(n17498), .B(sreg[1747]), .Z(n17502) );
  NAND U18567 ( .A(n17500), .B(n17499), .Z(n17501) );
  NAND U18568 ( .A(n17502), .B(n17501), .Z(n17520) );
  XOR U18569 ( .A(n17521), .B(n17520), .Z(c[1748]) );
  NANDN U18570 ( .A(n17504), .B(n17503), .Z(n17508) );
  OR U18571 ( .A(n17506), .B(n17505), .Z(n17507) );
  AND U18572 ( .A(n17508), .B(n17507), .Z(n17526) );
  XOR U18573 ( .A(a[727]), .B(n2280), .Z(n17530) );
  AND U18574 ( .A(a[729]), .B(b[0]), .Z(n17510) );
  XNOR U18575 ( .A(n17510), .B(n2175), .Z(n17512) );
  NANDN U18576 ( .A(b[0]), .B(a[728]), .Z(n17511) );
  NAND U18577 ( .A(n17512), .B(n17511), .Z(n17535) );
  AND U18578 ( .A(a[725]), .B(b[3]), .Z(n17534) );
  XOR U18579 ( .A(n17535), .B(n17534), .Z(n17537) );
  XOR U18580 ( .A(n17536), .B(n17537), .Z(n17525) );
  NANDN U18581 ( .A(n17514), .B(n17513), .Z(n17518) );
  OR U18582 ( .A(n17516), .B(n17515), .Z(n17517) );
  AND U18583 ( .A(n17518), .B(n17517), .Z(n17524) );
  XOR U18584 ( .A(n17525), .B(n17524), .Z(n17527) );
  XOR U18585 ( .A(n17526), .B(n17527), .Z(n17540) );
  XNOR U18586 ( .A(n17540), .B(sreg[1749]), .Z(n17542) );
  NANDN U18587 ( .A(n17519), .B(sreg[1748]), .Z(n17523) );
  NAND U18588 ( .A(n17521), .B(n17520), .Z(n17522) );
  NAND U18589 ( .A(n17523), .B(n17522), .Z(n17541) );
  XOR U18590 ( .A(n17542), .B(n17541), .Z(c[1749]) );
  NANDN U18591 ( .A(n17525), .B(n17524), .Z(n17529) );
  OR U18592 ( .A(n17527), .B(n17526), .Z(n17528) );
  AND U18593 ( .A(n17529), .B(n17528), .Z(n17547) );
  XOR U18594 ( .A(a[728]), .B(n2280), .Z(n17551) );
  AND U18595 ( .A(a[730]), .B(b[0]), .Z(n17531) );
  XNOR U18596 ( .A(n17531), .B(n2175), .Z(n17533) );
  NANDN U18597 ( .A(b[0]), .B(a[729]), .Z(n17532) );
  NAND U18598 ( .A(n17533), .B(n17532), .Z(n17556) );
  AND U18599 ( .A(a[726]), .B(b[3]), .Z(n17555) );
  XOR U18600 ( .A(n17556), .B(n17555), .Z(n17558) );
  XOR U18601 ( .A(n17557), .B(n17558), .Z(n17546) );
  NANDN U18602 ( .A(n17535), .B(n17534), .Z(n17539) );
  OR U18603 ( .A(n17537), .B(n17536), .Z(n17538) );
  AND U18604 ( .A(n17539), .B(n17538), .Z(n17545) );
  XOR U18605 ( .A(n17546), .B(n17545), .Z(n17548) );
  XOR U18606 ( .A(n17547), .B(n17548), .Z(n17561) );
  XNOR U18607 ( .A(n17561), .B(sreg[1750]), .Z(n17563) );
  NANDN U18608 ( .A(n17540), .B(sreg[1749]), .Z(n17544) );
  NAND U18609 ( .A(n17542), .B(n17541), .Z(n17543) );
  NAND U18610 ( .A(n17544), .B(n17543), .Z(n17562) );
  XOR U18611 ( .A(n17563), .B(n17562), .Z(c[1750]) );
  NANDN U18612 ( .A(n17546), .B(n17545), .Z(n17550) );
  OR U18613 ( .A(n17548), .B(n17547), .Z(n17549) );
  AND U18614 ( .A(n17550), .B(n17549), .Z(n17568) );
  XOR U18615 ( .A(a[729]), .B(n2280), .Z(n17572) );
  AND U18616 ( .A(a[731]), .B(b[0]), .Z(n17552) );
  XNOR U18617 ( .A(n17552), .B(n2175), .Z(n17554) );
  NANDN U18618 ( .A(b[0]), .B(a[730]), .Z(n17553) );
  NAND U18619 ( .A(n17554), .B(n17553), .Z(n17577) );
  AND U18620 ( .A(a[727]), .B(b[3]), .Z(n17576) );
  XOR U18621 ( .A(n17577), .B(n17576), .Z(n17579) );
  XOR U18622 ( .A(n17578), .B(n17579), .Z(n17567) );
  NANDN U18623 ( .A(n17556), .B(n17555), .Z(n17560) );
  OR U18624 ( .A(n17558), .B(n17557), .Z(n17559) );
  AND U18625 ( .A(n17560), .B(n17559), .Z(n17566) );
  XOR U18626 ( .A(n17567), .B(n17566), .Z(n17569) );
  XOR U18627 ( .A(n17568), .B(n17569), .Z(n17582) );
  XNOR U18628 ( .A(n17582), .B(sreg[1751]), .Z(n17584) );
  NANDN U18629 ( .A(n17561), .B(sreg[1750]), .Z(n17565) );
  NAND U18630 ( .A(n17563), .B(n17562), .Z(n17564) );
  NAND U18631 ( .A(n17565), .B(n17564), .Z(n17583) );
  XOR U18632 ( .A(n17584), .B(n17583), .Z(c[1751]) );
  NANDN U18633 ( .A(n17567), .B(n17566), .Z(n17571) );
  OR U18634 ( .A(n17569), .B(n17568), .Z(n17570) );
  AND U18635 ( .A(n17571), .B(n17570), .Z(n17589) );
  XOR U18636 ( .A(a[730]), .B(n2280), .Z(n17593) );
  AND U18637 ( .A(a[728]), .B(b[3]), .Z(n17597) );
  AND U18638 ( .A(a[732]), .B(b[0]), .Z(n17573) );
  XNOR U18639 ( .A(n17573), .B(n2175), .Z(n17575) );
  NANDN U18640 ( .A(b[0]), .B(a[731]), .Z(n17574) );
  NAND U18641 ( .A(n17575), .B(n17574), .Z(n17598) );
  XOR U18642 ( .A(n17597), .B(n17598), .Z(n17600) );
  XOR U18643 ( .A(n17599), .B(n17600), .Z(n17588) );
  NANDN U18644 ( .A(n17577), .B(n17576), .Z(n17581) );
  OR U18645 ( .A(n17579), .B(n17578), .Z(n17580) );
  AND U18646 ( .A(n17581), .B(n17580), .Z(n17587) );
  XOR U18647 ( .A(n17588), .B(n17587), .Z(n17590) );
  XOR U18648 ( .A(n17589), .B(n17590), .Z(n17603) );
  XNOR U18649 ( .A(n17603), .B(sreg[1752]), .Z(n17605) );
  NANDN U18650 ( .A(n17582), .B(sreg[1751]), .Z(n17586) );
  NAND U18651 ( .A(n17584), .B(n17583), .Z(n17585) );
  NAND U18652 ( .A(n17586), .B(n17585), .Z(n17604) );
  XOR U18653 ( .A(n17605), .B(n17604), .Z(c[1752]) );
  NANDN U18654 ( .A(n17588), .B(n17587), .Z(n17592) );
  OR U18655 ( .A(n17590), .B(n17589), .Z(n17591) );
  AND U18656 ( .A(n17592), .B(n17591), .Z(n17610) );
  XOR U18657 ( .A(a[731]), .B(n2280), .Z(n17614) );
  AND U18658 ( .A(a[733]), .B(b[0]), .Z(n17594) );
  XNOR U18659 ( .A(n17594), .B(n2175), .Z(n17596) );
  NANDN U18660 ( .A(b[0]), .B(a[732]), .Z(n17595) );
  NAND U18661 ( .A(n17596), .B(n17595), .Z(n17619) );
  AND U18662 ( .A(a[729]), .B(b[3]), .Z(n17618) );
  XOR U18663 ( .A(n17619), .B(n17618), .Z(n17621) );
  XOR U18664 ( .A(n17620), .B(n17621), .Z(n17609) );
  NANDN U18665 ( .A(n17598), .B(n17597), .Z(n17602) );
  OR U18666 ( .A(n17600), .B(n17599), .Z(n17601) );
  AND U18667 ( .A(n17602), .B(n17601), .Z(n17608) );
  XOR U18668 ( .A(n17609), .B(n17608), .Z(n17611) );
  XOR U18669 ( .A(n17610), .B(n17611), .Z(n17624) );
  XNOR U18670 ( .A(n17624), .B(sreg[1753]), .Z(n17626) );
  NANDN U18671 ( .A(n17603), .B(sreg[1752]), .Z(n17607) );
  NAND U18672 ( .A(n17605), .B(n17604), .Z(n17606) );
  NAND U18673 ( .A(n17607), .B(n17606), .Z(n17625) );
  XOR U18674 ( .A(n17626), .B(n17625), .Z(c[1753]) );
  NANDN U18675 ( .A(n17609), .B(n17608), .Z(n17613) );
  OR U18676 ( .A(n17611), .B(n17610), .Z(n17612) );
  AND U18677 ( .A(n17613), .B(n17612), .Z(n17631) );
  XOR U18678 ( .A(a[732]), .B(n2280), .Z(n17635) );
  AND U18679 ( .A(a[734]), .B(b[0]), .Z(n17615) );
  XNOR U18680 ( .A(n17615), .B(n2175), .Z(n17617) );
  NANDN U18681 ( .A(b[0]), .B(a[733]), .Z(n17616) );
  NAND U18682 ( .A(n17617), .B(n17616), .Z(n17640) );
  AND U18683 ( .A(a[730]), .B(b[3]), .Z(n17639) );
  XOR U18684 ( .A(n17640), .B(n17639), .Z(n17642) );
  XOR U18685 ( .A(n17641), .B(n17642), .Z(n17630) );
  NANDN U18686 ( .A(n17619), .B(n17618), .Z(n17623) );
  OR U18687 ( .A(n17621), .B(n17620), .Z(n17622) );
  AND U18688 ( .A(n17623), .B(n17622), .Z(n17629) );
  XOR U18689 ( .A(n17630), .B(n17629), .Z(n17632) );
  XOR U18690 ( .A(n17631), .B(n17632), .Z(n17645) );
  XNOR U18691 ( .A(n17645), .B(sreg[1754]), .Z(n17647) );
  NANDN U18692 ( .A(n17624), .B(sreg[1753]), .Z(n17628) );
  NAND U18693 ( .A(n17626), .B(n17625), .Z(n17627) );
  NAND U18694 ( .A(n17628), .B(n17627), .Z(n17646) );
  XOR U18695 ( .A(n17647), .B(n17646), .Z(c[1754]) );
  NANDN U18696 ( .A(n17630), .B(n17629), .Z(n17634) );
  OR U18697 ( .A(n17632), .B(n17631), .Z(n17633) );
  AND U18698 ( .A(n17634), .B(n17633), .Z(n17652) );
  XOR U18699 ( .A(a[733]), .B(n2280), .Z(n17656) );
  AND U18700 ( .A(a[731]), .B(b[3]), .Z(n17660) );
  AND U18701 ( .A(a[735]), .B(b[0]), .Z(n17636) );
  XNOR U18702 ( .A(n17636), .B(n2175), .Z(n17638) );
  NANDN U18703 ( .A(b[0]), .B(a[734]), .Z(n17637) );
  NAND U18704 ( .A(n17638), .B(n17637), .Z(n17661) );
  XOR U18705 ( .A(n17660), .B(n17661), .Z(n17663) );
  XOR U18706 ( .A(n17662), .B(n17663), .Z(n17651) );
  NANDN U18707 ( .A(n17640), .B(n17639), .Z(n17644) );
  OR U18708 ( .A(n17642), .B(n17641), .Z(n17643) );
  AND U18709 ( .A(n17644), .B(n17643), .Z(n17650) );
  XOR U18710 ( .A(n17651), .B(n17650), .Z(n17653) );
  XOR U18711 ( .A(n17652), .B(n17653), .Z(n17666) );
  XNOR U18712 ( .A(n17666), .B(sreg[1755]), .Z(n17668) );
  NANDN U18713 ( .A(n17645), .B(sreg[1754]), .Z(n17649) );
  NAND U18714 ( .A(n17647), .B(n17646), .Z(n17648) );
  NAND U18715 ( .A(n17649), .B(n17648), .Z(n17667) );
  XOR U18716 ( .A(n17668), .B(n17667), .Z(c[1755]) );
  NANDN U18717 ( .A(n17651), .B(n17650), .Z(n17655) );
  OR U18718 ( .A(n17653), .B(n17652), .Z(n17654) );
  AND U18719 ( .A(n17655), .B(n17654), .Z(n17673) );
  XOR U18720 ( .A(a[734]), .B(n2281), .Z(n17677) );
  AND U18721 ( .A(a[736]), .B(b[0]), .Z(n17657) );
  XNOR U18722 ( .A(n17657), .B(n2175), .Z(n17659) );
  NANDN U18723 ( .A(b[0]), .B(a[735]), .Z(n17658) );
  NAND U18724 ( .A(n17659), .B(n17658), .Z(n17682) );
  AND U18725 ( .A(a[732]), .B(b[3]), .Z(n17681) );
  XOR U18726 ( .A(n17682), .B(n17681), .Z(n17684) );
  XOR U18727 ( .A(n17683), .B(n17684), .Z(n17672) );
  NANDN U18728 ( .A(n17661), .B(n17660), .Z(n17665) );
  OR U18729 ( .A(n17663), .B(n17662), .Z(n17664) );
  AND U18730 ( .A(n17665), .B(n17664), .Z(n17671) );
  XOR U18731 ( .A(n17672), .B(n17671), .Z(n17674) );
  XOR U18732 ( .A(n17673), .B(n17674), .Z(n17687) );
  XNOR U18733 ( .A(n17687), .B(sreg[1756]), .Z(n17689) );
  NANDN U18734 ( .A(n17666), .B(sreg[1755]), .Z(n17670) );
  NAND U18735 ( .A(n17668), .B(n17667), .Z(n17669) );
  NAND U18736 ( .A(n17670), .B(n17669), .Z(n17688) );
  XOR U18737 ( .A(n17689), .B(n17688), .Z(c[1756]) );
  NANDN U18738 ( .A(n17672), .B(n17671), .Z(n17676) );
  OR U18739 ( .A(n17674), .B(n17673), .Z(n17675) );
  AND U18740 ( .A(n17676), .B(n17675), .Z(n17694) );
  XOR U18741 ( .A(a[735]), .B(n2281), .Z(n17698) );
  AND U18742 ( .A(a[737]), .B(b[0]), .Z(n17678) );
  XNOR U18743 ( .A(n17678), .B(n2175), .Z(n17680) );
  NANDN U18744 ( .A(b[0]), .B(a[736]), .Z(n17679) );
  NAND U18745 ( .A(n17680), .B(n17679), .Z(n17703) );
  AND U18746 ( .A(a[733]), .B(b[3]), .Z(n17702) );
  XOR U18747 ( .A(n17703), .B(n17702), .Z(n17705) );
  XOR U18748 ( .A(n17704), .B(n17705), .Z(n17693) );
  NANDN U18749 ( .A(n17682), .B(n17681), .Z(n17686) );
  OR U18750 ( .A(n17684), .B(n17683), .Z(n17685) );
  AND U18751 ( .A(n17686), .B(n17685), .Z(n17692) );
  XOR U18752 ( .A(n17693), .B(n17692), .Z(n17695) );
  XOR U18753 ( .A(n17694), .B(n17695), .Z(n17708) );
  XNOR U18754 ( .A(n17708), .B(sreg[1757]), .Z(n17710) );
  NANDN U18755 ( .A(n17687), .B(sreg[1756]), .Z(n17691) );
  NAND U18756 ( .A(n17689), .B(n17688), .Z(n17690) );
  NAND U18757 ( .A(n17691), .B(n17690), .Z(n17709) );
  XOR U18758 ( .A(n17710), .B(n17709), .Z(c[1757]) );
  NANDN U18759 ( .A(n17693), .B(n17692), .Z(n17697) );
  OR U18760 ( .A(n17695), .B(n17694), .Z(n17696) );
  AND U18761 ( .A(n17697), .B(n17696), .Z(n17715) );
  XOR U18762 ( .A(a[736]), .B(n2281), .Z(n17719) );
  AND U18763 ( .A(a[734]), .B(b[3]), .Z(n17723) );
  AND U18764 ( .A(a[738]), .B(b[0]), .Z(n17699) );
  XNOR U18765 ( .A(n17699), .B(n2175), .Z(n17701) );
  NANDN U18766 ( .A(b[0]), .B(a[737]), .Z(n17700) );
  NAND U18767 ( .A(n17701), .B(n17700), .Z(n17724) );
  XOR U18768 ( .A(n17723), .B(n17724), .Z(n17726) );
  XOR U18769 ( .A(n17725), .B(n17726), .Z(n17714) );
  NANDN U18770 ( .A(n17703), .B(n17702), .Z(n17707) );
  OR U18771 ( .A(n17705), .B(n17704), .Z(n17706) );
  AND U18772 ( .A(n17707), .B(n17706), .Z(n17713) );
  XOR U18773 ( .A(n17714), .B(n17713), .Z(n17716) );
  XOR U18774 ( .A(n17715), .B(n17716), .Z(n17729) );
  XNOR U18775 ( .A(n17729), .B(sreg[1758]), .Z(n17731) );
  NANDN U18776 ( .A(n17708), .B(sreg[1757]), .Z(n17712) );
  NAND U18777 ( .A(n17710), .B(n17709), .Z(n17711) );
  NAND U18778 ( .A(n17712), .B(n17711), .Z(n17730) );
  XOR U18779 ( .A(n17731), .B(n17730), .Z(c[1758]) );
  NANDN U18780 ( .A(n17714), .B(n17713), .Z(n17718) );
  OR U18781 ( .A(n17716), .B(n17715), .Z(n17717) );
  AND U18782 ( .A(n17718), .B(n17717), .Z(n17737) );
  XOR U18783 ( .A(a[737]), .B(n2281), .Z(n17738) );
  AND U18784 ( .A(b[0]), .B(a[739]), .Z(n17720) );
  XOR U18785 ( .A(b[1]), .B(n17720), .Z(n17722) );
  NANDN U18786 ( .A(b[0]), .B(a[738]), .Z(n17721) );
  AND U18787 ( .A(n17722), .B(n17721), .Z(n17742) );
  AND U18788 ( .A(a[735]), .B(b[3]), .Z(n17743) );
  XOR U18789 ( .A(n17742), .B(n17743), .Z(n17744) );
  XNOR U18790 ( .A(n17745), .B(n17744), .Z(n17734) );
  NANDN U18791 ( .A(n17724), .B(n17723), .Z(n17728) );
  OR U18792 ( .A(n17726), .B(n17725), .Z(n17727) );
  AND U18793 ( .A(n17728), .B(n17727), .Z(n17735) );
  XNOR U18794 ( .A(n17734), .B(n17735), .Z(n17736) );
  XNOR U18795 ( .A(n17737), .B(n17736), .Z(n17748) );
  XNOR U18796 ( .A(n17748), .B(sreg[1759]), .Z(n17750) );
  NANDN U18797 ( .A(n17729), .B(sreg[1758]), .Z(n17733) );
  NAND U18798 ( .A(n17731), .B(n17730), .Z(n17732) );
  NAND U18799 ( .A(n17733), .B(n17732), .Z(n17749) );
  XOR U18800 ( .A(n17750), .B(n17749), .Z(c[1759]) );
  XOR U18801 ( .A(a[738]), .B(n2281), .Z(n17757) );
  AND U18802 ( .A(a[740]), .B(b[0]), .Z(n17739) );
  XNOR U18803 ( .A(n17739), .B(n2175), .Z(n17741) );
  NANDN U18804 ( .A(b[0]), .B(a[739]), .Z(n17740) );
  NAND U18805 ( .A(n17741), .B(n17740), .Z(n17762) );
  AND U18806 ( .A(a[736]), .B(b[3]), .Z(n17761) );
  XOR U18807 ( .A(n17762), .B(n17761), .Z(n17764) );
  XOR U18808 ( .A(n17763), .B(n17764), .Z(n17752) );
  NAND U18809 ( .A(n17743), .B(n17742), .Z(n17747) );
  NANDN U18810 ( .A(n17745), .B(n17744), .Z(n17746) );
  AND U18811 ( .A(n17747), .B(n17746), .Z(n17751) );
  XOR U18812 ( .A(n17752), .B(n17751), .Z(n17754) );
  XOR U18813 ( .A(n17753), .B(n17754), .Z(n17767) );
  XNOR U18814 ( .A(n17767), .B(sreg[1760]), .Z(n17769) );
  XOR U18815 ( .A(n17769), .B(n17768), .Z(c[1760]) );
  NANDN U18816 ( .A(n17752), .B(n17751), .Z(n17756) );
  OR U18817 ( .A(n17754), .B(n17753), .Z(n17755) );
  AND U18818 ( .A(n17756), .B(n17755), .Z(n17775) );
  XOR U18819 ( .A(a[739]), .B(n2281), .Z(n17776) );
  AND U18820 ( .A(b[0]), .B(a[741]), .Z(n17758) );
  XOR U18821 ( .A(b[1]), .B(n17758), .Z(n17760) );
  NANDN U18822 ( .A(b[0]), .B(a[740]), .Z(n17759) );
  AND U18823 ( .A(n17760), .B(n17759), .Z(n17780) );
  AND U18824 ( .A(a[737]), .B(b[3]), .Z(n17781) );
  XOR U18825 ( .A(n17780), .B(n17781), .Z(n17782) );
  XNOR U18826 ( .A(n17783), .B(n17782), .Z(n17772) );
  NANDN U18827 ( .A(n17762), .B(n17761), .Z(n17766) );
  OR U18828 ( .A(n17764), .B(n17763), .Z(n17765) );
  AND U18829 ( .A(n17766), .B(n17765), .Z(n17773) );
  XNOR U18830 ( .A(n17772), .B(n17773), .Z(n17774) );
  XNOR U18831 ( .A(n17775), .B(n17774), .Z(n17786) );
  XNOR U18832 ( .A(n17786), .B(sreg[1761]), .Z(n17788) );
  NANDN U18833 ( .A(n17767), .B(sreg[1760]), .Z(n17771) );
  NAND U18834 ( .A(n17769), .B(n17768), .Z(n17770) );
  NAND U18835 ( .A(n17771), .B(n17770), .Z(n17787) );
  XOR U18836 ( .A(n17788), .B(n17787), .Z(c[1761]) );
  XOR U18837 ( .A(a[740]), .B(n2281), .Z(n17795) );
  AND U18838 ( .A(a[742]), .B(b[0]), .Z(n17777) );
  XNOR U18839 ( .A(n17777), .B(n2175), .Z(n17779) );
  NANDN U18840 ( .A(b[0]), .B(a[741]), .Z(n17778) );
  NAND U18841 ( .A(n17779), .B(n17778), .Z(n17800) );
  AND U18842 ( .A(a[738]), .B(b[3]), .Z(n17799) );
  XOR U18843 ( .A(n17800), .B(n17799), .Z(n17802) );
  XOR U18844 ( .A(n17801), .B(n17802), .Z(n17790) );
  NAND U18845 ( .A(n17781), .B(n17780), .Z(n17785) );
  NANDN U18846 ( .A(n17783), .B(n17782), .Z(n17784) );
  AND U18847 ( .A(n17785), .B(n17784), .Z(n17789) );
  XOR U18848 ( .A(n17790), .B(n17789), .Z(n17792) );
  XOR U18849 ( .A(n17791), .B(n17792), .Z(n17805) );
  XNOR U18850 ( .A(n17805), .B(sreg[1762]), .Z(n17807) );
  XOR U18851 ( .A(n17807), .B(n17806), .Z(c[1762]) );
  NANDN U18852 ( .A(n17790), .B(n17789), .Z(n17794) );
  OR U18853 ( .A(n17792), .B(n17791), .Z(n17793) );
  AND U18854 ( .A(n17794), .B(n17793), .Z(n17812) );
  XOR U18855 ( .A(a[741]), .B(n2282), .Z(n17816) );
  AND U18856 ( .A(a[743]), .B(b[0]), .Z(n17796) );
  XNOR U18857 ( .A(n17796), .B(n2175), .Z(n17798) );
  NANDN U18858 ( .A(b[0]), .B(a[742]), .Z(n17797) );
  NAND U18859 ( .A(n17798), .B(n17797), .Z(n17821) );
  AND U18860 ( .A(a[739]), .B(b[3]), .Z(n17820) );
  XOR U18861 ( .A(n17821), .B(n17820), .Z(n17823) );
  XOR U18862 ( .A(n17822), .B(n17823), .Z(n17811) );
  NANDN U18863 ( .A(n17800), .B(n17799), .Z(n17804) );
  OR U18864 ( .A(n17802), .B(n17801), .Z(n17803) );
  AND U18865 ( .A(n17804), .B(n17803), .Z(n17810) );
  XOR U18866 ( .A(n17811), .B(n17810), .Z(n17813) );
  XOR U18867 ( .A(n17812), .B(n17813), .Z(n17826) );
  XNOR U18868 ( .A(n17826), .B(sreg[1763]), .Z(n17828) );
  NANDN U18869 ( .A(n17805), .B(sreg[1762]), .Z(n17809) );
  NAND U18870 ( .A(n17807), .B(n17806), .Z(n17808) );
  NAND U18871 ( .A(n17809), .B(n17808), .Z(n17827) );
  XOR U18872 ( .A(n17828), .B(n17827), .Z(c[1763]) );
  NANDN U18873 ( .A(n17811), .B(n17810), .Z(n17815) );
  OR U18874 ( .A(n17813), .B(n17812), .Z(n17814) );
  AND U18875 ( .A(n17815), .B(n17814), .Z(n17833) );
  XOR U18876 ( .A(a[742]), .B(n2282), .Z(n17837) );
  AND U18877 ( .A(a[744]), .B(b[0]), .Z(n17817) );
  XNOR U18878 ( .A(n17817), .B(n2175), .Z(n17819) );
  NANDN U18879 ( .A(b[0]), .B(a[743]), .Z(n17818) );
  NAND U18880 ( .A(n17819), .B(n17818), .Z(n17842) );
  AND U18881 ( .A(a[740]), .B(b[3]), .Z(n17841) );
  XOR U18882 ( .A(n17842), .B(n17841), .Z(n17844) );
  XOR U18883 ( .A(n17843), .B(n17844), .Z(n17832) );
  NANDN U18884 ( .A(n17821), .B(n17820), .Z(n17825) );
  OR U18885 ( .A(n17823), .B(n17822), .Z(n17824) );
  AND U18886 ( .A(n17825), .B(n17824), .Z(n17831) );
  XOR U18887 ( .A(n17832), .B(n17831), .Z(n17834) );
  XOR U18888 ( .A(n17833), .B(n17834), .Z(n17847) );
  XNOR U18889 ( .A(n17847), .B(sreg[1764]), .Z(n17849) );
  NANDN U18890 ( .A(n17826), .B(sreg[1763]), .Z(n17830) );
  NAND U18891 ( .A(n17828), .B(n17827), .Z(n17829) );
  NAND U18892 ( .A(n17830), .B(n17829), .Z(n17848) );
  XOR U18893 ( .A(n17849), .B(n17848), .Z(c[1764]) );
  NANDN U18894 ( .A(n17832), .B(n17831), .Z(n17836) );
  OR U18895 ( .A(n17834), .B(n17833), .Z(n17835) );
  AND U18896 ( .A(n17836), .B(n17835), .Z(n17854) );
  XOR U18897 ( .A(a[743]), .B(n2282), .Z(n17858) );
  AND U18898 ( .A(a[745]), .B(b[0]), .Z(n17838) );
  XNOR U18899 ( .A(n17838), .B(n2175), .Z(n17840) );
  NANDN U18900 ( .A(b[0]), .B(a[744]), .Z(n17839) );
  NAND U18901 ( .A(n17840), .B(n17839), .Z(n17863) );
  AND U18902 ( .A(a[741]), .B(b[3]), .Z(n17862) );
  XOR U18903 ( .A(n17863), .B(n17862), .Z(n17865) );
  XOR U18904 ( .A(n17864), .B(n17865), .Z(n17853) );
  NANDN U18905 ( .A(n17842), .B(n17841), .Z(n17846) );
  OR U18906 ( .A(n17844), .B(n17843), .Z(n17845) );
  AND U18907 ( .A(n17846), .B(n17845), .Z(n17852) );
  XOR U18908 ( .A(n17853), .B(n17852), .Z(n17855) );
  XOR U18909 ( .A(n17854), .B(n17855), .Z(n17868) );
  XNOR U18910 ( .A(n17868), .B(sreg[1765]), .Z(n17870) );
  NANDN U18911 ( .A(n17847), .B(sreg[1764]), .Z(n17851) );
  NAND U18912 ( .A(n17849), .B(n17848), .Z(n17850) );
  NAND U18913 ( .A(n17851), .B(n17850), .Z(n17869) );
  XOR U18914 ( .A(n17870), .B(n17869), .Z(c[1765]) );
  NANDN U18915 ( .A(n17853), .B(n17852), .Z(n17857) );
  OR U18916 ( .A(n17855), .B(n17854), .Z(n17856) );
  AND U18917 ( .A(n17857), .B(n17856), .Z(n17875) );
  XOR U18918 ( .A(a[744]), .B(n2282), .Z(n17879) );
  AND U18919 ( .A(a[742]), .B(b[3]), .Z(n17883) );
  AND U18920 ( .A(a[746]), .B(b[0]), .Z(n17859) );
  XNOR U18921 ( .A(n17859), .B(n2175), .Z(n17861) );
  NANDN U18922 ( .A(b[0]), .B(a[745]), .Z(n17860) );
  NAND U18923 ( .A(n17861), .B(n17860), .Z(n17884) );
  XOR U18924 ( .A(n17883), .B(n17884), .Z(n17886) );
  XOR U18925 ( .A(n17885), .B(n17886), .Z(n17874) );
  NANDN U18926 ( .A(n17863), .B(n17862), .Z(n17867) );
  OR U18927 ( .A(n17865), .B(n17864), .Z(n17866) );
  AND U18928 ( .A(n17867), .B(n17866), .Z(n17873) );
  XOR U18929 ( .A(n17874), .B(n17873), .Z(n17876) );
  XOR U18930 ( .A(n17875), .B(n17876), .Z(n17889) );
  XNOR U18931 ( .A(n17889), .B(sreg[1766]), .Z(n17891) );
  NANDN U18932 ( .A(n17868), .B(sreg[1765]), .Z(n17872) );
  NAND U18933 ( .A(n17870), .B(n17869), .Z(n17871) );
  NAND U18934 ( .A(n17872), .B(n17871), .Z(n17890) );
  XOR U18935 ( .A(n17891), .B(n17890), .Z(c[1766]) );
  NANDN U18936 ( .A(n17874), .B(n17873), .Z(n17878) );
  OR U18937 ( .A(n17876), .B(n17875), .Z(n17877) );
  AND U18938 ( .A(n17878), .B(n17877), .Z(n17896) );
  XOR U18939 ( .A(a[745]), .B(n2282), .Z(n17900) );
  AND U18940 ( .A(a[743]), .B(b[3]), .Z(n17904) );
  AND U18941 ( .A(a[747]), .B(b[0]), .Z(n17880) );
  XNOR U18942 ( .A(n17880), .B(n2175), .Z(n17882) );
  NANDN U18943 ( .A(b[0]), .B(a[746]), .Z(n17881) );
  NAND U18944 ( .A(n17882), .B(n17881), .Z(n17905) );
  XOR U18945 ( .A(n17904), .B(n17905), .Z(n17907) );
  XOR U18946 ( .A(n17906), .B(n17907), .Z(n17895) );
  NANDN U18947 ( .A(n17884), .B(n17883), .Z(n17888) );
  OR U18948 ( .A(n17886), .B(n17885), .Z(n17887) );
  AND U18949 ( .A(n17888), .B(n17887), .Z(n17894) );
  XOR U18950 ( .A(n17895), .B(n17894), .Z(n17897) );
  XOR U18951 ( .A(n17896), .B(n17897), .Z(n17910) );
  XNOR U18952 ( .A(n17910), .B(sreg[1767]), .Z(n17912) );
  NANDN U18953 ( .A(n17889), .B(sreg[1766]), .Z(n17893) );
  NAND U18954 ( .A(n17891), .B(n17890), .Z(n17892) );
  NAND U18955 ( .A(n17893), .B(n17892), .Z(n17911) );
  XOR U18956 ( .A(n17912), .B(n17911), .Z(c[1767]) );
  NANDN U18957 ( .A(n17895), .B(n17894), .Z(n17899) );
  OR U18958 ( .A(n17897), .B(n17896), .Z(n17898) );
  AND U18959 ( .A(n17899), .B(n17898), .Z(n17917) );
  XOR U18960 ( .A(a[746]), .B(n2282), .Z(n17921) );
  AND U18961 ( .A(a[748]), .B(b[0]), .Z(n17901) );
  XNOR U18962 ( .A(n17901), .B(n2175), .Z(n17903) );
  NANDN U18963 ( .A(b[0]), .B(a[747]), .Z(n17902) );
  NAND U18964 ( .A(n17903), .B(n17902), .Z(n17926) );
  AND U18965 ( .A(a[744]), .B(b[3]), .Z(n17925) );
  XOR U18966 ( .A(n17926), .B(n17925), .Z(n17928) );
  XOR U18967 ( .A(n17927), .B(n17928), .Z(n17916) );
  NANDN U18968 ( .A(n17905), .B(n17904), .Z(n17909) );
  OR U18969 ( .A(n17907), .B(n17906), .Z(n17908) );
  AND U18970 ( .A(n17909), .B(n17908), .Z(n17915) );
  XOR U18971 ( .A(n17916), .B(n17915), .Z(n17918) );
  XOR U18972 ( .A(n17917), .B(n17918), .Z(n17931) );
  XNOR U18973 ( .A(n17931), .B(sreg[1768]), .Z(n17933) );
  NANDN U18974 ( .A(n17910), .B(sreg[1767]), .Z(n17914) );
  NAND U18975 ( .A(n17912), .B(n17911), .Z(n17913) );
  NAND U18976 ( .A(n17914), .B(n17913), .Z(n17932) );
  XOR U18977 ( .A(n17933), .B(n17932), .Z(c[1768]) );
  NANDN U18978 ( .A(n17916), .B(n17915), .Z(n17920) );
  OR U18979 ( .A(n17918), .B(n17917), .Z(n17919) );
  AND U18980 ( .A(n17920), .B(n17919), .Z(n17938) );
  XOR U18981 ( .A(a[747]), .B(n2282), .Z(n17942) );
  AND U18982 ( .A(a[745]), .B(b[3]), .Z(n17946) );
  AND U18983 ( .A(a[749]), .B(b[0]), .Z(n17922) );
  XNOR U18984 ( .A(n17922), .B(n2175), .Z(n17924) );
  NANDN U18985 ( .A(b[0]), .B(a[748]), .Z(n17923) );
  NAND U18986 ( .A(n17924), .B(n17923), .Z(n17947) );
  XOR U18987 ( .A(n17946), .B(n17947), .Z(n17949) );
  XOR U18988 ( .A(n17948), .B(n17949), .Z(n17937) );
  NANDN U18989 ( .A(n17926), .B(n17925), .Z(n17930) );
  OR U18990 ( .A(n17928), .B(n17927), .Z(n17929) );
  AND U18991 ( .A(n17930), .B(n17929), .Z(n17936) );
  XOR U18992 ( .A(n17937), .B(n17936), .Z(n17939) );
  XOR U18993 ( .A(n17938), .B(n17939), .Z(n17952) );
  XNOR U18994 ( .A(n17952), .B(sreg[1769]), .Z(n17954) );
  NANDN U18995 ( .A(n17931), .B(sreg[1768]), .Z(n17935) );
  NAND U18996 ( .A(n17933), .B(n17932), .Z(n17934) );
  NAND U18997 ( .A(n17935), .B(n17934), .Z(n17953) );
  XOR U18998 ( .A(n17954), .B(n17953), .Z(c[1769]) );
  NANDN U18999 ( .A(n17937), .B(n17936), .Z(n17941) );
  OR U19000 ( .A(n17939), .B(n17938), .Z(n17940) );
  AND U19001 ( .A(n17941), .B(n17940), .Z(n17959) );
  XOR U19002 ( .A(a[748]), .B(n2283), .Z(n17963) );
  AND U19003 ( .A(a[750]), .B(b[0]), .Z(n17943) );
  XNOR U19004 ( .A(n17943), .B(n2175), .Z(n17945) );
  NANDN U19005 ( .A(b[0]), .B(a[749]), .Z(n17944) );
  NAND U19006 ( .A(n17945), .B(n17944), .Z(n17968) );
  AND U19007 ( .A(a[746]), .B(b[3]), .Z(n17967) );
  XOR U19008 ( .A(n17968), .B(n17967), .Z(n17970) );
  XOR U19009 ( .A(n17969), .B(n17970), .Z(n17958) );
  NANDN U19010 ( .A(n17947), .B(n17946), .Z(n17951) );
  OR U19011 ( .A(n17949), .B(n17948), .Z(n17950) );
  AND U19012 ( .A(n17951), .B(n17950), .Z(n17957) );
  XOR U19013 ( .A(n17958), .B(n17957), .Z(n17960) );
  XOR U19014 ( .A(n17959), .B(n17960), .Z(n17973) );
  XNOR U19015 ( .A(n17973), .B(sreg[1770]), .Z(n17975) );
  NANDN U19016 ( .A(n17952), .B(sreg[1769]), .Z(n17956) );
  NAND U19017 ( .A(n17954), .B(n17953), .Z(n17955) );
  NAND U19018 ( .A(n17956), .B(n17955), .Z(n17974) );
  XOR U19019 ( .A(n17975), .B(n17974), .Z(c[1770]) );
  NANDN U19020 ( .A(n17958), .B(n17957), .Z(n17962) );
  OR U19021 ( .A(n17960), .B(n17959), .Z(n17961) );
  AND U19022 ( .A(n17962), .B(n17961), .Z(n17980) );
  XOR U19023 ( .A(a[749]), .B(n2283), .Z(n17984) );
  AND U19024 ( .A(a[751]), .B(b[0]), .Z(n17964) );
  XNOR U19025 ( .A(n17964), .B(n2175), .Z(n17966) );
  NANDN U19026 ( .A(b[0]), .B(a[750]), .Z(n17965) );
  NAND U19027 ( .A(n17966), .B(n17965), .Z(n17989) );
  AND U19028 ( .A(a[747]), .B(b[3]), .Z(n17988) );
  XOR U19029 ( .A(n17989), .B(n17988), .Z(n17991) );
  XOR U19030 ( .A(n17990), .B(n17991), .Z(n17979) );
  NANDN U19031 ( .A(n17968), .B(n17967), .Z(n17972) );
  OR U19032 ( .A(n17970), .B(n17969), .Z(n17971) );
  AND U19033 ( .A(n17972), .B(n17971), .Z(n17978) );
  XOR U19034 ( .A(n17979), .B(n17978), .Z(n17981) );
  XOR U19035 ( .A(n17980), .B(n17981), .Z(n17994) );
  XNOR U19036 ( .A(n17994), .B(sreg[1771]), .Z(n17996) );
  NANDN U19037 ( .A(n17973), .B(sreg[1770]), .Z(n17977) );
  NAND U19038 ( .A(n17975), .B(n17974), .Z(n17976) );
  NAND U19039 ( .A(n17977), .B(n17976), .Z(n17995) );
  XOR U19040 ( .A(n17996), .B(n17995), .Z(c[1771]) );
  NANDN U19041 ( .A(n17979), .B(n17978), .Z(n17983) );
  OR U19042 ( .A(n17981), .B(n17980), .Z(n17982) );
  AND U19043 ( .A(n17983), .B(n17982), .Z(n18001) );
  XOR U19044 ( .A(a[750]), .B(n2283), .Z(n18005) );
  AND U19045 ( .A(a[752]), .B(b[0]), .Z(n17985) );
  XNOR U19046 ( .A(n17985), .B(n2175), .Z(n17987) );
  NANDN U19047 ( .A(b[0]), .B(a[751]), .Z(n17986) );
  NAND U19048 ( .A(n17987), .B(n17986), .Z(n18010) );
  AND U19049 ( .A(a[748]), .B(b[3]), .Z(n18009) );
  XOR U19050 ( .A(n18010), .B(n18009), .Z(n18012) );
  XOR U19051 ( .A(n18011), .B(n18012), .Z(n18000) );
  NANDN U19052 ( .A(n17989), .B(n17988), .Z(n17993) );
  OR U19053 ( .A(n17991), .B(n17990), .Z(n17992) );
  AND U19054 ( .A(n17993), .B(n17992), .Z(n17999) );
  XOR U19055 ( .A(n18000), .B(n17999), .Z(n18002) );
  XOR U19056 ( .A(n18001), .B(n18002), .Z(n18015) );
  XNOR U19057 ( .A(n18015), .B(sreg[1772]), .Z(n18017) );
  NANDN U19058 ( .A(n17994), .B(sreg[1771]), .Z(n17998) );
  NAND U19059 ( .A(n17996), .B(n17995), .Z(n17997) );
  NAND U19060 ( .A(n17998), .B(n17997), .Z(n18016) );
  XOR U19061 ( .A(n18017), .B(n18016), .Z(c[1772]) );
  NANDN U19062 ( .A(n18000), .B(n17999), .Z(n18004) );
  OR U19063 ( .A(n18002), .B(n18001), .Z(n18003) );
  AND U19064 ( .A(n18004), .B(n18003), .Z(n18022) );
  XOR U19065 ( .A(a[751]), .B(n2283), .Z(n18026) );
  AND U19066 ( .A(a[753]), .B(b[0]), .Z(n18006) );
  XNOR U19067 ( .A(n18006), .B(n2175), .Z(n18008) );
  NANDN U19068 ( .A(b[0]), .B(a[752]), .Z(n18007) );
  NAND U19069 ( .A(n18008), .B(n18007), .Z(n18031) );
  AND U19070 ( .A(a[749]), .B(b[3]), .Z(n18030) );
  XOR U19071 ( .A(n18031), .B(n18030), .Z(n18033) );
  XOR U19072 ( .A(n18032), .B(n18033), .Z(n18021) );
  NANDN U19073 ( .A(n18010), .B(n18009), .Z(n18014) );
  OR U19074 ( .A(n18012), .B(n18011), .Z(n18013) );
  AND U19075 ( .A(n18014), .B(n18013), .Z(n18020) );
  XOR U19076 ( .A(n18021), .B(n18020), .Z(n18023) );
  XOR U19077 ( .A(n18022), .B(n18023), .Z(n18036) );
  XNOR U19078 ( .A(n18036), .B(sreg[1773]), .Z(n18038) );
  NANDN U19079 ( .A(n18015), .B(sreg[1772]), .Z(n18019) );
  NAND U19080 ( .A(n18017), .B(n18016), .Z(n18018) );
  NAND U19081 ( .A(n18019), .B(n18018), .Z(n18037) );
  XOR U19082 ( .A(n18038), .B(n18037), .Z(c[1773]) );
  NANDN U19083 ( .A(n18021), .B(n18020), .Z(n18025) );
  OR U19084 ( .A(n18023), .B(n18022), .Z(n18024) );
  AND U19085 ( .A(n18025), .B(n18024), .Z(n18043) );
  XOR U19086 ( .A(a[752]), .B(n2283), .Z(n18047) );
  AND U19087 ( .A(a[750]), .B(b[3]), .Z(n18051) );
  AND U19088 ( .A(a[754]), .B(b[0]), .Z(n18027) );
  XNOR U19089 ( .A(n18027), .B(n2175), .Z(n18029) );
  NANDN U19090 ( .A(b[0]), .B(a[753]), .Z(n18028) );
  NAND U19091 ( .A(n18029), .B(n18028), .Z(n18052) );
  XOR U19092 ( .A(n18051), .B(n18052), .Z(n18054) );
  XOR U19093 ( .A(n18053), .B(n18054), .Z(n18042) );
  NANDN U19094 ( .A(n18031), .B(n18030), .Z(n18035) );
  OR U19095 ( .A(n18033), .B(n18032), .Z(n18034) );
  AND U19096 ( .A(n18035), .B(n18034), .Z(n18041) );
  XOR U19097 ( .A(n18042), .B(n18041), .Z(n18044) );
  XOR U19098 ( .A(n18043), .B(n18044), .Z(n18057) );
  XNOR U19099 ( .A(n18057), .B(sreg[1774]), .Z(n18059) );
  NANDN U19100 ( .A(n18036), .B(sreg[1773]), .Z(n18040) );
  NAND U19101 ( .A(n18038), .B(n18037), .Z(n18039) );
  NAND U19102 ( .A(n18040), .B(n18039), .Z(n18058) );
  XOR U19103 ( .A(n18059), .B(n18058), .Z(c[1774]) );
  NANDN U19104 ( .A(n18042), .B(n18041), .Z(n18046) );
  OR U19105 ( .A(n18044), .B(n18043), .Z(n18045) );
  AND U19106 ( .A(n18046), .B(n18045), .Z(n18064) );
  XOR U19107 ( .A(a[753]), .B(n2283), .Z(n18068) );
  AND U19108 ( .A(a[751]), .B(b[3]), .Z(n18072) );
  AND U19109 ( .A(a[755]), .B(b[0]), .Z(n18048) );
  XNOR U19110 ( .A(n18048), .B(n2175), .Z(n18050) );
  NANDN U19111 ( .A(b[0]), .B(a[754]), .Z(n18049) );
  NAND U19112 ( .A(n18050), .B(n18049), .Z(n18073) );
  XOR U19113 ( .A(n18072), .B(n18073), .Z(n18075) );
  XOR U19114 ( .A(n18074), .B(n18075), .Z(n18063) );
  NANDN U19115 ( .A(n18052), .B(n18051), .Z(n18056) );
  OR U19116 ( .A(n18054), .B(n18053), .Z(n18055) );
  AND U19117 ( .A(n18056), .B(n18055), .Z(n18062) );
  XOR U19118 ( .A(n18063), .B(n18062), .Z(n18065) );
  XOR U19119 ( .A(n18064), .B(n18065), .Z(n18078) );
  XNOR U19120 ( .A(n18078), .B(sreg[1775]), .Z(n18080) );
  NANDN U19121 ( .A(n18057), .B(sreg[1774]), .Z(n18061) );
  NAND U19122 ( .A(n18059), .B(n18058), .Z(n18060) );
  NAND U19123 ( .A(n18061), .B(n18060), .Z(n18079) );
  XOR U19124 ( .A(n18080), .B(n18079), .Z(c[1775]) );
  NANDN U19125 ( .A(n18063), .B(n18062), .Z(n18067) );
  OR U19126 ( .A(n18065), .B(n18064), .Z(n18066) );
  AND U19127 ( .A(n18067), .B(n18066), .Z(n18085) );
  XOR U19128 ( .A(a[754]), .B(n2283), .Z(n18089) );
  AND U19129 ( .A(a[756]), .B(b[0]), .Z(n18069) );
  XNOR U19130 ( .A(n18069), .B(n2175), .Z(n18071) );
  NANDN U19131 ( .A(b[0]), .B(a[755]), .Z(n18070) );
  NAND U19132 ( .A(n18071), .B(n18070), .Z(n18094) );
  AND U19133 ( .A(a[752]), .B(b[3]), .Z(n18093) );
  XOR U19134 ( .A(n18094), .B(n18093), .Z(n18096) );
  XOR U19135 ( .A(n18095), .B(n18096), .Z(n18084) );
  NANDN U19136 ( .A(n18073), .B(n18072), .Z(n18077) );
  OR U19137 ( .A(n18075), .B(n18074), .Z(n18076) );
  AND U19138 ( .A(n18077), .B(n18076), .Z(n18083) );
  XOR U19139 ( .A(n18084), .B(n18083), .Z(n18086) );
  XOR U19140 ( .A(n18085), .B(n18086), .Z(n18099) );
  XNOR U19141 ( .A(n18099), .B(sreg[1776]), .Z(n18101) );
  NANDN U19142 ( .A(n18078), .B(sreg[1775]), .Z(n18082) );
  NAND U19143 ( .A(n18080), .B(n18079), .Z(n18081) );
  NAND U19144 ( .A(n18082), .B(n18081), .Z(n18100) );
  XOR U19145 ( .A(n18101), .B(n18100), .Z(c[1776]) );
  NANDN U19146 ( .A(n18084), .B(n18083), .Z(n18088) );
  OR U19147 ( .A(n18086), .B(n18085), .Z(n18087) );
  AND U19148 ( .A(n18088), .B(n18087), .Z(n18107) );
  XOR U19149 ( .A(a[755]), .B(n2284), .Z(n18108) );
  NAND U19150 ( .A(a[757]), .B(b[0]), .Z(n18090) );
  XNOR U19151 ( .A(b[1]), .B(n18090), .Z(n18092) );
  NANDN U19152 ( .A(b[0]), .B(a[756]), .Z(n18091) );
  AND U19153 ( .A(n18092), .B(n18091), .Z(n18112) );
  AND U19154 ( .A(a[753]), .B(b[3]), .Z(n18113) );
  XOR U19155 ( .A(n18112), .B(n18113), .Z(n18114) );
  XNOR U19156 ( .A(n18115), .B(n18114), .Z(n18104) );
  NANDN U19157 ( .A(n18094), .B(n18093), .Z(n18098) );
  OR U19158 ( .A(n18096), .B(n18095), .Z(n18097) );
  AND U19159 ( .A(n18098), .B(n18097), .Z(n18105) );
  XNOR U19160 ( .A(n18104), .B(n18105), .Z(n18106) );
  XNOR U19161 ( .A(n18107), .B(n18106), .Z(n18118) );
  XNOR U19162 ( .A(n18118), .B(sreg[1777]), .Z(n18120) );
  NANDN U19163 ( .A(n18099), .B(sreg[1776]), .Z(n18103) );
  NAND U19164 ( .A(n18101), .B(n18100), .Z(n18102) );
  NAND U19165 ( .A(n18103), .B(n18102), .Z(n18119) );
  XOR U19166 ( .A(n18120), .B(n18119), .Z(c[1777]) );
  XOR U19167 ( .A(a[756]), .B(n2284), .Z(n18127) );
  AND U19168 ( .A(a[758]), .B(b[0]), .Z(n18109) );
  XNOR U19169 ( .A(n18109), .B(n2175), .Z(n18111) );
  NANDN U19170 ( .A(b[0]), .B(a[757]), .Z(n18110) );
  NAND U19171 ( .A(n18111), .B(n18110), .Z(n18132) );
  AND U19172 ( .A(a[754]), .B(b[3]), .Z(n18131) );
  XOR U19173 ( .A(n18132), .B(n18131), .Z(n18134) );
  XOR U19174 ( .A(n18133), .B(n18134), .Z(n18122) );
  NAND U19175 ( .A(n18113), .B(n18112), .Z(n18117) );
  NANDN U19176 ( .A(n18115), .B(n18114), .Z(n18116) );
  AND U19177 ( .A(n18117), .B(n18116), .Z(n18121) );
  XOR U19178 ( .A(n18122), .B(n18121), .Z(n18124) );
  XOR U19179 ( .A(n18123), .B(n18124), .Z(n18137) );
  XNOR U19180 ( .A(n18137), .B(sreg[1778]), .Z(n18139) );
  XOR U19181 ( .A(n18139), .B(n18138), .Z(c[1778]) );
  NANDN U19182 ( .A(n18122), .B(n18121), .Z(n18126) );
  OR U19183 ( .A(n18124), .B(n18123), .Z(n18125) );
  AND U19184 ( .A(n18126), .B(n18125), .Z(n18144) );
  XOR U19185 ( .A(a[757]), .B(n2284), .Z(n18148) );
  AND U19186 ( .A(a[759]), .B(b[0]), .Z(n18128) );
  XNOR U19187 ( .A(n18128), .B(n2175), .Z(n18130) );
  NANDN U19188 ( .A(b[0]), .B(a[758]), .Z(n18129) );
  NAND U19189 ( .A(n18130), .B(n18129), .Z(n18153) );
  AND U19190 ( .A(a[755]), .B(b[3]), .Z(n18152) );
  XOR U19191 ( .A(n18153), .B(n18152), .Z(n18155) );
  XOR U19192 ( .A(n18154), .B(n18155), .Z(n18143) );
  NANDN U19193 ( .A(n18132), .B(n18131), .Z(n18136) );
  OR U19194 ( .A(n18134), .B(n18133), .Z(n18135) );
  AND U19195 ( .A(n18136), .B(n18135), .Z(n18142) );
  XOR U19196 ( .A(n18143), .B(n18142), .Z(n18145) );
  XOR U19197 ( .A(n18144), .B(n18145), .Z(n18158) );
  XNOR U19198 ( .A(n18158), .B(sreg[1779]), .Z(n18160) );
  NANDN U19199 ( .A(n18137), .B(sreg[1778]), .Z(n18141) );
  NAND U19200 ( .A(n18139), .B(n18138), .Z(n18140) );
  NAND U19201 ( .A(n18141), .B(n18140), .Z(n18159) );
  XOR U19202 ( .A(n18160), .B(n18159), .Z(c[1779]) );
  NANDN U19203 ( .A(n18143), .B(n18142), .Z(n18147) );
  OR U19204 ( .A(n18145), .B(n18144), .Z(n18146) );
  AND U19205 ( .A(n18147), .B(n18146), .Z(n18165) );
  XOR U19206 ( .A(a[758]), .B(n2284), .Z(n18169) );
  AND U19207 ( .A(a[756]), .B(b[3]), .Z(n18173) );
  AND U19208 ( .A(a[760]), .B(b[0]), .Z(n18149) );
  XNOR U19209 ( .A(n18149), .B(n2175), .Z(n18151) );
  NANDN U19210 ( .A(b[0]), .B(a[759]), .Z(n18150) );
  NAND U19211 ( .A(n18151), .B(n18150), .Z(n18174) );
  XOR U19212 ( .A(n18173), .B(n18174), .Z(n18176) );
  XOR U19213 ( .A(n18175), .B(n18176), .Z(n18164) );
  NANDN U19214 ( .A(n18153), .B(n18152), .Z(n18157) );
  OR U19215 ( .A(n18155), .B(n18154), .Z(n18156) );
  AND U19216 ( .A(n18157), .B(n18156), .Z(n18163) );
  XOR U19217 ( .A(n18164), .B(n18163), .Z(n18166) );
  XOR U19218 ( .A(n18165), .B(n18166), .Z(n18179) );
  XNOR U19219 ( .A(n18179), .B(sreg[1780]), .Z(n18181) );
  NANDN U19220 ( .A(n18158), .B(sreg[1779]), .Z(n18162) );
  NAND U19221 ( .A(n18160), .B(n18159), .Z(n18161) );
  NAND U19222 ( .A(n18162), .B(n18161), .Z(n18180) );
  XOR U19223 ( .A(n18181), .B(n18180), .Z(c[1780]) );
  NANDN U19224 ( .A(n18164), .B(n18163), .Z(n18168) );
  OR U19225 ( .A(n18166), .B(n18165), .Z(n18167) );
  AND U19226 ( .A(n18168), .B(n18167), .Z(n18186) );
  XOR U19227 ( .A(a[759]), .B(n2284), .Z(n18190) );
  AND U19228 ( .A(a[757]), .B(b[3]), .Z(n18194) );
  AND U19229 ( .A(a[761]), .B(b[0]), .Z(n18170) );
  XNOR U19230 ( .A(n18170), .B(n2175), .Z(n18172) );
  NANDN U19231 ( .A(b[0]), .B(a[760]), .Z(n18171) );
  NAND U19232 ( .A(n18172), .B(n18171), .Z(n18195) );
  XOR U19233 ( .A(n18194), .B(n18195), .Z(n18197) );
  XOR U19234 ( .A(n18196), .B(n18197), .Z(n18185) );
  NANDN U19235 ( .A(n18174), .B(n18173), .Z(n18178) );
  OR U19236 ( .A(n18176), .B(n18175), .Z(n18177) );
  AND U19237 ( .A(n18178), .B(n18177), .Z(n18184) );
  XOR U19238 ( .A(n18185), .B(n18184), .Z(n18187) );
  XOR U19239 ( .A(n18186), .B(n18187), .Z(n18200) );
  XNOR U19240 ( .A(n18200), .B(sreg[1781]), .Z(n18202) );
  NANDN U19241 ( .A(n18179), .B(sreg[1780]), .Z(n18183) );
  NAND U19242 ( .A(n18181), .B(n18180), .Z(n18182) );
  NAND U19243 ( .A(n18183), .B(n18182), .Z(n18201) );
  XOR U19244 ( .A(n18202), .B(n18201), .Z(c[1781]) );
  NANDN U19245 ( .A(n18185), .B(n18184), .Z(n18189) );
  OR U19246 ( .A(n18187), .B(n18186), .Z(n18188) );
  AND U19247 ( .A(n18189), .B(n18188), .Z(n18207) );
  XOR U19248 ( .A(a[760]), .B(n2284), .Z(n18211) );
  AND U19249 ( .A(a[762]), .B(b[0]), .Z(n18191) );
  XNOR U19250 ( .A(n18191), .B(n2175), .Z(n18193) );
  NANDN U19251 ( .A(b[0]), .B(a[761]), .Z(n18192) );
  NAND U19252 ( .A(n18193), .B(n18192), .Z(n18216) );
  AND U19253 ( .A(a[758]), .B(b[3]), .Z(n18215) );
  XOR U19254 ( .A(n18216), .B(n18215), .Z(n18218) );
  XOR U19255 ( .A(n18217), .B(n18218), .Z(n18206) );
  NANDN U19256 ( .A(n18195), .B(n18194), .Z(n18199) );
  OR U19257 ( .A(n18197), .B(n18196), .Z(n18198) );
  AND U19258 ( .A(n18199), .B(n18198), .Z(n18205) );
  XOR U19259 ( .A(n18206), .B(n18205), .Z(n18208) );
  XOR U19260 ( .A(n18207), .B(n18208), .Z(n18221) );
  XNOR U19261 ( .A(n18221), .B(sreg[1782]), .Z(n18223) );
  NANDN U19262 ( .A(n18200), .B(sreg[1781]), .Z(n18204) );
  NAND U19263 ( .A(n18202), .B(n18201), .Z(n18203) );
  NAND U19264 ( .A(n18204), .B(n18203), .Z(n18222) );
  XOR U19265 ( .A(n18223), .B(n18222), .Z(c[1782]) );
  NANDN U19266 ( .A(n18206), .B(n18205), .Z(n18210) );
  OR U19267 ( .A(n18208), .B(n18207), .Z(n18209) );
  AND U19268 ( .A(n18210), .B(n18209), .Z(n18228) );
  XOR U19269 ( .A(a[761]), .B(n2284), .Z(n18232) );
  AND U19270 ( .A(a[759]), .B(b[3]), .Z(n18236) );
  AND U19271 ( .A(a[763]), .B(b[0]), .Z(n18212) );
  XNOR U19272 ( .A(n18212), .B(n2175), .Z(n18214) );
  NANDN U19273 ( .A(b[0]), .B(a[762]), .Z(n18213) );
  NAND U19274 ( .A(n18214), .B(n18213), .Z(n18237) );
  XOR U19275 ( .A(n18236), .B(n18237), .Z(n18239) );
  XOR U19276 ( .A(n18238), .B(n18239), .Z(n18227) );
  NANDN U19277 ( .A(n18216), .B(n18215), .Z(n18220) );
  OR U19278 ( .A(n18218), .B(n18217), .Z(n18219) );
  AND U19279 ( .A(n18220), .B(n18219), .Z(n18226) );
  XOR U19280 ( .A(n18227), .B(n18226), .Z(n18229) );
  XOR U19281 ( .A(n18228), .B(n18229), .Z(n18242) );
  XNOR U19282 ( .A(n18242), .B(sreg[1783]), .Z(n18244) );
  NANDN U19283 ( .A(n18221), .B(sreg[1782]), .Z(n18225) );
  NAND U19284 ( .A(n18223), .B(n18222), .Z(n18224) );
  NAND U19285 ( .A(n18225), .B(n18224), .Z(n18243) );
  XOR U19286 ( .A(n18244), .B(n18243), .Z(c[1783]) );
  NANDN U19287 ( .A(n18227), .B(n18226), .Z(n18231) );
  OR U19288 ( .A(n18229), .B(n18228), .Z(n18230) );
  AND U19289 ( .A(n18231), .B(n18230), .Z(n18249) );
  XOR U19290 ( .A(a[762]), .B(n2285), .Z(n18253) );
  AND U19291 ( .A(a[764]), .B(b[0]), .Z(n18233) );
  XNOR U19292 ( .A(n18233), .B(n2175), .Z(n18235) );
  NANDN U19293 ( .A(b[0]), .B(a[763]), .Z(n18234) );
  NAND U19294 ( .A(n18235), .B(n18234), .Z(n18258) );
  AND U19295 ( .A(a[760]), .B(b[3]), .Z(n18257) );
  XOR U19296 ( .A(n18258), .B(n18257), .Z(n18260) );
  XOR U19297 ( .A(n18259), .B(n18260), .Z(n18248) );
  NANDN U19298 ( .A(n18237), .B(n18236), .Z(n18241) );
  OR U19299 ( .A(n18239), .B(n18238), .Z(n18240) );
  AND U19300 ( .A(n18241), .B(n18240), .Z(n18247) );
  XOR U19301 ( .A(n18248), .B(n18247), .Z(n18250) );
  XOR U19302 ( .A(n18249), .B(n18250), .Z(n18263) );
  XNOR U19303 ( .A(n18263), .B(sreg[1784]), .Z(n18265) );
  NANDN U19304 ( .A(n18242), .B(sreg[1783]), .Z(n18246) );
  NAND U19305 ( .A(n18244), .B(n18243), .Z(n18245) );
  NAND U19306 ( .A(n18246), .B(n18245), .Z(n18264) );
  XOR U19307 ( .A(n18265), .B(n18264), .Z(c[1784]) );
  NANDN U19308 ( .A(n18248), .B(n18247), .Z(n18252) );
  OR U19309 ( .A(n18250), .B(n18249), .Z(n18251) );
  AND U19310 ( .A(n18252), .B(n18251), .Z(n18270) );
  XOR U19311 ( .A(a[763]), .B(n2285), .Z(n18274) );
  AND U19312 ( .A(a[765]), .B(b[0]), .Z(n18254) );
  XNOR U19313 ( .A(n18254), .B(n2175), .Z(n18256) );
  NANDN U19314 ( .A(b[0]), .B(a[764]), .Z(n18255) );
  NAND U19315 ( .A(n18256), .B(n18255), .Z(n18279) );
  AND U19316 ( .A(a[761]), .B(b[3]), .Z(n18278) );
  XOR U19317 ( .A(n18279), .B(n18278), .Z(n18281) );
  XOR U19318 ( .A(n18280), .B(n18281), .Z(n18269) );
  NANDN U19319 ( .A(n18258), .B(n18257), .Z(n18262) );
  OR U19320 ( .A(n18260), .B(n18259), .Z(n18261) );
  AND U19321 ( .A(n18262), .B(n18261), .Z(n18268) );
  XOR U19322 ( .A(n18269), .B(n18268), .Z(n18271) );
  XOR U19323 ( .A(n18270), .B(n18271), .Z(n18284) );
  XNOR U19324 ( .A(n18284), .B(sreg[1785]), .Z(n18286) );
  NANDN U19325 ( .A(n18263), .B(sreg[1784]), .Z(n18267) );
  NAND U19326 ( .A(n18265), .B(n18264), .Z(n18266) );
  NAND U19327 ( .A(n18267), .B(n18266), .Z(n18285) );
  XOR U19328 ( .A(n18286), .B(n18285), .Z(c[1785]) );
  NANDN U19329 ( .A(n18269), .B(n18268), .Z(n18273) );
  OR U19330 ( .A(n18271), .B(n18270), .Z(n18272) );
  AND U19331 ( .A(n18273), .B(n18272), .Z(n18291) );
  XOR U19332 ( .A(a[764]), .B(n2285), .Z(n18295) );
  AND U19333 ( .A(a[766]), .B(b[0]), .Z(n18275) );
  XNOR U19334 ( .A(n18275), .B(n2175), .Z(n18277) );
  NANDN U19335 ( .A(b[0]), .B(a[765]), .Z(n18276) );
  NAND U19336 ( .A(n18277), .B(n18276), .Z(n18300) );
  AND U19337 ( .A(a[762]), .B(b[3]), .Z(n18299) );
  XOR U19338 ( .A(n18300), .B(n18299), .Z(n18302) );
  XOR U19339 ( .A(n18301), .B(n18302), .Z(n18290) );
  NANDN U19340 ( .A(n18279), .B(n18278), .Z(n18283) );
  OR U19341 ( .A(n18281), .B(n18280), .Z(n18282) );
  AND U19342 ( .A(n18283), .B(n18282), .Z(n18289) );
  XOR U19343 ( .A(n18290), .B(n18289), .Z(n18292) );
  XOR U19344 ( .A(n18291), .B(n18292), .Z(n18305) );
  XNOR U19345 ( .A(n18305), .B(sreg[1786]), .Z(n18307) );
  NANDN U19346 ( .A(n18284), .B(sreg[1785]), .Z(n18288) );
  NAND U19347 ( .A(n18286), .B(n18285), .Z(n18287) );
  NAND U19348 ( .A(n18288), .B(n18287), .Z(n18306) );
  XOR U19349 ( .A(n18307), .B(n18306), .Z(c[1786]) );
  NANDN U19350 ( .A(n18290), .B(n18289), .Z(n18294) );
  OR U19351 ( .A(n18292), .B(n18291), .Z(n18293) );
  AND U19352 ( .A(n18294), .B(n18293), .Z(n18312) );
  XOR U19353 ( .A(a[765]), .B(n2285), .Z(n18316) );
  AND U19354 ( .A(a[763]), .B(b[3]), .Z(n18320) );
  AND U19355 ( .A(a[767]), .B(b[0]), .Z(n18296) );
  XNOR U19356 ( .A(n18296), .B(n2175), .Z(n18298) );
  NANDN U19357 ( .A(b[0]), .B(a[766]), .Z(n18297) );
  NAND U19358 ( .A(n18298), .B(n18297), .Z(n18321) );
  XOR U19359 ( .A(n18320), .B(n18321), .Z(n18323) );
  XOR U19360 ( .A(n18322), .B(n18323), .Z(n18311) );
  NANDN U19361 ( .A(n18300), .B(n18299), .Z(n18304) );
  OR U19362 ( .A(n18302), .B(n18301), .Z(n18303) );
  AND U19363 ( .A(n18304), .B(n18303), .Z(n18310) );
  XOR U19364 ( .A(n18311), .B(n18310), .Z(n18313) );
  XOR U19365 ( .A(n18312), .B(n18313), .Z(n18326) );
  XNOR U19366 ( .A(n18326), .B(sreg[1787]), .Z(n18328) );
  NANDN U19367 ( .A(n18305), .B(sreg[1786]), .Z(n18309) );
  NAND U19368 ( .A(n18307), .B(n18306), .Z(n18308) );
  NAND U19369 ( .A(n18309), .B(n18308), .Z(n18327) );
  XOR U19370 ( .A(n18328), .B(n18327), .Z(c[1787]) );
  NANDN U19371 ( .A(n18311), .B(n18310), .Z(n18315) );
  OR U19372 ( .A(n18313), .B(n18312), .Z(n18314) );
  AND U19373 ( .A(n18315), .B(n18314), .Z(n18333) );
  XOR U19374 ( .A(a[766]), .B(n2285), .Z(n18337) );
  AND U19375 ( .A(a[768]), .B(b[0]), .Z(n18317) );
  XNOR U19376 ( .A(n18317), .B(n2175), .Z(n18319) );
  NANDN U19377 ( .A(b[0]), .B(a[767]), .Z(n18318) );
  NAND U19378 ( .A(n18319), .B(n18318), .Z(n18342) );
  AND U19379 ( .A(a[764]), .B(b[3]), .Z(n18341) );
  XOR U19380 ( .A(n18342), .B(n18341), .Z(n18344) );
  XOR U19381 ( .A(n18343), .B(n18344), .Z(n18332) );
  NANDN U19382 ( .A(n18321), .B(n18320), .Z(n18325) );
  OR U19383 ( .A(n18323), .B(n18322), .Z(n18324) );
  AND U19384 ( .A(n18325), .B(n18324), .Z(n18331) );
  XOR U19385 ( .A(n18332), .B(n18331), .Z(n18334) );
  XOR U19386 ( .A(n18333), .B(n18334), .Z(n18347) );
  XNOR U19387 ( .A(n18347), .B(sreg[1788]), .Z(n18349) );
  NANDN U19388 ( .A(n18326), .B(sreg[1787]), .Z(n18330) );
  NAND U19389 ( .A(n18328), .B(n18327), .Z(n18329) );
  NAND U19390 ( .A(n18330), .B(n18329), .Z(n18348) );
  XOR U19391 ( .A(n18349), .B(n18348), .Z(c[1788]) );
  NANDN U19392 ( .A(n18332), .B(n18331), .Z(n18336) );
  OR U19393 ( .A(n18334), .B(n18333), .Z(n18335) );
  AND U19394 ( .A(n18336), .B(n18335), .Z(n18354) );
  XOR U19395 ( .A(a[767]), .B(n2285), .Z(n18358) );
  AND U19396 ( .A(a[765]), .B(b[3]), .Z(n18362) );
  AND U19397 ( .A(a[769]), .B(b[0]), .Z(n18338) );
  XNOR U19398 ( .A(n18338), .B(n2175), .Z(n18340) );
  NANDN U19399 ( .A(b[0]), .B(a[768]), .Z(n18339) );
  NAND U19400 ( .A(n18340), .B(n18339), .Z(n18363) );
  XOR U19401 ( .A(n18362), .B(n18363), .Z(n18365) );
  XOR U19402 ( .A(n18364), .B(n18365), .Z(n18353) );
  NANDN U19403 ( .A(n18342), .B(n18341), .Z(n18346) );
  OR U19404 ( .A(n18344), .B(n18343), .Z(n18345) );
  AND U19405 ( .A(n18346), .B(n18345), .Z(n18352) );
  XOR U19406 ( .A(n18353), .B(n18352), .Z(n18355) );
  XOR U19407 ( .A(n18354), .B(n18355), .Z(n18368) );
  XNOR U19408 ( .A(n18368), .B(sreg[1789]), .Z(n18370) );
  NANDN U19409 ( .A(n18347), .B(sreg[1788]), .Z(n18351) );
  NAND U19410 ( .A(n18349), .B(n18348), .Z(n18350) );
  NAND U19411 ( .A(n18351), .B(n18350), .Z(n18369) );
  XOR U19412 ( .A(n18370), .B(n18369), .Z(c[1789]) );
  NANDN U19413 ( .A(n18353), .B(n18352), .Z(n18357) );
  OR U19414 ( .A(n18355), .B(n18354), .Z(n18356) );
  AND U19415 ( .A(n18357), .B(n18356), .Z(n18375) );
  XOR U19416 ( .A(a[768]), .B(n2285), .Z(n18379) );
  AND U19417 ( .A(a[766]), .B(b[3]), .Z(n18383) );
  AND U19418 ( .A(a[770]), .B(b[0]), .Z(n18359) );
  XNOR U19419 ( .A(n18359), .B(n2175), .Z(n18361) );
  NANDN U19420 ( .A(b[0]), .B(a[769]), .Z(n18360) );
  NAND U19421 ( .A(n18361), .B(n18360), .Z(n18384) );
  XOR U19422 ( .A(n18383), .B(n18384), .Z(n18386) );
  XOR U19423 ( .A(n18385), .B(n18386), .Z(n18374) );
  NANDN U19424 ( .A(n18363), .B(n18362), .Z(n18367) );
  OR U19425 ( .A(n18365), .B(n18364), .Z(n18366) );
  AND U19426 ( .A(n18367), .B(n18366), .Z(n18373) );
  XOR U19427 ( .A(n18374), .B(n18373), .Z(n18376) );
  XOR U19428 ( .A(n18375), .B(n18376), .Z(n18389) );
  XNOR U19429 ( .A(n18389), .B(sreg[1790]), .Z(n18391) );
  NANDN U19430 ( .A(n18368), .B(sreg[1789]), .Z(n18372) );
  NAND U19431 ( .A(n18370), .B(n18369), .Z(n18371) );
  NAND U19432 ( .A(n18372), .B(n18371), .Z(n18390) );
  XOR U19433 ( .A(n18391), .B(n18390), .Z(c[1790]) );
  NANDN U19434 ( .A(n18374), .B(n18373), .Z(n18378) );
  OR U19435 ( .A(n18376), .B(n18375), .Z(n18377) );
  AND U19436 ( .A(n18378), .B(n18377), .Z(n18396) );
  XOR U19437 ( .A(a[769]), .B(n2286), .Z(n18400) );
  AND U19438 ( .A(a[771]), .B(b[0]), .Z(n18380) );
  XNOR U19439 ( .A(n18380), .B(n2175), .Z(n18382) );
  NANDN U19440 ( .A(b[0]), .B(a[770]), .Z(n18381) );
  NAND U19441 ( .A(n18382), .B(n18381), .Z(n18405) );
  AND U19442 ( .A(a[767]), .B(b[3]), .Z(n18404) );
  XOR U19443 ( .A(n18405), .B(n18404), .Z(n18407) );
  XOR U19444 ( .A(n18406), .B(n18407), .Z(n18395) );
  NANDN U19445 ( .A(n18384), .B(n18383), .Z(n18388) );
  OR U19446 ( .A(n18386), .B(n18385), .Z(n18387) );
  AND U19447 ( .A(n18388), .B(n18387), .Z(n18394) );
  XOR U19448 ( .A(n18395), .B(n18394), .Z(n18397) );
  XOR U19449 ( .A(n18396), .B(n18397), .Z(n18410) );
  XNOR U19450 ( .A(n18410), .B(sreg[1791]), .Z(n18412) );
  NANDN U19451 ( .A(n18389), .B(sreg[1790]), .Z(n18393) );
  NAND U19452 ( .A(n18391), .B(n18390), .Z(n18392) );
  NAND U19453 ( .A(n18393), .B(n18392), .Z(n18411) );
  XOR U19454 ( .A(n18412), .B(n18411), .Z(c[1791]) );
  NANDN U19455 ( .A(n18395), .B(n18394), .Z(n18399) );
  OR U19456 ( .A(n18397), .B(n18396), .Z(n18398) );
  AND U19457 ( .A(n18399), .B(n18398), .Z(n18417) );
  XOR U19458 ( .A(a[770]), .B(n2286), .Z(n18421) );
  AND U19459 ( .A(a[772]), .B(b[0]), .Z(n18401) );
  XNOR U19460 ( .A(n18401), .B(n2175), .Z(n18403) );
  NANDN U19461 ( .A(b[0]), .B(a[771]), .Z(n18402) );
  NAND U19462 ( .A(n18403), .B(n18402), .Z(n18426) );
  AND U19463 ( .A(a[768]), .B(b[3]), .Z(n18425) );
  XOR U19464 ( .A(n18426), .B(n18425), .Z(n18428) );
  XOR U19465 ( .A(n18427), .B(n18428), .Z(n18416) );
  NANDN U19466 ( .A(n18405), .B(n18404), .Z(n18409) );
  OR U19467 ( .A(n18407), .B(n18406), .Z(n18408) );
  AND U19468 ( .A(n18409), .B(n18408), .Z(n18415) );
  XOR U19469 ( .A(n18416), .B(n18415), .Z(n18418) );
  XOR U19470 ( .A(n18417), .B(n18418), .Z(n18431) );
  XNOR U19471 ( .A(n18431), .B(sreg[1792]), .Z(n18433) );
  NANDN U19472 ( .A(n18410), .B(sreg[1791]), .Z(n18414) );
  NAND U19473 ( .A(n18412), .B(n18411), .Z(n18413) );
  NAND U19474 ( .A(n18414), .B(n18413), .Z(n18432) );
  XOR U19475 ( .A(n18433), .B(n18432), .Z(c[1792]) );
  NANDN U19476 ( .A(n18416), .B(n18415), .Z(n18420) );
  OR U19477 ( .A(n18418), .B(n18417), .Z(n18419) );
  AND U19478 ( .A(n18420), .B(n18419), .Z(n18438) );
  XOR U19479 ( .A(a[771]), .B(n2286), .Z(n18442) );
  AND U19480 ( .A(a[769]), .B(b[3]), .Z(n18446) );
  AND U19481 ( .A(a[773]), .B(b[0]), .Z(n18422) );
  XNOR U19482 ( .A(n18422), .B(n2175), .Z(n18424) );
  NANDN U19483 ( .A(b[0]), .B(a[772]), .Z(n18423) );
  NAND U19484 ( .A(n18424), .B(n18423), .Z(n18447) );
  XOR U19485 ( .A(n18446), .B(n18447), .Z(n18449) );
  XOR U19486 ( .A(n18448), .B(n18449), .Z(n18437) );
  NANDN U19487 ( .A(n18426), .B(n18425), .Z(n18430) );
  OR U19488 ( .A(n18428), .B(n18427), .Z(n18429) );
  AND U19489 ( .A(n18430), .B(n18429), .Z(n18436) );
  XOR U19490 ( .A(n18437), .B(n18436), .Z(n18439) );
  XOR U19491 ( .A(n18438), .B(n18439), .Z(n18452) );
  XNOR U19492 ( .A(n18452), .B(sreg[1793]), .Z(n18454) );
  NANDN U19493 ( .A(n18431), .B(sreg[1792]), .Z(n18435) );
  NAND U19494 ( .A(n18433), .B(n18432), .Z(n18434) );
  NAND U19495 ( .A(n18435), .B(n18434), .Z(n18453) );
  XOR U19496 ( .A(n18454), .B(n18453), .Z(c[1793]) );
  NANDN U19497 ( .A(n18437), .B(n18436), .Z(n18441) );
  OR U19498 ( .A(n18439), .B(n18438), .Z(n18440) );
  AND U19499 ( .A(n18441), .B(n18440), .Z(n18459) );
  XOR U19500 ( .A(a[772]), .B(n2286), .Z(n18463) );
  AND U19501 ( .A(a[774]), .B(b[0]), .Z(n18443) );
  XNOR U19502 ( .A(n18443), .B(n2175), .Z(n18445) );
  NANDN U19503 ( .A(b[0]), .B(a[773]), .Z(n18444) );
  NAND U19504 ( .A(n18445), .B(n18444), .Z(n18468) );
  AND U19505 ( .A(a[770]), .B(b[3]), .Z(n18467) );
  XOR U19506 ( .A(n18468), .B(n18467), .Z(n18470) );
  XOR U19507 ( .A(n18469), .B(n18470), .Z(n18458) );
  NANDN U19508 ( .A(n18447), .B(n18446), .Z(n18451) );
  OR U19509 ( .A(n18449), .B(n18448), .Z(n18450) );
  AND U19510 ( .A(n18451), .B(n18450), .Z(n18457) );
  XOR U19511 ( .A(n18458), .B(n18457), .Z(n18460) );
  XOR U19512 ( .A(n18459), .B(n18460), .Z(n18473) );
  XNOR U19513 ( .A(n18473), .B(sreg[1794]), .Z(n18475) );
  NANDN U19514 ( .A(n18452), .B(sreg[1793]), .Z(n18456) );
  NAND U19515 ( .A(n18454), .B(n18453), .Z(n18455) );
  NAND U19516 ( .A(n18456), .B(n18455), .Z(n18474) );
  XOR U19517 ( .A(n18475), .B(n18474), .Z(c[1794]) );
  NANDN U19518 ( .A(n18458), .B(n18457), .Z(n18462) );
  OR U19519 ( .A(n18460), .B(n18459), .Z(n18461) );
  AND U19520 ( .A(n18462), .B(n18461), .Z(n18480) );
  XOR U19521 ( .A(a[773]), .B(n2286), .Z(n18484) );
  AND U19522 ( .A(a[775]), .B(b[0]), .Z(n18464) );
  XNOR U19523 ( .A(n18464), .B(n2175), .Z(n18466) );
  NANDN U19524 ( .A(b[0]), .B(a[774]), .Z(n18465) );
  NAND U19525 ( .A(n18466), .B(n18465), .Z(n18489) );
  AND U19526 ( .A(a[771]), .B(b[3]), .Z(n18488) );
  XOR U19527 ( .A(n18489), .B(n18488), .Z(n18491) );
  XOR U19528 ( .A(n18490), .B(n18491), .Z(n18479) );
  NANDN U19529 ( .A(n18468), .B(n18467), .Z(n18472) );
  OR U19530 ( .A(n18470), .B(n18469), .Z(n18471) );
  AND U19531 ( .A(n18472), .B(n18471), .Z(n18478) );
  XOR U19532 ( .A(n18479), .B(n18478), .Z(n18481) );
  XOR U19533 ( .A(n18480), .B(n18481), .Z(n18494) );
  XNOR U19534 ( .A(n18494), .B(sreg[1795]), .Z(n18496) );
  NANDN U19535 ( .A(n18473), .B(sreg[1794]), .Z(n18477) );
  NAND U19536 ( .A(n18475), .B(n18474), .Z(n18476) );
  NAND U19537 ( .A(n18477), .B(n18476), .Z(n18495) );
  XOR U19538 ( .A(n18496), .B(n18495), .Z(c[1795]) );
  NANDN U19539 ( .A(n18479), .B(n18478), .Z(n18483) );
  OR U19540 ( .A(n18481), .B(n18480), .Z(n18482) );
  AND U19541 ( .A(n18483), .B(n18482), .Z(n18501) );
  XOR U19542 ( .A(a[774]), .B(n2286), .Z(n18505) );
  AND U19543 ( .A(a[772]), .B(b[3]), .Z(n18509) );
  AND U19544 ( .A(a[776]), .B(b[0]), .Z(n18485) );
  XNOR U19545 ( .A(n18485), .B(n2175), .Z(n18487) );
  NANDN U19546 ( .A(b[0]), .B(a[775]), .Z(n18486) );
  NAND U19547 ( .A(n18487), .B(n18486), .Z(n18510) );
  XOR U19548 ( .A(n18509), .B(n18510), .Z(n18512) );
  XOR U19549 ( .A(n18511), .B(n18512), .Z(n18500) );
  NANDN U19550 ( .A(n18489), .B(n18488), .Z(n18493) );
  OR U19551 ( .A(n18491), .B(n18490), .Z(n18492) );
  AND U19552 ( .A(n18493), .B(n18492), .Z(n18499) );
  XOR U19553 ( .A(n18500), .B(n18499), .Z(n18502) );
  XOR U19554 ( .A(n18501), .B(n18502), .Z(n18515) );
  XNOR U19555 ( .A(n18515), .B(sreg[1796]), .Z(n18517) );
  NANDN U19556 ( .A(n18494), .B(sreg[1795]), .Z(n18498) );
  NAND U19557 ( .A(n18496), .B(n18495), .Z(n18497) );
  NAND U19558 ( .A(n18498), .B(n18497), .Z(n18516) );
  XOR U19559 ( .A(n18517), .B(n18516), .Z(c[1796]) );
  NANDN U19560 ( .A(n18500), .B(n18499), .Z(n18504) );
  OR U19561 ( .A(n18502), .B(n18501), .Z(n18503) );
  AND U19562 ( .A(n18504), .B(n18503), .Z(n18522) );
  XOR U19563 ( .A(a[775]), .B(n2286), .Z(n18526) );
  AND U19564 ( .A(a[777]), .B(b[0]), .Z(n18506) );
  XNOR U19565 ( .A(n18506), .B(n2175), .Z(n18508) );
  NANDN U19566 ( .A(b[0]), .B(a[776]), .Z(n18507) );
  NAND U19567 ( .A(n18508), .B(n18507), .Z(n18531) );
  AND U19568 ( .A(a[773]), .B(b[3]), .Z(n18530) );
  XOR U19569 ( .A(n18531), .B(n18530), .Z(n18533) );
  XOR U19570 ( .A(n18532), .B(n18533), .Z(n18521) );
  NANDN U19571 ( .A(n18510), .B(n18509), .Z(n18514) );
  OR U19572 ( .A(n18512), .B(n18511), .Z(n18513) );
  AND U19573 ( .A(n18514), .B(n18513), .Z(n18520) );
  XOR U19574 ( .A(n18521), .B(n18520), .Z(n18523) );
  XOR U19575 ( .A(n18522), .B(n18523), .Z(n18536) );
  XNOR U19576 ( .A(n18536), .B(sreg[1797]), .Z(n18538) );
  NANDN U19577 ( .A(n18515), .B(sreg[1796]), .Z(n18519) );
  NAND U19578 ( .A(n18517), .B(n18516), .Z(n18518) );
  NAND U19579 ( .A(n18519), .B(n18518), .Z(n18537) );
  XOR U19580 ( .A(n18538), .B(n18537), .Z(c[1797]) );
  NANDN U19581 ( .A(n18521), .B(n18520), .Z(n18525) );
  OR U19582 ( .A(n18523), .B(n18522), .Z(n18524) );
  AND U19583 ( .A(n18525), .B(n18524), .Z(n18543) );
  XOR U19584 ( .A(a[776]), .B(n2287), .Z(n18547) );
  AND U19585 ( .A(a[778]), .B(b[0]), .Z(n18527) );
  XNOR U19586 ( .A(n18527), .B(n2175), .Z(n18529) );
  NANDN U19587 ( .A(b[0]), .B(a[777]), .Z(n18528) );
  NAND U19588 ( .A(n18529), .B(n18528), .Z(n18552) );
  AND U19589 ( .A(a[774]), .B(b[3]), .Z(n18551) );
  XOR U19590 ( .A(n18552), .B(n18551), .Z(n18554) );
  XOR U19591 ( .A(n18553), .B(n18554), .Z(n18542) );
  NANDN U19592 ( .A(n18531), .B(n18530), .Z(n18535) );
  OR U19593 ( .A(n18533), .B(n18532), .Z(n18534) );
  AND U19594 ( .A(n18535), .B(n18534), .Z(n18541) );
  XOR U19595 ( .A(n18542), .B(n18541), .Z(n18544) );
  XOR U19596 ( .A(n18543), .B(n18544), .Z(n18557) );
  XNOR U19597 ( .A(n18557), .B(sreg[1798]), .Z(n18559) );
  NANDN U19598 ( .A(n18536), .B(sreg[1797]), .Z(n18540) );
  NAND U19599 ( .A(n18538), .B(n18537), .Z(n18539) );
  NAND U19600 ( .A(n18540), .B(n18539), .Z(n18558) );
  XOR U19601 ( .A(n18559), .B(n18558), .Z(c[1798]) );
  NANDN U19602 ( .A(n18542), .B(n18541), .Z(n18546) );
  OR U19603 ( .A(n18544), .B(n18543), .Z(n18545) );
  AND U19604 ( .A(n18546), .B(n18545), .Z(n18564) );
  XOR U19605 ( .A(a[777]), .B(n2287), .Z(n18568) );
  AND U19606 ( .A(a[779]), .B(b[0]), .Z(n18548) );
  XNOR U19607 ( .A(n18548), .B(n2175), .Z(n18550) );
  NANDN U19608 ( .A(b[0]), .B(a[778]), .Z(n18549) );
  NAND U19609 ( .A(n18550), .B(n18549), .Z(n18573) );
  AND U19610 ( .A(a[775]), .B(b[3]), .Z(n18572) );
  XOR U19611 ( .A(n18573), .B(n18572), .Z(n18575) );
  XOR U19612 ( .A(n18574), .B(n18575), .Z(n18563) );
  NANDN U19613 ( .A(n18552), .B(n18551), .Z(n18556) );
  OR U19614 ( .A(n18554), .B(n18553), .Z(n18555) );
  AND U19615 ( .A(n18556), .B(n18555), .Z(n18562) );
  XOR U19616 ( .A(n18563), .B(n18562), .Z(n18565) );
  XOR U19617 ( .A(n18564), .B(n18565), .Z(n18578) );
  XNOR U19618 ( .A(n18578), .B(sreg[1799]), .Z(n18580) );
  NANDN U19619 ( .A(n18557), .B(sreg[1798]), .Z(n18561) );
  NAND U19620 ( .A(n18559), .B(n18558), .Z(n18560) );
  NAND U19621 ( .A(n18561), .B(n18560), .Z(n18579) );
  XOR U19622 ( .A(n18580), .B(n18579), .Z(c[1799]) );
  NANDN U19623 ( .A(n18563), .B(n18562), .Z(n18567) );
  OR U19624 ( .A(n18565), .B(n18564), .Z(n18566) );
  AND U19625 ( .A(n18567), .B(n18566), .Z(n18585) );
  XOR U19626 ( .A(a[778]), .B(n2287), .Z(n18589) );
  AND U19627 ( .A(a[780]), .B(b[0]), .Z(n18569) );
  XNOR U19628 ( .A(n18569), .B(n2175), .Z(n18571) );
  NANDN U19629 ( .A(b[0]), .B(a[779]), .Z(n18570) );
  NAND U19630 ( .A(n18571), .B(n18570), .Z(n18594) );
  AND U19631 ( .A(a[776]), .B(b[3]), .Z(n18593) );
  XOR U19632 ( .A(n18594), .B(n18593), .Z(n18596) );
  XOR U19633 ( .A(n18595), .B(n18596), .Z(n18584) );
  NANDN U19634 ( .A(n18573), .B(n18572), .Z(n18577) );
  OR U19635 ( .A(n18575), .B(n18574), .Z(n18576) );
  AND U19636 ( .A(n18577), .B(n18576), .Z(n18583) );
  XOR U19637 ( .A(n18584), .B(n18583), .Z(n18586) );
  XOR U19638 ( .A(n18585), .B(n18586), .Z(n18599) );
  XNOR U19639 ( .A(n18599), .B(sreg[1800]), .Z(n18601) );
  NANDN U19640 ( .A(n18578), .B(sreg[1799]), .Z(n18582) );
  NAND U19641 ( .A(n18580), .B(n18579), .Z(n18581) );
  NAND U19642 ( .A(n18582), .B(n18581), .Z(n18600) );
  XOR U19643 ( .A(n18601), .B(n18600), .Z(c[1800]) );
  NANDN U19644 ( .A(n18584), .B(n18583), .Z(n18588) );
  OR U19645 ( .A(n18586), .B(n18585), .Z(n18587) );
  AND U19646 ( .A(n18588), .B(n18587), .Z(n18606) );
  XOR U19647 ( .A(a[779]), .B(n2287), .Z(n18610) );
  AND U19648 ( .A(a[781]), .B(b[0]), .Z(n18590) );
  XNOR U19649 ( .A(n18590), .B(n2175), .Z(n18592) );
  NANDN U19650 ( .A(b[0]), .B(a[780]), .Z(n18591) );
  NAND U19651 ( .A(n18592), .B(n18591), .Z(n18615) );
  AND U19652 ( .A(a[777]), .B(b[3]), .Z(n18614) );
  XOR U19653 ( .A(n18615), .B(n18614), .Z(n18617) );
  XOR U19654 ( .A(n18616), .B(n18617), .Z(n18605) );
  NANDN U19655 ( .A(n18594), .B(n18593), .Z(n18598) );
  OR U19656 ( .A(n18596), .B(n18595), .Z(n18597) );
  AND U19657 ( .A(n18598), .B(n18597), .Z(n18604) );
  XOR U19658 ( .A(n18605), .B(n18604), .Z(n18607) );
  XOR U19659 ( .A(n18606), .B(n18607), .Z(n18620) );
  XNOR U19660 ( .A(n18620), .B(sreg[1801]), .Z(n18622) );
  NANDN U19661 ( .A(n18599), .B(sreg[1800]), .Z(n18603) );
  NAND U19662 ( .A(n18601), .B(n18600), .Z(n18602) );
  NAND U19663 ( .A(n18603), .B(n18602), .Z(n18621) );
  XOR U19664 ( .A(n18622), .B(n18621), .Z(c[1801]) );
  NANDN U19665 ( .A(n18605), .B(n18604), .Z(n18609) );
  OR U19666 ( .A(n18607), .B(n18606), .Z(n18608) );
  AND U19667 ( .A(n18609), .B(n18608), .Z(n18627) );
  XOR U19668 ( .A(a[780]), .B(n2287), .Z(n18631) );
  AND U19669 ( .A(a[782]), .B(b[0]), .Z(n18611) );
  XNOR U19670 ( .A(n18611), .B(n2175), .Z(n18613) );
  NANDN U19671 ( .A(b[0]), .B(a[781]), .Z(n18612) );
  NAND U19672 ( .A(n18613), .B(n18612), .Z(n18636) );
  AND U19673 ( .A(a[778]), .B(b[3]), .Z(n18635) );
  XOR U19674 ( .A(n18636), .B(n18635), .Z(n18638) );
  XOR U19675 ( .A(n18637), .B(n18638), .Z(n18626) );
  NANDN U19676 ( .A(n18615), .B(n18614), .Z(n18619) );
  OR U19677 ( .A(n18617), .B(n18616), .Z(n18618) );
  AND U19678 ( .A(n18619), .B(n18618), .Z(n18625) );
  XOR U19679 ( .A(n18626), .B(n18625), .Z(n18628) );
  XOR U19680 ( .A(n18627), .B(n18628), .Z(n18641) );
  XNOR U19681 ( .A(n18641), .B(sreg[1802]), .Z(n18643) );
  NANDN U19682 ( .A(n18620), .B(sreg[1801]), .Z(n18624) );
  NAND U19683 ( .A(n18622), .B(n18621), .Z(n18623) );
  NAND U19684 ( .A(n18624), .B(n18623), .Z(n18642) );
  XOR U19685 ( .A(n18643), .B(n18642), .Z(c[1802]) );
  NANDN U19686 ( .A(n18626), .B(n18625), .Z(n18630) );
  OR U19687 ( .A(n18628), .B(n18627), .Z(n18629) );
  AND U19688 ( .A(n18630), .B(n18629), .Z(n18648) );
  XOR U19689 ( .A(a[781]), .B(n2287), .Z(n18652) );
  AND U19690 ( .A(a[783]), .B(b[0]), .Z(n18632) );
  XNOR U19691 ( .A(n18632), .B(n2175), .Z(n18634) );
  NANDN U19692 ( .A(b[0]), .B(a[782]), .Z(n18633) );
  NAND U19693 ( .A(n18634), .B(n18633), .Z(n18657) );
  AND U19694 ( .A(a[779]), .B(b[3]), .Z(n18656) );
  XOR U19695 ( .A(n18657), .B(n18656), .Z(n18659) );
  XOR U19696 ( .A(n18658), .B(n18659), .Z(n18647) );
  NANDN U19697 ( .A(n18636), .B(n18635), .Z(n18640) );
  OR U19698 ( .A(n18638), .B(n18637), .Z(n18639) );
  AND U19699 ( .A(n18640), .B(n18639), .Z(n18646) );
  XOR U19700 ( .A(n18647), .B(n18646), .Z(n18649) );
  XOR U19701 ( .A(n18648), .B(n18649), .Z(n18662) );
  XNOR U19702 ( .A(n18662), .B(sreg[1803]), .Z(n18664) );
  NANDN U19703 ( .A(n18641), .B(sreg[1802]), .Z(n18645) );
  NAND U19704 ( .A(n18643), .B(n18642), .Z(n18644) );
  NAND U19705 ( .A(n18645), .B(n18644), .Z(n18663) );
  XOR U19706 ( .A(n18664), .B(n18663), .Z(c[1803]) );
  NANDN U19707 ( .A(n18647), .B(n18646), .Z(n18651) );
  OR U19708 ( .A(n18649), .B(n18648), .Z(n18650) );
  AND U19709 ( .A(n18651), .B(n18650), .Z(n18669) );
  XOR U19710 ( .A(a[782]), .B(n2287), .Z(n18673) );
  AND U19711 ( .A(a[784]), .B(b[0]), .Z(n18653) );
  XNOR U19712 ( .A(n18653), .B(n2175), .Z(n18655) );
  NANDN U19713 ( .A(b[0]), .B(a[783]), .Z(n18654) );
  NAND U19714 ( .A(n18655), .B(n18654), .Z(n18678) );
  AND U19715 ( .A(a[780]), .B(b[3]), .Z(n18677) );
  XOR U19716 ( .A(n18678), .B(n18677), .Z(n18680) );
  XOR U19717 ( .A(n18679), .B(n18680), .Z(n18668) );
  NANDN U19718 ( .A(n18657), .B(n18656), .Z(n18661) );
  OR U19719 ( .A(n18659), .B(n18658), .Z(n18660) );
  AND U19720 ( .A(n18661), .B(n18660), .Z(n18667) );
  XOR U19721 ( .A(n18668), .B(n18667), .Z(n18670) );
  XOR U19722 ( .A(n18669), .B(n18670), .Z(n18683) );
  XNOR U19723 ( .A(n18683), .B(sreg[1804]), .Z(n18685) );
  NANDN U19724 ( .A(n18662), .B(sreg[1803]), .Z(n18666) );
  NAND U19725 ( .A(n18664), .B(n18663), .Z(n18665) );
  NAND U19726 ( .A(n18666), .B(n18665), .Z(n18684) );
  XOR U19727 ( .A(n18685), .B(n18684), .Z(c[1804]) );
  NANDN U19728 ( .A(n18668), .B(n18667), .Z(n18672) );
  OR U19729 ( .A(n18670), .B(n18669), .Z(n18671) );
  AND U19730 ( .A(n18672), .B(n18671), .Z(n18690) );
  XOR U19731 ( .A(a[783]), .B(n2288), .Z(n18694) );
  AND U19732 ( .A(a[785]), .B(b[0]), .Z(n18674) );
  XNOR U19733 ( .A(n18674), .B(n2175), .Z(n18676) );
  NANDN U19734 ( .A(b[0]), .B(a[784]), .Z(n18675) );
  NAND U19735 ( .A(n18676), .B(n18675), .Z(n18699) );
  AND U19736 ( .A(a[781]), .B(b[3]), .Z(n18698) );
  XOR U19737 ( .A(n18699), .B(n18698), .Z(n18701) );
  XOR U19738 ( .A(n18700), .B(n18701), .Z(n18689) );
  NANDN U19739 ( .A(n18678), .B(n18677), .Z(n18682) );
  OR U19740 ( .A(n18680), .B(n18679), .Z(n18681) );
  AND U19741 ( .A(n18682), .B(n18681), .Z(n18688) );
  XOR U19742 ( .A(n18689), .B(n18688), .Z(n18691) );
  XOR U19743 ( .A(n18690), .B(n18691), .Z(n18704) );
  XNOR U19744 ( .A(n18704), .B(sreg[1805]), .Z(n18706) );
  NANDN U19745 ( .A(n18683), .B(sreg[1804]), .Z(n18687) );
  NAND U19746 ( .A(n18685), .B(n18684), .Z(n18686) );
  NAND U19747 ( .A(n18687), .B(n18686), .Z(n18705) );
  XOR U19748 ( .A(n18706), .B(n18705), .Z(c[1805]) );
  NANDN U19749 ( .A(n18689), .B(n18688), .Z(n18693) );
  OR U19750 ( .A(n18691), .B(n18690), .Z(n18692) );
  AND U19751 ( .A(n18693), .B(n18692), .Z(n18711) );
  XOR U19752 ( .A(a[784]), .B(n2288), .Z(n18715) );
  AND U19753 ( .A(a[782]), .B(b[3]), .Z(n18719) );
  AND U19754 ( .A(a[786]), .B(b[0]), .Z(n18695) );
  XNOR U19755 ( .A(n18695), .B(n2175), .Z(n18697) );
  NANDN U19756 ( .A(b[0]), .B(a[785]), .Z(n18696) );
  NAND U19757 ( .A(n18697), .B(n18696), .Z(n18720) );
  XOR U19758 ( .A(n18719), .B(n18720), .Z(n18722) );
  XOR U19759 ( .A(n18721), .B(n18722), .Z(n18710) );
  NANDN U19760 ( .A(n18699), .B(n18698), .Z(n18703) );
  OR U19761 ( .A(n18701), .B(n18700), .Z(n18702) );
  AND U19762 ( .A(n18703), .B(n18702), .Z(n18709) );
  XOR U19763 ( .A(n18710), .B(n18709), .Z(n18712) );
  XOR U19764 ( .A(n18711), .B(n18712), .Z(n18725) );
  XNOR U19765 ( .A(n18725), .B(sreg[1806]), .Z(n18727) );
  NANDN U19766 ( .A(n18704), .B(sreg[1805]), .Z(n18708) );
  NAND U19767 ( .A(n18706), .B(n18705), .Z(n18707) );
  NAND U19768 ( .A(n18708), .B(n18707), .Z(n18726) );
  XOR U19769 ( .A(n18727), .B(n18726), .Z(c[1806]) );
  NANDN U19770 ( .A(n18710), .B(n18709), .Z(n18714) );
  OR U19771 ( .A(n18712), .B(n18711), .Z(n18713) );
  AND U19772 ( .A(n18714), .B(n18713), .Z(n18732) );
  XOR U19773 ( .A(a[785]), .B(n2288), .Z(n18736) );
  AND U19774 ( .A(a[787]), .B(b[0]), .Z(n18716) );
  XNOR U19775 ( .A(n18716), .B(n2175), .Z(n18718) );
  NANDN U19776 ( .A(b[0]), .B(a[786]), .Z(n18717) );
  NAND U19777 ( .A(n18718), .B(n18717), .Z(n18741) );
  AND U19778 ( .A(a[783]), .B(b[3]), .Z(n18740) );
  XOR U19779 ( .A(n18741), .B(n18740), .Z(n18743) );
  XOR U19780 ( .A(n18742), .B(n18743), .Z(n18731) );
  NANDN U19781 ( .A(n18720), .B(n18719), .Z(n18724) );
  OR U19782 ( .A(n18722), .B(n18721), .Z(n18723) );
  AND U19783 ( .A(n18724), .B(n18723), .Z(n18730) );
  XOR U19784 ( .A(n18731), .B(n18730), .Z(n18733) );
  XOR U19785 ( .A(n18732), .B(n18733), .Z(n18746) );
  XNOR U19786 ( .A(n18746), .B(sreg[1807]), .Z(n18748) );
  NANDN U19787 ( .A(n18725), .B(sreg[1806]), .Z(n18729) );
  NAND U19788 ( .A(n18727), .B(n18726), .Z(n18728) );
  NAND U19789 ( .A(n18729), .B(n18728), .Z(n18747) );
  XOR U19790 ( .A(n18748), .B(n18747), .Z(c[1807]) );
  NANDN U19791 ( .A(n18731), .B(n18730), .Z(n18735) );
  OR U19792 ( .A(n18733), .B(n18732), .Z(n18734) );
  AND U19793 ( .A(n18735), .B(n18734), .Z(n18753) );
  XOR U19794 ( .A(a[786]), .B(n2288), .Z(n18757) );
  AND U19795 ( .A(a[784]), .B(b[3]), .Z(n18761) );
  AND U19796 ( .A(a[788]), .B(b[0]), .Z(n18737) );
  XNOR U19797 ( .A(n18737), .B(n2175), .Z(n18739) );
  NANDN U19798 ( .A(b[0]), .B(a[787]), .Z(n18738) );
  NAND U19799 ( .A(n18739), .B(n18738), .Z(n18762) );
  XOR U19800 ( .A(n18761), .B(n18762), .Z(n18764) );
  XOR U19801 ( .A(n18763), .B(n18764), .Z(n18752) );
  NANDN U19802 ( .A(n18741), .B(n18740), .Z(n18745) );
  OR U19803 ( .A(n18743), .B(n18742), .Z(n18744) );
  AND U19804 ( .A(n18745), .B(n18744), .Z(n18751) );
  XOR U19805 ( .A(n18752), .B(n18751), .Z(n18754) );
  XOR U19806 ( .A(n18753), .B(n18754), .Z(n18767) );
  XNOR U19807 ( .A(n18767), .B(sreg[1808]), .Z(n18769) );
  NANDN U19808 ( .A(n18746), .B(sreg[1807]), .Z(n18750) );
  NAND U19809 ( .A(n18748), .B(n18747), .Z(n18749) );
  NAND U19810 ( .A(n18750), .B(n18749), .Z(n18768) );
  XOR U19811 ( .A(n18769), .B(n18768), .Z(c[1808]) );
  NANDN U19812 ( .A(n18752), .B(n18751), .Z(n18756) );
  OR U19813 ( .A(n18754), .B(n18753), .Z(n18755) );
  AND U19814 ( .A(n18756), .B(n18755), .Z(n18774) );
  XOR U19815 ( .A(a[787]), .B(n2288), .Z(n18778) );
  AND U19816 ( .A(a[789]), .B(b[0]), .Z(n18758) );
  XNOR U19817 ( .A(n18758), .B(n2175), .Z(n18760) );
  NANDN U19818 ( .A(b[0]), .B(a[788]), .Z(n18759) );
  NAND U19819 ( .A(n18760), .B(n18759), .Z(n18783) );
  AND U19820 ( .A(a[785]), .B(b[3]), .Z(n18782) );
  XOR U19821 ( .A(n18783), .B(n18782), .Z(n18785) );
  XOR U19822 ( .A(n18784), .B(n18785), .Z(n18773) );
  NANDN U19823 ( .A(n18762), .B(n18761), .Z(n18766) );
  OR U19824 ( .A(n18764), .B(n18763), .Z(n18765) );
  AND U19825 ( .A(n18766), .B(n18765), .Z(n18772) );
  XOR U19826 ( .A(n18773), .B(n18772), .Z(n18775) );
  XOR U19827 ( .A(n18774), .B(n18775), .Z(n18788) );
  XNOR U19828 ( .A(n18788), .B(sreg[1809]), .Z(n18790) );
  NANDN U19829 ( .A(n18767), .B(sreg[1808]), .Z(n18771) );
  NAND U19830 ( .A(n18769), .B(n18768), .Z(n18770) );
  NAND U19831 ( .A(n18771), .B(n18770), .Z(n18789) );
  XOR U19832 ( .A(n18790), .B(n18789), .Z(c[1809]) );
  NANDN U19833 ( .A(n18773), .B(n18772), .Z(n18777) );
  OR U19834 ( .A(n18775), .B(n18774), .Z(n18776) );
  AND U19835 ( .A(n18777), .B(n18776), .Z(n18795) );
  XOR U19836 ( .A(a[788]), .B(n2288), .Z(n18799) );
  AND U19837 ( .A(a[790]), .B(b[0]), .Z(n18779) );
  XNOR U19838 ( .A(n18779), .B(n2175), .Z(n18781) );
  NANDN U19839 ( .A(b[0]), .B(a[789]), .Z(n18780) );
  NAND U19840 ( .A(n18781), .B(n18780), .Z(n18804) );
  AND U19841 ( .A(a[786]), .B(b[3]), .Z(n18803) );
  XOR U19842 ( .A(n18804), .B(n18803), .Z(n18806) );
  XOR U19843 ( .A(n18805), .B(n18806), .Z(n18794) );
  NANDN U19844 ( .A(n18783), .B(n18782), .Z(n18787) );
  OR U19845 ( .A(n18785), .B(n18784), .Z(n18786) );
  AND U19846 ( .A(n18787), .B(n18786), .Z(n18793) );
  XOR U19847 ( .A(n18794), .B(n18793), .Z(n18796) );
  XOR U19848 ( .A(n18795), .B(n18796), .Z(n18809) );
  XNOR U19849 ( .A(n18809), .B(sreg[1810]), .Z(n18811) );
  NANDN U19850 ( .A(n18788), .B(sreg[1809]), .Z(n18792) );
  NAND U19851 ( .A(n18790), .B(n18789), .Z(n18791) );
  NAND U19852 ( .A(n18792), .B(n18791), .Z(n18810) );
  XOR U19853 ( .A(n18811), .B(n18810), .Z(c[1810]) );
  NANDN U19854 ( .A(n18794), .B(n18793), .Z(n18798) );
  OR U19855 ( .A(n18796), .B(n18795), .Z(n18797) );
  AND U19856 ( .A(n18798), .B(n18797), .Z(n18816) );
  XOR U19857 ( .A(a[789]), .B(n2288), .Z(n18820) );
  AND U19858 ( .A(a[791]), .B(b[0]), .Z(n18800) );
  XNOR U19859 ( .A(n18800), .B(n2175), .Z(n18802) );
  NANDN U19860 ( .A(b[0]), .B(a[790]), .Z(n18801) );
  NAND U19861 ( .A(n18802), .B(n18801), .Z(n18825) );
  AND U19862 ( .A(a[787]), .B(b[3]), .Z(n18824) );
  XOR U19863 ( .A(n18825), .B(n18824), .Z(n18827) );
  XOR U19864 ( .A(n18826), .B(n18827), .Z(n18815) );
  NANDN U19865 ( .A(n18804), .B(n18803), .Z(n18808) );
  OR U19866 ( .A(n18806), .B(n18805), .Z(n18807) );
  AND U19867 ( .A(n18808), .B(n18807), .Z(n18814) );
  XOR U19868 ( .A(n18815), .B(n18814), .Z(n18817) );
  XOR U19869 ( .A(n18816), .B(n18817), .Z(n18830) );
  XNOR U19870 ( .A(n18830), .B(sreg[1811]), .Z(n18832) );
  NANDN U19871 ( .A(n18809), .B(sreg[1810]), .Z(n18813) );
  NAND U19872 ( .A(n18811), .B(n18810), .Z(n18812) );
  NAND U19873 ( .A(n18813), .B(n18812), .Z(n18831) );
  XOR U19874 ( .A(n18832), .B(n18831), .Z(c[1811]) );
  NANDN U19875 ( .A(n18815), .B(n18814), .Z(n18819) );
  OR U19876 ( .A(n18817), .B(n18816), .Z(n18818) );
  AND U19877 ( .A(n18819), .B(n18818), .Z(n18837) );
  XOR U19878 ( .A(a[790]), .B(n2289), .Z(n18841) );
  AND U19879 ( .A(a[792]), .B(b[0]), .Z(n18821) );
  XNOR U19880 ( .A(n18821), .B(n2175), .Z(n18823) );
  NANDN U19881 ( .A(b[0]), .B(a[791]), .Z(n18822) );
  NAND U19882 ( .A(n18823), .B(n18822), .Z(n18846) );
  AND U19883 ( .A(a[788]), .B(b[3]), .Z(n18845) );
  XOR U19884 ( .A(n18846), .B(n18845), .Z(n18848) );
  XOR U19885 ( .A(n18847), .B(n18848), .Z(n18836) );
  NANDN U19886 ( .A(n18825), .B(n18824), .Z(n18829) );
  OR U19887 ( .A(n18827), .B(n18826), .Z(n18828) );
  AND U19888 ( .A(n18829), .B(n18828), .Z(n18835) );
  XOR U19889 ( .A(n18836), .B(n18835), .Z(n18838) );
  XOR U19890 ( .A(n18837), .B(n18838), .Z(n18851) );
  XNOR U19891 ( .A(n18851), .B(sreg[1812]), .Z(n18853) );
  NANDN U19892 ( .A(n18830), .B(sreg[1811]), .Z(n18834) );
  NAND U19893 ( .A(n18832), .B(n18831), .Z(n18833) );
  NAND U19894 ( .A(n18834), .B(n18833), .Z(n18852) );
  XOR U19895 ( .A(n18853), .B(n18852), .Z(c[1812]) );
  NANDN U19896 ( .A(n18836), .B(n18835), .Z(n18840) );
  OR U19897 ( .A(n18838), .B(n18837), .Z(n18839) );
  AND U19898 ( .A(n18840), .B(n18839), .Z(n18858) );
  XOR U19899 ( .A(a[791]), .B(n2289), .Z(n18862) );
  AND U19900 ( .A(a[789]), .B(b[3]), .Z(n18866) );
  AND U19901 ( .A(a[793]), .B(b[0]), .Z(n18842) );
  XNOR U19902 ( .A(n18842), .B(n2175), .Z(n18844) );
  NANDN U19903 ( .A(b[0]), .B(a[792]), .Z(n18843) );
  NAND U19904 ( .A(n18844), .B(n18843), .Z(n18867) );
  XOR U19905 ( .A(n18866), .B(n18867), .Z(n18869) );
  XOR U19906 ( .A(n18868), .B(n18869), .Z(n18857) );
  NANDN U19907 ( .A(n18846), .B(n18845), .Z(n18850) );
  OR U19908 ( .A(n18848), .B(n18847), .Z(n18849) );
  AND U19909 ( .A(n18850), .B(n18849), .Z(n18856) );
  XOR U19910 ( .A(n18857), .B(n18856), .Z(n18859) );
  XOR U19911 ( .A(n18858), .B(n18859), .Z(n18872) );
  XNOR U19912 ( .A(n18872), .B(sreg[1813]), .Z(n18874) );
  NANDN U19913 ( .A(n18851), .B(sreg[1812]), .Z(n18855) );
  NAND U19914 ( .A(n18853), .B(n18852), .Z(n18854) );
  NAND U19915 ( .A(n18855), .B(n18854), .Z(n18873) );
  XOR U19916 ( .A(n18874), .B(n18873), .Z(c[1813]) );
  NANDN U19917 ( .A(n18857), .B(n18856), .Z(n18861) );
  OR U19918 ( .A(n18859), .B(n18858), .Z(n18860) );
  AND U19919 ( .A(n18861), .B(n18860), .Z(n18879) );
  XOR U19920 ( .A(a[792]), .B(n2289), .Z(n18883) );
  AND U19921 ( .A(a[794]), .B(b[0]), .Z(n18863) );
  XNOR U19922 ( .A(n18863), .B(n2175), .Z(n18865) );
  NANDN U19923 ( .A(b[0]), .B(a[793]), .Z(n18864) );
  NAND U19924 ( .A(n18865), .B(n18864), .Z(n18888) );
  AND U19925 ( .A(a[790]), .B(b[3]), .Z(n18887) );
  XOR U19926 ( .A(n18888), .B(n18887), .Z(n18890) );
  XOR U19927 ( .A(n18889), .B(n18890), .Z(n18878) );
  NANDN U19928 ( .A(n18867), .B(n18866), .Z(n18871) );
  OR U19929 ( .A(n18869), .B(n18868), .Z(n18870) );
  AND U19930 ( .A(n18871), .B(n18870), .Z(n18877) );
  XOR U19931 ( .A(n18878), .B(n18877), .Z(n18880) );
  XOR U19932 ( .A(n18879), .B(n18880), .Z(n18893) );
  XNOR U19933 ( .A(n18893), .B(sreg[1814]), .Z(n18895) );
  NANDN U19934 ( .A(n18872), .B(sreg[1813]), .Z(n18876) );
  NAND U19935 ( .A(n18874), .B(n18873), .Z(n18875) );
  NAND U19936 ( .A(n18876), .B(n18875), .Z(n18894) );
  XOR U19937 ( .A(n18895), .B(n18894), .Z(c[1814]) );
  NANDN U19938 ( .A(n18878), .B(n18877), .Z(n18882) );
  OR U19939 ( .A(n18880), .B(n18879), .Z(n18881) );
  AND U19940 ( .A(n18882), .B(n18881), .Z(n18900) );
  XOR U19941 ( .A(a[793]), .B(n2289), .Z(n18904) );
  AND U19942 ( .A(a[795]), .B(b[0]), .Z(n18884) );
  XNOR U19943 ( .A(n18884), .B(n2175), .Z(n18886) );
  NANDN U19944 ( .A(b[0]), .B(a[794]), .Z(n18885) );
  NAND U19945 ( .A(n18886), .B(n18885), .Z(n18909) );
  AND U19946 ( .A(a[791]), .B(b[3]), .Z(n18908) );
  XOR U19947 ( .A(n18909), .B(n18908), .Z(n18911) );
  XOR U19948 ( .A(n18910), .B(n18911), .Z(n18899) );
  NANDN U19949 ( .A(n18888), .B(n18887), .Z(n18892) );
  OR U19950 ( .A(n18890), .B(n18889), .Z(n18891) );
  AND U19951 ( .A(n18892), .B(n18891), .Z(n18898) );
  XOR U19952 ( .A(n18899), .B(n18898), .Z(n18901) );
  XOR U19953 ( .A(n18900), .B(n18901), .Z(n18914) );
  XNOR U19954 ( .A(n18914), .B(sreg[1815]), .Z(n18916) );
  NANDN U19955 ( .A(n18893), .B(sreg[1814]), .Z(n18897) );
  NAND U19956 ( .A(n18895), .B(n18894), .Z(n18896) );
  NAND U19957 ( .A(n18897), .B(n18896), .Z(n18915) );
  XOR U19958 ( .A(n18916), .B(n18915), .Z(c[1815]) );
  NANDN U19959 ( .A(n18899), .B(n18898), .Z(n18903) );
  OR U19960 ( .A(n18901), .B(n18900), .Z(n18902) );
  AND U19961 ( .A(n18903), .B(n18902), .Z(n18921) );
  XOR U19962 ( .A(a[794]), .B(n2289), .Z(n18925) );
  AND U19963 ( .A(a[792]), .B(b[3]), .Z(n18929) );
  AND U19964 ( .A(a[796]), .B(b[0]), .Z(n18905) );
  XNOR U19965 ( .A(n18905), .B(n2175), .Z(n18907) );
  NANDN U19966 ( .A(b[0]), .B(a[795]), .Z(n18906) );
  NAND U19967 ( .A(n18907), .B(n18906), .Z(n18930) );
  XOR U19968 ( .A(n18929), .B(n18930), .Z(n18932) );
  XOR U19969 ( .A(n18931), .B(n18932), .Z(n18920) );
  NANDN U19970 ( .A(n18909), .B(n18908), .Z(n18913) );
  OR U19971 ( .A(n18911), .B(n18910), .Z(n18912) );
  AND U19972 ( .A(n18913), .B(n18912), .Z(n18919) );
  XOR U19973 ( .A(n18920), .B(n18919), .Z(n18922) );
  XOR U19974 ( .A(n18921), .B(n18922), .Z(n18935) );
  XNOR U19975 ( .A(n18935), .B(sreg[1816]), .Z(n18937) );
  NANDN U19976 ( .A(n18914), .B(sreg[1815]), .Z(n18918) );
  NAND U19977 ( .A(n18916), .B(n18915), .Z(n18917) );
  NAND U19978 ( .A(n18918), .B(n18917), .Z(n18936) );
  XOR U19979 ( .A(n18937), .B(n18936), .Z(c[1816]) );
  NANDN U19980 ( .A(n18920), .B(n18919), .Z(n18924) );
  OR U19981 ( .A(n18922), .B(n18921), .Z(n18923) );
  AND U19982 ( .A(n18924), .B(n18923), .Z(n18942) );
  XOR U19983 ( .A(a[795]), .B(n2289), .Z(n18946) );
  AND U19984 ( .A(a[793]), .B(b[3]), .Z(n18950) );
  AND U19985 ( .A(a[797]), .B(b[0]), .Z(n18926) );
  XNOR U19986 ( .A(n18926), .B(n2175), .Z(n18928) );
  NANDN U19987 ( .A(b[0]), .B(a[796]), .Z(n18927) );
  NAND U19988 ( .A(n18928), .B(n18927), .Z(n18951) );
  XOR U19989 ( .A(n18950), .B(n18951), .Z(n18953) );
  XOR U19990 ( .A(n18952), .B(n18953), .Z(n18941) );
  NANDN U19991 ( .A(n18930), .B(n18929), .Z(n18934) );
  OR U19992 ( .A(n18932), .B(n18931), .Z(n18933) );
  AND U19993 ( .A(n18934), .B(n18933), .Z(n18940) );
  XOR U19994 ( .A(n18941), .B(n18940), .Z(n18943) );
  XOR U19995 ( .A(n18942), .B(n18943), .Z(n18956) );
  XNOR U19996 ( .A(n18956), .B(sreg[1817]), .Z(n18958) );
  NANDN U19997 ( .A(n18935), .B(sreg[1816]), .Z(n18939) );
  NAND U19998 ( .A(n18937), .B(n18936), .Z(n18938) );
  NAND U19999 ( .A(n18939), .B(n18938), .Z(n18957) );
  XOR U20000 ( .A(n18958), .B(n18957), .Z(c[1817]) );
  NANDN U20001 ( .A(n18941), .B(n18940), .Z(n18945) );
  OR U20002 ( .A(n18943), .B(n18942), .Z(n18944) );
  AND U20003 ( .A(n18945), .B(n18944), .Z(n18963) );
  XOR U20004 ( .A(a[796]), .B(n2289), .Z(n18967) );
  AND U20005 ( .A(a[794]), .B(b[3]), .Z(n18971) );
  AND U20006 ( .A(a[798]), .B(b[0]), .Z(n18947) );
  XNOR U20007 ( .A(n18947), .B(n2175), .Z(n18949) );
  NANDN U20008 ( .A(b[0]), .B(a[797]), .Z(n18948) );
  NAND U20009 ( .A(n18949), .B(n18948), .Z(n18972) );
  XOR U20010 ( .A(n18971), .B(n18972), .Z(n18974) );
  XOR U20011 ( .A(n18973), .B(n18974), .Z(n18962) );
  NANDN U20012 ( .A(n18951), .B(n18950), .Z(n18955) );
  OR U20013 ( .A(n18953), .B(n18952), .Z(n18954) );
  AND U20014 ( .A(n18955), .B(n18954), .Z(n18961) );
  XOR U20015 ( .A(n18962), .B(n18961), .Z(n18964) );
  XOR U20016 ( .A(n18963), .B(n18964), .Z(n18977) );
  XNOR U20017 ( .A(n18977), .B(sreg[1818]), .Z(n18979) );
  NANDN U20018 ( .A(n18956), .B(sreg[1817]), .Z(n18960) );
  NAND U20019 ( .A(n18958), .B(n18957), .Z(n18959) );
  NAND U20020 ( .A(n18960), .B(n18959), .Z(n18978) );
  XOR U20021 ( .A(n18979), .B(n18978), .Z(c[1818]) );
  NANDN U20022 ( .A(n18962), .B(n18961), .Z(n18966) );
  OR U20023 ( .A(n18964), .B(n18963), .Z(n18965) );
  AND U20024 ( .A(n18966), .B(n18965), .Z(n18984) );
  XOR U20025 ( .A(a[797]), .B(n2290), .Z(n18988) );
  AND U20026 ( .A(a[799]), .B(b[0]), .Z(n18968) );
  XNOR U20027 ( .A(n18968), .B(n2175), .Z(n18970) );
  NANDN U20028 ( .A(b[0]), .B(a[798]), .Z(n18969) );
  NAND U20029 ( .A(n18970), .B(n18969), .Z(n18993) );
  AND U20030 ( .A(a[795]), .B(b[3]), .Z(n18992) );
  XOR U20031 ( .A(n18993), .B(n18992), .Z(n18995) );
  XOR U20032 ( .A(n18994), .B(n18995), .Z(n18983) );
  NANDN U20033 ( .A(n18972), .B(n18971), .Z(n18976) );
  OR U20034 ( .A(n18974), .B(n18973), .Z(n18975) );
  AND U20035 ( .A(n18976), .B(n18975), .Z(n18982) );
  XOR U20036 ( .A(n18983), .B(n18982), .Z(n18985) );
  XOR U20037 ( .A(n18984), .B(n18985), .Z(n18998) );
  XNOR U20038 ( .A(n18998), .B(sreg[1819]), .Z(n19000) );
  NANDN U20039 ( .A(n18977), .B(sreg[1818]), .Z(n18981) );
  NAND U20040 ( .A(n18979), .B(n18978), .Z(n18980) );
  NAND U20041 ( .A(n18981), .B(n18980), .Z(n18999) );
  XOR U20042 ( .A(n19000), .B(n18999), .Z(c[1819]) );
  NANDN U20043 ( .A(n18983), .B(n18982), .Z(n18987) );
  OR U20044 ( .A(n18985), .B(n18984), .Z(n18986) );
  AND U20045 ( .A(n18987), .B(n18986), .Z(n19005) );
  XOR U20046 ( .A(a[798]), .B(n2290), .Z(n19009) );
  AND U20047 ( .A(a[800]), .B(b[0]), .Z(n18989) );
  XNOR U20048 ( .A(n18989), .B(n2175), .Z(n18991) );
  NANDN U20049 ( .A(b[0]), .B(a[799]), .Z(n18990) );
  NAND U20050 ( .A(n18991), .B(n18990), .Z(n19014) );
  AND U20051 ( .A(a[796]), .B(b[3]), .Z(n19013) );
  XOR U20052 ( .A(n19014), .B(n19013), .Z(n19016) );
  XOR U20053 ( .A(n19015), .B(n19016), .Z(n19004) );
  NANDN U20054 ( .A(n18993), .B(n18992), .Z(n18997) );
  OR U20055 ( .A(n18995), .B(n18994), .Z(n18996) );
  AND U20056 ( .A(n18997), .B(n18996), .Z(n19003) );
  XOR U20057 ( .A(n19004), .B(n19003), .Z(n19006) );
  XOR U20058 ( .A(n19005), .B(n19006), .Z(n19019) );
  XNOR U20059 ( .A(n19019), .B(sreg[1820]), .Z(n19021) );
  NANDN U20060 ( .A(n18998), .B(sreg[1819]), .Z(n19002) );
  NAND U20061 ( .A(n19000), .B(n18999), .Z(n19001) );
  NAND U20062 ( .A(n19002), .B(n19001), .Z(n19020) );
  XOR U20063 ( .A(n19021), .B(n19020), .Z(c[1820]) );
  NANDN U20064 ( .A(n19004), .B(n19003), .Z(n19008) );
  OR U20065 ( .A(n19006), .B(n19005), .Z(n19007) );
  AND U20066 ( .A(n19008), .B(n19007), .Z(n19026) );
  XOR U20067 ( .A(a[799]), .B(n2290), .Z(n19030) );
  AND U20068 ( .A(a[801]), .B(b[0]), .Z(n19010) );
  XNOR U20069 ( .A(n19010), .B(n2175), .Z(n19012) );
  NANDN U20070 ( .A(b[0]), .B(a[800]), .Z(n19011) );
  NAND U20071 ( .A(n19012), .B(n19011), .Z(n19035) );
  AND U20072 ( .A(a[797]), .B(b[3]), .Z(n19034) );
  XOR U20073 ( .A(n19035), .B(n19034), .Z(n19037) );
  XOR U20074 ( .A(n19036), .B(n19037), .Z(n19025) );
  NANDN U20075 ( .A(n19014), .B(n19013), .Z(n19018) );
  OR U20076 ( .A(n19016), .B(n19015), .Z(n19017) );
  AND U20077 ( .A(n19018), .B(n19017), .Z(n19024) );
  XOR U20078 ( .A(n19025), .B(n19024), .Z(n19027) );
  XOR U20079 ( .A(n19026), .B(n19027), .Z(n19040) );
  XNOR U20080 ( .A(n19040), .B(sreg[1821]), .Z(n19042) );
  NANDN U20081 ( .A(n19019), .B(sreg[1820]), .Z(n19023) );
  NAND U20082 ( .A(n19021), .B(n19020), .Z(n19022) );
  NAND U20083 ( .A(n19023), .B(n19022), .Z(n19041) );
  XOR U20084 ( .A(n19042), .B(n19041), .Z(c[1821]) );
  NANDN U20085 ( .A(n19025), .B(n19024), .Z(n19029) );
  OR U20086 ( .A(n19027), .B(n19026), .Z(n19028) );
  AND U20087 ( .A(n19029), .B(n19028), .Z(n19047) );
  XOR U20088 ( .A(a[800]), .B(n2290), .Z(n19051) );
  AND U20089 ( .A(a[798]), .B(b[3]), .Z(n19055) );
  AND U20090 ( .A(a[802]), .B(b[0]), .Z(n19031) );
  XNOR U20091 ( .A(n19031), .B(n2175), .Z(n19033) );
  NANDN U20092 ( .A(b[0]), .B(a[801]), .Z(n19032) );
  NAND U20093 ( .A(n19033), .B(n19032), .Z(n19056) );
  XOR U20094 ( .A(n19055), .B(n19056), .Z(n19058) );
  XOR U20095 ( .A(n19057), .B(n19058), .Z(n19046) );
  NANDN U20096 ( .A(n19035), .B(n19034), .Z(n19039) );
  OR U20097 ( .A(n19037), .B(n19036), .Z(n19038) );
  AND U20098 ( .A(n19039), .B(n19038), .Z(n19045) );
  XOR U20099 ( .A(n19046), .B(n19045), .Z(n19048) );
  XOR U20100 ( .A(n19047), .B(n19048), .Z(n19061) );
  XNOR U20101 ( .A(n19061), .B(sreg[1822]), .Z(n19063) );
  NANDN U20102 ( .A(n19040), .B(sreg[1821]), .Z(n19044) );
  NAND U20103 ( .A(n19042), .B(n19041), .Z(n19043) );
  NAND U20104 ( .A(n19044), .B(n19043), .Z(n19062) );
  XOR U20105 ( .A(n19063), .B(n19062), .Z(c[1822]) );
  NANDN U20106 ( .A(n19046), .B(n19045), .Z(n19050) );
  OR U20107 ( .A(n19048), .B(n19047), .Z(n19049) );
  AND U20108 ( .A(n19050), .B(n19049), .Z(n19068) );
  XOR U20109 ( .A(a[801]), .B(n2290), .Z(n19072) );
  AND U20110 ( .A(a[803]), .B(b[0]), .Z(n19052) );
  XNOR U20111 ( .A(n19052), .B(n2175), .Z(n19054) );
  NANDN U20112 ( .A(b[0]), .B(a[802]), .Z(n19053) );
  NAND U20113 ( .A(n19054), .B(n19053), .Z(n19077) );
  AND U20114 ( .A(a[799]), .B(b[3]), .Z(n19076) );
  XOR U20115 ( .A(n19077), .B(n19076), .Z(n19079) );
  XOR U20116 ( .A(n19078), .B(n19079), .Z(n19067) );
  NANDN U20117 ( .A(n19056), .B(n19055), .Z(n19060) );
  OR U20118 ( .A(n19058), .B(n19057), .Z(n19059) );
  AND U20119 ( .A(n19060), .B(n19059), .Z(n19066) );
  XOR U20120 ( .A(n19067), .B(n19066), .Z(n19069) );
  XOR U20121 ( .A(n19068), .B(n19069), .Z(n19082) );
  XNOR U20122 ( .A(n19082), .B(sreg[1823]), .Z(n19084) );
  NANDN U20123 ( .A(n19061), .B(sreg[1822]), .Z(n19065) );
  NAND U20124 ( .A(n19063), .B(n19062), .Z(n19064) );
  NAND U20125 ( .A(n19065), .B(n19064), .Z(n19083) );
  XOR U20126 ( .A(n19084), .B(n19083), .Z(c[1823]) );
  NANDN U20127 ( .A(n19067), .B(n19066), .Z(n19071) );
  OR U20128 ( .A(n19069), .B(n19068), .Z(n19070) );
  AND U20129 ( .A(n19071), .B(n19070), .Z(n19089) );
  XOR U20130 ( .A(a[802]), .B(n2290), .Z(n19093) );
  AND U20131 ( .A(a[800]), .B(b[3]), .Z(n19097) );
  AND U20132 ( .A(a[804]), .B(b[0]), .Z(n19073) );
  XNOR U20133 ( .A(n19073), .B(n2175), .Z(n19075) );
  NANDN U20134 ( .A(b[0]), .B(a[803]), .Z(n19074) );
  NAND U20135 ( .A(n19075), .B(n19074), .Z(n19098) );
  XOR U20136 ( .A(n19097), .B(n19098), .Z(n19100) );
  XOR U20137 ( .A(n19099), .B(n19100), .Z(n19088) );
  NANDN U20138 ( .A(n19077), .B(n19076), .Z(n19081) );
  OR U20139 ( .A(n19079), .B(n19078), .Z(n19080) );
  AND U20140 ( .A(n19081), .B(n19080), .Z(n19087) );
  XOR U20141 ( .A(n19088), .B(n19087), .Z(n19090) );
  XOR U20142 ( .A(n19089), .B(n19090), .Z(n19103) );
  XNOR U20143 ( .A(n19103), .B(sreg[1824]), .Z(n19105) );
  NANDN U20144 ( .A(n19082), .B(sreg[1823]), .Z(n19086) );
  NAND U20145 ( .A(n19084), .B(n19083), .Z(n19085) );
  NAND U20146 ( .A(n19086), .B(n19085), .Z(n19104) );
  XOR U20147 ( .A(n19105), .B(n19104), .Z(c[1824]) );
  NANDN U20148 ( .A(n19088), .B(n19087), .Z(n19092) );
  OR U20149 ( .A(n19090), .B(n19089), .Z(n19091) );
  AND U20150 ( .A(n19092), .B(n19091), .Z(n19110) );
  XOR U20151 ( .A(a[803]), .B(n2290), .Z(n19114) );
  AND U20152 ( .A(a[801]), .B(b[3]), .Z(n19118) );
  AND U20153 ( .A(a[805]), .B(b[0]), .Z(n19094) );
  XNOR U20154 ( .A(n19094), .B(n2175), .Z(n19096) );
  NANDN U20155 ( .A(b[0]), .B(a[804]), .Z(n19095) );
  NAND U20156 ( .A(n19096), .B(n19095), .Z(n19119) );
  XOR U20157 ( .A(n19118), .B(n19119), .Z(n19121) );
  XOR U20158 ( .A(n19120), .B(n19121), .Z(n19109) );
  NANDN U20159 ( .A(n19098), .B(n19097), .Z(n19102) );
  OR U20160 ( .A(n19100), .B(n19099), .Z(n19101) );
  AND U20161 ( .A(n19102), .B(n19101), .Z(n19108) );
  XOR U20162 ( .A(n19109), .B(n19108), .Z(n19111) );
  XOR U20163 ( .A(n19110), .B(n19111), .Z(n19124) );
  XNOR U20164 ( .A(n19124), .B(sreg[1825]), .Z(n19126) );
  NANDN U20165 ( .A(n19103), .B(sreg[1824]), .Z(n19107) );
  NAND U20166 ( .A(n19105), .B(n19104), .Z(n19106) );
  NAND U20167 ( .A(n19107), .B(n19106), .Z(n19125) );
  XOR U20168 ( .A(n19126), .B(n19125), .Z(c[1825]) );
  NANDN U20169 ( .A(n19109), .B(n19108), .Z(n19113) );
  OR U20170 ( .A(n19111), .B(n19110), .Z(n19112) );
  AND U20171 ( .A(n19113), .B(n19112), .Z(n19131) );
  XOR U20172 ( .A(a[804]), .B(n2291), .Z(n19135) );
  AND U20173 ( .A(a[806]), .B(b[0]), .Z(n19115) );
  XNOR U20174 ( .A(n19115), .B(n2175), .Z(n19117) );
  NANDN U20175 ( .A(b[0]), .B(a[805]), .Z(n19116) );
  NAND U20176 ( .A(n19117), .B(n19116), .Z(n19140) );
  AND U20177 ( .A(a[802]), .B(b[3]), .Z(n19139) );
  XOR U20178 ( .A(n19140), .B(n19139), .Z(n19142) );
  XOR U20179 ( .A(n19141), .B(n19142), .Z(n19130) );
  NANDN U20180 ( .A(n19119), .B(n19118), .Z(n19123) );
  OR U20181 ( .A(n19121), .B(n19120), .Z(n19122) );
  AND U20182 ( .A(n19123), .B(n19122), .Z(n19129) );
  XOR U20183 ( .A(n19130), .B(n19129), .Z(n19132) );
  XOR U20184 ( .A(n19131), .B(n19132), .Z(n19145) );
  XNOR U20185 ( .A(n19145), .B(sreg[1826]), .Z(n19147) );
  NANDN U20186 ( .A(n19124), .B(sreg[1825]), .Z(n19128) );
  NAND U20187 ( .A(n19126), .B(n19125), .Z(n19127) );
  NAND U20188 ( .A(n19128), .B(n19127), .Z(n19146) );
  XOR U20189 ( .A(n19147), .B(n19146), .Z(c[1826]) );
  NANDN U20190 ( .A(n19130), .B(n19129), .Z(n19134) );
  OR U20191 ( .A(n19132), .B(n19131), .Z(n19133) );
  AND U20192 ( .A(n19134), .B(n19133), .Z(n19152) );
  XOR U20193 ( .A(a[805]), .B(n2291), .Z(n19156) );
  AND U20194 ( .A(a[807]), .B(b[0]), .Z(n19136) );
  XNOR U20195 ( .A(n19136), .B(n2175), .Z(n19138) );
  NANDN U20196 ( .A(b[0]), .B(a[806]), .Z(n19137) );
  NAND U20197 ( .A(n19138), .B(n19137), .Z(n19161) );
  AND U20198 ( .A(a[803]), .B(b[3]), .Z(n19160) );
  XOR U20199 ( .A(n19161), .B(n19160), .Z(n19163) );
  XOR U20200 ( .A(n19162), .B(n19163), .Z(n19151) );
  NANDN U20201 ( .A(n19140), .B(n19139), .Z(n19144) );
  OR U20202 ( .A(n19142), .B(n19141), .Z(n19143) );
  AND U20203 ( .A(n19144), .B(n19143), .Z(n19150) );
  XOR U20204 ( .A(n19151), .B(n19150), .Z(n19153) );
  XOR U20205 ( .A(n19152), .B(n19153), .Z(n19166) );
  XNOR U20206 ( .A(n19166), .B(sreg[1827]), .Z(n19168) );
  NANDN U20207 ( .A(n19145), .B(sreg[1826]), .Z(n19149) );
  NAND U20208 ( .A(n19147), .B(n19146), .Z(n19148) );
  NAND U20209 ( .A(n19149), .B(n19148), .Z(n19167) );
  XOR U20210 ( .A(n19168), .B(n19167), .Z(c[1827]) );
  NANDN U20211 ( .A(n19151), .B(n19150), .Z(n19155) );
  OR U20212 ( .A(n19153), .B(n19152), .Z(n19154) );
  AND U20213 ( .A(n19155), .B(n19154), .Z(n19173) );
  XOR U20214 ( .A(a[806]), .B(n2291), .Z(n19177) );
  AND U20215 ( .A(a[808]), .B(b[0]), .Z(n19157) );
  XNOR U20216 ( .A(n19157), .B(n2175), .Z(n19159) );
  NANDN U20217 ( .A(b[0]), .B(a[807]), .Z(n19158) );
  NAND U20218 ( .A(n19159), .B(n19158), .Z(n19182) );
  AND U20219 ( .A(a[804]), .B(b[3]), .Z(n19181) );
  XOR U20220 ( .A(n19182), .B(n19181), .Z(n19184) );
  XOR U20221 ( .A(n19183), .B(n19184), .Z(n19172) );
  NANDN U20222 ( .A(n19161), .B(n19160), .Z(n19165) );
  OR U20223 ( .A(n19163), .B(n19162), .Z(n19164) );
  AND U20224 ( .A(n19165), .B(n19164), .Z(n19171) );
  XOR U20225 ( .A(n19172), .B(n19171), .Z(n19174) );
  XOR U20226 ( .A(n19173), .B(n19174), .Z(n19187) );
  XNOR U20227 ( .A(n19187), .B(sreg[1828]), .Z(n19189) );
  NANDN U20228 ( .A(n19166), .B(sreg[1827]), .Z(n19170) );
  NAND U20229 ( .A(n19168), .B(n19167), .Z(n19169) );
  NAND U20230 ( .A(n19170), .B(n19169), .Z(n19188) );
  XOR U20231 ( .A(n19189), .B(n19188), .Z(c[1828]) );
  NANDN U20232 ( .A(n19172), .B(n19171), .Z(n19176) );
  OR U20233 ( .A(n19174), .B(n19173), .Z(n19175) );
  AND U20234 ( .A(n19176), .B(n19175), .Z(n19194) );
  XOR U20235 ( .A(a[807]), .B(n2291), .Z(n19198) );
  AND U20236 ( .A(a[809]), .B(b[0]), .Z(n19178) );
  XNOR U20237 ( .A(n19178), .B(n2175), .Z(n19180) );
  NANDN U20238 ( .A(b[0]), .B(a[808]), .Z(n19179) );
  NAND U20239 ( .A(n19180), .B(n19179), .Z(n19203) );
  AND U20240 ( .A(a[805]), .B(b[3]), .Z(n19202) );
  XOR U20241 ( .A(n19203), .B(n19202), .Z(n19205) );
  XOR U20242 ( .A(n19204), .B(n19205), .Z(n19193) );
  NANDN U20243 ( .A(n19182), .B(n19181), .Z(n19186) );
  OR U20244 ( .A(n19184), .B(n19183), .Z(n19185) );
  AND U20245 ( .A(n19186), .B(n19185), .Z(n19192) );
  XOR U20246 ( .A(n19193), .B(n19192), .Z(n19195) );
  XOR U20247 ( .A(n19194), .B(n19195), .Z(n19208) );
  XNOR U20248 ( .A(n19208), .B(sreg[1829]), .Z(n19210) );
  NANDN U20249 ( .A(n19187), .B(sreg[1828]), .Z(n19191) );
  NAND U20250 ( .A(n19189), .B(n19188), .Z(n19190) );
  NAND U20251 ( .A(n19191), .B(n19190), .Z(n19209) );
  XOR U20252 ( .A(n19210), .B(n19209), .Z(c[1829]) );
  NANDN U20253 ( .A(n19193), .B(n19192), .Z(n19197) );
  OR U20254 ( .A(n19195), .B(n19194), .Z(n19196) );
  AND U20255 ( .A(n19197), .B(n19196), .Z(n19215) );
  XOR U20256 ( .A(a[808]), .B(n2291), .Z(n19219) );
  AND U20257 ( .A(a[806]), .B(b[3]), .Z(n19223) );
  AND U20258 ( .A(a[810]), .B(b[0]), .Z(n19199) );
  XNOR U20259 ( .A(n19199), .B(n2175), .Z(n19201) );
  NANDN U20260 ( .A(b[0]), .B(a[809]), .Z(n19200) );
  NAND U20261 ( .A(n19201), .B(n19200), .Z(n19224) );
  XOR U20262 ( .A(n19223), .B(n19224), .Z(n19226) );
  XOR U20263 ( .A(n19225), .B(n19226), .Z(n19214) );
  NANDN U20264 ( .A(n19203), .B(n19202), .Z(n19207) );
  OR U20265 ( .A(n19205), .B(n19204), .Z(n19206) );
  AND U20266 ( .A(n19207), .B(n19206), .Z(n19213) );
  XOR U20267 ( .A(n19214), .B(n19213), .Z(n19216) );
  XOR U20268 ( .A(n19215), .B(n19216), .Z(n19229) );
  XNOR U20269 ( .A(n19229), .B(sreg[1830]), .Z(n19231) );
  NANDN U20270 ( .A(n19208), .B(sreg[1829]), .Z(n19212) );
  NAND U20271 ( .A(n19210), .B(n19209), .Z(n19211) );
  NAND U20272 ( .A(n19212), .B(n19211), .Z(n19230) );
  XOR U20273 ( .A(n19231), .B(n19230), .Z(c[1830]) );
  NANDN U20274 ( .A(n19214), .B(n19213), .Z(n19218) );
  OR U20275 ( .A(n19216), .B(n19215), .Z(n19217) );
  AND U20276 ( .A(n19218), .B(n19217), .Z(n19236) );
  XOR U20277 ( .A(a[809]), .B(n2291), .Z(n19240) );
  AND U20278 ( .A(a[811]), .B(b[0]), .Z(n19220) );
  XNOR U20279 ( .A(n19220), .B(n2175), .Z(n19222) );
  NANDN U20280 ( .A(b[0]), .B(a[810]), .Z(n19221) );
  NAND U20281 ( .A(n19222), .B(n19221), .Z(n19245) );
  AND U20282 ( .A(a[807]), .B(b[3]), .Z(n19244) );
  XOR U20283 ( .A(n19245), .B(n19244), .Z(n19247) );
  XOR U20284 ( .A(n19246), .B(n19247), .Z(n19235) );
  NANDN U20285 ( .A(n19224), .B(n19223), .Z(n19228) );
  OR U20286 ( .A(n19226), .B(n19225), .Z(n19227) );
  AND U20287 ( .A(n19228), .B(n19227), .Z(n19234) );
  XOR U20288 ( .A(n19235), .B(n19234), .Z(n19237) );
  XOR U20289 ( .A(n19236), .B(n19237), .Z(n19250) );
  XNOR U20290 ( .A(n19250), .B(sreg[1831]), .Z(n19252) );
  NANDN U20291 ( .A(n19229), .B(sreg[1830]), .Z(n19233) );
  NAND U20292 ( .A(n19231), .B(n19230), .Z(n19232) );
  NAND U20293 ( .A(n19233), .B(n19232), .Z(n19251) );
  XOR U20294 ( .A(n19252), .B(n19251), .Z(c[1831]) );
  NANDN U20295 ( .A(n19235), .B(n19234), .Z(n19239) );
  OR U20296 ( .A(n19237), .B(n19236), .Z(n19238) );
  AND U20297 ( .A(n19239), .B(n19238), .Z(n19257) );
  XOR U20298 ( .A(a[810]), .B(n2291), .Z(n19261) );
  AND U20299 ( .A(a[808]), .B(b[3]), .Z(n19265) );
  AND U20300 ( .A(a[812]), .B(b[0]), .Z(n19241) );
  XNOR U20301 ( .A(n19241), .B(n2175), .Z(n19243) );
  NANDN U20302 ( .A(b[0]), .B(a[811]), .Z(n19242) );
  NAND U20303 ( .A(n19243), .B(n19242), .Z(n19266) );
  XOR U20304 ( .A(n19265), .B(n19266), .Z(n19268) );
  XOR U20305 ( .A(n19267), .B(n19268), .Z(n19256) );
  NANDN U20306 ( .A(n19245), .B(n19244), .Z(n19249) );
  OR U20307 ( .A(n19247), .B(n19246), .Z(n19248) );
  AND U20308 ( .A(n19249), .B(n19248), .Z(n19255) );
  XOR U20309 ( .A(n19256), .B(n19255), .Z(n19258) );
  XOR U20310 ( .A(n19257), .B(n19258), .Z(n19271) );
  XNOR U20311 ( .A(n19271), .B(sreg[1832]), .Z(n19273) );
  NANDN U20312 ( .A(n19250), .B(sreg[1831]), .Z(n19254) );
  NAND U20313 ( .A(n19252), .B(n19251), .Z(n19253) );
  NAND U20314 ( .A(n19254), .B(n19253), .Z(n19272) );
  XOR U20315 ( .A(n19273), .B(n19272), .Z(c[1832]) );
  NANDN U20316 ( .A(n19256), .B(n19255), .Z(n19260) );
  OR U20317 ( .A(n19258), .B(n19257), .Z(n19259) );
  AND U20318 ( .A(n19260), .B(n19259), .Z(n19278) );
  XOR U20319 ( .A(a[811]), .B(n2292), .Z(n19282) );
  AND U20320 ( .A(a[813]), .B(b[0]), .Z(n19262) );
  XNOR U20321 ( .A(n19262), .B(n2175), .Z(n19264) );
  NANDN U20322 ( .A(b[0]), .B(a[812]), .Z(n19263) );
  NAND U20323 ( .A(n19264), .B(n19263), .Z(n19287) );
  AND U20324 ( .A(a[809]), .B(b[3]), .Z(n19286) );
  XOR U20325 ( .A(n19287), .B(n19286), .Z(n19289) );
  XOR U20326 ( .A(n19288), .B(n19289), .Z(n19277) );
  NANDN U20327 ( .A(n19266), .B(n19265), .Z(n19270) );
  OR U20328 ( .A(n19268), .B(n19267), .Z(n19269) );
  AND U20329 ( .A(n19270), .B(n19269), .Z(n19276) );
  XOR U20330 ( .A(n19277), .B(n19276), .Z(n19279) );
  XOR U20331 ( .A(n19278), .B(n19279), .Z(n19292) );
  XNOR U20332 ( .A(n19292), .B(sreg[1833]), .Z(n19294) );
  NANDN U20333 ( .A(n19271), .B(sreg[1832]), .Z(n19275) );
  NAND U20334 ( .A(n19273), .B(n19272), .Z(n19274) );
  NAND U20335 ( .A(n19275), .B(n19274), .Z(n19293) );
  XOR U20336 ( .A(n19294), .B(n19293), .Z(c[1833]) );
  NANDN U20337 ( .A(n19277), .B(n19276), .Z(n19281) );
  OR U20338 ( .A(n19279), .B(n19278), .Z(n19280) );
  AND U20339 ( .A(n19281), .B(n19280), .Z(n19299) );
  XOR U20340 ( .A(a[812]), .B(n2292), .Z(n19303) );
  AND U20341 ( .A(a[814]), .B(b[0]), .Z(n19283) );
  XNOR U20342 ( .A(n19283), .B(n2175), .Z(n19285) );
  NANDN U20343 ( .A(b[0]), .B(a[813]), .Z(n19284) );
  NAND U20344 ( .A(n19285), .B(n19284), .Z(n19308) );
  AND U20345 ( .A(a[810]), .B(b[3]), .Z(n19307) );
  XOR U20346 ( .A(n19308), .B(n19307), .Z(n19310) );
  XOR U20347 ( .A(n19309), .B(n19310), .Z(n19298) );
  NANDN U20348 ( .A(n19287), .B(n19286), .Z(n19291) );
  OR U20349 ( .A(n19289), .B(n19288), .Z(n19290) );
  AND U20350 ( .A(n19291), .B(n19290), .Z(n19297) );
  XOR U20351 ( .A(n19298), .B(n19297), .Z(n19300) );
  XOR U20352 ( .A(n19299), .B(n19300), .Z(n19313) );
  XNOR U20353 ( .A(n19313), .B(sreg[1834]), .Z(n19315) );
  NANDN U20354 ( .A(n19292), .B(sreg[1833]), .Z(n19296) );
  NAND U20355 ( .A(n19294), .B(n19293), .Z(n19295) );
  NAND U20356 ( .A(n19296), .B(n19295), .Z(n19314) );
  XOR U20357 ( .A(n19315), .B(n19314), .Z(c[1834]) );
  NANDN U20358 ( .A(n19298), .B(n19297), .Z(n19302) );
  OR U20359 ( .A(n19300), .B(n19299), .Z(n19301) );
  AND U20360 ( .A(n19302), .B(n19301), .Z(n19320) );
  XOR U20361 ( .A(a[813]), .B(n2292), .Z(n19324) );
  AND U20362 ( .A(a[811]), .B(b[3]), .Z(n19328) );
  AND U20363 ( .A(a[815]), .B(b[0]), .Z(n19304) );
  XNOR U20364 ( .A(n19304), .B(n2175), .Z(n19306) );
  NANDN U20365 ( .A(b[0]), .B(a[814]), .Z(n19305) );
  NAND U20366 ( .A(n19306), .B(n19305), .Z(n19329) );
  XOR U20367 ( .A(n19328), .B(n19329), .Z(n19331) );
  XOR U20368 ( .A(n19330), .B(n19331), .Z(n19319) );
  NANDN U20369 ( .A(n19308), .B(n19307), .Z(n19312) );
  OR U20370 ( .A(n19310), .B(n19309), .Z(n19311) );
  AND U20371 ( .A(n19312), .B(n19311), .Z(n19318) );
  XOR U20372 ( .A(n19319), .B(n19318), .Z(n19321) );
  XOR U20373 ( .A(n19320), .B(n19321), .Z(n19334) );
  XNOR U20374 ( .A(n19334), .B(sreg[1835]), .Z(n19336) );
  NANDN U20375 ( .A(n19313), .B(sreg[1834]), .Z(n19317) );
  NAND U20376 ( .A(n19315), .B(n19314), .Z(n19316) );
  NAND U20377 ( .A(n19317), .B(n19316), .Z(n19335) );
  XOR U20378 ( .A(n19336), .B(n19335), .Z(c[1835]) );
  NANDN U20379 ( .A(n19319), .B(n19318), .Z(n19323) );
  OR U20380 ( .A(n19321), .B(n19320), .Z(n19322) );
  AND U20381 ( .A(n19323), .B(n19322), .Z(n19341) );
  XOR U20382 ( .A(a[814]), .B(n2292), .Z(n19345) );
  AND U20383 ( .A(a[816]), .B(b[0]), .Z(n19325) );
  XNOR U20384 ( .A(n19325), .B(n2175), .Z(n19327) );
  NANDN U20385 ( .A(b[0]), .B(a[815]), .Z(n19326) );
  NAND U20386 ( .A(n19327), .B(n19326), .Z(n19350) );
  AND U20387 ( .A(a[812]), .B(b[3]), .Z(n19349) );
  XOR U20388 ( .A(n19350), .B(n19349), .Z(n19352) );
  XOR U20389 ( .A(n19351), .B(n19352), .Z(n19340) );
  NANDN U20390 ( .A(n19329), .B(n19328), .Z(n19333) );
  OR U20391 ( .A(n19331), .B(n19330), .Z(n19332) );
  AND U20392 ( .A(n19333), .B(n19332), .Z(n19339) );
  XOR U20393 ( .A(n19340), .B(n19339), .Z(n19342) );
  XOR U20394 ( .A(n19341), .B(n19342), .Z(n19355) );
  XNOR U20395 ( .A(n19355), .B(sreg[1836]), .Z(n19357) );
  NANDN U20396 ( .A(n19334), .B(sreg[1835]), .Z(n19338) );
  NAND U20397 ( .A(n19336), .B(n19335), .Z(n19337) );
  NAND U20398 ( .A(n19338), .B(n19337), .Z(n19356) );
  XOR U20399 ( .A(n19357), .B(n19356), .Z(c[1836]) );
  NANDN U20400 ( .A(n19340), .B(n19339), .Z(n19344) );
  OR U20401 ( .A(n19342), .B(n19341), .Z(n19343) );
  AND U20402 ( .A(n19344), .B(n19343), .Z(n19362) );
  XOR U20403 ( .A(a[815]), .B(n2292), .Z(n19366) );
  AND U20404 ( .A(a[817]), .B(b[0]), .Z(n19346) );
  XNOR U20405 ( .A(n19346), .B(n2175), .Z(n19348) );
  NANDN U20406 ( .A(b[0]), .B(a[816]), .Z(n19347) );
  NAND U20407 ( .A(n19348), .B(n19347), .Z(n19371) );
  AND U20408 ( .A(a[813]), .B(b[3]), .Z(n19370) );
  XOR U20409 ( .A(n19371), .B(n19370), .Z(n19373) );
  XOR U20410 ( .A(n19372), .B(n19373), .Z(n19361) );
  NANDN U20411 ( .A(n19350), .B(n19349), .Z(n19354) );
  OR U20412 ( .A(n19352), .B(n19351), .Z(n19353) );
  AND U20413 ( .A(n19354), .B(n19353), .Z(n19360) );
  XOR U20414 ( .A(n19361), .B(n19360), .Z(n19363) );
  XOR U20415 ( .A(n19362), .B(n19363), .Z(n19376) );
  XNOR U20416 ( .A(n19376), .B(sreg[1837]), .Z(n19378) );
  NANDN U20417 ( .A(n19355), .B(sreg[1836]), .Z(n19359) );
  NAND U20418 ( .A(n19357), .B(n19356), .Z(n19358) );
  NAND U20419 ( .A(n19359), .B(n19358), .Z(n19377) );
  XOR U20420 ( .A(n19378), .B(n19377), .Z(c[1837]) );
  NANDN U20421 ( .A(n19361), .B(n19360), .Z(n19365) );
  OR U20422 ( .A(n19363), .B(n19362), .Z(n19364) );
  AND U20423 ( .A(n19365), .B(n19364), .Z(n19383) );
  XOR U20424 ( .A(a[816]), .B(n2292), .Z(n19387) );
  AND U20425 ( .A(a[818]), .B(b[0]), .Z(n19367) );
  XNOR U20426 ( .A(n19367), .B(n2175), .Z(n19369) );
  NANDN U20427 ( .A(b[0]), .B(a[817]), .Z(n19368) );
  NAND U20428 ( .A(n19369), .B(n19368), .Z(n19392) );
  AND U20429 ( .A(a[814]), .B(b[3]), .Z(n19391) );
  XOR U20430 ( .A(n19392), .B(n19391), .Z(n19394) );
  XOR U20431 ( .A(n19393), .B(n19394), .Z(n19382) );
  NANDN U20432 ( .A(n19371), .B(n19370), .Z(n19375) );
  OR U20433 ( .A(n19373), .B(n19372), .Z(n19374) );
  AND U20434 ( .A(n19375), .B(n19374), .Z(n19381) );
  XOR U20435 ( .A(n19382), .B(n19381), .Z(n19384) );
  XOR U20436 ( .A(n19383), .B(n19384), .Z(n19397) );
  XNOR U20437 ( .A(n19397), .B(sreg[1838]), .Z(n19399) );
  NANDN U20438 ( .A(n19376), .B(sreg[1837]), .Z(n19380) );
  NAND U20439 ( .A(n19378), .B(n19377), .Z(n19379) );
  NAND U20440 ( .A(n19380), .B(n19379), .Z(n19398) );
  XOR U20441 ( .A(n19399), .B(n19398), .Z(c[1838]) );
  NANDN U20442 ( .A(n19382), .B(n19381), .Z(n19386) );
  OR U20443 ( .A(n19384), .B(n19383), .Z(n19385) );
  AND U20444 ( .A(n19386), .B(n19385), .Z(n19404) );
  XOR U20445 ( .A(a[817]), .B(n2292), .Z(n19408) );
  AND U20446 ( .A(a[815]), .B(b[3]), .Z(n19412) );
  AND U20447 ( .A(a[819]), .B(b[0]), .Z(n19388) );
  XNOR U20448 ( .A(n19388), .B(n2175), .Z(n19390) );
  NANDN U20449 ( .A(b[0]), .B(a[818]), .Z(n19389) );
  NAND U20450 ( .A(n19390), .B(n19389), .Z(n19413) );
  XOR U20451 ( .A(n19412), .B(n19413), .Z(n19415) );
  XOR U20452 ( .A(n19414), .B(n19415), .Z(n19403) );
  NANDN U20453 ( .A(n19392), .B(n19391), .Z(n19396) );
  OR U20454 ( .A(n19394), .B(n19393), .Z(n19395) );
  AND U20455 ( .A(n19396), .B(n19395), .Z(n19402) );
  XOR U20456 ( .A(n19403), .B(n19402), .Z(n19405) );
  XOR U20457 ( .A(n19404), .B(n19405), .Z(n19418) );
  XNOR U20458 ( .A(n19418), .B(sreg[1839]), .Z(n19420) );
  NANDN U20459 ( .A(n19397), .B(sreg[1838]), .Z(n19401) );
  NAND U20460 ( .A(n19399), .B(n19398), .Z(n19400) );
  NAND U20461 ( .A(n19401), .B(n19400), .Z(n19419) );
  XOR U20462 ( .A(n19420), .B(n19419), .Z(c[1839]) );
  NANDN U20463 ( .A(n19403), .B(n19402), .Z(n19407) );
  OR U20464 ( .A(n19405), .B(n19404), .Z(n19406) );
  AND U20465 ( .A(n19407), .B(n19406), .Z(n19425) );
  XOR U20466 ( .A(a[818]), .B(n2293), .Z(n19429) );
  AND U20467 ( .A(a[820]), .B(b[0]), .Z(n19409) );
  XNOR U20468 ( .A(n19409), .B(n2175), .Z(n19411) );
  NANDN U20469 ( .A(b[0]), .B(a[819]), .Z(n19410) );
  NAND U20470 ( .A(n19411), .B(n19410), .Z(n19434) );
  AND U20471 ( .A(a[816]), .B(b[3]), .Z(n19433) );
  XOR U20472 ( .A(n19434), .B(n19433), .Z(n19436) );
  XOR U20473 ( .A(n19435), .B(n19436), .Z(n19424) );
  NANDN U20474 ( .A(n19413), .B(n19412), .Z(n19417) );
  OR U20475 ( .A(n19415), .B(n19414), .Z(n19416) );
  AND U20476 ( .A(n19417), .B(n19416), .Z(n19423) );
  XOR U20477 ( .A(n19424), .B(n19423), .Z(n19426) );
  XOR U20478 ( .A(n19425), .B(n19426), .Z(n19439) );
  XNOR U20479 ( .A(n19439), .B(sreg[1840]), .Z(n19441) );
  NANDN U20480 ( .A(n19418), .B(sreg[1839]), .Z(n19422) );
  NAND U20481 ( .A(n19420), .B(n19419), .Z(n19421) );
  NAND U20482 ( .A(n19422), .B(n19421), .Z(n19440) );
  XOR U20483 ( .A(n19441), .B(n19440), .Z(c[1840]) );
  NANDN U20484 ( .A(n19424), .B(n19423), .Z(n19428) );
  OR U20485 ( .A(n19426), .B(n19425), .Z(n19427) );
  AND U20486 ( .A(n19428), .B(n19427), .Z(n19446) );
  XOR U20487 ( .A(a[819]), .B(n2293), .Z(n19450) );
  AND U20488 ( .A(a[817]), .B(b[3]), .Z(n19454) );
  AND U20489 ( .A(a[821]), .B(b[0]), .Z(n19430) );
  XNOR U20490 ( .A(n19430), .B(n2175), .Z(n19432) );
  NANDN U20491 ( .A(b[0]), .B(a[820]), .Z(n19431) );
  NAND U20492 ( .A(n19432), .B(n19431), .Z(n19455) );
  XOR U20493 ( .A(n19454), .B(n19455), .Z(n19457) );
  XOR U20494 ( .A(n19456), .B(n19457), .Z(n19445) );
  NANDN U20495 ( .A(n19434), .B(n19433), .Z(n19438) );
  OR U20496 ( .A(n19436), .B(n19435), .Z(n19437) );
  AND U20497 ( .A(n19438), .B(n19437), .Z(n19444) );
  XOR U20498 ( .A(n19445), .B(n19444), .Z(n19447) );
  XOR U20499 ( .A(n19446), .B(n19447), .Z(n19460) );
  XNOR U20500 ( .A(n19460), .B(sreg[1841]), .Z(n19462) );
  NANDN U20501 ( .A(n19439), .B(sreg[1840]), .Z(n19443) );
  NAND U20502 ( .A(n19441), .B(n19440), .Z(n19442) );
  NAND U20503 ( .A(n19443), .B(n19442), .Z(n19461) );
  XOR U20504 ( .A(n19462), .B(n19461), .Z(c[1841]) );
  NANDN U20505 ( .A(n19445), .B(n19444), .Z(n19449) );
  OR U20506 ( .A(n19447), .B(n19446), .Z(n19448) );
  AND U20507 ( .A(n19449), .B(n19448), .Z(n19467) );
  XOR U20508 ( .A(a[820]), .B(n2293), .Z(n19471) );
  AND U20509 ( .A(a[822]), .B(b[0]), .Z(n19451) );
  XNOR U20510 ( .A(n19451), .B(n2175), .Z(n19453) );
  NANDN U20511 ( .A(b[0]), .B(a[821]), .Z(n19452) );
  NAND U20512 ( .A(n19453), .B(n19452), .Z(n19476) );
  AND U20513 ( .A(a[818]), .B(b[3]), .Z(n19475) );
  XOR U20514 ( .A(n19476), .B(n19475), .Z(n19478) );
  XOR U20515 ( .A(n19477), .B(n19478), .Z(n19466) );
  NANDN U20516 ( .A(n19455), .B(n19454), .Z(n19459) );
  OR U20517 ( .A(n19457), .B(n19456), .Z(n19458) );
  AND U20518 ( .A(n19459), .B(n19458), .Z(n19465) );
  XOR U20519 ( .A(n19466), .B(n19465), .Z(n19468) );
  XOR U20520 ( .A(n19467), .B(n19468), .Z(n19481) );
  XNOR U20521 ( .A(n19481), .B(sreg[1842]), .Z(n19483) );
  NANDN U20522 ( .A(n19460), .B(sreg[1841]), .Z(n19464) );
  NAND U20523 ( .A(n19462), .B(n19461), .Z(n19463) );
  NAND U20524 ( .A(n19464), .B(n19463), .Z(n19482) );
  XOR U20525 ( .A(n19483), .B(n19482), .Z(c[1842]) );
  NANDN U20526 ( .A(n19466), .B(n19465), .Z(n19470) );
  OR U20527 ( .A(n19468), .B(n19467), .Z(n19469) );
  AND U20528 ( .A(n19470), .B(n19469), .Z(n19488) );
  XOR U20529 ( .A(a[821]), .B(n2293), .Z(n19492) );
  AND U20530 ( .A(a[819]), .B(b[3]), .Z(n19496) );
  AND U20531 ( .A(a[823]), .B(b[0]), .Z(n19472) );
  XNOR U20532 ( .A(n19472), .B(n2175), .Z(n19474) );
  NANDN U20533 ( .A(b[0]), .B(a[822]), .Z(n19473) );
  NAND U20534 ( .A(n19474), .B(n19473), .Z(n19497) );
  XOR U20535 ( .A(n19496), .B(n19497), .Z(n19499) );
  XOR U20536 ( .A(n19498), .B(n19499), .Z(n19487) );
  NANDN U20537 ( .A(n19476), .B(n19475), .Z(n19480) );
  OR U20538 ( .A(n19478), .B(n19477), .Z(n19479) );
  AND U20539 ( .A(n19480), .B(n19479), .Z(n19486) );
  XOR U20540 ( .A(n19487), .B(n19486), .Z(n19489) );
  XOR U20541 ( .A(n19488), .B(n19489), .Z(n19502) );
  XNOR U20542 ( .A(n19502), .B(sreg[1843]), .Z(n19504) );
  NANDN U20543 ( .A(n19481), .B(sreg[1842]), .Z(n19485) );
  NAND U20544 ( .A(n19483), .B(n19482), .Z(n19484) );
  NAND U20545 ( .A(n19485), .B(n19484), .Z(n19503) );
  XOR U20546 ( .A(n19504), .B(n19503), .Z(c[1843]) );
  NANDN U20547 ( .A(n19487), .B(n19486), .Z(n19491) );
  OR U20548 ( .A(n19489), .B(n19488), .Z(n19490) );
  AND U20549 ( .A(n19491), .B(n19490), .Z(n19509) );
  XOR U20550 ( .A(a[822]), .B(n2293), .Z(n19513) );
  AND U20551 ( .A(a[824]), .B(b[0]), .Z(n19493) );
  XNOR U20552 ( .A(n19493), .B(n2175), .Z(n19495) );
  NANDN U20553 ( .A(b[0]), .B(a[823]), .Z(n19494) );
  NAND U20554 ( .A(n19495), .B(n19494), .Z(n19518) );
  AND U20555 ( .A(a[820]), .B(b[3]), .Z(n19517) );
  XOR U20556 ( .A(n19518), .B(n19517), .Z(n19520) );
  XOR U20557 ( .A(n19519), .B(n19520), .Z(n19508) );
  NANDN U20558 ( .A(n19497), .B(n19496), .Z(n19501) );
  OR U20559 ( .A(n19499), .B(n19498), .Z(n19500) );
  AND U20560 ( .A(n19501), .B(n19500), .Z(n19507) );
  XOR U20561 ( .A(n19508), .B(n19507), .Z(n19510) );
  XOR U20562 ( .A(n19509), .B(n19510), .Z(n19523) );
  XNOR U20563 ( .A(n19523), .B(sreg[1844]), .Z(n19525) );
  NANDN U20564 ( .A(n19502), .B(sreg[1843]), .Z(n19506) );
  NAND U20565 ( .A(n19504), .B(n19503), .Z(n19505) );
  NAND U20566 ( .A(n19506), .B(n19505), .Z(n19524) );
  XOR U20567 ( .A(n19525), .B(n19524), .Z(c[1844]) );
  NANDN U20568 ( .A(n19508), .B(n19507), .Z(n19512) );
  OR U20569 ( .A(n19510), .B(n19509), .Z(n19511) );
  AND U20570 ( .A(n19512), .B(n19511), .Z(n19530) );
  XOR U20571 ( .A(a[823]), .B(n2293), .Z(n19534) );
  AND U20572 ( .A(a[821]), .B(b[3]), .Z(n19538) );
  AND U20573 ( .A(a[825]), .B(b[0]), .Z(n19514) );
  XNOR U20574 ( .A(n19514), .B(n2175), .Z(n19516) );
  NANDN U20575 ( .A(b[0]), .B(a[824]), .Z(n19515) );
  NAND U20576 ( .A(n19516), .B(n19515), .Z(n19539) );
  XOR U20577 ( .A(n19538), .B(n19539), .Z(n19541) );
  XOR U20578 ( .A(n19540), .B(n19541), .Z(n19529) );
  NANDN U20579 ( .A(n19518), .B(n19517), .Z(n19522) );
  OR U20580 ( .A(n19520), .B(n19519), .Z(n19521) );
  AND U20581 ( .A(n19522), .B(n19521), .Z(n19528) );
  XOR U20582 ( .A(n19529), .B(n19528), .Z(n19531) );
  XOR U20583 ( .A(n19530), .B(n19531), .Z(n19544) );
  XNOR U20584 ( .A(n19544), .B(sreg[1845]), .Z(n19546) );
  NANDN U20585 ( .A(n19523), .B(sreg[1844]), .Z(n19527) );
  NAND U20586 ( .A(n19525), .B(n19524), .Z(n19526) );
  NAND U20587 ( .A(n19527), .B(n19526), .Z(n19545) );
  XOR U20588 ( .A(n19546), .B(n19545), .Z(c[1845]) );
  NANDN U20589 ( .A(n19529), .B(n19528), .Z(n19533) );
  OR U20590 ( .A(n19531), .B(n19530), .Z(n19532) );
  AND U20591 ( .A(n19533), .B(n19532), .Z(n19551) );
  XOR U20592 ( .A(a[824]), .B(n2293), .Z(n19555) );
  AND U20593 ( .A(a[826]), .B(b[0]), .Z(n19535) );
  XNOR U20594 ( .A(n19535), .B(n2175), .Z(n19537) );
  NANDN U20595 ( .A(b[0]), .B(a[825]), .Z(n19536) );
  NAND U20596 ( .A(n19537), .B(n19536), .Z(n19560) );
  AND U20597 ( .A(a[822]), .B(b[3]), .Z(n19559) );
  XOR U20598 ( .A(n19560), .B(n19559), .Z(n19562) );
  XOR U20599 ( .A(n19561), .B(n19562), .Z(n19550) );
  NANDN U20600 ( .A(n19539), .B(n19538), .Z(n19543) );
  OR U20601 ( .A(n19541), .B(n19540), .Z(n19542) );
  AND U20602 ( .A(n19543), .B(n19542), .Z(n19549) );
  XOR U20603 ( .A(n19550), .B(n19549), .Z(n19552) );
  XOR U20604 ( .A(n19551), .B(n19552), .Z(n19565) );
  XNOR U20605 ( .A(n19565), .B(sreg[1846]), .Z(n19567) );
  NANDN U20606 ( .A(n19544), .B(sreg[1845]), .Z(n19548) );
  NAND U20607 ( .A(n19546), .B(n19545), .Z(n19547) );
  NAND U20608 ( .A(n19548), .B(n19547), .Z(n19566) );
  XOR U20609 ( .A(n19567), .B(n19566), .Z(c[1846]) );
  NANDN U20610 ( .A(n19550), .B(n19549), .Z(n19554) );
  OR U20611 ( .A(n19552), .B(n19551), .Z(n19553) );
  AND U20612 ( .A(n19554), .B(n19553), .Z(n19572) );
  XOR U20613 ( .A(a[825]), .B(n2294), .Z(n19576) );
  AND U20614 ( .A(a[823]), .B(b[3]), .Z(n19580) );
  AND U20615 ( .A(a[827]), .B(b[0]), .Z(n19556) );
  XNOR U20616 ( .A(n19556), .B(n2175), .Z(n19558) );
  NANDN U20617 ( .A(b[0]), .B(a[826]), .Z(n19557) );
  NAND U20618 ( .A(n19558), .B(n19557), .Z(n19581) );
  XOR U20619 ( .A(n19580), .B(n19581), .Z(n19583) );
  XOR U20620 ( .A(n19582), .B(n19583), .Z(n19571) );
  NANDN U20621 ( .A(n19560), .B(n19559), .Z(n19564) );
  OR U20622 ( .A(n19562), .B(n19561), .Z(n19563) );
  AND U20623 ( .A(n19564), .B(n19563), .Z(n19570) );
  XOR U20624 ( .A(n19571), .B(n19570), .Z(n19573) );
  XOR U20625 ( .A(n19572), .B(n19573), .Z(n19586) );
  XNOR U20626 ( .A(n19586), .B(sreg[1847]), .Z(n19588) );
  NANDN U20627 ( .A(n19565), .B(sreg[1846]), .Z(n19569) );
  NAND U20628 ( .A(n19567), .B(n19566), .Z(n19568) );
  NAND U20629 ( .A(n19569), .B(n19568), .Z(n19587) );
  XOR U20630 ( .A(n19588), .B(n19587), .Z(c[1847]) );
  NANDN U20631 ( .A(n19571), .B(n19570), .Z(n19575) );
  OR U20632 ( .A(n19573), .B(n19572), .Z(n19574) );
  AND U20633 ( .A(n19575), .B(n19574), .Z(n19593) );
  XOR U20634 ( .A(a[826]), .B(n2294), .Z(n19597) );
  AND U20635 ( .A(a[828]), .B(b[0]), .Z(n19577) );
  XNOR U20636 ( .A(n19577), .B(n2175), .Z(n19579) );
  NANDN U20637 ( .A(b[0]), .B(a[827]), .Z(n19578) );
  NAND U20638 ( .A(n19579), .B(n19578), .Z(n19602) );
  AND U20639 ( .A(a[824]), .B(b[3]), .Z(n19601) );
  XOR U20640 ( .A(n19602), .B(n19601), .Z(n19604) );
  XOR U20641 ( .A(n19603), .B(n19604), .Z(n19592) );
  NANDN U20642 ( .A(n19581), .B(n19580), .Z(n19585) );
  OR U20643 ( .A(n19583), .B(n19582), .Z(n19584) );
  AND U20644 ( .A(n19585), .B(n19584), .Z(n19591) );
  XOR U20645 ( .A(n19592), .B(n19591), .Z(n19594) );
  XOR U20646 ( .A(n19593), .B(n19594), .Z(n19607) );
  XNOR U20647 ( .A(n19607), .B(sreg[1848]), .Z(n19609) );
  NANDN U20648 ( .A(n19586), .B(sreg[1847]), .Z(n19590) );
  NAND U20649 ( .A(n19588), .B(n19587), .Z(n19589) );
  NAND U20650 ( .A(n19590), .B(n19589), .Z(n19608) );
  XOR U20651 ( .A(n19609), .B(n19608), .Z(c[1848]) );
  NANDN U20652 ( .A(n19592), .B(n19591), .Z(n19596) );
  OR U20653 ( .A(n19594), .B(n19593), .Z(n19595) );
  AND U20654 ( .A(n19596), .B(n19595), .Z(n19614) );
  XOR U20655 ( .A(a[827]), .B(n2294), .Z(n19618) );
  AND U20656 ( .A(a[829]), .B(b[0]), .Z(n19598) );
  XNOR U20657 ( .A(n19598), .B(n2175), .Z(n19600) );
  NANDN U20658 ( .A(b[0]), .B(a[828]), .Z(n19599) );
  NAND U20659 ( .A(n19600), .B(n19599), .Z(n19623) );
  AND U20660 ( .A(a[825]), .B(b[3]), .Z(n19622) );
  XOR U20661 ( .A(n19623), .B(n19622), .Z(n19625) );
  XOR U20662 ( .A(n19624), .B(n19625), .Z(n19613) );
  NANDN U20663 ( .A(n19602), .B(n19601), .Z(n19606) );
  OR U20664 ( .A(n19604), .B(n19603), .Z(n19605) );
  AND U20665 ( .A(n19606), .B(n19605), .Z(n19612) );
  XOR U20666 ( .A(n19613), .B(n19612), .Z(n19615) );
  XOR U20667 ( .A(n19614), .B(n19615), .Z(n19628) );
  XNOR U20668 ( .A(n19628), .B(sreg[1849]), .Z(n19630) );
  NANDN U20669 ( .A(n19607), .B(sreg[1848]), .Z(n19611) );
  NAND U20670 ( .A(n19609), .B(n19608), .Z(n19610) );
  NAND U20671 ( .A(n19611), .B(n19610), .Z(n19629) );
  XOR U20672 ( .A(n19630), .B(n19629), .Z(c[1849]) );
  NANDN U20673 ( .A(n19613), .B(n19612), .Z(n19617) );
  OR U20674 ( .A(n19615), .B(n19614), .Z(n19616) );
  AND U20675 ( .A(n19617), .B(n19616), .Z(n19635) );
  XOR U20676 ( .A(a[828]), .B(n2294), .Z(n19639) );
  AND U20677 ( .A(a[830]), .B(b[0]), .Z(n19619) );
  XNOR U20678 ( .A(n19619), .B(n2175), .Z(n19621) );
  NANDN U20679 ( .A(b[0]), .B(a[829]), .Z(n19620) );
  NAND U20680 ( .A(n19621), .B(n19620), .Z(n19644) );
  AND U20681 ( .A(a[826]), .B(b[3]), .Z(n19643) );
  XOR U20682 ( .A(n19644), .B(n19643), .Z(n19646) );
  XOR U20683 ( .A(n19645), .B(n19646), .Z(n19634) );
  NANDN U20684 ( .A(n19623), .B(n19622), .Z(n19627) );
  OR U20685 ( .A(n19625), .B(n19624), .Z(n19626) );
  AND U20686 ( .A(n19627), .B(n19626), .Z(n19633) );
  XOR U20687 ( .A(n19634), .B(n19633), .Z(n19636) );
  XOR U20688 ( .A(n19635), .B(n19636), .Z(n19649) );
  XNOR U20689 ( .A(n19649), .B(sreg[1850]), .Z(n19651) );
  NANDN U20690 ( .A(n19628), .B(sreg[1849]), .Z(n19632) );
  NAND U20691 ( .A(n19630), .B(n19629), .Z(n19631) );
  NAND U20692 ( .A(n19632), .B(n19631), .Z(n19650) );
  XOR U20693 ( .A(n19651), .B(n19650), .Z(c[1850]) );
  NANDN U20694 ( .A(n19634), .B(n19633), .Z(n19638) );
  OR U20695 ( .A(n19636), .B(n19635), .Z(n19637) );
  AND U20696 ( .A(n19638), .B(n19637), .Z(n19656) );
  XOR U20697 ( .A(a[829]), .B(n2294), .Z(n19660) );
  AND U20698 ( .A(a[827]), .B(b[3]), .Z(n19664) );
  AND U20699 ( .A(a[831]), .B(b[0]), .Z(n19640) );
  XNOR U20700 ( .A(n19640), .B(n2175), .Z(n19642) );
  NANDN U20701 ( .A(b[0]), .B(a[830]), .Z(n19641) );
  NAND U20702 ( .A(n19642), .B(n19641), .Z(n19665) );
  XOR U20703 ( .A(n19664), .B(n19665), .Z(n19667) );
  XOR U20704 ( .A(n19666), .B(n19667), .Z(n19655) );
  NANDN U20705 ( .A(n19644), .B(n19643), .Z(n19648) );
  OR U20706 ( .A(n19646), .B(n19645), .Z(n19647) );
  AND U20707 ( .A(n19648), .B(n19647), .Z(n19654) );
  XOR U20708 ( .A(n19655), .B(n19654), .Z(n19657) );
  XOR U20709 ( .A(n19656), .B(n19657), .Z(n19670) );
  XNOR U20710 ( .A(n19670), .B(sreg[1851]), .Z(n19672) );
  NANDN U20711 ( .A(n19649), .B(sreg[1850]), .Z(n19653) );
  NAND U20712 ( .A(n19651), .B(n19650), .Z(n19652) );
  NAND U20713 ( .A(n19653), .B(n19652), .Z(n19671) );
  XOR U20714 ( .A(n19672), .B(n19671), .Z(c[1851]) );
  NANDN U20715 ( .A(n19655), .B(n19654), .Z(n19659) );
  OR U20716 ( .A(n19657), .B(n19656), .Z(n19658) );
  AND U20717 ( .A(n19659), .B(n19658), .Z(n19677) );
  XOR U20718 ( .A(a[830]), .B(n2294), .Z(n19681) );
  AND U20719 ( .A(a[832]), .B(b[0]), .Z(n19661) );
  XNOR U20720 ( .A(n19661), .B(n2175), .Z(n19663) );
  NANDN U20721 ( .A(b[0]), .B(a[831]), .Z(n19662) );
  NAND U20722 ( .A(n19663), .B(n19662), .Z(n19686) );
  AND U20723 ( .A(a[828]), .B(b[3]), .Z(n19685) );
  XOR U20724 ( .A(n19686), .B(n19685), .Z(n19688) );
  XOR U20725 ( .A(n19687), .B(n19688), .Z(n19676) );
  NANDN U20726 ( .A(n19665), .B(n19664), .Z(n19669) );
  OR U20727 ( .A(n19667), .B(n19666), .Z(n19668) );
  AND U20728 ( .A(n19669), .B(n19668), .Z(n19675) );
  XOR U20729 ( .A(n19676), .B(n19675), .Z(n19678) );
  XOR U20730 ( .A(n19677), .B(n19678), .Z(n19691) );
  XNOR U20731 ( .A(n19691), .B(sreg[1852]), .Z(n19693) );
  NANDN U20732 ( .A(n19670), .B(sreg[1851]), .Z(n19674) );
  NAND U20733 ( .A(n19672), .B(n19671), .Z(n19673) );
  NAND U20734 ( .A(n19674), .B(n19673), .Z(n19692) );
  XOR U20735 ( .A(n19693), .B(n19692), .Z(c[1852]) );
  NANDN U20736 ( .A(n19676), .B(n19675), .Z(n19680) );
  OR U20737 ( .A(n19678), .B(n19677), .Z(n19679) );
  AND U20738 ( .A(n19680), .B(n19679), .Z(n19699) );
  XOR U20739 ( .A(a[831]), .B(n2294), .Z(n19700) );
  AND U20740 ( .A(b[0]), .B(a[833]), .Z(n19682) );
  XOR U20741 ( .A(b[1]), .B(n19682), .Z(n19684) );
  NAND U20742 ( .A(n23588), .B(a[832]), .Z(n19683) );
  AND U20743 ( .A(n19684), .B(n19683), .Z(n19704) );
  AND U20744 ( .A(a[829]), .B(b[3]), .Z(n19705) );
  XOR U20745 ( .A(n19704), .B(n19705), .Z(n19706) );
  XNOR U20746 ( .A(n19707), .B(n19706), .Z(n19696) );
  NANDN U20747 ( .A(n19686), .B(n19685), .Z(n19690) );
  OR U20748 ( .A(n19688), .B(n19687), .Z(n19689) );
  AND U20749 ( .A(n19690), .B(n19689), .Z(n19697) );
  XNOR U20750 ( .A(n19696), .B(n19697), .Z(n19698) );
  XNOR U20751 ( .A(n19699), .B(n19698), .Z(n19710) );
  XNOR U20752 ( .A(n19710), .B(sreg[1853]), .Z(n19712) );
  NANDN U20753 ( .A(n19691), .B(sreg[1852]), .Z(n19695) );
  NAND U20754 ( .A(n19693), .B(n19692), .Z(n19694) );
  NAND U20755 ( .A(n19695), .B(n19694), .Z(n19711) );
  XOR U20756 ( .A(n19712), .B(n19711), .Z(c[1853]) );
  XOR U20757 ( .A(a[832]), .B(n2295), .Z(n19719) );
  AND U20758 ( .A(a[834]), .B(b[0]), .Z(n19701) );
  XNOR U20759 ( .A(n19701), .B(n2175), .Z(n19703) );
  NANDN U20760 ( .A(b[0]), .B(a[833]), .Z(n19702) );
  NAND U20761 ( .A(n19703), .B(n19702), .Z(n19724) );
  AND U20762 ( .A(a[830]), .B(b[3]), .Z(n19723) );
  XOR U20763 ( .A(n19724), .B(n19723), .Z(n19726) );
  XOR U20764 ( .A(n19725), .B(n19726), .Z(n19714) );
  NAND U20765 ( .A(n19705), .B(n19704), .Z(n19709) );
  NANDN U20766 ( .A(n19707), .B(n19706), .Z(n19708) );
  AND U20767 ( .A(n19709), .B(n19708), .Z(n19713) );
  XOR U20768 ( .A(n19714), .B(n19713), .Z(n19716) );
  XOR U20769 ( .A(n19715), .B(n19716), .Z(n19729) );
  XNOR U20770 ( .A(n19729), .B(sreg[1854]), .Z(n19731) );
  XOR U20771 ( .A(n19731), .B(n19730), .Z(c[1854]) );
  NANDN U20772 ( .A(n19714), .B(n19713), .Z(n19718) );
  OR U20773 ( .A(n19716), .B(n19715), .Z(n19717) );
  AND U20774 ( .A(n19718), .B(n19717), .Z(n19736) );
  XOR U20775 ( .A(a[833]), .B(n2295), .Z(n19740) );
  AND U20776 ( .A(a[831]), .B(b[3]), .Z(n19744) );
  AND U20777 ( .A(a[835]), .B(b[0]), .Z(n19720) );
  XNOR U20778 ( .A(n19720), .B(n2175), .Z(n19722) );
  NANDN U20779 ( .A(b[0]), .B(a[834]), .Z(n19721) );
  NAND U20780 ( .A(n19722), .B(n19721), .Z(n19745) );
  XOR U20781 ( .A(n19744), .B(n19745), .Z(n19747) );
  XOR U20782 ( .A(n19746), .B(n19747), .Z(n19735) );
  NANDN U20783 ( .A(n19724), .B(n19723), .Z(n19728) );
  OR U20784 ( .A(n19726), .B(n19725), .Z(n19727) );
  AND U20785 ( .A(n19728), .B(n19727), .Z(n19734) );
  XOR U20786 ( .A(n19735), .B(n19734), .Z(n19737) );
  XOR U20787 ( .A(n19736), .B(n19737), .Z(n19750) );
  XNOR U20788 ( .A(n19750), .B(sreg[1855]), .Z(n19752) );
  NANDN U20789 ( .A(n19729), .B(sreg[1854]), .Z(n19733) );
  NAND U20790 ( .A(n19731), .B(n19730), .Z(n19732) );
  NAND U20791 ( .A(n19733), .B(n19732), .Z(n19751) );
  XOR U20792 ( .A(n19752), .B(n19751), .Z(c[1855]) );
  NANDN U20793 ( .A(n19735), .B(n19734), .Z(n19739) );
  OR U20794 ( .A(n19737), .B(n19736), .Z(n19738) );
  AND U20795 ( .A(n19739), .B(n19738), .Z(n19757) );
  XOR U20796 ( .A(a[834]), .B(n2295), .Z(n19761) );
  AND U20797 ( .A(a[836]), .B(b[0]), .Z(n19741) );
  XNOR U20798 ( .A(n19741), .B(n2175), .Z(n19743) );
  NANDN U20799 ( .A(b[0]), .B(a[835]), .Z(n19742) );
  NAND U20800 ( .A(n19743), .B(n19742), .Z(n19766) );
  AND U20801 ( .A(a[832]), .B(b[3]), .Z(n19765) );
  XOR U20802 ( .A(n19766), .B(n19765), .Z(n19768) );
  XOR U20803 ( .A(n19767), .B(n19768), .Z(n19756) );
  NANDN U20804 ( .A(n19745), .B(n19744), .Z(n19749) );
  OR U20805 ( .A(n19747), .B(n19746), .Z(n19748) );
  AND U20806 ( .A(n19749), .B(n19748), .Z(n19755) );
  XOR U20807 ( .A(n19756), .B(n19755), .Z(n19758) );
  XOR U20808 ( .A(n19757), .B(n19758), .Z(n19771) );
  XNOR U20809 ( .A(n19771), .B(sreg[1856]), .Z(n19773) );
  NANDN U20810 ( .A(n19750), .B(sreg[1855]), .Z(n19754) );
  NAND U20811 ( .A(n19752), .B(n19751), .Z(n19753) );
  NAND U20812 ( .A(n19754), .B(n19753), .Z(n19772) );
  XOR U20813 ( .A(n19773), .B(n19772), .Z(c[1856]) );
  NANDN U20814 ( .A(n19756), .B(n19755), .Z(n19760) );
  OR U20815 ( .A(n19758), .B(n19757), .Z(n19759) );
  AND U20816 ( .A(n19760), .B(n19759), .Z(n19778) );
  XOR U20817 ( .A(a[835]), .B(n2295), .Z(n19782) );
  AND U20818 ( .A(a[837]), .B(b[0]), .Z(n19762) );
  XNOR U20819 ( .A(n19762), .B(n2175), .Z(n19764) );
  NANDN U20820 ( .A(b[0]), .B(a[836]), .Z(n19763) );
  NAND U20821 ( .A(n19764), .B(n19763), .Z(n19787) );
  AND U20822 ( .A(a[833]), .B(b[3]), .Z(n19786) );
  XOR U20823 ( .A(n19787), .B(n19786), .Z(n19789) );
  XOR U20824 ( .A(n19788), .B(n19789), .Z(n19777) );
  NANDN U20825 ( .A(n19766), .B(n19765), .Z(n19770) );
  OR U20826 ( .A(n19768), .B(n19767), .Z(n19769) );
  AND U20827 ( .A(n19770), .B(n19769), .Z(n19776) );
  XOR U20828 ( .A(n19777), .B(n19776), .Z(n19779) );
  XOR U20829 ( .A(n19778), .B(n19779), .Z(n19792) );
  XNOR U20830 ( .A(n19792), .B(sreg[1857]), .Z(n19794) );
  NANDN U20831 ( .A(n19771), .B(sreg[1856]), .Z(n19775) );
  NAND U20832 ( .A(n19773), .B(n19772), .Z(n19774) );
  NAND U20833 ( .A(n19775), .B(n19774), .Z(n19793) );
  XOR U20834 ( .A(n19794), .B(n19793), .Z(c[1857]) );
  NANDN U20835 ( .A(n19777), .B(n19776), .Z(n19781) );
  OR U20836 ( .A(n19779), .B(n19778), .Z(n19780) );
  AND U20837 ( .A(n19781), .B(n19780), .Z(n19799) );
  XOR U20838 ( .A(a[836]), .B(n2295), .Z(n19803) );
  AND U20839 ( .A(a[838]), .B(b[0]), .Z(n19783) );
  XNOR U20840 ( .A(n19783), .B(n2175), .Z(n19785) );
  NANDN U20841 ( .A(b[0]), .B(a[837]), .Z(n19784) );
  NAND U20842 ( .A(n19785), .B(n19784), .Z(n19808) );
  AND U20843 ( .A(a[834]), .B(b[3]), .Z(n19807) );
  XOR U20844 ( .A(n19808), .B(n19807), .Z(n19810) );
  XOR U20845 ( .A(n19809), .B(n19810), .Z(n19798) );
  NANDN U20846 ( .A(n19787), .B(n19786), .Z(n19791) );
  OR U20847 ( .A(n19789), .B(n19788), .Z(n19790) );
  AND U20848 ( .A(n19791), .B(n19790), .Z(n19797) );
  XOR U20849 ( .A(n19798), .B(n19797), .Z(n19800) );
  XOR U20850 ( .A(n19799), .B(n19800), .Z(n19813) );
  XNOR U20851 ( .A(n19813), .B(sreg[1858]), .Z(n19815) );
  NANDN U20852 ( .A(n19792), .B(sreg[1857]), .Z(n19796) );
  NAND U20853 ( .A(n19794), .B(n19793), .Z(n19795) );
  NAND U20854 ( .A(n19796), .B(n19795), .Z(n19814) );
  XOR U20855 ( .A(n19815), .B(n19814), .Z(c[1858]) );
  NANDN U20856 ( .A(n19798), .B(n19797), .Z(n19802) );
  OR U20857 ( .A(n19800), .B(n19799), .Z(n19801) );
  AND U20858 ( .A(n19802), .B(n19801), .Z(n19820) );
  XOR U20859 ( .A(a[837]), .B(n2295), .Z(n19824) );
  AND U20860 ( .A(a[835]), .B(b[3]), .Z(n19828) );
  AND U20861 ( .A(a[839]), .B(b[0]), .Z(n19804) );
  XNOR U20862 ( .A(n19804), .B(n2175), .Z(n19806) );
  NANDN U20863 ( .A(b[0]), .B(a[838]), .Z(n19805) );
  NAND U20864 ( .A(n19806), .B(n19805), .Z(n19829) );
  XOR U20865 ( .A(n19828), .B(n19829), .Z(n19831) );
  XOR U20866 ( .A(n19830), .B(n19831), .Z(n19819) );
  NANDN U20867 ( .A(n19808), .B(n19807), .Z(n19812) );
  OR U20868 ( .A(n19810), .B(n19809), .Z(n19811) );
  AND U20869 ( .A(n19812), .B(n19811), .Z(n19818) );
  XOR U20870 ( .A(n19819), .B(n19818), .Z(n19821) );
  XOR U20871 ( .A(n19820), .B(n19821), .Z(n19834) );
  XNOR U20872 ( .A(n19834), .B(sreg[1859]), .Z(n19836) );
  NANDN U20873 ( .A(n19813), .B(sreg[1858]), .Z(n19817) );
  NAND U20874 ( .A(n19815), .B(n19814), .Z(n19816) );
  NAND U20875 ( .A(n19817), .B(n19816), .Z(n19835) );
  XOR U20876 ( .A(n19836), .B(n19835), .Z(c[1859]) );
  NANDN U20877 ( .A(n19819), .B(n19818), .Z(n19823) );
  OR U20878 ( .A(n19821), .B(n19820), .Z(n19822) );
  AND U20879 ( .A(n19823), .B(n19822), .Z(n19841) );
  XOR U20880 ( .A(a[838]), .B(n2295), .Z(n19845) );
  AND U20881 ( .A(a[840]), .B(b[0]), .Z(n19825) );
  XNOR U20882 ( .A(n19825), .B(n2175), .Z(n19827) );
  NANDN U20883 ( .A(b[0]), .B(a[839]), .Z(n19826) );
  NAND U20884 ( .A(n19827), .B(n19826), .Z(n19850) );
  AND U20885 ( .A(a[836]), .B(b[3]), .Z(n19849) );
  XOR U20886 ( .A(n19850), .B(n19849), .Z(n19852) );
  XOR U20887 ( .A(n19851), .B(n19852), .Z(n19840) );
  NANDN U20888 ( .A(n19829), .B(n19828), .Z(n19833) );
  OR U20889 ( .A(n19831), .B(n19830), .Z(n19832) );
  AND U20890 ( .A(n19833), .B(n19832), .Z(n19839) );
  XOR U20891 ( .A(n19840), .B(n19839), .Z(n19842) );
  XOR U20892 ( .A(n19841), .B(n19842), .Z(n19855) );
  XNOR U20893 ( .A(n19855), .B(sreg[1860]), .Z(n19857) );
  NANDN U20894 ( .A(n19834), .B(sreg[1859]), .Z(n19838) );
  NAND U20895 ( .A(n19836), .B(n19835), .Z(n19837) );
  NAND U20896 ( .A(n19838), .B(n19837), .Z(n19856) );
  XOR U20897 ( .A(n19857), .B(n19856), .Z(c[1860]) );
  NANDN U20898 ( .A(n19840), .B(n19839), .Z(n19844) );
  OR U20899 ( .A(n19842), .B(n19841), .Z(n19843) );
  AND U20900 ( .A(n19844), .B(n19843), .Z(n19862) );
  XOR U20901 ( .A(a[839]), .B(n2296), .Z(n19866) );
  AND U20902 ( .A(a[841]), .B(b[0]), .Z(n19846) );
  XNOR U20903 ( .A(n19846), .B(n2175), .Z(n19848) );
  NANDN U20904 ( .A(b[0]), .B(a[840]), .Z(n19847) );
  NAND U20905 ( .A(n19848), .B(n19847), .Z(n19871) );
  AND U20906 ( .A(a[837]), .B(b[3]), .Z(n19870) );
  XOR U20907 ( .A(n19871), .B(n19870), .Z(n19873) );
  XOR U20908 ( .A(n19872), .B(n19873), .Z(n19861) );
  NANDN U20909 ( .A(n19850), .B(n19849), .Z(n19854) );
  OR U20910 ( .A(n19852), .B(n19851), .Z(n19853) );
  AND U20911 ( .A(n19854), .B(n19853), .Z(n19860) );
  XOR U20912 ( .A(n19861), .B(n19860), .Z(n19863) );
  XOR U20913 ( .A(n19862), .B(n19863), .Z(n19876) );
  XNOR U20914 ( .A(n19876), .B(sreg[1861]), .Z(n19878) );
  NANDN U20915 ( .A(n19855), .B(sreg[1860]), .Z(n19859) );
  NAND U20916 ( .A(n19857), .B(n19856), .Z(n19858) );
  NAND U20917 ( .A(n19859), .B(n19858), .Z(n19877) );
  XOR U20918 ( .A(n19878), .B(n19877), .Z(c[1861]) );
  NANDN U20919 ( .A(n19861), .B(n19860), .Z(n19865) );
  OR U20920 ( .A(n19863), .B(n19862), .Z(n19864) );
  AND U20921 ( .A(n19865), .B(n19864), .Z(n19883) );
  XOR U20922 ( .A(a[840]), .B(n2296), .Z(n19887) );
  AND U20923 ( .A(a[842]), .B(b[0]), .Z(n19867) );
  XNOR U20924 ( .A(n19867), .B(n2175), .Z(n19869) );
  NANDN U20925 ( .A(b[0]), .B(a[841]), .Z(n19868) );
  NAND U20926 ( .A(n19869), .B(n19868), .Z(n19892) );
  AND U20927 ( .A(a[838]), .B(b[3]), .Z(n19891) );
  XOR U20928 ( .A(n19892), .B(n19891), .Z(n19894) );
  XOR U20929 ( .A(n19893), .B(n19894), .Z(n19882) );
  NANDN U20930 ( .A(n19871), .B(n19870), .Z(n19875) );
  OR U20931 ( .A(n19873), .B(n19872), .Z(n19874) );
  AND U20932 ( .A(n19875), .B(n19874), .Z(n19881) );
  XOR U20933 ( .A(n19882), .B(n19881), .Z(n19884) );
  XOR U20934 ( .A(n19883), .B(n19884), .Z(n19897) );
  XNOR U20935 ( .A(n19897), .B(sreg[1862]), .Z(n19899) );
  NANDN U20936 ( .A(n19876), .B(sreg[1861]), .Z(n19880) );
  NAND U20937 ( .A(n19878), .B(n19877), .Z(n19879) );
  NAND U20938 ( .A(n19880), .B(n19879), .Z(n19898) );
  XOR U20939 ( .A(n19899), .B(n19898), .Z(c[1862]) );
  NANDN U20940 ( .A(n19882), .B(n19881), .Z(n19886) );
  OR U20941 ( .A(n19884), .B(n19883), .Z(n19885) );
  AND U20942 ( .A(n19886), .B(n19885), .Z(n19904) );
  XOR U20943 ( .A(a[841]), .B(n2296), .Z(n19908) );
  AND U20944 ( .A(a[843]), .B(b[0]), .Z(n19888) );
  XNOR U20945 ( .A(n19888), .B(n2175), .Z(n19890) );
  NANDN U20946 ( .A(b[0]), .B(a[842]), .Z(n19889) );
  NAND U20947 ( .A(n19890), .B(n19889), .Z(n19913) );
  AND U20948 ( .A(a[839]), .B(b[3]), .Z(n19912) );
  XOR U20949 ( .A(n19913), .B(n19912), .Z(n19915) );
  XOR U20950 ( .A(n19914), .B(n19915), .Z(n19903) );
  NANDN U20951 ( .A(n19892), .B(n19891), .Z(n19896) );
  OR U20952 ( .A(n19894), .B(n19893), .Z(n19895) );
  AND U20953 ( .A(n19896), .B(n19895), .Z(n19902) );
  XOR U20954 ( .A(n19903), .B(n19902), .Z(n19905) );
  XOR U20955 ( .A(n19904), .B(n19905), .Z(n19918) );
  XNOR U20956 ( .A(n19918), .B(sreg[1863]), .Z(n19920) );
  NANDN U20957 ( .A(n19897), .B(sreg[1862]), .Z(n19901) );
  NAND U20958 ( .A(n19899), .B(n19898), .Z(n19900) );
  NAND U20959 ( .A(n19901), .B(n19900), .Z(n19919) );
  XOR U20960 ( .A(n19920), .B(n19919), .Z(c[1863]) );
  NANDN U20961 ( .A(n19903), .B(n19902), .Z(n19907) );
  OR U20962 ( .A(n19905), .B(n19904), .Z(n19906) );
  AND U20963 ( .A(n19907), .B(n19906), .Z(n19925) );
  XOR U20964 ( .A(a[842]), .B(n2296), .Z(n19929) );
  AND U20965 ( .A(a[844]), .B(b[0]), .Z(n19909) );
  XNOR U20966 ( .A(n19909), .B(n2175), .Z(n19911) );
  NANDN U20967 ( .A(b[0]), .B(a[843]), .Z(n19910) );
  NAND U20968 ( .A(n19911), .B(n19910), .Z(n19934) );
  AND U20969 ( .A(a[840]), .B(b[3]), .Z(n19933) );
  XOR U20970 ( .A(n19934), .B(n19933), .Z(n19936) );
  XOR U20971 ( .A(n19935), .B(n19936), .Z(n19924) );
  NANDN U20972 ( .A(n19913), .B(n19912), .Z(n19917) );
  OR U20973 ( .A(n19915), .B(n19914), .Z(n19916) );
  AND U20974 ( .A(n19917), .B(n19916), .Z(n19923) );
  XOR U20975 ( .A(n19924), .B(n19923), .Z(n19926) );
  XOR U20976 ( .A(n19925), .B(n19926), .Z(n19939) );
  XNOR U20977 ( .A(n19939), .B(sreg[1864]), .Z(n19941) );
  NANDN U20978 ( .A(n19918), .B(sreg[1863]), .Z(n19922) );
  NAND U20979 ( .A(n19920), .B(n19919), .Z(n19921) );
  NAND U20980 ( .A(n19922), .B(n19921), .Z(n19940) );
  XOR U20981 ( .A(n19941), .B(n19940), .Z(c[1864]) );
  NANDN U20982 ( .A(n19924), .B(n19923), .Z(n19928) );
  OR U20983 ( .A(n19926), .B(n19925), .Z(n19927) );
  AND U20984 ( .A(n19928), .B(n19927), .Z(n19946) );
  XOR U20985 ( .A(a[843]), .B(n2296), .Z(n19950) );
  AND U20986 ( .A(a[841]), .B(b[3]), .Z(n19954) );
  AND U20987 ( .A(a[845]), .B(b[0]), .Z(n19930) );
  XNOR U20988 ( .A(n19930), .B(n2175), .Z(n19932) );
  NANDN U20989 ( .A(b[0]), .B(a[844]), .Z(n19931) );
  NAND U20990 ( .A(n19932), .B(n19931), .Z(n19955) );
  XOR U20991 ( .A(n19954), .B(n19955), .Z(n19957) );
  XOR U20992 ( .A(n19956), .B(n19957), .Z(n19945) );
  NANDN U20993 ( .A(n19934), .B(n19933), .Z(n19938) );
  OR U20994 ( .A(n19936), .B(n19935), .Z(n19937) );
  AND U20995 ( .A(n19938), .B(n19937), .Z(n19944) );
  XOR U20996 ( .A(n19945), .B(n19944), .Z(n19947) );
  XOR U20997 ( .A(n19946), .B(n19947), .Z(n19960) );
  XNOR U20998 ( .A(n19960), .B(sreg[1865]), .Z(n19962) );
  NANDN U20999 ( .A(n19939), .B(sreg[1864]), .Z(n19943) );
  NAND U21000 ( .A(n19941), .B(n19940), .Z(n19942) );
  NAND U21001 ( .A(n19943), .B(n19942), .Z(n19961) );
  XOR U21002 ( .A(n19962), .B(n19961), .Z(c[1865]) );
  NANDN U21003 ( .A(n19945), .B(n19944), .Z(n19949) );
  OR U21004 ( .A(n19947), .B(n19946), .Z(n19948) );
  AND U21005 ( .A(n19949), .B(n19948), .Z(n19967) );
  XOR U21006 ( .A(a[844]), .B(n2296), .Z(n19971) );
  AND U21007 ( .A(a[846]), .B(b[0]), .Z(n19951) );
  XNOR U21008 ( .A(n19951), .B(n2175), .Z(n19953) );
  NANDN U21009 ( .A(b[0]), .B(a[845]), .Z(n19952) );
  NAND U21010 ( .A(n19953), .B(n19952), .Z(n19976) );
  AND U21011 ( .A(a[842]), .B(b[3]), .Z(n19975) );
  XOR U21012 ( .A(n19976), .B(n19975), .Z(n19978) );
  XOR U21013 ( .A(n19977), .B(n19978), .Z(n19966) );
  NANDN U21014 ( .A(n19955), .B(n19954), .Z(n19959) );
  OR U21015 ( .A(n19957), .B(n19956), .Z(n19958) );
  AND U21016 ( .A(n19959), .B(n19958), .Z(n19965) );
  XOR U21017 ( .A(n19966), .B(n19965), .Z(n19968) );
  XOR U21018 ( .A(n19967), .B(n19968), .Z(n19981) );
  XNOR U21019 ( .A(n19981), .B(sreg[1866]), .Z(n19983) );
  NANDN U21020 ( .A(n19960), .B(sreg[1865]), .Z(n19964) );
  NAND U21021 ( .A(n19962), .B(n19961), .Z(n19963) );
  NAND U21022 ( .A(n19964), .B(n19963), .Z(n19982) );
  XOR U21023 ( .A(n19983), .B(n19982), .Z(c[1866]) );
  NANDN U21024 ( .A(n19966), .B(n19965), .Z(n19970) );
  OR U21025 ( .A(n19968), .B(n19967), .Z(n19969) );
  AND U21026 ( .A(n19970), .B(n19969), .Z(n19988) );
  XOR U21027 ( .A(a[845]), .B(n2296), .Z(n19992) );
  AND U21028 ( .A(a[847]), .B(b[0]), .Z(n19972) );
  XNOR U21029 ( .A(n19972), .B(n2175), .Z(n19974) );
  NANDN U21030 ( .A(b[0]), .B(a[846]), .Z(n19973) );
  NAND U21031 ( .A(n19974), .B(n19973), .Z(n19997) );
  AND U21032 ( .A(a[843]), .B(b[3]), .Z(n19996) );
  XOR U21033 ( .A(n19997), .B(n19996), .Z(n19999) );
  XOR U21034 ( .A(n19998), .B(n19999), .Z(n19987) );
  NANDN U21035 ( .A(n19976), .B(n19975), .Z(n19980) );
  OR U21036 ( .A(n19978), .B(n19977), .Z(n19979) );
  AND U21037 ( .A(n19980), .B(n19979), .Z(n19986) );
  XOR U21038 ( .A(n19987), .B(n19986), .Z(n19989) );
  XOR U21039 ( .A(n19988), .B(n19989), .Z(n20002) );
  XNOR U21040 ( .A(n20002), .B(sreg[1867]), .Z(n20004) );
  NANDN U21041 ( .A(n19981), .B(sreg[1866]), .Z(n19985) );
  NAND U21042 ( .A(n19983), .B(n19982), .Z(n19984) );
  NAND U21043 ( .A(n19985), .B(n19984), .Z(n20003) );
  XOR U21044 ( .A(n20004), .B(n20003), .Z(c[1867]) );
  NANDN U21045 ( .A(n19987), .B(n19986), .Z(n19991) );
  OR U21046 ( .A(n19989), .B(n19988), .Z(n19990) );
  AND U21047 ( .A(n19991), .B(n19990), .Z(n20009) );
  XOR U21048 ( .A(a[846]), .B(n2297), .Z(n20013) );
  AND U21049 ( .A(a[848]), .B(b[0]), .Z(n19993) );
  XNOR U21050 ( .A(n19993), .B(n2175), .Z(n19995) );
  NANDN U21051 ( .A(b[0]), .B(a[847]), .Z(n19994) );
  NAND U21052 ( .A(n19995), .B(n19994), .Z(n20018) );
  AND U21053 ( .A(a[844]), .B(b[3]), .Z(n20017) );
  XOR U21054 ( .A(n20018), .B(n20017), .Z(n20020) );
  XOR U21055 ( .A(n20019), .B(n20020), .Z(n20008) );
  NANDN U21056 ( .A(n19997), .B(n19996), .Z(n20001) );
  OR U21057 ( .A(n19999), .B(n19998), .Z(n20000) );
  AND U21058 ( .A(n20001), .B(n20000), .Z(n20007) );
  XOR U21059 ( .A(n20008), .B(n20007), .Z(n20010) );
  XOR U21060 ( .A(n20009), .B(n20010), .Z(n20023) );
  XNOR U21061 ( .A(n20023), .B(sreg[1868]), .Z(n20025) );
  NANDN U21062 ( .A(n20002), .B(sreg[1867]), .Z(n20006) );
  NAND U21063 ( .A(n20004), .B(n20003), .Z(n20005) );
  NAND U21064 ( .A(n20006), .B(n20005), .Z(n20024) );
  XOR U21065 ( .A(n20025), .B(n20024), .Z(c[1868]) );
  NANDN U21066 ( .A(n20008), .B(n20007), .Z(n20012) );
  OR U21067 ( .A(n20010), .B(n20009), .Z(n20011) );
  AND U21068 ( .A(n20012), .B(n20011), .Z(n20030) );
  XOR U21069 ( .A(a[847]), .B(n2297), .Z(n20034) );
  AND U21070 ( .A(a[845]), .B(b[3]), .Z(n20038) );
  AND U21071 ( .A(a[849]), .B(b[0]), .Z(n20014) );
  XNOR U21072 ( .A(n20014), .B(n2175), .Z(n20016) );
  NANDN U21073 ( .A(b[0]), .B(a[848]), .Z(n20015) );
  NAND U21074 ( .A(n20016), .B(n20015), .Z(n20039) );
  XOR U21075 ( .A(n20038), .B(n20039), .Z(n20041) );
  XOR U21076 ( .A(n20040), .B(n20041), .Z(n20029) );
  NANDN U21077 ( .A(n20018), .B(n20017), .Z(n20022) );
  OR U21078 ( .A(n20020), .B(n20019), .Z(n20021) );
  AND U21079 ( .A(n20022), .B(n20021), .Z(n20028) );
  XOR U21080 ( .A(n20029), .B(n20028), .Z(n20031) );
  XOR U21081 ( .A(n20030), .B(n20031), .Z(n20044) );
  XNOR U21082 ( .A(n20044), .B(sreg[1869]), .Z(n20046) );
  NANDN U21083 ( .A(n20023), .B(sreg[1868]), .Z(n20027) );
  NAND U21084 ( .A(n20025), .B(n20024), .Z(n20026) );
  NAND U21085 ( .A(n20027), .B(n20026), .Z(n20045) );
  XOR U21086 ( .A(n20046), .B(n20045), .Z(c[1869]) );
  NANDN U21087 ( .A(n20029), .B(n20028), .Z(n20033) );
  OR U21088 ( .A(n20031), .B(n20030), .Z(n20032) );
  AND U21089 ( .A(n20033), .B(n20032), .Z(n20051) );
  XOR U21090 ( .A(a[848]), .B(n2297), .Z(n20055) );
  AND U21091 ( .A(a[850]), .B(b[0]), .Z(n20035) );
  XNOR U21092 ( .A(n20035), .B(n2175), .Z(n20037) );
  NANDN U21093 ( .A(b[0]), .B(a[849]), .Z(n20036) );
  NAND U21094 ( .A(n20037), .B(n20036), .Z(n20060) );
  AND U21095 ( .A(a[846]), .B(b[3]), .Z(n20059) );
  XOR U21096 ( .A(n20060), .B(n20059), .Z(n20062) );
  XOR U21097 ( .A(n20061), .B(n20062), .Z(n20050) );
  NANDN U21098 ( .A(n20039), .B(n20038), .Z(n20043) );
  OR U21099 ( .A(n20041), .B(n20040), .Z(n20042) );
  AND U21100 ( .A(n20043), .B(n20042), .Z(n20049) );
  XOR U21101 ( .A(n20050), .B(n20049), .Z(n20052) );
  XOR U21102 ( .A(n20051), .B(n20052), .Z(n20065) );
  XNOR U21103 ( .A(n20065), .B(sreg[1870]), .Z(n20067) );
  NANDN U21104 ( .A(n20044), .B(sreg[1869]), .Z(n20048) );
  NAND U21105 ( .A(n20046), .B(n20045), .Z(n20047) );
  NAND U21106 ( .A(n20048), .B(n20047), .Z(n20066) );
  XOR U21107 ( .A(n20067), .B(n20066), .Z(c[1870]) );
  NANDN U21108 ( .A(n20050), .B(n20049), .Z(n20054) );
  OR U21109 ( .A(n20052), .B(n20051), .Z(n20053) );
  AND U21110 ( .A(n20054), .B(n20053), .Z(n20072) );
  XOR U21111 ( .A(a[849]), .B(n2297), .Z(n20076) );
  AND U21112 ( .A(a[851]), .B(b[0]), .Z(n20056) );
  XNOR U21113 ( .A(n20056), .B(n2175), .Z(n20058) );
  NANDN U21114 ( .A(b[0]), .B(a[850]), .Z(n20057) );
  NAND U21115 ( .A(n20058), .B(n20057), .Z(n20081) );
  AND U21116 ( .A(a[847]), .B(b[3]), .Z(n20080) );
  XOR U21117 ( .A(n20081), .B(n20080), .Z(n20083) );
  XOR U21118 ( .A(n20082), .B(n20083), .Z(n20071) );
  NANDN U21119 ( .A(n20060), .B(n20059), .Z(n20064) );
  OR U21120 ( .A(n20062), .B(n20061), .Z(n20063) );
  AND U21121 ( .A(n20064), .B(n20063), .Z(n20070) );
  XOR U21122 ( .A(n20071), .B(n20070), .Z(n20073) );
  XOR U21123 ( .A(n20072), .B(n20073), .Z(n20086) );
  XNOR U21124 ( .A(n20086), .B(sreg[1871]), .Z(n20088) );
  NANDN U21125 ( .A(n20065), .B(sreg[1870]), .Z(n20069) );
  NAND U21126 ( .A(n20067), .B(n20066), .Z(n20068) );
  NAND U21127 ( .A(n20069), .B(n20068), .Z(n20087) );
  XOR U21128 ( .A(n20088), .B(n20087), .Z(c[1871]) );
  NANDN U21129 ( .A(n20071), .B(n20070), .Z(n20075) );
  OR U21130 ( .A(n20073), .B(n20072), .Z(n20074) );
  AND U21131 ( .A(n20075), .B(n20074), .Z(n20093) );
  XOR U21132 ( .A(a[850]), .B(n2297), .Z(n20097) );
  AND U21133 ( .A(a[848]), .B(b[3]), .Z(n20101) );
  AND U21134 ( .A(a[852]), .B(b[0]), .Z(n20077) );
  XNOR U21135 ( .A(n20077), .B(n2175), .Z(n20079) );
  NANDN U21136 ( .A(b[0]), .B(a[851]), .Z(n20078) );
  NAND U21137 ( .A(n20079), .B(n20078), .Z(n20102) );
  XOR U21138 ( .A(n20101), .B(n20102), .Z(n20104) );
  XOR U21139 ( .A(n20103), .B(n20104), .Z(n20092) );
  NANDN U21140 ( .A(n20081), .B(n20080), .Z(n20085) );
  OR U21141 ( .A(n20083), .B(n20082), .Z(n20084) );
  AND U21142 ( .A(n20085), .B(n20084), .Z(n20091) );
  XOR U21143 ( .A(n20092), .B(n20091), .Z(n20094) );
  XOR U21144 ( .A(n20093), .B(n20094), .Z(n20107) );
  XNOR U21145 ( .A(n20107), .B(sreg[1872]), .Z(n20109) );
  NANDN U21146 ( .A(n20086), .B(sreg[1871]), .Z(n20090) );
  NAND U21147 ( .A(n20088), .B(n20087), .Z(n20089) );
  NAND U21148 ( .A(n20090), .B(n20089), .Z(n20108) );
  XOR U21149 ( .A(n20109), .B(n20108), .Z(c[1872]) );
  NANDN U21150 ( .A(n20092), .B(n20091), .Z(n20096) );
  OR U21151 ( .A(n20094), .B(n20093), .Z(n20095) );
  AND U21152 ( .A(n20096), .B(n20095), .Z(n20114) );
  XOR U21153 ( .A(a[851]), .B(n2297), .Z(n20118) );
  AND U21154 ( .A(a[853]), .B(b[0]), .Z(n20098) );
  XNOR U21155 ( .A(n20098), .B(n2175), .Z(n20100) );
  NANDN U21156 ( .A(b[0]), .B(a[852]), .Z(n20099) );
  NAND U21157 ( .A(n20100), .B(n20099), .Z(n20123) );
  AND U21158 ( .A(a[849]), .B(b[3]), .Z(n20122) );
  XOR U21159 ( .A(n20123), .B(n20122), .Z(n20125) );
  XOR U21160 ( .A(n20124), .B(n20125), .Z(n20113) );
  NANDN U21161 ( .A(n20102), .B(n20101), .Z(n20106) );
  OR U21162 ( .A(n20104), .B(n20103), .Z(n20105) );
  AND U21163 ( .A(n20106), .B(n20105), .Z(n20112) );
  XOR U21164 ( .A(n20113), .B(n20112), .Z(n20115) );
  XOR U21165 ( .A(n20114), .B(n20115), .Z(n20128) );
  XNOR U21166 ( .A(n20128), .B(sreg[1873]), .Z(n20130) );
  NANDN U21167 ( .A(n20107), .B(sreg[1872]), .Z(n20111) );
  NAND U21168 ( .A(n20109), .B(n20108), .Z(n20110) );
  NAND U21169 ( .A(n20111), .B(n20110), .Z(n20129) );
  XOR U21170 ( .A(n20130), .B(n20129), .Z(c[1873]) );
  NANDN U21171 ( .A(n20113), .B(n20112), .Z(n20117) );
  OR U21172 ( .A(n20115), .B(n20114), .Z(n20116) );
  AND U21173 ( .A(n20117), .B(n20116), .Z(n20136) );
  XOR U21174 ( .A(a[852]), .B(n2297), .Z(n20137) );
  AND U21175 ( .A(b[0]), .B(a[854]), .Z(n20119) );
  XOR U21176 ( .A(b[1]), .B(n20119), .Z(n20121) );
  NANDN U21177 ( .A(b[0]), .B(a[853]), .Z(n20120) );
  AND U21178 ( .A(n20121), .B(n20120), .Z(n20141) );
  AND U21179 ( .A(a[850]), .B(b[3]), .Z(n20142) );
  XOR U21180 ( .A(n20141), .B(n20142), .Z(n20143) );
  XNOR U21181 ( .A(n20144), .B(n20143), .Z(n20133) );
  NANDN U21182 ( .A(n20123), .B(n20122), .Z(n20127) );
  OR U21183 ( .A(n20125), .B(n20124), .Z(n20126) );
  AND U21184 ( .A(n20127), .B(n20126), .Z(n20134) );
  XNOR U21185 ( .A(n20133), .B(n20134), .Z(n20135) );
  XNOR U21186 ( .A(n20136), .B(n20135), .Z(n20147) );
  XNOR U21187 ( .A(n20147), .B(sreg[1874]), .Z(n20149) );
  NANDN U21188 ( .A(n20128), .B(sreg[1873]), .Z(n20132) );
  NAND U21189 ( .A(n20130), .B(n20129), .Z(n20131) );
  NAND U21190 ( .A(n20132), .B(n20131), .Z(n20148) );
  XOR U21191 ( .A(n20149), .B(n20148), .Z(c[1874]) );
  XOR U21192 ( .A(a[853]), .B(n2298), .Z(n20156) );
  AND U21193 ( .A(a[855]), .B(b[0]), .Z(n20138) );
  XNOR U21194 ( .A(n20138), .B(n2175), .Z(n20140) );
  NANDN U21195 ( .A(b[0]), .B(a[854]), .Z(n20139) );
  NAND U21196 ( .A(n20140), .B(n20139), .Z(n20161) );
  AND U21197 ( .A(a[851]), .B(b[3]), .Z(n20160) );
  XOR U21198 ( .A(n20161), .B(n20160), .Z(n20163) );
  XOR U21199 ( .A(n20162), .B(n20163), .Z(n20151) );
  NAND U21200 ( .A(n20142), .B(n20141), .Z(n20146) );
  NANDN U21201 ( .A(n20144), .B(n20143), .Z(n20145) );
  AND U21202 ( .A(n20146), .B(n20145), .Z(n20150) );
  XOR U21203 ( .A(n20151), .B(n20150), .Z(n20153) );
  XOR U21204 ( .A(n20152), .B(n20153), .Z(n20166) );
  XNOR U21205 ( .A(n20166), .B(sreg[1875]), .Z(n20168) );
  XOR U21206 ( .A(n20168), .B(n20167), .Z(c[1875]) );
  NANDN U21207 ( .A(n20151), .B(n20150), .Z(n20155) );
  OR U21208 ( .A(n20153), .B(n20152), .Z(n20154) );
  AND U21209 ( .A(n20155), .B(n20154), .Z(n20173) );
  XOR U21210 ( .A(a[854]), .B(n2298), .Z(n20177) );
  AND U21211 ( .A(a[856]), .B(b[0]), .Z(n20157) );
  XNOR U21212 ( .A(n20157), .B(n2175), .Z(n20159) );
  NANDN U21213 ( .A(b[0]), .B(a[855]), .Z(n20158) );
  NAND U21214 ( .A(n20159), .B(n20158), .Z(n20182) );
  AND U21215 ( .A(a[852]), .B(b[3]), .Z(n20181) );
  XOR U21216 ( .A(n20182), .B(n20181), .Z(n20184) );
  XOR U21217 ( .A(n20183), .B(n20184), .Z(n20172) );
  NANDN U21218 ( .A(n20161), .B(n20160), .Z(n20165) );
  OR U21219 ( .A(n20163), .B(n20162), .Z(n20164) );
  AND U21220 ( .A(n20165), .B(n20164), .Z(n20171) );
  XOR U21221 ( .A(n20172), .B(n20171), .Z(n20174) );
  XOR U21222 ( .A(n20173), .B(n20174), .Z(n20187) );
  XNOR U21223 ( .A(n20187), .B(sreg[1876]), .Z(n20189) );
  NANDN U21224 ( .A(n20166), .B(sreg[1875]), .Z(n20170) );
  NAND U21225 ( .A(n20168), .B(n20167), .Z(n20169) );
  NAND U21226 ( .A(n20170), .B(n20169), .Z(n20188) );
  XOR U21227 ( .A(n20189), .B(n20188), .Z(c[1876]) );
  NANDN U21228 ( .A(n20172), .B(n20171), .Z(n20176) );
  OR U21229 ( .A(n20174), .B(n20173), .Z(n20175) );
  AND U21230 ( .A(n20176), .B(n20175), .Z(n20194) );
  XOR U21231 ( .A(a[855]), .B(n2298), .Z(n20198) );
  AND U21232 ( .A(a[853]), .B(b[3]), .Z(n20202) );
  AND U21233 ( .A(a[857]), .B(b[0]), .Z(n20178) );
  XNOR U21234 ( .A(n20178), .B(n2175), .Z(n20180) );
  NANDN U21235 ( .A(b[0]), .B(a[856]), .Z(n20179) );
  NAND U21236 ( .A(n20180), .B(n20179), .Z(n20203) );
  XOR U21237 ( .A(n20202), .B(n20203), .Z(n20205) );
  XOR U21238 ( .A(n20204), .B(n20205), .Z(n20193) );
  NANDN U21239 ( .A(n20182), .B(n20181), .Z(n20186) );
  OR U21240 ( .A(n20184), .B(n20183), .Z(n20185) );
  AND U21241 ( .A(n20186), .B(n20185), .Z(n20192) );
  XOR U21242 ( .A(n20193), .B(n20192), .Z(n20195) );
  XOR U21243 ( .A(n20194), .B(n20195), .Z(n20208) );
  XNOR U21244 ( .A(n20208), .B(sreg[1877]), .Z(n20210) );
  NANDN U21245 ( .A(n20187), .B(sreg[1876]), .Z(n20191) );
  NAND U21246 ( .A(n20189), .B(n20188), .Z(n20190) );
  NAND U21247 ( .A(n20191), .B(n20190), .Z(n20209) );
  XOR U21248 ( .A(n20210), .B(n20209), .Z(c[1877]) );
  NANDN U21249 ( .A(n20193), .B(n20192), .Z(n20197) );
  OR U21250 ( .A(n20195), .B(n20194), .Z(n20196) );
  AND U21251 ( .A(n20197), .B(n20196), .Z(n20215) );
  XOR U21252 ( .A(a[856]), .B(n2298), .Z(n20219) );
  AND U21253 ( .A(a[858]), .B(b[0]), .Z(n20199) );
  XNOR U21254 ( .A(n20199), .B(n2175), .Z(n20201) );
  NANDN U21255 ( .A(b[0]), .B(a[857]), .Z(n20200) );
  NAND U21256 ( .A(n20201), .B(n20200), .Z(n20224) );
  AND U21257 ( .A(a[854]), .B(b[3]), .Z(n20223) );
  XOR U21258 ( .A(n20224), .B(n20223), .Z(n20226) );
  XOR U21259 ( .A(n20225), .B(n20226), .Z(n20214) );
  NANDN U21260 ( .A(n20203), .B(n20202), .Z(n20207) );
  OR U21261 ( .A(n20205), .B(n20204), .Z(n20206) );
  AND U21262 ( .A(n20207), .B(n20206), .Z(n20213) );
  XOR U21263 ( .A(n20214), .B(n20213), .Z(n20216) );
  XOR U21264 ( .A(n20215), .B(n20216), .Z(n20229) );
  XNOR U21265 ( .A(n20229), .B(sreg[1878]), .Z(n20231) );
  NANDN U21266 ( .A(n20208), .B(sreg[1877]), .Z(n20212) );
  NAND U21267 ( .A(n20210), .B(n20209), .Z(n20211) );
  NAND U21268 ( .A(n20212), .B(n20211), .Z(n20230) );
  XOR U21269 ( .A(n20231), .B(n20230), .Z(c[1878]) );
  NANDN U21270 ( .A(n20214), .B(n20213), .Z(n20218) );
  OR U21271 ( .A(n20216), .B(n20215), .Z(n20217) );
  AND U21272 ( .A(n20218), .B(n20217), .Z(n20236) );
  XOR U21273 ( .A(a[857]), .B(n2298), .Z(n20240) );
  AND U21274 ( .A(a[859]), .B(b[0]), .Z(n20220) );
  XNOR U21275 ( .A(n20220), .B(n2175), .Z(n20222) );
  NANDN U21276 ( .A(b[0]), .B(a[858]), .Z(n20221) );
  NAND U21277 ( .A(n20222), .B(n20221), .Z(n20245) );
  AND U21278 ( .A(a[855]), .B(b[3]), .Z(n20244) );
  XOR U21279 ( .A(n20245), .B(n20244), .Z(n20247) );
  XOR U21280 ( .A(n20246), .B(n20247), .Z(n20235) );
  NANDN U21281 ( .A(n20224), .B(n20223), .Z(n20228) );
  OR U21282 ( .A(n20226), .B(n20225), .Z(n20227) );
  AND U21283 ( .A(n20228), .B(n20227), .Z(n20234) );
  XOR U21284 ( .A(n20235), .B(n20234), .Z(n20237) );
  XOR U21285 ( .A(n20236), .B(n20237), .Z(n20250) );
  XNOR U21286 ( .A(n20250), .B(sreg[1879]), .Z(n20252) );
  NANDN U21287 ( .A(n20229), .B(sreg[1878]), .Z(n20233) );
  NAND U21288 ( .A(n20231), .B(n20230), .Z(n20232) );
  NAND U21289 ( .A(n20233), .B(n20232), .Z(n20251) );
  XOR U21290 ( .A(n20252), .B(n20251), .Z(c[1879]) );
  NANDN U21291 ( .A(n20235), .B(n20234), .Z(n20239) );
  OR U21292 ( .A(n20237), .B(n20236), .Z(n20238) );
  AND U21293 ( .A(n20239), .B(n20238), .Z(n20257) );
  XOR U21294 ( .A(a[858]), .B(n2298), .Z(n20261) );
  AND U21295 ( .A(a[856]), .B(b[3]), .Z(n20265) );
  AND U21296 ( .A(a[860]), .B(b[0]), .Z(n20241) );
  XNOR U21297 ( .A(n20241), .B(n2175), .Z(n20243) );
  NANDN U21298 ( .A(b[0]), .B(a[859]), .Z(n20242) );
  NAND U21299 ( .A(n20243), .B(n20242), .Z(n20266) );
  XOR U21300 ( .A(n20265), .B(n20266), .Z(n20268) );
  XOR U21301 ( .A(n20267), .B(n20268), .Z(n20256) );
  NANDN U21302 ( .A(n20245), .B(n20244), .Z(n20249) );
  OR U21303 ( .A(n20247), .B(n20246), .Z(n20248) );
  AND U21304 ( .A(n20249), .B(n20248), .Z(n20255) );
  XOR U21305 ( .A(n20256), .B(n20255), .Z(n20258) );
  XOR U21306 ( .A(n20257), .B(n20258), .Z(n20271) );
  XNOR U21307 ( .A(n20271), .B(sreg[1880]), .Z(n20273) );
  NANDN U21308 ( .A(n20250), .B(sreg[1879]), .Z(n20254) );
  NAND U21309 ( .A(n20252), .B(n20251), .Z(n20253) );
  NAND U21310 ( .A(n20254), .B(n20253), .Z(n20272) );
  XOR U21311 ( .A(n20273), .B(n20272), .Z(c[1880]) );
  NANDN U21312 ( .A(n20256), .B(n20255), .Z(n20260) );
  OR U21313 ( .A(n20258), .B(n20257), .Z(n20259) );
  AND U21314 ( .A(n20260), .B(n20259), .Z(n20278) );
  XOR U21315 ( .A(a[859]), .B(n2298), .Z(n20282) );
  AND U21316 ( .A(a[861]), .B(b[0]), .Z(n20262) );
  XNOR U21317 ( .A(n20262), .B(n2175), .Z(n20264) );
  NANDN U21318 ( .A(b[0]), .B(a[860]), .Z(n20263) );
  NAND U21319 ( .A(n20264), .B(n20263), .Z(n20287) );
  AND U21320 ( .A(a[857]), .B(b[3]), .Z(n20286) );
  XOR U21321 ( .A(n20287), .B(n20286), .Z(n20289) );
  XOR U21322 ( .A(n20288), .B(n20289), .Z(n20277) );
  NANDN U21323 ( .A(n20266), .B(n20265), .Z(n20270) );
  OR U21324 ( .A(n20268), .B(n20267), .Z(n20269) );
  AND U21325 ( .A(n20270), .B(n20269), .Z(n20276) );
  XOR U21326 ( .A(n20277), .B(n20276), .Z(n20279) );
  XOR U21327 ( .A(n20278), .B(n20279), .Z(n20292) );
  XNOR U21328 ( .A(n20292), .B(sreg[1881]), .Z(n20294) );
  NANDN U21329 ( .A(n20271), .B(sreg[1880]), .Z(n20275) );
  NAND U21330 ( .A(n20273), .B(n20272), .Z(n20274) );
  NAND U21331 ( .A(n20275), .B(n20274), .Z(n20293) );
  XOR U21332 ( .A(n20294), .B(n20293), .Z(c[1881]) );
  NANDN U21333 ( .A(n20277), .B(n20276), .Z(n20281) );
  OR U21334 ( .A(n20279), .B(n20278), .Z(n20280) );
  AND U21335 ( .A(n20281), .B(n20280), .Z(n20299) );
  XOR U21336 ( .A(a[860]), .B(n2299), .Z(n20303) );
  AND U21337 ( .A(a[858]), .B(b[3]), .Z(n20307) );
  AND U21338 ( .A(a[862]), .B(b[0]), .Z(n20283) );
  XNOR U21339 ( .A(n20283), .B(n2175), .Z(n20285) );
  NANDN U21340 ( .A(b[0]), .B(a[861]), .Z(n20284) );
  NAND U21341 ( .A(n20285), .B(n20284), .Z(n20308) );
  XOR U21342 ( .A(n20307), .B(n20308), .Z(n20310) );
  XOR U21343 ( .A(n20309), .B(n20310), .Z(n20298) );
  NANDN U21344 ( .A(n20287), .B(n20286), .Z(n20291) );
  OR U21345 ( .A(n20289), .B(n20288), .Z(n20290) );
  AND U21346 ( .A(n20291), .B(n20290), .Z(n20297) );
  XOR U21347 ( .A(n20298), .B(n20297), .Z(n20300) );
  XOR U21348 ( .A(n20299), .B(n20300), .Z(n20313) );
  XNOR U21349 ( .A(n20313), .B(sreg[1882]), .Z(n20315) );
  NANDN U21350 ( .A(n20292), .B(sreg[1881]), .Z(n20296) );
  NAND U21351 ( .A(n20294), .B(n20293), .Z(n20295) );
  NAND U21352 ( .A(n20296), .B(n20295), .Z(n20314) );
  XOR U21353 ( .A(n20315), .B(n20314), .Z(c[1882]) );
  NANDN U21354 ( .A(n20298), .B(n20297), .Z(n20302) );
  OR U21355 ( .A(n20300), .B(n20299), .Z(n20301) );
  AND U21356 ( .A(n20302), .B(n20301), .Z(n20320) );
  XOR U21357 ( .A(a[861]), .B(n2299), .Z(n20324) );
  AND U21358 ( .A(a[863]), .B(b[0]), .Z(n20304) );
  XNOR U21359 ( .A(n20304), .B(n2175), .Z(n20306) );
  NANDN U21360 ( .A(b[0]), .B(a[862]), .Z(n20305) );
  NAND U21361 ( .A(n20306), .B(n20305), .Z(n20329) );
  AND U21362 ( .A(a[859]), .B(b[3]), .Z(n20328) );
  XOR U21363 ( .A(n20329), .B(n20328), .Z(n20331) );
  XOR U21364 ( .A(n20330), .B(n20331), .Z(n20319) );
  NANDN U21365 ( .A(n20308), .B(n20307), .Z(n20312) );
  OR U21366 ( .A(n20310), .B(n20309), .Z(n20311) );
  AND U21367 ( .A(n20312), .B(n20311), .Z(n20318) );
  XOR U21368 ( .A(n20319), .B(n20318), .Z(n20321) );
  XOR U21369 ( .A(n20320), .B(n20321), .Z(n20334) );
  XNOR U21370 ( .A(n20334), .B(sreg[1883]), .Z(n20336) );
  NANDN U21371 ( .A(n20313), .B(sreg[1882]), .Z(n20317) );
  NAND U21372 ( .A(n20315), .B(n20314), .Z(n20316) );
  NAND U21373 ( .A(n20317), .B(n20316), .Z(n20335) );
  XOR U21374 ( .A(n20336), .B(n20335), .Z(c[1883]) );
  NANDN U21375 ( .A(n20319), .B(n20318), .Z(n20323) );
  OR U21376 ( .A(n20321), .B(n20320), .Z(n20322) );
  AND U21377 ( .A(n20323), .B(n20322), .Z(n20341) );
  XOR U21378 ( .A(a[862]), .B(n2299), .Z(n20345) );
  AND U21379 ( .A(a[860]), .B(b[3]), .Z(n20349) );
  AND U21380 ( .A(a[864]), .B(b[0]), .Z(n20325) );
  XNOR U21381 ( .A(n20325), .B(n2175), .Z(n20327) );
  NANDN U21382 ( .A(b[0]), .B(a[863]), .Z(n20326) );
  NAND U21383 ( .A(n20327), .B(n20326), .Z(n20350) );
  XOR U21384 ( .A(n20349), .B(n20350), .Z(n20352) );
  XOR U21385 ( .A(n20351), .B(n20352), .Z(n20340) );
  NANDN U21386 ( .A(n20329), .B(n20328), .Z(n20333) );
  OR U21387 ( .A(n20331), .B(n20330), .Z(n20332) );
  AND U21388 ( .A(n20333), .B(n20332), .Z(n20339) );
  XOR U21389 ( .A(n20340), .B(n20339), .Z(n20342) );
  XOR U21390 ( .A(n20341), .B(n20342), .Z(n20355) );
  XNOR U21391 ( .A(n20355), .B(sreg[1884]), .Z(n20357) );
  NANDN U21392 ( .A(n20334), .B(sreg[1883]), .Z(n20338) );
  NAND U21393 ( .A(n20336), .B(n20335), .Z(n20337) );
  NAND U21394 ( .A(n20338), .B(n20337), .Z(n20356) );
  XOR U21395 ( .A(n20357), .B(n20356), .Z(c[1884]) );
  NANDN U21396 ( .A(n20340), .B(n20339), .Z(n20344) );
  OR U21397 ( .A(n20342), .B(n20341), .Z(n20343) );
  AND U21398 ( .A(n20344), .B(n20343), .Z(n20362) );
  XOR U21399 ( .A(a[863]), .B(n2299), .Z(n20366) );
  AND U21400 ( .A(a[865]), .B(b[0]), .Z(n20346) );
  XNOR U21401 ( .A(n20346), .B(n2175), .Z(n20348) );
  NANDN U21402 ( .A(b[0]), .B(a[864]), .Z(n20347) );
  NAND U21403 ( .A(n20348), .B(n20347), .Z(n20371) );
  AND U21404 ( .A(a[861]), .B(b[3]), .Z(n20370) );
  XOR U21405 ( .A(n20371), .B(n20370), .Z(n20373) );
  XOR U21406 ( .A(n20372), .B(n20373), .Z(n20361) );
  NANDN U21407 ( .A(n20350), .B(n20349), .Z(n20354) );
  OR U21408 ( .A(n20352), .B(n20351), .Z(n20353) );
  AND U21409 ( .A(n20354), .B(n20353), .Z(n20360) );
  XOR U21410 ( .A(n20361), .B(n20360), .Z(n20363) );
  XOR U21411 ( .A(n20362), .B(n20363), .Z(n20376) );
  XNOR U21412 ( .A(n20376), .B(sreg[1885]), .Z(n20378) );
  NANDN U21413 ( .A(n20355), .B(sreg[1884]), .Z(n20359) );
  NAND U21414 ( .A(n20357), .B(n20356), .Z(n20358) );
  NAND U21415 ( .A(n20359), .B(n20358), .Z(n20377) );
  XOR U21416 ( .A(n20378), .B(n20377), .Z(c[1885]) );
  NANDN U21417 ( .A(n20361), .B(n20360), .Z(n20365) );
  OR U21418 ( .A(n20363), .B(n20362), .Z(n20364) );
  AND U21419 ( .A(n20365), .B(n20364), .Z(n20383) );
  XOR U21420 ( .A(a[864]), .B(n2299), .Z(n20387) );
  AND U21421 ( .A(a[866]), .B(b[0]), .Z(n20367) );
  XNOR U21422 ( .A(n20367), .B(n2175), .Z(n20369) );
  NANDN U21423 ( .A(b[0]), .B(a[865]), .Z(n20368) );
  NAND U21424 ( .A(n20369), .B(n20368), .Z(n20392) );
  AND U21425 ( .A(a[862]), .B(b[3]), .Z(n20391) );
  XOR U21426 ( .A(n20392), .B(n20391), .Z(n20394) );
  XOR U21427 ( .A(n20393), .B(n20394), .Z(n20382) );
  NANDN U21428 ( .A(n20371), .B(n20370), .Z(n20375) );
  OR U21429 ( .A(n20373), .B(n20372), .Z(n20374) );
  AND U21430 ( .A(n20375), .B(n20374), .Z(n20381) );
  XOR U21431 ( .A(n20382), .B(n20381), .Z(n20384) );
  XOR U21432 ( .A(n20383), .B(n20384), .Z(n20397) );
  XNOR U21433 ( .A(n20397), .B(sreg[1886]), .Z(n20399) );
  NANDN U21434 ( .A(n20376), .B(sreg[1885]), .Z(n20380) );
  NAND U21435 ( .A(n20378), .B(n20377), .Z(n20379) );
  NAND U21436 ( .A(n20380), .B(n20379), .Z(n20398) );
  XOR U21437 ( .A(n20399), .B(n20398), .Z(c[1886]) );
  NANDN U21438 ( .A(n20382), .B(n20381), .Z(n20386) );
  OR U21439 ( .A(n20384), .B(n20383), .Z(n20385) );
  AND U21440 ( .A(n20386), .B(n20385), .Z(n20404) );
  XOR U21441 ( .A(a[865]), .B(n2299), .Z(n20408) );
  AND U21442 ( .A(a[867]), .B(b[0]), .Z(n20388) );
  XNOR U21443 ( .A(n20388), .B(n2175), .Z(n20390) );
  NANDN U21444 ( .A(b[0]), .B(a[866]), .Z(n20389) );
  NAND U21445 ( .A(n20390), .B(n20389), .Z(n20413) );
  AND U21446 ( .A(a[863]), .B(b[3]), .Z(n20412) );
  XOR U21447 ( .A(n20413), .B(n20412), .Z(n20415) );
  XOR U21448 ( .A(n20414), .B(n20415), .Z(n20403) );
  NANDN U21449 ( .A(n20392), .B(n20391), .Z(n20396) );
  OR U21450 ( .A(n20394), .B(n20393), .Z(n20395) );
  AND U21451 ( .A(n20396), .B(n20395), .Z(n20402) );
  XOR U21452 ( .A(n20403), .B(n20402), .Z(n20405) );
  XOR U21453 ( .A(n20404), .B(n20405), .Z(n20418) );
  XNOR U21454 ( .A(n20418), .B(sreg[1887]), .Z(n20420) );
  NANDN U21455 ( .A(n20397), .B(sreg[1886]), .Z(n20401) );
  NAND U21456 ( .A(n20399), .B(n20398), .Z(n20400) );
  NAND U21457 ( .A(n20401), .B(n20400), .Z(n20419) );
  XOR U21458 ( .A(n20420), .B(n20419), .Z(c[1887]) );
  NANDN U21459 ( .A(n20403), .B(n20402), .Z(n20407) );
  OR U21460 ( .A(n20405), .B(n20404), .Z(n20406) );
  AND U21461 ( .A(n20407), .B(n20406), .Z(n20425) );
  XOR U21462 ( .A(a[866]), .B(n2299), .Z(n20429) );
  AND U21463 ( .A(a[868]), .B(b[0]), .Z(n20409) );
  XNOR U21464 ( .A(n20409), .B(n2175), .Z(n20411) );
  NANDN U21465 ( .A(b[0]), .B(a[867]), .Z(n20410) );
  NAND U21466 ( .A(n20411), .B(n20410), .Z(n20434) );
  AND U21467 ( .A(a[864]), .B(b[3]), .Z(n20433) );
  XOR U21468 ( .A(n20434), .B(n20433), .Z(n20436) );
  XOR U21469 ( .A(n20435), .B(n20436), .Z(n20424) );
  NANDN U21470 ( .A(n20413), .B(n20412), .Z(n20417) );
  OR U21471 ( .A(n20415), .B(n20414), .Z(n20416) );
  AND U21472 ( .A(n20417), .B(n20416), .Z(n20423) );
  XOR U21473 ( .A(n20424), .B(n20423), .Z(n20426) );
  XOR U21474 ( .A(n20425), .B(n20426), .Z(n20439) );
  XNOR U21475 ( .A(n20439), .B(sreg[1888]), .Z(n20441) );
  NANDN U21476 ( .A(n20418), .B(sreg[1887]), .Z(n20422) );
  NAND U21477 ( .A(n20420), .B(n20419), .Z(n20421) );
  NAND U21478 ( .A(n20422), .B(n20421), .Z(n20440) );
  XOR U21479 ( .A(n20441), .B(n20440), .Z(c[1888]) );
  NANDN U21480 ( .A(n20424), .B(n20423), .Z(n20428) );
  OR U21481 ( .A(n20426), .B(n20425), .Z(n20427) );
  AND U21482 ( .A(n20428), .B(n20427), .Z(n20446) );
  XOR U21483 ( .A(a[867]), .B(n2300), .Z(n20450) );
  AND U21484 ( .A(a[869]), .B(b[0]), .Z(n20430) );
  XNOR U21485 ( .A(n20430), .B(n2175), .Z(n20432) );
  NANDN U21486 ( .A(b[0]), .B(a[868]), .Z(n20431) );
  NAND U21487 ( .A(n20432), .B(n20431), .Z(n20455) );
  AND U21488 ( .A(a[865]), .B(b[3]), .Z(n20454) );
  XOR U21489 ( .A(n20455), .B(n20454), .Z(n20457) );
  XOR U21490 ( .A(n20456), .B(n20457), .Z(n20445) );
  NANDN U21491 ( .A(n20434), .B(n20433), .Z(n20438) );
  OR U21492 ( .A(n20436), .B(n20435), .Z(n20437) );
  AND U21493 ( .A(n20438), .B(n20437), .Z(n20444) );
  XOR U21494 ( .A(n20445), .B(n20444), .Z(n20447) );
  XOR U21495 ( .A(n20446), .B(n20447), .Z(n20460) );
  XNOR U21496 ( .A(n20460), .B(sreg[1889]), .Z(n20462) );
  NANDN U21497 ( .A(n20439), .B(sreg[1888]), .Z(n20443) );
  NAND U21498 ( .A(n20441), .B(n20440), .Z(n20442) );
  NAND U21499 ( .A(n20443), .B(n20442), .Z(n20461) );
  XOR U21500 ( .A(n20462), .B(n20461), .Z(c[1889]) );
  NANDN U21501 ( .A(n20445), .B(n20444), .Z(n20449) );
  OR U21502 ( .A(n20447), .B(n20446), .Z(n20448) );
  AND U21503 ( .A(n20449), .B(n20448), .Z(n20467) );
  XOR U21504 ( .A(a[868]), .B(n2300), .Z(n20471) );
  AND U21505 ( .A(a[870]), .B(b[0]), .Z(n20451) );
  XNOR U21506 ( .A(n20451), .B(n2175), .Z(n20453) );
  NANDN U21507 ( .A(b[0]), .B(a[869]), .Z(n20452) );
  NAND U21508 ( .A(n20453), .B(n20452), .Z(n20476) );
  AND U21509 ( .A(a[866]), .B(b[3]), .Z(n20475) );
  XOR U21510 ( .A(n20476), .B(n20475), .Z(n20478) );
  XOR U21511 ( .A(n20477), .B(n20478), .Z(n20466) );
  NANDN U21512 ( .A(n20455), .B(n20454), .Z(n20459) );
  OR U21513 ( .A(n20457), .B(n20456), .Z(n20458) );
  AND U21514 ( .A(n20459), .B(n20458), .Z(n20465) );
  XOR U21515 ( .A(n20466), .B(n20465), .Z(n20468) );
  XOR U21516 ( .A(n20467), .B(n20468), .Z(n20481) );
  XNOR U21517 ( .A(n20481), .B(sreg[1890]), .Z(n20483) );
  NANDN U21518 ( .A(n20460), .B(sreg[1889]), .Z(n20464) );
  NAND U21519 ( .A(n20462), .B(n20461), .Z(n20463) );
  NAND U21520 ( .A(n20464), .B(n20463), .Z(n20482) );
  XOR U21521 ( .A(n20483), .B(n20482), .Z(c[1890]) );
  NANDN U21522 ( .A(n20466), .B(n20465), .Z(n20470) );
  OR U21523 ( .A(n20468), .B(n20467), .Z(n20469) );
  AND U21524 ( .A(n20470), .B(n20469), .Z(n20488) );
  XOR U21525 ( .A(a[869]), .B(n2300), .Z(n20492) );
  AND U21526 ( .A(a[871]), .B(b[0]), .Z(n20472) );
  XNOR U21527 ( .A(n20472), .B(n2175), .Z(n20474) );
  NANDN U21528 ( .A(b[0]), .B(a[870]), .Z(n20473) );
  NAND U21529 ( .A(n20474), .B(n20473), .Z(n20497) );
  AND U21530 ( .A(a[867]), .B(b[3]), .Z(n20496) );
  XOR U21531 ( .A(n20497), .B(n20496), .Z(n20499) );
  XOR U21532 ( .A(n20498), .B(n20499), .Z(n20487) );
  NANDN U21533 ( .A(n20476), .B(n20475), .Z(n20480) );
  OR U21534 ( .A(n20478), .B(n20477), .Z(n20479) );
  AND U21535 ( .A(n20480), .B(n20479), .Z(n20486) );
  XOR U21536 ( .A(n20487), .B(n20486), .Z(n20489) );
  XOR U21537 ( .A(n20488), .B(n20489), .Z(n20502) );
  XNOR U21538 ( .A(n20502), .B(sreg[1891]), .Z(n20504) );
  NANDN U21539 ( .A(n20481), .B(sreg[1890]), .Z(n20485) );
  NAND U21540 ( .A(n20483), .B(n20482), .Z(n20484) );
  NAND U21541 ( .A(n20485), .B(n20484), .Z(n20503) );
  XOR U21542 ( .A(n20504), .B(n20503), .Z(c[1891]) );
  NANDN U21543 ( .A(n20487), .B(n20486), .Z(n20491) );
  OR U21544 ( .A(n20489), .B(n20488), .Z(n20490) );
  AND U21545 ( .A(n20491), .B(n20490), .Z(n20509) );
  XOR U21546 ( .A(a[870]), .B(n2300), .Z(n20513) );
  AND U21547 ( .A(a[872]), .B(b[0]), .Z(n20493) );
  XNOR U21548 ( .A(n20493), .B(n2175), .Z(n20495) );
  NANDN U21549 ( .A(b[0]), .B(a[871]), .Z(n20494) );
  NAND U21550 ( .A(n20495), .B(n20494), .Z(n20518) );
  AND U21551 ( .A(a[868]), .B(b[3]), .Z(n20517) );
  XOR U21552 ( .A(n20518), .B(n20517), .Z(n20520) );
  XOR U21553 ( .A(n20519), .B(n20520), .Z(n20508) );
  NANDN U21554 ( .A(n20497), .B(n20496), .Z(n20501) );
  OR U21555 ( .A(n20499), .B(n20498), .Z(n20500) );
  AND U21556 ( .A(n20501), .B(n20500), .Z(n20507) );
  XOR U21557 ( .A(n20508), .B(n20507), .Z(n20510) );
  XOR U21558 ( .A(n20509), .B(n20510), .Z(n20523) );
  XNOR U21559 ( .A(n20523), .B(sreg[1892]), .Z(n20525) );
  NANDN U21560 ( .A(n20502), .B(sreg[1891]), .Z(n20506) );
  NAND U21561 ( .A(n20504), .B(n20503), .Z(n20505) );
  NAND U21562 ( .A(n20506), .B(n20505), .Z(n20524) );
  XOR U21563 ( .A(n20525), .B(n20524), .Z(c[1892]) );
  NANDN U21564 ( .A(n20508), .B(n20507), .Z(n20512) );
  OR U21565 ( .A(n20510), .B(n20509), .Z(n20511) );
  AND U21566 ( .A(n20512), .B(n20511), .Z(n20530) );
  XOR U21567 ( .A(a[871]), .B(n2300), .Z(n20534) );
  AND U21568 ( .A(a[869]), .B(b[3]), .Z(n20538) );
  AND U21569 ( .A(a[873]), .B(b[0]), .Z(n20514) );
  XNOR U21570 ( .A(n20514), .B(n2175), .Z(n20516) );
  NANDN U21571 ( .A(b[0]), .B(a[872]), .Z(n20515) );
  NAND U21572 ( .A(n20516), .B(n20515), .Z(n20539) );
  XOR U21573 ( .A(n20538), .B(n20539), .Z(n20541) );
  XOR U21574 ( .A(n20540), .B(n20541), .Z(n20529) );
  NANDN U21575 ( .A(n20518), .B(n20517), .Z(n20522) );
  OR U21576 ( .A(n20520), .B(n20519), .Z(n20521) );
  AND U21577 ( .A(n20522), .B(n20521), .Z(n20528) );
  XOR U21578 ( .A(n20529), .B(n20528), .Z(n20531) );
  XOR U21579 ( .A(n20530), .B(n20531), .Z(n20544) );
  XNOR U21580 ( .A(n20544), .B(sreg[1893]), .Z(n20546) );
  NANDN U21581 ( .A(n20523), .B(sreg[1892]), .Z(n20527) );
  NAND U21582 ( .A(n20525), .B(n20524), .Z(n20526) );
  NAND U21583 ( .A(n20527), .B(n20526), .Z(n20545) );
  XOR U21584 ( .A(n20546), .B(n20545), .Z(c[1893]) );
  NANDN U21585 ( .A(n20529), .B(n20528), .Z(n20533) );
  OR U21586 ( .A(n20531), .B(n20530), .Z(n20532) );
  AND U21587 ( .A(n20533), .B(n20532), .Z(n20551) );
  XOR U21588 ( .A(a[872]), .B(n2300), .Z(n20555) );
  AND U21589 ( .A(a[874]), .B(b[0]), .Z(n20535) );
  XNOR U21590 ( .A(n20535), .B(n2175), .Z(n20537) );
  NANDN U21591 ( .A(b[0]), .B(a[873]), .Z(n20536) );
  NAND U21592 ( .A(n20537), .B(n20536), .Z(n20560) );
  AND U21593 ( .A(a[870]), .B(b[3]), .Z(n20559) );
  XOR U21594 ( .A(n20560), .B(n20559), .Z(n20562) );
  XOR U21595 ( .A(n20561), .B(n20562), .Z(n20550) );
  NANDN U21596 ( .A(n20539), .B(n20538), .Z(n20543) );
  OR U21597 ( .A(n20541), .B(n20540), .Z(n20542) );
  AND U21598 ( .A(n20543), .B(n20542), .Z(n20549) );
  XOR U21599 ( .A(n20550), .B(n20549), .Z(n20552) );
  XOR U21600 ( .A(n20551), .B(n20552), .Z(n20565) );
  XNOR U21601 ( .A(n20565), .B(sreg[1894]), .Z(n20567) );
  NANDN U21602 ( .A(n20544), .B(sreg[1893]), .Z(n20548) );
  NAND U21603 ( .A(n20546), .B(n20545), .Z(n20547) );
  NAND U21604 ( .A(n20548), .B(n20547), .Z(n20566) );
  XOR U21605 ( .A(n20567), .B(n20566), .Z(c[1894]) );
  NANDN U21606 ( .A(n20550), .B(n20549), .Z(n20554) );
  OR U21607 ( .A(n20552), .B(n20551), .Z(n20553) );
  AND U21608 ( .A(n20554), .B(n20553), .Z(n20572) );
  XOR U21609 ( .A(a[873]), .B(n2300), .Z(n20576) );
  AND U21610 ( .A(a[875]), .B(b[0]), .Z(n20556) );
  XNOR U21611 ( .A(n20556), .B(n2175), .Z(n20558) );
  NANDN U21612 ( .A(b[0]), .B(a[874]), .Z(n20557) );
  NAND U21613 ( .A(n20558), .B(n20557), .Z(n20581) );
  AND U21614 ( .A(a[871]), .B(b[3]), .Z(n20580) );
  XOR U21615 ( .A(n20581), .B(n20580), .Z(n20583) );
  XOR U21616 ( .A(n20582), .B(n20583), .Z(n20571) );
  NANDN U21617 ( .A(n20560), .B(n20559), .Z(n20564) );
  OR U21618 ( .A(n20562), .B(n20561), .Z(n20563) );
  AND U21619 ( .A(n20564), .B(n20563), .Z(n20570) );
  XOR U21620 ( .A(n20571), .B(n20570), .Z(n20573) );
  XOR U21621 ( .A(n20572), .B(n20573), .Z(n20586) );
  XNOR U21622 ( .A(n20586), .B(sreg[1895]), .Z(n20588) );
  NANDN U21623 ( .A(n20565), .B(sreg[1894]), .Z(n20569) );
  NAND U21624 ( .A(n20567), .B(n20566), .Z(n20568) );
  NAND U21625 ( .A(n20569), .B(n20568), .Z(n20587) );
  XOR U21626 ( .A(n20588), .B(n20587), .Z(c[1895]) );
  NANDN U21627 ( .A(n20571), .B(n20570), .Z(n20575) );
  OR U21628 ( .A(n20573), .B(n20572), .Z(n20574) );
  AND U21629 ( .A(n20575), .B(n20574), .Z(n20593) );
  XOR U21630 ( .A(a[874]), .B(n2301), .Z(n20597) );
  AND U21631 ( .A(a[872]), .B(b[3]), .Z(n20601) );
  AND U21632 ( .A(a[876]), .B(b[0]), .Z(n20577) );
  XNOR U21633 ( .A(n20577), .B(n2175), .Z(n20579) );
  NANDN U21634 ( .A(b[0]), .B(a[875]), .Z(n20578) );
  NAND U21635 ( .A(n20579), .B(n20578), .Z(n20602) );
  XOR U21636 ( .A(n20601), .B(n20602), .Z(n20604) );
  XOR U21637 ( .A(n20603), .B(n20604), .Z(n20592) );
  NANDN U21638 ( .A(n20581), .B(n20580), .Z(n20585) );
  OR U21639 ( .A(n20583), .B(n20582), .Z(n20584) );
  AND U21640 ( .A(n20585), .B(n20584), .Z(n20591) );
  XOR U21641 ( .A(n20592), .B(n20591), .Z(n20594) );
  XOR U21642 ( .A(n20593), .B(n20594), .Z(n20607) );
  XNOR U21643 ( .A(n20607), .B(sreg[1896]), .Z(n20609) );
  NANDN U21644 ( .A(n20586), .B(sreg[1895]), .Z(n20590) );
  NAND U21645 ( .A(n20588), .B(n20587), .Z(n20589) );
  NAND U21646 ( .A(n20590), .B(n20589), .Z(n20608) );
  XOR U21647 ( .A(n20609), .B(n20608), .Z(c[1896]) );
  NANDN U21648 ( .A(n20592), .B(n20591), .Z(n20596) );
  OR U21649 ( .A(n20594), .B(n20593), .Z(n20595) );
  AND U21650 ( .A(n20596), .B(n20595), .Z(n20614) );
  XOR U21651 ( .A(a[875]), .B(n2301), .Z(n20618) );
  AND U21652 ( .A(a[877]), .B(b[0]), .Z(n20598) );
  XNOR U21653 ( .A(n20598), .B(n2175), .Z(n20600) );
  NANDN U21654 ( .A(b[0]), .B(a[876]), .Z(n20599) );
  NAND U21655 ( .A(n20600), .B(n20599), .Z(n20623) );
  AND U21656 ( .A(a[873]), .B(b[3]), .Z(n20622) );
  XOR U21657 ( .A(n20623), .B(n20622), .Z(n20625) );
  XOR U21658 ( .A(n20624), .B(n20625), .Z(n20613) );
  NANDN U21659 ( .A(n20602), .B(n20601), .Z(n20606) );
  OR U21660 ( .A(n20604), .B(n20603), .Z(n20605) );
  AND U21661 ( .A(n20606), .B(n20605), .Z(n20612) );
  XOR U21662 ( .A(n20613), .B(n20612), .Z(n20615) );
  XOR U21663 ( .A(n20614), .B(n20615), .Z(n20628) );
  XNOR U21664 ( .A(n20628), .B(sreg[1897]), .Z(n20630) );
  NANDN U21665 ( .A(n20607), .B(sreg[1896]), .Z(n20611) );
  NAND U21666 ( .A(n20609), .B(n20608), .Z(n20610) );
  NAND U21667 ( .A(n20611), .B(n20610), .Z(n20629) );
  XOR U21668 ( .A(n20630), .B(n20629), .Z(c[1897]) );
  NANDN U21669 ( .A(n20613), .B(n20612), .Z(n20617) );
  OR U21670 ( .A(n20615), .B(n20614), .Z(n20616) );
  AND U21671 ( .A(n20617), .B(n20616), .Z(n20635) );
  XOR U21672 ( .A(a[876]), .B(n2301), .Z(n20639) );
  AND U21673 ( .A(a[874]), .B(b[3]), .Z(n20643) );
  AND U21674 ( .A(a[878]), .B(b[0]), .Z(n20619) );
  XNOR U21675 ( .A(n20619), .B(n2175), .Z(n20621) );
  NANDN U21676 ( .A(b[0]), .B(a[877]), .Z(n20620) );
  NAND U21677 ( .A(n20621), .B(n20620), .Z(n20644) );
  XOR U21678 ( .A(n20643), .B(n20644), .Z(n20646) );
  XOR U21679 ( .A(n20645), .B(n20646), .Z(n20634) );
  NANDN U21680 ( .A(n20623), .B(n20622), .Z(n20627) );
  OR U21681 ( .A(n20625), .B(n20624), .Z(n20626) );
  AND U21682 ( .A(n20627), .B(n20626), .Z(n20633) );
  XOR U21683 ( .A(n20634), .B(n20633), .Z(n20636) );
  XOR U21684 ( .A(n20635), .B(n20636), .Z(n20649) );
  XNOR U21685 ( .A(n20649), .B(sreg[1898]), .Z(n20651) );
  NANDN U21686 ( .A(n20628), .B(sreg[1897]), .Z(n20632) );
  NAND U21687 ( .A(n20630), .B(n20629), .Z(n20631) );
  NAND U21688 ( .A(n20632), .B(n20631), .Z(n20650) );
  XOR U21689 ( .A(n20651), .B(n20650), .Z(c[1898]) );
  NANDN U21690 ( .A(n20634), .B(n20633), .Z(n20638) );
  OR U21691 ( .A(n20636), .B(n20635), .Z(n20637) );
  AND U21692 ( .A(n20638), .B(n20637), .Z(n20656) );
  XOR U21693 ( .A(a[877]), .B(n2301), .Z(n20660) );
  AND U21694 ( .A(a[879]), .B(b[0]), .Z(n20640) );
  XNOR U21695 ( .A(n20640), .B(n2175), .Z(n20642) );
  NANDN U21696 ( .A(b[0]), .B(a[878]), .Z(n20641) );
  NAND U21697 ( .A(n20642), .B(n20641), .Z(n20665) );
  AND U21698 ( .A(a[875]), .B(b[3]), .Z(n20664) );
  XOR U21699 ( .A(n20665), .B(n20664), .Z(n20667) );
  XOR U21700 ( .A(n20666), .B(n20667), .Z(n20655) );
  NANDN U21701 ( .A(n20644), .B(n20643), .Z(n20648) );
  OR U21702 ( .A(n20646), .B(n20645), .Z(n20647) );
  AND U21703 ( .A(n20648), .B(n20647), .Z(n20654) );
  XOR U21704 ( .A(n20655), .B(n20654), .Z(n20657) );
  XOR U21705 ( .A(n20656), .B(n20657), .Z(n20670) );
  XNOR U21706 ( .A(n20670), .B(sreg[1899]), .Z(n20672) );
  NANDN U21707 ( .A(n20649), .B(sreg[1898]), .Z(n20653) );
  NAND U21708 ( .A(n20651), .B(n20650), .Z(n20652) );
  NAND U21709 ( .A(n20653), .B(n20652), .Z(n20671) );
  XOR U21710 ( .A(n20672), .B(n20671), .Z(c[1899]) );
  NANDN U21711 ( .A(n20655), .B(n20654), .Z(n20659) );
  OR U21712 ( .A(n20657), .B(n20656), .Z(n20658) );
  AND U21713 ( .A(n20659), .B(n20658), .Z(n20677) );
  XOR U21714 ( .A(a[878]), .B(n2301), .Z(n20681) );
  AND U21715 ( .A(a[876]), .B(b[3]), .Z(n20685) );
  AND U21716 ( .A(a[880]), .B(b[0]), .Z(n20661) );
  XNOR U21717 ( .A(n20661), .B(n2175), .Z(n20663) );
  NANDN U21718 ( .A(b[0]), .B(a[879]), .Z(n20662) );
  NAND U21719 ( .A(n20663), .B(n20662), .Z(n20686) );
  XOR U21720 ( .A(n20685), .B(n20686), .Z(n20688) );
  XOR U21721 ( .A(n20687), .B(n20688), .Z(n20676) );
  NANDN U21722 ( .A(n20665), .B(n20664), .Z(n20669) );
  OR U21723 ( .A(n20667), .B(n20666), .Z(n20668) );
  AND U21724 ( .A(n20669), .B(n20668), .Z(n20675) );
  XOR U21725 ( .A(n20676), .B(n20675), .Z(n20678) );
  XOR U21726 ( .A(n20677), .B(n20678), .Z(n20691) );
  XNOR U21727 ( .A(n20691), .B(sreg[1900]), .Z(n20693) );
  NANDN U21728 ( .A(n20670), .B(sreg[1899]), .Z(n20674) );
  NAND U21729 ( .A(n20672), .B(n20671), .Z(n20673) );
  NAND U21730 ( .A(n20674), .B(n20673), .Z(n20692) );
  XOR U21731 ( .A(n20693), .B(n20692), .Z(c[1900]) );
  NANDN U21732 ( .A(n20676), .B(n20675), .Z(n20680) );
  OR U21733 ( .A(n20678), .B(n20677), .Z(n20679) );
  AND U21734 ( .A(n20680), .B(n20679), .Z(n20698) );
  XOR U21735 ( .A(a[879]), .B(n2301), .Z(n20702) );
  AND U21736 ( .A(a[881]), .B(b[0]), .Z(n20682) );
  XNOR U21737 ( .A(n20682), .B(n2175), .Z(n20684) );
  NANDN U21738 ( .A(b[0]), .B(a[880]), .Z(n20683) );
  NAND U21739 ( .A(n20684), .B(n20683), .Z(n20707) );
  AND U21740 ( .A(a[877]), .B(b[3]), .Z(n20706) );
  XOR U21741 ( .A(n20707), .B(n20706), .Z(n20709) );
  XOR U21742 ( .A(n20708), .B(n20709), .Z(n20697) );
  NANDN U21743 ( .A(n20686), .B(n20685), .Z(n20690) );
  OR U21744 ( .A(n20688), .B(n20687), .Z(n20689) );
  AND U21745 ( .A(n20690), .B(n20689), .Z(n20696) );
  XOR U21746 ( .A(n20697), .B(n20696), .Z(n20699) );
  XOR U21747 ( .A(n20698), .B(n20699), .Z(n20712) );
  XNOR U21748 ( .A(n20712), .B(sreg[1901]), .Z(n20714) );
  NANDN U21749 ( .A(n20691), .B(sreg[1900]), .Z(n20695) );
  NAND U21750 ( .A(n20693), .B(n20692), .Z(n20694) );
  NAND U21751 ( .A(n20695), .B(n20694), .Z(n20713) );
  XOR U21752 ( .A(n20714), .B(n20713), .Z(c[1901]) );
  NANDN U21753 ( .A(n20697), .B(n20696), .Z(n20701) );
  OR U21754 ( .A(n20699), .B(n20698), .Z(n20700) );
  AND U21755 ( .A(n20701), .B(n20700), .Z(n20719) );
  XOR U21756 ( .A(a[880]), .B(n2301), .Z(n20723) );
  AND U21757 ( .A(a[882]), .B(b[0]), .Z(n20703) );
  XNOR U21758 ( .A(n20703), .B(n2175), .Z(n20705) );
  NANDN U21759 ( .A(b[0]), .B(a[881]), .Z(n20704) );
  NAND U21760 ( .A(n20705), .B(n20704), .Z(n20728) );
  AND U21761 ( .A(a[878]), .B(b[3]), .Z(n20727) );
  XOR U21762 ( .A(n20728), .B(n20727), .Z(n20730) );
  XOR U21763 ( .A(n20729), .B(n20730), .Z(n20718) );
  NANDN U21764 ( .A(n20707), .B(n20706), .Z(n20711) );
  OR U21765 ( .A(n20709), .B(n20708), .Z(n20710) );
  AND U21766 ( .A(n20711), .B(n20710), .Z(n20717) );
  XOR U21767 ( .A(n20718), .B(n20717), .Z(n20720) );
  XOR U21768 ( .A(n20719), .B(n20720), .Z(n20733) );
  XNOR U21769 ( .A(n20733), .B(sreg[1902]), .Z(n20735) );
  NANDN U21770 ( .A(n20712), .B(sreg[1901]), .Z(n20716) );
  NAND U21771 ( .A(n20714), .B(n20713), .Z(n20715) );
  NAND U21772 ( .A(n20716), .B(n20715), .Z(n20734) );
  XOR U21773 ( .A(n20735), .B(n20734), .Z(c[1902]) );
  NANDN U21774 ( .A(n20718), .B(n20717), .Z(n20722) );
  OR U21775 ( .A(n20720), .B(n20719), .Z(n20721) );
  AND U21776 ( .A(n20722), .B(n20721), .Z(n20740) );
  XOR U21777 ( .A(a[881]), .B(n2302), .Z(n20744) );
  AND U21778 ( .A(a[883]), .B(b[0]), .Z(n20724) );
  XNOR U21779 ( .A(n20724), .B(n2175), .Z(n20726) );
  NANDN U21780 ( .A(b[0]), .B(a[882]), .Z(n20725) );
  NAND U21781 ( .A(n20726), .B(n20725), .Z(n20749) );
  AND U21782 ( .A(a[879]), .B(b[3]), .Z(n20748) );
  XOR U21783 ( .A(n20749), .B(n20748), .Z(n20751) );
  XOR U21784 ( .A(n20750), .B(n20751), .Z(n20739) );
  NANDN U21785 ( .A(n20728), .B(n20727), .Z(n20732) );
  OR U21786 ( .A(n20730), .B(n20729), .Z(n20731) );
  AND U21787 ( .A(n20732), .B(n20731), .Z(n20738) );
  XOR U21788 ( .A(n20739), .B(n20738), .Z(n20741) );
  XOR U21789 ( .A(n20740), .B(n20741), .Z(n20754) );
  XNOR U21790 ( .A(n20754), .B(sreg[1903]), .Z(n20756) );
  NANDN U21791 ( .A(n20733), .B(sreg[1902]), .Z(n20737) );
  NAND U21792 ( .A(n20735), .B(n20734), .Z(n20736) );
  NAND U21793 ( .A(n20737), .B(n20736), .Z(n20755) );
  XOR U21794 ( .A(n20756), .B(n20755), .Z(c[1903]) );
  NANDN U21795 ( .A(n20739), .B(n20738), .Z(n20743) );
  OR U21796 ( .A(n20741), .B(n20740), .Z(n20742) );
  AND U21797 ( .A(n20743), .B(n20742), .Z(n20761) );
  XOR U21798 ( .A(a[882]), .B(n2302), .Z(n20765) );
  AND U21799 ( .A(a[884]), .B(b[0]), .Z(n20745) );
  XNOR U21800 ( .A(n20745), .B(n2175), .Z(n20747) );
  NANDN U21801 ( .A(b[0]), .B(a[883]), .Z(n20746) );
  NAND U21802 ( .A(n20747), .B(n20746), .Z(n20770) );
  AND U21803 ( .A(a[880]), .B(b[3]), .Z(n20769) );
  XOR U21804 ( .A(n20770), .B(n20769), .Z(n20772) );
  XOR U21805 ( .A(n20771), .B(n20772), .Z(n20760) );
  NANDN U21806 ( .A(n20749), .B(n20748), .Z(n20753) );
  OR U21807 ( .A(n20751), .B(n20750), .Z(n20752) );
  AND U21808 ( .A(n20753), .B(n20752), .Z(n20759) );
  XOR U21809 ( .A(n20760), .B(n20759), .Z(n20762) );
  XOR U21810 ( .A(n20761), .B(n20762), .Z(n20775) );
  XNOR U21811 ( .A(n20775), .B(sreg[1904]), .Z(n20777) );
  NANDN U21812 ( .A(n20754), .B(sreg[1903]), .Z(n20758) );
  NAND U21813 ( .A(n20756), .B(n20755), .Z(n20757) );
  NAND U21814 ( .A(n20758), .B(n20757), .Z(n20776) );
  XOR U21815 ( .A(n20777), .B(n20776), .Z(c[1904]) );
  NANDN U21816 ( .A(n20760), .B(n20759), .Z(n20764) );
  OR U21817 ( .A(n20762), .B(n20761), .Z(n20763) );
  AND U21818 ( .A(n20764), .B(n20763), .Z(n20782) );
  XOR U21819 ( .A(a[883]), .B(n2302), .Z(n20786) );
  AND U21820 ( .A(a[881]), .B(b[3]), .Z(n20790) );
  AND U21821 ( .A(a[885]), .B(b[0]), .Z(n20766) );
  XNOR U21822 ( .A(n20766), .B(n2175), .Z(n20768) );
  NANDN U21823 ( .A(b[0]), .B(a[884]), .Z(n20767) );
  NAND U21824 ( .A(n20768), .B(n20767), .Z(n20791) );
  XOR U21825 ( .A(n20790), .B(n20791), .Z(n20793) );
  XOR U21826 ( .A(n20792), .B(n20793), .Z(n20781) );
  NANDN U21827 ( .A(n20770), .B(n20769), .Z(n20774) );
  OR U21828 ( .A(n20772), .B(n20771), .Z(n20773) );
  AND U21829 ( .A(n20774), .B(n20773), .Z(n20780) );
  XOR U21830 ( .A(n20781), .B(n20780), .Z(n20783) );
  XOR U21831 ( .A(n20782), .B(n20783), .Z(n20796) );
  XNOR U21832 ( .A(n20796), .B(sreg[1905]), .Z(n20798) );
  NANDN U21833 ( .A(n20775), .B(sreg[1904]), .Z(n20779) );
  NAND U21834 ( .A(n20777), .B(n20776), .Z(n20778) );
  NAND U21835 ( .A(n20779), .B(n20778), .Z(n20797) );
  XOR U21836 ( .A(n20798), .B(n20797), .Z(c[1905]) );
  NANDN U21837 ( .A(n20781), .B(n20780), .Z(n20785) );
  OR U21838 ( .A(n20783), .B(n20782), .Z(n20784) );
  AND U21839 ( .A(n20785), .B(n20784), .Z(n20803) );
  XOR U21840 ( .A(a[884]), .B(n2302), .Z(n20807) );
  AND U21841 ( .A(a[886]), .B(b[0]), .Z(n20787) );
  XNOR U21842 ( .A(n20787), .B(n2175), .Z(n20789) );
  NANDN U21843 ( .A(b[0]), .B(a[885]), .Z(n20788) );
  NAND U21844 ( .A(n20789), .B(n20788), .Z(n20812) );
  AND U21845 ( .A(a[882]), .B(b[3]), .Z(n20811) );
  XOR U21846 ( .A(n20812), .B(n20811), .Z(n20814) );
  XOR U21847 ( .A(n20813), .B(n20814), .Z(n20802) );
  NANDN U21848 ( .A(n20791), .B(n20790), .Z(n20795) );
  OR U21849 ( .A(n20793), .B(n20792), .Z(n20794) );
  AND U21850 ( .A(n20795), .B(n20794), .Z(n20801) );
  XOR U21851 ( .A(n20802), .B(n20801), .Z(n20804) );
  XOR U21852 ( .A(n20803), .B(n20804), .Z(n20817) );
  XNOR U21853 ( .A(n20817), .B(sreg[1906]), .Z(n20819) );
  NANDN U21854 ( .A(n20796), .B(sreg[1905]), .Z(n20800) );
  NAND U21855 ( .A(n20798), .B(n20797), .Z(n20799) );
  NAND U21856 ( .A(n20800), .B(n20799), .Z(n20818) );
  XOR U21857 ( .A(n20819), .B(n20818), .Z(c[1906]) );
  NANDN U21858 ( .A(n20802), .B(n20801), .Z(n20806) );
  OR U21859 ( .A(n20804), .B(n20803), .Z(n20805) );
  AND U21860 ( .A(n20806), .B(n20805), .Z(n20824) );
  XOR U21861 ( .A(a[885]), .B(n2302), .Z(n20828) );
  AND U21862 ( .A(a[883]), .B(b[3]), .Z(n20832) );
  AND U21863 ( .A(a[887]), .B(b[0]), .Z(n20808) );
  XNOR U21864 ( .A(n20808), .B(n2175), .Z(n20810) );
  NANDN U21865 ( .A(b[0]), .B(a[886]), .Z(n20809) );
  NAND U21866 ( .A(n20810), .B(n20809), .Z(n20833) );
  XOR U21867 ( .A(n20832), .B(n20833), .Z(n20835) );
  XOR U21868 ( .A(n20834), .B(n20835), .Z(n20823) );
  NANDN U21869 ( .A(n20812), .B(n20811), .Z(n20816) );
  OR U21870 ( .A(n20814), .B(n20813), .Z(n20815) );
  AND U21871 ( .A(n20816), .B(n20815), .Z(n20822) );
  XOR U21872 ( .A(n20823), .B(n20822), .Z(n20825) );
  XOR U21873 ( .A(n20824), .B(n20825), .Z(n20838) );
  XNOR U21874 ( .A(n20838), .B(sreg[1907]), .Z(n20840) );
  NANDN U21875 ( .A(n20817), .B(sreg[1906]), .Z(n20821) );
  NAND U21876 ( .A(n20819), .B(n20818), .Z(n20820) );
  NAND U21877 ( .A(n20821), .B(n20820), .Z(n20839) );
  XOR U21878 ( .A(n20840), .B(n20839), .Z(c[1907]) );
  NANDN U21879 ( .A(n20823), .B(n20822), .Z(n20827) );
  OR U21880 ( .A(n20825), .B(n20824), .Z(n20826) );
  AND U21881 ( .A(n20827), .B(n20826), .Z(n20845) );
  XOR U21882 ( .A(a[886]), .B(n2302), .Z(n20849) );
  AND U21883 ( .A(a[884]), .B(b[3]), .Z(n20853) );
  AND U21884 ( .A(a[888]), .B(b[0]), .Z(n20829) );
  XNOR U21885 ( .A(n20829), .B(n2175), .Z(n20831) );
  NANDN U21886 ( .A(b[0]), .B(a[887]), .Z(n20830) );
  NAND U21887 ( .A(n20831), .B(n20830), .Z(n20854) );
  XOR U21888 ( .A(n20853), .B(n20854), .Z(n20856) );
  XOR U21889 ( .A(n20855), .B(n20856), .Z(n20844) );
  NANDN U21890 ( .A(n20833), .B(n20832), .Z(n20837) );
  OR U21891 ( .A(n20835), .B(n20834), .Z(n20836) );
  AND U21892 ( .A(n20837), .B(n20836), .Z(n20843) );
  XOR U21893 ( .A(n20844), .B(n20843), .Z(n20846) );
  XOR U21894 ( .A(n20845), .B(n20846), .Z(n20859) );
  XNOR U21895 ( .A(n20859), .B(sreg[1908]), .Z(n20861) );
  NANDN U21896 ( .A(n20838), .B(sreg[1907]), .Z(n20842) );
  NAND U21897 ( .A(n20840), .B(n20839), .Z(n20841) );
  NAND U21898 ( .A(n20842), .B(n20841), .Z(n20860) );
  XOR U21899 ( .A(n20861), .B(n20860), .Z(c[1908]) );
  NANDN U21900 ( .A(n20844), .B(n20843), .Z(n20848) );
  OR U21901 ( .A(n20846), .B(n20845), .Z(n20847) );
  AND U21902 ( .A(n20848), .B(n20847), .Z(n20866) );
  XOR U21903 ( .A(a[887]), .B(n2302), .Z(n20870) );
  AND U21904 ( .A(a[889]), .B(b[0]), .Z(n20850) );
  XNOR U21905 ( .A(n20850), .B(n2175), .Z(n20852) );
  NANDN U21906 ( .A(b[0]), .B(a[888]), .Z(n20851) );
  NAND U21907 ( .A(n20852), .B(n20851), .Z(n20875) );
  AND U21908 ( .A(a[885]), .B(b[3]), .Z(n20874) );
  XOR U21909 ( .A(n20875), .B(n20874), .Z(n20877) );
  XOR U21910 ( .A(n20876), .B(n20877), .Z(n20865) );
  NANDN U21911 ( .A(n20854), .B(n20853), .Z(n20858) );
  OR U21912 ( .A(n20856), .B(n20855), .Z(n20857) );
  AND U21913 ( .A(n20858), .B(n20857), .Z(n20864) );
  XOR U21914 ( .A(n20865), .B(n20864), .Z(n20867) );
  XOR U21915 ( .A(n20866), .B(n20867), .Z(n20880) );
  XNOR U21916 ( .A(n20880), .B(sreg[1909]), .Z(n20882) );
  NANDN U21917 ( .A(n20859), .B(sreg[1908]), .Z(n20863) );
  NAND U21918 ( .A(n20861), .B(n20860), .Z(n20862) );
  NAND U21919 ( .A(n20863), .B(n20862), .Z(n20881) );
  XOR U21920 ( .A(n20882), .B(n20881), .Z(c[1909]) );
  NANDN U21921 ( .A(n20865), .B(n20864), .Z(n20869) );
  OR U21922 ( .A(n20867), .B(n20866), .Z(n20868) );
  AND U21923 ( .A(n20869), .B(n20868), .Z(n20887) );
  XOR U21924 ( .A(a[888]), .B(n2303), .Z(n20891) );
  AND U21925 ( .A(a[886]), .B(b[3]), .Z(n20895) );
  AND U21926 ( .A(a[890]), .B(b[0]), .Z(n20871) );
  XNOR U21927 ( .A(n20871), .B(n2175), .Z(n20873) );
  NANDN U21928 ( .A(b[0]), .B(a[889]), .Z(n20872) );
  NAND U21929 ( .A(n20873), .B(n20872), .Z(n20896) );
  XOR U21930 ( .A(n20895), .B(n20896), .Z(n20898) );
  XOR U21931 ( .A(n20897), .B(n20898), .Z(n20886) );
  NANDN U21932 ( .A(n20875), .B(n20874), .Z(n20879) );
  OR U21933 ( .A(n20877), .B(n20876), .Z(n20878) );
  AND U21934 ( .A(n20879), .B(n20878), .Z(n20885) );
  XOR U21935 ( .A(n20886), .B(n20885), .Z(n20888) );
  XOR U21936 ( .A(n20887), .B(n20888), .Z(n20901) );
  XNOR U21937 ( .A(n20901), .B(sreg[1910]), .Z(n20903) );
  NANDN U21938 ( .A(n20880), .B(sreg[1909]), .Z(n20884) );
  NAND U21939 ( .A(n20882), .B(n20881), .Z(n20883) );
  NAND U21940 ( .A(n20884), .B(n20883), .Z(n20902) );
  XOR U21941 ( .A(n20903), .B(n20902), .Z(c[1910]) );
  NANDN U21942 ( .A(n20886), .B(n20885), .Z(n20890) );
  OR U21943 ( .A(n20888), .B(n20887), .Z(n20889) );
  AND U21944 ( .A(n20890), .B(n20889), .Z(n20908) );
  XOR U21945 ( .A(a[889]), .B(n2303), .Z(n20912) );
  AND U21946 ( .A(a[891]), .B(b[0]), .Z(n20892) );
  XNOR U21947 ( .A(n20892), .B(n2175), .Z(n20894) );
  NANDN U21948 ( .A(b[0]), .B(a[890]), .Z(n20893) );
  NAND U21949 ( .A(n20894), .B(n20893), .Z(n20917) );
  AND U21950 ( .A(a[887]), .B(b[3]), .Z(n20916) );
  XOR U21951 ( .A(n20917), .B(n20916), .Z(n20919) );
  XOR U21952 ( .A(n20918), .B(n20919), .Z(n20907) );
  NANDN U21953 ( .A(n20896), .B(n20895), .Z(n20900) );
  OR U21954 ( .A(n20898), .B(n20897), .Z(n20899) );
  AND U21955 ( .A(n20900), .B(n20899), .Z(n20906) );
  XOR U21956 ( .A(n20907), .B(n20906), .Z(n20909) );
  XOR U21957 ( .A(n20908), .B(n20909), .Z(n20922) );
  XNOR U21958 ( .A(n20922), .B(sreg[1911]), .Z(n20924) );
  NANDN U21959 ( .A(n20901), .B(sreg[1910]), .Z(n20905) );
  NAND U21960 ( .A(n20903), .B(n20902), .Z(n20904) );
  NAND U21961 ( .A(n20905), .B(n20904), .Z(n20923) );
  XOR U21962 ( .A(n20924), .B(n20923), .Z(c[1911]) );
  NANDN U21963 ( .A(n20907), .B(n20906), .Z(n20911) );
  OR U21964 ( .A(n20909), .B(n20908), .Z(n20910) );
  AND U21965 ( .A(n20911), .B(n20910), .Z(n20929) );
  XOR U21966 ( .A(a[890]), .B(n2303), .Z(n20933) );
  AND U21967 ( .A(a[892]), .B(b[0]), .Z(n20913) );
  XNOR U21968 ( .A(n20913), .B(n2175), .Z(n20915) );
  NANDN U21969 ( .A(b[0]), .B(a[891]), .Z(n20914) );
  NAND U21970 ( .A(n20915), .B(n20914), .Z(n20938) );
  AND U21971 ( .A(a[888]), .B(b[3]), .Z(n20937) );
  XOR U21972 ( .A(n20938), .B(n20937), .Z(n20940) );
  XOR U21973 ( .A(n20939), .B(n20940), .Z(n20928) );
  NANDN U21974 ( .A(n20917), .B(n20916), .Z(n20921) );
  OR U21975 ( .A(n20919), .B(n20918), .Z(n20920) );
  AND U21976 ( .A(n20921), .B(n20920), .Z(n20927) );
  XOR U21977 ( .A(n20928), .B(n20927), .Z(n20930) );
  XOR U21978 ( .A(n20929), .B(n20930), .Z(n20943) );
  XNOR U21979 ( .A(n20943), .B(sreg[1912]), .Z(n20945) );
  NANDN U21980 ( .A(n20922), .B(sreg[1911]), .Z(n20926) );
  NAND U21981 ( .A(n20924), .B(n20923), .Z(n20925) );
  NAND U21982 ( .A(n20926), .B(n20925), .Z(n20944) );
  XOR U21983 ( .A(n20945), .B(n20944), .Z(c[1912]) );
  NANDN U21984 ( .A(n20928), .B(n20927), .Z(n20932) );
  OR U21985 ( .A(n20930), .B(n20929), .Z(n20931) );
  AND U21986 ( .A(n20932), .B(n20931), .Z(n20950) );
  XOR U21987 ( .A(a[891]), .B(n2303), .Z(n20954) );
  AND U21988 ( .A(a[889]), .B(b[3]), .Z(n20958) );
  AND U21989 ( .A(a[893]), .B(b[0]), .Z(n20934) );
  XNOR U21990 ( .A(n20934), .B(n2175), .Z(n20936) );
  NANDN U21991 ( .A(b[0]), .B(a[892]), .Z(n20935) );
  NAND U21992 ( .A(n20936), .B(n20935), .Z(n20959) );
  XOR U21993 ( .A(n20958), .B(n20959), .Z(n20961) );
  XOR U21994 ( .A(n20960), .B(n20961), .Z(n20949) );
  NANDN U21995 ( .A(n20938), .B(n20937), .Z(n20942) );
  OR U21996 ( .A(n20940), .B(n20939), .Z(n20941) );
  AND U21997 ( .A(n20942), .B(n20941), .Z(n20948) );
  XOR U21998 ( .A(n20949), .B(n20948), .Z(n20951) );
  XOR U21999 ( .A(n20950), .B(n20951), .Z(n20964) );
  XNOR U22000 ( .A(n20964), .B(sreg[1913]), .Z(n20966) );
  NANDN U22001 ( .A(n20943), .B(sreg[1912]), .Z(n20947) );
  NAND U22002 ( .A(n20945), .B(n20944), .Z(n20946) );
  NAND U22003 ( .A(n20947), .B(n20946), .Z(n20965) );
  XOR U22004 ( .A(n20966), .B(n20965), .Z(c[1913]) );
  NANDN U22005 ( .A(n20949), .B(n20948), .Z(n20953) );
  OR U22006 ( .A(n20951), .B(n20950), .Z(n20952) );
  AND U22007 ( .A(n20953), .B(n20952), .Z(n20971) );
  XOR U22008 ( .A(a[892]), .B(n2303), .Z(n20975) );
  AND U22009 ( .A(a[894]), .B(b[0]), .Z(n20955) );
  XNOR U22010 ( .A(n20955), .B(n2175), .Z(n20957) );
  NANDN U22011 ( .A(b[0]), .B(a[893]), .Z(n20956) );
  NAND U22012 ( .A(n20957), .B(n20956), .Z(n20980) );
  AND U22013 ( .A(a[890]), .B(b[3]), .Z(n20979) );
  XOR U22014 ( .A(n20980), .B(n20979), .Z(n20982) );
  XOR U22015 ( .A(n20981), .B(n20982), .Z(n20970) );
  NANDN U22016 ( .A(n20959), .B(n20958), .Z(n20963) );
  OR U22017 ( .A(n20961), .B(n20960), .Z(n20962) );
  AND U22018 ( .A(n20963), .B(n20962), .Z(n20969) );
  XOR U22019 ( .A(n20970), .B(n20969), .Z(n20972) );
  XOR U22020 ( .A(n20971), .B(n20972), .Z(n20985) );
  XNOR U22021 ( .A(n20985), .B(sreg[1914]), .Z(n20987) );
  NANDN U22022 ( .A(n20964), .B(sreg[1913]), .Z(n20968) );
  NAND U22023 ( .A(n20966), .B(n20965), .Z(n20967) );
  NAND U22024 ( .A(n20968), .B(n20967), .Z(n20986) );
  XOR U22025 ( .A(n20987), .B(n20986), .Z(c[1914]) );
  NANDN U22026 ( .A(n20970), .B(n20969), .Z(n20974) );
  OR U22027 ( .A(n20972), .B(n20971), .Z(n20973) );
  AND U22028 ( .A(n20974), .B(n20973), .Z(n20992) );
  XOR U22029 ( .A(a[893]), .B(n2303), .Z(n20996) );
  AND U22030 ( .A(a[895]), .B(b[0]), .Z(n20976) );
  XNOR U22031 ( .A(n20976), .B(n2175), .Z(n20978) );
  NANDN U22032 ( .A(b[0]), .B(a[894]), .Z(n20977) );
  NAND U22033 ( .A(n20978), .B(n20977), .Z(n21001) );
  AND U22034 ( .A(a[891]), .B(b[3]), .Z(n21000) );
  XOR U22035 ( .A(n21001), .B(n21000), .Z(n21003) );
  XOR U22036 ( .A(n21002), .B(n21003), .Z(n20991) );
  NANDN U22037 ( .A(n20980), .B(n20979), .Z(n20984) );
  OR U22038 ( .A(n20982), .B(n20981), .Z(n20983) );
  AND U22039 ( .A(n20984), .B(n20983), .Z(n20990) );
  XOR U22040 ( .A(n20991), .B(n20990), .Z(n20993) );
  XOR U22041 ( .A(n20992), .B(n20993), .Z(n21006) );
  XNOR U22042 ( .A(n21006), .B(sreg[1915]), .Z(n21008) );
  NANDN U22043 ( .A(n20985), .B(sreg[1914]), .Z(n20989) );
  NAND U22044 ( .A(n20987), .B(n20986), .Z(n20988) );
  NAND U22045 ( .A(n20989), .B(n20988), .Z(n21007) );
  XOR U22046 ( .A(n21008), .B(n21007), .Z(c[1915]) );
  NANDN U22047 ( .A(n20991), .B(n20990), .Z(n20995) );
  OR U22048 ( .A(n20993), .B(n20992), .Z(n20994) );
  AND U22049 ( .A(n20995), .B(n20994), .Z(n21013) );
  XOR U22050 ( .A(a[894]), .B(n2303), .Z(n21017) );
  AND U22051 ( .A(a[896]), .B(b[0]), .Z(n20997) );
  XNOR U22052 ( .A(n20997), .B(n2175), .Z(n20999) );
  NANDN U22053 ( .A(b[0]), .B(a[895]), .Z(n20998) );
  NAND U22054 ( .A(n20999), .B(n20998), .Z(n21022) );
  AND U22055 ( .A(a[892]), .B(b[3]), .Z(n21021) );
  XOR U22056 ( .A(n21022), .B(n21021), .Z(n21024) );
  XOR U22057 ( .A(n21023), .B(n21024), .Z(n21012) );
  NANDN U22058 ( .A(n21001), .B(n21000), .Z(n21005) );
  OR U22059 ( .A(n21003), .B(n21002), .Z(n21004) );
  AND U22060 ( .A(n21005), .B(n21004), .Z(n21011) );
  XOR U22061 ( .A(n21012), .B(n21011), .Z(n21014) );
  XOR U22062 ( .A(n21013), .B(n21014), .Z(n21027) );
  XNOR U22063 ( .A(n21027), .B(sreg[1916]), .Z(n21029) );
  NANDN U22064 ( .A(n21006), .B(sreg[1915]), .Z(n21010) );
  NAND U22065 ( .A(n21008), .B(n21007), .Z(n21009) );
  NAND U22066 ( .A(n21010), .B(n21009), .Z(n21028) );
  XOR U22067 ( .A(n21029), .B(n21028), .Z(c[1916]) );
  NANDN U22068 ( .A(n21012), .B(n21011), .Z(n21016) );
  OR U22069 ( .A(n21014), .B(n21013), .Z(n21015) );
  AND U22070 ( .A(n21016), .B(n21015), .Z(n21035) );
  XOR U22071 ( .A(a[895]), .B(n2304), .Z(n21036) );
  AND U22072 ( .A(b[0]), .B(a[897]), .Z(n21018) );
  XOR U22073 ( .A(b[1]), .B(n21018), .Z(n21020) );
  NANDN U22074 ( .A(b[0]), .B(a[896]), .Z(n21019) );
  AND U22075 ( .A(n21020), .B(n21019), .Z(n21040) );
  AND U22076 ( .A(a[893]), .B(b[3]), .Z(n21041) );
  XOR U22077 ( .A(n21040), .B(n21041), .Z(n21042) );
  XNOR U22078 ( .A(n21043), .B(n21042), .Z(n21032) );
  NANDN U22079 ( .A(n21022), .B(n21021), .Z(n21026) );
  OR U22080 ( .A(n21024), .B(n21023), .Z(n21025) );
  AND U22081 ( .A(n21026), .B(n21025), .Z(n21033) );
  XNOR U22082 ( .A(n21032), .B(n21033), .Z(n21034) );
  XNOR U22083 ( .A(n21035), .B(n21034), .Z(n21046) );
  XNOR U22084 ( .A(n21046), .B(sreg[1917]), .Z(n21048) );
  NANDN U22085 ( .A(n21027), .B(sreg[1916]), .Z(n21031) );
  NAND U22086 ( .A(n21029), .B(n21028), .Z(n21030) );
  NAND U22087 ( .A(n21031), .B(n21030), .Z(n21047) );
  XOR U22088 ( .A(n21048), .B(n21047), .Z(c[1917]) );
  XOR U22089 ( .A(a[896]), .B(n2304), .Z(n21055) );
  AND U22090 ( .A(a[898]), .B(b[0]), .Z(n21037) );
  XNOR U22091 ( .A(n21037), .B(n2175), .Z(n21039) );
  NANDN U22092 ( .A(b[0]), .B(a[897]), .Z(n21038) );
  NAND U22093 ( .A(n21039), .B(n21038), .Z(n21060) );
  AND U22094 ( .A(a[894]), .B(b[3]), .Z(n21059) );
  XOR U22095 ( .A(n21060), .B(n21059), .Z(n21062) );
  XOR U22096 ( .A(n21061), .B(n21062), .Z(n21050) );
  NAND U22097 ( .A(n21041), .B(n21040), .Z(n21045) );
  NANDN U22098 ( .A(n21043), .B(n21042), .Z(n21044) );
  AND U22099 ( .A(n21045), .B(n21044), .Z(n21049) );
  XOR U22100 ( .A(n21050), .B(n21049), .Z(n21052) );
  XOR U22101 ( .A(n21051), .B(n21052), .Z(n21065) );
  XNOR U22102 ( .A(n21065), .B(sreg[1918]), .Z(n21067) );
  XOR U22103 ( .A(n21067), .B(n21066), .Z(c[1918]) );
  NANDN U22104 ( .A(n21050), .B(n21049), .Z(n21054) );
  OR U22105 ( .A(n21052), .B(n21051), .Z(n21053) );
  AND U22106 ( .A(n21054), .B(n21053), .Z(n21072) );
  XOR U22107 ( .A(a[897]), .B(n2304), .Z(n21076) );
  AND U22108 ( .A(a[899]), .B(b[0]), .Z(n21056) );
  XNOR U22109 ( .A(n21056), .B(n2175), .Z(n21058) );
  NANDN U22110 ( .A(b[0]), .B(a[898]), .Z(n21057) );
  NAND U22111 ( .A(n21058), .B(n21057), .Z(n21081) );
  AND U22112 ( .A(a[895]), .B(b[3]), .Z(n21080) );
  XOR U22113 ( .A(n21081), .B(n21080), .Z(n21083) );
  XOR U22114 ( .A(n21082), .B(n21083), .Z(n21071) );
  NANDN U22115 ( .A(n21060), .B(n21059), .Z(n21064) );
  OR U22116 ( .A(n21062), .B(n21061), .Z(n21063) );
  AND U22117 ( .A(n21064), .B(n21063), .Z(n21070) );
  XOR U22118 ( .A(n21071), .B(n21070), .Z(n21073) );
  XOR U22119 ( .A(n21072), .B(n21073), .Z(n21086) );
  XNOR U22120 ( .A(n21086), .B(sreg[1919]), .Z(n21088) );
  NANDN U22121 ( .A(n21065), .B(sreg[1918]), .Z(n21069) );
  NAND U22122 ( .A(n21067), .B(n21066), .Z(n21068) );
  NAND U22123 ( .A(n21069), .B(n21068), .Z(n21087) );
  XOR U22124 ( .A(n21088), .B(n21087), .Z(c[1919]) );
  NANDN U22125 ( .A(n21071), .B(n21070), .Z(n21075) );
  OR U22126 ( .A(n21073), .B(n21072), .Z(n21074) );
  AND U22127 ( .A(n21075), .B(n21074), .Z(n21093) );
  XOR U22128 ( .A(a[898]), .B(n2304), .Z(n21097) );
  AND U22129 ( .A(a[896]), .B(b[3]), .Z(n21101) );
  AND U22130 ( .A(a[900]), .B(b[0]), .Z(n21077) );
  XNOR U22131 ( .A(n21077), .B(n2175), .Z(n21079) );
  NANDN U22132 ( .A(b[0]), .B(a[899]), .Z(n21078) );
  NAND U22133 ( .A(n21079), .B(n21078), .Z(n21102) );
  XOR U22134 ( .A(n21101), .B(n21102), .Z(n21104) );
  XOR U22135 ( .A(n21103), .B(n21104), .Z(n21092) );
  NANDN U22136 ( .A(n21081), .B(n21080), .Z(n21085) );
  OR U22137 ( .A(n21083), .B(n21082), .Z(n21084) );
  AND U22138 ( .A(n21085), .B(n21084), .Z(n21091) );
  XOR U22139 ( .A(n21092), .B(n21091), .Z(n21094) );
  XOR U22140 ( .A(n21093), .B(n21094), .Z(n21107) );
  XNOR U22141 ( .A(n21107), .B(sreg[1920]), .Z(n21109) );
  NANDN U22142 ( .A(n21086), .B(sreg[1919]), .Z(n21090) );
  NAND U22143 ( .A(n21088), .B(n21087), .Z(n21089) );
  NAND U22144 ( .A(n21090), .B(n21089), .Z(n21108) );
  XOR U22145 ( .A(n21109), .B(n21108), .Z(c[1920]) );
  NANDN U22146 ( .A(n21092), .B(n21091), .Z(n21096) );
  OR U22147 ( .A(n21094), .B(n21093), .Z(n21095) );
  AND U22148 ( .A(n21096), .B(n21095), .Z(n21114) );
  XOR U22149 ( .A(a[899]), .B(n2304), .Z(n21118) );
  AND U22150 ( .A(a[901]), .B(b[0]), .Z(n21098) );
  XNOR U22151 ( .A(n21098), .B(n2175), .Z(n21100) );
  NANDN U22152 ( .A(b[0]), .B(a[900]), .Z(n21099) );
  NAND U22153 ( .A(n21100), .B(n21099), .Z(n21123) );
  AND U22154 ( .A(a[897]), .B(b[3]), .Z(n21122) );
  XOR U22155 ( .A(n21123), .B(n21122), .Z(n21125) );
  XOR U22156 ( .A(n21124), .B(n21125), .Z(n21113) );
  NANDN U22157 ( .A(n21102), .B(n21101), .Z(n21106) );
  OR U22158 ( .A(n21104), .B(n21103), .Z(n21105) );
  AND U22159 ( .A(n21106), .B(n21105), .Z(n21112) );
  XOR U22160 ( .A(n21113), .B(n21112), .Z(n21115) );
  XOR U22161 ( .A(n21114), .B(n21115), .Z(n21128) );
  XNOR U22162 ( .A(n21128), .B(sreg[1921]), .Z(n21130) );
  NANDN U22163 ( .A(n21107), .B(sreg[1920]), .Z(n21111) );
  NAND U22164 ( .A(n21109), .B(n21108), .Z(n21110) );
  NAND U22165 ( .A(n21111), .B(n21110), .Z(n21129) );
  XOR U22166 ( .A(n21130), .B(n21129), .Z(c[1921]) );
  NANDN U22167 ( .A(n21113), .B(n21112), .Z(n21117) );
  OR U22168 ( .A(n21115), .B(n21114), .Z(n21116) );
  AND U22169 ( .A(n21117), .B(n21116), .Z(n21135) );
  XOR U22170 ( .A(a[900]), .B(n2304), .Z(n21139) );
  AND U22171 ( .A(a[902]), .B(b[0]), .Z(n21119) );
  XNOR U22172 ( .A(n21119), .B(n2175), .Z(n21121) );
  NANDN U22173 ( .A(b[0]), .B(a[901]), .Z(n21120) );
  NAND U22174 ( .A(n21121), .B(n21120), .Z(n21144) );
  AND U22175 ( .A(a[898]), .B(b[3]), .Z(n21143) );
  XOR U22176 ( .A(n21144), .B(n21143), .Z(n21146) );
  XOR U22177 ( .A(n21145), .B(n21146), .Z(n21134) );
  NANDN U22178 ( .A(n21123), .B(n21122), .Z(n21127) );
  OR U22179 ( .A(n21125), .B(n21124), .Z(n21126) );
  AND U22180 ( .A(n21127), .B(n21126), .Z(n21133) );
  XOR U22181 ( .A(n21134), .B(n21133), .Z(n21136) );
  XOR U22182 ( .A(n21135), .B(n21136), .Z(n21149) );
  XNOR U22183 ( .A(n21149), .B(sreg[1922]), .Z(n21151) );
  NANDN U22184 ( .A(n21128), .B(sreg[1921]), .Z(n21132) );
  NAND U22185 ( .A(n21130), .B(n21129), .Z(n21131) );
  NAND U22186 ( .A(n21132), .B(n21131), .Z(n21150) );
  XOR U22187 ( .A(n21151), .B(n21150), .Z(c[1922]) );
  NANDN U22188 ( .A(n21134), .B(n21133), .Z(n21138) );
  OR U22189 ( .A(n21136), .B(n21135), .Z(n21137) );
  AND U22190 ( .A(n21138), .B(n21137), .Z(n21156) );
  XOR U22191 ( .A(a[901]), .B(n2304), .Z(n21160) );
  AND U22192 ( .A(a[903]), .B(b[0]), .Z(n21140) );
  XNOR U22193 ( .A(n21140), .B(n2175), .Z(n21142) );
  NANDN U22194 ( .A(b[0]), .B(a[902]), .Z(n21141) );
  NAND U22195 ( .A(n21142), .B(n21141), .Z(n21165) );
  AND U22196 ( .A(a[899]), .B(b[3]), .Z(n21164) );
  XOR U22197 ( .A(n21165), .B(n21164), .Z(n21167) );
  XOR U22198 ( .A(n21166), .B(n21167), .Z(n21155) );
  NANDN U22199 ( .A(n21144), .B(n21143), .Z(n21148) );
  OR U22200 ( .A(n21146), .B(n21145), .Z(n21147) );
  AND U22201 ( .A(n21148), .B(n21147), .Z(n21154) );
  XOR U22202 ( .A(n21155), .B(n21154), .Z(n21157) );
  XOR U22203 ( .A(n21156), .B(n21157), .Z(n21170) );
  XNOR U22204 ( .A(n21170), .B(sreg[1923]), .Z(n21172) );
  NANDN U22205 ( .A(n21149), .B(sreg[1922]), .Z(n21153) );
  NAND U22206 ( .A(n21151), .B(n21150), .Z(n21152) );
  NAND U22207 ( .A(n21153), .B(n21152), .Z(n21171) );
  XOR U22208 ( .A(n21172), .B(n21171), .Z(c[1923]) );
  NANDN U22209 ( .A(n21155), .B(n21154), .Z(n21159) );
  OR U22210 ( .A(n21157), .B(n21156), .Z(n21158) );
  AND U22211 ( .A(n21159), .B(n21158), .Z(n21177) );
  XOR U22212 ( .A(a[902]), .B(n2305), .Z(n21181) );
  AND U22213 ( .A(a[900]), .B(b[3]), .Z(n21185) );
  AND U22214 ( .A(a[904]), .B(b[0]), .Z(n21161) );
  XNOR U22215 ( .A(n21161), .B(n2175), .Z(n21163) );
  NANDN U22216 ( .A(b[0]), .B(a[903]), .Z(n21162) );
  NAND U22217 ( .A(n21163), .B(n21162), .Z(n21186) );
  XOR U22218 ( .A(n21185), .B(n21186), .Z(n21188) );
  XOR U22219 ( .A(n21187), .B(n21188), .Z(n21176) );
  NANDN U22220 ( .A(n21165), .B(n21164), .Z(n21169) );
  OR U22221 ( .A(n21167), .B(n21166), .Z(n21168) );
  AND U22222 ( .A(n21169), .B(n21168), .Z(n21175) );
  XOR U22223 ( .A(n21176), .B(n21175), .Z(n21178) );
  XOR U22224 ( .A(n21177), .B(n21178), .Z(n21191) );
  XNOR U22225 ( .A(n21191), .B(sreg[1924]), .Z(n21193) );
  NANDN U22226 ( .A(n21170), .B(sreg[1923]), .Z(n21174) );
  NAND U22227 ( .A(n21172), .B(n21171), .Z(n21173) );
  NAND U22228 ( .A(n21174), .B(n21173), .Z(n21192) );
  XOR U22229 ( .A(n21193), .B(n21192), .Z(c[1924]) );
  NANDN U22230 ( .A(n21176), .B(n21175), .Z(n21180) );
  OR U22231 ( .A(n21178), .B(n21177), .Z(n21179) );
  AND U22232 ( .A(n21180), .B(n21179), .Z(n21198) );
  XOR U22233 ( .A(a[903]), .B(n2305), .Z(n21202) );
  AND U22234 ( .A(a[901]), .B(b[3]), .Z(n21206) );
  AND U22235 ( .A(a[905]), .B(b[0]), .Z(n21182) );
  XNOR U22236 ( .A(n21182), .B(n2175), .Z(n21184) );
  NANDN U22237 ( .A(b[0]), .B(a[904]), .Z(n21183) );
  NAND U22238 ( .A(n21184), .B(n21183), .Z(n21207) );
  XOR U22239 ( .A(n21206), .B(n21207), .Z(n21209) );
  XOR U22240 ( .A(n21208), .B(n21209), .Z(n21197) );
  NANDN U22241 ( .A(n21186), .B(n21185), .Z(n21190) );
  OR U22242 ( .A(n21188), .B(n21187), .Z(n21189) );
  AND U22243 ( .A(n21190), .B(n21189), .Z(n21196) );
  XOR U22244 ( .A(n21197), .B(n21196), .Z(n21199) );
  XOR U22245 ( .A(n21198), .B(n21199), .Z(n21212) );
  XNOR U22246 ( .A(n21212), .B(sreg[1925]), .Z(n21214) );
  NANDN U22247 ( .A(n21191), .B(sreg[1924]), .Z(n21195) );
  NAND U22248 ( .A(n21193), .B(n21192), .Z(n21194) );
  NAND U22249 ( .A(n21195), .B(n21194), .Z(n21213) );
  XOR U22250 ( .A(n21214), .B(n21213), .Z(c[1925]) );
  NANDN U22251 ( .A(n21197), .B(n21196), .Z(n21201) );
  OR U22252 ( .A(n21199), .B(n21198), .Z(n21200) );
  AND U22253 ( .A(n21201), .B(n21200), .Z(n21219) );
  XOR U22254 ( .A(a[904]), .B(n2305), .Z(n21223) );
  AND U22255 ( .A(a[906]), .B(b[0]), .Z(n21203) );
  XNOR U22256 ( .A(n21203), .B(n2175), .Z(n21205) );
  NANDN U22257 ( .A(b[0]), .B(a[905]), .Z(n21204) );
  NAND U22258 ( .A(n21205), .B(n21204), .Z(n21228) );
  AND U22259 ( .A(a[902]), .B(b[3]), .Z(n21227) );
  XOR U22260 ( .A(n21228), .B(n21227), .Z(n21230) );
  XOR U22261 ( .A(n21229), .B(n21230), .Z(n21218) );
  NANDN U22262 ( .A(n21207), .B(n21206), .Z(n21211) );
  OR U22263 ( .A(n21209), .B(n21208), .Z(n21210) );
  AND U22264 ( .A(n21211), .B(n21210), .Z(n21217) );
  XOR U22265 ( .A(n21218), .B(n21217), .Z(n21220) );
  XOR U22266 ( .A(n21219), .B(n21220), .Z(n21233) );
  XNOR U22267 ( .A(n21233), .B(sreg[1926]), .Z(n21235) );
  NANDN U22268 ( .A(n21212), .B(sreg[1925]), .Z(n21216) );
  NAND U22269 ( .A(n21214), .B(n21213), .Z(n21215) );
  NAND U22270 ( .A(n21216), .B(n21215), .Z(n21234) );
  XOR U22271 ( .A(n21235), .B(n21234), .Z(c[1926]) );
  NANDN U22272 ( .A(n21218), .B(n21217), .Z(n21222) );
  OR U22273 ( .A(n21220), .B(n21219), .Z(n21221) );
  AND U22274 ( .A(n21222), .B(n21221), .Z(n21240) );
  XOR U22275 ( .A(a[905]), .B(n2305), .Z(n21244) );
  AND U22276 ( .A(a[907]), .B(b[0]), .Z(n21224) );
  XNOR U22277 ( .A(n21224), .B(n2175), .Z(n21226) );
  NANDN U22278 ( .A(b[0]), .B(a[906]), .Z(n21225) );
  NAND U22279 ( .A(n21226), .B(n21225), .Z(n21249) );
  AND U22280 ( .A(a[903]), .B(b[3]), .Z(n21248) );
  XOR U22281 ( .A(n21249), .B(n21248), .Z(n21251) );
  XOR U22282 ( .A(n21250), .B(n21251), .Z(n21239) );
  NANDN U22283 ( .A(n21228), .B(n21227), .Z(n21232) );
  OR U22284 ( .A(n21230), .B(n21229), .Z(n21231) );
  AND U22285 ( .A(n21232), .B(n21231), .Z(n21238) );
  XOR U22286 ( .A(n21239), .B(n21238), .Z(n21241) );
  XOR U22287 ( .A(n21240), .B(n21241), .Z(n21254) );
  XNOR U22288 ( .A(n21254), .B(sreg[1927]), .Z(n21256) );
  NANDN U22289 ( .A(n21233), .B(sreg[1926]), .Z(n21237) );
  NAND U22290 ( .A(n21235), .B(n21234), .Z(n21236) );
  NAND U22291 ( .A(n21237), .B(n21236), .Z(n21255) );
  XOR U22292 ( .A(n21256), .B(n21255), .Z(c[1927]) );
  NANDN U22293 ( .A(n21239), .B(n21238), .Z(n21243) );
  OR U22294 ( .A(n21241), .B(n21240), .Z(n21242) );
  AND U22295 ( .A(n21243), .B(n21242), .Z(n21261) );
  XOR U22296 ( .A(a[906]), .B(n2305), .Z(n21265) );
  AND U22297 ( .A(a[908]), .B(b[0]), .Z(n21245) );
  XNOR U22298 ( .A(n21245), .B(n2175), .Z(n21247) );
  NANDN U22299 ( .A(b[0]), .B(a[907]), .Z(n21246) );
  NAND U22300 ( .A(n21247), .B(n21246), .Z(n21270) );
  AND U22301 ( .A(a[904]), .B(b[3]), .Z(n21269) );
  XOR U22302 ( .A(n21270), .B(n21269), .Z(n21272) );
  XOR U22303 ( .A(n21271), .B(n21272), .Z(n21260) );
  NANDN U22304 ( .A(n21249), .B(n21248), .Z(n21253) );
  OR U22305 ( .A(n21251), .B(n21250), .Z(n21252) );
  AND U22306 ( .A(n21253), .B(n21252), .Z(n21259) );
  XOR U22307 ( .A(n21260), .B(n21259), .Z(n21262) );
  XOR U22308 ( .A(n21261), .B(n21262), .Z(n21275) );
  XNOR U22309 ( .A(n21275), .B(sreg[1928]), .Z(n21277) );
  NANDN U22310 ( .A(n21254), .B(sreg[1927]), .Z(n21258) );
  NAND U22311 ( .A(n21256), .B(n21255), .Z(n21257) );
  NAND U22312 ( .A(n21258), .B(n21257), .Z(n21276) );
  XOR U22313 ( .A(n21277), .B(n21276), .Z(c[1928]) );
  NANDN U22314 ( .A(n21260), .B(n21259), .Z(n21264) );
  OR U22315 ( .A(n21262), .B(n21261), .Z(n21263) );
  AND U22316 ( .A(n21264), .B(n21263), .Z(n21283) );
  XOR U22317 ( .A(a[907]), .B(n2305), .Z(n21284) );
  NAND U22318 ( .A(a[909]), .B(b[0]), .Z(n21266) );
  XNOR U22319 ( .A(b[1]), .B(n21266), .Z(n21268) );
  NANDN U22320 ( .A(b[0]), .B(a[908]), .Z(n21267) );
  AND U22321 ( .A(n21268), .B(n21267), .Z(n21288) );
  AND U22322 ( .A(a[905]), .B(b[3]), .Z(n21289) );
  XOR U22323 ( .A(n21288), .B(n21289), .Z(n21290) );
  XNOR U22324 ( .A(n21291), .B(n21290), .Z(n21280) );
  NANDN U22325 ( .A(n21270), .B(n21269), .Z(n21274) );
  OR U22326 ( .A(n21272), .B(n21271), .Z(n21273) );
  AND U22327 ( .A(n21274), .B(n21273), .Z(n21281) );
  XNOR U22328 ( .A(n21280), .B(n21281), .Z(n21282) );
  XNOR U22329 ( .A(n21283), .B(n21282), .Z(n21294) );
  XNOR U22330 ( .A(n21294), .B(sreg[1929]), .Z(n21296) );
  NANDN U22331 ( .A(n21275), .B(sreg[1928]), .Z(n21279) );
  NAND U22332 ( .A(n21277), .B(n21276), .Z(n21278) );
  NAND U22333 ( .A(n21279), .B(n21278), .Z(n21295) );
  XOR U22334 ( .A(n21296), .B(n21295), .Z(c[1929]) );
  XOR U22335 ( .A(a[908]), .B(n2305), .Z(n21303) );
  AND U22336 ( .A(a[910]), .B(b[0]), .Z(n21285) );
  XNOR U22337 ( .A(n21285), .B(n2175), .Z(n21287) );
  NANDN U22338 ( .A(b[0]), .B(a[909]), .Z(n21286) );
  NAND U22339 ( .A(n21287), .B(n21286), .Z(n21308) );
  AND U22340 ( .A(a[906]), .B(b[3]), .Z(n21307) );
  XOR U22341 ( .A(n21308), .B(n21307), .Z(n21310) );
  XOR U22342 ( .A(n21309), .B(n21310), .Z(n21298) );
  NAND U22343 ( .A(n21289), .B(n21288), .Z(n21293) );
  NANDN U22344 ( .A(n21291), .B(n21290), .Z(n21292) );
  AND U22345 ( .A(n21293), .B(n21292), .Z(n21297) );
  XOR U22346 ( .A(n21298), .B(n21297), .Z(n21300) );
  XOR U22347 ( .A(n21299), .B(n21300), .Z(n21313) );
  XNOR U22348 ( .A(n21313), .B(sreg[1930]), .Z(n21315) );
  XOR U22349 ( .A(n21315), .B(n21314), .Z(c[1930]) );
  NANDN U22350 ( .A(n21298), .B(n21297), .Z(n21302) );
  OR U22351 ( .A(n21300), .B(n21299), .Z(n21301) );
  AND U22352 ( .A(n21302), .B(n21301), .Z(n21320) );
  XOR U22353 ( .A(a[909]), .B(n2306), .Z(n21324) );
  AND U22354 ( .A(a[911]), .B(b[0]), .Z(n21304) );
  XNOR U22355 ( .A(n21304), .B(n2175), .Z(n21306) );
  NANDN U22356 ( .A(b[0]), .B(a[910]), .Z(n21305) );
  NAND U22357 ( .A(n21306), .B(n21305), .Z(n21329) );
  AND U22358 ( .A(a[907]), .B(b[3]), .Z(n21328) );
  XOR U22359 ( .A(n21329), .B(n21328), .Z(n21331) );
  XOR U22360 ( .A(n21330), .B(n21331), .Z(n21319) );
  NANDN U22361 ( .A(n21308), .B(n21307), .Z(n21312) );
  OR U22362 ( .A(n21310), .B(n21309), .Z(n21311) );
  AND U22363 ( .A(n21312), .B(n21311), .Z(n21318) );
  XOR U22364 ( .A(n21319), .B(n21318), .Z(n21321) );
  XOR U22365 ( .A(n21320), .B(n21321), .Z(n21334) );
  XNOR U22366 ( .A(n21334), .B(sreg[1931]), .Z(n21336) );
  NANDN U22367 ( .A(n21313), .B(sreg[1930]), .Z(n21317) );
  NAND U22368 ( .A(n21315), .B(n21314), .Z(n21316) );
  NAND U22369 ( .A(n21317), .B(n21316), .Z(n21335) );
  XOR U22370 ( .A(n21336), .B(n21335), .Z(c[1931]) );
  NANDN U22371 ( .A(n21319), .B(n21318), .Z(n21323) );
  OR U22372 ( .A(n21321), .B(n21320), .Z(n21322) );
  AND U22373 ( .A(n21323), .B(n21322), .Z(n21341) );
  XOR U22374 ( .A(a[910]), .B(n2306), .Z(n21345) );
  AND U22375 ( .A(a[908]), .B(b[3]), .Z(n21349) );
  AND U22376 ( .A(a[912]), .B(b[0]), .Z(n21325) );
  XNOR U22377 ( .A(n21325), .B(n2175), .Z(n21327) );
  NANDN U22378 ( .A(b[0]), .B(a[911]), .Z(n21326) );
  NAND U22379 ( .A(n21327), .B(n21326), .Z(n21350) );
  XOR U22380 ( .A(n21349), .B(n21350), .Z(n21352) );
  XOR U22381 ( .A(n21351), .B(n21352), .Z(n21340) );
  NANDN U22382 ( .A(n21329), .B(n21328), .Z(n21333) );
  OR U22383 ( .A(n21331), .B(n21330), .Z(n21332) );
  AND U22384 ( .A(n21333), .B(n21332), .Z(n21339) );
  XOR U22385 ( .A(n21340), .B(n21339), .Z(n21342) );
  XOR U22386 ( .A(n21341), .B(n21342), .Z(n21355) );
  XNOR U22387 ( .A(n21355), .B(sreg[1932]), .Z(n21357) );
  NANDN U22388 ( .A(n21334), .B(sreg[1931]), .Z(n21338) );
  NAND U22389 ( .A(n21336), .B(n21335), .Z(n21337) );
  NAND U22390 ( .A(n21338), .B(n21337), .Z(n21356) );
  XOR U22391 ( .A(n21357), .B(n21356), .Z(c[1932]) );
  NANDN U22392 ( .A(n21340), .B(n21339), .Z(n21344) );
  OR U22393 ( .A(n21342), .B(n21341), .Z(n21343) );
  AND U22394 ( .A(n21344), .B(n21343), .Z(n21362) );
  XOR U22395 ( .A(a[911]), .B(n2306), .Z(n21366) );
  AND U22396 ( .A(a[913]), .B(b[0]), .Z(n21346) );
  XNOR U22397 ( .A(n21346), .B(n2175), .Z(n21348) );
  NANDN U22398 ( .A(b[0]), .B(a[912]), .Z(n21347) );
  NAND U22399 ( .A(n21348), .B(n21347), .Z(n21371) );
  AND U22400 ( .A(a[909]), .B(b[3]), .Z(n21370) );
  XOR U22401 ( .A(n21371), .B(n21370), .Z(n21373) );
  XOR U22402 ( .A(n21372), .B(n21373), .Z(n21361) );
  NANDN U22403 ( .A(n21350), .B(n21349), .Z(n21354) );
  OR U22404 ( .A(n21352), .B(n21351), .Z(n21353) );
  AND U22405 ( .A(n21354), .B(n21353), .Z(n21360) );
  XOR U22406 ( .A(n21361), .B(n21360), .Z(n21363) );
  XOR U22407 ( .A(n21362), .B(n21363), .Z(n21376) );
  XNOR U22408 ( .A(n21376), .B(sreg[1933]), .Z(n21378) );
  NANDN U22409 ( .A(n21355), .B(sreg[1932]), .Z(n21359) );
  NAND U22410 ( .A(n21357), .B(n21356), .Z(n21358) );
  NAND U22411 ( .A(n21359), .B(n21358), .Z(n21377) );
  XOR U22412 ( .A(n21378), .B(n21377), .Z(c[1933]) );
  NANDN U22413 ( .A(n21361), .B(n21360), .Z(n21365) );
  OR U22414 ( .A(n21363), .B(n21362), .Z(n21364) );
  AND U22415 ( .A(n21365), .B(n21364), .Z(n21383) );
  XOR U22416 ( .A(a[912]), .B(n2306), .Z(n21387) );
  AND U22417 ( .A(a[914]), .B(b[0]), .Z(n21367) );
  XNOR U22418 ( .A(n21367), .B(n2175), .Z(n21369) );
  NANDN U22419 ( .A(b[0]), .B(a[913]), .Z(n21368) );
  NAND U22420 ( .A(n21369), .B(n21368), .Z(n21392) );
  AND U22421 ( .A(a[910]), .B(b[3]), .Z(n21391) );
  XOR U22422 ( .A(n21392), .B(n21391), .Z(n21394) );
  XOR U22423 ( .A(n21393), .B(n21394), .Z(n21382) );
  NANDN U22424 ( .A(n21371), .B(n21370), .Z(n21375) );
  OR U22425 ( .A(n21373), .B(n21372), .Z(n21374) );
  AND U22426 ( .A(n21375), .B(n21374), .Z(n21381) );
  XOR U22427 ( .A(n21382), .B(n21381), .Z(n21384) );
  XOR U22428 ( .A(n21383), .B(n21384), .Z(n21397) );
  XNOR U22429 ( .A(n21397), .B(sreg[1934]), .Z(n21399) );
  NANDN U22430 ( .A(n21376), .B(sreg[1933]), .Z(n21380) );
  NAND U22431 ( .A(n21378), .B(n21377), .Z(n21379) );
  NAND U22432 ( .A(n21380), .B(n21379), .Z(n21398) );
  XOR U22433 ( .A(n21399), .B(n21398), .Z(c[1934]) );
  NANDN U22434 ( .A(n21382), .B(n21381), .Z(n21386) );
  OR U22435 ( .A(n21384), .B(n21383), .Z(n21385) );
  AND U22436 ( .A(n21386), .B(n21385), .Z(n21404) );
  XOR U22437 ( .A(a[913]), .B(n2306), .Z(n21408) );
  AND U22438 ( .A(a[915]), .B(b[0]), .Z(n21388) );
  XNOR U22439 ( .A(n21388), .B(n2175), .Z(n21390) );
  NANDN U22440 ( .A(b[0]), .B(a[914]), .Z(n21389) );
  NAND U22441 ( .A(n21390), .B(n21389), .Z(n21413) );
  AND U22442 ( .A(a[911]), .B(b[3]), .Z(n21412) );
  XOR U22443 ( .A(n21413), .B(n21412), .Z(n21415) );
  XOR U22444 ( .A(n21414), .B(n21415), .Z(n21403) );
  NANDN U22445 ( .A(n21392), .B(n21391), .Z(n21396) );
  OR U22446 ( .A(n21394), .B(n21393), .Z(n21395) );
  AND U22447 ( .A(n21396), .B(n21395), .Z(n21402) );
  XOR U22448 ( .A(n21403), .B(n21402), .Z(n21405) );
  XOR U22449 ( .A(n21404), .B(n21405), .Z(n21418) );
  XNOR U22450 ( .A(n21418), .B(sreg[1935]), .Z(n21420) );
  NANDN U22451 ( .A(n21397), .B(sreg[1934]), .Z(n21401) );
  NAND U22452 ( .A(n21399), .B(n21398), .Z(n21400) );
  NAND U22453 ( .A(n21401), .B(n21400), .Z(n21419) );
  XOR U22454 ( .A(n21420), .B(n21419), .Z(c[1935]) );
  NANDN U22455 ( .A(n21403), .B(n21402), .Z(n21407) );
  OR U22456 ( .A(n21405), .B(n21404), .Z(n21406) );
  AND U22457 ( .A(n21407), .B(n21406), .Z(n21425) );
  XOR U22458 ( .A(a[914]), .B(n2306), .Z(n21429) );
  AND U22459 ( .A(a[916]), .B(b[0]), .Z(n21409) );
  XNOR U22460 ( .A(n21409), .B(n2175), .Z(n21411) );
  NANDN U22461 ( .A(b[0]), .B(a[915]), .Z(n21410) );
  NAND U22462 ( .A(n21411), .B(n21410), .Z(n21434) );
  AND U22463 ( .A(a[912]), .B(b[3]), .Z(n21433) );
  XOR U22464 ( .A(n21434), .B(n21433), .Z(n21436) );
  XOR U22465 ( .A(n21435), .B(n21436), .Z(n21424) );
  NANDN U22466 ( .A(n21413), .B(n21412), .Z(n21417) );
  OR U22467 ( .A(n21415), .B(n21414), .Z(n21416) );
  AND U22468 ( .A(n21417), .B(n21416), .Z(n21423) );
  XOR U22469 ( .A(n21424), .B(n21423), .Z(n21426) );
  XOR U22470 ( .A(n21425), .B(n21426), .Z(n21439) );
  XNOR U22471 ( .A(n21439), .B(sreg[1936]), .Z(n21441) );
  NANDN U22472 ( .A(n21418), .B(sreg[1935]), .Z(n21422) );
  NAND U22473 ( .A(n21420), .B(n21419), .Z(n21421) );
  NAND U22474 ( .A(n21422), .B(n21421), .Z(n21440) );
  XOR U22475 ( .A(n21441), .B(n21440), .Z(c[1936]) );
  NANDN U22476 ( .A(n21424), .B(n21423), .Z(n21428) );
  OR U22477 ( .A(n21426), .B(n21425), .Z(n21427) );
  AND U22478 ( .A(n21428), .B(n21427), .Z(n21446) );
  XOR U22479 ( .A(a[915]), .B(n2306), .Z(n21450) );
  AND U22480 ( .A(a[917]), .B(b[0]), .Z(n21430) );
  XNOR U22481 ( .A(n21430), .B(n2175), .Z(n21432) );
  NANDN U22482 ( .A(b[0]), .B(a[916]), .Z(n21431) );
  NAND U22483 ( .A(n21432), .B(n21431), .Z(n21455) );
  AND U22484 ( .A(a[913]), .B(b[3]), .Z(n21454) );
  XOR U22485 ( .A(n21455), .B(n21454), .Z(n21457) );
  XOR U22486 ( .A(n21456), .B(n21457), .Z(n21445) );
  NANDN U22487 ( .A(n21434), .B(n21433), .Z(n21438) );
  OR U22488 ( .A(n21436), .B(n21435), .Z(n21437) );
  AND U22489 ( .A(n21438), .B(n21437), .Z(n21444) );
  XOR U22490 ( .A(n21445), .B(n21444), .Z(n21447) );
  XOR U22491 ( .A(n21446), .B(n21447), .Z(n21460) );
  XNOR U22492 ( .A(n21460), .B(sreg[1937]), .Z(n21462) );
  NANDN U22493 ( .A(n21439), .B(sreg[1936]), .Z(n21443) );
  NAND U22494 ( .A(n21441), .B(n21440), .Z(n21442) );
  NAND U22495 ( .A(n21443), .B(n21442), .Z(n21461) );
  XOR U22496 ( .A(n21462), .B(n21461), .Z(c[1937]) );
  NANDN U22497 ( .A(n21445), .B(n21444), .Z(n21449) );
  OR U22498 ( .A(n21447), .B(n21446), .Z(n21448) );
  AND U22499 ( .A(n21449), .B(n21448), .Z(n21467) );
  XOR U22500 ( .A(a[916]), .B(n2307), .Z(n21471) );
  AND U22501 ( .A(a[918]), .B(b[0]), .Z(n21451) );
  XNOR U22502 ( .A(n21451), .B(n2175), .Z(n21453) );
  NANDN U22503 ( .A(b[0]), .B(a[917]), .Z(n21452) );
  NAND U22504 ( .A(n21453), .B(n21452), .Z(n21476) );
  AND U22505 ( .A(a[914]), .B(b[3]), .Z(n21475) );
  XOR U22506 ( .A(n21476), .B(n21475), .Z(n21478) );
  XOR U22507 ( .A(n21477), .B(n21478), .Z(n21466) );
  NANDN U22508 ( .A(n21455), .B(n21454), .Z(n21459) );
  OR U22509 ( .A(n21457), .B(n21456), .Z(n21458) );
  AND U22510 ( .A(n21459), .B(n21458), .Z(n21465) );
  XOR U22511 ( .A(n21466), .B(n21465), .Z(n21468) );
  XOR U22512 ( .A(n21467), .B(n21468), .Z(n21481) );
  XNOR U22513 ( .A(n21481), .B(sreg[1938]), .Z(n21483) );
  NANDN U22514 ( .A(n21460), .B(sreg[1937]), .Z(n21464) );
  NAND U22515 ( .A(n21462), .B(n21461), .Z(n21463) );
  NAND U22516 ( .A(n21464), .B(n21463), .Z(n21482) );
  XOR U22517 ( .A(n21483), .B(n21482), .Z(c[1938]) );
  NANDN U22518 ( .A(n21466), .B(n21465), .Z(n21470) );
  OR U22519 ( .A(n21468), .B(n21467), .Z(n21469) );
  AND U22520 ( .A(n21470), .B(n21469), .Z(n21488) );
  XOR U22521 ( .A(a[917]), .B(n2307), .Z(n21492) );
  AND U22522 ( .A(a[919]), .B(b[0]), .Z(n21472) );
  XNOR U22523 ( .A(n21472), .B(n2175), .Z(n21474) );
  NANDN U22524 ( .A(b[0]), .B(a[918]), .Z(n21473) );
  NAND U22525 ( .A(n21474), .B(n21473), .Z(n21497) );
  AND U22526 ( .A(a[915]), .B(b[3]), .Z(n21496) );
  XOR U22527 ( .A(n21497), .B(n21496), .Z(n21499) );
  XOR U22528 ( .A(n21498), .B(n21499), .Z(n21487) );
  NANDN U22529 ( .A(n21476), .B(n21475), .Z(n21480) );
  OR U22530 ( .A(n21478), .B(n21477), .Z(n21479) );
  AND U22531 ( .A(n21480), .B(n21479), .Z(n21486) );
  XOR U22532 ( .A(n21487), .B(n21486), .Z(n21489) );
  XOR U22533 ( .A(n21488), .B(n21489), .Z(n21502) );
  XNOR U22534 ( .A(n21502), .B(sreg[1939]), .Z(n21504) );
  NANDN U22535 ( .A(n21481), .B(sreg[1938]), .Z(n21485) );
  NAND U22536 ( .A(n21483), .B(n21482), .Z(n21484) );
  NAND U22537 ( .A(n21485), .B(n21484), .Z(n21503) );
  XOR U22538 ( .A(n21504), .B(n21503), .Z(c[1939]) );
  NANDN U22539 ( .A(n21487), .B(n21486), .Z(n21491) );
  OR U22540 ( .A(n21489), .B(n21488), .Z(n21490) );
  AND U22541 ( .A(n21491), .B(n21490), .Z(n21509) );
  XOR U22542 ( .A(a[918]), .B(n2307), .Z(n21513) );
  AND U22543 ( .A(a[920]), .B(b[0]), .Z(n21493) );
  XNOR U22544 ( .A(n21493), .B(n2175), .Z(n21495) );
  NANDN U22545 ( .A(b[0]), .B(a[919]), .Z(n21494) );
  NAND U22546 ( .A(n21495), .B(n21494), .Z(n21518) );
  AND U22547 ( .A(a[916]), .B(b[3]), .Z(n21517) );
  XOR U22548 ( .A(n21518), .B(n21517), .Z(n21520) );
  XOR U22549 ( .A(n21519), .B(n21520), .Z(n21508) );
  NANDN U22550 ( .A(n21497), .B(n21496), .Z(n21501) );
  OR U22551 ( .A(n21499), .B(n21498), .Z(n21500) );
  AND U22552 ( .A(n21501), .B(n21500), .Z(n21507) );
  XOR U22553 ( .A(n21508), .B(n21507), .Z(n21510) );
  XOR U22554 ( .A(n21509), .B(n21510), .Z(n21523) );
  XNOR U22555 ( .A(n21523), .B(sreg[1940]), .Z(n21525) );
  NANDN U22556 ( .A(n21502), .B(sreg[1939]), .Z(n21506) );
  NAND U22557 ( .A(n21504), .B(n21503), .Z(n21505) );
  NAND U22558 ( .A(n21506), .B(n21505), .Z(n21524) );
  XOR U22559 ( .A(n21525), .B(n21524), .Z(c[1940]) );
  NANDN U22560 ( .A(n21508), .B(n21507), .Z(n21512) );
  OR U22561 ( .A(n21510), .B(n21509), .Z(n21511) );
  AND U22562 ( .A(n21512), .B(n21511), .Z(n21530) );
  XOR U22563 ( .A(a[919]), .B(n2307), .Z(n21534) );
  AND U22564 ( .A(a[921]), .B(b[0]), .Z(n21514) );
  XNOR U22565 ( .A(n21514), .B(n2175), .Z(n21516) );
  NANDN U22566 ( .A(b[0]), .B(a[920]), .Z(n21515) );
  NAND U22567 ( .A(n21516), .B(n21515), .Z(n21539) );
  AND U22568 ( .A(a[917]), .B(b[3]), .Z(n21538) );
  XOR U22569 ( .A(n21539), .B(n21538), .Z(n21541) );
  XOR U22570 ( .A(n21540), .B(n21541), .Z(n21529) );
  NANDN U22571 ( .A(n21518), .B(n21517), .Z(n21522) );
  OR U22572 ( .A(n21520), .B(n21519), .Z(n21521) );
  AND U22573 ( .A(n21522), .B(n21521), .Z(n21528) );
  XOR U22574 ( .A(n21529), .B(n21528), .Z(n21531) );
  XOR U22575 ( .A(n21530), .B(n21531), .Z(n21544) );
  XNOR U22576 ( .A(n21544), .B(sreg[1941]), .Z(n21546) );
  NANDN U22577 ( .A(n21523), .B(sreg[1940]), .Z(n21527) );
  NAND U22578 ( .A(n21525), .B(n21524), .Z(n21526) );
  NAND U22579 ( .A(n21527), .B(n21526), .Z(n21545) );
  XOR U22580 ( .A(n21546), .B(n21545), .Z(c[1941]) );
  NANDN U22581 ( .A(n21529), .B(n21528), .Z(n21533) );
  OR U22582 ( .A(n21531), .B(n21530), .Z(n21532) );
  AND U22583 ( .A(n21533), .B(n21532), .Z(n21551) );
  XOR U22584 ( .A(a[920]), .B(n2307), .Z(n21555) );
  AND U22585 ( .A(a[922]), .B(b[0]), .Z(n21535) );
  XNOR U22586 ( .A(n21535), .B(n2175), .Z(n21537) );
  NANDN U22587 ( .A(b[0]), .B(a[921]), .Z(n21536) );
  NAND U22588 ( .A(n21537), .B(n21536), .Z(n21560) );
  AND U22589 ( .A(a[918]), .B(b[3]), .Z(n21559) );
  XOR U22590 ( .A(n21560), .B(n21559), .Z(n21562) );
  XOR U22591 ( .A(n21561), .B(n21562), .Z(n21550) );
  NANDN U22592 ( .A(n21539), .B(n21538), .Z(n21543) );
  OR U22593 ( .A(n21541), .B(n21540), .Z(n21542) );
  AND U22594 ( .A(n21543), .B(n21542), .Z(n21549) );
  XOR U22595 ( .A(n21550), .B(n21549), .Z(n21552) );
  XOR U22596 ( .A(n21551), .B(n21552), .Z(n21565) );
  XNOR U22597 ( .A(n21565), .B(sreg[1942]), .Z(n21567) );
  NANDN U22598 ( .A(n21544), .B(sreg[1941]), .Z(n21548) );
  NAND U22599 ( .A(n21546), .B(n21545), .Z(n21547) );
  NAND U22600 ( .A(n21548), .B(n21547), .Z(n21566) );
  XOR U22601 ( .A(n21567), .B(n21566), .Z(c[1942]) );
  NANDN U22602 ( .A(n21550), .B(n21549), .Z(n21554) );
  OR U22603 ( .A(n21552), .B(n21551), .Z(n21553) );
  AND U22604 ( .A(n21554), .B(n21553), .Z(n21572) );
  XOR U22605 ( .A(a[921]), .B(n2307), .Z(n21576) );
  AND U22606 ( .A(a[923]), .B(b[0]), .Z(n21556) );
  XNOR U22607 ( .A(n21556), .B(n2175), .Z(n21558) );
  NANDN U22608 ( .A(b[0]), .B(a[922]), .Z(n21557) );
  NAND U22609 ( .A(n21558), .B(n21557), .Z(n21581) );
  AND U22610 ( .A(a[919]), .B(b[3]), .Z(n21580) );
  XOR U22611 ( .A(n21581), .B(n21580), .Z(n21583) );
  XOR U22612 ( .A(n21582), .B(n21583), .Z(n21571) );
  NANDN U22613 ( .A(n21560), .B(n21559), .Z(n21564) );
  OR U22614 ( .A(n21562), .B(n21561), .Z(n21563) );
  AND U22615 ( .A(n21564), .B(n21563), .Z(n21570) );
  XOR U22616 ( .A(n21571), .B(n21570), .Z(n21573) );
  XOR U22617 ( .A(n21572), .B(n21573), .Z(n21586) );
  XNOR U22618 ( .A(n21586), .B(sreg[1943]), .Z(n21588) );
  NANDN U22619 ( .A(n21565), .B(sreg[1942]), .Z(n21569) );
  NAND U22620 ( .A(n21567), .B(n21566), .Z(n21568) );
  NAND U22621 ( .A(n21569), .B(n21568), .Z(n21587) );
  XOR U22622 ( .A(n21588), .B(n21587), .Z(c[1943]) );
  NANDN U22623 ( .A(n21571), .B(n21570), .Z(n21575) );
  OR U22624 ( .A(n21573), .B(n21572), .Z(n21574) );
  AND U22625 ( .A(n21575), .B(n21574), .Z(n21593) );
  XOR U22626 ( .A(a[922]), .B(n2307), .Z(n21597) );
  AND U22627 ( .A(a[924]), .B(b[0]), .Z(n21577) );
  XNOR U22628 ( .A(n21577), .B(n2175), .Z(n21579) );
  NANDN U22629 ( .A(b[0]), .B(a[923]), .Z(n21578) );
  NAND U22630 ( .A(n21579), .B(n21578), .Z(n21602) );
  AND U22631 ( .A(a[920]), .B(b[3]), .Z(n21601) );
  XOR U22632 ( .A(n21602), .B(n21601), .Z(n21604) );
  XOR U22633 ( .A(n21603), .B(n21604), .Z(n21592) );
  NANDN U22634 ( .A(n21581), .B(n21580), .Z(n21585) );
  OR U22635 ( .A(n21583), .B(n21582), .Z(n21584) );
  AND U22636 ( .A(n21585), .B(n21584), .Z(n21591) );
  XOR U22637 ( .A(n21592), .B(n21591), .Z(n21594) );
  XOR U22638 ( .A(n21593), .B(n21594), .Z(n21607) );
  XNOR U22639 ( .A(n21607), .B(sreg[1944]), .Z(n21609) );
  NANDN U22640 ( .A(n21586), .B(sreg[1943]), .Z(n21590) );
  NAND U22641 ( .A(n21588), .B(n21587), .Z(n21589) );
  NAND U22642 ( .A(n21590), .B(n21589), .Z(n21608) );
  XOR U22643 ( .A(n21609), .B(n21608), .Z(c[1944]) );
  NANDN U22644 ( .A(n21592), .B(n21591), .Z(n21596) );
  OR U22645 ( .A(n21594), .B(n21593), .Z(n21595) );
  AND U22646 ( .A(n21596), .B(n21595), .Z(n21614) );
  XOR U22647 ( .A(a[923]), .B(n2308), .Z(n21618) );
  AND U22648 ( .A(a[921]), .B(b[3]), .Z(n21622) );
  AND U22649 ( .A(a[925]), .B(b[0]), .Z(n21598) );
  XNOR U22650 ( .A(n21598), .B(n2175), .Z(n21600) );
  NANDN U22651 ( .A(b[0]), .B(a[924]), .Z(n21599) );
  NAND U22652 ( .A(n21600), .B(n21599), .Z(n21623) );
  XOR U22653 ( .A(n21622), .B(n21623), .Z(n21625) );
  XOR U22654 ( .A(n21624), .B(n21625), .Z(n21613) );
  NANDN U22655 ( .A(n21602), .B(n21601), .Z(n21606) );
  OR U22656 ( .A(n21604), .B(n21603), .Z(n21605) );
  AND U22657 ( .A(n21606), .B(n21605), .Z(n21612) );
  XOR U22658 ( .A(n21613), .B(n21612), .Z(n21615) );
  XOR U22659 ( .A(n21614), .B(n21615), .Z(n21628) );
  XNOR U22660 ( .A(n21628), .B(sreg[1945]), .Z(n21630) );
  NANDN U22661 ( .A(n21607), .B(sreg[1944]), .Z(n21611) );
  NAND U22662 ( .A(n21609), .B(n21608), .Z(n21610) );
  NAND U22663 ( .A(n21611), .B(n21610), .Z(n21629) );
  XOR U22664 ( .A(n21630), .B(n21629), .Z(c[1945]) );
  NANDN U22665 ( .A(n21613), .B(n21612), .Z(n21617) );
  OR U22666 ( .A(n21615), .B(n21614), .Z(n21616) );
  AND U22667 ( .A(n21617), .B(n21616), .Z(n21635) );
  XOR U22668 ( .A(a[924]), .B(n2308), .Z(n21639) );
  AND U22669 ( .A(a[926]), .B(b[0]), .Z(n21619) );
  XNOR U22670 ( .A(n21619), .B(n2175), .Z(n21621) );
  NANDN U22671 ( .A(b[0]), .B(a[925]), .Z(n21620) );
  NAND U22672 ( .A(n21621), .B(n21620), .Z(n21644) );
  AND U22673 ( .A(a[922]), .B(b[3]), .Z(n21643) );
  XOR U22674 ( .A(n21644), .B(n21643), .Z(n21646) );
  XOR U22675 ( .A(n21645), .B(n21646), .Z(n21634) );
  NANDN U22676 ( .A(n21623), .B(n21622), .Z(n21627) );
  OR U22677 ( .A(n21625), .B(n21624), .Z(n21626) );
  AND U22678 ( .A(n21627), .B(n21626), .Z(n21633) );
  XOR U22679 ( .A(n21634), .B(n21633), .Z(n21636) );
  XOR U22680 ( .A(n21635), .B(n21636), .Z(n21649) );
  XNOR U22681 ( .A(n21649), .B(sreg[1946]), .Z(n21651) );
  NANDN U22682 ( .A(n21628), .B(sreg[1945]), .Z(n21632) );
  NAND U22683 ( .A(n21630), .B(n21629), .Z(n21631) );
  NAND U22684 ( .A(n21632), .B(n21631), .Z(n21650) );
  XOR U22685 ( .A(n21651), .B(n21650), .Z(c[1946]) );
  NANDN U22686 ( .A(n21634), .B(n21633), .Z(n21638) );
  OR U22687 ( .A(n21636), .B(n21635), .Z(n21637) );
  AND U22688 ( .A(n21638), .B(n21637), .Z(n21656) );
  XOR U22689 ( .A(a[925]), .B(n2308), .Z(n21660) );
  AND U22690 ( .A(a[927]), .B(b[0]), .Z(n21640) );
  XNOR U22691 ( .A(n21640), .B(n2175), .Z(n21642) );
  NANDN U22692 ( .A(b[0]), .B(a[926]), .Z(n21641) );
  NAND U22693 ( .A(n21642), .B(n21641), .Z(n21665) );
  AND U22694 ( .A(a[923]), .B(b[3]), .Z(n21664) );
  XOR U22695 ( .A(n21665), .B(n21664), .Z(n21667) );
  XOR U22696 ( .A(n21666), .B(n21667), .Z(n21655) );
  NANDN U22697 ( .A(n21644), .B(n21643), .Z(n21648) );
  OR U22698 ( .A(n21646), .B(n21645), .Z(n21647) );
  AND U22699 ( .A(n21648), .B(n21647), .Z(n21654) );
  XOR U22700 ( .A(n21655), .B(n21654), .Z(n21657) );
  XOR U22701 ( .A(n21656), .B(n21657), .Z(n21670) );
  XNOR U22702 ( .A(n21670), .B(sreg[1947]), .Z(n21672) );
  NANDN U22703 ( .A(n21649), .B(sreg[1946]), .Z(n21653) );
  NAND U22704 ( .A(n21651), .B(n21650), .Z(n21652) );
  NAND U22705 ( .A(n21653), .B(n21652), .Z(n21671) );
  XOR U22706 ( .A(n21672), .B(n21671), .Z(c[1947]) );
  NANDN U22707 ( .A(n21655), .B(n21654), .Z(n21659) );
  OR U22708 ( .A(n21657), .B(n21656), .Z(n21658) );
  AND U22709 ( .A(n21659), .B(n21658), .Z(n21677) );
  XOR U22710 ( .A(a[926]), .B(n2308), .Z(n21681) );
  AND U22711 ( .A(a[928]), .B(b[0]), .Z(n21661) );
  XNOR U22712 ( .A(n21661), .B(n2175), .Z(n21663) );
  NANDN U22713 ( .A(b[0]), .B(a[927]), .Z(n21662) );
  NAND U22714 ( .A(n21663), .B(n21662), .Z(n21686) );
  AND U22715 ( .A(a[924]), .B(b[3]), .Z(n21685) );
  XOR U22716 ( .A(n21686), .B(n21685), .Z(n21688) );
  XOR U22717 ( .A(n21687), .B(n21688), .Z(n21676) );
  NANDN U22718 ( .A(n21665), .B(n21664), .Z(n21669) );
  OR U22719 ( .A(n21667), .B(n21666), .Z(n21668) );
  AND U22720 ( .A(n21669), .B(n21668), .Z(n21675) );
  XOR U22721 ( .A(n21676), .B(n21675), .Z(n21678) );
  XOR U22722 ( .A(n21677), .B(n21678), .Z(n21691) );
  XNOR U22723 ( .A(n21691), .B(sreg[1948]), .Z(n21693) );
  NANDN U22724 ( .A(n21670), .B(sreg[1947]), .Z(n21674) );
  NAND U22725 ( .A(n21672), .B(n21671), .Z(n21673) );
  NAND U22726 ( .A(n21674), .B(n21673), .Z(n21692) );
  XOR U22727 ( .A(n21693), .B(n21692), .Z(c[1948]) );
  NANDN U22728 ( .A(n21676), .B(n21675), .Z(n21680) );
  OR U22729 ( .A(n21678), .B(n21677), .Z(n21679) );
  AND U22730 ( .A(n21680), .B(n21679), .Z(n21698) );
  XOR U22731 ( .A(a[927]), .B(n2308), .Z(n21702) );
  AND U22732 ( .A(a[925]), .B(b[3]), .Z(n21706) );
  AND U22733 ( .A(a[929]), .B(b[0]), .Z(n21682) );
  XNOR U22734 ( .A(n21682), .B(n2175), .Z(n21684) );
  NANDN U22735 ( .A(b[0]), .B(a[928]), .Z(n21683) );
  NAND U22736 ( .A(n21684), .B(n21683), .Z(n21707) );
  XOR U22737 ( .A(n21706), .B(n21707), .Z(n21709) );
  XOR U22738 ( .A(n21708), .B(n21709), .Z(n21697) );
  NANDN U22739 ( .A(n21686), .B(n21685), .Z(n21690) );
  OR U22740 ( .A(n21688), .B(n21687), .Z(n21689) );
  AND U22741 ( .A(n21690), .B(n21689), .Z(n21696) );
  XOR U22742 ( .A(n21697), .B(n21696), .Z(n21699) );
  XOR U22743 ( .A(n21698), .B(n21699), .Z(n21712) );
  XNOR U22744 ( .A(n21712), .B(sreg[1949]), .Z(n21714) );
  NANDN U22745 ( .A(n21691), .B(sreg[1948]), .Z(n21695) );
  NAND U22746 ( .A(n21693), .B(n21692), .Z(n21694) );
  NAND U22747 ( .A(n21695), .B(n21694), .Z(n21713) );
  XOR U22748 ( .A(n21714), .B(n21713), .Z(c[1949]) );
  NANDN U22749 ( .A(n21697), .B(n21696), .Z(n21701) );
  OR U22750 ( .A(n21699), .B(n21698), .Z(n21700) );
  AND U22751 ( .A(n21701), .B(n21700), .Z(n21719) );
  XOR U22752 ( .A(a[928]), .B(n2308), .Z(n21723) );
  AND U22753 ( .A(a[930]), .B(b[0]), .Z(n21703) );
  XNOR U22754 ( .A(n21703), .B(n2175), .Z(n21705) );
  NANDN U22755 ( .A(b[0]), .B(a[929]), .Z(n21704) );
  NAND U22756 ( .A(n21705), .B(n21704), .Z(n21728) );
  AND U22757 ( .A(a[926]), .B(b[3]), .Z(n21727) );
  XOR U22758 ( .A(n21728), .B(n21727), .Z(n21730) );
  XOR U22759 ( .A(n21729), .B(n21730), .Z(n21718) );
  NANDN U22760 ( .A(n21707), .B(n21706), .Z(n21711) );
  OR U22761 ( .A(n21709), .B(n21708), .Z(n21710) );
  AND U22762 ( .A(n21711), .B(n21710), .Z(n21717) );
  XOR U22763 ( .A(n21718), .B(n21717), .Z(n21720) );
  XOR U22764 ( .A(n21719), .B(n21720), .Z(n21733) );
  XNOR U22765 ( .A(n21733), .B(sreg[1950]), .Z(n21735) );
  NANDN U22766 ( .A(n21712), .B(sreg[1949]), .Z(n21716) );
  NAND U22767 ( .A(n21714), .B(n21713), .Z(n21715) );
  NAND U22768 ( .A(n21716), .B(n21715), .Z(n21734) );
  XOR U22769 ( .A(n21735), .B(n21734), .Z(c[1950]) );
  NANDN U22770 ( .A(n21718), .B(n21717), .Z(n21722) );
  OR U22771 ( .A(n21720), .B(n21719), .Z(n21721) );
  AND U22772 ( .A(n21722), .B(n21721), .Z(n21740) );
  XOR U22773 ( .A(a[929]), .B(n2308), .Z(n21744) );
  AND U22774 ( .A(a[931]), .B(b[0]), .Z(n21724) );
  XNOR U22775 ( .A(n21724), .B(n2175), .Z(n21726) );
  NANDN U22776 ( .A(b[0]), .B(a[930]), .Z(n21725) );
  NAND U22777 ( .A(n21726), .B(n21725), .Z(n21749) );
  AND U22778 ( .A(a[927]), .B(b[3]), .Z(n21748) );
  XOR U22779 ( .A(n21749), .B(n21748), .Z(n21751) );
  XOR U22780 ( .A(n21750), .B(n21751), .Z(n21739) );
  NANDN U22781 ( .A(n21728), .B(n21727), .Z(n21732) );
  OR U22782 ( .A(n21730), .B(n21729), .Z(n21731) );
  AND U22783 ( .A(n21732), .B(n21731), .Z(n21738) );
  XOR U22784 ( .A(n21739), .B(n21738), .Z(n21741) );
  XOR U22785 ( .A(n21740), .B(n21741), .Z(n21754) );
  XNOR U22786 ( .A(n21754), .B(sreg[1951]), .Z(n21756) );
  NANDN U22787 ( .A(n21733), .B(sreg[1950]), .Z(n21737) );
  NAND U22788 ( .A(n21735), .B(n21734), .Z(n21736) );
  NAND U22789 ( .A(n21737), .B(n21736), .Z(n21755) );
  XOR U22790 ( .A(n21756), .B(n21755), .Z(c[1951]) );
  NANDN U22791 ( .A(n21739), .B(n21738), .Z(n21743) );
  OR U22792 ( .A(n21741), .B(n21740), .Z(n21742) );
  AND U22793 ( .A(n21743), .B(n21742), .Z(n21761) );
  XOR U22794 ( .A(a[930]), .B(n2309), .Z(n21765) );
  AND U22795 ( .A(a[928]), .B(b[3]), .Z(n21769) );
  AND U22796 ( .A(a[932]), .B(b[0]), .Z(n21745) );
  XNOR U22797 ( .A(n21745), .B(n2175), .Z(n21747) );
  NANDN U22798 ( .A(b[0]), .B(a[931]), .Z(n21746) );
  NAND U22799 ( .A(n21747), .B(n21746), .Z(n21770) );
  XOR U22800 ( .A(n21769), .B(n21770), .Z(n21772) );
  XOR U22801 ( .A(n21771), .B(n21772), .Z(n21760) );
  NANDN U22802 ( .A(n21749), .B(n21748), .Z(n21753) );
  OR U22803 ( .A(n21751), .B(n21750), .Z(n21752) );
  AND U22804 ( .A(n21753), .B(n21752), .Z(n21759) );
  XOR U22805 ( .A(n21760), .B(n21759), .Z(n21762) );
  XOR U22806 ( .A(n21761), .B(n21762), .Z(n21775) );
  XNOR U22807 ( .A(n21775), .B(sreg[1952]), .Z(n21777) );
  NANDN U22808 ( .A(n21754), .B(sreg[1951]), .Z(n21758) );
  NAND U22809 ( .A(n21756), .B(n21755), .Z(n21757) );
  NAND U22810 ( .A(n21758), .B(n21757), .Z(n21776) );
  XOR U22811 ( .A(n21777), .B(n21776), .Z(c[1952]) );
  NANDN U22812 ( .A(n21760), .B(n21759), .Z(n21764) );
  OR U22813 ( .A(n21762), .B(n21761), .Z(n21763) );
  AND U22814 ( .A(n21764), .B(n21763), .Z(n21782) );
  XOR U22815 ( .A(a[931]), .B(n2309), .Z(n21786) );
  AND U22816 ( .A(a[933]), .B(b[0]), .Z(n21766) );
  XNOR U22817 ( .A(n21766), .B(n2175), .Z(n21768) );
  NANDN U22818 ( .A(b[0]), .B(a[932]), .Z(n21767) );
  NAND U22819 ( .A(n21768), .B(n21767), .Z(n21791) );
  AND U22820 ( .A(a[929]), .B(b[3]), .Z(n21790) );
  XOR U22821 ( .A(n21791), .B(n21790), .Z(n21793) );
  XOR U22822 ( .A(n21792), .B(n21793), .Z(n21781) );
  NANDN U22823 ( .A(n21770), .B(n21769), .Z(n21774) );
  OR U22824 ( .A(n21772), .B(n21771), .Z(n21773) );
  AND U22825 ( .A(n21774), .B(n21773), .Z(n21780) );
  XOR U22826 ( .A(n21781), .B(n21780), .Z(n21783) );
  XOR U22827 ( .A(n21782), .B(n21783), .Z(n21796) );
  XNOR U22828 ( .A(n21796), .B(sreg[1953]), .Z(n21798) );
  NANDN U22829 ( .A(n21775), .B(sreg[1952]), .Z(n21779) );
  NAND U22830 ( .A(n21777), .B(n21776), .Z(n21778) );
  NAND U22831 ( .A(n21779), .B(n21778), .Z(n21797) );
  XOR U22832 ( .A(n21798), .B(n21797), .Z(c[1953]) );
  NANDN U22833 ( .A(n21781), .B(n21780), .Z(n21785) );
  OR U22834 ( .A(n21783), .B(n21782), .Z(n21784) );
  AND U22835 ( .A(n21785), .B(n21784), .Z(n21803) );
  XOR U22836 ( .A(a[932]), .B(n2309), .Z(n21807) );
  AND U22837 ( .A(a[930]), .B(b[3]), .Z(n21811) );
  AND U22838 ( .A(a[934]), .B(b[0]), .Z(n21787) );
  XNOR U22839 ( .A(n21787), .B(n2175), .Z(n21789) );
  NANDN U22840 ( .A(b[0]), .B(a[933]), .Z(n21788) );
  NAND U22841 ( .A(n21789), .B(n21788), .Z(n21812) );
  XOR U22842 ( .A(n21811), .B(n21812), .Z(n21814) );
  XOR U22843 ( .A(n21813), .B(n21814), .Z(n21802) );
  NANDN U22844 ( .A(n21791), .B(n21790), .Z(n21795) );
  OR U22845 ( .A(n21793), .B(n21792), .Z(n21794) );
  AND U22846 ( .A(n21795), .B(n21794), .Z(n21801) );
  XOR U22847 ( .A(n21802), .B(n21801), .Z(n21804) );
  XOR U22848 ( .A(n21803), .B(n21804), .Z(n21817) );
  XNOR U22849 ( .A(n21817), .B(sreg[1954]), .Z(n21819) );
  NANDN U22850 ( .A(n21796), .B(sreg[1953]), .Z(n21800) );
  NAND U22851 ( .A(n21798), .B(n21797), .Z(n21799) );
  NAND U22852 ( .A(n21800), .B(n21799), .Z(n21818) );
  XOR U22853 ( .A(n21819), .B(n21818), .Z(c[1954]) );
  NANDN U22854 ( .A(n21802), .B(n21801), .Z(n21806) );
  OR U22855 ( .A(n21804), .B(n21803), .Z(n21805) );
  AND U22856 ( .A(n21806), .B(n21805), .Z(n21824) );
  XOR U22857 ( .A(a[933]), .B(n2309), .Z(n21828) );
  AND U22858 ( .A(a[935]), .B(b[0]), .Z(n21808) );
  XNOR U22859 ( .A(n21808), .B(n2175), .Z(n21810) );
  NANDN U22860 ( .A(b[0]), .B(a[934]), .Z(n21809) );
  NAND U22861 ( .A(n21810), .B(n21809), .Z(n21833) );
  AND U22862 ( .A(a[931]), .B(b[3]), .Z(n21832) );
  XOR U22863 ( .A(n21833), .B(n21832), .Z(n21835) );
  XOR U22864 ( .A(n21834), .B(n21835), .Z(n21823) );
  NANDN U22865 ( .A(n21812), .B(n21811), .Z(n21816) );
  OR U22866 ( .A(n21814), .B(n21813), .Z(n21815) );
  AND U22867 ( .A(n21816), .B(n21815), .Z(n21822) );
  XOR U22868 ( .A(n21823), .B(n21822), .Z(n21825) );
  XOR U22869 ( .A(n21824), .B(n21825), .Z(n21838) );
  XNOR U22870 ( .A(n21838), .B(sreg[1955]), .Z(n21840) );
  NANDN U22871 ( .A(n21817), .B(sreg[1954]), .Z(n21821) );
  NAND U22872 ( .A(n21819), .B(n21818), .Z(n21820) );
  NAND U22873 ( .A(n21821), .B(n21820), .Z(n21839) );
  XOR U22874 ( .A(n21840), .B(n21839), .Z(c[1955]) );
  NANDN U22875 ( .A(n21823), .B(n21822), .Z(n21827) );
  OR U22876 ( .A(n21825), .B(n21824), .Z(n21826) );
  AND U22877 ( .A(n21827), .B(n21826), .Z(n21845) );
  XOR U22878 ( .A(a[934]), .B(n2309), .Z(n21849) );
  AND U22879 ( .A(a[936]), .B(b[0]), .Z(n21829) );
  XNOR U22880 ( .A(n21829), .B(n2175), .Z(n21831) );
  NANDN U22881 ( .A(b[0]), .B(a[935]), .Z(n21830) );
  NAND U22882 ( .A(n21831), .B(n21830), .Z(n21854) );
  AND U22883 ( .A(a[932]), .B(b[3]), .Z(n21853) );
  XOR U22884 ( .A(n21854), .B(n21853), .Z(n21856) );
  XOR U22885 ( .A(n21855), .B(n21856), .Z(n21844) );
  NANDN U22886 ( .A(n21833), .B(n21832), .Z(n21837) );
  OR U22887 ( .A(n21835), .B(n21834), .Z(n21836) );
  AND U22888 ( .A(n21837), .B(n21836), .Z(n21843) );
  XOR U22889 ( .A(n21844), .B(n21843), .Z(n21846) );
  XOR U22890 ( .A(n21845), .B(n21846), .Z(n21859) );
  XNOR U22891 ( .A(n21859), .B(sreg[1956]), .Z(n21861) );
  NANDN U22892 ( .A(n21838), .B(sreg[1955]), .Z(n21842) );
  NAND U22893 ( .A(n21840), .B(n21839), .Z(n21841) );
  NAND U22894 ( .A(n21842), .B(n21841), .Z(n21860) );
  XOR U22895 ( .A(n21861), .B(n21860), .Z(c[1956]) );
  NANDN U22896 ( .A(n21844), .B(n21843), .Z(n21848) );
  OR U22897 ( .A(n21846), .B(n21845), .Z(n21847) );
  AND U22898 ( .A(n21848), .B(n21847), .Z(n21866) );
  XOR U22899 ( .A(a[935]), .B(n2309), .Z(n21870) );
  AND U22900 ( .A(a[937]), .B(b[0]), .Z(n21850) );
  XNOR U22901 ( .A(n21850), .B(n2175), .Z(n21852) );
  NANDN U22902 ( .A(b[0]), .B(a[936]), .Z(n21851) );
  NAND U22903 ( .A(n21852), .B(n21851), .Z(n21875) );
  AND U22904 ( .A(a[933]), .B(b[3]), .Z(n21874) );
  XOR U22905 ( .A(n21875), .B(n21874), .Z(n21877) );
  XOR U22906 ( .A(n21876), .B(n21877), .Z(n21865) );
  NANDN U22907 ( .A(n21854), .B(n21853), .Z(n21858) );
  OR U22908 ( .A(n21856), .B(n21855), .Z(n21857) );
  AND U22909 ( .A(n21858), .B(n21857), .Z(n21864) );
  XOR U22910 ( .A(n21865), .B(n21864), .Z(n21867) );
  XOR U22911 ( .A(n21866), .B(n21867), .Z(n21880) );
  XNOR U22912 ( .A(n21880), .B(sreg[1957]), .Z(n21882) );
  NANDN U22913 ( .A(n21859), .B(sreg[1956]), .Z(n21863) );
  NAND U22914 ( .A(n21861), .B(n21860), .Z(n21862) );
  NAND U22915 ( .A(n21863), .B(n21862), .Z(n21881) );
  XOR U22916 ( .A(n21882), .B(n21881), .Z(c[1957]) );
  NANDN U22917 ( .A(n21865), .B(n21864), .Z(n21869) );
  OR U22918 ( .A(n21867), .B(n21866), .Z(n21868) );
  AND U22919 ( .A(n21869), .B(n21868), .Z(n21887) );
  XOR U22920 ( .A(a[936]), .B(n2309), .Z(n21891) );
  AND U22921 ( .A(a[934]), .B(b[3]), .Z(n21895) );
  AND U22922 ( .A(a[938]), .B(b[0]), .Z(n21871) );
  XNOR U22923 ( .A(n21871), .B(n2175), .Z(n21873) );
  NANDN U22924 ( .A(b[0]), .B(a[937]), .Z(n21872) );
  NAND U22925 ( .A(n21873), .B(n21872), .Z(n21896) );
  XOR U22926 ( .A(n21895), .B(n21896), .Z(n21898) );
  XOR U22927 ( .A(n21897), .B(n21898), .Z(n21886) );
  NANDN U22928 ( .A(n21875), .B(n21874), .Z(n21879) );
  OR U22929 ( .A(n21877), .B(n21876), .Z(n21878) );
  AND U22930 ( .A(n21879), .B(n21878), .Z(n21885) );
  XOR U22931 ( .A(n21886), .B(n21885), .Z(n21888) );
  XOR U22932 ( .A(n21887), .B(n21888), .Z(n21901) );
  XNOR U22933 ( .A(n21901), .B(sreg[1958]), .Z(n21903) );
  NANDN U22934 ( .A(n21880), .B(sreg[1957]), .Z(n21884) );
  NAND U22935 ( .A(n21882), .B(n21881), .Z(n21883) );
  NAND U22936 ( .A(n21884), .B(n21883), .Z(n21902) );
  XOR U22937 ( .A(n21903), .B(n21902), .Z(c[1958]) );
  NANDN U22938 ( .A(n21886), .B(n21885), .Z(n21890) );
  OR U22939 ( .A(n21888), .B(n21887), .Z(n21889) );
  AND U22940 ( .A(n21890), .B(n21889), .Z(n21908) );
  XOR U22941 ( .A(a[937]), .B(n2310), .Z(n21912) );
  AND U22942 ( .A(a[939]), .B(b[0]), .Z(n21892) );
  XNOR U22943 ( .A(n21892), .B(n2175), .Z(n21894) );
  NANDN U22944 ( .A(b[0]), .B(a[938]), .Z(n21893) );
  NAND U22945 ( .A(n21894), .B(n21893), .Z(n21917) );
  AND U22946 ( .A(a[935]), .B(b[3]), .Z(n21916) );
  XOR U22947 ( .A(n21917), .B(n21916), .Z(n21919) );
  XOR U22948 ( .A(n21918), .B(n21919), .Z(n21907) );
  NANDN U22949 ( .A(n21896), .B(n21895), .Z(n21900) );
  OR U22950 ( .A(n21898), .B(n21897), .Z(n21899) );
  AND U22951 ( .A(n21900), .B(n21899), .Z(n21906) );
  XOR U22952 ( .A(n21907), .B(n21906), .Z(n21909) );
  XOR U22953 ( .A(n21908), .B(n21909), .Z(n21922) );
  XNOR U22954 ( .A(n21922), .B(sreg[1959]), .Z(n21924) );
  NANDN U22955 ( .A(n21901), .B(sreg[1958]), .Z(n21905) );
  NAND U22956 ( .A(n21903), .B(n21902), .Z(n21904) );
  NAND U22957 ( .A(n21905), .B(n21904), .Z(n21923) );
  XOR U22958 ( .A(n21924), .B(n21923), .Z(c[1959]) );
  NANDN U22959 ( .A(n21907), .B(n21906), .Z(n21911) );
  OR U22960 ( .A(n21909), .B(n21908), .Z(n21910) );
  AND U22961 ( .A(n21911), .B(n21910), .Z(n21929) );
  XOR U22962 ( .A(a[938]), .B(n2310), .Z(n21933) );
  AND U22963 ( .A(a[940]), .B(b[0]), .Z(n21913) );
  XNOR U22964 ( .A(n21913), .B(n2175), .Z(n21915) );
  NANDN U22965 ( .A(b[0]), .B(a[939]), .Z(n21914) );
  NAND U22966 ( .A(n21915), .B(n21914), .Z(n21938) );
  AND U22967 ( .A(a[936]), .B(b[3]), .Z(n21937) );
  XOR U22968 ( .A(n21938), .B(n21937), .Z(n21940) );
  XOR U22969 ( .A(n21939), .B(n21940), .Z(n21928) );
  NANDN U22970 ( .A(n21917), .B(n21916), .Z(n21921) );
  OR U22971 ( .A(n21919), .B(n21918), .Z(n21920) );
  AND U22972 ( .A(n21921), .B(n21920), .Z(n21927) );
  XOR U22973 ( .A(n21928), .B(n21927), .Z(n21930) );
  XOR U22974 ( .A(n21929), .B(n21930), .Z(n21943) );
  XNOR U22975 ( .A(n21943), .B(sreg[1960]), .Z(n21945) );
  NANDN U22976 ( .A(n21922), .B(sreg[1959]), .Z(n21926) );
  NAND U22977 ( .A(n21924), .B(n21923), .Z(n21925) );
  NAND U22978 ( .A(n21926), .B(n21925), .Z(n21944) );
  XOR U22979 ( .A(n21945), .B(n21944), .Z(c[1960]) );
  NANDN U22980 ( .A(n21928), .B(n21927), .Z(n21932) );
  OR U22981 ( .A(n21930), .B(n21929), .Z(n21931) );
  AND U22982 ( .A(n21932), .B(n21931), .Z(n21950) );
  XOR U22983 ( .A(a[939]), .B(n2310), .Z(n21954) );
  AND U22984 ( .A(a[941]), .B(b[0]), .Z(n21934) );
  XNOR U22985 ( .A(n21934), .B(n2175), .Z(n21936) );
  NANDN U22986 ( .A(b[0]), .B(a[940]), .Z(n21935) );
  NAND U22987 ( .A(n21936), .B(n21935), .Z(n21959) );
  AND U22988 ( .A(a[937]), .B(b[3]), .Z(n21958) );
  XOR U22989 ( .A(n21959), .B(n21958), .Z(n21961) );
  XOR U22990 ( .A(n21960), .B(n21961), .Z(n21949) );
  NANDN U22991 ( .A(n21938), .B(n21937), .Z(n21942) );
  OR U22992 ( .A(n21940), .B(n21939), .Z(n21941) );
  AND U22993 ( .A(n21942), .B(n21941), .Z(n21948) );
  XOR U22994 ( .A(n21949), .B(n21948), .Z(n21951) );
  XOR U22995 ( .A(n21950), .B(n21951), .Z(n21964) );
  XNOR U22996 ( .A(n21964), .B(sreg[1961]), .Z(n21966) );
  NANDN U22997 ( .A(n21943), .B(sreg[1960]), .Z(n21947) );
  NAND U22998 ( .A(n21945), .B(n21944), .Z(n21946) );
  NAND U22999 ( .A(n21947), .B(n21946), .Z(n21965) );
  XOR U23000 ( .A(n21966), .B(n21965), .Z(c[1961]) );
  NANDN U23001 ( .A(n21949), .B(n21948), .Z(n21953) );
  OR U23002 ( .A(n21951), .B(n21950), .Z(n21952) );
  AND U23003 ( .A(n21953), .B(n21952), .Z(n21971) );
  XOR U23004 ( .A(a[940]), .B(n2310), .Z(n21975) );
  AND U23005 ( .A(a[942]), .B(b[0]), .Z(n21955) );
  XNOR U23006 ( .A(n21955), .B(n2175), .Z(n21957) );
  NANDN U23007 ( .A(b[0]), .B(a[941]), .Z(n21956) );
  NAND U23008 ( .A(n21957), .B(n21956), .Z(n21980) );
  AND U23009 ( .A(a[938]), .B(b[3]), .Z(n21979) );
  XOR U23010 ( .A(n21980), .B(n21979), .Z(n21982) );
  XOR U23011 ( .A(n21981), .B(n21982), .Z(n21970) );
  NANDN U23012 ( .A(n21959), .B(n21958), .Z(n21963) );
  OR U23013 ( .A(n21961), .B(n21960), .Z(n21962) );
  AND U23014 ( .A(n21963), .B(n21962), .Z(n21969) );
  XOR U23015 ( .A(n21970), .B(n21969), .Z(n21972) );
  XOR U23016 ( .A(n21971), .B(n21972), .Z(n21985) );
  XNOR U23017 ( .A(n21985), .B(sreg[1962]), .Z(n21987) );
  NANDN U23018 ( .A(n21964), .B(sreg[1961]), .Z(n21968) );
  NAND U23019 ( .A(n21966), .B(n21965), .Z(n21967) );
  NAND U23020 ( .A(n21968), .B(n21967), .Z(n21986) );
  XOR U23021 ( .A(n21987), .B(n21986), .Z(c[1962]) );
  NANDN U23022 ( .A(n21970), .B(n21969), .Z(n21974) );
  OR U23023 ( .A(n21972), .B(n21971), .Z(n21973) );
  AND U23024 ( .A(n21974), .B(n21973), .Z(n21992) );
  XOR U23025 ( .A(a[941]), .B(n2310), .Z(n21996) );
  AND U23026 ( .A(a[939]), .B(b[3]), .Z(n22000) );
  AND U23027 ( .A(a[943]), .B(b[0]), .Z(n21976) );
  XNOR U23028 ( .A(n21976), .B(n2175), .Z(n21978) );
  NANDN U23029 ( .A(b[0]), .B(a[942]), .Z(n21977) );
  NAND U23030 ( .A(n21978), .B(n21977), .Z(n22001) );
  XOR U23031 ( .A(n22000), .B(n22001), .Z(n22003) );
  XOR U23032 ( .A(n22002), .B(n22003), .Z(n21991) );
  NANDN U23033 ( .A(n21980), .B(n21979), .Z(n21984) );
  OR U23034 ( .A(n21982), .B(n21981), .Z(n21983) );
  AND U23035 ( .A(n21984), .B(n21983), .Z(n21990) );
  XOR U23036 ( .A(n21991), .B(n21990), .Z(n21993) );
  XOR U23037 ( .A(n21992), .B(n21993), .Z(n22006) );
  XNOR U23038 ( .A(n22006), .B(sreg[1963]), .Z(n22008) );
  NANDN U23039 ( .A(n21985), .B(sreg[1962]), .Z(n21989) );
  NAND U23040 ( .A(n21987), .B(n21986), .Z(n21988) );
  NAND U23041 ( .A(n21989), .B(n21988), .Z(n22007) );
  XOR U23042 ( .A(n22008), .B(n22007), .Z(c[1963]) );
  NANDN U23043 ( .A(n21991), .B(n21990), .Z(n21995) );
  OR U23044 ( .A(n21993), .B(n21992), .Z(n21994) );
  AND U23045 ( .A(n21995), .B(n21994), .Z(n22013) );
  XOR U23046 ( .A(a[942]), .B(n2310), .Z(n22017) );
  AND U23047 ( .A(a[944]), .B(b[0]), .Z(n21997) );
  XNOR U23048 ( .A(n21997), .B(n2175), .Z(n21999) );
  NANDN U23049 ( .A(b[0]), .B(a[943]), .Z(n21998) );
  NAND U23050 ( .A(n21999), .B(n21998), .Z(n22022) );
  AND U23051 ( .A(a[940]), .B(b[3]), .Z(n22021) );
  XOR U23052 ( .A(n22022), .B(n22021), .Z(n22024) );
  XOR U23053 ( .A(n22023), .B(n22024), .Z(n22012) );
  NANDN U23054 ( .A(n22001), .B(n22000), .Z(n22005) );
  OR U23055 ( .A(n22003), .B(n22002), .Z(n22004) );
  AND U23056 ( .A(n22005), .B(n22004), .Z(n22011) );
  XOR U23057 ( .A(n22012), .B(n22011), .Z(n22014) );
  XOR U23058 ( .A(n22013), .B(n22014), .Z(n22027) );
  XNOR U23059 ( .A(n22027), .B(sreg[1964]), .Z(n22029) );
  NANDN U23060 ( .A(n22006), .B(sreg[1963]), .Z(n22010) );
  NAND U23061 ( .A(n22008), .B(n22007), .Z(n22009) );
  NAND U23062 ( .A(n22010), .B(n22009), .Z(n22028) );
  XOR U23063 ( .A(n22029), .B(n22028), .Z(c[1964]) );
  NANDN U23064 ( .A(n22012), .B(n22011), .Z(n22016) );
  OR U23065 ( .A(n22014), .B(n22013), .Z(n22015) );
  AND U23066 ( .A(n22016), .B(n22015), .Z(n22034) );
  XOR U23067 ( .A(a[943]), .B(n2310), .Z(n22038) );
  AND U23068 ( .A(a[945]), .B(b[0]), .Z(n22018) );
  XNOR U23069 ( .A(n22018), .B(n2175), .Z(n22020) );
  NANDN U23070 ( .A(b[0]), .B(a[944]), .Z(n22019) );
  NAND U23071 ( .A(n22020), .B(n22019), .Z(n22043) );
  AND U23072 ( .A(a[941]), .B(b[3]), .Z(n22042) );
  XOR U23073 ( .A(n22043), .B(n22042), .Z(n22045) );
  XOR U23074 ( .A(n22044), .B(n22045), .Z(n22033) );
  NANDN U23075 ( .A(n22022), .B(n22021), .Z(n22026) );
  OR U23076 ( .A(n22024), .B(n22023), .Z(n22025) );
  AND U23077 ( .A(n22026), .B(n22025), .Z(n22032) );
  XOR U23078 ( .A(n22033), .B(n22032), .Z(n22035) );
  XOR U23079 ( .A(n22034), .B(n22035), .Z(n22048) );
  XNOR U23080 ( .A(n22048), .B(sreg[1965]), .Z(n22050) );
  NANDN U23081 ( .A(n22027), .B(sreg[1964]), .Z(n22031) );
  NAND U23082 ( .A(n22029), .B(n22028), .Z(n22030) );
  NAND U23083 ( .A(n22031), .B(n22030), .Z(n22049) );
  XOR U23084 ( .A(n22050), .B(n22049), .Z(c[1965]) );
  NANDN U23085 ( .A(n22033), .B(n22032), .Z(n22037) );
  OR U23086 ( .A(n22035), .B(n22034), .Z(n22036) );
  AND U23087 ( .A(n22037), .B(n22036), .Z(n22055) );
  XOR U23088 ( .A(a[944]), .B(n2311), .Z(n22059) );
  AND U23089 ( .A(a[946]), .B(b[0]), .Z(n22039) );
  XNOR U23090 ( .A(n22039), .B(n2175), .Z(n22041) );
  NANDN U23091 ( .A(b[0]), .B(a[945]), .Z(n22040) );
  NAND U23092 ( .A(n22041), .B(n22040), .Z(n22064) );
  AND U23093 ( .A(a[942]), .B(b[3]), .Z(n22063) );
  XOR U23094 ( .A(n22064), .B(n22063), .Z(n22066) );
  XOR U23095 ( .A(n22065), .B(n22066), .Z(n22054) );
  NANDN U23096 ( .A(n22043), .B(n22042), .Z(n22047) );
  OR U23097 ( .A(n22045), .B(n22044), .Z(n22046) );
  AND U23098 ( .A(n22047), .B(n22046), .Z(n22053) );
  XOR U23099 ( .A(n22054), .B(n22053), .Z(n22056) );
  XOR U23100 ( .A(n22055), .B(n22056), .Z(n22069) );
  XNOR U23101 ( .A(n22069), .B(sreg[1966]), .Z(n22071) );
  NANDN U23102 ( .A(n22048), .B(sreg[1965]), .Z(n22052) );
  NAND U23103 ( .A(n22050), .B(n22049), .Z(n22051) );
  NAND U23104 ( .A(n22052), .B(n22051), .Z(n22070) );
  XOR U23105 ( .A(n22071), .B(n22070), .Z(c[1966]) );
  NANDN U23106 ( .A(n22054), .B(n22053), .Z(n22058) );
  OR U23107 ( .A(n22056), .B(n22055), .Z(n22057) );
  AND U23108 ( .A(n22058), .B(n22057), .Z(n22076) );
  XOR U23109 ( .A(a[945]), .B(n2311), .Z(n22080) );
  AND U23110 ( .A(a[947]), .B(b[0]), .Z(n22060) );
  XNOR U23111 ( .A(n22060), .B(n2175), .Z(n22062) );
  NANDN U23112 ( .A(b[0]), .B(a[946]), .Z(n22061) );
  NAND U23113 ( .A(n22062), .B(n22061), .Z(n22085) );
  AND U23114 ( .A(a[943]), .B(b[3]), .Z(n22084) );
  XOR U23115 ( .A(n22085), .B(n22084), .Z(n22087) );
  XOR U23116 ( .A(n22086), .B(n22087), .Z(n22075) );
  NANDN U23117 ( .A(n22064), .B(n22063), .Z(n22068) );
  OR U23118 ( .A(n22066), .B(n22065), .Z(n22067) );
  AND U23119 ( .A(n22068), .B(n22067), .Z(n22074) );
  XOR U23120 ( .A(n22075), .B(n22074), .Z(n22077) );
  XOR U23121 ( .A(n22076), .B(n22077), .Z(n22090) );
  XNOR U23122 ( .A(n22090), .B(sreg[1967]), .Z(n22092) );
  NANDN U23123 ( .A(n22069), .B(sreg[1966]), .Z(n22073) );
  NAND U23124 ( .A(n22071), .B(n22070), .Z(n22072) );
  NAND U23125 ( .A(n22073), .B(n22072), .Z(n22091) );
  XOR U23126 ( .A(n22092), .B(n22091), .Z(c[1967]) );
  NANDN U23127 ( .A(n22075), .B(n22074), .Z(n22079) );
  OR U23128 ( .A(n22077), .B(n22076), .Z(n22078) );
  AND U23129 ( .A(n22079), .B(n22078), .Z(n22097) );
  XOR U23130 ( .A(a[946]), .B(n2311), .Z(n22101) );
  AND U23131 ( .A(a[948]), .B(b[0]), .Z(n22081) );
  XNOR U23132 ( .A(n22081), .B(n2175), .Z(n22083) );
  NANDN U23133 ( .A(b[0]), .B(a[947]), .Z(n22082) );
  NAND U23134 ( .A(n22083), .B(n22082), .Z(n22106) );
  AND U23135 ( .A(a[944]), .B(b[3]), .Z(n22105) );
  XOR U23136 ( .A(n22106), .B(n22105), .Z(n22108) );
  XOR U23137 ( .A(n22107), .B(n22108), .Z(n22096) );
  NANDN U23138 ( .A(n22085), .B(n22084), .Z(n22089) );
  OR U23139 ( .A(n22087), .B(n22086), .Z(n22088) );
  AND U23140 ( .A(n22089), .B(n22088), .Z(n22095) );
  XOR U23141 ( .A(n22096), .B(n22095), .Z(n22098) );
  XOR U23142 ( .A(n22097), .B(n22098), .Z(n22111) );
  XNOR U23143 ( .A(n22111), .B(sreg[1968]), .Z(n22113) );
  NANDN U23144 ( .A(n22090), .B(sreg[1967]), .Z(n22094) );
  NAND U23145 ( .A(n22092), .B(n22091), .Z(n22093) );
  NAND U23146 ( .A(n22094), .B(n22093), .Z(n22112) );
  XOR U23147 ( .A(n22113), .B(n22112), .Z(c[1968]) );
  NANDN U23148 ( .A(n22096), .B(n22095), .Z(n22100) );
  OR U23149 ( .A(n22098), .B(n22097), .Z(n22099) );
  AND U23150 ( .A(n22100), .B(n22099), .Z(n22118) );
  XOR U23151 ( .A(a[947]), .B(n2311), .Z(n22122) );
  AND U23152 ( .A(a[949]), .B(b[0]), .Z(n22102) );
  XNOR U23153 ( .A(n22102), .B(n2175), .Z(n22104) );
  NANDN U23154 ( .A(b[0]), .B(a[948]), .Z(n22103) );
  NAND U23155 ( .A(n22104), .B(n22103), .Z(n22127) );
  AND U23156 ( .A(a[945]), .B(b[3]), .Z(n22126) );
  XOR U23157 ( .A(n22127), .B(n22126), .Z(n22129) );
  XOR U23158 ( .A(n22128), .B(n22129), .Z(n22117) );
  NANDN U23159 ( .A(n22106), .B(n22105), .Z(n22110) );
  OR U23160 ( .A(n22108), .B(n22107), .Z(n22109) );
  AND U23161 ( .A(n22110), .B(n22109), .Z(n22116) );
  XOR U23162 ( .A(n22117), .B(n22116), .Z(n22119) );
  XOR U23163 ( .A(n22118), .B(n22119), .Z(n22132) );
  XNOR U23164 ( .A(n22132), .B(sreg[1969]), .Z(n22134) );
  NANDN U23165 ( .A(n22111), .B(sreg[1968]), .Z(n22115) );
  NAND U23166 ( .A(n22113), .B(n22112), .Z(n22114) );
  NAND U23167 ( .A(n22115), .B(n22114), .Z(n22133) );
  XOR U23168 ( .A(n22134), .B(n22133), .Z(c[1969]) );
  NANDN U23169 ( .A(n22117), .B(n22116), .Z(n22121) );
  OR U23170 ( .A(n22119), .B(n22118), .Z(n22120) );
  AND U23171 ( .A(n22121), .B(n22120), .Z(n22139) );
  XOR U23172 ( .A(a[948]), .B(n2311), .Z(n22143) );
  AND U23173 ( .A(a[950]), .B(b[0]), .Z(n22123) );
  XNOR U23174 ( .A(n22123), .B(n2175), .Z(n22125) );
  NANDN U23175 ( .A(b[0]), .B(a[949]), .Z(n22124) );
  NAND U23176 ( .A(n22125), .B(n22124), .Z(n22148) );
  AND U23177 ( .A(a[946]), .B(b[3]), .Z(n22147) );
  XOR U23178 ( .A(n22148), .B(n22147), .Z(n22150) );
  XOR U23179 ( .A(n22149), .B(n22150), .Z(n22138) );
  NANDN U23180 ( .A(n22127), .B(n22126), .Z(n22131) );
  OR U23181 ( .A(n22129), .B(n22128), .Z(n22130) );
  AND U23182 ( .A(n22131), .B(n22130), .Z(n22137) );
  XOR U23183 ( .A(n22138), .B(n22137), .Z(n22140) );
  XOR U23184 ( .A(n22139), .B(n22140), .Z(n22153) );
  XNOR U23185 ( .A(n22153), .B(sreg[1970]), .Z(n22155) );
  NANDN U23186 ( .A(n22132), .B(sreg[1969]), .Z(n22136) );
  NAND U23187 ( .A(n22134), .B(n22133), .Z(n22135) );
  NAND U23188 ( .A(n22136), .B(n22135), .Z(n22154) );
  XOR U23189 ( .A(n22155), .B(n22154), .Z(c[1970]) );
  NANDN U23190 ( .A(n22138), .B(n22137), .Z(n22142) );
  OR U23191 ( .A(n22140), .B(n22139), .Z(n22141) );
  AND U23192 ( .A(n22142), .B(n22141), .Z(n22160) );
  XOR U23193 ( .A(a[949]), .B(n2311), .Z(n22164) );
  AND U23194 ( .A(a[951]), .B(b[0]), .Z(n22144) );
  XNOR U23195 ( .A(n22144), .B(n2175), .Z(n22146) );
  NANDN U23196 ( .A(b[0]), .B(a[950]), .Z(n22145) );
  NAND U23197 ( .A(n22146), .B(n22145), .Z(n22169) );
  AND U23198 ( .A(a[947]), .B(b[3]), .Z(n22168) );
  XOR U23199 ( .A(n22169), .B(n22168), .Z(n22171) );
  XOR U23200 ( .A(n22170), .B(n22171), .Z(n22159) );
  NANDN U23201 ( .A(n22148), .B(n22147), .Z(n22152) );
  OR U23202 ( .A(n22150), .B(n22149), .Z(n22151) );
  AND U23203 ( .A(n22152), .B(n22151), .Z(n22158) );
  XOR U23204 ( .A(n22159), .B(n22158), .Z(n22161) );
  XOR U23205 ( .A(n22160), .B(n22161), .Z(n22174) );
  XNOR U23206 ( .A(n22174), .B(sreg[1971]), .Z(n22176) );
  NANDN U23207 ( .A(n22153), .B(sreg[1970]), .Z(n22157) );
  NAND U23208 ( .A(n22155), .B(n22154), .Z(n22156) );
  NAND U23209 ( .A(n22157), .B(n22156), .Z(n22175) );
  XOR U23210 ( .A(n22176), .B(n22175), .Z(c[1971]) );
  NANDN U23211 ( .A(n22159), .B(n22158), .Z(n22163) );
  OR U23212 ( .A(n22161), .B(n22160), .Z(n22162) );
  AND U23213 ( .A(n22163), .B(n22162), .Z(n22181) );
  XOR U23214 ( .A(a[950]), .B(n2311), .Z(n22185) );
  AND U23215 ( .A(a[952]), .B(b[0]), .Z(n22165) );
  XNOR U23216 ( .A(n22165), .B(n2175), .Z(n22167) );
  NANDN U23217 ( .A(b[0]), .B(a[951]), .Z(n22166) );
  NAND U23218 ( .A(n22167), .B(n22166), .Z(n22190) );
  AND U23219 ( .A(a[948]), .B(b[3]), .Z(n22189) );
  XOR U23220 ( .A(n22190), .B(n22189), .Z(n22192) );
  XOR U23221 ( .A(n22191), .B(n22192), .Z(n22180) );
  NANDN U23222 ( .A(n22169), .B(n22168), .Z(n22173) );
  OR U23223 ( .A(n22171), .B(n22170), .Z(n22172) );
  AND U23224 ( .A(n22173), .B(n22172), .Z(n22179) );
  XOR U23225 ( .A(n22180), .B(n22179), .Z(n22182) );
  XOR U23226 ( .A(n22181), .B(n22182), .Z(n22195) );
  XNOR U23227 ( .A(n22195), .B(sreg[1972]), .Z(n22197) );
  NANDN U23228 ( .A(n22174), .B(sreg[1971]), .Z(n22178) );
  NAND U23229 ( .A(n22176), .B(n22175), .Z(n22177) );
  NAND U23230 ( .A(n22178), .B(n22177), .Z(n22196) );
  XOR U23231 ( .A(n22197), .B(n22196), .Z(c[1972]) );
  NANDN U23232 ( .A(n22180), .B(n22179), .Z(n22184) );
  OR U23233 ( .A(n22182), .B(n22181), .Z(n22183) );
  AND U23234 ( .A(n22184), .B(n22183), .Z(n22202) );
  XOR U23235 ( .A(a[951]), .B(n2312), .Z(n22206) );
  AND U23236 ( .A(a[949]), .B(b[3]), .Z(n22210) );
  AND U23237 ( .A(a[953]), .B(b[0]), .Z(n22186) );
  XNOR U23238 ( .A(n22186), .B(n2175), .Z(n22188) );
  NANDN U23239 ( .A(b[0]), .B(a[952]), .Z(n22187) );
  NAND U23240 ( .A(n22188), .B(n22187), .Z(n22211) );
  XOR U23241 ( .A(n22210), .B(n22211), .Z(n22213) );
  XOR U23242 ( .A(n22212), .B(n22213), .Z(n22201) );
  NANDN U23243 ( .A(n22190), .B(n22189), .Z(n22194) );
  OR U23244 ( .A(n22192), .B(n22191), .Z(n22193) );
  AND U23245 ( .A(n22194), .B(n22193), .Z(n22200) );
  XOR U23246 ( .A(n22201), .B(n22200), .Z(n22203) );
  XOR U23247 ( .A(n22202), .B(n22203), .Z(n22216) );
  XNOR U23248 ( .A(n22216), .B(sreg[1973]), .Z(n22218) );
  NANDN U23249 ( .A(n22195), .B(sreg[1972]), .Z(n22199) );
  NAND U23250 ( .A(n22197), .B(n22196), .Z(n22198) );
  NAND U23251 ( .A(n22199), .B(n22198), .Z(n22217) );
  XOR U23252 ( .A(n22218), .B(n22217), .Z(c[1973]) );
  NANDN U23253 ( .A(n22201), .B(n22200), .Z(n22205) );
  OR U23254 ( .A(n22203), .B(n22202), .Z(n22204) );
  AND U23255 ( .A(n22205), .B(n22204), .Z(n22223) );
  XOR U23256 ( .A(a[952]), .B(n2312), .Z(n22227) );
  AND U23257 ( .A(a[950]), .B(b[3]), .Z(n22231) );
  AND U23258 ( .A(a[954]), .B(b[0]), .Z(n22207) );
  XNOR U23259 ( .A(n22207), .B(n2175), .Z(n22209) );
  NANDN U23260 ( .A(b[0]), .B(a[953]), .Z(n22208) );
  NAND U23261 ( .A(n22209), .B(n22208), .Z(n22232) );
  XOR U23262 ( .A(n22231), .B(n22232), .Z(n22234) );
  XOR U23263 ( .A(n22233), .B(n22234), .Z(n22222) );
  NANDN U23264 ( .A(n22211), .B(n22210), .Z(n22215) );
  OR U23265 ( .A(n22213), .B(n22212), .Z(n22214) );
  AND U23266 ( .A(n22215), .B(n22214), .Z(n22221) );
  XOR U23267 ( .A(n22222), .B(n22221), .Z(n22224) );
  XOR U23268 ( .A(n22223), .B(n22224), .Z(n22237) );
  XNOR U23269 ( .A(n22237), .B(sreg[1974]), .Z(n22239) );
  NANDN U23270 ( .A(n22216), .B(sreg[1973]), .Z(n22220) );
  NAND U23271 ( .A(n22218), .B(n22217), .Z(n22219) );
  NAND U23272 ( .A(n22220), .B(n22219), .Z(n22238) );
  XOR U23273 ( .A(n22239), .B(n22238), .Z(c[1974]) );
  NANDN U23274 ( .A(n22222), .B(n22221), .Z(n22226) );
  OR U23275 ( .A(n22224), .B(n22223), .Z(n22225) );
  AND U23276 ( .A(n22226), .B(n22225), .Z(n22244) );
  XOR U23277 ( .A(a[953]), .B(n2312), .Z(n22248) );
  AND U23278 ( .A(a[955]), .B(b[0]), .Z(n22228) );
  XNOR U23279 ( .A(n22228), .B(n2175), .Z(n22230) );
  NANDN U23280 ( .A(b[0]), .B(a[954]), .Z(n22229) );
  NAND U23281 ( .A(n22230), .B(n22229), .Z(n22253) );
  AND U23282 ( .A(a[951]), .B(b[3]), .Z(n22252) );
  XOR U23283 ( .A(n22253), .B(n22252), .Z(n22255) );
  XOR U23284 ( .A(n22254), .B(n22255), .Z(n22243) );
  NANDN U23285 ( .A(n22232), .B(n22231), .Z(n22236) );
  OR U23286 ( .A(n22234), .B(n22233), .Z(n22235) );
  AND U23287 ( .A(n22236), .B(n22235), .Z(n22242) );
  XOR U23288 ( .A(n22243), .B(n22242), .Z(n22245) );
  XOR U23289 ( .A(n22244), .B(n22245), .Z(n22258) );
  XNOR U23290 ( .A(n22258), .B(sreg[1975]), .Z(n22260) );
  NANDN U23291 ( .A(n22237), .B(sreg[1974]), .Z(n22241) );
  NAND U23292 ( .A(n22239), .B(n22238), .Z(n22240) );
  NAND U23293 ( .A(n22241), .B(n22240), .Z(n22259) );
  XOR U23294 ( .A(n22260), .B(n22259), .Z(c[1975]) );
  NANDN U23295 ( .A(n22243), .B(n22242), .Z(n22247) );
  OR U23296 ( .A(n22245), .B(n22244), .Z(n22246) );
  AND U23297 ( .A(n22247), .B(n22246), .Z(n22265) );
  XOR U23298 ( .A(a[954]), .B(n2312), .Z(n22269) );
  AND U23299 ( .A(a[956]), .B(b[0]), .Z(n22249) );
  XNOR U23300 ( .A(n22249), .B(n2175), .Z(n22251) );
  NANDN U23301 ( .A(b[0]), .B(a[955]), .Z(n22250) );
  NAND U23302 ( .A(n22251), .B(n22250), .Z(n22274) );
  AND U23303 ( .A(a[952]), .B(b[3]), .Z(n22273) );
  XOR U23304 ( .A(n22274), .B(n22273), .Z(n22276) );
  XOR U23305 ( .A(n22275), .B(n22276), .Z(n22264) );
  NANDN U23306 ( .A(n22253), .B(n22252), .Z(n22257) );
  OR U23307 ( .A(n22255), .B(n22254), .Z(n22256) );
  AND U23308 ( .A(n22257), .B(n22256), .Z(n22263) );
  XOR U23309 ( .A(n22264), .B(n22263), .Z(n22266) );
  XOR U23310 ( .A(n22265), .B(n22266), .Z(n22279) );
  XNOR U23311 ( .A(n22279), .B(sreg[1976]), .Z(n22281) );
  NANDN U23312 ( .A(n22258), .B(sreg[1975]), .Z(n22262) );
  NAND U23313 ( .A(n22260), .B(n22259), .Z(n22261) );
  NAND U23314 ( .A(n22262), .B(n22261), .Z(n22280) );
  XOR U23315 ( .A(n22281), .B(n22280), .Z(c[1976]) );
  NANDN U23316 ( .A(n22264), .B(n22263), .Z(n22268) );
  OR U23317 ( .A(n22266), .B(n22265), .Z(n22267) );
  AND U23318 ( .A(n22268), .B(n22267), .Z(n22286) );
  XOR U23319 ( .A(a[955]), .B(n2312), .Z(n22290) );
  AND U23320 ( .A(a[957]), .B(b[0]), .Z(n22270) );
  XNOR U23321 ( .A(n22270), .B(n2175), .Z(n22272) );
  NANDN U23322 ( .A(b[0]), .B(a[956]), .Z(n22271) );
  NAND U23323 ( .A(n22272), .B(n22271), .Z(n22295) );
  AND U23324 ( .A(a[953]), .B(b[3]), .Z(n22294) );
  XOR U23325 ( .A(n22295), .B(n22294), .Z(n22297) );
  XOR U23326 ( .A(n22296), .B(n22297), .Z(n22285) );
  NANDN U23327 ( .A(n22274), .B(n22273), .Z(n22278) );
  OR U23328 ( .A(n22276), .B(n22275), .Z(n22277) );
  AND U23329 ( .A(n22278), .B(n22277), .Z(n22284) );
  XOR U23330 ( .A(n22285), .B(n22284), .Z(n22287) );
  XOR U23331 ( .A(n22286), .B(n22287), .Z(n22300) );
  XNOR U23332 ( .A(n22300), .B(sreg[1977]), .Z(n22302) );
  NANDN U23333 ( .A(n22279), .B(sreg[1976]), .Z(n22283) );
  NAND U23334 ( .A(n22281), .B(n22280), .Z(n22282) );
  NAND U23335 ( .A(n22283), .B(n22282), .Z(n22301) );
  XOR U23336 ( .A(n22302), .B(n22301), .Z(c[1977]) );
  NANDN U23337 ( .A(n22285), .B(n22284), .Z(n22289) );
  OR U23338 ( .A(n22287), .B(n22286), .Z(n22288) );
  AND U23339 ( .A(n22289), .B(n22288), .Z(n22307) );
  XOR U23340 ( .A(a[956]), .B(n2312), .Z(n22311) );
  AND U23341 ( .A(a[954]), .B(b[3]), .Z(n22315) );
  AND U23342 ( .A(a[958]), .B(b[0]), .Z(n22291) );
  XNOR U23343 ( .A(n22291), .B(n2175), .Z(n22293) );
  NANDN U23344 ( .A(b[0]), .B(a[957]), .Z(n22292) );
  NAND U23345 ( .A(n22293), .B(n22292), .Z(n22316) );
  XOR U23346 ( .A(n22315), .B(n22316), .Z(n22318) );
  XOR U23347 ( .A(n22317), .B(n22318), .Z(n22306) );
  NANDN U23348 ( .A(n22295), .B(n22294), .Z(n22299) );
  OR U23349 ( .A(n22297), .B(n22296), .Z(n22298) );
  AND U23350 ( .A(n22299), .B(n22298), .Z(n22305) );
  XOR U23351 ( .A(n22306), .B(n22305), .Z(n22308) );
  XOR U23352 ( .A(n22307), .B(n22308), .Z(n22321) );
  XNOR U23353 ( .A(n22321), .B(sreg[1978]), .Z(n22323) );
  NANDN U23354 ( .A(n22300), .B(sreg[1977]), .Z(n22304) );
  NAND U23355 ( .A(n22302), .B(n22301), .Z(n22303) );
  NAND U23356 ( .A(n22304), .B(n22303), .Z(n22322) );
  XOR U23357 ( .A(n22323), .B(n22322), .Z(c[1978]) );
  NANDN U23358 ( .A(n22306), .B(n22305), .Z(n22310) );
  OR U23359 ( .A(n22308), .B(n22307), .Z(n22309) );
  AND U23360 ( .A(n22310), .B(n22309), .Z(n22329) );
  XOR U23361 ( .A(a[957]), .B(n2312), .Z(n22330) );
  NAND U23362 ( .A(a[959]), .B(b[0]), .Z(n22312) );
  XNOR U23363 ( .A(b[1]), .B(n22312), .Z(n22314) );
  NANDN U23364 ( .A(b[0]), .B(a[958]), .Z(n22313) );
  AND U23365 ( .A(n22314), .B(n22313), .Z(n22334) );
  AND U23366 ( .A(a[955]), .B(b[3]), .Z(n22335) );
  XOR U23367 ( .A(n22334), .B(n22335), .Z(n22336) );
  XNOR U23368 ( .A(n22337), .B(n22336), .Z(n22326) );
  NANDN U23369 ( .A(n22316), .B(n22315), .Z(n22320) );
  OR U23370 ( .A(n22318), .B(n22317), .Z(n22319) );
  AND U23371 ( .A(n22320), .B(n22319), .Z(n22327) );
  XNOR U23372 ( .A(n22326), .B(n22327), .Z(n22328) );
  XNOR U23373 ( .A(n22329), .B(n22328), .Z(n22340) );
  XNOR U23374 ( .A(n22340), .B(sreg[1979]), .Z(n22342) );
  NANDN U23375 ( .A(n22321), .B(sreg[1978]), .Z(n22325) );
  NAND U23376 ( .A(n22323), .B(n22322), .Z(n22324) );
  NAND U23377 ( .A(n22325), .B(n22324), .Z(n22341) );
  XOR U23378 ( .A(n22342), .B(n22341), .Z(c[1979]) );
  XOR U23379 ( .A(a[958]), .B(n2313), .Z(n22349) );
  AND U23380 ( .A(a[960]), .B(b[0]), .Z(n22331) );
  XNOR U23381 ( .A(n22331), .B(n2175), .Z(n22333) );
  NANDN U23382 ( .A(b[0]), .B(a[959]), .Z(n22332) );
  NAND U23383 ( .A(n22333), .B(n22332), .Z(n22354) );
  AND U23384 ( .A(a[956]), .B(b[3]), .Z(n22353) );
  XOR U23385 ( .A(n22354), .B(n22353), .Z(n22356) );
  XOR U23386 ( .A(n22355), .B(n22356), .Z(n22344) );
  NAND U23387 ( .A(n22335), .B(n22334), .Z(n22339) );
  NANDN U23388 ( .A(n22337), .B(n22336), .Z(n22338) );
  AND U23389 ( .A(n22339), .B(n22338), .Z(n22343) );
  XOR U23390 ( .A(n22344), .B(n22343), .Z(n22346) );
  XOR U23391 ( .A(n22345), .B(n22346), .Z(n22359) );
  XNOR U23392 ( .A(n22359), .B(sreg[1980]), .Z(n22361) );
  XOR U23393 ( .A(n22361), .B(n22360), .Z(c[1980]) );
  NANDN U23394 ( .A(n22344), .B(n22343), .Z(n22348) );
  OR U23395 ( .A(n22346), .B(n22345), .Z(n22347) );
  AND U23396 ( .A(n22348), .B(n22347), .Z(n22366) );
  XOR U23397 ( .A(a[959]), .B(n2313), .Z(n22370) );
  AND U23398 ( .A(a[961]), .B(b[0]), .Z(n22350) );
  XNOR U23399 ( .A(n22350), .B(n2175), .Z(n22352) );
  NANDN U23400 ( .A(b[0]), .B(a[960]), .Z(n22351) );
  NAND U23401 ( .A(n22352), .B(n22351), .Z(n22375) );
  AND U23402 ( .A(a[957]), .B(b[3]), .Z(n22374) );
  XOR U23403 ( .A(n22375), .B(n22374), .Z(n22377) );
  XOR U23404 ( .A(n22376), .B(n22377), .Z(n22365) );
  NANDN U23405 ( .A(n22354), .B(n22353), .Z(n22358) );
  OR U23406 ( .A(n22356), .B(n22355), .Z(n22357) );
  AND U23407 ( .A(n22358), .B(n22357), .Z(n22364) );
  XOR U23408 ( .A(n22365), .B(n22364), .Z(n22367) );
  XOR U23409 ( .A(n22366), .B(n22367), .Z(n22380) );
  XNOR U23410 ( .A(n22380), .B(sreg[1981]), .Z(n22382) );
  NANDN U23411 ( .A(n22359), .B(sreg[1980]), .Z(n22363) );
  NAND U23412 ( .A(n22361), .B(n22360), .Z(n22362) );
  NAND U23413 ( .A(n22363), .B(n22362), .Z(n22381) );
  XOR U23414 ( .A(n22382), .B(n22381), .Z(c[1981]) );
  NANDN U23415 ( .A(n22365), .B(n22364), .Z(n22369) );
  OR U23416 ( .A(n22367), .B(n22366), .Z(n22368) );
  AND U23417 ( .A(n22369), .B(n22368), .Z(n22387) );
  XOR U23418 ( .A(a[960]), .B(n2313), .Z(n22391) );
  AND U23419 ( .A(a[962]), .B(b[0]), .Z(n22371) );
  XNOR U23420 ( .A(n22371), .B(n2175), .Z(n22373) );
  NANDN U23421 ( .A(b[0]), .B(a[961]), .Z(n22372) );
  NAND U23422 ( .A(n22373), .B(n22372), .Z(n22396) );
  AND U23423 ( .A(a[958]), .B(b[3]), .Z(n22395) );
  XOR U23424 ( .A(n22396), .B(n22395), .Z(n22398) );
  XOR U23425 ( .A(n22397), .B(n22398), .Z(n22386) );
  NANDN U23426 ( .A(n22375), .B(n22374), .Z(n22379) );
  OR U23427 ( .A(n22377), .B(n22376), .Z(n22378) );
  AND U23428 ( .A(n22379), .B(n22378), .Z(n22385) );
  XOR U23429 ( .A(n22386), .B(n22385), .Z(n22388) );
  XOR U23430 ( .A(n22387), .B(n22388), .Z(n22401) );
  XNOR U23431 ( .A(n22401), .B(sreg[1982]), .Z(n22403) );
  NANDN U23432 ( .A(n22380), .B(sreg[1981]), .Z(n22384) );
  NAND U23433 ( .A(n22382), .B(n22381), .Z(n22383) );
  NAND U23434 ( .A(n22384), .B(n22383), .Z(n22402) );
  XOR U23435 ( .A(n22403), .B(n22402), .Z(c[1982]) );
  NANDN U23436 ( .A(n22386), .B(n22385), .Z(n22390) );
  OR U23437 ( .A(n22388), .B(n22387), .Z(n22389) );
  AND U23438 ( .A(n22390), .B(n22389), .Z(n22408) );
  XOR U23439 ( .A(a[961]), .B(n2313), .Z(n22412) );
  AND U23440 ( .A(a[959]), .B(b[3]), .Z(n22416) );
  AND U23441 ( .A(a[963]), .B(b[0]), .Z(n22392) );
  XNOR U23442 ( .A(n22392), .B(n2175), .Z(n22394) );
  NANDN U23443 ( .A(b[0]), .B(a[962]), .Z(n22393) );
  NAND U23444 ( .A(n22394), .B(n22393), .Z(n22417) );
  XOR U23445 ( .A(n22416), .B(n22417), .Z(n22419) );
  XOR U23446 ( .A(n22418), .B(n22419), .Z(n22407) );
  NANDN U23447 ( .A(n22396), .B(n22395), .Z(n22400) );
  OR U23448 ( .A(n22398), .B(n22397), .Z(n22399) );
  AND U23449 ( .A(n22400), .B(n22399), .Z(n22406) );
  XOR U23450 ( .A(n22407), .B(n22406), .Z(n22409) );
  XOR U23451 ( .A(n22408), .B(n22409), .Z(n22422) );
  XNOR U23452 ( .A(n22422), .B(sreg[1983]), .Z(n22424) );
  NANDN U23453 ( .A(n22401), .B(sreg[1982]), .Z(n22405) );
  NAND U23454 ( .A(n22403), .B(n22402), .Z(n22404) );
  NAND U23455 ( .A(n22405), .B(n22404), .Z(n22423) );
  XOR U23456 ( .A(n22424), .B(n22423), .Z(c[1983]) );
  NANDN U23457 ( .A(n22407), .B(n22406), .Z(n22411) );
  OR U23458 ( .A(n22409), .B(n22408), .Z(n22410) );
  AND U23459 ( .A(n22411), .B(n22410), .Z(n22429) );
  XOR U23460 ( .A(a[962]), .B(n2313), .Z(n22433) );
  AND U23461 ( .A(a[960]), .B(b[3]), .Z(n22437) );
  AND U23462 ( .A(a[964]), .B(b[0]), .Z(n22413) );
  XNOR U23463 ( .A(n22413), .B(n2175), .Z(n22415) );
  NANDN U23464 ( .A(b[0]), .B(a[963]), .Z(n22414) );
  NAND U23465 ( .A(n22415), .B(n22414), .Z(n22438) );
  XOR U23466 ( .A(n22437), .B(n22438), .Z(n22440) );
  XOR U23467 ( .A(n22439), .B(n22440), .Z(n22428) );
  NANDN U23468 ( .A(n22417), .B(n22416), .Z(n22421) );
  OR U23469 ( .A(n22419), .B(n22418), .Z(n22420) );
  AND U23470 ( .A(n22421), .B(n22420), .Z(n22427) );
  XOR U23471 ( .A(n22428), .B(n22427), .Z(n22430) );
  XOR U23472 ( .A(n22429), .B(n22430), .Z(n22443) );
  XNOR U23473 ( .A(n22443), .B(sreg[1984]), .Z(n22445) );
  NANDN U23474 ( .A(n22422), .B(sreg[1983]), .Z(n22426) );
  NAND U23475 ( .A(n22424), .B(n22423), .Z(n22425) );
  NAND U23476 ( .A(n22426), .B(n22425), .Z(n22444) );
  XOR U23477 ( .A(n22445), .B(n22444), .Z(c[1984]) );
  NANDN U23478 ( .A(n22428), .B(n22427), .Z(n22432) );
  OR U23479 ( .A(n22430), .B(n22429), .Z(n22431) );
  AND U23480 ( .A(n22432), .B(n22431), .Z(n22450) );
  XOR U23481 ( .A(a[963]), .B(n2313), .Z(n22454) );
  AND U23482 ( .A(a[965]), .B(b[0]), .Z(n22434) );
  XNOR U23483 ( .A(n22434), .B(n2175), .Z(n22436) );
  NANDN U23484 ( .A(b[0]), .B(a[964]), .Z(n22435) );
  NAND U23485 ( .A(n22436), .B(n22435), .Z(n22459) );
  AND U23486 ( .A(a[961]), .B(b[3]), .Z(n22458) );
  XOR U23487 ( .A(n22459), .B(n22458), .Z(n22461) );
  XOR U23488 ( .A(n22460), .B(n22461), .Z(n22449) );
  NANDN U23489 ( .A(n22438), .B(n22437), .Z(n22442) );
  OR U23490 ( .A(n22440), .B(n22439), .Z(n22441) );
  AND U23491 ( .A(n22442), .B(n22441), .Z(n22448) );
  XOR U23492 ( .A(n22449), .B(n22448), .Z(n22451) );
  XOR U23493 ( .A(n22450), .B(n22451), .Z(n22464) );
  XNOR U23494 ( .A(n22464), .B(sreg[1985]), .Z(n22466) );
  NANDN U23495 ( .A(n22443), .B(sreg[1984]), .Z(n22447) );
  NAND U23496 ( .A(n22445), .B(n22444), .Z(n22446) );
  NAND U23497 ( .A(n22447), .B(n22446), .Z(n22465) );
  XOR U23498 ( .A(n22466), .B(n22465), .Z(c[1985]) );
  NANDN U23499 ( .A(n22449), .B(n22448), .Z(n22453) );
  OR U23500 ( .A(n22451), .B(n22450), .Z(n22452) );
  AND U23501 ( .A(n22453), .B(n22452), .Z(n22471) );
  XOR U23502 ( .A(a[964]), .B(n2313), .Z(n22475) );
  AND U23503 ( .A(a[966]), .B(b[0]), .Z(n22455) );
  XNOR U23504 ( .A(n22455), .B(n2175), .Z(n22457) );
  NANDN U23505 ( .A(b[0]), .B(a[965]), .Z(n22456) );
  NAND U23506 ( .A(n22457), .B(n22456), .Z(n22480) );
  AND U23507 ( .A(a[962]), .B(b[3]), .Z(n22479) );
  XOR U23508 ( .A(n22480), .B(n22479), .Z(n22482) );
  XOR U23509 ( .A(n22481), .B(n22482), .Z(n22470) );
  NANDN U23510 ( .A(n22459), .B(n22458), .Z(n22463) );
  OR U23511 ( .A(n22461), .B(n22460), .Z(n22462) );
  AND U23512 ( .A(n22463), .B(n22462), .Z(n22469) );
  XOR U23513 ( .A(n22470), .B(n22469), .Z(n22472) );
  XOR U23514 ( .A(n22471), .B(n22472), .Z(n22485) );
  XNOR U23515 ( .A(n22485), .B(sreg[1986]), .Z(n22487) );
  NANDN U23516 ( .A(n22464), .B(sreg[1985]), .Z(n22468) );
  NAND U23517 ( .A(n22466), .B(n22465), .Z(n22467) );
  NAND U23518 ( .A(n22468), .B(n22467), .Z(n22486) );
  XOR U23519 ( .A(n22487), .B(n22486), .Z(c[1986]) );
  NANDN U23520 ( .A(n22470), .B(n22469), .Z(n22474) );
  OR U23521 ( .A(n22472), .B(n22471), .Z(n22473) );
  AND U23522 ( .A(n22474), .B(n22473), .Z(n22492) );
  XOR U23523 ( .A(a[965]), .B(n2314), .Z(n22496) );
  AND U23524 ( .A(a[963]), .B(b[3]), .Z(n22500) );
  AND U23525 ( .A(a[967]), .B(b[0]), .Z(n22476) );
  XNOR U23526 ( .A(n22476), .B(n2175), .Z(n22478) );
  NANDN U23527 ( .A(b[0]), .B(a[966]), .Z(n22477) );
  NAND U23528 ( .A(n22478), .B(n22477), .Z(n22501) );
  XOR U23529 ( .A(n22500), .B(n22501), .Z(n22503) );
  XOR U23530 ( .A(n22502), .B(n22503), .Z(n22491) );
  NANDN U23531 ( .A(n22480), .B(n22479), .Z(n22484) );
  OR U23532 ( .A(n22482), .B(n22481), .Z(n22483) );
  AND U23533 ( .A(n22484), .B(n22483), .Z(n22490) );
  XOR U23534 ( .A(n22491), .B(n22490), .Z(n22493) );
  XOR U23535 ( .A(n22492), .B(n22493), .Z(n22506) );
  XNOR U23536 ( .A(n22506), .B(sreg[1987]), .Z(n22508) );
  NANDN U23537 ( .A(n22485), .B(sreg[1986]), .Z(n22489) );
  NAND U23538 ( .A(n22487), .B(n22486), .Z(n22488) );
  NAND U23539 ( .A(n22489), .B(n22488), .Z(n22507) );
  XOR U23540 ( .A(n22508), .B(n22507), .Z(c[1987]) );
  NANDN U23541 ( .A(n22491), .B(n22490), .Z(n22495) );
  OR U23542 ( .A(n22493), .B(n22492), .Z(n22494) );
  AND U23543 ( .A(n22495), .B(n22494), .Z(n22513) );
  XOR U23544 ( .A(a[966]), .B(n2314), .Z(n22517) );
  AND U23545 ( .A(a[968]), .B(b[0]), .Z(n22497) );
  XNOR U23546 ( .A(n22497), .B(n2175), .Z(n22499) );
  NANDN U23547 ( .A(b[0]), .B(a[967]), .Z(n22498) );
  NAND U23548 ( .A(n22499), .B(n22498), .Z(n22522) );
  AND U23549 ( .A(a[964]), .B(b[3]), .Z(n22521) );
  XOR U23550 ( .A(n22522), .B(n22521), .Z(n22524) );
  XOR U23551 ( .A(n22523), .B(n22524), .Z(n22512) );
  NANDN U23552 ( .A(n22501), .B(n22500), .Z(n22505) );
  OR U23553 ( .A(n22503), .B(n22502), .Z(n22504) );
  AND U23554 ( .A(n22505), .B(n22504), .Z(n22511) );
  XOR U23555 ( .A(n22512), .B(n22511), .Z(n22514) );
  XOR U23556 ( .A(n22513), .B(n22514), .Z(n22527) );
  XNOR U23557 ( .A(n22527), .B(sreg[1988]), .Z(n22529) );
  NANDN U23558 ( .A(n22506), .B(sreg[1987]), .Z(n22510) );
  NAND U23559 ( .A(n22508), .B(n22507), .Z(n22509) );
  NAND U23560 ( .A(n22510), .B(n22509), .Z(n22528) );
  XOR U23561 ( .A(n22529), .B(n22528), .Z(c[1988]) );
  NANDN U23562 ( .A(n22512), .B(n22511), .Z(n22516) );
  OR U23563 ( .A(n22514), .B(n22513), .Z(n22515) );
  AND U23564 ( .A(n22516), .B(n22515), .Z(n22534) );
  XOR U23565 ( .A(a[967]), .B(n2314), .Z(n22538) );
  AND U23566 ( .A(a[969]), .B(b[0]), .Z(n22518) );
  XNOR U23567 ( .A(n22518), .B(n2175), .Z(n22520) );
  NANDN U23568 ( .A(b[0]), .B(a[968]), .Z(n22519) );
  NAND U23569 ( .A(n22520), .B(n22519), .Z(n22543) );
  AND U23570 ( .A(a[965]), .B(b[3]), .Z(n22542) );
  XOR U23571 ( .A(n22543), .B(n22542), .Z(n22545) );
  XOR U23572 ( .A(n22544), .B(n22545), .Z(n22533) );
  NANDN U23573 ( .A(n22522), .B(n22521), .Z(n22526) );
  OR U23574 ( .A(n22524), .B(n22523), .Z(n22525) );
  AND U23575 ( .A(n22526), .B(n22525), .Z(n22532) );
  XOR U23576 ( .A(n22533), .B(n22532), .Z(n22535) );
  XOR U23577 ( .A(n22534), .B(n22535), .Z(n22548) );
  XNOR U23578 ( .A(n22548), .B(sreg[1989]), .Z(n22550) );
  NANDN U23579 ( .A(n22527), .B(sreg[1988]), .Z(n22531) );
  NAND U23580 ( .A(n22529), .B(n22528), .Z(n22530) );
  NAND U23581 ( .A(n22531), .B(n22530), .Z(n22549) );
  XOR U23582 ( .A(n22550), .B(n22549), .Z(c[1989]) );
  NANDN U23583 ( .A(n22533), .B(n22532), .Z(n22537) );
  OR U23584 ( .A(n22535), .B(n22534), .Z(n22536) );
  AND U23585 ( .A(n22537), .B(n22536), .Z(n22555) );
  XOR U23586 ( .A(a[968]), .B(n2314), .Z(n22559) );
  AND U23587 ( .A(a[970]), .B(b[0]), .Z(n22539) );
  XNOR U23588 ( .A(n22539), .B(n2175), .Z(n22541) );
  NANDN U23589 ( .A(b[0]), .B(a[969]), .Z(n22540) );
  NAND U23590 ( .A(n22541), .B(n22540), .Z(n22564) );
  AND U23591 ( .A(a[966]), .B(b[3]), .Z(n22563) );
  XOR U23592 ( .A(n22564), .B(n22563), .Z(n22566) );
  XOR U23593 ( .A(n22565), .B(n22566), .Z(n22554) );
  NANDN U23594 ( .A(n22543), .B(n22542), .Z(n22547) );
  OR U23595 ( .A(n22545), .B(n22544), .Z(n22546) );
  AND U23596 ( .A(n22547), .B(n22546), .Z(n22553) );
  XOR U23597 ( .A(n22554), .B(n22553), .Z(n22556) );
  XOR U23598 ( .A(n22555), .B(n22556), .Z(n22569) );
  XNOR U23599 ( .A(n22569), .B(sreg[1990]), .Z(n22571) );
  NANDN U23600 ( .A(n22548), .B(sreg[1989]), .Z(n22552) );
  NAND U23601 ( .A(n22550), .B(n22549), .Z(n22551) );
  NAND U23602 ( .A(n22552), .B(n22551), .Z(n22570) );
  XOR U23603 ( .A(n22571), .B(n22570), .Z(c[1990]) );
  NANDN U23604 ( .A(n22554), .B(n22553), .Z(n22558) );
  OR U23605 ( .A(n22556), .B(n22555), .Z(n22557) );
  AND U23606 ( .A(n22558), .B(n22557), .Z(n22576) );
  XOR U23607 ( .A(a[969]), .B(n2314), .Z(n22580) );
  AND U23608 ( .A(a[967]), .B(b[3]), .Z(n22584) );
  AND U23609 ( .A(a[971]), .B(b[0]), .Z(n22560) );
  XNOR U23610 ( .A(n22560), .B(n2175), .Z(n22562) );
  NANDN U23611 ( .A(b[0]), .B(a[970]), .Z(n22561) );
  NAND U23612 ( .A(n22562), .B(n22561), .Z(n22585) );
  XOR U23613 ( .A(n22584), .B(n22585), .Z(n22587) );
  XOR U23614 ( .A(n22586), .B(n22587), .Z(n22575) );
  NANDN U23615 ( .A(n22564), .B(n22563), .Z(n22568) );
  OR U23616 ( .A(n22566), .B(n22565), .Z(n22567) );
  AND U23617 ( .A(n22568), .B(n22567), .Z(n22574) );
  XOR U23618 ( .A(n22575), .B(n22574), .Z(n22577) );
  XOR U23619 ( .A(n22576), .B(n22577), .Z(n22590) );
  XNOR U23620 ( .A(n22590), .B(sreg[1991]), .Z(n22592) );
  NANDN U23621 ( .A(n22569), .B(sreg[1990]), .Z(n22573) );
  NAND U23622 ( .A(n22571), .B(n22570), .Z(n22572) );
  NAND U23623 ( .A(n22573), .B(n22572), .Z(n22591) );
  XOR U23624 ( .A(n22592), .B(n22591), .Z(c[1991]) );
  NANDN U23625 ( .A(n22575), .B(n22574), .Z(n22579) );
  OR U23626 ( .A(n22577), .B(n22576), .Z(n22578) );
  AND U23627 ( .A(n22579), .B(n22578), .Z(n22597) );
  XOR U23628 ( .A(a[970]), .B(n2314), .Z(n22601) );
  AND U23629 ( .A(a[972]), .B(b[0]), .Z(n22581) );
  XNOR U23630 ( .A(n22581), .B(n2175), .Z(n22583) );
  NANDN U23631 ( .A(b[0]), .B(a[971]), .Z(n22582) );
  NAND U23632 ( .A(n22583), .B(n22582), .Z(n22606) );
  AND U23633 ( .A(a[968]), .B(b[3]), .Z(n22605) );
  XOR U23634 ( .A(n22606), .B(n22605), .Z(n22608) );
  XOR U23635 ( .A(n22607), .B(n22608), .Z(n22596) );
  NANDN U23636 ( .A(n22585), .B(n22584), .Z(n22589) );
  OR U23637 ( .A(n22587), .B(n22586), .Z(n22588) );
  AND U23638 ( .A(n22589), .B(n22588), .Z(n22595) );
  XOR U23639 ( .A(n22596), .B(n22595), .Z(n22598) );
  XOR U23640 ( .A(n22597), .B(n22598), .Z(n22611) );
  XNOR U23641 ( .A(n22611), .B(sreg[1992]), .Z(n22613) );
  NANDN U23642 ( .A(n22590), .B(sreg[1991]), .Z(n22594) );
  NAND U23643 ( .A(n22592), .B(n22591), .Z(n22593) );
  NAND U23644 ( .A(n22594), .B(n22593), .Z(n22612) );
  XOR U23645 ( .A(n22613), .B(n22612), .Z(c[1992]) );
  NANDN U23646 ( .A(n22596), .B(n22595), .Z(n22600) );
  OR U23647 ( .A(n22598), .B(n22597), .Z(n22599) );
  AND U23648 ( .A(n22600), .B(n22599), .Z(n22618) );
  XOR U23649 ( .A(a[971]), .B(n2314), .Z(n22622) );
  AND U23650 ( .A(a[973]), .B(b[0]), .Z(n22602) );
  XNOR U23651 ( .A(n22602), .B(n2175), .Z(n22604) );
  NANDN U23652 ( .A(b[0]), .B(a[972]), .Z(n22603) );
  NAND U23653 ( .A(n22604), .B(n22603), .Z(n22627) );
  AND U23654 ( .A(a[969]), .B(b[3]), .Z(n22626) );
  XOR U23655 ( .A(n22627), .B(n22626), .Z(n22629) );
  XOR U23656 ( .A(n22628), .B(n22629), .Z(n22617) );
  NANDN U23657 ( .A(n22606), .B(n22605), .Z(n22610) );
  OR U23658 ( .A(n22608), .B(n22607), .Z(n22609) );
  AND U23659 ( .A(n22610), .B(n22609), .Z(n22616) );
  XOR U23660 ( .A(n22617), .B(n22616), .Z(n22619) );
  XOR U23661 ( .A(n22618), .B(n22619), .Z(n22632) );
  XNOR U23662 ( .A(n22632), .B(sreg[1993]), .Z(n22634) );
  NANDN U23663 ( .A(n22611), .B(sreg[1992]), .Z(n22615) );
  NAND U23664 ( .A(n22613), .B(n22612), .Z(n22614) );
  NAND U23665 ( .A(n22615), .B(n22614), .Z(n22633) );
  XOR U23666 ( .A(n22634), .B(n22633), .Z(c[1993]) );
  NANDN U23667 ( .A(n22617), .B(n22616), .Z(n22621) );
  OR U23668 ( .A(n22619), .B(n22618), .Z(n22620) );
  AND U23669 ( .A(n22621), .B(n22620), .Z(n22639) );
  XOR U23670 ( .A(a[972]), .B(n2315), .Z(n22643) );
  AND U23671 ( .A(a[970]), .B(b[3]), .Z(n22647) );
  AND U23672 ( .A(a[974]), .B(b[0]), .Z(n22623) );
  XNOR U23673 ( .A(n22623), .B(n2175), .Z(n22625) );
  NANDN U23674 ( .A(b[0]), .B(a[973]), .Z(n22624) );
  NAND U23675 ( .A(n22625), .B(n22624), .Z(n22648) );
  XOR U23676 ( .A(n22647), .B(n22648), .Z(n22650) );
  XOR U23677 ( .A(n22649), .B(n22650), .Z(n22638) );
  NANDN U23678 ( .A(n22627), .B(n22626), .Z(n22631) );
  OR U23679 ( .A(n22629), .B(n22628), .Z(n22630) );
  AND U23680 ( .A(n22631), .B(n22630), .Z(n22637) );
  XOR U23681 ( .A(n22638), .B(n22637), .Z(n22640) );
  XOR U23682 ( .A(n22639), .B(n22640), .Z(n22653) );
  XNOR U23683 ( .A(n22653), .B(sreg[1994]), .Z(n22655) );
  NANDN U23684 ( .A(n22632), .B(sreg[1993]), .Z(n22636) );
  NAND U23685 ( .A(n22634), .B(n22633), .Z(n22635) );
  NAND U23686 ( .A(n22636), .B(n22635), .Z(n22654) );
  XOR U23687 ( .A(n22655), .B(n22654), .Z(c[1994]) );
  NANDN U23688 ( .A(n22638), .B(n22637), .Z(n22642) );
  OR U23689 ( .A(n22640), .B(n22639), .Z(n22641) );
  AND U23690 ( .A(n22642), .B(n22641), .Z(n22660) );
  XOR U23691 ( .A(a[973]), .B(n2315), .Z(n22664) );
  AND U23692 ( .A(a[971]), .B(b[3]), .Z(n22668) );
  AND U23693 ( .A(a[975]), .B(b[0]), .Z(n22644) );
  XNOR U23694 ( .A(n22644), .B(n2175), .Z(n22646) );
  NANDN U23695 ( .A(b[0]), .B(a[974]), .Z(n22645) );
  NAND U23696 ( .A(n22646), .B(n22645), .Z(n22669) );
  XOR U23697 ( .A(n22668), .B(n22669), .Z(n22671) );
  XOR U23698 ( .A(n22670), .B(n22671), .Z(n22659) );
  NANDN U23699 ( .A(n22648), .B(n22647), .Z(n22652) );
  OR U23700 ( .A(n22650), .B(n22649), .Z(n22651) );
  AND U23701 ( .A(n22652), .B(n22651), .Z(n22658) );
  XOR U23702 ( .A(n22659), .B(n22658), .Z(n22661) );
  XOR U23703 ( .A(n22660), .B(n22661), .Z(n22674) );
  XNOR U23704 ( .A(n22674), .B(sreg[1995]), .Z(n22676) );
  NANDN U23705 ( .A(n22653), .B(sreg[1994]), .Z(n22657) );
  NAND U23706 ( .A(n22655), .B(n22654), .Z(n22656) );
  NAND U23707 ( .A(n22657), .B(n22656), .Z(n22675) );
  XOR U23708 ( .A(n22676), .B(n22675), .Z(c[1995]) );
  NANDN U23709 ( .A(n22659), .B(n22658), .Z(n22663) );
  OR U23710 ( .A(n22661), .B(n22660), .Z(n22662) );
  AND U23711 ( .A(n22663), .B(n22662), .Z(n22681) );
  XOR U23712 ( .A(a[974]), .B(n2315), .Z(n22685) );
  AND U23713 ( .A(a[972]), .B(b[3]), .Z(n22689) );
  AND U23714 ( .A(a[976]), .B(b[0]), .Z(n22665) );
  XNOR U23715 ( .A(n22665), .B(n2175), .Z(n22667) );
  NANDN U23716 ( .A(b[0]), .B(a[975]), .Z(n22666) );
  NAND U23717 ( .A(n22667), .B(n22666), .Z(n22690) );
  XOR U23718 ( .A(n22689), .B(n22690), .Z(n22692) );
  XOR U23719 ( .A(n22691), .B(n22692), .Z(n22680) );
  NANDN U23720 ( .A(n22669), .B(n22668), .Z(n22673) );
  OR U23721 ( .A(n22671), .B(n22670), .Z(n22672) );
  AND U23722 ( .A(n22673), .B(n22672), .Z(n22679) );
  XOR U23723 ( .A(n22680), .B(n22679), .Z(n22682) );
  XOR U23724 ( .A(n22681), .B(n22682), .Z(n22695) );
  XNOR U23725 ( .A(n22695), .B(sreg[1996]), .Z(n22697) );
  NANDN U23726 ( .A(n22674), .B(sreg[1995]), .Z(n22678) );
  NAND U23727 ( .A(n22676), .B(n22675), .Z(n22677) );
  NAND U23728 ( .A(n22678), .B(n22677), .Z(n22696) );
  XOR U23729 ( .A(n22697), .B(n22696), .Z(c[1996]) );
  NANDN U23730 ( .A(n22680), .B(n22679), .Z(n22684) );
  OR U23731 ( .A(n22682), .B(n22681), .Z(n22683) );
  AND U23732 ( .A(n22684), .B(n22683), .Z(n22702) );
  XOR U23733 ( .A(a[975]), .B(n2315), .Z(n22706) );
  AND U23734 ( .A(a[973]), .B(b[3]), .Z(n22710) );
  AND U23735 ( .A(a[977]), .B(b[0]), .Z(n22686) );
  XNOR U23736 ( .A(n22686), .B(n2175), .Z(n22688) );
  NANDN U23737 ( .A(b[0]), .B(a[976]), .Z(n22687) );
  NAND U23738 ( .A(n22688), .B(n22687), .Z(n22711) );
  XOR U23739 ( .A(n22710), .B(n22711), .Z(n22713) );
  XOR U23740 ( .A(n22712), .B(n22713), .Z(n22701) );
  NANDN U23741 ( .A(n22690), .B(n22689), .Z(n22694) );
  OR U23742 ( .A(n22692), .B(n22691), .Z(n22693) );
  AND U23743 ( .A(n22694), .B(n22693), .Z(n22700) );
  XOR U23744 ( .A(n22701), .B(n22700), .Z(n22703) );
  XOR U23745 ( .A(n22702), .B(n22703), .Z(n22716) );
  XNOR U23746 ( .A(n22716), .B(sreg[1997]), .Z(n22718) );
  NANDN U23747 ( .A(n22695), .B(sreg[1996]), .Z(n22699) );
  NAND U23748 ( .A(n22697), .B(n22696), .Z(n22698) );
  NAND U23749 ( .A(n22699), .B(n22698), .Z(n22717) );
  XOR U23750 ( .A(n22718), .B(n22717), .Z(c[1997]) );
  NANDN U23751 ( .A(n22701), .B(n22700), .Z(n22705) );
  OR U23752 ( .A(n22703), .B(n22702), .Z(n22704) );
  AND U23753 ( .A(n22705), .B(n22704), .Z(n22723) );
  XOR U23754 ( .A(a[976]), .B(n2315), .Z(n22727) );
  AND U23755 ( .A(a[978]), .B(b[0]), .Z(n22707) );
  XNOR U23756 ( .A(n22707), .B(n2175), .Z(n22709) );
  NANDN U23757 ( .A(b[0]), .B(a[977]), .Z(n22708) );
  NAND U23758 ( .A(n22709), .B(n22708), .Z(n22732) );
  AND U23759 ( .A(a[974]), .B(b[3]), .Z(n22731) );
  XOR U23760 ( .A(n22732), .B(n22731), .Z(n22734) );
  XOR U23761 ( .A(n22733), .B(n22734), .Z(n22722) );
  NANDN U23762 ( .A(n22711), .B(n22710), .Z(n22715) );
  OR U23763 ( .A(n22713), .B(n22712), .Z(n22714) );
  AND U23764 ( .A(n22715), .B(n22714), .Z(n22721) );
  XOR U23765 ( .A(n22722), .B(n22721), .Z(n22724) );
  XOR U23766 ( .A(n22723), .B(n22724), .Z(n22737) );
  XNOR U23767 ( .A(n22737), .B(sreg[1998]), .Z(n22739) );
  NANDN U23768 ( .A(n22716), .B(sreg[1997]), .Z(n22720) );
  NAND U23769 ( .A(n22718), .B(n22717), .Z(n22719) );
  NAND U23770 ( .A(n22720), .B(n22719), .Z(n22738) );
  XOR U23771 ( .A(n22739), .B(n22738), .Z(c[1998]) );
  NANDN U23772 ( .A(n22722), .B(n22721), .Z(n22726) );
  OR U23773 ( .A(n22724), .B(n22723), .Z(n22725) );
  AND U23774 ( .A(n22726), .B(n22725), .Z(n22744) );
  XOR U23775 ( .A(a[977]), .B(n2315), .Z(n22748) );
  AND U23776 ( .A(a[975]), .B(b[3]), .Z(n22752) );
  AND U23777 ( .A(a[979]), .B(b[0]), .Z(n22728) );
  XNOR U23778 ( .A(n22728), .B(n2175), .Z(n22730) );
  NANDN U23779 ( .A(b[0]), .B(a[978]), .Z(n22729) );
  NAND U23780 ( .A(n22730), .B(n22729), .Z(n22753) );
  XOR U23781 ( .A(n22752), .B(n22753), .Z(n22755) );
  XOR U23782 ( .A(n22754), .B(n22755), .Z(n22743) );
  NANDN U23783 ( .A(n22732), .B(n22731), .Z(n22736) );
  OR U23784 ( .A(n22734), .B(n22733), .Z(n22735) );
  AND U23785 ( .A(n22736), .B(n22735), .Z(n22742) );
  XOR U23786 ( .A(n22743), .B(n22742), .Z(n22745) );
  XOR U23787 ( .A(n22744), .B(n22745), .Z(n22758) );
  XNOR U23788 ( .A(n22758), .B(sreg[1999]), .Z(n22760) );
  NANDN U23789 ( .A(n22737), .B(sreg[1998]), .Z(n22741) );
  NAND U23790 ( .A(n22739), .B(n22738), .Z(n22740) );
  NAND U23791 ( .A(n22741), .B(n22740), .Z(n22759) );
  XOR U23792 ( .A(n22760), .B(n22759), .Z(c[1999]) );
  NANDN U23793 ( .A(n22743), .B(n22742), .Z(n22747) );
  OR U23794 ( .A(n22745), .B(n22744), .Z(n22746) );
  AND U23795 ( .A(n22747), .B(n22746), .Z(n22765) );
  XOR U23796 ( .A(a[978]), .B(n2315), .Z(n22769) );
  AND U23797 ( .A(a[980]), .B(b[0]), .Z(n22749) );
  XNOR U23798 ( .A(n22749), .B(n2175), .Z(n22751) );
  NANDN U23799 ( .A(b[0]), .B(a[979]), .Z(n22750) );
  NAND U23800 ( .A(n22751), .B(n22750), .Z(n22774) );
  AND U23801 ( .A(a[976]), .B(b[3]), .Z(n22773) );
  XOR U23802 ( .A(n22774), .B(n22773), .Z(n22776) );
  XOR U23803 ( .A(n22775), .B(n22776), .Z(n22764) );
  NANDN U23804 ( .A(n22753), .B(n22752), .Z(n22757) );
  OR U23805 ( .A(n22755), .B(n22754), .Z(n22756) );
  AND U23806 ( .A(n22757), .B(n22756), .Z(n22763) );
  XOR U23807 ( .A(n22764), .B(n22763), .Z(n22766) );
  XOR U23808 ( .A(n22765), .B(n22766), .Z(n22779) );
  XNOR U23809 ( .A(n22779), .B(sreg[2000]), .Z(n22781) );
  NANDN U23810 ( .A(n22758), .B(sreg[1999]), .Z(n22762) );
  NAND U23811 ( .A(n22760), .B(n22759), .Z(n22761) );
  NAND U23812 ( .A(n22762), .B(n22761), .Z(n22780) );
  XOR U23813 ( .A(n22781), .B(n22780), .Z(c[2000]) );
  NANDN U23814 ( .A(n22764), .B(n22763), .Z(n22768) );
  OR U23815 ( .A(n22766), .B(n22765), .Z(n22767) );
  AND U23816 ( .A(n22768), .B(n22767), .Z(n22786) );
  XOR U23817 ( .A(a[979]), .B(n2316), .Z(n22790) );
  AND U23818 ( .A(a[981]), .B(b[0]), .Z(n22770) );
  XNOR U23819 ( .A(n22770), .B(n2175), .Z(n22772) );
  NANDN U23820 ( .A(b[0]), .B(a[980]), .Z(n22771) );
  NAND U23821 ( .A(n22772), .B(n22771), .Z(n22795) );
  AND U23822 ( .A(a[977]), .B(b[3]), .Z(n22794) );
  XOR U23823 ( .A(n22795), .B(n22794), .Z(n22797) );
  XOR U23824 ( .A(n22796), .B(n22797), .Z(n22785) );
  NANDN U23825 ( .A(n22774), .B(n22773), .Z(n22778) );
  OR U23826 ( .A(n22776), .B(n22775), .Z(n22777) );
  AND U23827 ( .A(n22778), .B(n22777), .Z(n22784) );
  XOR U23828 ( .A(n22785), .B(n22784), .Z(n22787) );
  XOR U23829 ( .A(n22786), .B(n22787), .Z(n22800) );
  XNOR U23830 ( .A(n22800), .B(sreg[2001]), .Z(n22802) );
  NANDN U23831 ( .A(n22779), .B(sreg[2000]), .Z(n22783) );
  NAND U23832 ( .A(n22781), .B(n22780), .Z(n22782) );
  NAND U23833 ( .A(n22783), .B(n22782), .Z(n22801) );
  XOR U23834 ( .A(n22802), .B(n22801), .Z(c[2001]) );
  NANDN U23835 ( .A(n22785), .B(n22784), .Z(n22789) );
  OR U23836 ( .A(n22787), .B(n22786), .Z(n22788) );
  AND U23837 ( .A(n22789), .B(n22788), .Z(n22807) );
  XOR U23838 ( .A(a[980]), .B(n2316), .Z(n22811) );
  AND U23839 ( .A(a[982]), .B(b[0]), .Z(n22791) );
  XNOR U23840 ( .A(n22791), .B(n2175), .Z(n22793) );
  NANDN U23841 ( .A(b[0]), .B(a[981]), .Z(n22792) );
  NAND U23842 ( .A(n22793), .B(n22792), .Z(n22816) );
  AND U23843 ( .A(a[978]), .B(b[3]), .Z(n22815) );
  XOR U23844 ( .A(n22816), .B(n22815), .Z(n22818) );
  XOR U23845 ( .A(n22817), .B(n22818), .Z(n22806) );
  NANDN U23846 ( .A(n22795), .B(n22794), .Z(n22799) );
  OR U23847 ( .A(n22797), .B(n22796), .Z(n22798) );
  AND U23848 ( .A(n22799), .B(n22798), .Z(n22805) );
  XOR U23849 ( .A(n22806), .B(n22805), .Z(n22808) );
  XOR U23850 ( .A(n22807), .B(n22808), .Z(n22821) );
  XNOR U23851 ( .A(n22821), .B(sreg[2002]), .Z(n22823) );
  NANDN U23852 ( .A(n22800), .B(sreg[2001]), .Z(n22804) );
  NAND U23853 ( .A(n22802), .B(n22801), .Z(n22803) );
  NAND U23854 ( .A(n22804), .B(n22803), .Z(n22822) );
  XOR U23855 ( .A(n22823), .B(n22822), .Z(c[2002]) );
  NANDN U23856 ( .A(n22806), .B(n22805), .Z(n22810) );
  OR U23857 ( .A(n22808), .B(n22807), .Z(n22809) );
  AND U23858 ( .A(n22810), .B(n22809), .Z(n22828) );
  XOR U23859 ( .A(a[981]), .B(n2316), .Z(n22832) );
  AND U23860 ( .A(a[979]), .B(b[3]), .Z(n22836) );
  AND U23861 ( .A(a[983]), .B(b[0]), .Z(n22812) );
  XNOR U23862 ( .A(n22812), .B(n2175), .Z(n22814) );
  NANDN U23863 ( .A(b[0]), .B(a[982]), .Z(n22813) );
  NAND U23864 ( .A(n22814), .B(n22813), .Z(n22837) );
  XOR U23865 ( .A(n22836), .B(n22837), .Z(n22839) );
  XOR U23866 ( .A(n22838), .B(n22839), .Z(n22827) );
  NANDN U23867 ( .A(n22816), .B(n22815), .Z(n22820) );
  OR U23868 ( .A(n22818), .B(n22817), .Z(n22819) );
  AND U23869 ( .A(n22820), .B(n22819), .Z(n22826) );
  XOR U23870 ( .A(n22827), .B(n22826), .Z(n22829) );
  XOR U23871 ( .A(n22828), .B(n22829), .Z(n22842) );
  XNOR U23872 ( .A(n22842), .B(sreg[2003]), .Z(n22844) );
  NANDN U23873 ( .A(n22821), .B(sreg[2002]), .Z(n22825) );
  NAND U23874 ( .A(n22823), .B(n22822), .Z(n22824) );
  NAND U23875 ( .A(n22825), .B(n22824), .Z(n22843) );
  XOR U23876 ( .A(n22844), .B(n22843), .Z(c[2003]) );
  NANDN U23877 ( .A(n22827), .B(n22826), .Z(n22831) );
  OR U23878 ( .A(n22829), .B(n22828), .Z(n22830) );
  AND U23879 ( .A(n22831), .B(n22830), .Z(n22849) );
  XOR U23880 ( .A(a[982]), .B(n2316), .Z(n22853) );
  AND U23881 ( .A(a[984]), .B(b[0]), .Z(n22833) );
  XNOR U23882 ( .A(n22833), .B(n2175), .Z(n22835) );
  NANDN U23883 ( .A(b[0]), .B(a[983]), .Z(n22834) );
  NAND U23884 ( .A(n22835), .B(n22834), .Z(n22858) );
  AND U23885 ( .A(a[980]), .B(b[3]), .Z(n22857) );
  XOR U23886 ( .A(n22858), .B(n22857), .Z(n22860) );
  XOR U23887 ( .A(n22859), .B(n22860), .Z(n22848) );
  NANDN U23888 ( .A(n22837), .B(n22836), .Z(n22841) );
  OR U23889 ( .A(n22839), .B(n22838), .Z(n22840) );
  AND U23890 ( .A(n22841), .B(n22840), .Z(n22847) );
  XOR U23891 ( .A(n22848), .B(n22847), .Z(n22850) );
  XOR U23892 ( .A(n22849), .B(n22850), .Z(n22863) );
  XNOR U23893 ( .A(n22863), .B(sreg[2004]), .Z(n22865) );
  NANDN U23894 ( .A(n22842), .B(sreg[2003]), .Z(n22846) );
  NAND U23895 ( .A(n22844), .B(n22843), .Z(n22845) );
  NAND U23896 ( .A(n22846), .B(n22845), .Z(n22864) );
  XOR U23897 ( .A(n22865), .B(n22864), .Z(c[2004]) );
  NANDN U23898 ( .A(n22848), .B(n22847), .Z(n22852) );
  OR U23899 ( .A(n22850), .B(n22849), .Z(n22851) );
  AND U23900 ( .A(n22852), .B(n22851), .Z(n22870) );
  XOR U23901 ( .A(a[983]), .B(n2316), .Z(n22874) );
  AND U23902 ( .A(a[981]), .B(b[3]), .Z(n22878) );
  AND U23903 ( .A(a[985]), .B(b[0]), .Z(n22854) );
  XNOR U23904 ( .A(n22854), .B(n2175), .Z(n22856) );
  NANDN U23905 ( .A(b[0]), .B(a[984]), .Z(n22855) );
  NAND U23906 ( .A(n22856), .B(n22855), .Z(n22879) );
  XOR U23907 ( .A(n22878), .B(n22879), .Z(n22881) );
  XOR U23908 ( .A(n22880), .B(n22881), .Z(n22869) );
  NANDN U23909 ( .A(n22858), .B(n22857), .Z(n22862) );
  OR U23910 ( .A(n22860), .B(n22859), .Z(n22861) );
  AND U23911 ( .A(n22862), .B(n22861), .Z(n22868) );
  XOR U23912 ( .A(n22869), .B(n22868), .Z(n22871) );
  XOR U23913 ( .A(n22870), .B(n22871), .Z(n22884) );
  XNOR U23914 ( .A(n22884), .B(sreg[2005]), .Z(n22886) );
  NANDN U23915 ( .A(n22863), .B(sreg[2004]), .Z(n22867) );
  NAND U23916 ( .A(n22865), .B(n22864), .Z(n22866) );
  NAND U23917 ( .A(n22867), .B(n22866), .Z(n22885) );
  XOR U23918 ( .A(n22886), .B(n22885), .Z(c[2005]) );
  NANDN U23919 ( .A(n22869), .B(n22868), .Z(n22873) );
  OR U23920 ( .A(n22871), .B(n22870), .Z(n22872) );
  AND U23921 ( .A(n22873), .B(n22872), .Z(n22891) );
  XOR U23922 ( .A(a[984]), .B(n2316), .Z(n22895) );
  AND U23923 ( .A(a[986]), .B(b[0]), .Z(n22875) );
  XNOR U23924 ( .A(n22875), .B(n2175), .Z(n22877) );
  NANDN U23925 ( .A(b[0]), .B(a[985]), .Z(n22876) );
  NAND U23926 ( .A(n22877), .B(n22876), .Z(n22900) );
  AND U23927 ( .A(a[982]), .B(b[3]), .Z(n22899) );
  XOR U23928 ( .A(n22900), .B(n22899), .Z(n22902) );
  XOR U23929 ( .A(n22901), .B(n22902), .Z(n22890) );
  NANDN U23930 ( .A(n22879), .B(n22878), .Z(n22883) );
  OR U23931 ( .A(n22881), .B(n22880), .Z(n22882) );
  AND U23932 ( .A(n22883), .B(n22882), .Z(n22889) );
  XOR U23933 ( .A(n22890), .B(n22889), .Z(n22892) );
  XOR U23934 ( .A(n22891), .B(n22892), .Z(n22905) );
  XNOR U23935 ( .A(n22905), .B(sreg[2006]), .Z(n22907) );
  NANDN U23936 ( .A(n22884), .B(sreg[2005]), .Z(n22888) );
  NAND U23937 ( .A(n22886), .B(n22885), .Z(n22887) );
  NAND U23938 ( .A(n22888), .B(n22887), .Z(n22906) );
  XOR U23939 ( .A(n22907), .B(n22906), .Z(c[2006]) );
  NANDN U23940 ( .A(n22890), .B(n22889), .Z(n22894) );
  OR U23941 ( .A(n22892), .B(n22891), .Z(n22893) );
  AND U23942 ( .A(n22894), .B(n22893), .Z(n22912) );
  XOR U23943 ( .A(a[985]), .B(n2316), .Z(n22916) );
  AND U23944 ( .A(a[987]), .B(b[0]), .Z(n22896) );
  XNOR U23945 ( .A(n22896), .B(n2175), .Z(n22898) );
  NANDN U23946 ( .A(b[0]), .B(a[986]), .Z(n22897) );
  NAND U23947 ( .A(n22898), .B(n22897), .Z(n22921) );
  AND U23948 ( .A(a[983]), .B(b[3]), .Z(n22920) );
  XOR U23949 ( .A(n22921), .B(n22920), .Z(n22923) );
  XOR U23950 ( .A(n22922), .B(n22923), .Z(n22911) );
  NANDN U23951 ( .A(n22900), .B(n22899), .Z(n22904) );
  OR U23952 ( .A(n22902), .B(n22901), .Z(n22903) );
  AND U23953 ( .A(n22904), .B(n22903), .Z(n22910) );
  XOR U23954 ( .A(n22911), .B(n22910), .Z(n22913) );
  XOR U23955 ( .A(n22912), .B(n22913), .Z(n22926) );
  XNOR U23956 ( .A(n22926), .B(sreg[2007]), .Z(n22928) );
  NANDN U23957 ( .A(n22905), .B(sreg[2006]), .Z(n22909) );
  NAND U23958 ( .A(n22907), .B(n22906), .Z(n22908) );
  NAND U23959 ( .A(n22909), .B(n22908), .Z(n22927) );
  XOR U23960 ( .A(n22928), .B(n22927), .Z(c[2007]) );
  NANDN U23961 ( .A(n22911), .B(n22910), .Z(n22915) );
  OR U23962 ( .A(n22913), .B(n22912), .Z(n22914) );
  AND U23963 ( .A(n22915), .B(n22914), .Z(n22933) );
  XOR U23964 ( .A(a[986]), .B(n2317), .Z(n22937) );
  AND U23965 ( .A(a[988]), .B(b[0]), .Z(n22917) );
  XNOR U23966 ( .A(n22917), .B(n2175), .Z(n22919) );
  NANDN U23967 ( .A(b[0]), .B(a[987]), .Z(n22918) );
  NAND U23968 ( .A(n22919), .B(n22918), .Z(n22942) );
  AND U23969 ( .A(a[984]), .B(b[3]), .Z(n22941) );
  XOR U23970 ( .A(n22942), .B(n22941), .Z(n22944) );
  XOR U23971 ( .A(n22943), .B(n22944), .Z(n22932) );
  NANDN U23972 ( .A(n22921), .B(n22920), .Z(n22925) );
  OR U23973 ( .A(n22923), .B(n22922), .Z(n22924) );
  AND U23974 ( .A(n22925), .B(n22924), .Z(n22931) );
  XOR U23975 ( .A(n22932), .B(n22931), .Z(n22934) );
  XOR U23976 ( .A(n22933), .B(n22934), .Z(n22947) );
  XNOR U23977 ( .A(n22947), .B(sreg[2008]), .Z(n22949) );
  NANDN U23978 ( .A(n22926), .B(sreg[2007]), .Z(n22930) );
  NAND U23979 ( .A(n22928), .B(n22927), .Z(n22929) );
  NAND U23980 ( .A(n22930), .B(n22929), .Z(n22948) );
  XOR U23981 ( .A(n22949), .B(n22948), .Z(c[2008]) );
  NANDN U23982 ( .A(n22932), .B(n22931), .Z(n22936) );
  OR U23983 ( .A(n22934), .B(n22933), .Z(n22935) );
  AND U23984 ( .A(n22936), .B(n22935), .Z(n22954) );
  XOR U23985 ( .A(a[987]), .B(n2317), .Z(n22958) );
  AND U23986 ( .A(a[985]), .B(b[3]), .Z(n22962) );
  AND U23987 ( .A(a[989]), .B(b[0]), .Z(n22938) );
  XNOR U23988 ( .A(n22938), .B(n2175), .Z(n22940) );
  NANDN U23989 ( .A(b[0]), .B(a[988]), .Z(n22939) );
  NAND U23990 ( .A(n22940), .B(n22939), .Z(n22963) );
  XOR U23991 ( .A(n22962), .B(n22963), .Z(n22965) );
  XOR U23992 ( .A(n22964), .B(n22965), .Z(n22953) );
  NANDN U23993 ( .A(n22942), .B(n22941), .Z(n22946) );
  OR U23994 ( .A(n22944), .B(n22943), .Z(n22945) );
  AND U23995 ( .A(n22946), .B(n22945), .Z(n22952) );
  XOR U23996 ( .A(n22953), .B(n22952), .Z(n22955) );
  XOR U23997 ( .A(n22954), .B(n22955), .Z(n22968) );
  XNOR U23998 ( .A(n22968), .B(sreg[2009]), .Z(n22970) );
  NANDN U23999 ( .A(n22947), .B(sreg[2008]), .Z(n22951) );
  NAND U24000 ( .A(n22949), .B(n22948), .Z(n22950) );
  NAND U24001 ( .A(n22951), .B(n22950), .Z(n22969) );
  XOR U24002 ( .A(n22970), .B(n22969), .Z(c[2009]) );
  NANDN U24003 ( .A(n22953), .B(n22952), .Z(n22957) );
  OR U24004 ( .A(n22955), .B(n22954), .Z(n22956) );
  AND U24005 ( .A(n22957), .B(n22956), .Z(n22975) );
  XOR U24006 ( .A(a[988]), .B(n2317), .Z(n22979) );
  AND U24007 ( .A(a[990]), .B(b[0]), .Z(n22959) );
  XNOR U24008 ( .A(n22959), .B(n2175), .Z(n22961) );
  NANDN U24009 ( .A(b[0]), .B(a[989]), .Z(n22960) );
  NAND U24010 ( .A(n22961), .B(n22960), .Z(n22984) );
  AND U24011 ( .A(a[986]), .B(b[3]), .Z(n22983) );
  XOR U24012 ( .A(n22984), .B(n22983), .Z(n22986) );
  XOR U24013 ( .A(n22985), .B(n22986), .Z(n22974) );
  NANDN U24014 ( .A(n22963), .B(n22962), .Z(n22967) );
  OR U24015 ( .A(n22965), .B(n22964), .Z(n22966) );
  AND U24016 ( .A(n22967), .B(n22966), .Z(n22973) );
  XOR U24017 ( .A(n22974), .B(n22973), .Z(n22976) );
  XOR U24018 ( .A(n22975), .B(n22976), .Z(n22989) );
  XNOR U24019 ( .A(n22989), .B(sreg[2010]), .Z(n22991) );
  NANDN U24020 ( .A(n22968), .B(sreg[2009]), .Z(n22972) );
  NAND U24021 ( .A(n22970), .B(n22969), .Z(n22971) );
  NAND U24022 ( .A(n22972), .B(n22971), .Z(n22990) );
  XOR U24023 ( .A(n22991), .B(n22990), .Z(c[2010]) );
  NANDN U24024 ( .A(n22974), .B(n22973), .Z(n22978) );
  OR U24025 ( .A(n22976), .B(n22975), .Z(n22977) );
  AND U24026 ( .A(n22978), .B(n22977), .Z(n22996) );
  XOR U24027 ( .A(a[989]), .B(n2317), .Z(n23000) );
  AND U24028 ( .A(a[987]), .B(b[3]), .Z(n23004) );
  AND U24029 ( .A(a[991]), .B(b[0]), .Z(n22980) );
  XNOR U24030 ( .A(n22980), .B(n2175), .Z(n22982) );
  NANDN U24031 ( .A(b[0]), .B(a[990]), .Z(n22981) );
  NAND U24032 ( .A(n22982), .B(n22981), .Z(n23005) );
  XOR U24033 ( .A(n23004), .B(n23005), .Z(n23007) );
  XOR U24034 ( .A(n23006), .B(n23007), .Z(n22995) );
  NANDN U24035 ( .A(n22984), .B(n22983), .Z(n22988) );
  OR U24036 ( .A(n22986), .B(n22985), .Z(n22987) );
  AND U24037 ( .A(n22988), .B(n22987), .Z(n22994) );
  XOR U24038 ( .A(n22995), .B(n22994), .Z(n22997) );
  XOR U24039 ( .A(n22996), .B(n22997), .Z(n23010) );
  XNOR U24040 ( .A(n23010), .B(sreg[2011]), .Z(n23012) );
  NANDN U24041 ( .A(n22989), .B(sreg[2010]), .Z(n22993) );
  NAND U24042 ( .A(n22991), .B(n22990), .Z(n22992) );
  NAND U24043 ( .A(n22993), .B(n22992), .Z(n23011) );
  XOR U24044 ( .A(n23012), .B(n23011), .Z(c[2011]) );
  NANDN U24045 ( .A(n22995), .B(n22994), .Z(n22999) );
  OR U24046 ( .A(n22997), .B(n22996), .Z(n22998) );
  AND U24047 ( .A(n22999), .B(n22998), .Z(n23017) );
  XOR U24048 ( .A(a[990]), .B(n2317), .Z(n23021) );
  AND U24049 ( .A(a[988]), .B(b[3]), .Z(n23025) );
  AND U24050 ( .A(a[992]), .B(b[0]), .Z(n23001) );
  XNOR U24051 ( .A(n23001), .B(n2175), .Z(n23003) );
  NANDN U24052 ( .A(b[0]), .B(a[991]), .Z(n23002) );
  NAND U24053 ( .A(n23003), .B(n23002), .Z(n23026) );
  XOR U24054 ( .A(n23025), .B(n23026), .Z(n23028) );
  XOR U24055 ( .A(n23027), .B(n23028), .Z(n23016) );
  NANDN U24056 ( .A(n23005), .B(n23004), .Z(n23009) );
  OR U24057 ( .A(n23007), .B(n23006), .Z(n23008) );
  AND U24058 ( .A(n23009), .B(n23008), .Z(n23015) );
  XOR U24059 ( .A(n23016), .B(n23015), .Z(n23018) );
  XOR U24060 ( .A(n23017), .B(n23018), .Z(n23031) );
  XNOR U24061 ( .A(n23031), .B(sreg[2012]), .Z(n23033) );
  NANDN U24062 ( .A(n23010), .B(sreg[2011]), .Z(n23014) );
  NAND U24063 ( .A(n23012), .B(n23011), .Z(n23013) );
  NAND U24064 ( .A(n23014), .B(n23013), .Z(n23032) );
  XOR U24065 ( .A(n23033), .B(n23032), .Z(c[2012]) );
  NANDN U24066 ( .A(n23016), .B(n23015), .Z(n23020) );
  OR U24067 ( .A(n23018), .B(n23017), .Z(n23019) );
  AND U24068 ( .A(n23020), .B(n23019), .Z(n23038) );
  XOR U24069 ( .A(a[991]), .B(n2317), .Z(n23042) );
  AND U24070 ( .A(a[993]), .B(b[0]), .Z(n23022) );
  XNOR U24071 ( .A(n23022), .B(n2175), .Z(n23024) );
  NANDN U24072 ( .A(b[0]), .B(a[992]), .Z(n23023) );
  NAND U24073 ( .A(n23024), .B(n23023), .Z(n23047) );
  AND U24074 ( .A(a[989]), .B(b[3]), .Z(n23046) );
  XOR U24075 ( .A(n23047), .B(n23046), .Z(n23049) );
  XOR U24076 ( .A(n23048), .B(n23049), .Z(n23037) );
  NANDN U24077 ( .A(n23026), .B(n23025), .Z(n23030) );
  OR U24078 ( .A(n23028), .B(n23027), .Z(n23029) );
  AND U24079 ( .A(n23030), .B(n23029), .Z(n23036) );
  XOR U24080 ( .A(n23037), .B(n23036), .Z(n23039) );
  XOR U24081 ( .A(n23038), .B(n23039), .Z(n23052) );
  XNOR U24082 ( .A(n23052), .B(sreg[2013]), .Z(n23054) );
  NANDN U24083 ( .A(n23031), .B(sreg[2012]), .Z(n23035) );
  NAND U24084 ( .A(n23033), .B(n23032), .Z(n23034) );
  NAND U24085 ( .A(n23035), .B(n23034), .Z(n23053) );
  XOR U24086 ( .A(n23054), .B(n23053), .Z(c[2013]) );
  NANDN U24087 ( .A(n23037), .B(n23036), .Z(n23041) );
  OR U24088 ( .A(n23039), .B(n23038), .Z(n23040) );
  AND U24089 ( .A(n23041), .B(n23040), .Z(n23059) );
  XOR U24090 ( .A(a[992]), .B(n2317), .Z(n23063) );
  AND U24091 ( .A(a[990]), .B(b[3]), .Z(n23067) );
  AND U24092 ( .A(a[994]), .B(b[0]), .Z(n23043) );
  XNOR U24093 ( .A(n23043), .B(n2175), .Z(n23045) );
  NANDN U24094 ( .A(b[0]), .B(a[993]), .Z(n23044) );
  NAND U24095 ( .A(n23045), .B(n23044), .Z(n23068) );
  XOR U24096 ( .A(n23067), .B(n23068), .Z(n23070) );
  XOR U24097 ( .A(n23069), .B(n23070), .Z(n23058) );
  NANDN U24098 ( .A(n23047), .B(n23046), .Z(n23051) );
  OR U24099 ( .A(n23049), .B(n23048), .Z(n23050) );
  AND U24100 ( .A(n23051), .B(n23050), .Z(n23057) );
  XOR U24101 ( .A(n23058), .B(n23057), .Z(n23060) );
  XOR U24102 ( .A(n23059), .B(n23060), .Z(n23073) );
  XNOR U24103 ( .A(n23073), .B(sreg[2014]), .Z(n23075) );
  NANDN U24104 ( .A(n23052), .B(sreg[2013]), .Z(n23056) );
  NAND U24105 ( .A(n23054), .B(n23053), .Z(n23055) );
  NAND U24106 ( .A(n23056), .B(n23055), .Z(n23074) );
  XOR U24107 ( .A(n23075), .B(n23074), .Z(c[2014]) );
  NANDN U24108 ( .A(n23058), .B(n23057), .Z(n23062) );
  OR U24109 ( .A(n23060), .B(n23059), .Z(n23061) );
  AND U24110 ( .A(n23062), .B(n23061), .Z(n23080) );
  XOR U24111 ( .A(a[993]), .B(n2318), .Z(n23084) );
  AND U24112 ( .A(a[991]), .B(b[3]), .Z(n23088) );
  AND U24113 ( .A(a[995]), .B(b[0]), .Z(n23064) );
  XNOR U24114 ( .A(n23064), .B(n2175), .Z(n23066) );
  NANDN U24115 ( .A(b[0]), .B(a[994]), .Z(n23065) );
  NAND U24116 ( .A(n23066), .B(n23065), .Z(n23089) );
  XOR U24117 ( .A(n23088), .B(n23089), .Z(n23091) );
  XOR U24118 ( .A(n23090), .B(n23091), .Z(n23079) );
  NANDN U24119 ( .A(n23068), .B(n23067), .Z(n23072) );
  OR U24120 ( .A(n23070), .B(n23069), .Z(n23071) );
  AND U24121 ( .A(n23072), .B(n23071), .Z(n23078) );
  XOR U24122 ( .A(n23079), .B(n23078), .Z(n23081) );
  XOR U24123 ( .A(n23080), .B(n23081), .Z(n23094) );
  XNOR U24124 ( .A(n23094), .B(sreg[2015]), .Z(n23096) );
  NANDN U24125 ( .A(n23073), .B(sreg[2014]), .Z(n23077) );
  NAND U24126 ( .A(n23075), .B(n23074), .Z(n23076) );
  NAND U24127 ( .A(n23077), .B(n23076), .Z(n23095) );
  XOR U24128 ( .A(n23096), .B(n23095), .Z(c[2015]) );
  NANDN U24129 ( .A(n23079), .B(n23078), .Z(n23083) );
  OR U24130 ( .A(n23081), .B(n23080), .Z(n23082) );
  AND U24131 ( .A(n23083), .B(n23082), .Z(n23101) );
  XOR U24132 ( .A(a[994]), .B(n2318), .Z(n23105) );
  AND U24133 ( .A(a[996]), .B(b[0]), .Z(n23085) );
  XNOR U24134 ( .A(n23085), .B(n2175), .Z(n23087) );
  NANDN U24135 ( .A(b[0]), .B(a[995]), .Z(n23086) );
  NAND U24136 ( .A(n23087), .B(n23086), .Z(n23110) );
  AND U24137 ( .A(a[992]), .B(b[3]), .Z(n23109) );
  XOR U24138 ( .A(n23110), .B(n23109), .Z(n23112) );
  XOR U24139 ( .A(n23111), .B(n23112), .Z(n23100) );
  NANDN U24140 ( .A(n23089), .B(n23088), .Z(n23093) );
  OR U24141 ( .A(n23091), .B(n23090), .Z(n23092) );
  AND U24142 ( .A(n23093), .B(n23092), .Z(n23099) );
  XOR U24143 ( .A(n23100), .B(n23099), .Z(n23102) );
  XOR U24144 ( .A(n23101), .B(n23102), .Z(n23115) );
  XNOR U24145 ( .A(n23115), .B(sreg[2016]), .Z(n23117) );
  NANDN U24146 ( .A(n23094), .B(sreg[2015]), .Z(n23098) );
  NAND U24147 ( .A(n23096), .B(n23095), .Z(n23097) );
  NAND U24148 ( .A(n23098), .B(n23097), .Z(n23116) );
  XOR U24149 ( .A(n23117), .B(n23116), .Z(c[2016]) );
  NANDN U24150 ( .A(n23100), .B(n23099), .Z(n23104) );
  OR U24151 ( .A(n23102), .B(n23101), .Z(n23103) );
  AND U24152 ( .A(n23104), .B(n23103), .Z(n23122) );
  XOR U24153 ( .A(a[995]), .B(n2318), .Z(n23126) );
  AND U24154 ( .A(a[997]), .B(b[0]), .Z(n23106) );
  XNOR U24155 ( .A(n23106), .B(n2175), .Z(n23108) );
  NANDN U24156 ( .A(b[0]), .B(a[996]), .Z(n23107) );
  NAND U24157 ( .A(n23108), .B(n23107), .Z(n23131) );
  AND U24158 ( .A(a[993]), .B(b[3]), .Z(n23130) );
  XOR U24159 ( .A(n23131), .B(n23130), .Z(n23133) );
  XOR U24160 ( .A(n23132), .B(n23133), .Z(n23121) );
  NANDN U24161 ( .A(n23110), .B(n23109), .Z(n23114) );
  OR U24162 ( .A(n23112), .B(n23111), .Z(n23113) );
  AND U24163 ( .A(n23114), .B(n23113), .Z(n23120) );
  XOR U24164 ( .A(n23121), .B(n23120), .Z(n23123) );
  XOR U24165 ( .A(n23122), .B(n23123), .Z(n23136) );
  XNOR U24166 ( .A(n23136), .B(sreg[2017]), .Z(n23138) );
  NANDN U24167 ( .A(n23115), .B(sreg[2016]), .Z(n23119) );
  NAND U24168 ( .A(n23117), .B(n23116), .Z(n23118) );
  NAND U24169 ( .A(n23119), .B(n23118), .Z(n23137) );
  XOR U24170 ( .A(n23138), .B(n23137), .Z(c[2017]) );
  NANDN U24171 ( .A(n23121), .B(n23120), .Z(n23125) );
  OR U24172 ( .A(n23123), .B(n23122), .Z(n23124) );
  AND U24173 ( .A(n23125), .B(n23124), .Z(n23143) );
  XOR U24174 ( .A(a[996]), .B(n2318), .Z(n23147) );
  AND U24175 ( .A(a[994]), .B(b[3]), .Z(n23151) );
  AND U24176 ( .A(a[998]), .B(b[0]), .Z(n23127) );
  XNOR U24177 ( .A(n23127), .B(n2175), .Z(n23129) );
  NANDN U24178 ( .A(b[0]), .B(a[997]), .Z(n23128) );
  NAND U24179 ( .A(n23129), .B(n23128), .Z(n23152) );
  XOR U24180 ( .A(n23151), .B(n23152), .Z(n23154) );
  XOR U24181 ( .A(n23153), .B(n23154), .Z(n23142) );
  NANDN U24182 ( .A(n23131), .B(n23130), .Z(n23135) );
  OR U24183 ( .A(n23133), .B(n23132), .Z(n23134) );
  AND U24184 ( .A(n23135), .B(n23134), .Z(n23141) );
  XOR U24185 ( .A(n23142), .B(n23141), .Z(n23144) );
  XOR U24186 ( .A(n23143), .B(n23144), .Z(n23157) );
  XNOR U24187 ( .A(n23157), .B(sreg[2018]), .Z(n23159) );
  NANDN U24188 ( .A(n23136), .B(sreg[2017]), .Z(n23140) );
  NAND U24189 ( .A(n23138), .B(n23137), .Z(n23139) );
  NAND U24190 ( .A(n23140), .B(n23139), .Z(n23158) );
  XOR U24191 ( .A(n23159), .B(n23158), .Z(c[2018]) );
  NANDN U24192 ( .A(n23142), .B(n23141), .Z(n23146) );
  OR U24193 ( .A(n23144), .B(n23143), .Z(n23145) );
  AND U24194 ( .A(n23146), .B(n23145), .Z(n23164) );
  XOR U24195 ( .A(a[997]), .B(n2318), .Z(n23168) );
  AND U24196 ( .A(a[995]), .B(b[3]), .Z(n23172) );
  AND U24197 ( .A(a[999]), .B(b[0]), .Z(n23148) );
  XNOR U24198 ( .A(n23148), .B(n2175), .Z(n23150) );
  NANDN U24199 ( .A(b[0]), .B(a[998]), .Z(n23149) );
  NAND U24200 ( .A(n23150), .B(n23149), .Z(n23173) );
  XOR U24201 ( .A(n23172), .B(n23173), .Z(n23175) );
  XOR U24202 ( .A(n23174), .B(n23175), .Z(n23163) );
  NANDN U24203 ( .A(n23152), .B(n23151), .Z(n23156) );
  OR U24204 ( .A(n23154), .B(n23153), .Z(n23155) );
  AND U24205 ( .A(n23156), .B(n23155), .Z(n23162) );
  XOR U24206 ( .A(n23163), .B(n23162), .Z(n23165) );
  XOR U24207 ( .A(n23164), .B(n23165), .Z(n23178) );
  XNOR U24208 ( .A(n23178), .B(sreg[2019]), .Z(n23180) );
  NANDN U24209 ( .A(n23157), .B(sreg[2018]), .Z(n23161) );
  NAND U24210 ( .A(n23159), .B(n23158), .Z(n23160) );
  NAND U24211 ( .A(n23161), .B(n23160), .Z(n23179) );
  XOR U24212 ( .A(n23180), .B(n23179), .Z(c[2019]) );
  NANDN U24213 ( .A(n23163), .B(n23162), .Z(n23167) );
  OR U24214 ( .A(n23165), .B(n23164), .Z(n23166) );
  AND U24215 ( .A(n23167), .B(n23166), .Z(n23185) );
  XOR U24216 ( .A(a[998]), .B(n2318), .Z(n23189) );
  AND U24217 ( .A(a[1000]), .B(b[0]), .Z(n23169) );
  XNOR U24218 ( .A(n23169), .B(n2175), .Z(n23171) );
  NANDN U24219 ( .A(b[0]), .B(a[999]), .Z(n23170) );
  NAND U24220 ( .A(n23171), .B(n23170), .Z(n23194) );
  AND U24221 ( .A(a[996]), .B(b[3]), .Z(n23193) );
  XOR U24222 ( .A(n23194), .B(n23193), .Z(n23196) );
  XOR U24223 ( .A(n23195), .B(n23196), .Z(n23184) );
  NANDN U24224 ( .A(n23173), .B(n23172), .Z(n23177) );
  OR U24225 ( .A(n23175), .B(n23174), .Z(n23176) );
  AND U24226 ( .A(n23177), .B(n23176), .Z(n23183) );
  XOR U24227 ( .A(n23184), .B(n23183), .Z(n23186) );
  XOR U24228 ( .A(n23185), .B(n23186), .Z(n23199) );
  XNOR U24229 ( .A(n23199), .B(sreg[2020]), .Z(n23201) );
  NANDN U24230 ( .A(n23178), .B(sreg[2019]), .Z(n23182) );
  NAND U24231 ( .A(n23180), .B(n23179), .Z(n23181) );
  NAND U24232 ( .A(n23182), .B(n23181), .Z(n23200) );
  XOR U24233 ( .A(n23201), .B(n23200), .Z(c[2020]) );
  NANDN U24234 ( .A(n23184), .B(n23183), .Z(n23188) );
  OR U24235 ( .A(n23186), .B(n23185), .Z(n23187) );
  AND U24236 ( .A(n23188), .B(n23187), .Z(n23206) );
  XOR U24237 ( .A(a[999]), .B(n2318), .Z(n23210) );
  AND U24238 ( .A(a[1001]), .B(b[0]), .Z(n23190) );
  XNOR U24239 ( .A(n23190), .B(n2175), .Z(n23192) );
  NANDN U24240 ( .A(b[0]), .B(a[1000]), .Z(n23191) );
  NAND U24241 ( .A(n23192), .B(n23191), .Z(n23215) );
  AND U24242 ( .A(a[997]), .B(b[3]), .Z(n23214) );
  XOR U24243 ( .A(n23215), .B(n23214), .Z(n23217) );
  XOR U24244 ( .A(n23216), .B(n23217), .Z(n23205) );
  NANDN U24245 ( .A(n23194), .B(n23193), .Z(n23198) );
  OR U24246 ( .A(n23196), .B(n23195), .Z(n23197) );
  AND U24247 ( .A(n23198), .B(n23197), .Z(n23204) );
  XOR U24248 ( .A(n23205), .B(n23204), .Z(n23207) );
  XOR U24249 ( .A(n23206), .B(n23207), .Z(n23220) );
  XNOR U24250 ( .A(n23220), .B(sreg[2021]), .Z(n23222) );
  NANDN U24251 ( .A(n23199), .B(sreg[2020]), .Z(n23203) );
  NAND U24252 ( .A(n23201), .B(n23200), .Z(n23202) );
  NAND U24253 ( .A(n23203), .B(n23202), .Z(n23221) );
  XOR U24254 ( .A(n23222), .B(n23221), .Z(c[2021]) );
  NANDN U24255 ( .A(n23205), .B(n23204), .Z(n23209) );
  OR U24256 ( .A(n23207), .B(n23206), .Z(n23208) );
  AND U24257 ( .A(n23209), .B(n23208), .Z(n23227) );
  XOR U24258 ( .A(a[1000]), .B(n2319), .Z(n23231) );
  AND U24259 ( .A(a[1002]), .B(b[0]), .Z(n23211) );
  XNOR U24260 ( .A(n23211), .B(n2175), .Z(n23213) );
  NANDN U24261 ( .A(b[0]), .B(a[1001]), .Z(n23212) );
  NAND U24262 ( .A(n23213), .B(n23212), .Z(n23236) );
  AND U24263 ( .A(a[998]), .B(b[3]), .Z(n23235) );
  XOR U24264 ( .A(n23236), .B(n23235), .Z(n23238) );
  XOR U24265 ( .A(n23237), .B(n23238), .Z(n23226) );
  NANDN U24266 ( .A(n23215), .B(n23214), .Z(n23219) );
  OR U24267 ( .A(n23217), .B(n23216), .Z(n23218) );
  AND U24268 ( .A(n23219), .B(n23218), .Z(n23225) );
  XOR U24269 ( .A(n23226), .B(n23225), .Z(n23228) );
  XOR U24270 ( .A(n23227), .B(n23228), .Z(n23241) );
  XNOR U24271 ( .A(n23241), .B(sreg[2022]), .Z(n23243) );
  NANDN U24272 ( .A(n23220), .B(sreg[2021]), .Z(n23224) );
  NAND U24273 ( .A(n23222), .B(n23221), .Z(n23223) );
  NAND U24274 ( .A(n23224), .B(n23223), .Z(n23242) );
  XOR U24275 ( .A(n23243), .B(n23242), .Z(c[2022]) );
  NANDN U24276 ( .A(n23226), .B(n23225), .Z(n23230) );
  OR U24277 ( .A(n23228), .B(n23227), .Z(n23229) );
  AND U24278 ( .A(n23230), .B(n23229), .Z(n23248) );
  XOR U24279 ( .A(a[1001]), .B(n2319), .Z(n23252) );
  AND U24280 ( .A(a[1003]), .B(b[0]), .Z(n23232) );
  XNOR U24281 ( .A(n23232), .B(n2175), .Z(n23234) );
  NANDN U24282 ( .A(b[0]), .B(a[1002]), .Z(n23233) );
  NAND U24283 ( .A(n23234), .B(n23233), .Z(n23257) );
  AND U24284 ( .A(a[999]), .B(b[3]), .Z(n23256) );
  XOR U24285 ( .A(n23257), .B(n23256), .Z(n23259) );
  XOR U24286 ( .A(n23258), .B(n23259), .Z(n23247) );
  NANDN U24287 ( .A(n23236), .B(n23235), .Z(n23240) );
  OR U24288 ( .A(n23238), .B(n23237), .Z(n23239) );
  AND U24289 ( .A(n23240), .B(n23239), .Z(n23246) );
  XOR U24290 ( .A(n23247), .B(n23246), .Z(n23249) );
  XOR U24291 ( .A(n23248), .B(n23249), .Z(n23262) );
  XNOR U24292 ( .A(n23262), .B(sreg[2023]), .Z(n23264) );
  NANDN U24293 ( .A(n23241), .B(sreg[2022]), .Z(n23245) );
  NAND U24294 ( .A(n23243), .B(n23242), .Z(n23244) );
  NAND U24295 ( .A(n23245), .B(n23244), .Z(n23263) );
  XOR U24296 ( .A(n23264), .B(n23263), .Z(c[2023]) );
  NANDN U24297 ( .A(n23247), .B(n23246), .Z(n23251) );
  OR U24298 ( .A(n23249), .B(n23248), .Z(n23250) );
  AND U24299 ( .A(n23251), .B(n23250), .Z(n23269) );
  XOR U24300 ( .A(a[1002]), .B(n2319), .Z(n23273) );
  AND U24301 ( .A(a[1004]), .B(b[0]), .Z(n23253) );
  XNOR U24302 ( .A(n23253), .B(n2175), .Z(n23255) );
  NANDN U24303 ( .A(b[0]), .B(a[1003]), .Z(n23254) );
  NAND U24304 ( .A(n23255), .B(n23254), .Z(n23278) );
  AND U24305 ( .A(a[1000]), .B(b[3]), .Z(n23277) );
  XOR U24306 ( .A(n23278), .B(n23277), .Z(n23280) );
  XOR U24307 ( .A(n23279), .B(n23280), .Z(n23268) );
  NANDN U24308 ( .A(n23257), .B(n23256), .Z(n23261) );
  OR U24309 ( .A(n23259), .B(n23258), .Z(n23260) );
  AND U24310 ( .A(n23261), .B(n23260), .Z(n23267) );
  XOR U24311 ( .A(n23268), .B(n23267), .Z(n23270) );
  XOR U24312 ( .A(n23269), .B(n23270), .Z(n23283) );
  XNOR U24313 ( .A(n23283), .B(sreg[2024]), .Z(n23285) );
  NANDN U24314 ( .A(n23262), .B(sreg[2023]), .Z(n23266) );
  NAND U24315 ( .A(n23264), .B(n23263), .Z(n23265) );
  NAND U24316 ( .A(n23266), .B(n23265), .Z(n23284) );
  XOR U24317 ( .A(n23285), .B(n23284), .Z(c[2024]) );
  NANDN U24318 ( .A(n23268), .B(n23267), .Z(n23272) );
  OR U24319 ( .A(n23270), .B(n23269), .Z(n23271) );
  AND U24320 ( .A(n23272), .B(n23271), .Z(n23290) );
  XOR U24321 ( .A(a[1003]), .B(n2319), .Z(n23294) );
  AND U24322 ( .A(a[1005]), .B(b[0]), .Z(n23274) );
  XNOR U24323 ( .A(n23274), .B(n2175), .Z(n23276) );
  NANDN U24324 ( .A(b[0]), .B(a[1004]), .Z(n23275) );
  NAND U24325 ( .A(n23276), .B(n23275), .Z(n23299) );
  AND U24326 ( .A(a[1001]), .B(b[3]), .Z(n23298) );
  XOR U24327 ( .A(n23299), .B(n23298), .Z(n23301) );
  XOR U24328 ( .A(n23300), .B(n23301), .Z(n23289) );
  NANDN U24329 ( .A(n23278), .B(n23277), .Z(n23282) );
  OR U24330 ( .A(n23280), .B(n23279), .Z(n23281) );
  AND U24331 ( .A(n23282), .B(n23281), .Z(n23288) );
  XOR U24332 ( .A(n23289), .B(n23288), .Z(n23291) );
  XOR U24333 ( .A(n23290), .B(n23291), .Z(n23304) );
  XNOR U24334 ( .A(n23304), .B(sreg[2025]), .Z(n23306) );
  NANDN U24335 ( .A(n23283), .B(sreg[2024]), .Z(n23287) );
  NAND U24336 ( .A(n23285), .B(n23284), .Z(n23286) );
  NAND U24337 ( .A(n23287), .B(n23286), .Z(n23305) );
  XOR U24338 ( .A(n23306), .B(n23305), .Z(c[2025]) );
  NANDN U24339 ( .A(n23289), .B(n23288), .Z(n23293) );
  OR U24340 ( .A(n23291), .B(n23290), .Z(n23292) );
  AND U24341 ( .A(n23293), .B(n23292), .Z(n23311) );
  XOR U24342 ( .A(a[1004]), .B(n2319), .Z(n23315) );
  AND U24343 ( .A(a[1002]), .B(b[3]), .Z(n23319) );
  AND U24344 ( .A(a[1006]), .B(b[0]), .Z(n23295) );
  XNOR U24345 ( .A(n23295), .B(n2175), .Z(n23297) );
  NANDN U24346 ( .A(b[0]), .B(a[1005]), .Z(n23296) );
  NAND U24347 ( .A(n23297), .B(n23296), .Z(n23320) );
  XOR U24348 ( .A(n23319), .B(n23320), .Z(n23322) );
  XOR U24349 ( .A(n23321), .B(n23322), .Z(n23310) );
  NANDN U24350 ( .A(n23299), .B(n23298), .Z(n23303) );
  OR U24351 ( .A(n23301), .B(n23300), .Z(n23302) );
  AND U24352 ( .A(n23303), .B(n23302), .Z(n23309) );
  XOR U24353 ( .A(n23310), .B(n23309), .Z(n23312) );
  XOR U24354 ( .A(n23311), .B(n23312), .Z(n23325) );
  XNOR U24355 ( .A(n23325), .B(sreg[2026]), .Z(n23327) );
  NANDN U24356 ( .A(n23304), .B(sreg[2025]), .Z(n23308) );
  NAND U24357 ( .A(n23306), .B(n23305), .Z(n23307) );
  NAND U24358 ( .A(n23308), .B(n23307), .Z(n23326) );
  XOR U24359 ( .A(n23327), .B(n23326), .Z(c[2026]) );
  NANDN U24360 ( .A(n23310), .B(n23309), .Z(n23314) );
  OR U24361 ( .A(n23312), .B(n23311), .Z(n23313) );
  AND U24362 ( .A(n23314), .B(n23313), .Z(n23332) );
  XOR U24363 ( .A(a[1005]), .B(n2319), .Z(n23336) );
  AND U24364 ( .A(a[1007]), .B(b[0]), .Z(n23316) );
  XNOR U24365 ( .A(n23316), .B(n2175), .Z(n23318) );
  NANDN U24366 ( .A(b[0]), .B(a[1006]), .Z(n23317) );
  NAND U24367 ( .A(n23318), .B(n23317), .Z(n23341) );
  AND U24368 ( .A(a[1003]), .B(b[3]), .Z(n23340) );
  XOR U24369 ( .A(n23341), .B(n23340), .Z(n23343) );
  XOR U24370 ( .A(n23342), .B(n23343), .Z(n23331) );
  NANDN U24371 ( .A(n23320), .B(n23319), .Z(n23324) );
  OR U24372 ( .A(n23322), .B(n23321), .Z(n23323) );
  AND U24373 ( .A(n23324), .B(n23323), .Z(n23330) );
  XOR U24374 ( .A(n23331), .B(n23330), .Z(n23333) );
  XOR U24375 ( .A(n23332), .B(n23333), .Z(n23346) );
  XNOR U24376 ( .A(n23346), .B(sreg[2027]), .Z(n23348) );
  NANDN U24377 ( .A(n23325), .B(sreg[2026]), .Z(n23329) );
  NAND U24378 ( .A(n23327), .B(n23326), .Z(n23328) );
  NAND U24379 ( .A(n23329), .B(n23328), .Z(n23347) );
  XOR U24380 ( .A(n23348), .B(n23347), .Z(c[2027]) );
  NANDN U24381 ( .A(n23331), .B(n23330), .Z(n23335) );
  OR U24382 ( .A(n23333), .B(n23332), .Z(n23334) );
  AND U24383 ( .A(n23335), .B(n23334), .Z(n23353) );
  XOR U24384 ( .A(a[1006]), .B(n2319), .Z(n23357) );
  AND U24385 ( .A(a[1008]), .B(b[0]), .Z(n23337) );
  XNOR U24386 ( .A(n23337), .B(n2175), .Z(n23339) );
  NANDN U24387 ( .A(b[0]), .B(a[1007]), .Z(n23338) );
  NAND U24388 ( .A(n23339), .B(n23338), .Z(n23362) );
  AND U24389 ( .A(a[1004]), .B(b[3]), .Z(n23361) );
  XOR U24390 ( .A(n23362), .B(n23361), .Z(n23364) );
  XOR U24391 ( .A(n23363), .B(n23364), .Z(n23352) );
  NANDN U24392 ( .A(n23341), .B(n23340), .Z(n23345) );
  OR U24393 ( .A(n23343), .B(n23342), .Z(n23344) );
  AND U24394 ( .A(n23345), .B(n23344), .Z(n23351) );
  XOR U24395 ( .A(n23352), .B(n23351), .Z(n23354) );
  XOR U24396 ( .A(n23353), .B(n23354), .Z(n23367) );
  XNOR U24397 ( .A(n23367), .B(sreg[2028]), .Z(n23369) );
  NANDN U24398 ( .A(n23346), .B(sreg[2027]), .Z(n23350) );
  NAND U24399 ( .A(n23348), .B(n23347), .Z(n23349) );
  NAND U24400 ( .A(n23350), .B(n23349), .Z(n23368) );
  XOR U24401 ( .A(n23369), .B(n23368), .Z(c[2028]) );
  NANDN U24402 ( .A(n23352), .B(n23351), .Z(n23356) );
  OR U24403 ( .A(n23354), .B(n23353), .Z(n23355) );
  AND U24404 ( .A(n23356), .B(n23355), .Z(n23374) );
  XOR U24405 ( .A(a[1007]), .B(n2320), .Z(n23378) );
  AND U24406 ( .A(a[1005]), .B(b[3]), .Z(n23382) );
  AND U24407 ( .A(a[1009]), .B(b[0]), .Z(n23358) );
  XNOR U24408 ( .A(n23358), .B(n2175), .Z(n23360) );
  NANDN U24409 ( .A(b[0]), .B(a[1008]), .Z(n23359) );
  NAND U24410 ( .A(n23360), .B(n23359), .Z(n23383) );
  XOR U24411 ( .A(n23382), .B(n23383), .Z(n23385) );
  XOR U24412 ( .A(n23384), .B(n23385), .Z(n23373) );
  NANDN U24413 ( .A(n23362), .B(n23361), .Z(n23366) );
  OR U24414 ( .A(n23364), .B(n23363), .Z(n23365) );
  AND U24415 ( .A(n23366), .B(n23365), .Z(n23372) );
  XOR U24416 ( .A(n23373), .B(n23372), .Z(n23375) );
  XOR U24417 ( .A(n23374), .B(n23375), .Z(n23388) );
  XNOR U24418 ( .A(n23388), .B(sreg[2029]), .Z(n23390) );
  NANDN U24419 ( .A(n23367), .B(sreg[2028]), .Z(n23371) );
  NAND U24420 ( .A(n23369), .B(n23368), .Z(n23370) );
  NAND U24421 ( .A(n23371), .B(n23370), .Z(n23389) );
  XOR U24422 ( .A(n23390), .B(n23389), .Z(c[2029]) );
  NANDN U24423 ( .A(n23373), .B(n23372), .Z(n23377) );
  OR U24424 ( .A(n23375), .B(n23374), .Z(n23376) );
  AND U24425 ( .A(n23377), .B(n23376), .Z(n23395) );
  XOR U24426 ( .A(a[1008]), .B(n2320), .Z(n23399) );
  AND U24427 ( .A(a[1006]), .B(b[3]), .Z(n23403) );
  AND U24428 ( .A(a[1010]), .B(b[0]), .Z(n23379) );
  XNOR U24429 ( .A(n23379), .B(n2175), .Z(n23381) );
  NANDN U24430 ( .A(b[0]), .B(a[1009]), .Z(n23380) );
  NAND U24431 ( .A(n23381), .B(n23380), .Z(n23404) );
  XOR U24432 ( .A(n23403), .B(n23404), .Z(n23406) );
  XOR U24433 ( .A(n23405), .B(n23406), .Z(n23394) );
  NANDN U24434 ( .A(n23383), .B(n23382), .Z(n23387) );
  OR U24435 ( .A(n23385), .B(n23384), .Z(n23386) );
  AND U24436 ( .A(n23387), .B(n23386), .Z(n23393) );
  XOR U24437 ( .A(n23394), .B(n23393), .Z(n23396) );
  XOR U24438 ( .A(n23395), .B(n23396), .Z(n23409) );
  XNOR U24439 ( .A(n23409), .B(sreg[2030]), .Z(n23411) );
  NANDN U24440 ( .A(n23388), .B(sreg[2029]), .Z(n23392) );
  NAND U24441 ( .A(n23390), .B(n23389), .Z(n23391) );
  NAND U24442 ( .A(n23392), .B(n23391), .Z(n23410) );
  XOR U24443 ( .A(n23411), .B(n23410), .Z(c[2030]) );
  NANDN U24444 ( .A(n23394), .B(n23393), .Z(n23398) );
  OR U24445 ( .A(n23396), .B(n23395), .Z(n23397) );
  AND U24446 ( .A(n23398), .B(n23397), .Z(n23416) );
  XOR U24447 ( .A(a[1009]), .B(n2320), .Z(n23420) );
  AND U24448 ( .A(a[1011]), .B(b[0]), .Z(n23400) );
  XNOR U24449 ( .A(n23400), .B(n2175), .Z(n23402) );
  NANDN U24450 ( .A(b[0]), .B(a[1010]), .Z(n23401) );
  NAND U24451 ( .A(n23402), .B(n23401), .Z(n23425) );
  AND U24452 ( .A(a[1007]), .B(b[3]), .Z(n23424) );
  XOR U24453 ( .A(n23425), .B(n23424), .Z(n23427) );
  XOR U24454 ( .A(n23426), .B(n23427), .Z(n23415) );
  NANDN U24455 ( .A(n23404), .B(n23403), .Z(n23408) );
  OR U24456 ( .A(n23406), .B(n23405), .Z(n23407) );
  AND U24457 ( .A(n23408), .B(n23407), .Z(n23414) );
  XOR U24458 ( .A(n23415), .B(n23414), .Z(n23417) );
  XOR U24459 ( .A(n23416), .B(n23417), .Z(n23430) );
  XNOR U24460 ( .A(n23430), .B(sreg[2031]), .Z(n23432) );
  NANDN U24461 ( .A(n23409), .B(sreg[2030]), .Z(n23413) );
  NAND U24462 ( .A(n23411), .B(n23410), .Z(n23412) );
  NAND U24463 ( .A(n23413), .B(n23412), .Z(n23431) );
  XOR U24464 ( .A(n23432), .B(n23431), .Z(c[2031]) );
  NANDN U24465 ( .A(n23415), .B(n23414), .Z(n23419) );
  OR U24466 ( .A(n23417), .B(n23416), .Z(n23418) );
  AND U24467 ( .A(n23419), .B(n23418), .Z(n23437) );
  XOR U24468 ( .A(a[1010]), .B(n2320), .Z(n23441) );
  AND U24469 ( .A(a[1012]), .B(b[0]), .Z(n23421) );
  XNOR U24470 ( .A(n23421), .B(n2175), .Z(n23423) );
  NANDN U24471 ( .A(b[0]), .B(a[1011]), .Z(n23422) );
  NAND U24472 ( .A(n23423), .B(n23422), .Z(n23446) );
  AND U24473 ( .A(a[1008]), .B(b[3]), .Z(n23445) );
  XOR U24474 ( .A(n23446), .B(n23445), .Z(n23448) );
  XOR U24475 ( .A(n23447), .B(n23448), .Z(n23436) );
  NANDN U24476 ( .A(n23425), .B(n23424), .Z(n23429) );
  OR U24477 ( .A(n23427), .B(n23426), .Z(n23428) );
  AND U24478 ( .A(n23429), .B(n23428), .Z(n23435) );
  XOR U24479 ( .A(n23436), .B(n23435), .Z(n23438) );
  XOR U24480 ( .A(n23437), .B(n23438), .Z(n23451) );
  XNOR U24481 ( .A(n23451), .B(sreg[2032]), .Z(n23453) );
  NANDN U24482 ( .A(n23430), .B(sreg[2031]), .Z(n23434) );
  NAND U24483 ( .A(n23432), .B(n23431), .Z(n23433) );
  NAND U24484 ( .A(n23434), .B(n23433), .Z(n23452) );
  XOR U24485 ( .A(n23453), .B(n23452), .Z(c[2032]) );
  NANDN U24486 ( .A(n23436), .B(n23435), .Z(n23440) );
  OR U24487 ( .A(n23438), .B(n23437), .Z(n23439) );
  AND U24488 ( .A(n23440), .B(n23439), .Z(n23458) );
  XOR U24489 ( .A(a[1011]), .B(n2320), .Z(n23462) );
  AND U24490 ( .A(a[1009]), .B(b[3]), .Z(n23466) );
  AND U24491 ( .A(a[1013]), .B(b[0]), .Z(n23442) );
  XNOR U24492 ( .A(n23442), .B(n2175), .Z(n23444) );
  NANDN U24493 ( .A(b[0]), .B(a[1012]), .Z(n23443) );
  NAND U24494 ( .A(n23444), .B(n23443), .Z(n23467) );
  XOR U24495 ( .A(n23466), .B(n23467), .Z(n23469) );
  XOR U24496 ( .A(n23468), .B(n23469), .Z(n23457) );
  NANDN U24497 ( .A(n23446), .B(n23445), .Z(n23450) );
  OR U24498 ( .A(n23448), .B(n23447), .Z(n23449) );
  AND U24499 ( .A(n23450), .B(n23449), .Z(n23456) );
  XOR U24500 ( .A(n23457), .B(n23456), .Z(n23459) );
  XOR U24501 ( .A(n23458), .B(n23459), .Z(n23472) );
  XNOR U24502 ( .A(n23472), .B(sreg[2033]), .Z(n23474) );
  NANDN U24503 ( .A(n23451), .B(sreg[2032]), .Z(n23455) );
  NAND U24504 ( .A(n23453), .B(n23452), .Z(n23454) );
  NAND U24505 ( .A(n23455), .B(n23454), .Z(n23473) );
  XOR U24506 ( .A(n23474), .B(n23473), .Z(c[2033]) );
  NANDN U24507 ( .A(n23457), .B(n23456), .Z(n23461) );
  OR U24508 ( .A(n23459), .B(n23458), .Z(n23460) );
  AND U24509 ( .A(n23461), .B(n23460), .Z(n23479) );
  XOR U24510 ( .A(a[1012]), .B(n2320), .Z(n23483) );
  AND U24511 ( .A(a[1014]), .B(b[0]), .Z(n23463) );
  XNOR U24512 ( .A(n23463), .B(n2175), .Z(n23465) );
  NANDN U24513 ( .A(b[0]), .B(a[1013]), .Z(n23464) );
  NAND U24514 ( .A(n23465), .B(n23464), .Z(n23488) );
  AND U24515 ( .A(a[1010]), .B(b[3]), .Z(n23487) );
  XOR U24516 ( .A(n23488), .B(n23487), .Z(n23490) );
  XOR U24517 ( .A(n23489), .B(n23490), .Z(n23478) );
  NANDN U24518 ( .A(n23467), .B(n23466), .Z(n23471) );
  OR U24519 ( .A(n23469), .B(n23468), .Z(n23470) );
  AND U24520 ( .A(n23471), .B(n23470), .Z(n23477) );
  XOR U24521 ( .A(n23478), .B(n23477), .Z(n23480) );
  XOR U24522 ( .A(n23479), .B(n23480), .Z(n23493) );
  XNOR U24523 ( .A(n23493), .B(sreg[2034]), .Z(n23495) );
  NANDN U24524 ( .A(n23472), .B(sreg[2033]), .Z(n23476) );
  NAND U24525 ( .A(n23474), .B(n23473), .Z(n23475) );
  NAND U24526 ( .A(n23476), .B(n23475), .Z(n23494) );
  XOR U24527 ( .A(n23495), .B(n23494), .Z(c[2034]) );
  NANDN U24528 ( .A(n23478), .B(n23477), .Z(n23482) );
  OR U24529 ( .A(n23480), .B(n23479), .Z(n23481) );
  AND U24530 ( .A(n23482), .B(n23481), .Z(n23500) );
  XOR U24531 ( .A(a[1013]), .B(n2320), .Z(n23504) );
  AND U24532 ( .A(a[1011]), .B(b[3]), .Z(n23508) );
  AND U24533 ( .A(a[1015]), .B(b[0]), .Z(n23484) );
  XNOR U24534 ( .A(n23484), .B(n2175), .Z(n23486) );
  NANDN U24535 ( .A(b[0]), .B(a[1014]), .Z(n23485) );
  NAND U24536 ( .A(n23486), .B(n23485), .Z(n23509) );
  XOR U24537 ( .A(n23508), .B(n23509), .Z(n23511) );
  XOR U24538 ( .A(n23510), .B(n23511), .Z(n23499) );
  NANDN U24539 ( .A(n23488), .B(n23487), .Z(n23492) );
  OR U24540 ( .A(n23490), .B(n23489), .Z(n23491) );
  AND U24541 ( .A(n23492), .B(n23491), .Z(n23498) );
  XOR U24542 ( .A(n23499), .B(n23498), .Z(n23501) );
  XOR U24543 ( .A(n23500), .B(n23501), .Z(n23514) );
  XNOR U24544 ( .A(n23514), .B(sreg[2035]), .Z(n23516) );
  NANDN U24545 ( .A(n23493), .B(sreg[2034]), .Z(n23497) );
  NAND U24546 ( .A(n23495), .B(n23494), .Z(n23496) );
  NAND U24547 ( .A(n23497), .B(n23496), .Z(n23515) );
  XOR U24548 ( .A(n23516), .B(n23515), .Z(c[2035]) );
  NANDN U24549 ( .A(n23499), .B(n23498), .Z(n23503) );
  OR U24550 ( .A(n23501), .B(n23500), .Z(n23502) );
  AND U24551 ( .A(n23503), .B(n23502), .Z(n23521) );
  XOR U24552 ( .A(a[1014]), .B(n2321), .Z(n23525) );
  AND U24553 ( .A(a[1016]), .B(b[0]), .Z(n23505) );
  XNOR U24554 ( .A(n23505), .B(n2175), .Z(n23507) );
  NANDN U24555 ( .A(b[0]), .B(a[1015]), .Z(n23506) );
  NAND U24556 ( .A(n23507), .B(n23506), .Z(n23530) );
  AND U24557 ( .A(a[1012]), .B(b[3]), .Z(n23529) );
  XOR U24558 ( .A(n23530), .B(n23529), .Z(n23532) );
  XOR U24559 ( .A(n23531), .B(n23532), .Z(n23520) );
  NANDN U24560 ( .A(n23509), .B(n23508), .Z(n23513) );
  OR U24561 ( .A(n23511), .B(n23510), .Z(n23512) );
  AND U24562 ( .A(n23513), .B(n23512), .Z(n23519) );
  XOR U24563 ( .A(n23520), .B(n23519), .Z(n23522) );
  XOR U24564 ( .A(n23521), .B(n23522), .Z(n23535) );
  XNOR U24565 ( .A(n23535), .B(sreg[2036]), .Z(n23537) );
  NANDN U24566 ( .A(n23514), .B(sreg[2035]), .Z(n23518) );
  NAND U24567 ( .A(n23516), .B(n23515), .Z(n23517) );
  NAND U24568 ( .A(n23518), .B(n23517), .Z(n23536) );
  XOR U24569 ( .A(n23537), .B(n23536), .Z(c[2036]) );
  NANDN U24570 ( .A(n23520), .B(n23519), .Z(n23524) );
  OR U24571 ( .A(n23522), .B(n23521), .Z(n23523) );
  AND U24572 ( .A(n23524), .B(n23523), .Z(n23542) );
  XOR U24573 ( .A(a[1015]), .B(n2321), .Z(n23546) );
  AND U24574 ( .A(a[1017]), .B(b[0]), .Z(n23526) );
  XNOR U24575 ( .A(n23526), .B(n2175), .Z(n23528) );
  NANDN U24576 ( .A(b[0]), .B(a[1016]), .Z(n23527) );
  NAND U24577 ( .A(n23528), .B(n23527), .Z(n23551) );
  AND U24578 ( .A(a[1013]), .B(b[3]), .Z(n23550) );
  XOR U24579 ( .A(n23551), .B(n23550), .Z(n23553) );
  XOR U24580 ( .A(n23552), .B(n23553), .Z(n23541) );
  NANDN U24581 ( .A(n23530), .B(n23529), .Z(n23534) );
  OR U24582 ( .A(n23532), .B(n23531), .Z(n23533) );
  AND U24583 ( .A(n23534), .B(n23533), .Z(n23540) );
  XOR U24584 ( .A(n23541), .B(n23540), .Z(n23543) );
  XOR U24585 ( .A(n23542), .B(n23543), .Z(n23556) );
  XNOR U24586 ( .A(n23556), .B(sreg[2037]), .Z(n23558) );
  NANDN U24587 ( .A(n23535), .B(sreg[2036]), .Z(n23539) );
  NAND U24588 ( .A(n23537), .B(n23536), .Z(n23538) );
  NAND U24589 ( .A(n23539), .B(n23538), .Z(n23557) );
  XOR U24590 ( .A(n23558), .B(n23557), .Z(c[2037]) );
  NANDN U24591 ( .A(n23541), .B(n23540), .Z(n23545) );
  OR U24592 ( .A(n23543), .B(n23542), .Z(n23544) );
  AND U24593 ( .A(n23545), .B(n23544), .Z(n23563) );
  XOR U24594 ( .A(a[1016]), .B(n2321), .Z(n23567) );
  AND U24595 ( .A(a[1018]), .B(b[0]), .Z(n23547) );
  XNOR U24596 ( .A(n23547), .B(n2175), .Z(n23549) );
  NANDN U24597 ( .A(b[0]), .B(a[1017]), .Z(n23548) );
  NAND U24598 ( .A(n23549), .B(n23548), .Z(n23572) );
  AND U24599 ( .A(a[1014]), .B(b[3]), .Z(n23571) );
  XOR U24600 ( .A(n23572), .B(n23571), .Z(n23574) );
  XOR U24601 ( .A(n23573), .B(n23574), .Z(n23562) );
  NANDN U24602 ( .A(n23551), .B(n23550), .Z(n23555) );
  OR U24603 ( .A(n23553), .B(n23552), .Z(n23554) );
  AND U24604 ( .A(n23555), .B(n23554), .Z(n23561) );
  XOR U24605 ( .A(n23562), .B(n23561), .Z(n23564) );
  XOR U24606 ( .A(n23563), .B(n23564), .Z(n23577) );
  XNOR U24607 ( .A(n23577), .B(sreg[2038]), .Z(n23579) );
  NANDN U24608 ( .A(n23556), .B(sreg[2037]), .Z(n23560) );
  NAND U24609 ( .A(n23558), .B(n23557), .Z(n23559) );
  NAND U24610 ( .A(n23560), .B(n23559), .Z(n23578) );
  XOR U24611 ( .A(n23579), .B(n23578), .Z(c[2038]) );
  NANDN U24612 ( .A(n23562), .B(n23561), .Z(n23566) );
  OR U24613 ( .A(n23564), .B(n23563), .Z(n23565) );
  AND U24614 ( .A(n23566), .B(n23565), .Z(n23585) );
  XOR U24615 ( .A(a[1017]), .B(n2321), .Z(n23586) );
  AND U24616 ( .A(b[0]), .B(a[1019]), .Z(n23568) );
  XOR U24617 ( .A(b[1]), .B(n23568), .Z(n23570) );
  NANDN U24618 ( .A(b[0]), .B(a[1018]), .Z(n23569) );
  AND U24619 ( .A(n23570), .B(n23569), .Z(n23591) );
  AND U24620 ( .A(a[1015]), .B(b[3]), .Z(n23592) );
  XOR U24621 ( .A(n23591), .B(n23592), .Z(n23593) );
  XNOR U24622 ( .A(n23594), .B(n23593), .Z(n23582) );
  NANDN U24623 ( .A(n23572), .B(n23571), .Z(n23576) );
  OR U24624 ( .A(n23574), .B(n23573), .Z(n23575) );
  AND U24625 ( .A(n23576), .B(n23575), .Z(n23583) );
  XNOR U24626 ( .A(n23582), .B(n23583), .Z(n23584) );
  XNOR U24627 ( .A(n23585), .B(n23584), .Z(n23597) );
  XNOR U24628 ( .A(n23597), .B(sreg[2039]), .Z(n23599) );
  NANDN U24629 ( .A(n23577), .B(sreg[2038]), .Z(n23581) );
  NAND U24630 ( .A(n23579), .B(n23578), .Z(n23580) );
  NAND U24631 ( .A(n23581), .B(n23580), .Z(n23598) );
  XOR U24632 ( .A(n23599), .B(n23598), .Z(c[2039]) );
  XOR U24633 ( .A(a[1018]), .B(n2321), .Z(n23604) );
  AND U24634 ( .A(b[0]), .B(a[1020]), .Z(n23587) );
  XOR U24635 ( .A(b[1]), .B(n23587), .Z(n23590) );
  NAND U24636 ( .A(n23588), .B(a[1019]), .Z(n23589) );
  AND U24637 ( .A(n23590), .B(n23589), .Z(n23608) );
  AND U24638 ( .A(a[1016]), .B(b[3]), .Z(n23609) );
  XOR U24639 ( .A(n23608), .B(n23609), .Z(n23610) );
  XNOR U24640 ( .A(n23611), .B(n23610), .Z(n23600) );
  NAND U24641 ( .A(n23592), .B(n23591), .Z(n23596) );
  NANDN U24642 ( .A(n23594), .B(n23593), .Z(n23595) );
  AND U24643 ( .A(n23596), .B(n23595), .Z(n23601) );
  XNOR U24644 ( .A(n23600), .B(n23601), .Z(n23602) );
  XNOR U24645 ( .A(n23603), .B(n23602), .Z(n23614) );
  XNOR U24646 ( .A(n23614), .B(sreg[2040]), .Z(n23616) );
  XOR U24647 ( .A(n23616), .B(n23615), .Z(c[2040]) );
  XOR U24648 ( .A(a[1019]), .B(n2321), .Z(n23623) );
  AND U24649 ( .A(a[1021]), .B(b[0]), .Z(n23605) );
  XNOR U24650 ( .A(n23605), .B(n2175), .Z(n23607) );
  NANDN U24651 ( .A(b[0]), .B(a[1020]), .Z(n23606) );
  NAND U24652 ( .A(n23607), .B(n23606), .Z(n23628) );
  AND U24653 ( .A(a[1017]), .B(b[3]), .Z(n23627) );
  XOR U24654 ( .A(n23628), .B(n23627), .Z(n23630) );
  XOR U24655 ( .A(n23629), .B(n23630), .Z(n23618) );
  NAND U24656 ( .A(n23609), .B(n23608), .Z(n23613) );
  NANDN U24657 ( .A(n23611), .B(n23610), .Z(n23612) );
  AND U24658 ( .A(n23613), .B(n23612), .Z(n23617) );
  XOR U24659 ( .A(n23618), .B(n23617), .Z(n23620) );
  XOR U24660 ( .A(n23619), .B(n23620), .Z(n23633) );
  XNOR U24661 ( .A(n23633), .B(sreg[2041]), .Z(n23635) );
  XOR U24662 ( .A(n23635), .B(n23634), .Z(c[2041]) );
  NANDN U24663 ( .A(n23618), .B(n23617), .Z(n23622) );
  OR U24664 ( .A(n23620), .B(n23619), .Z(n23621) );
  AND U24665 ( .A(n23622), .B(n23621), .Z(n23640) );
  XNOR U24666 ( .A(b[3]), .B(a[1020]), .Z(n23644) );
  AND U24667 ( .A(a[1022]), .B(b[0]), .Z(n23624) );
  XNOR U24668 ( .A(n23624), .B(n2175), .Z(n23626) );
  NANDN U24669 ( .A(b[0]), .B(a[1021]), .Z(n23625) );
  NAND U24670 ( .A(n23626), .B(n23625), .Z(n23651) );
  AND U24671 ( .A(a[1018]), .B(b[3]), .Z(n23650) );
  XOR U24672 ( .A(n23651), .B(n23650), .Z(n23653) );
  XOR U24673 ( .A(n23652), .B(n23653), .Z(n23639) );
  NANDN U24674 ( .A(n23628), .B(n23627), .Z(n23632) );
  OR U24675 ( .A(n23630), .B(n23629), .Z(n23631) );
  AND U24676 ( .A(n23632), .B(n23631), .Z(n23638) );
  XOR U24677 ( .A(n23639), .B(n23638), .Z(n23641) );
  XOR U24678 ( .A(n23640), .B(n23641), .Z(n23656) );
  XNOR U24679 ( .A(n23656), .B(sreg[2042]), .Z(n23658) );
  NANDN U24680 ( .A(n23633), .B(sreg[2041]), .Z(n23637) );
  NAND U24681 ( .A(n23635), .B(n23634), .Z(n23636) );
  NAND U24682 ( .A(n23637), .B(n23636), .Z(n23657) );
  XOR U24683 ( .A(n23658), .B(n23657), .Z(c[2042]) );
  NANDN U24684 ( .A(n23639), .B(n23638), .Z(n23643) );
  OR U24685 ( .A(n23641), .B(n23640), .Z(n23642) );
  AND U24686 ( .A(n23643), .B(n23642), .Z(n23664) );
  OR U24687 ( .A(n23644), .B(n2172), .Z(n23646) );
  XNOR U24688 ( .A(b[3]), .B(a[1021]), .Z(n23667) );
  OR U24689 ( .A(n23667), .B(n2171), .Z(n23645) );
  NAND U24690 ( .A(n23646), .B(n23645), .Z(n23672) );
  AND U24691 ( .A(a[1023]), .B(b[0]), .Z(n23647) );
  XNOR U24692 ( .A(n23647), .B(n2175), .Z(n23649) );
  NANDN U24693 ( .A(b[0]), .B(a[1022]), .Z(n23648) );
  NAND U24694 ( .A(n23649), .B(n23648), .Z(n23671) );
  AND U24695 ( .A(a[1019]), .B(b[3]), .Z(n23670) );
  XOR U24696 ( .A(n23671), .B(n23670), .Z(n23673) );
  XNOR U24697 ( .A(n23672), .B(n23673), .Z(n23661) );
  NANDN U24698 ( .A(n23651), .B(n23650), .Z(n23655) );
  OR U24699 ( .A(n23653), .B(n23652), .Z(n23654) );
  AND U24700 ( .A(n23655), .B(n23654), .Z(n23662) );
  XNOR U24701 ( .A(n23661), .B(n23662), .Z(n23663) );
  XNOR U24702 ( .A(n23664), .B(n23663), .Z(n23676) );
  XNOR U24703 ( .A(n23676), .B(sreg[2043]), .Z(n23678) );
  NANDN U24704 ( .A(n23656), .B(sreg[2042]), .Z(n23660) );
  NAND U24705 ( .A(n23658), .B(n23657), .Z(n23659) );
  NAND U24706 ( .A(n23660), .B(n23659), .Z(n23677) );
  XOR U24707 ( .A(n23678), .B(n23677), .Z(c[2043]) );
  NANDN U24708 ( .A(a[1023]), .B(b[1]), .Z(n23666) );
  NAND U24709 ( .A(b[1]), .B(b[0]), .Z(n23665) );
  AND U24710 ( .A(n23666), .B(n23665), .Z(n23689) );
  OR U24711 ( .A(n23667), .B(n2172), .Z(n23669) );
  XNOR U24712 ( .A(b[3]), .B(a[1022]), .Z(n23691) );
  OR U24713 ( .A(n23691), .B(n2171), .Z(n23668) );
  AND U24714 ( .A(n23669), .B(n23668), .Z(n23687) );
  AND U24715 ( .A(a[1020]), .B(b[3]), .Z(n23688) );
  XNOR U24716 ( .A(n23687), .B(n23688), .Z(n23690) );
  XNOR U24717 ( .A(n23689), .B(n23690), .Z(n23682) );
  NANDN U24718 ( .A(n23671), .B(n23670), .Z(n23675) );
  NANDN U24719 ( .A(n23673), .B(n23672), .Z(n23674) );
  AND U24720 ( .A(n23675), .B(n23674), .Z(n23681) );
  XOR U24721 ( .A(n23682), .B(n23681), .Z(n23684) );
  XOR U24722 ( .A(n23683), .B(n23684), .Z(n23680) );
  XOR U24723 ( .A(n23680), .B(n23679), .Z(c[2044]) );
  AND U24724 ( .A(n23680), .B(n23679), .Z(n23709) );
  NANDN U24725 ( .A(n23682), .B(n23681), .Z(n23686) );
  NANDN U24726 ( .A(n23684), .B(n23683), .Z(n23685) );
  NAND U24727 ( .A(n23686), .B(n23685), .Z(n23696) );
  OR U24728 ( .A(n23691), .B(n2172), .Z(n23693) );
  XNOR U24729 ( .A(a[1023]), .B(b[3]), .Z(n23705) );
  OR U24730 ( .A(n23705), .B(n2171), .Z(n23692) );
  AND U24731 ( .A(n23693), .B(n23692), .Z(n23700) );
  AND U24732 ( .A(a[1021]), .B(b[3]), .Z(n23716) );
  XNOR U24733 ( .A(b[1]), .B(n23716), .Z(n23701) );
  XNOR U24734 ( .A(n23700), .B(n23701), .Z(n23694) );
  XNOR U24735 ( .A(n23695), .B(n23694), .Z(n23697) );
  XOR U24736 ( .A(n23696), .B(n23697), .Z(n23708) );
  XOR U24737 ( .A(n23709), .B(n23708), .Z(c[2045]) );
  NAND U24738 ( .A(n23695), .B(n23694), .Z(n23699) );
  NANDN U24739 ( .A(n23697), .B(n23696), .Z(n23698) );
  AND U24740 ( .A(n23699), .B(n23698), .Z(n23715) );
  NAND U24741 ( .A(b[1]), .B(n23716), .Z(n23703) );
  NANDN U24742 ( .A(n23701), .B(n23700), .Z(n23702) );
  AND U24743 ( .A(n23703), .B(n23702), .Z(n23714) );
  XOR U24744 ( .A(n23715), .B(n23714), .Z(n23711) );
  XNOR U24745 ( .A(b[2]), .B(n2175), .Z(n23704) );
  NANDN U24746 ( .A(n2321), .B(n23704), .Z(n23707) );
  OR U24747 ( .A(n23705), .B(n2172), .Z(n23706) );
  NAND U24748 ( .A(n23707), .B(n23706), .Z(n23719) );
  AND U24749 ( .A(a[1022]), .B(b[3]), .Z(n23717) );
  XOR U24750 ( .A(n23716), .B(n23717), .Z(n23718) );
  XNOR U24751 ( .A(n23719), .B(n23718), .Z(n23713) );
  NAND U24752 ( .A(n23709), .B(n23708), .Z(n23712) );
  XOR U24753 ( .A(n23713), .B(n23712), .Z(n23710) );
  XNOR U24754 ( .A(n23711), .B(n23710), .Z(c[2046]) );
endmodule

