
module mult_N128_CC2 ( clk, rst, a, b, c );
  input [127:0] a;
  input [63:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305;
  wire   [255:0] sreg;

  DFF \sreg_reg[191]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U67 ( .A(n5614), .B(n5613), .Z(n5538) );
  NAND U68 ( .A(n38260), .B(n38261), .Z(n1) );
  NAND U69 ( .A(n38259), .B(n38275), .Z(n2) );
  NAND U70 ( .A(n1), .B(n2), .Z(n38286) );
  XNOR U71 ( .A(n11349), .B(n11348), .Z(n11457) );
  XNOR U72 ( .A(n13141), .B(n13140), .Z(n13249) );
  XNOR U73 ( .A(n14568), .B(n14567), .Z(n14676) );
  XNOR U74 ( .A(n15163), .B(n15162), .Z(n15271) );
  XNOR U75 ( .A(n15772), .B(n15771), .Z(n15880) );
  XNOR U76 ( .A(n16032), .B(n16031), .Z(n16140) );
  XNOR U77 ( .A(n20436), .B(n20435), .Z(n20544) );
  XNOR U78 ( .A(n20745), .B(n20744), .Z(n20853) );
  XNOR U79 ( .A(n21622), .B(n21621), .Z(n21730) );
  XNOR U80 ( .A(n22726), .B(n22725), .Z(n22864) );
  XNOR U81 ( .A(n25340), .B(n25339), .Z(n25499) );
  XNOR U82 ( .A(n5602), .B(n5601), .Z(n5539) );
  NAND U83 ( .A(n27668), .B(n27667), .Z(n3) );
  NAND U84 ( .A(n27666), .B(n27665), .Z(n4) );
  AND U85 ( .A(n3), .B(n4), .Z(n28141) );
  NAND U86 ( .A(n37179), .B(n37077), .Z(n5) );
  NANDN U87 ( .A(n37079), .B(n37078), .Z(n6) );
  AND U88 ( .A(n5), .B(n6), .Z(n37193) );
  NAND U89 ( .A(n37870), .B(n37869), .Z(n7) );
  NANDN U90 ( .A(n37868), .B(n37867), .Z(n8) );
  NAND U91 ( .A(n7), .B(n8), .Z(n37890) );
  NAND U92 ( .A(n38273), .B(n38274), .Z(n9) );
  NANDN U93 ( .A(n38275), .B(n38276), .Z(n10) );
  AND U94 ( .A(n9), .B(n10), .Z(n38299) );
  XOR U95 ( .A(n11080), .B(n11079), .Z(n11144) );
  XOR U96 ( .A(n12782), .B(n12781), .Z(n12894) );
  XOR U97 ( .A(n14293), .B(n14292), .Z(n14357) );
  XOR U98 ( .A(n14889), .B(n14888), .Z(n14953) );
  XOR U99 ( .A(n15425), .B(n15424), .Z(n15537) );
  XOR U100 ( .A(n15766), .B(n15765), .Z(n15788) );
  XOR U101 ( .A(n20077), .B(n20076), .Z(n20189) );
  XOR U102 ( .A(n20430), .B(n20429), .Z(n20494) );
  XOR U103 ( .A(n21299), .B(n21298), .Z(n21321) );
  XOR U104 ( .A(n22493), .B(n22492), .Z(n22515) );
  XOR U105 ( .A(n25128), .B(n25127), .Z(n25192) );
  XOR U106 ( .A(n10021), .B(n10020), .Z(n9816) );
  XNOR U107 ( .A(n11319), .B(n11318), .Z(n11458) );
  XNOR U108 ( .A(n13042), .B(n13041), .Z(n13250) );
  XNOR U109 ( .A(n14463), .B(n14462), .Z(n14677) );
  XNOR U110 ( .A(n15112), .B(n15111), .Z(n15272) );
  XNOR U111 ( .A(n15721), .B(n15720), .Z(n15881) );
  XNOR U112 ( .A(n15927), .B(n15926), .Z(n16141) );
  XNOR U113 ( .A(n20385), .B(n20384), .Z(n20545) );
  XNOR U114 ( .A(n20715), .B(n20714), .Z(n20854) );
  XNOR U115 ( .A(n21571), .B(n21570), .Z(n21731) );
  XNOR U116 ( .A(n22756), .B(n22755), .Z(n22865) );
  XNOR U117 ( .A(n25391), .B(n25390), .Z(n25500) );
  NAND U118 ( .A(n6170), .B(n6169), .Z(n11) );
  NANDN U119 ( .A(n6168), .B(n6167), .Z(n12) );
  NAND U120 ( .A(n11), .B(n12), .Z(n6448) );
  NAND U121 ( .A(n28833), .B(b[1]), .Z(n13) );
  XOR U122 ( .A(n28833), .B(b[1]), .Z(n14) );
  NANDN U123 ( .A(n29147), .B(n14), .Z(n15) );
  NAND U124 ( .A(n13), .B(n15), .Z(n29187) );
  XNOR U125 ( .A(n29448), .B(n29447), .Z(n29449) );
  NAND U126 ( .A(n27784), .B(n27785), .Z(n16) );
  NANDN U127 ( .A(n27787), .B(n27786), .Z(n17) );
  AND U128 ( .A(n16), .B(n17), .Z(n28132) );
  NAND U129 ( .A(n30116), .B(n30117), .Z(n18) );
  XOR U130 ( .A(n30116), .B(n30117), .Z(n19) );
  NANDN U131 ( .A(n30115), .B(n19), .Z(n20) );
  NAND U132 ( .A(n18), .B(n20), .Z(n30172) );
  NAND U133 ( .A(n36185), .B(n36114), .Z(n21) );
  NANDN U134 ( .A(n36116), .B(n36115), .Z(n22) );
  AND U135 ( .A(n21), .B(n22), .Z(n36155) );
  NAND U136 ( .A(n4543), .B(n4542), .Z(n23) );
  NAND U137 ( .A(n4541), .B(n4540), .Z(n24) );
  AND U138 ( .A(n23), .B(n24), .Z(n4796) );
  NAND U139 ( .A(n5447), .B(n5446), .Z(n25) );
  NANDN U140 ( .A(n5445), .B(n5444), .Z(n26) );
  AND U141 ( .A(n25), .B(n26), .Z(n5860) );
  NAND U142 ( .A(n8062), .B(n8061), .Z(n27) );
  NANDN U143 ( .A(n8060), .B(n8059), .Z(n28) );
  AND U144 ( .A(n27), .B(n28), .Z(n8335) );
  NAND U145 ( .A(n9378), .B(n9379), .Z(n29) );
  NANDN U146 ( .A(n9381), .B(n9380), .Z(n30) );
  AND U147 ( .A(n29), .B(n30), .Z(n9490) );
  NAND U148 ( .A(n27661), .B(n27662), .Z(n31) );
  NANDN U149 ( .A(n27664), .B(n27663), .Z(n32) );
  AND U150 ( .A(n31), .B(n32), .Z(n28165) );
  NAND U151 ( .A(n31376), .B(n31375), .Z(n33) );
  NANDN U152 ( .A(n31374), .B(n31373), .Z(n34) );
  AND U153 ( .A(n33), .B(n34), .Z(n31697) );
  NAND U154 ( .A(n37196), .B(n37197), .Z(n35) );
  NANDN U155 ( .A(n37199), .B(n37198), .Z(n36) );
  AND U156 ( .A(n35), .B(n36), .Z(n37253) );
  NAND U157 ( .A(n37337), .B(n37300), .Z(n37) );
  NANDN U158 ( .A(n37302), .B(n37301), .Z(n38) );
  AND U159 ( .A(n37), .B(n38), .Z(n37387) );
  NAND U160 ( .A(n37830), .B(n37763), .Z(n39) );
  NANDN U161 ( .A(n37765), .B(n37764), .Z(n40) );
  NAND U162 ( .A(n39), .B(n40), .Z(n37871) );
  NAND U163 ( .A(n29343), .B(n29342), .Z(n41) );
  NANDN U164 ( .A(n29341), .B(n29340), .Z(n42) );
  AND U165 ( .A(n41), .B(n42), .Z(n29620) );
  NAND U166 ( .A(n35395), .B(n35396), .Z(n43) );
  NANDN U167 ( .A(n35398), .B(n35397), .Z(n44) );
  AND U168 ( .A(n43), .B(n44), .Z(n35693) );
  NAND U169 ( .A(n37889), .B(n37890), .Z(n45) );
  NANDN U170 ( .A(n37892), .B(n37891), .Z(n46) );
  AND U171 ( .A(n45), .B(n46), .Z(n37944) );
  NAND U172 ( .A(n261), .B(n262), .Z(n47) );
  NANDN U173 ( .A(n264), .B(n263), .Z(n48) );
  AND U174 ( .A(n47), .B(n48), .Z(n297) );
  NAND U175 ( .A(sreg[105]), .B(n4225), .Z(n49) );
  XOR U176 ( .A(sreg[105]), .B(n4225), .Z(n50) );
  NANDN U177 ( .A(n4224), .B(n50), .Z(n51) );
  NAND U178 ( .A(n49), .B(n51), .Z(n4604) );
  XOR U179 ( .A(n3678), .B(sreg[102]), .Z(n52) );
  NANDN U180 ( .A(n3679), .B(n52), .Z(n53) );
  NAND U181 ( .A(n3678), .B(sreg[102]), .Z(n54) );
  AND U182 ( .A(n53), .B(n54), .Z(n4035) );
  NAND U183 ( .A(n38290), .B(n38291), .Z(n55) );
  NANDN U184 ( .A(n38293), .B(n38292), .Z(n56) );
  NAND U185 ( .A(n55), .B(n56), .Z(n38305) );
  NANDN U186 ( .A(b[0]), .B(a[127]), .Z(n57) );
  NAND U187 ( .A(b[1]), .B(n57), .Z(n28574) );
  NAND U188 ( .A(b[0]), .B(a[41]), .Z(n58) );
  XNOR U189 ( .A(b[1]), .B(n58), .Z(n59) );
  NANDN U190 ( .A(b[0]), .B(a[40]), .Z(n60) );
  AND U191 ( .A(n59), .B(n60), .Z(n4346) );
  XOR U192 ( .A(n5388), .B(n5387), .Z(n5362) );
  XOR U193 ( .A(n5400), .B(n5399), .Z(n5356) );
  NAND U194 ( .A(n9367), .B(n9366), .Z(n61) );
  NANDN U195 ( .A(n9365), .B(n9364), .Z(n62) );
  AND U196 ( .A(n61), .B(n62), .Z(n9514) );
  NAND U197 ( .A(n9812), .B(n9811), .Z(n63) );
  NANDN U198 ( .A(n9810), .B(n9809), .Z(n64) );
  AND U199 ( .A(n63), .B(n64), .Z(n10293) );
  NAND U200 ( .A(n11457), .B(n11458), .Z(n65) );
  NANDN U201 ( .A(n11460), .B(n11459), .Z(n66) );
  AND U202 ( .A(n65), .B(n66), .Z(n11568) );
  NAND U203 ( .A(n13249), .B(n13250), .Z(n67) );
  NANDN U204 ( .A(n13252), .B(n13251), .Z(n68) );
  AND U205 ( .A(n67), .B(n68), .Z(n13318) );
  NAND U206 ( .A(n14676), .B(n14677), .Z(n69) );
  NANDN U207 ( .A(n14679), .B(n14678), .Z(n70) );
  AND U208 ( .A(n69), .B(n70), .Z(n14781) );
  NAND U209 ( .A(n15271), .B(n15272), .Z(n71) );
  NANDN U210 ( .A(n15274), .B(n15273), .Z(n72) );
  AND U211 ( .A(n71), .B(n72), .Z(n15365) );
  NAND U212 ( .A(n15880), .B(n15881), .Z(n73) );
  NANDN U213 ( .A(n15883), .B(n15882), .Z(n74) );
  AND U214 ( .A(n73), .B(n74), .Z(n15918) );
  NAND U215 ( .A(n16140), .B(n16141), .Z(n75) );
  NANDN U216 ( .A(n16143), .B(n16142), .Z(n76) );
  AND U217 ( .A(n75), .B(n76), .Z(n16240) );
  NAND U218 ( .A(n20544), .B(n20545), .Z(n77) );
  NANDN U219 ( .A(n20547), .B(n20546), .Z(n78) );
  AND U220 ( .A(n77), .B(n78), .Z(n20631) );
  NAND U221 ( .A(n20853), .B(n20854), .Z(n79) );
  NANDN U222 ( .A(n20856), .B(n20855), .Z(n80) );
  AND U223 ( .A(n79), .B(n80), .Z(n20922) );
  NAND U224 ( .A(n21730), .B(n21731), .Z(n81) );
  NANDN U225 ( .A(n21733), .B(n21732), .Z(n82) );
  AND U226 ( .A(n81), .B(n82), .Z(n21775) );
  NAND U227 ( .A(n22864), .B(n22865), .Z(n83) );
  NANDN U228 ( .A(n22867), .B(n22866), .Z(n84) );
  AND U229 ( .A(n83), .B(n84), .Z(n22957) );
  NAND U230 ( .A(n25499), .B(n25500), .Z(n85) );
  NANDN U231 ( .A(n25502), .B(n25501), .Z(n86) );
  AND U232 ( .A(n85), .B(n86), .Z(n25610) );
  NAND U233 ( .A(n29374), .B(n29373), .Z(n87) );
  NANDN U234 ( .A(n29372), .B(n29371), .Z(n88) );
  AND U235 ( .A(n87), .B(n88), .Z(n29820) );
  NAND U236 ( .A(n2499), .B(n2498), .Z(n89) );
  NANDN U237 ( .A(n2497), .B(n2496), .Z(n90) );
  AND U238 ( .A(n89), .B(n90), .Z(n2584) );
  XOR U239 ( .A(n3901), .B(n3900), .Z(n3927) );
  NAND U240 ( .A(n4509), .B(n4508), .Z(n91) );
  NANDN U241 ( .A(n4507), .B(n4506), .Z(n92) );
  NAND U242 ( .A(n91), .B(n92), .Z(n4636) );
  NAND U243 ( .A(n4843), .B(n4842), .Z(n93) );
  NANDN U244 ( .A(n4841), .B(n4840), .Z(n94) );
  NAND U245 ( .A(n93), .B(n94), .Z(n5050) );
  XNOR U246 ( .A(n5266), .B(n5265), .Z(n5415) );
  NAND U247 ( .A(n5188), .B(n5189), .Z(n95) );
  NANDN U248 ( .A(n5191), .B(n5190), .Z(n96) );
  NAND U249 ( .A(n95), .B(n96), .Z(n5422) );
  NAND U250 ( .A(n6451), .B(n6450), .Z(n97) );
  NANDN U251 ( .A(n6449), .B(n6448), .Z(n98) );
  NAND U252 ( .A(n97), .B(n98), .Z(n6650) );
  NAND U253 ( .A(n27783), .B(n27782), .Z(n99) );
  NANDN U254 ( .A(n27781), .B(n27780), .Z(n100) );
  AND U255 ( .A(n99), .B(n100), .Z(n28151) );
  NAND U256 ( .A(n31345), .B(n31346), .Z(n101) );
  NANDN U257 ( .A(n31348), .B(n31347), .Z(n102) );
  AND U258 ( .A(n101), .B(n102), .Z(n31648) );
  NAND U259 ( .A(n33775), .B(n33776), .Z(n103) );
  NANDN U260 ( .A(n33778), .B(n33777), .Z(n104) );
  NAND U261 ( .A(n103), .B(n104), .Z(n34094) );
  NAND U262 ( .A(n34266), .B(n34031), .Z(n105) );
  NANDN U263 ( .A(n34033), .B(n34032), .Z(n106) );
  AND U264 ( .A(n105), .B(n106), .Z(n34162) );
  NAND U265 ( .A(n34256), .B(n34255), .Z(n107) );
  NANDN U266 ( .A(n34254), .B(n34253), .Z(n108) );
  NAND U267 ( .A(n107), .B(n108), .Z(n34481) );
  NAND U268 ( .A(n35340), .B(n35341), .Z(n109) );
  NANDN U269 ( .A(n35342), .B(n35343), .Z(n110) );
  AND U270 ( .A(n109), .B(n110), .Z(n35430) );
  NAND U271 ( .A(n1723), .B(n1722), .Z(n111) );
  NANDN U272 ( .A(n1721), .B(n1720), .Z(n112) );
  AND U273 ( .A(n111), .B(n112), .Z(n1878) );
  NAND U274 ( .A(n2106), .B(n2105), .Z(n113) );
  NANDN U275 ( .A(n2104), .B(n2103), .Z(n114) );
  AND U276 ( .A(n113), .B(n114), .Z(n2226) );
  NAND U277 ( .A(n4881), .B(n4880), .Z(n115) );
  NANDN U278 ( .A(n4879), .B(n4878), .Z(n116) );
  NAND U279 ( .A(n115), .B(n116), .Z(n5047) );
  NAND U280 ( .A(n5538), .B(n5539), .Z(n117) );
  NANDN U281 ( .A(n5541), .B(n5540), .Z(n118) );
  NAND U282 ( .A(n117), .B(n118), .Z(n5857) );
  NAND U283 ( .A(n28796), .B(n28795), .Z(n119) );
  NAND U284 ( .A(n28793), .B(n28794), .Z(n120) );
  AND U285 ( .A(n119), .B(n120), .Z(n29318) );
  NAND U286 ( .A(n30139), .B(n30138), .Z(n121) );
  NANDN U287 ( .A(n30137), .B(n30136), .Z(n122) );
  NAND U288 ( .A(n121), .B(n122), .Z(n30407) );
  NAND U289 ( .A(n33085), .B(n33084), .Z(n123) );
  NAND U290 ( .A(n33082), .B(n33083), .Z(n124) );
  NAND U291 ( .A(n123), .B(n124), .Z(n33112) );
  NAND U292 ( .A(n33517), .B(n33516), .Z(n125) );
  NANDN U293 ( .A(n33515), .B(n33514), .Z(n126) );
  AND U294 ( .A(n125), .B(n126), .Z(n33698) );
  NAND U295 ( .A(n34933), .B(n34932), .Z(n127) );
  NANDN U296 ( .A(n34931), .B(n34930), .Z(n128) );
  NAND U297 ( .A(n127), .B(n128), .Z(n35082) );
  NAND U298 ( .A(n36031), .B(n36032), .Z(n129) );
  NANDN U299 ( .A(n36034), .B(n36033), .Z(n130) );
  AND U300 ( .A(n129), .B(n130), .Z(n36261) );
  NAND U301 ( .A(n36942), .B(n36855), .Z(n131) );
  NANDN U302 ( .A(n36857), .B(n36856), .Z(n132) );
  NAND U303 ( .A(n131), .B(n132), .Z(n37006) );
  NAND U304 ( .A(n36957), .B(n36956), .Z(n133) );
  NANDN U305 ( .A(n36955), .B(n36954), .Z(n134) );
  AND U306 ( .A(n133), .B(n134), .Z(n37040) );
  NAND U307 ( .A(n37348), .B(n37349), .Z(n135) );
  NANDN U308 ( .A(n37351), .B(n37350), .Z(n136) );
  NAND U309 ( .A(n135), .B(n136), .Z(n37481) );
  NAND U310 ( .A(n790), .B(n789), .Z(n137) );
  NANDN U311 ( .A(n788), .B(n787), .Z(n138) );
  NAND U312 ( .A(n137), .B(n138), .Z(n813) );
  NAND U313 ( .A(n1666), .B(n1665), .Z(n139) );
  NANDN U314 ( .A(n1664), .B(n1663), .Z(n140) );
  AND U315 ( .A(n139), .B(n140), .Z(n1786) );
  NAND U316 ( .A(n5632), .B(n5631), .Z(n141) );
  NANDN U317 ( .A(n5630), .B(n5629), .Z(n142) );
  NAND U318 ( .A(n141), .B(n142), .Z(n5651) );
  NAND U319 ( .A(n8078), .B(n8077), .Z(n143) );
  NANDN U320 ( .A(n8076), .B(n8075), .Z(n144) );
  NAND U321 ( .A(n143), .B(n144), .Z(n8340) );
  NAND U322 ( .A(n8938), .B(n8939), .Z(n145) );
  NANDN U323 ( .A(n8941), .B(n8940), .Z(n146) );
  AND U324 ( .A(n145), .B(n146), .Z(n9207) );
  NAND U325 ( .A(n9374), .B(n9375), .Z(n147) );
  NANDN U326 ( .A(n9377), .B(n9376), .Z(n148) );
  AND U327 ( .A(n147), .B(n148), .Z(n9483) );
  NAND U328 ( .A(n10059), .B(n10060), .Z(n149) );
  NANDN U329 ( .A(n10062), .B(n10061), .Z(n150) );
  AND U330 ( .A(n149), .B(n150), .Z(n10628) );
  NAND U331 ( .A(n28162), .B(n28163), .Z(n151) );
  NANDN U332 ( .A(n28165), .B(n28164), .Z(n152) );
  AND U333 ( .A(n151), .B(n152), .Z(n28195) );
  NAND U334 ( .A(n31380), .B(n31379), .Z(n153) );
  NANDN U335 ( .A(n31378), .B(n31377), .Z(n154) );
  AND U336 ( .A(n153), .B(n154), .Z(n31477) );
  NAND U337 ( .A(n35526), .B(n35527), .Z(n155) );
  NANDN U338 ( .A(n35529), .B(n35528), .Z(n156) );
  NAND U339 ( .A(n155), .B(n156), .Z(n35545) );
  NAND U340 ( .A(n37217), .B(n37216), .Z(n157) );
  NAND U341 ( .A(n37215), .B(n37214), .Z(n158) );
  AND U342 ( .A(n157), .B(n158), .Z(n37310) );
  NAND U343 ( .A(n37250), .B(n37251), .Z(n159) );
  NANDN U344 ( .A(n37253), .B(n37252), .Z(n160) );
  NAND U345 ( .A(n159), .B(n160), .Z(n37324) );
  NAND U346 ( .A(n37831), .B(n37832), .Z(n161) );
  NANDN U347 ( .A(n37830), .B(n37829), .Z(n162) );
  AND U348 ( .A(n161), .B(n162), .Z(n37893) );
  NAND U349 ( .A(n37963), .B(n37962), .Z(n163) );
  NANDN U350 ( .A(n37961), .B(n37960), .Z(n164) );
  AND U351 ( .A(n163), .B(n164), .Z(n38008) );
  NAND U352 ( .A(n1341), .B(n1340), .Z(n165) );
  NAND U353 ( .A(n1338), .B(n1339), .Z(n166) );
  AND U354 ( .A(n165), .B(n166), .Z(n1525) );
  NAND U355 ( .A(n4623), .B(n4622), .Z(n167) );
  NAND U356 ( .A(n4620), .B(n4621), .Z(n168) );
  AND U357 ( .A(n167), .B(n168), .Z(n5006) );
  NAND U358 ( .A(n6826), .B(n6825), .Z(n169) );
  NANDN U359 ( .A(n6824), .B(n6823), .Z(n170) );
  AND U360 ( .A(n169), .B(n170), .Z(n7068) );
  XOR U361 ( .A(n17373), .B(n17371), .Z(n171) );
  NANDN U362 ( .A(n17372), .B(n171), .Z(n172) );
  NAND U363 ( .A(n17373), .B(n17371), .Z(n173) );
  AND U364 ( .A(n172), .B(n173), .Z(n17656) );
  NAND U365 ( .A(n29339), .B(n29338), .Z(n174) );
  NAND U366 ( .A(n29337), .B(n29336), .Z(n175) );
  AND U367 ( .A(n174), .B(n175), .Z(n29612) );
  NAND U368 ( .A(n35394), .B(n35393), .Z(n176) );
  NAND U369 ( .A(n35392), .B(n35391), .Z(n177) );
  AND U370 ( .A(n176), .B(n177), .Z(n35539) );
  NAND U371 ( .A(n37885), .B(n37886), .Z(n178) );
  NANDN U372 ( .A(n37888), .B(n37887), .Z(n179) );
  AND U373 ( .A(n178), .B(n179), .Z(n37937) );
  XOR U374 ( .A(n251), .B(n249), .Z(n180) );
  NANDN U375 ( .A(n250), .B(n180), .Z(n181) );
  NAND U376 ( .A(n251), .B(n249), .Z(n182) );
  AND U377 ( .A(n181), .B(n182), .Z(n264) );
  NAND U378 ( .A(sreg[99]), .B(n3172), .Z(n183) );
  XOR U379 ( .A(sreg[99]), .B(n3172), .Z(n184) );
  NANDN U380 ( .A(n3171), .B(n184), .Z(n185) );
  NAND U381 ( .A(n183), .B(n185), .Z(n3499) );
  XOR U382 ( .A(n2699), .B(sreg[96]), .Z(n186) );
  NANDN U383 ( .A(n2700), .B(n186), .Z(n187) );
  NAND U384 ( .A(n2699), .B(sreg[96]), .Z(n188) );
  AND U385 ( .A(n187), .B(n188), .Z(n2852) );
  NAND U386 ( .A(sreg[104]), .B(n4222), .Z(n189) );
  XOR U387 ( .A(sreg[104]), .B(n4222), .Z(n190) );
  NANDN U388 ( .A(n4221), .B(n190), .Z(n191) );
  NAND U389 ( .A(n189), .B(n191), .Z(n4225) );
  XOR U390 ( .A(n4808), .B(sreg[108]), .Z(n192) );
  NANDN U391 ( .A(n4809), .B(n192), .Z(n193) );
  NAND U392 ( .A(n4808), .B(sreg[108]), .Z(n194) );
  AND U393 ( .A(n193), .B(n194), .Z(n5011) );
  XNOR U394 ( .A(a[127]), .B(a[126]), .Z(n195) );
  XNOR U395 ( .A(n38296), .B(n195), .Z(n196) );
  AND U396 ( .A(n196), .B(b[63]), .Z(n197) );
  NANDN U397 ( .A(n38299), .B(n38300), .Z(n198) );
  NANDN U398 ( .A(n38297), .B(n38298), .Z(n199) );
  AND U399 ( .A(n198), .B(n199), .Z(n200) );
  NOR U400 ( .A(n38305), .B(n38304), .Z(n201) );
  NANDN U401 ( .A(n38301), .B(n38304), .Z(n202) );
  OR U402 ( .A(n201), .B(n38302), .Z(n203) );
  NAND U403 ( .A(n202), .B(n203), .Z(n204) );
  OR U404 ( .A(n38302), .B(n202), .Z(n205) );
  NANDN U405 ( .A(n38303), .B(n205), .Z(n206) );
  NAND U406 ( .A(n204), .B(n206), .Z(n207) );
  XNOR U407 ( .A(n197), .B(n200), .Z(n208) );
  XNOR U408 ( .A(n207), .B(n208), .Z(c[255]) );
  IV U409 ( .A(n9942), .Z(n209) );
  IV U410 ( .A(n30627), .Z(n210) );
  IV U411 ( .A(n37294), .Z(n211) );
  IV U412 ( .A(n37536), .Z(n212) );
  AND U413 ( .A(b[0]), .B(a[0]), .Z(n214) );
  XOR U414 ( .A(n214), .B(sreg[64]), .Z(c[64]) );
  AND U415 ( .A(b[0]), .B(a[1]), .Z(n221) );
  NAND U416 ( .A(a[0]), .B(b[1]), .Z(n213) );
  XOR U417 ( .A(n221), .B(n213), .Z(n215) );
  XNOR U418 ( .A(sreg[65]), .B(n215), .Z(n217) );
  AND U419 ( .A(n214), .B(sreg[64]), .Z(n216) );
  XOR U420 ( .A(n217), .B(n216), .Z(c[65]) );
  NANDN U421 ( .A(n215), .B(sreg[65]), .Z(n219) );
  NAND U422 ( .A(n217), .B(n216), .Z(n218) );
  AND U423 ( .A(n219), .B(n218), .Z(n239) );
  XNOR U424 ( .A(n239), .B(sreg[66]), .Z(n241) );
  NAND U425 ( .A(a[0]), .B(b[2]), .Z(n220) );
  XNOR U426 ( .A(b[1]), .B(n220), .Z(n223) );
  NANDN U427 ( .A(a[0]), .B(n221), .Z(n222) );
  NAND U428 ( .A(n223), .B(n222), .Z(n228) );
  NAND U429 ( .A(b[0]), .B(a[2]), .Z(n224) );
  XNOR U430 ( .A(b[1]), .B(n224), .Z(n226) );
  NANDN U431 ( .A(b[0]), .B(a[1]), .Z(n225) );
  NAND U432 ( .A(n226), .B(n225), .Z(n227) );
  XOR U433 ( .A(n228), .B(n227), .Z(n240) );
  XOR U434 ( .A(n241), .B(n240), .Z(c[66]) );
  NOR U435 ( .A(n228), .B(n227), .Z(n251) );
  XOR U436 ( .A(b[3]), .B(b[2]), .Z(n252) );
  XOR U437 ( .A(b[3]), .B(a[0]), .Z(n229) );
  NAND U438 ( .A(n252), .B(n229), .Z(n230) );
  XOR U439 ( .A(b[1]), .B(b[2]), .Z(n9653) );
  OR U440 ( .A(n230), .B(n9653), .Z(n232) );
  XOR U441 ( .A(b[3]), .B(a[1]), .Z(n253) );
  NAND U442 ( .A(n9653), .B(n253), .Z(n231) );
  AND U443 ( .A(n232), .B(n231), .Z(n260) );
  NAND U444 ( .A(b[0]), .B(a[3]), .Z(n233) );
  XNOR U445 ( .A(b[1]), .B(n233), .Z(n235) );
  NANDN U446 ( .A(b[0]), .B(a[2]), .Z(n234) );
  NAND U447 ( .A(n235), .B(n234), .Z(n259) );
  XNOR U448 ( .A(n260), .B(n259), .Z(n250) );
  NAND U449 ( .A(b[1]), .B(b[2]), .Z(n236) );
  AND U450 ( .A(b[3]), .B(n236), .Z(n29556) );
  IV U451 ( .A(n9653), .Z(n28941) );
  NANDN U452 ( .A(n28941), .B(a[0]), .Z(n237) );
  AND U453 ( .A(n29556), .B(n237), .Z(n249) );
  XOR U454 ( .A(n250), .B(n249), .Z(n238) );
  XOR U455 ( .A(n251), .B(n238), .Z(n244) );
  XNOR U456 ( .A(sreg[67]), .B(n244), .Z(n246) );
  NANDN U457 ( .A(n239), .B(sreg[66]), .Z(n243) );
  NAND U458 ( .A(n241), .B(n240), .Z(n242) );
  NAND U459 ( .A(n243), .B(n242), .Z(n245) );
  XOR U460 ( .A(n246), .B(n245), .Z(c[67]) );
  NANDN U461 ( .A(n244), .B(sreg[67]), .Z(n248) );
  NAND U462 ( .A(n246), .B(n245), .Z(n247) );
  AND U463 ( .A(n248), .B(n247), .Z(n284) );
  XNOR U464 ( .A(n284), .B(sreg[68]), .Z(n286) );
  ANDN U465 ( .B(n252), .A(n9653), .Z(n9942) );
  NANDN U466 ( .A(n209), .B(n253), .Z(n255) );
  XOR U467 ( .A(b[3]), .B(a[2]), .Z(n265) );
  NANDN U468 ( .A(n28941), .B(n265), .Z(n254) );
  AND U469 ( .A(n255), .B(n254), .Z(n281) );
  XOR U470 ( .A(b[4]), .B(b[3]), .Z(n29552) );
  IV U471 ( .A(n29552), .Z(n29138) );
  ANDN U472 ( .B(a[0]), .A(n29138), .Z(n278) );
  NAND U473 ( .A(b[0]), .B(a[4]), .Z(n256) );
  XNOR U474 ( .A(b[1]), .B(n256), .Z(n258) );
  NANDN U475 ( .A(b[0]), .B(a[3]), .Z(n257) );
  NAND U476 ( .A(n258), .B(n257), .Z(n279) );
  XNOR U477 ( .A(n278), .B(n279), .Z(n280) );
  XNOR U478 ( .A(n281), .B(n280), .Z(n262) );
  NOR U479 ( .A(n260), .B(n259), .Z(n261) );
  XOR U480 ( .A(n262), .B(n261), .Z(n263) );
  XNOR U481 ( .A(n264), .B(n263), .Z(n285) );
  XOR U482 ( .A(n286), .B(n285), .Z(c[68]) );
  NANDN U483 ( .A(n209), .B(n265), .Z(n267) );
  XOR U484 ( .A(b[3]), .B(a[3]), .Z(n306) );
  NANDN U485 ( .A(n28941), .B(n306), .Z(n266) );
  AND U486 ( .A(n267), .B(n266), .Z(n313) );
  NAND U487 ( .A(b[3]), .B(b[4]), .Z(n268) );
  AND U488 ( .A(b[5]), .B(n268), .Z(n30104) );
  ANDN U489 ( .B(n30104), .A(n278), .Z(n312) );
  XNOR U490 ( .A(n313), .B(n312), .Z(n315) );
  XOR U491 ( .A(b[5]), .B(a[1]), .Z(n301) );
  NANDN U492 ( .A(n29138), .B(n301), .Z(n274) );
  ANDN U493 ( .B(b[4]), .A(b[5]), .Z(n269) );
  NAND U494 ( .A(n269), .B(a[0]), .Z(n271) );
  NANDN U495 ( .A(a[0]), .B(n30104), .Z(n270) );
  NAND U496 ( .A(n271), .B(n270), .Z(n272) );
  NAND U497 ( .A(n29138), .B(n272), .Z(n273) );
  NAND U498 ( .A(n274), .B(n273), .Z(n305) );
  NAND U499 ( .A(b[0]), .B(a[5]), .Z(n275) );
  XNOR U500 ( .A(b[1]), .B(n275), .Z(n277) );
  NANDN U501 ( .A(b[0]), .B(a[4]), .Z(n276) );
  NAND U502 ( .A(n277), .B(n276), .Z(n304) );
  XNOR U503 ( .A(n305), .B(n304), .Z(n314) );
  XOR U504 ( .A(n315), .B(n314), .Z(n295) );
  NANDN U505 ( .A(n279), .B(n278), .Z(n283) );
  NANDN U506 ( .A(n281), .B(n280), .Z(n282) );
  AND U507 ( .A(n283), .B(n282), .Z(n294) );
  XNOR U508 ( .A(n295), .B(n294), .Z(n296) );
  XOR U509 ( .A(n297), .B(n296), .Z(n289) );
  XNOR U510 ( .A(n289), .B(sreg[69]), .Z(n291) );
  NANDN U511 ( .A(n284), .B(sreg[68]), .Z(n288) );
  NAND U512 ( .A(n286), .B(n285), .Z(n287) );
  NAND U513 ( .A(n288), .B(n287), .Z(n290) );
  XOR U514 ( .A(n291), .B(n290), .Z(c[69]) );
  NANDN U515 ( .A(n289), .B(sreg[69]), .Z(n293) );
  NAND U516 ( .A(n291), .B(n290), .Z(n292) );
  AND U517 ( .A(n293), .B(n292), .Z(n350) );
  XNOR U518 ( .A(n350), .B(sreg[70]), .Z(n352) );
  NANDN U519 ( .A(n295), .B(n294), .Z(n299) );
  NAND U520 ( .A(n297), .B(n296), .Z(n298) );
  AND U521 ( .A(n299), .B(n298), .Z(n320) );
  XOR U522 ( .A(b[4]), .B(b[5]), .Z(n300) );
  ANDN U523 ( .B(n300), .A(n29552), .Z(n29551) );
  IV U524 ( .A(n29551), .Z(n28889) );
  NANDN U525 ( .A(n28889), .B(n301), .Z(n303) );
  XOR U526 ( .A(b[5]), .B(a[2]), .Z(n328) );
  NANDN U527 ( .A(n29138), .B(n328), .Z(n302) );
  AND U528 ( .A(n303), .B(n302), .Z(n345) );
  ANDN U529 ( .B(n305), .A(n304), .Z(n344) );
  XNOR U530 ( .A(n345), .B(n344), .Z(n347) );
  NANDN U531 ( .A(n209), .B(n306), .Z(n308) );
  XOR U532 ( .A(b[3]), .B(a[4]), .Z(n335) );
  NANDN U533 ( .A(n28941), .B(n335), .Z(n307) );
  AND U534 ( .A(n308), .B(n307), .Z(n341) );
  XOR U535 ( .A(b[6]), .B(b[5]), .Z(n30004) );
  IV U536 ( .A(n30004), .Z(n29735) );
  ANDN U537 ( .B(a[0]), .A(n29735), .Z(n338) );
  NAND U538 ( .A(b[0]), .B(a[6]), .Z(n309) );
  XNOR U539 ( .A(b[1]), .B(n309), .Z(n311) );
  NANDN U540 ( .A(b[0]), .B(a[5]), .Z(n310) );
  NAND U541 ( .A(n311), .B(n310), .Z(n339) );
  XNOR U542 ( .A(n338), .B(n339), .Z(n340) );
  XNOR U543 ( .A(n341), .B(n340), .Z(n346) );
  XOR U544 ( .A(n347), .B(n346), .Z(n319) );
  NANDN U545 ( .A(n313), .B(n312), .Z(n317) );
  NAND U546 ( .A(n315), .B(n314), .Z(n316) );
  AND U547 ( .A(n317), .B(n316), .Z(n318) );
  XOR U548 ( .A(n319), .B(n318), .Z(n321) );
  XNOR U549 ( .A(n320), .B(n321), .Z(n351) );
  XOR U550 ( .A(n352), .B(n351), .Z(c[70]) );
  NANDN U551 ( .A(n319), .B(n318), .Z(n323) );
  OR U552 ( .A(n321), .B(n320), .Z(n322) );
  AND U553 ( .A(n323), .B(n322), .Z(n362) );
  XOR U554 ( .A(b[7]), .B(b[6]), .Z(n378) );
  XOR U555 ( .A(b[7]), .B(a[0]), .Z(n324) );
  NAND U556 ( .A(n378), .B(n324), .Z(n325) );
  OR U557 ( .A(n325), .B(n30004), .Z(n327) );
  XOR U558 ( .A(b[7]), .B(a[1]), .Z(n379) );
  NAND U559 ( .A(n30004), .B(n379), .Z(n326) );
  AND U560 ( .A(n327), .B(n326), .Z(n386) );
  NANDN U561 ( .A(n28889), .B(n328), .Z(n330) );
  XOR U562 ( .A(b[5]), .B(a[3]), .Z(n390) );
  NANDN U563 ( .A(n29138), .B(n390), .Z(n329) );
  AND U564 ( .A(n330), .B(n329), .Z(n385) );
  XOR U565 ( .A(n386), .B(n385), .Z(n375) );
  NAND U566 ( .A(b[5]), .B(b[6]), .Z(n331) );
  AND U567 ( .A(b[7]), .B(n331), .Z(n30514) );
  ANDN U568 ( .B(n30514), .A(n338), .Z(n373) );
  NAND U569 ( .A(b[0]), .B(a[7]), .Z(n332) );
  XNOR U570 ( .A(b[1]), .B(n332), .Z(n334) );
  NANDN U571 ( .A(b[0]), .B(a[6]), .Z(n333) );
  NAND U572 ( .A(n334), .B(n333), .Z(n372) );
  XNOR U573 ( .A(n373), .B(n372), .Z(n374) );
  XNOR U574 ( .A(n375), .B(n374), .Z(n366) );
  NAND U575 ( .A(n9942), .B(n335), .Z(n337) );
  XNOR U576 ( .A(b[3]), .B(a[5]), .Z(n382) );
  NANDN U577 ( .A(n382), .B(n9653), .Z(n336) );
  NAND U578 ( .A(n337), .B(n336), .Z(n367) );
  XNOR U579 ( .A(n366), .B(n367), .Z(n368) );
  NANDN U580 ( .A(n339), .B(n338), .Z(n343) );
  NANDN U581 ( .A(n341), .B(n340), .Z(n342) );
  NAND U582 ( .A(n343), .B(n342), .Z(n369) );
  XNOR U583 ( .A(n368), .B(n369), .Z(n360) );
  NANDN U584 ( .A(n345), .B(n344), .Z(n349) );
  NAND U585 ( .A(n347), .B(n346), .Z(n348) );
  NAND U586 ( .A(n349), .B(n348), .Z(n361) );
  XOR U587 ( .A(n360), .B(n361), .Z(n363) );
  XOR U588 ( .A(n362), .B(n363), .Z(n355) );
  XNOR U589 ( .A(n355), .B(sreg[71]), .Z(n357) );
  NANDN U590 ( .A(n350), .B(sreg[70]), .Z(n354) );
  NAND U591 ( .A(n352), .B(n351), .Z(n353) );
  NAND U592 ( .A(n354), .B(n353), .Z(n356) );
  XOR U593 ( .A(n357), .B(n356), .Z(c[71]) );
  NANDN U594 ( .A(n355), .B(sreg[71]), .Z(n359) );
  NAND U595 ( .A(n357), .B(n356), .Z(n358) );
  AND U596 ( .A(n359), .B(n358), .Z(n436) );
  XNOR U597 ( .A(n436), .B(sreg[72]), .Z(n438) );
  NANDN U598 ( .A(n361), .B(n360), .Z(n365) );
  OR U599 ( .A(n363), .B(n362), .Z(n364) );
  AND U600 ( .A(n365), .B(n364), .Z(n432) );
  NANDN U601 ( .A(n367), .B(n366), .Z(n371) );
  NANDN U602 ( .A(n369), .B(n368), .Z(n370) );
  AND U603 ( .A(n371), .B(n370), .Z(n431) );
  NANDN U604 ( .A(n373), .B(n372), .Z(n377) );
  NANDN U605 ( .A(n375), .B(n374), .Z(n376) );
  AND U606 ( .A(n377), .B(n376), .Z(n396) );
  ANDN U607 ( .B(n378), .A(n30004), .Z(n30003) );
  IV U608 ( .A(n30003), .Z(n29499) );
  NANDN U609 ( .A(n29499), .B(n379), .Z(n381) );
  XOR U610 ( .A(b[7]), .B(a[2]), .Z(n410) );
  NANDN U611 ( .A(n29735), .B(n410), .Z(n380) );
  AND U612 ( .A(n381), .B(n380), .Z(n400) );
  NANDN U613 ( .A(n382), .B(n9942), .Z(n384) );
  XOR U614 ( .A(b[3]), .B(a[6]), .Z(n427) );
  NANDN U615 ( .A(n28941), .B(n427), .Z(n383) );
  NAND U616 ( .A(n384), .B(n383), .Z(n399) );
  XNOR U617 ( .A(n400), .B(n399), .Z(n402) );
  NOR U618 ( .A(n386), .B(n385), .Z(n401) );
  XOR U619 ( .A(n402), .B(n401), .Z(n394) );
  NAND U620 ( .A(b[0]), .B(a[8]), .Z(n387) );
  XNOR U621 ( .A(b[1]), .B(n387), .Z(n389) );
  NANDN U622 ( .A(b[0]), .B(a[7]), .Z(n388) );
  NAND U623 ( .A(n389), .B(n388), .Z(n407) );
  XOR U624 ( .A(b[8]), .B(b[7]), .Z(n30628) );
  IV U625 ( .A(n30628), .Z(n30267) );
  ANDN U626 ( .B(a[0]), .A(n30267), .Z(n420) );
  NANDN U627 ( .A(n28889), .B(n390), .Z(n392) );
  XOR U628 ( .A(b[5]), .B(a[4]), .Z(n421) );
  NANDN U629 ( .A(n29138), .B(n421), .Z(n391) );
  AND U630 ( .A(n392), .B(n391), .Z(n405) );
  XOR U631 ( .A(n420), .B(n405), .Z(n406) );
  XNOR U632 ( .A(n407), .B(n406), .Z(n393) );
  XNOR U633 ( .A(n394), .B(n393), .Z(n395) );
  XNOR U634 ( .A(n396), .B(n395), .Z(n430) );
  XOR U635 ( .A(n431), .B(n430), .Z(n433) );
  XNOR U636 ( .A(n432), .B(n433), .Z(n437) );
  XOR U637 ( .A(n438), .B(n437), .Z(c[72]) );
  NANDN U638 ( .A(n394), .B(n393), .Z(n398) );
  NANDN U639 ( .A(n396), .B(n395), .Z(n397) );
  AND U640 ( .A(n398), .B(n397), .Z(n446) );
  NANDN U641 ( .A(n400), .B(n399), .Z(n404) );
  NAND U642 ( .A(n402), .B(n401), .Z(n403) );
  AND U643 ( .A(n404), .B(n403), .Z(n485) );
  NANDN U644 ( .A(n405), .B(n420), .Z(n409) );
  OR U645 ( .A(n407), .B(n406), .Z(n408) );
  AND U646 ( .A(n409), .B(n408), .Z(n483) );
  NANDN U647 ( .A(n29499), .B(n410), .Z(n412) );
  XOR U648 ( .A(b[7]), .B(a[3]), .Z(n467) );
  NANDN U649 ( .A(n29735), .B(n467), .Z(n411) );
  AND U650 ( .A(n412), .B(n411), .Z(n477) );
  XOR U651 ( .A(b[9]), .B(a[1]), .Z(n474) );
  NANDN U652 ( .A(n30267), .B(n474), .Z(n419) );
  ANDN U653 ( .B(b[8]), .A(b[9]), .Z(n413) );
  NAND U654 ( .A(n413), .B(a[0]), .Z(n416) );
  NAND U655 ( .A(b[7]), .B(b[8]), .Z(n414) );
  NAND U656 ( .A(b[9]), .B(n414), .Z(n30898) );
  OR U657 ( .A(a[0]), .B(n30898), .Z(n415) );
  NAND U658 ( .A(n416), .B(n415), .Z(n417) );
  NAND U659 ( .A(n30267), .B(n417), .Z(n418) );
  NAND U660 ( .A(n419), .B(n418), .Z(n478) );
  XOR U661 ( .A(n477), .B(n478), .Z(n454) );
  NOR U662 ( .A(n30898), .B(n420), .Z(n453) );
  NANDN U663 ( .A(n28889), .B(n421), .Z(n423) );
  XOR U664 ( .A(b[5]), .B(a[5]), .Z(n470) );
  NANDN U665 ( .A(n29138), .B(n470), .Z(n422) );
  AND U666 ( .A(n423), .B(n422), .Z(n452) );
  XOR U667 ( .A(n453), .B(n452), .Z(n455) );
  XOR U668 ( .A(n454), .B(n455), .Z(n461) );
  NAND U669 ( .A(b[0]), .B(a[9]), .Z(n424) );
  XNOR U670 ( .A(b[1]), .B(n424), .Z(n426) );
  NANDN U671 ( .A(b[0]), .B(a[8]), .Z(n425) );
  NAND U672 ( .A(n426), .B(n425), .Z(n459) );
  NANDN U673 ( .A(n209), .B(n427), .Z(n429) );
  XOR U674 ( .A(b[3]), .B(a[7]), .Z(n479) );
  NANDN U675 ( .A(n28941), .B(n479), .Z(n428) );
  NAND U676 ( .A(n429), .B(n428), .Z(n458) );
  XNOR U677 ( .A(n459), .B(n458), .Z(n460) );
  XOR U678 ( .A(n461), .B(n460), .Z(n482) );
  XNOR U679 ( .A(n483), .B(n482), .Z(n484) );
  XOR U680 ( .A(n485), .B(n484), .Z(n447) );
  XNOR U681 ( .A(n446), .B(n447), .Z(n448) );
  NANDN U682 ( .A(n431), .B(n430), .Z(n435) );
  OR U683 ( .A(n433), .B(n432), .Z(n434) );
  NAND U684 ( .A(n435), .B(n434), .Z(n449) );
  XOR U685 ( .A(n448), .B(n449), .Z(n441) );
  XNOR U686 ( .A(sreg[73]), .B(n441), .Z(n443) );
  NANDN U687 ( .A(n436), .B(sreg[72]), .Z(n440) );
  NAND U688 ( .A(n438), .B(n437), .Z(n439) );
  NAND U689 ( .A(n440), .B(n439), .Z(n442) );
  XOR U690 ( .A(n443), .B(n442), .Z(c[73]) );
  NANDN U691 ( .A(n441), .B(sreg[73]), .Z(n445) );
  NAND U692 ( .A(n443), .B(n442), .Z(n444) );
  AND U693 ( .A(n445), .B(n444), .Z(n488) );
  XNOR U694 ( .A(n488), .B(sreg[74]), .Z(n490) );
  NANDN U695 ( .A(n447), .B(n446), .Z(n451) );
  NANDN U696 ( .A(n449), .B(n448), .Z(n450) );
  AND U697 ( .A(n451), .B(n450), .Z(n496) );
  NANDN U698 ( .A(n453), .B(n452), .Z(n457) );
  NANDN U699 ( .A(n455), .B(n454), .Z(n456) );
  AND U700 ( .A(n457), .B(n456), .Z(n540) );
  NANDN U701 ( .A(n459), .B(n458), .Z(n463) );
  NAND U702 ( .A(n461), .B(n460), .Z(n462) );
  AND U703 ( .A(n463), .B(n462), .Z(n539) );
  XNOR U704 ( .A(n540), .B(n539), .Z(n541) );
  NAND U705 ( .A(b[0]), .B(a[10]), .Z(n464) );
  XNOR U706 ( .A(b[1]), .B(n464), .Z(n466) );
  NANDN U707 ( .A(b[0]), .B(a[9]), .Z(n465) );
  NAND U708 ( .A(n466), .B(n465), .Z(n507) );
  XOR U709 ( .A(b[10]), .B(b[9]), .Z(n31060) );
  IV U710 ( .A(n31060), .Z(n30891) );
  ANDN U711 ( .B(a[0]), .A(n30891), .Z(n538) );
  NANDN U712 ( .A(n29499), .B(n467), .Z(n469) );
  XOR U713 ( .A(b[7]), .B(a[4]), .Z(n535) );
  NANDN U714 ( .A(n29735), .B(n535), .Z(n468) );
  AND U715 ( .A(n469), .B(n468), .Z(n505) );
  XOR U716 ( .A(n538), .B(n505), .Z(n506) );
  XOR U717 ( .A(n507), .B(n506), .Z(n502) );
  NANDN U718 ( .A(n28889), .B(n470), .Z(n472) );
  XOR U719 ( .A(b[5]), .B(a[6]), .Z(n529) );
  NANDN U720 ( .A(n29138), .B(n529), .Z(n471) );
  AND U721 ( .A(n472), .B(n471), .Z(n511) );
  XOR U722 ( .A(b[8]), .B(b[9]), .Z(n473) );
  ANDN U723 ( .B(n473), .A(n30628), .Z(n30627) );
  NANDN U724 ( .A(n210), .B(n474), .Z(n476) );
  XOR U725 ( .A(b[9]), .B(a[2]), .Z(n516) );
  NANDN U726 ( .A(n30267), .B(n516), .Z(n475) );
  NAND U727 ( .A(n476), .B(n475), .Z(n510) );
  XNOR U728 ( .A(n511), .B(n510), .Z(n513) );
  ANDN U729 ( .B(n478), .A(n477), .Z(n512) );
  XOR U730 ( .A(n513), .B(n512), .Z(n500) );
  NAND U731 ( .A(n9942), .B(n479), .Z(n481) );
  XNOR U732 ( .A(b[3]), .B(a[8]), .Z(n532) );
  NANDN U733 ( .A(n532), .B(n9653), .Z(n480) );
  AND U734 ( .A(n481), .B(n480), .Z(n499) );
  XNOR U735 ( .A(n500), .B(n499), .Z(n501) );
  XOR U736 ( .A(n502), .B(n501), .Z(n542) );
  XNOR U737 ( .A(n541), .B(n542), .Z(n493) );
  NANDN U738 ( .A(n483), .B(n482), .Z(n487) );
  NANDN U739 ( .A(n485), .B(n484), .Z(n486) );
  NAND U740 ( .A(n487), .B(n486), .Z(n494) );
  XNOR U741 ( .A(n493), .B(n494), .Z(n495) );
  XNOR U742 ( .A(n496), .B(n495), .Z(n489) );
  XOR U743 ( .A(n490), .B(n489), .Z(c[74]) );
  NANDN U744 ( .A(n488), .B(sreg[74]), .Z(n492) );
  NAND U745 ( .A(n490), .B(n489), .Z(n491) );
  AND U746 ( .A(n492), .B(n491), .Z(n547) );
  NANDN U747 ( .A(n494), .B(n493), .Z(n498) );
  NAND U748 ( .A(n496), .B(n495), .Z(n497) );
  AND U749 ( .A(n498), .B(n497), .Z(n553) );
  NANDN U750 ( .A(n500), .B(n499), .Z(n504) );
  NANDN U751 ( .A(n502), .B(n501), .Z(n503) );
  AND U752 ( .A(n504), .B(n503), .Z(n598) );
  NANDN U753 ( .A(n505), .B(n538), .Z(n509) );
  OR U754 ( .A(n507), .B(n506), .Z(n508) );
  AND U755 ( .A(n509), .B(n508), .Z(n596) );
  NANDN U756 ( .A(n511), .B(n510), .Z(n515) );
  NAND U757 ( .A(n513), .B(n512), .Z(n514) );
  AND U758 ( .A(n515), .B(n514), .Z(n592) );
  NANDN U759 ( .A(n210), .B(n516), .Z(n518) );
  XOR U760 ( .A(b[9]), .B(a[3]), .Z(n571) );
  NANDN U761 ( .A(n30267), .B(n571), .Z(n517) );
  AND U762 ( .A(n518), .B(n517), .Z(n556) );
  XOR U763 ( .A(b[11]), .B(a[1]), .Z(n568) );
  NANDN U764 ( .A(n30891), .B(n568), .Z(n525) );
  ANDN U765 ( .B(b[10]), .A(b[11]), .Z(n519) );
  NAND U766 ( .A(n519), .B(a[0]), .Z(n522) );
  NAND U767 ( .A(b[9]), .B(b[10]), .Z(n520) );
  AND U768 ( .A(b[11]), .B(n520), .Z(n31512) );
  NANDN U769 ( .A(a[0]), .B(n31512), .Z(n521) );
  NAND U770 ( .A(n522), .B(n521), .Z(n523) );
  NAND U771 ( .A(n30891), .B(n523), .Z(n524) );
  AND U772 ( .A(n525), .B(n524), .Z(n557) );
  XOR U773 ( .A(n556), .B(n557), .Z(n579) );
  NAND U774 ( .A(b[0]), .B(a[11]), .Z(n526) );
  XNOR U775 ( .A(b[1]), .B(n526), .Z(n528) );
  NANDN U776 ( .A(b[0]), .B(a[10]), .Z(n527) );
  NAND U777 ( .A(n528), .B(n527), .Z(n577) );
  NAND U778 ( .A(n29551), .B(n529), .Z(n531) );
  XNOR U779 ( .A(b[5]), .B(a[7]), .Z(n564) );
  NANDN U780 ( .A(n564), .B(n29552), .Z(n530) );
  NAND U781 ( .A(n531), .B(n530), .Z(n578) );
  XOR U782 ( .A(n577), .B(n578), .Z(n580) );
  XOR U783 ( .A(n579), .B(n580), .Z(n590) );
  NANDN U784 ( .A(n532), .B(n9942), .Z(n534) );
  XOR U785 ( .A(b[3]), .B(a[9]), .Z(n558) );
  NANDN U786 ( .A(n28941), .B(n558), .Z(n533) );
  AND U787 ( .A(n534), .B(n533), .Z(n586) );
  NANDN U788 ( .A(n29499), .B(n535), .Z(n537) );
  XOR U789 ( .A(b[7]), .B(a[5]), .Z(n561) );
  NANDN U790 ( .A(n29735), .B(n561), .Z(n536) );
  AND U791 ( .A(n537), .B(n536), .Z(n584) );
  ANDN U792 ( .B(n31512), .A(n538), .Z(n583) );
  XNOR U793 ( .A(n584), .B(n583), .Z(n585) );
  XNOR U794 ( .A(n586), .B(n585), .Z(n589) );
  XNOR U795 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U796 ( .A(n592), .B(n591), .Z(n595) );
  XNOR U797 ( .A(n596), .B(n595), .Z(n597) );
  XOR U798 ( .A(n598), .B(n597), .Z(n551) );
  NANDN U799 ( .A(n540), .B(n539), .Z(n544) );
  NANDN U800 ( .A(n542), .B(n541), .Z(n543) );
  NAND U801 ( .A(n544), .B(n543), .Z(n550) );
  XNOR U802 ( .A(n551), .B(n550), .Z(n552) );
  XNOR U803 ( .A(n553), .B(n552), .Z(n545) );
  XNOR U804 ( .A(sreg[75]), .B(n545), .Z(n546) );
  XNOR U805 ( .A(n547), .B(n546), .Z(c[75]) );
  NANDN U806 ( .A(sreg[75]), .B(n545), .Z(n549) );
  NAND U807 ( .A(n547), .B(n546), .Z(n548) );
  NAND U808 ( .A(n549), .B(n548), .Z(n660) );
  XNOR U809 ( .A(sreg[76]), .B(n660), .Z(n662) );
  NANDN U810 ( .A(n551), .B(n550), .Z(n555) );
  NANDN U811 ( .A(n553), .B(n552), .Z(n554) );
  AND U812 ( .A(n555), .B(n554), .Z(n603) );
  NOR U813 ( .A(n557), .B(n556), .Z(n650) );
  NAND U814 ( .A(n9942), .B(n558), .Z(n560) );
  XNOR U815 ( .A(b[3]), .B(a[10]), .Z(n632) );
  NANDN U816 ( .A(n632), .B(n9653), .Z(n559) );
  AND U817 ( .A(n560), .B(n559), .Z(n648) );
  NAND U818 ( .A(n30003), .B(n561), .Z(n563) );
  XNOR U819 ( .A(b[7]), .B(a[6]), .Z(n622) );
  NANDN U820 ( .A(n622), .B(n30004), .Z(n562) );
  NAND U821 ( .A(n563), .B(n562), .Z(n649) );
  XOR U822 ( .A(n648), .B(n649), .Z(n651) );
  XOR U823 ( .A(n650), .B(n651), .Z(n616) );
  NANDN U824 ( .A(n564), .B(n29551), .Z(n566) );
  XOR U825 ( .A(b[5]), .B(a[8]), .Z(n639) );
  NANDN U826 ( .A(n29138), .B(n639), .Z(n565) );
  AND U827 ( .A(n566), .B(n565), .Z(n614) );
  XOR U828 ( .A(b[10]), .B(b[11]), .Z(n567) );
  ANDN U829 ( .B(n567), .A(n31060), .Z(n31059) );
  IV U830 ( .A(n31059), .Z(n30482) );
  NANDN U831 ( .A(n30482), .B(n568), .Z(n570) );
  XOR U832 ( .A(b[11]), .B(a[2]), .Z(n625) );
  NANDN U833 ( .A(n30891), .B(n625), .Z(n569) );
  NAND U834 ( .A(n570), .B(n569), .Z(n613) );
  XNOR U835 ( .A(n614), .B(n613), .Z(n615) );
  XNOR U836 ( .A(n616), .B(n615), .Z(n610) );
  XOR U837 ( .A(b[12]), .B(b[11]), .Z(n31508) );
  IV U838 ( .A(n31508), .Z(n31293) );
  ANDN U839 ( .B(a[0]), .A(n31293), .Z(n642) );
  NANDN U840 ( .A(n210), .B(n571), .Z(n573) );
  XOR U841 ( .A(b[9]), .B(a[4]), .Z(n635) );
  NANDN U842 ( .A(n30267), .B(n635), .Z(n572) );
  AND U843 ( .A(n573), .B(n572), .Z(n643) );
  XNOR U844 ( .A(n642), .B(n643), .Z(n644) );
  NAND U845 ( .A(b[0]), .B(a[12]), .Z(n574) );
  XNOR U846 ( .A(b[1]), .B(n574), .Z(n576) );
  NANDN U847 ( .A(b[0]), .B(a[11]), .Z(n575) );
  NAND U848 ( .A(n576), .B(n575), .Z(n645) );
  XNOR U849 ( .A(n644), .B(n645), .Z(n607) );
  NANDN U850 ( .A(n578), .B(n577), .Z(n582) );
  OR U851 ( .A(n580), .B(n579), .Z(n581) );
  NAND U852 ( .A(n582), .B(n581), .Z(n608) );
  XNOR U853 ( .A(n607), .B(n608), .Z(n609) );
  XOR U854 ( .A(n610), .B(n609), .Z(n657) );
  NANDN U855 ( .A(n584), .B(n583), .Z(n588) );
  NANDN U856 ( .A(n586), .B(n585), .Z(n587) );
  AND U857 ( .A(n588), .B(n587), .Z(n654) );
  NANDN U858 ( .A(n590), .B(n589), .Z(n594) );
  NANDN U859 ( .A(n592), .B(n591), .Z(n593) );
  NAND U860 ( .A(n594), .B(n593), .Z(n655) );
  XNOR U861 ( .A(n654), .B(n655), .Z(n656) );
  XNOR U862 ( .A(n657), .B(n656), .Z(n601) );
  NANDN U863 ( .A(n596), .B(n595), .Z(n600) );
  NAND U864 ( .A(n598), .B(n597), .Z(n599) );
  NAND U865 ( .A(n600), .B(n599), .Z(n602) );
  XOR U866 ( .A(n601), .B(n602), .Z(n604) );
  XNOR U867 ( .A(n603), .B(n604), .Z(n661) );
  XOR U868 ( .A(n662), .B(n661), .Z(c[76]) );
  NANDN U869 ( .A(n602), .B(n601), .Z(n606) );
  OR U870 ( .A(n604), .B(n603), .Z(n605) );
  AND U871 ( .A(n606), .B(n605), .Z(n672) );
  NANDN U872 ( .A(n608), .B(n607), .Z(n612) );
  NAND U873 ( .A(n610), .B(n609), .Z(n611) );
  AND U874 ( .A(n612), .B(n611), .Z(n726) );
  NANDN U875 ( .A(n614), .B(n613), .Z(n618) );
  NANDN U876 ( .A(n616), .B(n615), .Z(n617) );
  AND U877 ( .A(n618), .B(n617), .Z(n725) );
  NAND U878 ( .A(b[0]), .B(a[13]), .Z(n619) );
  XNOR U879 ( .A(b[1]), .B(n619), .Z(n621) );
  NANDN U880 ( .A(b[0]), .B(a[12]), .Z(n620) );
  NAND U881 ( .A(n621), .B(n620), .Z(n710) );
  NANDN U882 ( .A(n622), .B(n30003), .Z(n624) );
  XOR U883 ( .A(b[7]), .B(a[7]), .Z(n703) );
  NANDN U884 ( .A(n29735), .B(n703), .Z(n623) );
  NAND U885 ( .A(n624), .B(n623), .Z(n709) );
  XNOR U886 ( .A(n710), .B(n709), .Z(n712) );
  NANDN U887 ( .A(n30482), .B(n625), .Z(n627) );
  XOR U888 ( .A(b[11]), .B(a[3]), .Z(n697) );
  NANDN U889 ( .A(n30891), .B(n697), .Z(n626) );
  AND U890 ( .A(n627), .B(n626), .Z(n722) );
  XOR U891 ( .A(b[13]), .B(b[12]), .Z(n715) );
  XOR U892 ( .A(b[13]), .B(a[0]), .Z(n628) );
  NAND U893 ( .A(n715), .B(n628), .Z(n629) );
  OR U894 ( .A(n629), .B(n31508), .Z(n631) );
  XOR U895 ( .A(b[13]), .B(a[1]), .Z(n716) );
  NAND U896 ( .A(n31508), .B(n716), .Z(n630) );
  NAND U897 ( .A(n631), .B(n630), .Z(n723) );
  XNOR U898 ( .A(n722), .B(n723), .Z(n711) );
  XOR U899 ( .A(n712), .B(n711), .Z(n684) );
  NANDN U900 ( .A(n632), .B(n9942), .Z(n634) );
  XOR U901 ( .A(b[3]), .B(a[11]), .Z(n706) );
  NANDN U902 ( .A(n28941), .B(n706), .Z(n633) );
  AND U903 ( .A(n634), .B(n633), .Z(n689) );
  NANDN U904 ( .A(n210), .B(n635), .Z(n637) );
  XOR U905 ( .A(b[9]), .B(a[5]), .Z(n719) );
  NANDN U906 ( .A(n30267), .B(n719), .Z(n636) );
  NAND U907 ( .A(n637), .B(n636), .Z(n688) );
  XNOR U908 ( .A(n689), .B(n688), .Z(n691) );
  NAND U909 ( .A(b[11]), .B(b[12]), .Z(n638) );
  AND U910 ( .A(b[13]), .B(n638), .Z(n32142) );
  ANDN U911 ( .B(n32142), .A(n642), .Z(n690) );
  XOR U912 ( .A(n691), .B(n690), .Z(n683) );
  NAND U913 ( .A(n29551), .B(n639), .Z(n641) );
  XNOR U914 ( .A(b[5]), .B(a[9]), .Z(n700) );
  NANDN U915 ( .A(n700), .B(n29552), .Z(n640) );
  AND U916 ( .A(n641), .B(n640), .Z(n682) );
  XOR U917 ( .A(n683), .B(n682), .Z(n685) );
  XOR U918 ( .A(n684), .B(n685), .Z(n679) );
  NANDN U919 ( .A(n643), .B(n642), .Z(n647) );
  NANDN U920 ( .A(n645), .B(n644), .Z(n646) );
  AND U921 ( .A(n647), .B(n646), .Z(n677) );
  NANDN U922 ( .A(n649), .B(n648), .Z(n653) );
  OR U923 ( .A(n651), .B(n650), .Z(n652) );
  AND U924 ( .A(n653), .B(n652), .Z(n676) );
  XNOR U925 ( .A(n677), .B(n676), .Z(n678) );
  XNOR U926 ( .A(n679), .B(n678), .Z(n724) );
  XOR U927 ( .A(n725), .B(n724), .Z(n727) );
  XOR U928 ( .A(n726), .B(n727), .Z(n671) );
  NANDN U929 ( .A(n655), .B(n654), .Z(n659) );
  NANDN U930 ( .A(n657), .B(n656), .Z(n658) );
  NAND U931 ( .A(n659), .B(n658), .Z(n670) );
  XOR U932 ( .A(n671), .B(n670), .Z(n673) );
  XOR U933 ( .A(n672), .B(n673), .Z(n665) );
  XNOR U934 ( .A(n665), .B(sreg[77]), .Z(n667) );
  NANDN U935 ( .A(n660), .B(sreg[76]), .Z(n664) );
  NAND U936 ( .A(n662), .B(n661), .Z(n663) );
  NAND U937 ( .A(n664), .B(n663), .Z(n666) );
  XOR U938 ( .A(n667), .B(n666), .Z(c[77]) );
  NANDN U939 ( .A(n665), .B(sreg[77]), .Z(n669) );
  NAND U940 ( .A(n667), .B(n666), .Z(n668) );
  AND U941 ( .A(n669), .B(n668), .Z(n797) );
  XNOR U942 ( .A(sreg[78]), .B(n797), .Z(n799) );
  NANDN U943 ( .A(n671), .B(n670), .Z(n675) );
  OR U944 ( .A(n673), .B(n672), .Z(n674) );
  AND U945 ( .A(n675), .B(n674), .Z(n733) );
  NANDN U946 ( .A(n677), .B(n676), .Z(n681) );
  NANDN U947 ( .A(n679), .B(n678), .Z(n680) );
  AND U948 ( .A(n681), .B(n680), .Z(n793) );
  NANDN U949 ( .A(n683), .B(n682), .Z(n687) );
  OR U950 ( .A(n685), .B(n684), .Z(n686) );
  AND U951 ( .A(n687), .B(n686), .Z(n791) );
  NANDN U952 ( .A(n689), .B(n688), .Z(n693) );
  NAND U953 ( .A(n691), .B(n690), .Z(n692) );
  AND U954 ( .A(n693), .B(n692), .Z(n778) );
  NAND U955 ( .A(b[0]), .B(a[14]), .Z(n694) );
  XNOR U956 ( .A(b[1]), .B(n694), .Z(n696) );
  NANDN U957 ( .A(b[0]), .B(a[13]), .Z(n695) );
  NAND U958 ( .A(n696), .B(n695), .Z(n784) );
  XOR U959 ( .A(b[14]), .B(b[13]), .Z(n32024) );
  IV U960 ( .A(n32024), .Z(n31925) );
  ANDN U961 ( .B(a[0]), .A(n31925), .Z(n781) );
  NANDN U962 ( .A(n30482), .B(n697), .Z(n699) );
  XOR U963 ( .A(b[11]), .B(a[4]), .Z(n751) );
  NANDN U964 ( .A(n30891), .B(n751), .Z(n698) );
  AND U965 ( .A(n699), .B(n698), .Z(n782) );
  XNOR U966 ( .A(n781), .B(n782), .Z(n783) );
  XNOR U967 ( .A(n784), .B(n783), .Z(n775) );
  NANDN U968 ( .A(n700), .B(n29551), .Z(n702) );
  XOR U969 ( .A(b[5]), .B(a[10]), .Z(n745) );
  NANDN U970 ( .A(n29138), .B(n745), .Z(n701) );
  AND U971 ( .A(n702), .B(n701), .Z(n772) );
  NANDN U972 ( .A(n29499), .B(n703), .Z(n705) );
  XOR U973 ( .A(b[7]), .B(a[8]), .Z(n742) );
  NANDN U974 ( .A(n29735), .B(n742), .Z(n704) );
  AND U975 ( .A(n705), .B(n704), .Z(n770) );
  NANDN U976 ( .A(n209), .B(n706), .Z(n708) );
  XOR U977 ( .A(b[3]), .B(a[12]), .Z(n748) );
  NANDN U978 ( .A(n28941), .B(n748), .Z(n707) );
  NAND U979 ( .A(n708), .B(n707), .Z(n769) );
  XNOR U980 ( .A(n770), .B(n769), .Z(n771) );
  XOR U981 ( .A(n772), .B(n771), .Z(n776) );
  XNOR U982 ( .A(n775), .B(n776), .Z(n777) );
  XNOR U983 ( .A(n778), .B(n777), .Z(n738) );
  NANDN U984 ( .A(n710), .B(n709), .Z(n714) );
  NAND U985 ( .A(n712), .B(n711), .Z(n713) );
  AND U986 ( .A(n714), .B(n713), .Z(n737) );
  ANDN U987 ( .B(n715), .A(n31508), .Z(n31507) );
  IV U988 ( .A(n31507), .Z(n31055) );
  NANDN U989 ( .A(n31055), .B(n716), .Z(n718) );
  XOR U990 ( .A(b[13]), .B(a[2]), .Z(n766) );
  NANDN U991 ( .A(n31293), .B(n766), .Z(n717) );
  AND U992 ( .A(n718), .B(n717), .Z(n788) );
  NANDN U993 ( .A(n210), .B(n719), .Z(n721) );
  XOR U994 ( .A(b[9]), .B(a[6]), .Z(n758) );
  NANDN U995 ( .A(n30267), .B(n758), .Z(n720) );
  NAND U996 ( .A(n721), .B(n720), .Z(n787) );
  XNOR U997 ( .A(n788), .B(n787), .Z(n790) );
  ANDN U998 ( .B(n723), .A(n722), .Z(n789) );
  XOR U999 ( .A(n790), .B(n789), .Z(n736) );
  XOR U1000 ( .A(n737), .B(n736), .Z(n739) );
  XOR U1001 ( .A(n738), .B(n739), .Z(n792) );
  XOR U1002 ( .A(n791), .B(n792), .Z(n794) );
  XOR U1003 ( .A(n793), .B(n794), .Z(n731) );
  NANDN U1004 ( .A(n725), .B(n724), .Z(n729) );
  OR U1005 ( .A(n727), .B(n726), .Z(n728) );
  AND U1006 ( .A(n729), .B(n728), .Z(n730) );
  XNOR U1007 ( .A(n731), .B(n730), .Z(n732) );
  XNOR U1008 ( .A(n733), .B(n732), .Z(n798) );
  XNOR U1009 ( .A(n799), .B(n798), .Z(c[78]) );
  NANDN U1010 ( .A(n731), .B(n730), .Z(n735) );
  NANDN U1011 ( .A(n733), .B(n732), .Z(n734) );
  AND U1012 ( .A(n735), .B(n734), .Z(n809) );
  NANDN U1013 ( .A(n737), .B(n736), .Z(n741) );
  NANDN U1014 ( .A(n739), .B(n738), .Z(n740) );
  AND U1015 ( .A(n741), .B(n740), .Z(n871) );
  NANDN U1016 ( .A(n29499), .B(n742), .Z(n744) );
  XOR U1017 ( .A(b[7]), .B(a[9]), .Z(n851) );
  NANDN U1018 ( .A(n29735), .B(n851), .Z(n743) );
  AND U1019 ( .A(n744), .B(n743), .Z(n838) );
  NANDN U1020 ( .A(n28889), .B(n745), .Z(n747) );
  XOR U1021 ( .A(b[5]), .B(a[11]), .Z(n861) );
  NANDN U1022 ( .A(n29138), .B(n861), .Z(n746) );
  AND U1023 ( .A(n747), .B(n746), .Z(n834) );
  NANDN U1024 ( .A(n209), .B(n748), .Z(n750) );
  XOR U1025 ( .A(b[3]), .B(a[13]), .Z(n845) );
  NANDN U1026 ( .A(n28941), .B(n845), .Z(n749) );
  AND U1027 ( .A(n750), .B(n749), .Z(n832) );
  NANDN U1028 ( .A(n30482), .B(n751), .Z(n753) );
  XOR U1029 ( .A(b[11]), .B(a[5]), .Z(n854) );
  NANDN U1030 ( .A(n30891), .B(n854), .Z(n752) );
  NAND U1031 ( .A(n753), .B(n752), .Z(n831) );
  XNOR U1032 ( .A(n832), .B(n831), .Z(n833) );
  XNOR U1033 ( .A(n834), .B(n833), .Z(n837) );
  XNOR U1034 ( .A(n838), .B(n837), .Z(n840) );
  NAND U1035 ( .A(b[13]), .B(b[14]), .Z(n754) );
  AND U1036 ( .A(b[15]), .B(n754), .Z(n32535) );
  ANDN U1037 ( .B(n32535), .A(n781), .Z(n839) );
  XOR U1038 ( .A(n840), .B(n839), .Z(n866) );
  NAND U1039 ( .A(b[0]), .B(a[15]), .Z(n755) );
  XNOR U1040 ( .A(b[1]), .B(n755), .Z(n757) );
  NANDN U1041 ( .A(b[0]), .B(a[14]), .Z(n756) );
  NAND U1042 ( .A(n757), .B(n756), .Z(n826) );
  NANDN U1043 ( .A(n210), .B(n758), .Z(n760) );
  XOR U1044 ( .A(b[9]), .B(a[7]), .Z(n848) );
  NANDN U1045 ( .A(n30267), .B(n848), .Z(n759) );
  NAND U1046 ( .A(n760), .B(n759), .Z(n825) );
  XNOR U1047 ( .A(n826), .B(n825), .Z(n828) );
  XOR U1048 ( .A(b[15]), .B(a[0]), .Z(n763) );
  XOR U1049 ( .A(b[15]), .B(b[13]), .Z(n761) );
  XOR U1050 ( .A(b[15]), .B(b[14]), .Z(n857) );
  AND U1051 ( .A(n761), .B(n857), .Z(n762) );
  NAND U1052 ( .A(n763), .B(n762), .Z(n765) );
  XOR U1053 ( .A(b[15]), .B(a[1]), .Z(n858) );
  NANDN U1054 ( .A(n31925), .B(n858), .Z(n764) );
  AND U1055 ( .A(n765), .B(n764), .Z(n843) );
  NANDN U1056 ( .A(n31055), .B(n766), .Z(n768) );
  XOR U1057 ( .A(b[13]), .B(a[3]), .Z(n822) );
  NANDN U1058 ( .A(n31293), .B(n822), .Z(n767) );
  NAND U1059 ( .A(n768), .B(n767), .Z(n844) );
  XNOR U1060 ( .A(n843), .B(n844), .Z(n827) );
  XOR U1061 ( .A(n828), .B(n827), .Z(n865) );
  NANDN U1062 ( .A(n770), .B(n769), .Z(n774) );
  NANDN U1063 ( .A(n772), .B(n771), .Z(n773) );
  AND U1064 ( .A(n774), .B(n773), .Z(n864) );
  XOR U1065 ( .A(n865), .B(n864), .Z(n867) );
  XNOR U1066 ( .A(n866), .B(n867), .Z(n870) );
  XNOR U1067 ( .A(n871), .B(n870), .Z(n873) );
  NANDN U1068 ( .A(n776), .B(n775), .Z(n780) );
  NANDN U1069 ( .A(n778), .B(n777), .Z(n779) );
  AND U1070 ( .A(n780), .B(n779), .Z(n816) );
  NANDN U1071 ( .A(n782), .B(n781), .Z(n786) );
  NANDN U1072 ( .A(n784), .B(n783), .Z(n785) );
  AND U1073 ( .A(n786), .B(n785), .Z(n814) );
  XNOR U1074 ( .A(n814), .B(n813), .Z(n815) );
  XNOR U1075 ( .A(n816), .B(n815), .Z(n872) );
  XOR U1076 ( .A(n873), .B(n872), .Z(n808) );
  NANDN U1077 ( .A(n792), .B(n791), .Z(n796) );
  OR U1078 ( .A(n794), .B(n793), .Z(n795) );
  AND U1079 ( .A(n796), .B(n795), .Z(n807) );
  XOR U1080 ( .A(n808), .B(n807), .Z(n810) );
  XOR U1081 ( .A(n809), .B(n810), .Z(n802) );
  XNOR U1082 ( .A(n802), .B(sreg[79]), .Z(n804) );
  NANDN U1083 ( .A(sreg[78]), .B(n797), .Z(n801) );
  NAND U1084 ( .A(n799), .B(n798), .Z(n800) );
  AND U1085 ( .A(n801), .B(n800), .Z(n803) );
  XOR U1086 ( .A(n804), .B(n803), .Z(c[79]) );
  NANDN U1087 ( .A(n802), .B(sreg[79]), .Z(n806) );
  NAND U1088 ( .A(n804), .B(n803), .Z(n805) );
  AND U1089 ( .A(n806), .B(n805), .Z(n876) );
  XNOR U1090 ( .A(n876), .B(sreg[80]), .Z(n878) );
  NANDN U1091 ( .A(n808), .B(n807), .Z(n812) );
  OR U1092 ( .A(n810), .B(n809), .Z(n811) );
  AND U1093 ( .A(n812), .B(n811), .Z(n883) );
  NANDN U1094 ( .A(n814), .B(n813), .Z(n818) );
  NANDN U1095 ( .A(n816), .B(n815), .Z(n817) );
  AND U1096 ( .A(n818), .B(n817), .Z(n954) );
  NAND U1097 ( .A(b[0]), .B(a[16]), .Z(n819) );
  XNOR U1098 ( .A(b[1]), .B(n819), .Z(n821) );
  NANDN U1099 ( .A(b[0]), .B(a[15]), .Z(n820) );
  NAND U1100 ( .A(n821), .B(n820), .Z(n889) );
  XOR U1101 ( .A(b[16]), .B(b[15]), .Z(n32545) );
  IV U1102 ( .A(n32545), .Z(n32292) );
  ANDN U1103 ( .B(a[0]), .A(n32292), .Z(n900) );
  NANDN U1104 ( .A(n31055), .B(n822), .Z(n824) );
  XOR U1105 ( .A(b[13]), .B(a[4]), .Z(n928) );
  NANDN U1106 ( .A(n31293), .B(n928), .Z(n823) );
  AND U1107 ( .A(n824), .B(n823), .Z(n887) );
  XOR U1108 ( .A(n900), .B(n887), .Z(n888) );
  XOR U1109 ( .A(n889), .B(n888), .Z(n947) );
  NANDN U1110 ( .A(n826), .B(n825), .Z(n830) );
  NAND U1111 ( .A(n828), .B(n827), .Z(n829) );
  AND U1112 ( .A(n830), .B(n829), .Z(n946) );
  XNOR U1113 ( .A(n947), .B(n946), .Z(n949) );
  NANDN U1114 ( .A(n832), .B(n831), .Z(n836) );
  NANDN U1115 ( .A(n834), .B(n833), .Z(n835) );
  AND U1116 ( .A(n836), .B(n835), .Z(n948) );
  XOR U1117 ( .A(n949), .B(n948), .Z(n943) );
  NANDN U1118 ( .A(n838), .B(n837), .Z(n842) );
  NAND U1119 ( .A(n840), .B(n839), .Z(n841) );
  AND U1120 ( .A(n842), .B(n841), .Z(n941) );
  ANDN U1121 ( .B(n844), .A(n843), .Z(n921) );
  NAND U1122 ( .A(n9942), .B(n845), .Z(n847) );
  XNOR U1123 ( .A(b[3]), .B(a[14]), .Z(n910) );
  NANDN U1124 ( .A(n910), .B(n9653), .Z(n846) );
  AND U1125 ( .A(n847), .B(n846), .Z(n919) );
  NAND U1126 ( .A(n30627), .B(n848), .Z(n850) );
  XNOR U1127 ( .A(b[9]), .B(a[8]), .Z(n901) );
  NANDN U1128 ( .A(n901), .B(n30628), .Z(n849) );
  NAND U1129 ( .A(n850), .B(n849), .Z(n920) );
  XOR U1130 ( .A(n919), .B(n920), .Z(n922) );
  XOR U1131 ( .A(n921), .B(n922), .Z(n916) );
  NANDN U1132 ( .A(n29499), .B(n851), .Z(n853) );
  XOR U1133 ( .A(b[7]), .B(a[10]), .Z(n931) );
  NANDN U1134 ( .A(n29735), .B(n931), .Z(n852) );
  AND U1135 ( .A(n853), .B(n852), .Z(n914) );
  NANDN U1136 ( .A(n30482), .B(n854), .Z(n856) );
  XOR U1137 ( .A(b[11]), .B(a[6]), .Z(n925) );
  NANDN U1138 ( .A(n30891), .B(n925), .Z(n855) );
  AND U1139 ( .A(n856), .B(n855), .Z(n937) );
  ANDN U1140 ( .B(n857), .A(n32024), .Z(n32023) );
  IV U1141 ( .A(n32023), .Z(n31536) );
  NANDN U1142 ( .A(n31536), .B(n858), .Z(n860) );
  XOR U1143 ( .A(b[15]), .B(a[2]), .Z(n896) );
  NANDN U1144 ( .A(n31925), .B(n896), .Z(n859) );
  AND U1145 ( .A(n860), .B(n859), .Z(n935) );
  NANDN U1146 ( .A(n28889), .B(n861), .Z(n863) );
  XOR U1147 ( .A(b[5]), .B(a[12]), .Z(n907) );
  NANDN U1148 ( .A(n29138), .B(n907), .Z(n862) );
  NAND U1149 ( .A(n863), .B(n862), .Z(n934) );
  XNOR U1150 ( .A(n935), .B(n934), .Z(n936) );
  XNOR U1151 ( .A(n937), .B(n936), .Z(n913) );
  XNOR U1152 ( .A(n914), .B(n913), .Z(n915) );
  XNOR U1153 ( .A(n916), .B(n915), .Z(n940) );
  XNOR U1154 ( .A(n941), .B(n940), .Z(n942) );
  XNOR U1155 ( .A(n943), .B(n942), .Z(n952) );
  NANDN U1156 ( .A(n865), .B(n864), .Z(n869) );
  OR U1157 ( .A(n867), .B(n866), .Z(n868) );
  NAND U1158 ( .A(n869), .B(n868), .Z(n953) );
  XOR U1159 ( .A(n952), .B(n953), .Z(n955) );
  XOR U1160 ( .A(n954), .B(n955), .Z(n882) );
  NANDN U1161 ( .A(n871), .B(n870), .Z(n875) );
  NAND U1162 ( .A(n873), .B(n872), .Z(n874) );
  AND U1163 ( .A(n875), .B(n874), .Z(n881) );
  XOR U1164 ( .A(n882), .B(n881), .Z(n884) );
  XNOR U1165 ( .A(n883), .B(n884), .Z(n877) );
  XOR U1166 ( .A(n878), .B(n877), .Z(c[80]) );
  NANDN U1167 ( .A(n876), .B(sreg[80]), .Z(n880) );
  NAND U1168 ( .A(n878), .B(n877), .Z(n879) );
  AND U1169 ( .A(n880), .B(n879), .Z(n960) );
  NANDN U1170 ( .A(n882), .B(n881), .Z(n886) );
  OR U1171 ( .A(n884), .B(n883), .Z(n885) );
  AND U1172 ( .A(n886), .B(n885), .Z(n966) );
  NANDN U1173 ( .A(n887), .B(n900), .Z(n891) );
  OR U1174 ( .A(n889), .B(n888), .Z(n890) );
  AND U1175 ( .A(n891), .B(n890), .Z(n983) );
  XOR U1176 ( .A(b[17]), .B(b[16]), .Z(n1010) );
  XOR U1177 ( .A(b[17]), .B(a[0]), .Z(n892) );
  NAND U1178 ( .A(n1010), .B(n892), .Z(n893) );
  OR U1179 ( .A(n893), .B(n32545), .Z(n895) );
  XOR U1180 ( .A(b[17]), .B(a[1]), .Z(n1011) );
  NAND U1181 ( .A(n32545), .B(n1011), .Z(n894) );
  AND U1182 ( .A(n895), .B(n894), .Z(n1006) );
  NANDN U1183 ( .A(n31536), .B(n896), .Z(n898) );
  XOR U1184 ( .A(b[15]), .B(a[3]), .Z(n1002) );
  NANDN U1185 ( .A(n31925), .B(n1002), .Z(n897) );
  AND U1186 ( .A(n898), .B(n897), .Z(n1005) );
  XOR U1187 ( .A(n1006), .B(n1005), .Z(n995) );
  NAND U1188 ( .A(b[15]), .B(b[16]), .Z(n899) );
  NAND U1189 ( .A(b[17]), .B(n899), .Z(n32830) );
  NOR U1190 ( .A(n32830), .B(n900), .Z(n994) );
  NANDN U1191 ( .A(n901), .B(n30627), .Z(n903) );
  XNOR U1192 ( .A(b[9]), .B(a[9]), .Z(n1026) );
  NANDN U1193 ( .A(n1026), .B(n30628), .Z(n902) );
  AND U1194 ( .A(n903), .B(n902), .Z(n993) );
  XOR U1195 ( .A(n994), .B(n993), .Z(n996) );
  XOR U1196 ( .A(n995), .B(n996), .Z(n982) );
  NAND U1197 ( .A(b[0]), .B(a[17]), .Z(n904) );
  XNOR U1198 ( .A(b[1]), .B(n904), .Z(n906) );
  NANDN U1199 ( .A(b[0]), .B(a[16]), .Z(n905) );
  NAND U1200 ( .A(n906), .B(n905), .Z(n988) );
  NANDN U1201 ( .A(n28889), .B(n907), .Z(n909) );
  XOR U1202 ( .A(b[5]), .B(a[13]), .Z(n1020) );
  NANDN U1203 ( .A(n29138), .B(n1020), .Z(n908) );
  NAND U1204 ( .A(n909), .B(n908), .Z(n987) );
  XNOR U1205 ( .A(n988), .B(n987), .Z(n990) );
  NANDN U1206 ( .A(n910), .B(n9942), .Z(n912) );
  XNOR U1207 ( .A(b[3]), .B(a[15]), .Z(n1032) );
  NANDN U1208 ( .A(n1032), .B(n9653), .Z(n911) );
  NAND U1209 ( .A(n912), .B(n911), .Z(n989) );
  XOR U1210 ( .A(n990), .B(n989), .Z(n981) );
  XOR U1211 ( .A(n982), .B(n981), .Z(n984) );
  XOR U1212 ( .A(n983), .B(n984), .Z(n970) );
  NANDN U1213 ( .A(n914), .B(n913), .Z(n918) );
  NANDN U1214 ( .A(n916), .B(n915), .Z(n917) );
  AND U1215 ( .A(n918), .B(n917), .Z(n969) );
  XNOR U1216 ( .A(n970), .B(n969), .Z(n972) );
  NANDN U1217 ( .A(n920), .B(n919), .Z(n924) );
  OR U1218 ( .A(n922), .B(n921), .Z(n923) );
  AND U1219 ( .A(n924), .B(n923), .Z(n976) );
  NANDN U1220 ( .A(n30482), .B(n925), .Z(n927) );
  XOR U1221 ( .A(b[11]), .B(a[7]), .Z(n1007) );
  NANDN U1222 ( .A(n30891), .B(n1007), .Z(n926) );
  AND U1223 ( .A(n927), .B(n926), .Z(n1016) );
  NANDN U1224 ( .A(n31055), .B(n928), .Z(n930) );
  XOR U1225 ( .A(b[13]), .B(a[5]), .Z(n1029) );
  NANDN U1226 ( .A(n31293), .B(n1029), .Z(n929) );
  AND U1227 ( .A(n930), .B(n929), .Z(n1015) );
  NANDN U1228 ( .A(n29499), .B(n931), .Z(n933) );
  XOR U1229 ( .A(b[7]), .B(a[11]), .Z(n1023) );
  NANDN U1230 ( .A(n29735), .B(n1023), .Z(n932) );
  NAND U1231 ( .A(n933), .B(n932), .Z(n1014) );
  XOR U1232 ( .A(n1015), .B(n1014), .Z(n1017) );
  XNOR U1233 ( .A(n1016), .B(n1017), .Z(n975) );
  XNOR U1234 ( .A(n976), .B(n975), .Z(n977) );
  NANDN U1235 ( .A(n935), .B(n934), .Z(n939) );
  NANDN U1236 ( .A(n937), .B(n936), .Z(n938) );
  NAND U1237 ( .A(n939), .B(n938), .Z(n978) );
  XNOR U1238 ( .A(n977), .B(n978), .Z(n971) );
  XOR U1239 ( .A(n972), .B(n971), .Z(n1037) );
  NANDN U1240 ( .A(n941), .B(n940), .Z(n945) );
  NANDN U1241 ( .A(n943), .B(n942), .Z(n944) );
  AND U1242 ( .A(n945), .B(n944), .Z(n1036) );
  NANDN U1243 ( .A(n947), .B(n946), .Z(n951) );
  NAND U1244 ( .A(n949), .B(n948), .Z(n950) );
  AND U1245 ( .A(n951), .B(n950), .Z(n1035) );
  XOR U1246 ( .A(n1036), .B(n1035), .Z(n1038) );
  XOR U1247 ( .A(n1037), .B(n1038), .Z(n964) );
  NANDN U1248 ( .A(n953), .B(n952), .Z(n957) );
  OR U1249 ( .A(n955), .B(n954), .Z(n956) );
  AND U1250 ( .A(n957), .B(n956), .Z(n963) );
  XNOR U1251 ( .A(n964), .B(n963), .Z(n965) );
  XNOR U1252 ( .A(n966), .B(n965), .Z(n958) );
  XNOR U1253 ( .A(sreg[81]), .B(n958), .Z(n959) );
  XNOR U1254 ( .A(n960), .B(n959), .Z(c[81]) );
  NANDN U1255 ( .A(sreg[81]), .B(n958), .Z(n962) );
  NAND U1256 ( .A(n960), .B(n959), .Z(n961) );
  NAND U1257 ( .A(n962), .B(n961), .Z(n1128) );
  XNOR U1258 ( .A(sreg[82]), .B(n1128), .Z(n1130) );
  NANDN U1259 ( .A(n964), .B(n963), .Z(n968) );
  NANDN U1260 ( .A(n966), .B(n965), .Z(n967) );
  AND U1261 ( .A(n968), .B(n967), .Z(n1043) );
  NANDN U1262 ( .A(n970), .B(n969), .Z(n974) );
  NAND U1263 ( .A(n972), .B(n971), .Z(n973) );
  AND U1264 ( .A(n974), .B(n973), .Z(n1125) );
  NANDN U1265 ( .A(n976), .B(n975), .Z(n980) );
  NANDN U1266 ( .A(n978), .B(n977), .Z(n979) );
  AND U1267 ( .A(n980), .B(n979), .Z(n1122) );
  NANDN U1268 ( .A(n982), .B(n981), .Z(n986) );
  OR U1269 ( .A(n984), .B(n983), .Z(n985) );
  AND U1270 ( .A(n986), .B(n985), .Z(n1117) );
  NANDN U1271 ( .A(n988), .B(n987), .Z(n992) );
  NAND U1272 ( .A(n990), .B(n989), .Z(n991) );
  NAND U1273 ( .A(n992), .B(n991), .Z(n1116) );
  XNOR U1274 ( .A(n1117), .B(n1116), .Z(n1118) );
  NANDN U1275 ( .A(n994), .B(n993), .Z(n998) );
  OR U1276 ( .A(n996), .B(n995), .Z(n997) );
  AND U1277 ( .A(n998), .B(n997), .Z(n1049) );
  NAND U1278 ( .A(b[0]), .B(a[18]), .Z(n999) );
  XNOR U1279 ( .A(b[1]), .B(n999), .Z(n1001) );
  NANDN U1280 ( .A(b[0]), .B(a[17]), .Z(n1000) );
  NAND U1281 ( .A(n1001), .B(n1000), .Z(n1086) );
  XOR U1282 ( .A(b[18]), .B(b[17]), .Z(n33001) );
  IV U1283 ( .A(n33001), .Z(n32823) );
  ANDN U1284 ( .B(a[0]), .A(n32823), .Z(n1083) );
  NANDN U1285 ( .A(n31536), .B(n1002), .Z(n1004) );
  XOR U1286 ( .A(b[15]), .B(a[4]), .Z(n1095) );
  NANDN U1287 ( .A(n31925), .B(n1095), .Z(n1003) );
  AND U1288 ( .A(n1004), .B(n1003), .Z(n1084) );
  XOR U1289 ( .A(n1083), .B(n1084), .Z(n1085) );
  XOR U1290 ( .A(n1086), .B(n1085), .Z(n1048) );
  NOR U1291 ( .A(n1006), .B(n1005), .Z(n1074) );
  NAND U1292 ( .A(n31059), .B(n1007), .Z(n1009) );
  XNOR U1293 ( .A(b[11]), .B(a[8]), .Z(n1107) );
  NANDN U1294 ( .A(n1107), .B(n31060), .Z(n1008) );
  AND U1295 ( .A(n1009), .B(n1008), .Z(n1071) );
  ANDN U1296 ( .B(n1010), .A(n32545), .Z(n32544) );
  NAND U1297 ( .A(n32544), .B(n1011), .Z(n1013) );
  XNOR U1298 ( .A(b[17]), .B(a[2]), .Z(n1058) );
  NANDN U1299 ( .A(n1058), .B(n32545), .Z(n1012) );
  NAND U1300 ( .A(n1013), .B(n1012), .Z(n1072) );
  XNOR U1301 ( .A(n1071), .B(n1072), .Z(n1073) );
  XNOR U1302 ( .A(n1074), .B(n1073), .Z(n1047) );
  XOR U1303 ( .A(n1048), .B(n1047), .Z(n1050) );
  XOR U1304 ( .A(n1049), .B(n1050), .Z(n1113) );
  NANDN U1305 ( .A(n1015), .B(n1014), .Z(n1019) );
  OR U1306 ( .A(n1017), .B(n1016), .Z(n1018) );
  AND U1307 ( .A(n1019), .B(n1018), .Z(n1111) );
  NANDN U1308 ( .A(n28889), .B(n1020), .Z(n1022) );
  XOR U1309 ( .A(b[5]), .B(a[14]), .Z(n1098) );
  NANDN U1310 ( .A(n29138), .B(n1098), .Z(n1021) );
  AND U1311 ( .A(n1022), .B(n1021), .Z(n1078) );
  NANDN U1312 ( .A(n29499), .B(n1023), .Z(n1025) );
  XOR U1313 ( .A(b[7]), .B(a[12]), .Z(n1089) );
  NANDN U1314 ( .A(n29735), .B(n1089), .Z(n1024) );
  NAND U1315 ( .A(n1025), .B(n1024), .Z(n1077) );
  XNOR U1316 ( .A(n1078), .B(n1077), .Z(n1079) );
  NANDN U1317 ( .A(n1026), .B(n30627), .Z(n1028) );
  XOR U1318 ( .A(b[9]), .B(a[10]), .Z(n1062) );
  NANDN U1319 ( .A(n30267), .B(n1062), .Z(n1027) );
  AND U1320 ( .A(n1028), .B(n1027), .Z(n1068) );
  NANDN U1321 ( .A(n31055), .B(n1029), .Z(n1031) );
  XOR U1322 ( .A(b[13]), .B(a[6]), .Z(n1092) );
  NANDN U1323 ( .A(n31293), .B(n1092), .Z(n1030) );
  AND U1324 ( .A(n1031), .B(n1030), .Z(n1066) );
  NANDN U1325 ( .A(n1032), .B(n9942), .Z(n1034) );
  XOR U1326 ( .A(b[3]), .B(a[16]), .Z(n1101) );
  NANDN U1327 ( .A(n28941), .B(n1101), .Z(n1033) );
  NAND U1328 ( .A(n1034), .B(n1033), .Z(n1065) );
  XNOR U1329 ( .A(n1066), .B(n1065), .Z(n1067) );
  XOR U1330 ( .A(n1068), .B(n1067), .Z(n1080) );
  XNOR U1331 ( .A(n1079), .B(n1080), .Z(n1110) );
  XNOR U1332 ( .A(n1111), .B(n1110), .Z(n1112) );
  XOR U1333 ( .A(n1113), .B(n1112), .Z(n1119) );
  XOR U1334 ( .A(n1118), .B(n1119), .Z(n1123) );
  XNOR U1335 ( .A(n1122), .B(n1123), .Z(n1124) );
  XOR U1336 ( .A(n1125), .B(n1124), .Z(n1042) );
  NANDN U1337 ( .A(n1036), .B(n1035), .Z(n1040) );
  OR U1338 ( .A(n1038), .B(n1037), .Z(n1039) );
  AND U1339 ( .A(n1040), .B(n1039), .Z(n1041) );
  XOR U1340 ( .A(n1042), .B(n1041), .Z(n1044) );
  XNOR U1341 ( .A(n1043), .B(n1044), .Z(n1129) );
  XOR U1342 ( .A(n1130), .B(n1129), .Z(c[82]) );
  NANDN U1343 ( .A(n1042), .B(n1041), .Z(n1046) );
  OR U1344 ( .A(n1044), .B(n1043), .Z(n1045) );
  AND U1345 ( .A(n1046), .B(n1045), .Z(n1140) );
  NANDN U1346 ( .A(n1048), .B(n1047), .Z(n1052) );
  OR U1347 ( .A(n1050), .B(n1049), .Z(n1051) );
  AND U1348 ( .A(n1052), .B(n1051), .Z(n1150) );
  XOR U1349 ( .A(b[19]), .B(a[0]), .Z(n1055) );
  XOR U1350 ( .A(b[19]), .B(b[17]), .Z(n1053) );
  XOR U1351 ( .A(b[19]), .B(b[18]), .Z(n1194) );
  AND U1352 ( .A(n1053), .B(n1194), .Z(n1054) );
  NAND U1353 ( .A(n1055), .B(n1054), .Z(n1057) );
  XOR U1354 ( .A(b[19]), .B(a[1]), .Z(n1195) );
  NANDN U1355 ( .A(n32823), .B(n1195), .Z(n1056) );
  AND U1356 ( .A(n1057), .B(n1056), .Z(n1190) );
  NANDN U1357 ( .A(n1058), .B(n32544), .Z(n1060) );
  XOR U1358 ( .A(b[17]), .B(a[3]), .Z(n1162) );
  NANDN U1359 ( .A(n32292), .B(n1162), .Z(n1059) );
  AND U1360 ( .A(n1060), .B(n1059), .Z(n1189) );
  XOR U1361 ( .A(n1190), .B(n1189), .Z(n1179) );
  NAND U1362 ( .A(b[17]), .B(b[18]), .Z(n1061) );
  AND U1363 ( .A(b[19]), .B(n1061), .Z(n33509) );
  ANDN U1364 ( .B(n33509), .A(n1083), .Z(n1178) );
  NAND U1365 ( .A(n30627), .B(n1062), .Z(n1064) );
  XNOR U1366 ( .A(b[9]), .B(a[11]), .Z(n1198) );
  NANDN U1367 ( .A(n1198), .B(n30628), .Z(n1063) );
  AND U1368 ( .A(n1064), .B(n1063), .Z(n1177) );
  XOR U1369 ( .A(n1178), .B(n1177), .Z(n1180) );
  XOR U1370 ( .A(n1179), .B(n1180), .Z(n1208) );
  NANDN U1371 ( .A(n1066), .B(n1065), .Z(n1070) );
  NANDN U1372 ( .A(n1068), .B(n1067), .Z(n1069) );
  NAND U1373 ( .A(n1070), .B(n1069), .Z(n1207) );
  XNOR U1374 ( .A(n1208), .B(n1207), .Z(n1209) );
  NANDN U1375 ( .A(n1072), .B(n1071), .Z(n1076) );
  NANDN U1376 ( .A(n1074), .B(n1073), .Z(n1075) );
  NAND U1377 ( .A(n1076), .B(n1075), .Z(n1210) );
  XOR U1378 ( .A(n1209), .B(n1210), .Z(n1151) );
  XNOR U1379 ( .A(n1150), .B(n1151), .Z(n1153) );
  NANDN U1380 ( .A(n1078), .B(n1077), .Z(n1082) );
  NANDN U1381 ( .A(n1080), .B(n1079), .Z(n1081) );
  AND U1382 ( .A(n1082), .B(n1081), .Z(n1145) );
  NANDN U1383 ( .A(n1084), .B(n1083), .Z(n1088) );
  OR U1384 ( .A(n1086), .B(n1085), .Z(n1087) );
  NAND U1385 ( .A(n1088), .B(n1087), .Z(n1144) );
  XNOR U1386 ( .A(n1145), .B(n1144), .Z(n1146) );
  NANDN U1387 ( .A(n29499), .B(n1089), .Z(n1091) );
  XOR U1388 ( .A(b[7]), .B(a[13]), .Z(n1171) );
  NANDN U1389 ( .A(n29735), .B(n1171), .Z(n1090) );
  AND U1390 ( .A(n1091), .B(n1090), .Z(n1214) );
  NANDN U1391 ( .A(n31055), .B(n1092), .Z(n1094) );
  XOR U1392 ( .A(b[13]), .B(a[7]), .Z(n1204) );
  NANDN U1393 ( .A(n31293), .B(n1204), .Z(n1093) );
  AND U1394 ( .A(n1094), .B(n1093), .Z(n1159) );
  NANDN U1395 ( .A(n31536), .B(n1095), .Z(n1097) );
  XOR U1396 ( .A(b[15]), .B(a[5]), .Z(n1201) );
  NANDN U1397 ( .A(n31925), .B(n1201), .Z(n1096) );
  AND U1398 ( .A(n1097), .B(n1096), .Z(n1157) );
  NANDN U1399 ( .A(n28889), .B(n1098), .Z(n1100) );
  XOR U1400 ( .A(b[5]), .B(a[15]), .Z(n1168) );
  NANDN U1401 ( .A(n29138), .B(n1168), .Z(n1099) );
  NAND U1402 ( .A(n1100), .B(n1099), .Z(n1156) );
  XNOR U1403 ( .A(n1157), .B(n1156), .Z(n1158) );
  XNOR U1404 ( .A(n1159), .B(n1158), .Z(n1213) );
  XNOR U1405 ( .A(n1214), .B(n1213), .Z(n1215) );
  NANDN U1406 ( .A(n209), .B(n1101), .Z(n1103) );
  XOR U1407 ( .A(b[3]), .B(a[17]), .Z(n1174) );
  NANDN U1408 ( .A(n28941), .B(n1174), .Z(n1102) );
  AND U1409 ( .A(n1103), .B(n1102), .Z(n1186) );
  NAND U1410 ( .A(b[0]), .B(a[19]), .Z(n1104) );
  XNOR U1411 ( .A(b[1]), .B(n1104), .Z(n1106) );
  NANDN U1412 ( .A(b[0]), .B(a[18]), .Z(n1105) );
  NAND U1413 ( .A(n1106), .B(n1105), .Z(n1184) );
  NANDN U1414 ( .A(n1107), .B(n31059), .Z(n1109) );
  XOR U1415 ( .A(b[11]), .B(a[9]), .Z(n1191) );
  NANDN U1416 ( .A(n30891), .B(n1191), .Z(n1108) );
  NAND U1417 ( .A(n1109), .B(n1108), .Z(n1183) );
  XNOR U1418 ( .A(n1184), .B(n1183), .Z(n1185) );
  XOR U1419 ( .A(n1186), .B(n1185), .Z(n1216) );
  XOR U1420 ( .A(n1215), .B(n1216), .Z(n1147) );
  XNOR U1421 ( .A(n1146), .B(n1147), .Z(n1152) );
  XOR U1422 ( .A(n1153), .B(n1152), .Z(n1220) );
  NANDN U1423 ( .A(n1111), .B(n1110), .Z(n1115) );
  NANDN U1424 ( .A(n1113), .B(n1112), .Z(n1114) );
  AND U1425 ( .A(n1115), .B(n1114), .Z(n1219) );
  XNOR U1426 ( .A(n1220), .B(n1219), .Z(n1221) );
  NANDN U1427 ( .A(n1117), .B(n1116), .Z(n1121) );
  NANDN U1428 ( .A(n1119), .B(n1118), .Z(n1120) );
  NAND U1429 ( .A(n1121), .B(n1120), .Z(n1222) );
  XNOR U1430 ( .A(n1221), .B(n1222), .Z(n1138) );
  NANDN U1431 ( .A(n1123), .B(n1122), .Z(n1127) );
  NAND U1432 ( .A(n1125), .B(n1124), .Z(n1126) );
  NAND U1433 ( .A(n1127), .B(n1126), .Z(n1139) );
  XOR U1434 ( .A(n1138), .B(n1139), .Z(n1141) );
  XOR U1435 ( .A(n1140), .B(n1141), .Z(n1133) );
  XNOR U1436 ( .A(n1133), .B(sreg[83]), .Z(n1135) );
  NANDN U1437 ( .A(n1128), .B(sreg[82]), .Z(n1132) );
  NAND U1438 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U1439 ( .A(n1132), .B(n1131), .Z(n1134) );
  XOR U1440 ( .A(n1135), .B(n1134), .Z(c[83]) );
  NANDN U1441 ( .A(n1133), .B(sreg[83]), .Z(n1137) );
  NAND U1442 ( .A(n1135), .B(n1134), .Z(n1136) );
  AND U1443 ( .A(n1137), .B(n1136), .Z(n1322) );
  XNOR U1444 ( .A(sreg[84]), .B(n1322), .Z(n1324) );
  NANDN U1445 ( .A(n1139), .B(n1138), .Z(n1143) );
  OR U1446 ( .A(n1141), .B(n1140), .Z(n1142) );
  AND U1447 ( .A(n1143), .B(n1142), .Z(n1228) );
  NANDN U1448 ( .A(n1145), .B(n1144), .Z(n1149) );
  NANDN U1449 ( .A(n1147), .B(n1146), .Z(n1148) );
  AND U1450 ( .A(n1149), .B(n1148), .Z(n1317) );
  NANDN U1451 ( .A(n1151), .B(n1150), .Z(n1155) );
  NAND U1452 ( .A(n1153), .B(n1152), .Z(n1154) );
  NAND U1453 ( .A(n1155), .B(n1154), .Z(n1316) );
  XNOR U1454 ( .A(n1317), .B(n1316), .Z(n1319) );
  NANDN U1455 ( .A(n1157), .B(n1156), .Z(n1161) );
  NANDN U1456 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1457 ( .A(n1161), .B(n1160), .Z(n1300) );
  XOR U1458 ( .A(b[20]), .B(b[19]), .Z(n33414) );
  IV U1459 ( .A(n33414), .Z(n33271) );
  ANDN U1460 ( .B(a[0]), .A(n33271), .Z(n1246) );
  IV U1461 ( .A(n32544), .Z(n32013) );
  NANDN U1462 ( .A(n32013), .B(n1162), .Z(n1164) );
  XOR U1463 ( .A(b[17]), .B(a[4]), .Z(n1274) );
  NANDN U1464 ( .A(n32292), .B(n1274), .Z(n1163) );
  AND U1465 ( .A(n1164), .B(n1163), .Z(n1231) );
  XNOR U1466 ( .A(n1246), .B(n1231), .Z(n1232) );
  NAND U1467 ( .A(b[0]), .B(a[20]), .Z(n1165) );
  XNOR U1468 ( .A(b[1]), .B(n1165), .Z(n1167) );
  NANDN U1469 ( .A(b[0]), .B(a[19]), .Z(n1166) );
  NAND U1470 ( .A(n1167), .B(n1166), .Z(n1233) );
  XNOR U1471 ( .A(n1232), .B(n1233), .Z(n1298) );
  NANDN U1472 ( .A(n28889), .B(n1168), .Z(n1170) );
  XOR U1473 ( .A(b[5]), .B(a[16]), .Z(n1268) );
  NANDN U1474 ( .A(n29138), .B(n1268), .Z(n1169) );
  AND U1475 ( .A(n1170), .B(n1169), .Z(n1295) );
  NANDN U1476 ( .A(n29499), .B(n1171), .Z(n1173) );
  XOR U1477 ( .A(b[7]), .B(a[14]), .Z(n1265) );
  NANDN U1478 ( .A(n29735), .B(n1265), .Z(n1172) );
  AND U1479 ( .A(n1173), .B(n1172), .Z(n1293) );
  NANDN U1480 ( .A(n209), .B(n1174), .Z(n1176) );
  XOR U1481 ( .A(b[3]), .B(a[18]), .Z(n1250) );
  NANDN U1482 ( .A(n28941), .B(n1250), .Z(n1175) );
  NAND U1483 ( .A(n1176), .B(n1175), .Z(n1292) );
  XNOR U1484 ( .A(n1293), .B(n1292), .Z(n1294) );
  XOR U1485 ( .A(n1295), .B(n1294), .Z(n1299) );
  XOR U1486 ( .A(n1298), .B(n1299), .Z(n1301) );
  XOR U1487 ( .A(n1300), .B(n1301), .Z(n1306) );
  NANDN U1488 ( .A(n1178), .B(n1177), .Z(n1182) );
  OR U1489 ( .A(n1180), .B(n1179), .Z(n1181) );
  AND U1490 ( .A(n1182), .B(n1181), .Z(n1305) );
  NANDN U1491 ( .A(n1184), .B(n1183), .Z(n1188) );
  NANDN U1492 ( .A(n1186), .B(n1185), .Z(n1187) );
  AND U1493 ( .A(n1188), .B(n1187), .Z(n1282) );
  NOR U1494 ( .A(n1190), .B(n1189), .Z(n1261) );
  NAND U1495 ( .A(n31059), .B(n1191), .Z(n1193) );
  XNOR U1496 ( .A(b[11]), .B(a[10]), .Z(n1247) );
  NANDN U1497 ( .A(n1247), .B(n31060), .Z(n1192) );
  AND U1498 ( .A(n1193), .B(n1192), .Z(n1259) );
  ANDN U1499 ( .B(n1194), .A(n33001), .Z(n33000) );
  NAND U1500 ( .A(n33000), .B(n1195), .Z(n1197) );
  XNOR U1501 ( .A(b[19]), .B(a[2]), .Z(n1236) );
  NANDN U1502 ( .A(n1236), .B(n33001), .Z(n1196) );
  NAND U1503 ( .A(n1197), .B(n1196), .Z(n1260) );
  XOR U1504 ( .A(n1259), .B(n1260), .Z(n1262) );
  XOR U1505 ( .A(n1261), .B(n1262), .Z(n1281) );
  NANDN U1506 ( .A(n1198), .B(n30627), .Z(n1200) );
  XNOR U1507 ( .A(b[9]), .B(a[12]), .Z(n1256) );
  NANDN U1508 ( .A(n1256), .B(n30628), .Z(n1199) );
  NAND U1509 ( .A(n1200), .B(n1199), .Z(n1287) );
  NANDN U1510 ( .A(n31536), .B(n1201), .Z(n1203) );
  XOR U1511 ( .A(b[15]), .B(a[6]), .Z(n1277) );
  NANDN U1512 ( .A(n31925), .B(n1277), .Z(n1202) );
  NAND U1513 ( .A(n1203), .B(n1202), .Z(n1286) );
  XOR U1514 ( .A(n1287), .B(n1286), .Z(n1289) );
  NAND U1515 ( .A(n31507), .B(n1204), .Z(n1206) );
  XNOR U1516 ( .A(b[13]), .B(a[8]), .Z(n1271) );
  NANDN U1517 ( .A(n1271), .B(n31508), .Z(n1205) );
  NAND U1518 ( .A(n1206), .B(n1205), .Z(n1288) );
  XOR U1519 ( .A(n1289), .B(n1288), .Z(n1280) );
  XOR U1520 ( .A(n1281), .B(n1280), .Z(n1283) );
  XNOR U1521 ( .A(n1282), .B(n1283), .Z(n1304) );
  XOR U1522 ( .A(n1305), .B(n1304), .Z(n1307) );
  XOR U1523 ( .A(n1306), .B(n1307), .Z(n1313) );
  NANDN U1524 ( .A(n1208), .B(n1207), .Z(n1212) );
  NANDN U1525 ( .A(n1210), .B(n1209), .Z(n1211) );
  AND U1526 ( .A(n1212), .B(n1211), .Z(n1311) );
  NANDN U1527 ( .A(n1214), .B(n1213), .Z(n1218) );
  NANDN U1528 ( .A(n1216), .B(n1215), .Z(n1217) );
  NAND U1529 ( .A(n1218), .B(n1217), .Z(n1310) );
  XNOR U1530 ( .A(n1311), .B(n1310), .Z(n1312) );
  XNOR U1531 ( .A(n1313), .B(n1312), .Z(n1318) );
  XOR U1532 ( .A(n1319), .B(n1318), .Z(n1226) );
  NANDN U1533 ( .A(n1220), .B(n1219), .Z(n1224) );
  NANDN U1534 ( .A(n1222), .B(n1221), .Z(n1223) );
  NAND U1535 ( .A(n1224), .B(n1223), .Z(n1225) );
  XNOR U1536 ( .A(n1226), .B(n1225), .Z(n1227) );
  XNOR U1537 ( .A(n1228), .B(n1227), .Z(n1323) );
  XNOR U1538 ( .A(n1324), .B(n1323), .Z(c[84]) );
  NANDN U1539 ( .A(n1226), .B(n1225), .Z(n1230) );
  NANDN U1540 ( .A(n1228), .B(n1227), .Z(n1229) );
  AND U1541 ( .A(n1230), .B(n1229), .Z(n1334) );
  NANDN U1542 ( .A(n1231), .B(n1246), .Z(n1235) );
  NANDN U1543 ( .A(n1233), .B(n1232), .Z(n1234) );
  NAND U1544 ( .A(n1235), .B(n1234), .Z(n1350) );
  NANDN U1545 ( .A(n1236), .B(n33000), .Z(n1238) );
  XOR U1546 ( .A(b[19]), .B(a[3]), .Z(n1383) );
  NANDN U1547 ( .A(n32823), .B(n1383), .Z(n1237) );
  AND U1548 ( .A(n1238), .B(n1237), .Z(n1378) );
  XOR U1549 ( .A(b[21]), .B(a[1]), .Z(n1399) );
  NANDN U1550 ( .A(n33271), .B(n1399), .Z(n1245) );
  ANDN U1551 ( .B(b[20]), .A(b[21]), .Z(n1239) );
  NAND U1552 ( .A(n1239), .B(a[0]), .Z(n1242) );
  NAND U1553 ( .A(b[19]), .B(b[20]), .Z(n1240) );
  NAND U1554 ( .A(b[21]), .B(n1240), .Z(n33775) );
  OR U1555 ( .A(a[0]), .B(n33775), .Z(n1241) );
  NAND U1556 ( .A(n1242), .B(n1241), .Z(n1243) );
  NAND U1557 ( .A(n33271), .B(n1243), .Z(n1244) );
  AND U1558 ( .A(n1245), .B(n1244), .Z(n1379) );
  XOR U1559 ( .A(n1378), .B(n1379), .Z(n1369) );
  NOR U1560 ( .A(n33775), .B(n1246), .Z(n1367) );
  NANDN U1561 ( .A(n1247), .B(n31059), .Z(n1249) );
  XNOR U1562 ( .A(b[11]), .B(a[11]), .Z(n1405) );
  NANDN U1563 ( .A(n1405), .B(n31060), .Z(n1248) );
  AND U1564 ( .A(n1249), .B(n1248), .Z(n1366) );
  XNOR U1565 ( .A(n1367), .B(n1366), .Z(n1368) );
  XOR U1566 ( .A(n1369), .B(n1368), .Z(n1348) );
  NANDN U1567 ( .A(n209), .B(n1250), .Z(n1252) );
  XOR U1568 ( .A(b[3]), .B(a[19]), .Z(n1372) );
  NANDN U1569 ( .A(n28941), .B(n1372), .Z(n1251) );
  AND U1570 ( .A(n1252), .B(n1251), .Z(n1416) );
  NAND U1571 ( .A(b[0]), .B(a[21]), .Z(n1253) );
  XNOR U1572 ( .A(b[1]), .B(n1253), .Z(n1255) );
  NANDN U1573 ( .A(b[0]), .B(a[20]), .Z(n1254) );
  NAND U1574 ( .A(n1255), .B(n1254), .Z(n1415) );
  NANDN U1575 ( .A(n1256), .B(n30627), .Z(n1258) );
  XOR U1576 ( .A(b[9]), .B(a[13]), .Z(n1402) );
  NANDN U1577 ( .A(n30267), .B(n1402), .Z(n1257) );
  NAND U1578 ( .A(n1258), .B(n1257), .Z(n1414) );
  XOR U1579 ( .A(n1415), .B(n1414), .Z(n1417) );
  XOR U1580 ( .A(n1416), .B(n1417), .Z(n1349) );
  XOR U1581 ( .A(n1348), .B(n1349), .Z(n1351) );
  XNOR U1582 ( .A(n1350), .B(n1351), .Z(n1356) );
  NANDN U1583 ( .A(n1260), .B(n1259), .Z(n1264) );
  OR U1584 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U1585 ( .A(n1264), .B(n1263), .Z(n1355) );
  NANDN U1586 ( .A(n29499), .B(n1265), .Z(n1267) );
  XOR U1587 ( .A(b[7]), .B(a[15]), .Z(n1386) );
  NANDN U1588 ( .A(n29735), .B(n1386), .Z(n1266) );
  AND U1589 ( .A(n1267), .B(n1266), .Z(n1361) );
  NANDN U1590 ( .A(n28889), .B(n1268), .Z(n1270) );
  XOR U1591 ( .A(b[5]), .B(a[17]), .Z(n1389) );
  NANDN U1592 ( .A(n29138), .B(n1389), .Z(n1269) );
  NAND U1593 ( .A(n1270), .B(n1269), .Z(n1360) );
  XNOR U1594 ( .A(n1361), .B(n1360), .Z(n1363) );
  NANDN U1595 ( .A(n1271), .B(n31507), .Z(n1273) );
  XOR U1596 ( .A(b[13]), .B(a[9]), .Z(n1375) );
  NANDN U1597 ( .A(n31293), .B(n1375), .Z(n1272) );
  AND U1598 ( .A(n1273), .B(n1272), .Z(n1411) );
  NANDN U1599 ( .A(n32013), .B(n1274), .Z(n1276) );
  XOR U1600 ( .A(b[17]), .B(a[5]), .Z(n1395) );
  NANDN U1601 ( .A(n32292), .B(n1395), .Z(n1275) );
  AND U1602 ( .A(n1276), .B(n1275), .Z(n1409) );
  NANDN U1603 ( .A(n31536), .B(n1277), .Z(n1279) );
  XOR U1604 ( .A(b[15]), .B(a[7]), .Z(n1392) );
  NANDN U1605 ( .A(n31925), .B(n1392), .Z(n1278) );
  NAND U1606 ( .A(n1279), .B(n1278), .Z(n1408) );
  XNOR U1607 ( .A(n1409), .B(n1408), .Z(n1410) );
  XNOR U1608 ( .A(n1411), .B(n1410), .Z(n1362) );
  XNOR U1609 ( .A(n1363), .B(n1362), .Z(n1354) );
  XOR U1610 ( .A(n1355), .B(n1354), .Z(n1357) );
  XOR U1611 ( .A(n1356), .B(n1357), .Z(n1338) );
  NANDN U1612 ( .A(n1281), .B(n1280), .Z(n1285) );
  OR U1613 ( .A(n1283), .B(n1282), .Z(n1284) );
  NAND U1614 ( .A(n1285), .B(n1284), .Z(n1339) );
  XOR U1615 ( .A(n1338), .B(n1339), .Z(n1341) );
  NAND U1616 ( .A(n1287), .B(n1286), .Z(n1291) );
  NAND U1617 ( .A(n1289), .B(n1288), .Z(n1290) );
  NAND U1618 ( .A(n1291), .B(n1290), .Z(n1343) );
  NANDN U1619 ( .A(n1293), .B(n1292), .Z(n1297) );
  NANDN U1620 ( .A(n1295), .B(n1294), .Z(n1296) );
  NAND U1621 ( .A(n1297), .B(n1296), .Z(n1342) );
  XOR U1622 ( .A(n1343), .B(n1342), .Z(n1345) );
  NANDN U1623 ( .A(n1299), .B(n1298), .Z(n1303) );
  OR U1624 ( .A(n1301), .B(n1300), .Z(n1302) );
  NAND U1625 ( .A(n1303), .B(n1302), .Z(n1344) );
  XOR U1626 ( .A(n1345), .B(n1344), .Z(n1340) );
  XOR U1627 ( .A(n1341), .B(n1340), .Z(n1421) );
  NANDN U1628 ( .A(n1305), .B(n1304), .Z(n1309) );
  OR U1629 ( .A(n1307), .B(n1306), .Z(n1308) );
  NAND U1630 ( .A(n1309), .B(n1308), .Z(n1420) );
  XNOR U1631 ( .A(n1421), .B(n1420), .Z(n1422) );
  NANDN U1632 ( .A(n1311), .B(n1310), .Z(n1315) );
  NANDN U1633 ( .A(n1313), .B(n1312), .Z(n1314) );
  NAND U1634 ( .A(n1315), .B(n1314), .Z(n1423) );
  XNOR U1635 ( .A(n1422), .B(n1423), .Z(n1332) );
  NANDN U1636 ( .A(n1317), .B(n1316), .Z(n1321) );
  NAND U1637 ( .A(n1319), .B(n1318), .Z(n1320) );
  NAND U1638 ( .A(n1321), .B(n1320), .Z(n1333) );
  XOR U1639 ( .A(n1332), .B(n1333), .Z(n1335) );
  XOR U1640 ( .A(n1334), .B(n1335), .Z(n1327) );
  XNOR U1641 ( .A(n1327), .B(sreg[85]), .Z(n1329) );
  NANDN U1642 ( .A(sreg[84]), .B(n1322), .Z(n1326) );
  NAND U1643 ( .A(n1324), .B(n1323), .Z(n1325) );
  AND U1644 ( .A(n1326), .B(n1325), .Z(n1328) );
  XOR U1645 ( .A(n1329), .B(n1328), .Z(c[85]) );
  NANDN U1646 ( .A(n1327), .B(sreg[85]), .Z(n1331) );
  NAND U1647 ( .A(n1329), .B(n1328), .Z(n1330) );
  AND U1648 ( .A(n1331), .B(n1330), .Z(n1530) );
  XNOR U1649 ( .A(sreg[86]), .B(n1530), .Z(n1532) );
  NANDN U1650 ( .A(n1333), .B(n1332), .Z(n1337) );
  OR U1651 ( .A(n1335), .B(n1334), .Z(n1336) );
  AND U1652 ( .A(n1337), .B(n1336), .Z(n1429) );
  NAND U1653 ( .A(n1343), .B(n1342), .Z(n1347) );
  NAND U1654 ( .A(n1345), .B(n1344), .Z(n1346) );
  NAND U1655 ( .A(n1347), .B(n1346), .Z(n1524) );
  XNOR U1656 ( .A(n1525), .B(n1524), .Z(n1527) );
  NAND U1657 ( .A(n1349), .B(n1348), .Z(n1353) );
  NAND U1658 ( .A(n1351), .B(n1350), .Z(n1352) );
  AND U1659 ( .A(n1353), .B(n1352), .Z(n1433) );
  NANDN U1660 ( .A(n1355), .B(n1354), .Z(n1359) );
  NANDN U1661 ( .A(n1357), .B(n1356), .Z(n1358) );
  AND U1662 ( .A(n1359), .B(n1358), .Z(n1432) );
  XNOR U1663 ( .A(n1433), .B(n1432), .Z(n1434) );
  NANDN U1664 ( .A(n1361), .B(n1360), .Z(n1365) );
  NAND U1665 ( .A(n1363), .B(n1362), .Z(n1364) );
  AND U1666 ( .A(n1365), .B(n1364), .Z(n1439) );
  NANDN U1667 ( .A(n1367), .B(n1366), .Z(n1371) );
  NANDN U1668 ( .A(n1369), .B(n1368), .Z(n1370) );
  AND U1669 ( .A(n1371), .B(n1370), .Z(n1446) );
  NANDN U1670 ( .A(n209), .B(n1372), .Z(n1374) );
  XOR U1671 ( .A(b[3]), .B(a[20]), .Z(n1467) );
  NANDN U1672 ( .A(n28941), .B(n1467), .Z(n1373) );
  AND U1673 ( .A(n1374), .B(n1373), .Z(n1507) );
  NANDN U1674 ( .A(n31055), .B(n1375), .Z(n1377) );
  XOR U1675 ( .A(b[13]), .B(a[10]), .Z(n1481) );
  NANDN U1676 ( .A(n31293), .B(n1481), .Z(n1376) );
  NAND U1677 ( .A(n1377), .B(n1376), .Z(n1506) );
  XNOR U1678 ( .A(n1507), .B(n1506), .Z(n1509) );
  NOR U1679 ( .A(n1379), .B(n1378), .Z(n1508) );
  XOR U1680 ( .A(n1509), .B(n1508), .Z(n1445) );
  NAND U1681 ( .A(b[0]), .B(a[22]), .Z(n1380) );
  XNOR U1682 ( .A(b[1]), .B(n1380), .Z(n1382) );
  NANDN U1683 ( .A(b[0]), .B(a[21]), .Z(n1381) );
  NAND U1684 ( .A(n1382), .B(n1381), .Z(n1464) );
  XOR U1685 ( .A(b[22]), .B(b[21]), .Z(n33868) );
  IV U1686 ( .A(n33868), .Z(n33644) );
  ANDN U1687 ( .B(a[0]), .A(n33644), .Z(n1474) );
  IV U1688 ( .A(n33000), .Z(n32483) );
  NANDN U1689 ( .A(n32483), .B(n1383), .Z(n1385) );
  XOR U1690 ( .A(b[19]), .B(a[4]), .Z(n1478) );
  NANDN U1691 ( .A(n32823), .B(n1478), .Z(n1384) );
  AND U1692 ( .A(n1385), .B(n1384), .Z(n1462) );
  XOR U1693 ( .A(n1474), .B(n1462), .Z(n1463) );
  XNOR U1694 ( .A(n1464), .B(n1463), .Z(n1444) );
  XOR U1695 ( .A(n1445), .B(n1444), .Z(n1447) );
  XNOR U1696 ( .A(n1446), .B(n1447), .Z(n1438) );
  XNOR U1697 ( .A(n1439), .B(n1438), .Z(n1440) );
  NANDN U1698 ( .A(n29499), .B(n1386), .Z(n1388) );
  XOR U1699 ( .A(b[7]), .B(a[16]), .Z(n1497) );
  NANDN U1700 ( .A(n29735), .B(n1497), .Z(n1387) );
  AND U1701 ( .A(n1388), .B(n1387), .Z(n1520) );
  NANDN U1702 ( .A(n28889), .B(n1389), .Z(n1391) );
  XOR U1703 ( .A(b[5]), .B(a[18]), .Z(n1503) );
  NANDN U1704 ( .A(n29138), .B(n1503), .Z(n1390) );
  AND U1705 ( .A(n1391), .B(n1390), .Z(n1519) );
  NANDN U1706 ( .A(n31536), .B(n1392), .Z(n1394) );
  XOR U1707 ( .A(b[15]), .B(a[8]), .Z(n1470) );
  NANDN U1708 ( .A(n31925), .B(n1470), .Z(n1393) );
  NAND U1709 ( .A(n1394), .B(n1393), .Z(n1518) );
  XOR U1710 ( .A(n1519), .B(n1518), .Z(n1521) );
  XOR U1711 ( .A(n1520), .B(n1521), .Z(n1458) );
  NANDN U1712 ( .A(n32013), .B(n1395), .Z(n1397) );
  XOR U1713 ( .A(b[17]), .B(a[6]), .Z(n1475) );
  NANDN U1714 ( .A(n32292), .B(n1475), .Z(n1396) );
  AND U1715 ( .A(n1397), .B(n1396), .Z(n1514) );
  XOR U1716 ( .A(b[20]), .B(b[21]), .Z(n1398) );
  ANDN U1717 ( .B(n1398), .A(n33414), .Z(n33413) );
  IV U1718 ( .A(n33413), .Z(n32996) );
  NANDN U1719 ( .A(n32996), .B(n1399), .Z(n1401) );
  XOR U1720 ( .A(b[21]), .B(a[2]), .Z(n1490) );
  NANDN U1721 ( .A(n33271), .B(n1490), .Z(n1400) );
  AND U1722 ( .A(n1401), .B(n1400), .Z(n1513) );
  NANDN U1723 ( .A(n210), .B(n1402), .Z(n1404) );
  XOR U1724 ( .A(b[9]), .B(a[14]), .Z(n1500) );
  NANDN U1725 ( .A(n30267), .B(n1500), .Z(n1403) );
  NAND U1726 ( .A(n1404), .B(n1403), .Z(n1512) );
  XOR U1727 ( .A(n1513), .B(n1512), .Z(n1515) );
  XOR U1728 ( .A(n1514), .B(n1515), .Z(n1457) );
  NANDN U1729 ( .A(n1405), .B(n31059), .Z(n1407) );
  XNOR U1730 ( .A(b[11]), .B(a[12]), .Z(n1487) );
  NANDN U1731 ( .A(n1487), .B(n31060), .Z(n1406) );
  AND U1732 ( .A(n1407), .B(n1406), .Z(n1456) );
  XOR U1733 ( .A(n1457), .B(n1456), .Z(n1459) );
  XOR U1734 ( .A(n1458), .B(n1459), .Z(n1453) );
  NANDN U1735 ( .A(n1409), .B(n1408), .Z(n1413) );
  NANDN U1736 ( .A(n1411), .B(n1410), .Z(n1412) );
  AND U1737 ( .A(n1413), .B(n1412), .Z(n1451) );
  NANDN U1738 ( .A(n1415), .B(n1414), .Z(n1419) );
  OR U1739 ( .A(n1417), .B(n1416), .Z(n1418) );
  NAND U1740 ( .A(n1419), .B(n1418), .Z(n1450) );
  XNOR U1741 ( .A(n1451), .B(n1450), .Z(n1452) );
  XOR U1742 ( .A(n1453), .B(n1452), .Z(n1441) );
  XOR U1743 ( .A(n1440), .B(n1441), .Z(n1435) );
  XNOR U1744 ( .A(n1434), .B(n1435), .Z(n1526) );
  XOR U1745 ( .A(n1527), .B(n1526), .Z(n1427) );
  NANDN U1746 ( .A(n1421), .B(n1420), .Z(n1425) );
  NANDN U1747 ( .A(n1423), .B(n1422), .Z(n1424) );
  NAND U1748 ( .A(n1425), .B(n1424), .Z(n1426) );
  XNOR U1749 ( .A(n1427), .B(n1426), .Z(n1428) );
  XNOR U1750 ( .A(n1429), .B(n1428), .Z(n1531) );
  XNOR U1751 ( .A(n1532), .B(n1531), .Z(c[86]) );
  NANDN U1752 ( .A(n1427), .B(n1426), .Z(n1431) );
  NANDN U1753 ( .A(n1429), .B(n1428), .Z(n1430) );
  AND U1754 ( .A(n1431), .B(n1430), .Z(n1543) );
  NANDN U1755 ( .A(n1433), .B(n1432), .Z(n1437) );
  NANDN U1756 ( .A(n1435), .B(n1434), .Z(n1436) );
  AND U1757 ( .A(n1437), .B(n1436), .Z(n1641) );
  NANDN U1758 ( .A(n1439), .B(n1438), .Z(n1443) );
  NANDN U1759 ( .A(n1441), .B(n1440), .Z(n1442) );
  AND U1760 ( .A(n1443), .B(n1442), .Z(n1549) );
  NANDN U1761 ( .A(n1445), .B(n1444), .Z(n1449) );
  OR U1762 ( .A(n1447), .B(n1446), .Z(n1448) );
  AND U1763 ( .A(n1449), .B(n1448), .Z(n1547) );
  NANDN U1764 ( .A(n1451), .B(n1450), .Z(n1455) );
  NANDN U1765 ( .A(n1453), .B(n1452), .Z(n1454) );
  AND U1766 ( .A(n1455), .B(n1454), .Z(n1546) );
  XNOR U1767 ( .A(n1547), .B(n1546), .Z(n1548) );
  XOR U1768 ( .A(n1549), .B(n1548), .Z(n1640) );
  NANDN U1769 ( .A(n1457), .B(n1456), .Z(n1461) );
  OR U1770 ( .A(n1459), .B(n1458), .Z(n1460) );
  AND U1771 ( .A(n1461), .B(n1460), .Z(n1552) );
  NANDN U1772 ( .A(n1462), .B(n1474), .Z(n1466) );
  OR U1773 ( .A(n1464), .B(n1463), .Z(n1465) );
  AND U1774 ( .A(n1466), .B(n1465), .Z(n1636) );
  NANDN U1775 ( .A(n209), .B(n1467), .Z(n1469) );
  XOR U1776 ( .A(b[3]), .B(a[21]), .Z(n1575) );
  NANDN U1777 ( .A(n28941), .B(n1575), .Z(n1468) );
  AND U1778 ( .A(n1469), .B(n1468), .Z(n1587) );
  NANDN U1779 ( .A(n31536), .B(n1470), .Z(n1472) );
  XOR U1780 ( .A(b[15]), .B(a[9]), .Z(n1611) );
  NANDN U1781 ( .A(n31925), .B(n1611), .Z(n1471) );
  AND U1782 ( .A(n1472), .B(n1471), .Z(n1585) );
  NAND U1783 ( .A(b[21]), .B(b[22]), .Z(n1473) );
  AND U1784 ( .A(b[23]), .B(n1473), .Z(n34267) );
  ANDN U1785 ( .B(n34267), .A(n1474), .Z(n1584) );
  XNOR U1786 ( .A(n1585), .B(n1584), .Z(n1586) );
  XNOR U1787 ( .A(n1587), .B(n1586), .Z(n1633) );
  NANDN U1788 ( .A(n32013), .B(n1475), .Z(n1477) );
  XOR U1789 ( .A(b[17]), .B(a[7]), .Z(n1608) );
  NANDN U1790 ( .A(n32292), .B(n1608), .Z(n1476) );
  AND U1791 ( .A(n1477), .B(n1476), .Z(n1567) );
  NANDN U1792 ( .A(n32483), .B(n1478), .Z(n1480) );
  XOR U1793 ( .A(b[19]), .B(a[5]), .Z(n1617) );
  NANDN U1794 ( .A(n32823), .B(n1617), .Z(n1479) );
  AND U1795 ( .A(n1480), .B(n1479), .Z(n1565) );
  NANDN U1796 ( .A(n31055), .B(n1481), .Z(n1483) );
  XOR U1797 ( .A(b[13]), .B(a[11]), .Z(n1572) );
  NANDN U1798 ( .A(n31293), .B(n1572), .Z(n1482) );
  NAND U1799 ( .A(n1483), .B(n1482), .Z(n1564) );
  XNOR U1800 ( .A(n1565), .B(n1564), .Z(n1566) );
  XOR U1801 ( .A(n1567), .B(n1566), .Z(n1634) );
  XNOR U1802 ( .A(n1633), .B(n1634), .Z(n1635) );
  XOR U1803 ( .A(n1636), .B(n1635), .Z(n1553) );
  XNOR U1804 ( .A(n1552), .B(n1553), .Z(n1554) );
  NAND U1805 ( .A(b[0]), .B(a[23]), .Z(n1484) );
  XNOR U1806 ( .A(b[1]), .B(n1484), .Z(n1486) );
  NANDN U1807 ( .A(b[0]), .B(a[22]), .Z(n1485) );
  NAND U1808 ( .A(n1486), .B(n1485), .Z(n1579) );
  NANDN U1809 ( .A(n1487), .B(n31059), .Z(n1489) );
  XOR U1810 ( .A(b[11]), .B(a[13]), .Z(n1614) );
  NANDN U1811 ( .A(n30891), .B(n1614), .Z(n1488) );
  NAND U1812 ( .A(n1489), .B(n1488), .Z(n1578) );
  XNOR U1813 ( .A(n1579), .B(n1578), .Z(n1580) );
  NANDN U1814 ( .A(n32996), .B(n1490), .Z(n1492) );
  XOR U1815 ( .A(b[21]), .B(a[3]), .Z(n1599) );
  NANDN U1816 ( .A(n33271), .B(n1599), .Z(n1491) );
  AND U1817 ( .A(n1492), .B(n1491), .Z(n1570) );
  XOR U1818 ( .A(b[23]), .B(b[22]), .Z(n1620) );
  XOR U1819 ( .A(b[23]), .B(a[0]), .Z(n1493) );
  NAND U1820 ( .A(n1620), .B(n1493), .Z(n1494) );
  OR U1821 ( .A(n1494), .B(n33868), .Z(n1496) );
  XOR U1822 ( .A(b[23]), .B(a[1]), .Z(n1621) );
  NAND U1823 ( .A(n33868), .B(n1621), .Z(n1495) );
  NAND U1824 ( .A(n1496), .B(n1495), .Z(n1571) );
  XOR U1825 ( .A(n1570), .B(n1571), .Z(n1581) );
  XNOR U1826 ( .A(n1580), .B(n1581), .Z(n1628) );
  NANDN U1827 ( .A(n29499), .B(n1497), .Z(n1499) );
  XOR U1828 ( .A(b[7]), .B(a[17]), .Z(n1602) );
  NANDN U1829 ( .A(n29735), .B(n1602), .Z(n1498) );
  AND U1830 ( .A(n1499), .B(n1498), .Z(n1592) );
  NANDN U1831 ( .A(n210), .B(n1500), .Z(n1502) );
  XOR U1832 ( .A(b[9]), .B(a[15]), .Z(n1624) );
  NANDN U1833 ( .A(n30267), .B(n1624), .Z(n1501) );
  AND U1834 ( .A(n1502), .B(n1501), .Z(n1591) );
  NANDN U1835 ( .A(n28889), .B(n1503), .Z(n1505) );
  XOR U1836 ( .A(b[5]), .B(a[19]), .Z(n1605) );
  NANDN U1837 ( .A(n29138), .B(n1605), .Z(n1504) );
  NAND U1838 ( .A(n1505), .B(n1504), .Z(n1590) );
  XOR U1839 ( .A(n1591), .B(n1590), .Z(n1593) );
  XOR U1840 ( .A(n1592), .B(n1593), .Z(n1627) );
  XOR U1841 ( .A(n1628), .B(n1627), .Z(n1630) );
  NANDN U1842 ( .A(n1507), .B(n1506), .Z(n1511) );
  NAND U1843 ( .A(n1509), .B(n1508), .Z(n1510) );
  NAND U1844 ( .A(n1511), .B(n1510), .Z(n1629) );
  XOR U1845 ( .A(n1630), .B(n1629), .Z(n1560) );
  NANDN U1846 ( .A(n1513), .B(n1512), .Z(n1517) );
  OR U1847 ( .A(n1515), .B(n1514), .Z(n1516) );
  AND U1848 ( .A(n1517), .B(n1516), .Z(n1559) );
  NANDN U1849 ( .A(n1519), .B(n1518), .Z(n1523) );
  OR U1850 ( .A(n1521), .B(n1520), .Z(n1522) );
  NAND U1851 ( .A(n1523), .B(n1522), .Z(n1558) );
  XOR U1852 ( .A(n1559), .B(n1558), .Z(n1561) );
  XOR U1853 ( .A(n1560), .B(n1561), .Z(n1555) );
  XNOR U1854 ( .A(n1554), .B(n1555), .Z(n1639) );
  XOR U1855 ( .A(n1640), .B(n1639), .Z(n1642) );
  XOR U1856 ( .A(n1641), .B(n1642), .Z(n1541) );
  NANDN U1857 ( .A(n1525), .B(n1524), .Z(n1529) );
  NAND U1858 ( .A(n1527), .B(n1526), .Z(n1528) );
  AND U1859 ( .A(n1529), .B(n1528), .Z(n1540) );
  XNOR U1860 ( .A(n1541), .B(n1540), .Z(n1542) );
  XNOR U1861 ( .A(n1543), .B(n1542), .Z(n1535) );
  XNOR U1862 ( .A(sreg[87]), .B(n1535), .Z(n1537) );
  NANDN U1863 ( .A(sreg[86]), .B(n1530), .Z(n1534) );
  NAND U1864 ( .A(n1532), .B(n1531), .Z(n1533) );
  NAND U1865 ( .A(n1534), .B(n1533), .Z(n1536) );
  XNOR U1866 ( .A(n1537), .B(n1536), .Z(c[87]) );
  NANDN U1867 ( .A(sreg[87]), .B(n1535), .Z(n1539) );
  NAND U1868 ( .A(n1537), .B(n1536), .Z(n1538) );
  NAND U1869 ( .A(n1539), .B(n1538), .Z(n1757) );
  XNOR U1870 ( .A(sreg[88]), .B(n1757), .Z(n1759) );
  NANDN U1871 ( .A(n1541), .B(n1540), .Z(n1545) );
  NANDN U1872 ( .A(n1543), .B(n1542), .Z(n1544) );
  AND U1873 ( .A(n1545), .B(n1544), .Z(n1648) );
  NANDN U1874 ( .A(n1547), .B(n1546), .Z(n1551) );
  NAND U1875 ( .A(n1549), .B(n1548), .Z(n1550) );
  AND U1876 ( .A(n1551), .B(n1550), .Z(n1654) );
  NANDN U1877 ( .A(n1553), .B(n1552), .Z(n1557) );
  NANDN U1878 ( .A(n1555), .B(n1554), .Z(n1556) );
  AND U1879 ( .A(n1557), .B(n1556), .Z(n1651) );
  NANDN U1880 ( .A(n1559), .B(n1558), .Z(n1563) );
  NANDN U1881 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U1882 ( .A(n1563), .B(n1562), .Z(n1753) );
  NANDN U1883 ( .A(n1565), .B(n1564), .Z(n1569) );
  NANDN U1884 ( .A(n1567), .B(n1566), .Z(n1568) );
  AND U1885 ( .A(n1569), .B(n1568), .Z(n1667) );
  ANDN U1886 ( .B(n1571), .A(n1570), .Z(n1711) );
  NAND U1887 ( .A(n31507), .B(n1572), .Z(n1574) );
  XNOR U1888 ( .A(b[13]), .B(a[12]), .Z(n1697) );
  NANDN U1889 ( .A(n1697), .B(n31508), .Z(n1573) );
  AND U1890 ( .A(n1574), .B(n1573), .Z(n1708) );
  NAND U1891 ( .A(n9942), .B(n1575), .Z(n1577) );
  XNOR U1892 ( .A(b[3]), .B(a[22]), .Z(n1700) );
  NANDN U1893 ( .A(n1700), .B(n9653), .Z(n1576) );
  NAND U1894 ( .A(n1577), .B(n1576), .Z(n1709) );
  XNOR U1895 ( .A(n1708), .B(n1709), .Z(n1710) );
  XOR U1896 ( .A(n1711), .B(n1710), .Z(n1668) );
  XNOR U1897 ( .A(n1667), .B(n1668), .Z(n1670) );
  NANDN U1898 ( .A(n1579), .B(n1578), .Z(n1583) );
  NANDN U1899 ( .A(n1581), .B(n1580), .Z(n1582) );
  AND U1900 ( .A(n1583), .B(n1582), .Z(n1669) );
  XOR U1901 ( .A(n1670), .B(n1669), .Z(n1752) );
  NANDN U1902 ( .A(n1585), .B(n1584), .Z(n1589) );
  NANDN U1903 ( .A(n1587), .B(n1586), .Z(n1588) );
  AND U1904 ( .A(n1589), .B(n1588), .Z(n1664) );
  NANDN U1905 ( .A(n1591), .B(n1590), .Z(n1595) );
  OR U1906 ( .A(n1593), .B(n1592), .Z(n1594) );
  NAND U1907 ( .A(n1595), .B(n1594), .Z(n1663) );
  XNOR U1908 ( .A(n1664), .B(n1663), .Z(n1666) );
  AND U1909 ( .A(b[0]), .B(a[24]), .Z(n1596) );
  XOR U1910 ( .A(b[1]), .B(n1596), .Z(n1598) );
  NANDN U1911 ( .A(b[0]), .B(a[23]), .Z(n1597) );
  AND U1912 ( .A(n1598), .B(n1597), .Z(n1680) );
  XOR U1913 ( .A(b[24]), .B(b[23]), .Z(n34298) );
  IV U1914 ( .A(n34298), .Z(n33994) );
  ANDN U1915 ( .B(a[0]), .A(n33994), .Z(n1707) );
  NANDN U1916 ( .A(n32996), .B(n1599), .Z(n1601) );
  XOR U1917 ( .A(b[21]), .B(a[4]), .Z(n1742) );
  NANDN U1918 ( .A(n33271), .B(n1742), .Z(n1600) );
  AND U1919 ( .A(n1601), .B(n1600), .Z(n1679) );
  XOR U1920 ( .A(n1707), .B(n1679), .Z(n1681) );
  XNOR U1921 ( .A(n1680), .B(n1681), .Z(n1673) );
  NANDN U1922 ( .A(n29499), .B(n1602), .Z(n1604) );
  XOR U1923 ( .A(b[7]), .B(a[18]), .Z(n1730) );
  NANDN U1924 ( .A(n29735), .B(n1730), .Z(n1603) );
  AND U1925 ( .A(n1604), .B(n1603), .Z(n1727) );
  NANDN U1926 ( .A(n28889), .B(n1605), .Z(n1607) );
  XOR U1927 ( .A(b[5]), .B(a[20]), .Z(n1733) );
  NANDN U1928 ( .A(n29138), .B(n1733), .Z(n1606) );
  AND U1929 ( .A(n1607), .B(n1606), .Z(n1725) );
  NANDN U1930 ( .A(n32013), .B(n1608), .Z(n1610) );
  XOR U1931 ( .A(b[17]), .B(a[8]), .Z(n1736) );
  NANDN U1932 ( .A(n32292), .B(n1736), .Z(n1609) );
  NAND U1933 ( .A(n1610), .B(n1609), .Z(n1724) );
  XNOR U1934 ( .A(n1725), .B(n1724), .Z(n1726) );
  XOR U1935 ( .A(n1727), .B(n1726), .Z(n1674) );
  XNOR U1936 ( .A(n1673), .B(n1674), .Z(n1675) );
  NANDN U1937 ( .A(n31536), .B(n1611), .Z(n1613) );
  XOR U1938 ( .A(b[15]), .B(a[10]), .Z(n1703) );
  NANDN U1939 ( .A(n31925), .B(n1703), .Z(n1612) );
  AND U1940 ( .A(n1613), .B(n1612), .Z(n1721) );
  NANDN U1941 ( .A(n30482), .B(n1614), .Z(n1616) );
  XOR U1942 ( .A(b[11]), .B(a[14]), .Z(n1748) );
  NANDN U1943 ( .A(n30891), .B(n1748), .Z(n1615) );
  NAND U1944 ( .A(n1616), .B(n1615), .Z(n1720) );
  XNOR U1945 ( .A(n1721), .B(n1720), .Z(n1723) );
  NAND U1946 ( .A(n33000), .B(n1617), .Z(n1619) );
  XNOR U1947 ( .A(b[19]), .B(a[6]), .Z(n1739) );
  NANDN U1948 ( .A(n1739), .B(n33001), .Z(n1618) );
  NAND U1949 ( .A(n1619), .B(n1618), .Z(n1716) );
  ANDN U1950 ( .B(n1620), .A(n33868), .Z(n33492) );
  NAND U1951 ( .A(n33492), .B(n1621), .Z(n1623) );
  XNOR U1952 ( .A(b[23]), .B(a[2]), .Z(n1684) );
  NANDN U1953 ( .A(n1684), .B(n33868), .Z(n1622) );
  NAND U1954 ( .A(n1623), .B(n1622), .Z(n1715) );
  NANDN U1955 ( .A(n210), .B(n1624), .Z(n1626) );
  XOR U1956 ( .A(b[9]), .B(a[16]), .Z(n1745) );
  NANDN U1957 ( .A(n30267), .B(n1745), .Z(n1625) );
  NAND U1958 ( .A(n1626), .B(n1625), .Z(n1714) );
  XOR U1959 ( .A(n1715), .B(n1714), .Z(n1717) );
  XOR U1960 ( .A(n1716), .B(n1717), .Z(n1722) );
  XNOR U1961 ( .A(n1723), .B(n1722), .Z(n1676) );
  XNOR U1962 ( .A(n1675), .B(n1676), .Z(n1665) );
  XOR U1963 ( .A(n1666), .B(n1665), .Z(n1751) );
  XOR U1964 ( .A(n1752), .B(n1751), .Z(n1754) );
  XOR U1965 ( .A(n1753), .B(n1754), .Z(n1660) );
  NAND U1966 ( .A(n1628), .B(n1627), .Z(n1632) );
  NAND U1967 ( .A(n1630), .B(n1629), .Z(n1631) );
  AND U1968 ( .A(n1632), .B(n1631), .Z(n1657) );
  NANDN U1969 ( .A(n1634), .B(n1633), .Z(n1638) );
  NANDN U1970 ( .A(n1636), .B(n1635), .Z(n1637) );
  NAND U1971 ( .A(n1638), .B(n1637), .Z(n1658) );
  XNOR U1972 ( .A(n1657), .B(n1658), .Z(n1659) );
  XOR U1973 ( .A(n1660), .B(n1659), .Z(n1652) );
  XNOR U1974 ( .A(n1651), .B(n1652), .Z(n1653) );
  XNOR U1975 ( .A(n1654), .B(n1653), .Z(n1645) );
  NANDN U1976 ( .A(n1640), .B(n1639), .Z(n1644) );
  OR U1977 ( .A(n1642), .B(n1641), .Z(n1643) );
  NAND U1978 ( .A(n1644), .B(n1643), .Z(n1646) );
  XNOR U1979 ( .A(n1645), .B(n1646), .Z(n1647) );
  XNOR U1980 ( .A(n1648), .B(n1647), .Z(n1758) );
  XNOR U1981 ( .A(n1759), .B(n1758), .Z(c[88]) );
  NANDN U1982 ( .A(n1646), .B(n1645), .Z(n1650) );
  NANDN U1983 ( .A(n1648), .B(n1647), .Z(n1649) );
  AND U1984 ( .A(n1650), .B(n1649), .Z(n1770) );
  NANDN U1985 ( .A(n1652), .B(n1651), .Z(n1656) );
  NANDN U1986 ( .A(n1654), .B(n1653), .Z(n1655) );
  AND U1987 ( .A(n1656), .B(n1655), .Z(n1768) );
  NANDN U1988 ( .A(n1658), .B(n1657), .Z(n1662) );
  NANDN U1989 ( .A(n1660), .B(n1659), .Z(n1661) );
  AND U1990 ( .A(n1662), .B(n1661), .Z(n1776) );
  NANDN U1991 ( .A(n1668), .B(n1667), .Z(n1672) );
  NAND U1992 ( .A(n1670), .B(n1669), .Z(n1671) );
  AND U1993 ( .A(n1672), .B(n1671), .Z(n1785) );
  XNOR U1994 ( .A(n1786), .B(n1785), .Z(n1788) );
  NANDN U1995 ( .A(n1674), .B(n1673), .Z(n1678) );
  NANDN U1996 ( .A(n1676), .B(n1675), .Z(n1677) );
  AND U1997 ( .A(n1678), .B(n1677), .Z(n1780) );
  NANDN U1998 ( .A(n1679), .B(n1707), .Z(n1683) );
  NANDN U1999 ( .A(n1681), .B(n1680), .Z(n1682) );
  AND U2000 ( .A(n1683), .B(n1682), .Z(n1793) );
  NANDN U2001 ( .A(n1684), .B(n33492), .Z(n1686) );
  XOR U2002 ( .A(b[23]), .B(a[3]), .Z(n1828) );
  NANDN U2003 ( .A(n33644), .B(n1828), .Z(n1685) );
  AND U2004 ( .A(n1686), .B(n1685), .Z(n1846) );
  XOR U2005 ( .A(b[25]), .B(a[1]), .Z(n1807) );
  NANDN U2006 ( .A(n33994), .B(n1807), .Z(n1693) );
  ANDN U2007 ( .B(b[24]), .A(b[25]), .Z(n1687) );
  NAND U2008 ( .A(n1687), .B(a[0]), .Z(n1690) );
  NAND U2009 ( .A(b[23]), .B(b[24]), .Z(n1688) );
  NAND U2010 ( .A(b[25]), .B(n1688), .Z(n1706) );
  OR U2011 ( .A(a[0]), .B(n1706), .Z(n1689) );
  NAND U2012 ( .A(n1690), .B(n1689), .Z(n1691) );
  NAND U2013 ( .A(n33994), .B(n1691), .Z(n1692) );
  AND U2014 ( .A(n1693), .B(n1692), .Z(n1847) );
  XOR U2015 ( .A(n1846), .B(n1847), .Z(n1799) );
  NAND U2016 ( .A(b[0]), .B(a[25]), .Z(n1694) );
  XNOR U2017 ( .A(b[1]), .B(n1694), .Z(n1696) );
  NANDN U2018 ( .A(b[0]), .B(a[24]), .Z(n1695) );
  NAND U2019 ( .A(n1696), .B(n1695), .Z(n1797) );
  NANDN U2020 ( .A(n1697), .B(n31507), .Z(n1699) );
  XNOR U2021 ( .A(b[13]), .B(a[13]), .Z(n1854) );
  NANDN U2022 ( .A(n1854), .B(n31508), .Z(n1698) );
  NAND U2023 ( .A(n1699), .B(n1698), .Z(n1798) );
  XOR U2024 ( .A(n1797), .B(n1798), .Z(n1800) );
  XOR U2025 ( .A(n1799), .B(n1800), .Z(n1792) );
  NANDN U2026 ( .A(n1700), .B(n9942), .Z(n1702) );
  XOR U2027 ( .A(b[3]), .B(a[23]), .Z(n1851) );
  NANDN U2028 ( .A(n28941), .B(n1851), .Z(n1701) );
  AND U2029 ( .A(n1702), .B(n1701), .Z(n1816) );
  NANDN U2030 ( .A(n31536), .B(n1703), .Z(n1705) );
  XOR U2031 ( .A(b[15]), .B(a[11]), .Z(n1848) );
  NANDN U2032 ( .A(n31925), .B(n1848), .Z(n1704) );
  AND U2033 ( .A(n1705), .B(n1704), .Z(n1814) );
  IV U2034 ( .A(n1706), .Z(n34619) );
  ANDN U2035 ( .B(n34619), .A(n1707), .Z(n1813) );
  XNOR U2036 ( .A(n1814), .B(n1813), .Z(n1815) );
  XNOR U2037 ( .A(n1816), .B(n1815), .Z(n1791) );
  XOR U2038 ( .A(n1792), .B(n1791), .Z(n1794) );
  XOR U2039 ( .A(n1793), .B(n1794), .Z(n1871) );
  NANDN U2040 ( .A(n1709), .B(n1708), .Z(n1713) );
  NANDN U2041 ( .A(n1711), .B(n1710), .Z(n1712) );
  AND U2042 ( .A(n1713), .B(n1712), .Z(n1870) );
  NAND U2043 ( .A(n1715), .B(n1714), .Z(n1719) );
  NAND U2044 ( .A(n1717), .B(n1716), .Z(n1718) );
  AND U2045 ( .A(n1719), .B(n1718), .Z(n1869) );
  XOR U2046 ( .A(n1870), .B(n1869), .Z(n1872) );
  XNOR U2047 ( .A(n1871), .B(n1872), .Z(n1779) );
  XNOR U2048 ( .A(n1780), .B(n1779), .Z(n1781) );
  NANDN U2049 ( .A(n1725), .B(n1724), .Z(n1729) );
  NANDN U2050 ( .A(n1727), .B(n1726), .Z(n1728) );
  AND U2051 ( .A(n1729), .B(n1728), .Z(n1876) );
  NANDN U2052 ( .A(n29499), .B(n1730), .Z(n1732) );
  XOR U2053 ( .A(b[7]), .B(a[19]), .Z(n1837) );
  NANDN U2054 ( .A(n29735), .B(n1837), .Z(n1731) );
  AND U2055 ( .A(n1732), .B(n1731), .Z(n1842) );
  NANDN U2056 ( .A(n28889), .B(n1733), .Z(n1735) );
  XOR U2057 ( .A(b[5]), .B(a[21]), .Z(n1860) );
  NANDN U2058 ( .A(n29138), .B(n1860), .Z(n1734) );
  AND U2059 ( .A(n1735), .B(n1734), .Z(n1841) );
  NANDN U2060 ( .A(n32013), .B(n1736), .Z(n1738) );
  XOR U2061 ( .A(b[17]), .B(a[9]), .Z(n1810) );
  NANDN U2062 ( .A(n32292), .B(n1810), .Z(n1737) );
  NAND U2063 ( .A(n1738), .B(n1737), .Z(n1840) );
  XOR U2064 ( .A(n1841), .B(n1840), .Z(n1843) );
  XOR U2065 ( .A(n1842), .B(n1843), .Z(n1865) );
  NANDN U2066 ( .A(n1739), .B(n33000), .Z(n1741) );
  XOR U2067 ( .A(b[19]), .B(a[7]), .Z(n1857) );
  NANDN U2068 ( .A(n32823), .B(n1857), .Z(n1740) );
  AND U2069 ( .A(n1741), .B(n1740), .Z(n1821) );
  NANDN U2070 ( .A(n32996), .B(n1742), .Z(n1744) );
  XOR U2071 ( .A(b[21]), .B(a[5]), .Z(n1803) );
  NANDN U2072 ( .A(n33271), .B(n1803), .Z(n1743) );
  AND U2073 ( .A(n1744), .B(n1743), .Z(n1820) );
  NANDN U2074 ( .A(n210), .B(n1745), .Z(n1747) );
  XOR U2075 ( .A(b[9]), .B(a[17]), .Z(n1831) );
  NANDN U2076 ( .A(n30267), .B(n1831), .Z(n1746) );
  NAND U2077 ( .A(n1747), .B(n1746), .Z(n1819) );
  XOR U2078 ( .A(n1820), .B(n1819), .Z(n1822) );
  XOR U2079 ( .A(n1821), .B(n1822), .Z(n1864) );
  NAND U2080 ( .A(n31059), .B(n1748), .Z(n1750) );
  XNOR U2081 ( .A(b[11]), .B(a[15]), .Z(n1834) );
  NANDN U2082 ( .A(n1834), .B(n31060), .Z(n1749) );
  AND U2083 ( .A(n1750), .B(n1749), .Z(n1863) );
  XOR U2084 ( .A(n1864), .B(n1863), .Z(n1866) );
  XNOR U2085 ( .A(n1865), .B(n1866), .Z(n1875) );
  XNOR U2086 ( .A(n1876), .B(n1875), .Z(n1877) );
  XOR U2087 ( .A(n1878), .B(n1877), .Z(n1782) );
  XNOR U2088 ( .A(n1781), .B(n1782), .Z(n1787) );
  XOR U2089 ( .A(n1788), .B(n1787), .Z(n1774) );
  NANDN U2090 ( .A(n1752), .B(n1751), .Z(n1756) );
  OR U2091 ( .A(n1754), .B(n1753), .Z(n1755) );
  AND U2092 ( .A(n1756), .B(n1755), .Z(n1773) );
  XNOR U2093 ( .A(n1774), .B(n1773), .Z(n1775) );
  XNOR U2094 ( .A(n1776), .B(n1775), .Z(n1767) );
  XNOR U2095 ( .A(n1768), .B(n1767), .Z(n1769) );
  XNOR U2096 ( .A(n1770), .B(n1769), .Z(n1762) );
  XNOR U2097 ( .A(sreg[89]), .B(n1762), .Z(n1764) );
  NANDN U2098 ( .A(sreg[88]), .B(n1757), .Z(n1761) );
  NAND U2099 ( .A(n1759), .B(n1758), .Z(n1760) );
  NAND U2100 ( .A(n1761), .B(n1760), .Z(n1763) );
  XNOR U2101 ( .A(n1764), .B(n1763), .Z(c[89]) );
  NANDN U2102 ( .A(sreg[89]), .B(n1762), .Z(n1766) );
  NAND U2103 ( .A(n1764), .B(n1763), .Z(n1765) );
  NAND U2104 ( .A(n1766), .B(n1765), .Z(n2003) );
  XNOR U2105 ( .A(sreg[90]), .B(n2003), .Z(n2005) );
  NANDN U2106 ( .A(n1768), .B(n1767), .Z(n1772) );
  NANDN U2107 ( .A(n1770), .B(n1769), .Z(n1771) );
  AND U2108 ( .A(n1772), .B(n1771), .Z(n1884) );
  NANDN U2109 ( .A(n1774), .B(n1773), .Z(n1778) );
  NANDN U2110 ( .A(n1776), .B(n1775), .Z(n1777) );
  AND U2111 ( .A(n1778), .B(n1777), .Z(n1882) );
  NANDN U2112 ( .A(n1780), .B(n1779), .Z(n1784) );
  NANDN U2113 ( .A(n1782), .B(n1781), .Z(n1783) );
  AND U2114 ( .A(n1784), .B(n1783), .Z(n1887) );
  NANDN U2115 ( .A(n1786), .B(n1785), .Z(n1790) );
  NAND U2116 ( .A(n1788), .B(n1787), .Z(n1789) );
  NAND U2117 ( .A(n1790), .B(n1789), .Z(n1888) );
  XNOR U2118 ( .A(n1887), .B(n1888), .Z(n1889) );
  NANDN U2119 ( .A(n1792), .B(n1791), .Z(n1796) );
  OR U2120 ( .A(n1794), .B(n1793), .Z(n1795) );
  AND U2121 ( .A(n1796), .B(n1795), .Z(n1906) );
  NANDN U2122 ( .A(n1798), .B(n1797), .Z(n1802) );
  OR U2123 ( .A(n1800), .B(n1799), .Z(n1801) );
  AND U2124 ( .A(n1802), .B(n1801), .Z(n1986) );
  NANDN U2125 ( .A(n32996), .B(n1803), .Z(n1805) );
  XOR U2126 ( .A(b[21]), .B(a[6]), .Z(n1970) );
  NANDN U2127 ( .A(n33271), .B(n1970), .Z(n1804) );
  AND U2128 ( .A(n1805), .B(n1804), .Z(n1941) );
  XOR U2129 ( .A(b[24]), .B(b[25]), .Z(n1806) );
  ANDN U2130 ( .B(n1806), .A(n34298), .Z(n34297) );
  IV U2131 ( .A(n34297), .Z(n33875) );
  NANDN U2132 ( .A(n33875), .B(n1807), .Z(n1809) );
  XOR U2133 ( .A(b[25]), .B(a[2]), .Z(n1921) );
  NANDN U2134 ( .A(n33994), .B(n1921), .Z(n1808) );
  AND U2135 ( .A(n1809), .B(n1808), .Z(n1940) );
  NANDN U2136 ( .A(n32013), .B(n1810), .Z(n1812) );
  XOR U2137 ( .A(b[17]), .B(a[10]), .Z(n1967) );
  NANDN U2138 ( .A(n32292), .B(n1967), .Z(n1811) );
  NAND U2139 ( .A(n1812), .B(n1811), .Z(n1939) );
  XOR U2140 ( .A(n1940), .B(n1939), .Z(n1942) );
  XNOR U2141 ( .A(n1941), .B(n1942), .Z(n1985) );
  XNOR U2142 ( .A(n1986), .B(n1985), .Z(n1988) );
  NANDN U2143 ( .A(n1814), .B(n1813), .Z(n1818) );
  NANDN U2144 ( .A(n1816), .B(n1815), .Z(n1817) );
  AND U2145 ( .A(n1818), .B(n1817), .Z(n1987) );
  XNOR U2146 ( .A(n1988), .B(n1987), .Z(n1905) );
  XNOR U2147 ( .A(n1906), .B(n1905), .Z(n1908) );
  NANDN U2148 ( .A(n1820), .B(n1819), .Z(n1824) );
  OR U2149 ( .A(n1822), .B(n1821), .Z(n1823) );
  AND U2150 ( .A(n1824), .B(n1823), .Z(n1994) );
  NAND U2151 ( .A(b[0]), .B(a[26]), .Z(n1825) );
  XNOR U2152 ( .A(b[1]), .B(n1825), .Z(n1827) );
  NANDN U2153 ( .A(b[0]), .B(a[25]), .Z(n1826) );
  NAND U2154 ( .A(n1827), .B(n1826), .Z(n1953) );
  XOR U2155 ( .A(b[26]), .B(b[25]), .Z(n34648) );
  IV U2156 ( .A(n34648), .Z(n34458) );
  ANDN U2157 ( .B(a[0]), .A(n34458), .Z(n1963) );
  IV U2158 ( .A(n33492), .Z(n33866) );
  NANDN U2159 ( .A(n33866), .B(n1828), .Z(n1830) );
  XOR U2160 ( .A(b[23]), .B(a[4]), .Z(n1973) );
  NANDN U2161 ( .A(n33644), .B(n1973), .Z(n1829) );
  AND U2162 ( .A(n1830), .B(n1829), .Z(n1951) );
  XNOR U2163 ( .A(n1963), .B(n1951), .Z(n1952) );
  XNOR U2164 ( .A(n1953), .B(n1952), .Z(n1991) );
  NANDN U2165 ( .A(n210), .B(n1831), .Z(n1833) );
  XOR U2166 ( .A(b[9]), .B(a[18]), .Z(n1976) );
  NANDN U2167 ( .A(n30267), .B(n1976), .Z(n1832) );
  AND U2168 ( .A(n1833), .B(n1832), .Z(n1948) );
  NANDN U2169 ( .A(n1834), .B(n31059), .Z(n1836) );
  XOR U2170 ( .A(b[11]), .B(a[16]), .Z(n1964) );
  NANDN U2171 ( .A(n30891), .B(n1964), .Z(n1835) );
  AND U2172 ( .A(n1836), .B(n1835), .Z(n1946) );
  NANDN U2173 ( .A(n29499), .B(n1837), .Z(n1839) );
  XOR U2174 ( .A(b[7]), .B(a[20]), .Z(n1924) );
  NANDN U2175 ( .A(n29735), .B(n1924), .Z(n1838) );
  NAND U2176 ( .A(n1839), .B(n1838), .Z(n1945) );
  XNOR U2177 ( .A(n1946), .B(n1945), .Z(n1947) );
  XOR U2178 ( .A(n1948), .B(n1947), .Z(n1992) );
  XNOR U2179 ( .A(n1991), .B(n1992), .Z(n1993) );
  XNOR U2180 ( .A(n1994), .B(n1993), .Z(n1900) );
  NANDN U2181 ( .A(n1841), .B(n1840), .Z(n1845) );
  OR U2182 ( .A(n1843), .B(n1842), .Z(n1844) );
  AND U2183 ( .A(n1845), .B(n1844), .Z(n1999) );
  NOR U2184 ( .A(n1847), .B(n1846), .Z(n1935) );
  NAND U2185 ( .A(n32023), .B(n1848), .Z(n1850) );
  XNOR U2186 ( .A(b[15]), .B(a[12]), .Z(n1959) );
  NANDN U2187 ( .A(n1959), .B(n32024), .Z(n1849) );
  AND U2188 ( .A(n1850), .B(n1849), .Z(n1933) );
  NAND U2189 ( .A(n9942), .B(n1851), .Z(n1853) );
  XNOR U2190 ( .A(b[3]), .B(a[24]), .Z(n1956) );
  NANDN U2191 ( .A(n1956), .B(n9653), .Z(n1852) );
  NAND U2192 ( .A(n1853), .B(n1852), .Z(n1934) );
  XOR U2193 ( .A(n1933), .B(n1934), .Z(n1936) );
  XOR U2194 ( .A(n1935), .B(n1936), .Z(n1998) );
  NANDN U2195 ( .A(n1854), .B(n31507), .Z(n1856) );
  XOR U2196 ( .A(b[13]), .B(a[14]), .Z(n1914) );
  NANDN U2197 ( .A(n31293), .B(n1914), .Z(n1855) );
  AND U2198 ( .A(n1856), .B(n1855), .Z(n1982) );
  NANDN U2199 ( .A(n32483), .B(n1857), .Z(n1859) );
  XOR U2200 ( .A(b[19]), .B(a[8]), .Z(n1930) );
  NANDN U2201 ( .A(n32823), .B(n1930), .Z(n1858) );
  AND U2202 ( .A(n1859), .B(n1858), .Z(n1980) );
  NANDN U2203 ( .A(n28889), .B(n1860), .Z(n1862) );
  XOR U2204 ( .A(b[5]), .B(a[22]), .Z(n1927) );
  NANDN U2205 ( .A(n29138), .B(n1927), .Z(n1861) );
  NAND U2206 ( .A(n1862), .B(n1861), .Z(n1979) );
  XNOR U2207 ( .A(n1980), .B(n1979), .Z(n1981) );
  XNOR U2208 ( .A(n1982), .B(n1981), .Z(n1997) );
  XOR U2209 ( .A(n1998), .B(n1997), .Z(n2000) );
  XOR U2210 ( .A(n1999), .B(n2000), .Z(n1899) );
  XOR U2211 ( .A(n1900), .B(n1899), .Z(n1902) );
  NANDN U2212 ( .A(n1864), .B(n1863), .Z(n1868) );
  OR U2213 ( .A(n1866), .B(n1865), .Z(n1867) );
  AND U2214 ( .A(n1868), .B(n1867), .Z(n1901) );
  XOR U2215 ( .A(n1902), .B(n1901), .Z(n1907) );
  XOR U2216 ( .A(n1908), .B(n1907), .Z(n1896) );
  NANDN U2217 ( .A(n1870), .B(n1869), .Z(n1874) );
  OR U2218 ( .A(n1872), .B(n1871), .Z(n1873) );
  AND U2219 ( .A(n1874), .B(n1873), .Z(n1894) );
  NANDN U2220 ( .A(n1876), .B(n1875), .Z(n1880) );
  NANDN U2221 ( .A(n1878), .B(n1877), .Z(n1879) );
  AND U2222 ( .A(n1880), .B(n1879), .Z(n1893) );
  XNOR U2223 ( .A(n1894), .B(n1893), .Z(n1895) );
  XOR U2224 ( .A(n1896), .B(n1895), .Z(n1890) );
  XNOR U2225 ( .A(n1889), .B(n1890), .Z(n1881) );
  XNOR U2226 ( .A(n1882), .B(n1881), .Z(n1883) );
  XNOR U2227 ( .A(n1884), .B(n1883), .Z(n2004) );
  XNOR U2228 ( .A(n2005), .B(n2004), .Z(c[90]) );
  NANDN U2229 ( .A(n1882), .B(n1881), .Z(n1886) );
  NANDN U2230 ( .A(n1884), .B(n1883), .Z(n1885) );
  AND U2231 ( .A(n1886), .B(n1885), .Z(n2016) );
  NANDN U2232 ( .A(n1888), .B(n1887), .Z(n1892) );
  NANDN U2233 ( .A(n1890), .B(n1889), .Z(n1891) );
  AND U2234 ( .A(n1892), .B(n1891), .Z(n2014) );
  NANDN U2235 ( .A(n1894), .B(n1893), .Z(n1898) );
  NANDN U2236 ( .A(n1896), .B(n1895), .Z(n1897) );
  AND U2237 ( .A(n1898), .B(n1897), .Z(n2022) );
  NAND U2238 ( .A(n1900), .B(n1899), .Z(n1904) );
  NAND U2239 ( .A(n1902), .B(n1901), .Z(n1903) );
  AND U2240 ( .A(n1904), .B(n1903), .Z(n2019) );
  NANDN U2241 ( .A(n1906), .B(n1905), .Z(n1910) );
  NAND U2242 ( .A(n1908), .B(n1907), .Z(n1909) );
  AND U2243 ( .A(n1910), .B(n1909), .Z(n2130) );
  NAND U2244 ( .A(b[0]), .B(a[27]), .Z(n1911) );
  XNOR U2245 ( .A(b[1]), .B(n1911), .Z(n1913) );
  NANDN U2246 ( .A(b[0]), .B(a[26]), .Z(n1912) );
  NAND U2247 ( .A(n1913), .B(n1912), .Z(n2080) );
  NANDN U2248 ( .A(n31055), .B(n1914), .Z(n1916) );
  XOR U2249 ( .A(b[13]), .B(a[15]), .Z(n2076) );
  NANDN U2250 ( .A(n31293), .B(n2076), .Z(n1915) );
  NAND U2251 ( .A(n1916), .B(n1915), .Z(n2079) );
  XNOR U2252 ( .A(n2080), .B(n2079), .Z(n2081) );
  XOR U2253 ( .A(b[27]), .B(b[26]), .Z(n2118) );
  XOR U2254 ( .A(b[27]), .B(a[0]), .Z(n1917) );
  NAND U2255 ( .A(n2118), .B(n1917), .Z(n1918) );
  OR U2256 ( .A(n1918), .B(n34648), .Z(n1920) );
  XOR U2257 ( .A(b[27]), .B(a[1]), .Z(n2119) );
  NAND U2258 ( .A(n34648), .B(n2119), .Z(n1919) );
  AND U2259 ( .A(n1920), .B(n1919), .Z(n2113) );
  NANDN U2260 ( .A(n33875), .B(n1921), .Z(n1923) );
  XOR U2261 ( .A(b[25]), .B(a[3]), .Z(n2110) );
  NANDN U2262 ( .A(n33994), .B(n2110), .Z(n1922) );
  NAND U2263 ( .A(n1923), .B(n1922), .Z(n2114) );
  XOR U2264 ( .A(n2113), .B(n2114), .Z(n2082) );
  XNOR U2265 ( .A(n2081), .B(n2082), .Z(n2043) );
  NANDN U2266 ( .A(n29499), .B(n1924), .Z(n1926) );
  XOR U2267 ( .A(b[7]), .B(a[21]), .Z(n2064) );
  NANDN U2268 ( .A(n29735), .B(n2064), .Z(n1925) );
  AND U2269 ( .A(n1926), .B(n1925), .Z(n2125) );
  NANDN U2270 ( .A(n28889), .B(n1927), .Z(n1929) );
  XOR U2271 ( .A(b[5]), .B(a[23]), .Z(n2055) );
  NANDN U2272 ( .A(n29138), .B(n2055), .Z(n1928) );
  AND U2273 ( .A(n1929), .B(n1928), .Z(n2123) );
  NANDN U2274 ( .A(n32483), .B(n1930), .Z(n1932) );
  XOR U2275 ( .A(b[19]), .B(a[9]), .Z(n2049) );
  NANDN U2276 ( .A(n32823), .B(n2049), .Z(n1931) );
  NAND U2277 ( .A(n1932), .B(n1931), .Z(n2122) );
  XNOR U2278 ( .A(n2123), .B(n2122), .Z(n2124) );
  XOR U2279 ( .A(n2125), .B(n2124), .Z(n2044) );
  XNOR U2280 ( .A(n2043), .B(n2044), .Z(n2045) );
  NANDN U2281 ( .A(n1934), .B(n1933), .Z(n1938) );
  OR U2282 ( .A(n1936), .B(n1935), .Z(n1937) );
  NAND U2283 ( .A(n1938), .B(n1937), .Z(n2046) );
  XNOR U2284 ( .A(n2045), .B(n2046), .Z(n2034) );
  NANDN U2285 ( .A(n1940), .B(n1939), .Z(n1944) );
  OR U2286 ( .A(n1942), .B(n1941), .Z(n1943) );
  NAND U2287 ( .A(n1944), .B(n1943), .Z(n2032) );
  NANDN U2288 ( .A(n1946), .B(n1945), .Z(n1950) );
  NANDN U2289 ( .A(n1948), .B(n1947), .Z(n1949) );
  NAND U2290 ( .A(n1950), .B(n1949), .Z(n2031) );
  XOR U2291 ( .A(n2032), .B(n2031), .Z(n2033) );
  XOR U2292 ( .A(n2034), .B(n2033), .Z(n2040) );
  NANDN U2293 ( .A(n1951), .B(n1963), .Z(n1955) );
  NANDN U2294 ( .A(n1953), .B(n1952), .Z(n1954) );
  AND U2295 ( .A(n1955), .B(n1954), .Z(n2092) );
  NANDN U2296 ( .A(n1956), .B(n9942), .Z(n1958) );
  XOR U2297 ( .A(b[3]), .B(a[25]), .Z(n2070) );
  NANDN U2298 ( .A(n28941), .B(n2070), .Z(n1957) );
  AND U2299 ( .A(n1958), .B(n1957), .Z(n2104) );
  NANDN U2300 ( .A(n1959), .B(n32023), .Z(n1961) );
  XOR U2301 ( .A(b[15]), .B(a[13]), .Z(n2115) );
  NANDN U2302 ( .A(n31925), .B(n2115), .Z(n1960) );
  NAND U2303 ( .A(n1961), .B(n1960), .Z(n2103) );
  XNOR U2304 ( .A(n2104), .B(n2103), .Z(n2106) );
  NAND U2305 ( .A(b[25]), .B(b[26]), .Z(n1962) );
  AND U2306 ( .A(b[27]), .B(n1962), .Z(n34992) );
  ANDN U2307 ( .B(n34992), .A(n1963), .Z(n2105) );
  XOR U2308 ( .A(n2106), .B(n2105), .Z(n2091) );
  XNOR U2309 ( .A(n2092), .B(n2091), .Z(n2094) );
  NANDN U2310 ( .A(n30482), .B(n1964), .Z(n1966) );
  XOR U2311 ( .A(b[11]), .B(a[17]), .Z(n2058) );
  NANDN U2312 ( .A(n30891), .B(n2058), .Z(n1965) );
  AND U2313 ( .A(n1966), .B(n1965), .Z(n2098) );
  NANDN U2314 ( .A(n32013), .B(n1967), .Z(n1969) );
  XOR U2315 ( .A(b[17]), .B(a[11]), .Z(n2061) );
  NANDN U2316 ( .A(n32292), .B(n2061), .Z(n1968) );
  NAND U2317 ( .A(n1969), .B(n1968), .Z(n2097) );
  XNOR U2318 ( .A(n2098), .B(n2097), .Z(n2099) );
  NANDN U2319 ( .A(n32996), .B(n1970), .Z(n1972) );
  XOR U2320 ( .A(b[21]), .B(a[7]), .Z(n2052) );
  NANDN U2321 ( .A(n33271), .B(n2052), .Z(n1971) );
  AND U2322 ( .A(n1972), .B(n1971), .Z(n2088) );
  NANDN U2323 ( .A(n33866), .B(n1973), .Z(n1975) );
  XOR U2324 ( .A(b[23]), .B(a[5]), .Z(n2073) );
  NANDN U2325 ( .A(n33644), .B(n2073), .Z(n1974) );
  AND U2326 ( .A(n1975), .B(n1974), .Z(n2086) );
  NANDN U2327 ( .A(n210), .B(n1976), .Z(n1978) );
  XOR U2328 ( .A(b[9]), .B(a[19]), .Z(n2067) );
  NANDN U2329 ( .A(n30267), .B(n2067), .Z(n1977) );
  NAND U2330 ( .A(n1978), .B(n1977), .Z(n2085) );
  XNOR U2331 ( .A(n2086), .B(n2085), .Z(n2087) );
  XOR U2332 ( .A(n2088), .B(n2087), .Z(n2100) );
  XNOR U2333 ( .A(n2099), .B(n2100), .Z(n2093) );
  XOR U2334 ( .A(n2094), .B(n2093), .Z(n2038) );
  NANDN U2335 ( .A(n1980), .B(n1979), .Z(n1984) );
  NANDN U2336 ( .A(n1982), .B(n1981), .Z(n1983) );
  AND U2337 ( .A(n1984), .B(n1983), .Z(n2037) );
  XNOR U2338 ( .A(n2038), .B(n2037), .Z(n2039) );
  XNOR U2339 ( .A(n2040), .B(n2039), .Z(n2128) );
  NANDN U2340 ( .A(n1986), .B(n1985), .Z(n1990) );
  NAND U2341 ( .A(n1988), .B(n1987), .Z(n1989) );
  AND U2342 ( .A(n1990), .B(n1989), .Z(n2028) );
  NANDN U2343 ( .A(n1992), .B(n1991), .Z(n1996) );
  NANDN U2344 ( .A(n1994), .B(n1993), .Z(n1995) );
  AND U2345 ( .A(n1996), .B(n1995), .Z(n2025) );
  NANDN U2346 ( .A(n1998), .B(n1997), .Z(n2002) );
  OR U2347 ( .A(n2000), .B(n1999), .Z(n2001) );
  NAND U2348 ( .A(n2002), .B(n2001), .Z(n2026) );
  XNOR U2349 ( .A(n2025), .B(n2026), .Z(n2027) );
  XOR U2350 ( .A(n2028), .B(n2027), .Z(n2129) );
  XOR U2351 ( .A(n2128), .B(n2129), .Z(n2131) );
  XOR U2352 ( .A(n2130), .B(n2131), .Z(n2020) );
  XNOR U2353 ( .A(n2019), .B(n2020), .Z(n2021) );
  XNOR U2354 ( .A(n2022), .B(n2021), .Z(n2013) );
  XNOR U2355 ( .A(n2014), .B(n2013), .Z(n2015) );
  XNOR U2356 ( .A(n2016), .B(n2015), .Z(n2008) );
  XNOR U2357 ( .A(sreg[91]), .B(n2008), .Z(n2010) );
  NANDN U2358 ( .A(sreg[90]), .B(n2003), .Z(n2007) );
  NAND U2359 ( .A(n2005), .B(n2004), .Z(n2006) );
  NAND U2360 ( .A(n2007), .B(n2006), .Z(n2009) );
  XNOR U2361 ( .A(n2010), .B(n2009), .Z(c[91]) );
  NANDN U2362 ( .A(sreg[91]), .B(n2008), .Z(n2012) );
  NAND U2363 ( .A(n2010), .B(n2009), .Z(n2011) );
  NAND U2364 ( .A(n2012), .B(n2011), .Z(n2267) );
  XNOR U2365 ( .A(sreg[92]), .B(n2267), .Z(n2269) );
  NANDN U2366 ( .A(n2014), .B(n2013), .Z(n2018) );
  NANDN U2367 ( .A(n2016), .B(n2015), .Z(n2017) );
  AND U2368 ( .A(n2018), .B(n2017), .Z(n2137) );
  NANDN U2369 ( .A(n2020), .B(n2019), .Z(n2024) );
  NANDN U2370 ( .A(n2022), .B(n2021), .Z(n2023) );
  AND U2371 ( .A(n2024), .B(n2023), .Z(n2135) );
  NANDN U2372 ( .A(n2026), .B(n2025), .Z(n2030) );
  NANDN U2373 ( .A(n2028), .B(n2027), .Z(n2029) );
  AND U2374 ( .A(n2030), .B(n2029), .Z(n2143) );
  NAND U2375 ( .A(n2032), .B(n2031), .Z(n2036) );
  NAND U2376 ( .A(n2034), .B(n2033), .Z(n2035) );
  AND U2377 ( .A(n2036), .B(n2035), .Z(n2141) );
  NANDN U2378 ( .A(n2038), .B(n2037), .Z(n2042) );
  NANDN U2379 ( .A(n2040), .B(n2039), .Z(n2041) );
  AND U2380 ( .A(n2042), .B(n2041), .Z(n2140) );
  XNOR U2381 ( .A(n2141), .B(n2140), .Z(n2142) );
  XOR U2382 ( .A(n2143), .B(n2142), .Z(n2264) );
  NANDN U2383 ( .A(n2044), .B(n2043), .Z(n2048) );
  NANDN U2384 ( .A(n2046), .B(n2045), .Z(n2047) );
  AND U2385 ( .A(n2048), .B(n2047), .Z(n2234) );
  NANDN U2386 ( .A(n32483), .B(n2049), .Z(n2051) );
  XOR U2387 ( .A(b[19]), .B(a[10]), .Z(n2165) );
  NANDN U2388 ( .A(n32823), .B(n2165), .Z(n2050) );
  AND U2389 ( .A(n2051), .B(n2050), .Z(n2185) );
  NANDN U2390 ( .A(n32996), .B(n2052), .Z(n2054) );
  XOR U2391 ( .A(b[21]), .B(a[8]), .Z(n2192) );
  NANDN U2392 ( .A(n33271), .B(n2192), .Z(n2053) );
  AND U2393 ( .A(n2054), .B(n2053), .Z(n2184) );
  NANDN U2394 ( .A(n28889), .B(n2055), .Z(n2057) );
  XOR U2395 ( .A(b[5]), .B(a[24]), .Z(n2195) );
  NANDN U2396 ( .A(n29138), .B(n2195), .Z(n2056) );
  NAND U2397 ( .A(n2057), .B(n2056), .Z(n2183) );
  XOR U2398 ( .A(n2184), .B(n2183), .Z(n2186) );
  XOR U2399 ( .A(n2185), .B(n2186), .Z(n2252) );
  NANDN U2400 ( .A(n30482), .B(n2058), .Z(n2060) );
  XOR U2401 ( .A(b[11]), .B(a[18]), .Z(n2168) );
  NANDN U2402 ( .A(n30891), .B(n2168), .Z(n2059) );
  AND U2403 ( .A(n2060), .B(n2059), .Z(n2221) );
  NANDN U2404 ( .A(n32013), .B(n2061), .Z(n2063) );
  XOR U2405 ( .A(b[17]), .B(a[12]), .Z(n2201) );
  NANDN U2406 ( .A(n32292), .B(n2201), .Z(n2062) );
  AND U2407 ( .A(n2063), .B(n2062), .Z(n2220) );
  NANDN U2408 ( .A(n29499), .B(n2064), .Z(n2066) );
  XOR U2409 ( .A(b[7]), .B(a[22]), .Z(n2189) );
  NANDN U2410 ( .A(n29735), .B(n2189), .Z(n2065) );
  NAND U2411 ( .A(n2066), .B(n2065), .Z(n2219) );
  XOR U2412 ( .A(n2220), .B(n2219), .Z(n2222) );
  XOR U2413 ( .A(n2221), .B(n2222), .Z(n2250) );
  NAND U2414 ( .A(n30627), .B(n2067), .Z(n2069) );
  XNOR U2415 ( .A(b[9]), .B(a[20]), .Z(n2210) );
  NANDN U2416 ( .A(n2210), .B(n30628), .Z(n2068) );
  AND U2417 ( .A(n2069), .B(n2068), .Z(n2249) );
  XNOR U2418 ( .A(n2250), .B(n2249), .Z(n2251) );
  XNOR U2419 ( .A(n2252), .B(n2251), .Z(n2231) );
  NANDN U2420 ( .A(n209), .B(n2070), .Z(n2072) );
  XOR U2421 ( .A(b[3]), .B(a[26]), .Z(n2198) );
  NANDN U2422 ( .A(n28941), .B(n2198), .Z(n2071) );
  AND U2423 ( .A(n2072), .B(n2071), .Z(n2179) );
  NANDN U2424 ( .A(n33866), .B(n2073), .Z(n2075) );
  XOR U2425 ( .A(b[23]), .B(a[6]), .Z(n2204) );
  NANDN U2426 ( .A(n33644), .B(n2204), .Z(n2074) );
  AND U2427 ( .A(n2075), .B(n2074), .Z(n2178) );
  NANDN U2428 ( .A(n31055), .B(n2076), .Z(n2078) );
  XOR U2429 ( .A(b[13]), .B(a[16]), .Z(n2162) );
  NANDN U2430 ( .A(n31293), .B(n2162), .Z(n2077) );
  NAND U2431 ( .A(n2078), .B(n2077), .Z(n2177) );
  XOR U2432 ( .A(n2178), .B(n2177), .Z(n2180) );
  XOR U2433 ( .A(n2179), .B(n2180), .Z(n2238) );
  NANDN U2434 ( .A(n2080), .B(n2079), .Z(n2084) );
  NANDN U2435 ( .A(n2082), .B(n2081), .Z(n2083) );
  AND U2436 ( .A(n2084), .B(n2083), .Z(n2237) );
  XNOR U2437 ( .A(n2238), .B(n2237), .Z(n2239) );
  NANDN U2438 ( .A(n2086), .B(n2085), .Z(n2090) );
  NANDN U2439 ( .A(n2088), .B(n2087), .Z(n2089) );
  NAND U2440 ( .A(n2090), .B(n2089), .Z(n2240) );
  XOR U2441 ( .A(n2239), .B(n2240), .Z(n2232) );
  XNOR U2442 ( .A(n2231), .B(n2232), .Z(n2233) );
  XOR U2443 ( .A(n2234), .B(n2233), .Z(n2257) );
  NANDN U2444 ( .A(n2092), .B(n2091), .Z(n2096) );
  NAND U2445 ( .A(n2094), .B(n2093), .Z(n2095) );
  AND U2446 ( .A(n2096), .B(n2095), .Z(n2256) );
  NANDN U2447 ( .A(n2098), .B(n2097), .Z(n2102) );
  NANDN U2448 ( .A(n2100), .B(n2099), .Z(n2101) );
  AND U2449 ( .A(n2102), .B(n2101), .Z(n2228) );
  NAND U2450 ( .A(b[0]), .B(a[28]), .Z(n2107) );
  XNOR U2451 ( .A(b[1]), .B(n2107), .Z(n2109) );
  NANDN U2452 ( .A(b[0]), .B(a[27]), .Z(n2108) );
  NAND U2453 ( .A(n2109), .B(n2108), .Z(n2216) );
  XOR U2454 ( .A(b[28]), .B(b[27]), .Z(n35002) );
  IV U2455 ( .A(n35002), .Z(n34722) );
  ANDN U2456 ( .B(a[0]), .A(n34722), .Z(n2213) );
  NANDN U2457 ( .A(n33875), .B(n2110), .Z(n2112) );
  XOR U2458 ( .A(b[25]), .B(a[4]), .Z(n2207) );
  NANDN U2459 ( .A(n33994), .B(n2207), .Z(n2111) );
  AND U2460 ( .A(n2112), .B(n2111), .Z(n2214) );
  XOR U2461 ( .A(n2213), .B(n2214), .Z(n2215) );
  XOR U2462 ( .A(n2216), .B(n2215), .Z(n2244) );
  ANDN U2463 ( .B(n2114), .A(n2113), .Z(n2174) );
  NAND U2464 ( .A(n32023), .B(n2115), .Z(n2117) );
  XNOR U2465 ( .A(b[15]), .B(a[14]), .Z(n2159) );
  NANDN U2466 ( .A(n2159), .B(n32024), .Z(n2116) );
  AND U2467 ( .A(n2117), .B(n2116), .Z(n2171) );
  ANDN U2468 ( .B(n2118), .A(n34648), .Z(n34647) );
  NAND U2469 ( .A(n34647), .B(n2119), .Z(n2121) );
  XNOR U2470 ( .A(b[27]), .B(a[2]), .Z(n2146) );
  NANDN U2471 ( .A(n2146), .B(n34648), .Z(n2120) );
  NAND U2472 ( .A(n2121), .B(n2120), .Z(n2172) );
  XNOR U2473 ( .A(n2171), .B(n2172), .Z(n2173) );
  XNOR U2474 ( .A(n2174), .B(n2173), .Z(n2243) );
  XNOR U2475 ( .A(n2244), .B(n2243), .Z(n2246) );
  NANDN U2476 ( .A(n2123), .B(n2122), .Z(n2127) );
  NANDN U2477 ( .A(n2125), .B(n2124), .Z(n2126) );
  AND U2478 ( .A(n2127), .B(n2126), .Z(n2245) );
  XNOR U2479 ( .A(n2246), .B(n2245), .Z(n2225) );
  XNOR U2480 ( .A(n2226), .B(n2225), .Z(n2227) );
  XNOR U2481 ( .A(n2228), .B(n2227), .Z(n2255) );
  XOR U2482 ( .A(n2256), .B(n2255), .Z(n2258) );
  XOR U2483 ( .A(n2257), .B(n2258), .Z(n2262) );
  NANDN U2484 ( .A(n2129), .B(n2128), .Z(n2133) );
  NANDN U2485 ( .A(n2131), .B(n2130), .Z(n2132) );
  NAND U2486 ( .A(n2133), .B(n2132), .Z(n2261) );
  XNOR U2487 ( .A(n2262), .B(n2261), .Z(n2263) );
  XNOR U2488 ( .A(n2264), .B(n2263), .Z(n2134) );
  XNOR U2489 ( .A(n2135), .B(n2134), .Z(n2136) );
  XNOR U2490 ( .A(n2137), .B(n2136), .Z(n2268) );
  XNOR U2491 ( .A(n2269), .B(n2268), .Z(c[92]) );
  NANDN U2492 ( .A(n2135), .B(n2134), .Z(n2139) );
  NANDN U2493 ( .A(n2137), .B(n2136), .Z(n2138) );
  AND U2494 ( .A(n2139), .B(n2138), .Z(n2280) );
  NANDN U2495 ( .A(n2141), .B(n2140), .Z(n2145) );
  NAND U2496 ( .A(n2143), .B(n2142), .Z(n2144) );
  AND U2497 ( .A(n2145), .B(n2144), .Z(n2405) );
  NANDN U2498 ( .A(n2146), .B(n34647), .Z(n2148) );
  XOR U2499 ( .A(b[27]), .B(a[3]), .Z(n2322) );
  NANDN U2500 ( .A(n34458), .B(n2322), .Z(n2147) );
  AND U2501 ( .A(n2148), .B(n2147), .Z(n2353) );
  XOR U2502 ( .A(b[29]), .B(a[1]), .Z(n2347) );
  NANDN U2503 ( .A(n34722), .B(n2347), .Z(n2155) );
  ANDN U2504 ( .B(b[28]), .A(b[29]), .Z(n2149) );
  NAND U2505 ( .A(n2149), .B(a[0]), .Z(n2152) );
  NAND U2506 ( .A(b[27]), .B(b[28]), .Z(n2150) );
  NAND U2507 ( .A(b[29]), .B(n2150), .Z(n35340) );
  OR U2508 ( .A(a[0]), .B(n35340), .Z(n2151) );
  NAND U2509 ( .A(n2152), .B(n2151), .Z(n2153) );
  NAND U2510 ( .A(n34722), .B(n2153), .Z(n2154) );
  AND U2511 ( .A(n2155), .B(n2154), .Z(n2354) );
  XOR U2512 ( .A(n2353), .B(n2354), .Z(n2387) );
  NAND U2513 ( .A(b[0]), .B(a[29]), .Z(n2156) );
  XNOR U2514 ( .A(b[1]), .B(n2156), .Z(n2158) );
  NANDN U2515 ( .A(b[0]), .B(a[28]), .Z(n2157) );
  NAND U2516 ( .A(n2158), .B(n2157), .Z(n2385) );
  NANDN U2517 ( .A(n2159), .B(n32023), .Z(n2161) );
  XNOR U2518 ( .A(b[15]), .B(a[15]), .Z(n2361) );
  NANDN U2519 ( .A(n2361), .B(n32024), .Z(n2160) );
  NAND U2520 ( .A(n2161), .B(n2160), .Z(n2386) );
  XOR U2521 ( .A(n2385), .B(n2386), .Z(n2388) );
  XOR U2522 ( .A(n2387), .B(n2388), .Z(n2392) );
  NANDN U2523 ( .A(n31055), .B(n2162), .Z(n2164) );
  XOR U2524 ( .A(b[13]), .B(a[17]), .Z(n2370) );
  NANDN U2525 ( .A(n31293), .B(n2370), .Z(n2163) );
  AND U2526 ( .A(n2164), .B(n2163), .Z(n2382) );
  NANDN U2527 ( .A(n32483), .B(n2165), .Z(n2167) );
  XOR U2528 ( .A(b[19]), .B(a[11]), .Z(n2373) );
  NANDN U2529 ( .A(n32823), .B(n2373), .Z(n2166) );
  AND U2530 ( .A(n2167), .B(n2166), .Z(n2380) );
  NANDN U2531 ( .A(n30482), .B(n2168), .Z(n2170) );
  XOR U2532 ( .A(b[11]), .B(a[19]), .Z(n2367) );
  NANDN U2533 ( .A(n30891), .B(n2367), .Z(n2169) );
  NAND U2534 ( .A(n2170), .B(n2169), .Z(n2379) );
  XNOR U2535 ( .A(n2380), .B(n2379), .Z(n2381) );
  XNOR U2536 ( .A(n2382), .B(n2381), .Z(n2391) );
  XNOR U2537 ( .A(n2392), .B(n2391), .Z(n2393) );
  NANDN U2538 ( .A(n2172), .B(n2171), .Z(n2176) );
  NANDN U2539 ( .A(n2174), .B(n2173), .Z(n2175) );
  NAND U2540 ( .A(n2176), .B(n2175), .Z(n2394) );
  XNOR U2541 ( .A(n2393), .B(n2394), .Z(n2292) );
  NANDN U2542 ( .A(n2178), .B(n2177), .Z(n2182) );
  OR U2543 ( .A(n2180), .B(n2179), .Z(n2181) );
  AND U2544 ( .A(n2182), .B(n2181), .Z(n2290) );
  NANDN U2545 ( .A(n2184), .B(n2183), .Z(n2188) );
  OR U2546 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U2547 ( .A(n2188), .B(n2187), .Z(n2298) );
  NANDN U2548 ( .A(n29499), .B(n2189), .Z(n2191) );
  XOR U2549 ( .A(b[7]), .B(a[23]), .Z(n2376) );
  NANDN U2550 ( .A(n29735), .B(n2376), .Z(n2190) );
  AND U2551 ( .A(n2191), .B(n2190), .Z(n2308) );
  NANDN U2552 ( .A(n32996), .B(n2192), .Z(n2194) );
  XOR U2553 ( .A(b[21]), .B(a[9]), .Z(n2331) );
  NANDN U2554 ( .A(n33271), .B(n2331), .Z(n2193) );
  NAND U2555 ( .A(n2194), .B(n2193), .Z(n2307) );
  XNOR U2556 ( .A(n2308), .B(n2307), .Z(n2309) );
  NOR U2557 ( .A(n35340), .B(n2213), .Z(n2310) );
  XOR U2558 ( .A(n2309), .B(n2310), .Z(n2295) );
  NANDN U2559 ( .A(n28889), .B(n2195), .Z(n2197) );
  XOR U2560 ( .A(b[5]), .B(a[25]), .Z(n2355) );
  NANDN U2561 ( .A(n29138), .B(n2355), .Z(n2196) );
  AND U2562 ( .A(n2197), .B(n2196), .Z(n2316) );
  NANDN U2563 ( .A(n209), .B(n2198), .Z(n2200) );
  XOR U2564 ( .A(b[3]), .B(a[27]), .Z(n2358) );
  NANDN U2565 ( .A(n28941), .B(n2358), .Z(n2199) );
  AND U2566 ( .A(n2200), .B(n2199), .Z(n2314) );
  NANDN U2567 ( .A(n32013), .B(n2201), .Z(n2203) );
  XOR U2568 ( .A(b[17]), .B(a[13]), .Z(n2350) );
  NANDN U2569 ( .A(n32292), .B(n2350), .Z(n2202) );
  NAND U2570 ( .A(n2203), .B(n2202), .Z(n2313) );
  XNOR U2571 ( .A(n2314), .B(n2313), .Z(n2315) );
  XOR U2572 ( .A(n2316), .B(n2315), .Z(n2296) );
  XNOR U2573 ( .A(n2295), .B(n2296), .Z(n2297) );
  XNOR U2574 ( .A(n2298), .B(n2297), .Z(n2289) );
  XNOR U2575 ( .A(n2290), .B(n2289), .Z(n2291) );
  XOR U2576 ( .A(n2292), .B(n2291), .Z(n2398) );
  NANDN U2577 ( .A(n33866), .B(n2204), .Z(n2206) );
  XOR U2578 ( .A(b[23]), .B(a[7]), .Z(n2325) );
  NANDN U2579 ( .A(n33644), .B(n2325), .Z(n2205) );
  AND U2580 ( .A(n2206), .B(n2205), .Z(n2303) );
  NANDN U2581 ( .A(n33875), .B(n2207), .Z(n2209) );
  XOR U2582 ( .A(b[25]), .B(a[5]), .Z(n2328) );
  NANDN U2583 ( .A(n33994), .B(n2328), .Z(n2208) );
  AND U2584 ( .A(n2209), .B(n2208), .Z(n2302) );
  NANDN U2585 ( .A(n2210), .B(n30627), .Z(n2212) );
  XOR U2586 ( .A(b[9]), .B(a[21]), .Z(n2364) );
  NANDN U2587 ( .A(n30267), .B(n2364), .Z(n2211) );
  NAND U2588 ( .A(n2212), .B(n2211), .Z(n2301) );
  XOR U2589 ( .A(n2302), .B(n2301), .Z(n2304) );
  XOR U2590 ( .A(n2303), .B(n2304), .Z(n2341) );
  NANDN U2591 ( .A(n2214), .B(n2213), .Z(n2218) );
  OR U2592 ( .A(n2216), .B(n2215), .Z(n2217) );
  AND U2593 ( .A(n2218), .B(n2217), .Z(n2340) );
  XNOR U2594 ( .A(n2341), .B(n2340), .Z(n2342) );
  NANDN U2595 ( .A(n2220), .B(n2219), .Z(n2224) );
  OR U2596 ( .A(n2222), .B(n2221), .Z(n2223) );
  NAND U2597 ( .A(n2224), .B(n2223), .Z(n2343) );
  XNOR U2598 ( .A(n2342), .B(n2343), .Z(n2397) );
  XNOR U2599 ( .A(n2398), .B(n2397), .Z(n2399) );
  NANDN U2600 ( .A(n2226), .B(n2225), .Z(n2230) );
  NANDN U2601 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U2602 ( .A(n2230), .B(n2229), .Z(n2400) );
  XNOR U2603 ( .A(n2399), .B(n2400), .Z(n2286) );
  NANDN U2604 ( .A(n2232), .B(n2231), .Z(n2236) );
  NAND U2605 ( .A(n2234), .B(n2233), .Z(n2235) );
  AND U2606 ( .A(n2236), .B(n2235), .Z(n2284) );
  NANDN U2607 ( .A(n2238), .B(n2237), .Z(n2242) );
  NANDN U2608 ( .A(n2240), .B(n2239), .Z(n2241) );
  AND U2609 ( .A(n2242), .B(n2241), .Z(n2337) );
  NANDN U2610 ( .A(n2244), .B(n2243), .Z(n2248) );
  NAND U2611 ( .A(n2246), .B(n2245), .Z(n2247) );
  AND U2612 ( .A(n2248), .B(n2247), .Z(n2335) );
  NANDN U2613 ( .A(n2250), .B(n2249), .Z(n2254) );
  NANDN U2614 ( .A(n2252), .B(n2251), .Z(n2253) );
  NAND U2615 ( .A(n2254), .B(n2253), .Z(n2334) );
  XNOR U2616 ( .A(n2335), .B(n2334), .Z(n2336) );
  XNOR U2617 ( .A(n2337), .B(n2336), .Z(n2283) );
  XNOR U2618 ( .A(n2284), .B(n2283), .Z(n2285) );
  XOR U2619 ( .A(n2286), .B(n2285), .Z(n2404) );
  NANDN U2620 ( .A(n2256), .B(n2255), .Z(n2260) );
  OR U2621 ( .A(n2258), .B(n2257), .Z(n2259) );
  NAND U2622 ( .A(n2260), .B(n2259), .Z(n2403) );
  XOR U2623 ( .A(n2404), .B(n2403), .Z(n2406) );
  XOR U2624 ( .A(n2405), .B(n2406), .Z(n2278) );
  NANDN U2625 ( .A(n2262), .B(n2261), .Z(n2266) );
  NANDN U2626 ( .A(n2264), .B(n2263), .Z(n2265) );
  NAND U2627 ( .A(n2266), .B(n2265), .Z(n2277) );
  XNOR U2628 ( .A(n2278), .B(n2277), .Z(n2279) );
  XNOR U2629 ( .A(n2280), .B(n2279), .Z(n2272) );
  XNOR U2630 ( .A(sreg[93]), .B(n2272), .Z(n2274) );
  NANDN U2631 ( .A(sreg[92]), .B(n2267), .Z(n2271) );
  NAND U2632 ( .A(n2269), .B(n2268), .Z(n2270) );
  NAND U2633 ( .A(n2271), .B(n2270), .Z(n2273) );
  XNOR U2634 ( .A(n2274), .B(n2273), .Z(c[93]) );
  NANDN U2635 ( .A(sreg[93]), .B(n2272), .Z(n2276) );
  NAND U2636 ( .A(n2274), .B(n2273), .Z(n2275) );
  NAND U2637 ( .A(n2276), .B(n2275), .Z(n2547) );
  XNOR U2638 ( .A(sreg[94]), .B(n2547), .Z(n2549) );
  NANDN U2639 ( .A(n2278), .B(n2277), .Z(n2282) );
  NANDN U2640 ( .A(n2280), .B(n2279), .Z(n2281) );
  AND U2641 ( .A(n2282), .B(n2281), .Z(n2412) );
  NANDN U2642 ( .A(n2284), .B(n2283), .Z(n2288) );
  NAND U2643 ( .A(n2286), .B(n2285), .Z(n2287) );
  AND U2644 ( .A(n2288), .B(n2287), .Z(n2544) );
  NANDN U2645 ( .A(n2290), .B(n2289), .Z(n2294) );
  NAND U2646 ( .A(n2292), .B(n2291), .Z(n2293) );
  AND U2647 ( .A(n2294), .B(n2293), .Z(n2537) );
  NANDN U2648 ( .A(n2296), .B(n2295), .Z(n2300) );
  NANDN U2649 ( .A(n2298), .B(n2297), .Z(n2299) );
  AND U2650 ( .A(n2300), .B(n2299), .Z(n2536) );
  NANDN U2651 ( .A(n2302), .B(n2301), .Z(n2306) );
  OR U2652 ( .A(n2304), .B(n2303), .Z(n2305) );
  AND U2653 ( .A(n2306), .B(n2305), .Z(n2422) );
  NANDN U2654 ( .A(n2308), .B(n2307), .Z(n2312) );
  NAND U2655 ( .A(n2310), .B(n2309), .Z(n2311) );
  NAND U2656 ( .A(n2312), .B(n2311), .Z(n2421) );
  XNOR U2657 ( .A(n2422), .B(n2421), .Z(n2423) );
  NANDN U2658 ( .A(n2314), .B(n2313), .Z(n2318) );
  NANDN U2659 ( .A(n2316), .B(n2315), .Z(n2317) );
  AND U2660 ( .A(n2318), .B(n2317), .Z(n2466) );
  NAND U2661 ( .A(b[0]), .B(a[30]), .Z(n2319) );
  XNOR U2662 ( .A(b[1]), .B(n2319), .Z(n2321) );
  NANDN U2663 ( .A(b[0]), .B(a[29]), .Z(n2320) );
  NAND U2664 ( .A(n2321), .B(n2320), .Z(n2448) );
  XOR U2665 ( .A(b[30]), .B(b[29]), .Z(n35310) );
  IV U2666 ( .A(n35310), .Z(n35145) );
  ANDN U2667 ( .B(a[0]), .A(n35145), .Z(n2516) );
  IV U2668 ( .A(n34647), .Z(n34223) );
  NANDN U2669 ( .A(n34223), .B(n2322), .Z(n2324) );
  XOR U2670 ( .A(b[27]), .B(a[4]), .Z(n2481) );
  NANDN U2671 ( .A(n34458), .B(n2481), .Z(n2323) );
  AND U2672 ( .A(n2324), .B(n2323), .Z(n2446) );
  XNOR U2673 ( .A(n2516), .B(n2446), .Z(n2447) );
  XNOR U2674 ( .A(n2448), .B(n2447), .Z(n2463) );
  NANDN U2675 ( .A(n33866), .B(n2325), .Z(n2327) );
  XOR U2676 ( .A(b[23]), .B(a[8]), .Z(n2475) );
  NANDN U2677 ( .A(n33644), .B(n2475), .Z(n2326) );
  AND U2678 ( .A(n2327), .B(n2326), .Z(n2526) );
  NANDN U2679 ( .A(n33875), .B(n2328), .Z(n2330) );
  XOR U2680 ( .A(b[25]), .B(a[6]), .Z(n2478) );
  NANDN U2681 ( .A(n33994), .B(n2478), .Z(n2329) );
  AND U2682 ( .A(n2330), .B(n2329), .Z(n2524) );
  NANDN U2683 ( .A(n32996), .B(n2331), .Z(n2333) );
  XOR U2684 ( .A(b[21]), .B(a[10]), .Z(n2487) );
  NANDN U2685 ( .A(n33271), .B(n2487), .Z(n2332) );
  NAND U2686 ( .A(n2333), .B(n2332), .Z(n2523) );
  XNOR U2687 ( .A(n2524), .B(n2523), .Z(n2525) );
  XOR U2688 ( .A(n2526), .B(n2525), .Z(n2464) );
  XNOR U2689 ( .A(n2463), .B(n2464), .Z(n2465) );
  XOR U2690 ( .A(n2466), .B(n2465), .Z(n2424) );
  XNOR U2691 ( .A(n2423), .B(n2424), .Z(n2535) );
  XOR U2692 ( .A(n2536), .B(n2535), .Z(n2538) );
  XOR U2693 ( .A(n2537), .B(n2538), .Z(n2417) );
  NANDN U2694 ( .A(n2335), .B(n2334), .Z(n2339) );
  NANDN U2695 ( .A(n2337), .B(n2336), .Z(n2338) );
  AND U2696 ( .A(n2339), .B(n2338), .Z(n2416) );
  NANDN U2697 ( .A(n2341), .B(n2340), .Z(n2345) );
  NANDN U2698 ( .A(n2343), .B(n2342), .Z(n2344) );
  AND U2699 ( .A(n2345), .B(n2344), .Z(n2460) );
  XOR U2700 ( .A(b[28]), .B(b[29]), .Z(n2346) );
  ANDN U2701 ( .B(n2346), .A(n35002), .Z(n35001) );
  IV U2702 ( .A(n35001), .Z(n34634) );
  NANDN U2703 ( .A(n34634), .B(n2347), .Z(n2349) );
  XOR U2704 ( .A(b[29]), .B(a[2]), .Z(n2433) );
  NANDN U2705 ( .A(n34722), .B(n2433), .Z(n2348) );
  AND U2706 ( .A(n2349), .B(n2348), .Z(n2497) );
  NANDN U2707 ( .A(n32013), .B(n2350), .Z(n2352) );
  XOR U2708 ( .A(b[17]), .B(a[14]), .Z(n2512) );
  NANDN U2709 ( .A(n32292), .B(n2512), .Z(n2351) );
  NAND U2710 ( .A(n2352), .B(n2351), .Z(n2496) );
  XNOR U2711 ( .A(n2497), .B(n2496), .Z(n2499) );
  NOR U2712 ( .A(n2354), .B(n2353), .Z(n2498) );
  XOR U2713 ( .A(n2499), .B(n2498), .Z(n2469) );
  NANDN U2714 ( .A(n28889), .B(n2355), .Z(n2357) );
  XOR U2715 ( .A(b[5]), .B(a[26]), .Z(n2503) );
  NANDN U2716 ( .A(n29138), .B(n2503), .Z(n2356) );
  AND U2717 ( .A(n2357), .B(n2356), .Z(n2532) );
  NANDN U2718 ( .A(n209), .B(n2358), .Z(n2360) );
  XOR U2719 ( .A(b[3]), .B(a[28]), .Z(n2509) );
  NANDN U2720 ( .A(n28941), .B(n2509), .Z(n2359) );
  AND U2721 ( .A(n2360), .B(n2359), .Z(n2530) );
  NANDN U2722 ( .A(n2361), .B(n32023), .Z(n2363) );
  XOR U2723 ( .A(b[15]), .B(a[16]), .Z(n2443) );
  NANDN U2724 ( .A(n31925), .B(n2443), .Z(n2362) );
  NAND U2725 ( .A(n2363), .B(n2362), .Z(n2529) );
  XNOR U2726 ( .A(n2530), .B(n2529), .Z(n2531) );
  XOR U2727 ( .A(n2532), .B(n2531), .Z(n2470) );
  XNOR U2728 ( .A(n2469), .B(n2470), .Z(n2471) );
  NANDN U2729 ( .A(n210), .B(n2364), .Z(n2366) );
  XOR U2730 ( .A(b[9]), .B(a[22]), .Z(n2490) );
  NANDN U2731 ( .A(n30267), .B(n2490), .Z(n2365) );
  AND U2732 ( .A(n2366), .B(n2365), .Z(n2518) );
  NANDN U2733 ( .A(n30482), .B(n2367), .Z(n2369) );
  XOR U2734 ( .A(b[11]), .B(a[20]), .Z(n2493) );
  NANDN U2735 ( .A(n30891), .B(n2493), .Z(n2368) );
  NAND U2736 ( .A(n2369), .B(n2368), .Z(n2517) );
  XNOR U2737 ( .A(n2518), .B(n2517), .Z(n2519) );
  NANDN U2738 ( .A(n31055), .B(n2370), .Z(n2372) );
  XOR U2739 ( .A(b[13]), .B(a[18]), .Z(n2484) );
  NANDN U2740 ( .A(n31293), .B(n2484), .Z(n2371) );
  AND U2741 ( .A(n2372), .B(n2371), .Z(n2430) );
  NANDN U2742 ( .A(n32483), .B(n2373), .Z(n2375) );
  XOR U2743 ( .A(b[19]), .B(a[12]), .Z(n2506) );
  NANDN U2744 ( .A(n32823), .B(n2506), .Z(n2374) );
  AND U2745 ( .A(n2375), .B(n2374), .Z(n2428) );
  NANDN U2746 ( .A(n29499), .B(n2376), .Z(n2378) );
  XOR U2747 ( .A(b[7]), .B(a[24]), .Z(n2500) );
  NANDN U2748 ( .A(n29735), .B(n2500), .Z(n2377) );
  NAND U2749 ( .A(n2378), .B(n2377), .Z(n2427) );
  XNOR U2750 ( .A(n2428), .B(n2427), .Z(n2429) );
  XOR U2751 ( .A(n2430), .B(n2429), .Z(n2520) );
  XOR U2752 ( .A(n2519), .B(n2520), .Z(n2472) );
  XNOR U2753 ( .A(n2471), .B(n2472), .Z(n2454) );
  NANDN U2754 ( .A(n2380), .B(n2379), .Z(n2384) );
  NANDN U2755 ( .A(n2382), .B(n2381), .Z(n2383) );
  AND U2756 ( .A(n2384), .B(n2383), .Z(n2452) );
  NANDN U2757 ( .A(n2386), .B(n2385), .Z(n2390) );
  OR U2758 ( .A(n2388), .B(n2387), .Z(n2389) );
  AND U2759 ( .A(n2390), .B(n2389), .Z(n2451) );
  XNOR U2760 ( .A(n2452), .B(n2451), .Z(n2453) );
  XOR U2761 ( .A(n2454), .B(n2453), .Z(n2458) );
  NANDN U2762 ( .A(n2392), .B(n2391), .Z(n2396) );
  NANDN U2763 ( .A(n2394), .B(n2393), .Z(n2395) );
  AND U2764 ( .A(n2396), .B(n2395), .Z(n2457) );
  XNOR U2765 ( .A(n2458), .B(n2457), .Z(n2459) );
  XNOR U2766 ( .A(n2460), .B(n2459), .Z(n2415) );
  XOR U2767 ( .A(n2416), .B(n2415), .Z(n2418) );
  XOR U2768 ( .A(n2417), .B(n2418), .Z(n2542) );
  NANDN U2769 ( .A(n2398), .B(n2397), .Z(n2402) );
  NANDN U2770 ( .A(n2400), .B(n2399), .Z(n2401) );
  AND U2771 ( .A(n2402), .B(n2401), .Z(n2541) );
  XNOR U2772 ( .A(n2542), .B(n2541), .Z(n2543) );
  XOR U2773 ( .A(n2544), .B(n2543), .Z(n2410) );
  NANDN U2774 ( .A(n2404), .B(n2403), .Z(n2408) );
  OR U2775 ( .A(n2406), .B(n2405), .Z(n2407) );
  AND U2776 ( .A(n2408), .B(n2407), .Z(n2409) );
  XNOR U2777 ( .A(n2410), .B(n2409), .Z(n2411) );
  XNOR U2778 ( .A(n2412), .B(n2411), .Z(n2548) );
  XNOR U2779 ( .A(n2549), .B(n2548), .Z(c[94]) );
  NANDN U2780 ( .A(n2410), .B(n2409), .Z(n2414) );
  NANDN U2781 ( .A(n2412), .B(n2411), .Z(n2413) );
  AND U2782 ( .A(n2414), .B(n2413), .Z(n2560) );
  NANDN U2783 ( .A(n2416), .B(n2415), .Z(n2420) );
  OR U2784 ( .A(n2418), .B(n2417), .Z(n2419) );
  AND U2785 ( .A(n2420), .B(n2419), .Z(n2695) );
  NANDN U2786 ( .A(n2422), .B(n2421), .Z(n2426) );
  NANDN U2787 ( .A(n2424), .B(n2423), .Z(n2425) );
  AND U2788 ( .A(n2426), .B(n2425), .Z(n2572) );
  NANDN U2789 ( .A(n2428), .B(n2427), .Z(n2432) );
  NANDN U2790 ( .A(n2430), .B(n2429), .Z(n2431) );
  AND U2791 ( .A(n2432), .B(n2431), .Z(n2577) );
  NANDN U2792 ( .A(n34634), .B(n2433), .Z(n2435) );
  XOR U2793 ( .A(b[29]), .B(a[3]), .Z(n2587) );
  NANDN U2794 ( .A(n34722), .B(n2587), .Z(n2434) );
  AND U2795 ( .A(n2435), .B(n2434), .Z(n2662) );
  XOR U2796 ( .A(b[31]), .B(b[30]), .Z(n2667) );
  XOR U2797 ( .A(b[31]), .B(a[0]), .Z(n2436) );
  NAND U2798 ( .A(n2667), .B(n2436), .Z(n2437) );
  OR U2799 ( .A(n2437), .B(n35310), .Z(n2439) );
  XOR U2800 ( .A(b[31]), .B(a[1]), .Z(n2668) );
  NAND U2801 ( .A(n35310), .B(n2668), .Z(n2438) );
  AND U2802 ( .A(n2439), .B(n2438), .Z(n2663) );
  XOR U2803 ( .A(n2662), .B(n2663), .Z(n2616) );
  NAND U2804 ( .A(b[0]), .B(a[31]), .Z(n2440) );
  XNOR U2805 ( .A(b[1]), .B(n2440), .Z(n2442) );
  NANDN U2806 ( .A(b[0]), .B(a[30]), .Z(n2441) );
  NAND U2807 ( .A(n2442), .B(n2441), .Z(n2614) );
  NAND U2808 ( .A(n32023), .B(n2443), .Z(n2445) );
  XNOR U2809 ( .A(b[15]), .B(a[17]), .Z(n2596) );
  NANDN U2810 ( .A(n2596), .B(n32024), .Z(n2444) );
  NAND U2811 ( .A(n2445), .B(n2444), .Z(n2615) );
  XOR U2812 ( .A(n2614), .B(n2615), .Z(n2617) );
  XOR U2813 ( .A(n2616), .B(n2617), .Z(n2576) );
  NANDN U2814 ( .A(n2446), .B(n2516), .Z(n2450) );
  NANDN U2815 ( .A(n2448), .B(n2447), .Z(n2449) );
  NAND U2816 ( .A(n2450), .B(n2449), .Z(n2575) );
  XOR U2817 ( .A(n2576), .B(n2575), .Z(n2578) );
  XOR U2818 ( .A(n2577), .B(n2578), .Z(n2570) );
  NANDN U2819 ( .A(n2452), .B(n2451), .Z(n2456) );
  NAND U2820 ( .A(n2454), .B(n2453), .Z(n2455) );
  AND U2821 ( .A(n2456), .B(n2455), .Z(n2569) );
  XNOR U2822 ( .A(n2570), .B(n2569), .Z(n2571) );
  XOR U2823 ( .A(n2572), .B(n2571), .Z(n2565) );
  NANDN U2824 ( .A(n2458), .B(n2457), .Z(n2462) );
  NANDN U2825 ( .A(n2460), .B(n2459), .Z(n2461) );
  AND U2826 ( .A(n2462), .B(n2461), .Z(n2563) );
  NANDN U2827 ( .A(n2464), .B(n2463), .Z(n2468) );
  NANDN U2828 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U2829 ( .A(n2468), .B(n2467), .Z(n2687) );
  NANDN U2830 ( .A(n2470), .B(n2469), .Z(n2474) );
  NANDN U2831 ( .A(n2472), .B(n2471), .Z(n2473) );
  NAND U2832 ( .A(n2474), .B(n2473), .Z(n2686) );
  XNOR U2833 ( .A(n2687), .B(n2686), .Z(n2688) );
  NANDN U2834 ( .A(n33866), .B(n2475), .Z(n2477) );
  XOR U2835 ( .A(b[23]), .B(a[9]), .Z(n2671) );
  NANDN U2836 ( .A(n33644), .B(n2671), .Z(n2476) );
  AND U2837 ( .A(n2477), .B(n2476), .Z(n2646) );
  NANDN U2838 ( .A(n33875), .B(n2478), .Z(n2480) );
  XOR U2839 ( .A(b[25]), .B(a[7]), .Z(n2626) );
  NANDN U2840 ( .A(n33994), .B(n2626), .Z(n2479) );
  AND U2841 ( .A(n2480), .B(n2479), .Z(n2645) );
  NANDN U2842 ( .A(n34223), .B(n2481), .Z(n2483) );
  XOR U2843 ( .A(b[27]), .B(a[5]), .Z(n2629) );
  NANDN U2844 ( .A(n34458), .B(n2629), .Z(n2482) );
  NAND U2845 ( .A(n2483), .B(n2482), .Z(n2644) );
  XOR U2846 ( .A(n2645), .B(n2644), .Z(n2647) );
  XOR U2847 ( .A(n2646), .B(n2647), .Z(n2622) );
  NANDN U2848 ( .A(n31055), .B(n2484), .Z(n2486) );
  XOR U2849 ( .A(b[13]), .B(a[19]), .Z(n2599) );
  NANDN U2850 ( .A(n31293), .B(n2599), .Z(n2485) );
  AND U2851 ( .A(n2486), .B(n2485), .Z(n2604) );
  NANDN U2852 ( .A(n32996), .B(n2487), .Z(n2489) );
  XOR U2853 ( .A(b[21]), .B(a[11]), .Z(n2593) );
  NANDN U2854 ( .A(n33271), .B(n2593), .Z(n2488) );
  AND U2855 ( .A(n2489), .B(n2488), .Z(n2603) );
  NANDN U2856 ( .A(n210), .B(n2490), .Z(n2492) );
  XOR U2857 ( .A(b[9]), .B(a[23]), .Z(n2664) );
  NANDN U2858 ( .A(n30267), .B(n2664), .Z(n2491) );
  NAND U2859 ( .A(n2492), .B(n2491), .Z(n2602) );
  XOR U2860 ( .A(n2603), .B(n2602), .Z(n2605) );
  XOR U2861 ( .A(n2604), .B(n2605), .Z(n2621) );
  NAND U2862 ( .A(n31059), .B(n2493), .Z(n2495) );
  XNOR U2863 ( .A(b[11]), .B(a[21]), .Z(n2632) );
  NANDN U2864 ( .A(n2632), .B(n31060), .Z(n2494) );
  AND U2865 ( .A(n2495), .B(n2494), .Z(n2620) );
  XOR U2866 ( .A(n2621), .B(n2620), .Z(n2623) );
  XOR U2867 ( .A(n2622), .B(n2623), .Z(n2681) );
  NANDN U2868 ( .A(n29499), .B(n2500), .Z(n2502) );
  XOR U2869 ( .A(b[7]), .B(a[25]), .Z(n2635) );
  NANDN U2870 ( .A(n29735), .B(n2635), .Z(n2501) );
  AND U2871 ( .A(n2502), .B(n2501), .Z(n2653) );
  NANDN U2872 ( .A(n28889), .B(n2503), .Z(n2505) );
  XOR U2873 ( .A(b[5]), .B(a[27]), .Z(n2638) );
  NANDN U2874 ( .A(n29138), .B(n2638), .Z(n2504) );
  AND U2875 ( .A(n2505), .B(n2504), .Z(n2651) );
  NANDN U2876 ( .A(n32483), .B(n2506), .Z(n2508) );
  XOR U2877 ( .A(b[19]), .B(a[13]), .Z(n2641) );
  NANDN U2878 ( .A(n32823), .B(n2641), .Z(n2507) );
  NAND U2879 ( .A(n2508), .B(n2507), .Z(n2650) );
  XNOR U2880 ( .A(n2651), .B(n2650), .Z(n2652) );
  XNOR U2881 ( .A(n2653), .B(n2652), .Z(n2581) );
  NANDN U2882 ( .A(n209), .B(n2509), .Z(n2511) );
  XOR U2883 ( .A(b[3]), .B(a[29]), .Z(n2656) );
  NANDN U2884 ( .A(n28941), .B(n2656), .Z(n2510) );
  AND U2885 ( .A(n2511), .B(n2510), .Z(n2611) );
  NANDN U2886 ( .A(n32013), .B(n2512), .Z(n2514) );
  XOR U2887 ( .A(b[17]), .B(a[15]), .Z(n2659) );
  NANDN U2888 ( .A(n32292), .B(n2659), .Z(n2513) );
  AND U2889 ( .A(n2514), .B(n2513), .Z(n2609) );
  NAND U2890 ( .A(b[29]), .B(b[30]), .Z(n2515) );
  AND U2891 ( .A(b[31]), .B(n2515), .Z(n35581) );
  ANDN U2892 ( .B(n35581), .A(n2516), .Z(n2608) );
  XNOR U2893 ( .A(n2609), .B(n2608), .Z(n2610) );
  XOR U2894 ( .A(n2611), .B(n2610), .Z(n2582) );
  XNOR U2895 ( .A(n2581), .B(n2582), .Z(n2583) );
  XNOR U2896 ( .A(n2584), .B(n2583), .Z(n2680) );
  XNOR U2897 ( .A(n2681), .B(n2680), .Z(n2682) );
  NANDN U2898 ( .A(n2518), .B(n2517), .Z(n2522) );
  NANDN U2899 ( .A(n2520), .B(n2519), .Z(n2521) );
  AND U2900 ( .A(n2522), .B(n2521), .Z(n2677) );
  NANDN U2901 ( .A(n2524), .B(n2523), .Z(n2528) );
  NANDN U2902 ( .A(n2526), .B(n2525), .Z(n2527) );
  AND U2903 ( .A(n2528), .B(n2527), .Z(n2675) );
  NANDN U2904 ( .A(n2530), .B(n2529), .Z(n2534) );
  NANDN U2905 ( .A(n2532), .B(n2531), .Z(n2533) );
  NAND U2906 ( .A(n2534), .B(n2533), .Z(n2674) );
  XNOR U2907 ( .A(n2675), .B(n2674), .Z(n2676) );
  XOR U2908 ( .A(n2677), .B(n2676), .Z(n2683) );
  XOR U2909 ( .A(n2682), .B(n2683), .Z(n2689) );
  XOR U2910 ( .A(n2688), .B(n2689), .Z(n2564) );
  XOR U2911 ( .A(n2563), .B(n2564), .Z(n2566) );
  XOR U2912 ( .A(n2565), .B(n2566), .Z(n2693) );
  NANDN U2913 ( .A(n2536), .B(n2535), .Z(n2540) );
  OR U2914 ( .A(n2538), .B(n2537), .Z(n2539) );
  AND U2915 ( .A(n2540), .B(n2539), .Z(n2692) );
  XNOR U2916 ( .A(n2693), .B(n2692), .Z(n2694) );
  XNOR U2917 ( .A(n2695), .B(n2694), .Z(n2557) );
  NANDN U2918 ( .A(n2542), .B(n2541), .Z(n2546) );
  NAND U2919 ( .A(n2544), .B(n2543), .Z(n2545) );
  NAND U2920 ( .A(n2546), .B(n2545), .Z(n2558) );
  XNOR U2921 ( .A(n2557), .B(n2558), .Z(n2559) );
  XNOR U2922 ( .A(n2560), .B(n2559), .Z(n2552) );
  XNOR U2923 ( .A(sreg[95]), .B(n2552), .Z(n2554) );
  NANDN U2924 ( .A(sreg[94]), .B(n2547), .Z(n2551) );
  NAND U2925 ( .A(n2549), .B(n2548), .Z(n2550) );
  NAND U2926 ( .A(n2551), .B(n2550), .Z(n2553) );
  XNOR U2927 ( .A(n2554), .B(n2553), .Z(c[95]) );
  NANDN U2928 ( .A(sreg[95]), .B(n2552), .Z(n2556) );
  NAND U2929 ( .A(n2554), .B(n2553), .Z(n2555) );
  AND U2930 ( .A(n2556), .B(n2555), .Z(n2699) );
  NANDN U2931 ( .A(n2558), .B(n2557), .Z(n2562) );
  NANDN U2932 ( .A(n2560), .B(n2559), .Z(n2561) );
  AND U2933 ( .A(n2562), .B(n2561), .Z(n2704) );
  NANDN U2934 ( .A(n2564), .B(n2563), .Z(n2568) );
  OR U2935 ( .A(n2566), .B(n2565), .Z(n2567) );
  AND U2936 ( .A(n2568), .B(n2567), .Z(n2846) );
  NANDN U2937 ( .A(n2570), .B(n2569), .Z(n2574) );
  NAND U2938 ( .A(n2572), .B(n2571), .Z(n2573) );
  AND U2939 ( .A(n2574), .B(n2573), .Z(n2844) );
  NANDN U2940 ( .A(n2576), .B(n2575), .Z(n2580) );
  OR U2941 ( .A(n2578), .B(n2577), .Z(n2579) );
  AND U2942 ( .A(n2580), .B(n2579), .Z(n2739) );
  NANDN U2943 ( .A(n2582), .B(n2581), .Z(n2586) );
  NANDN U2944 ( .A(n2584), .B(n2583), .Z(n2585) );
  AND U2945 ( .A(n2586), .B(n2585), .Z(n2738) );
  XOR U2946 ( .A(b[32]), .B(b[31]), .Z(n35655) );
  IV U2947 ( .A(n35655), .Z(n35456) );
  ANDN U2948 ( .B(a[0]), .A(n35456), .Z(n2819) );
  NANDN U2949 ( .A(n34634), .B(n2587), .Z(n2589) );
  XOR U2950 ( .A(b[29]), .B(a[4]), .Z(n2823) );
  NANDN U2951 ( .A(n34722), .B(n2823), .Z(n2588) );
  AND U2952 ( .A(n2589), .B(n2588), .Z(n2755) );
  XNOR U2953 ( .A(n2819), .B(n2755), .Z(n2756) );
  NAND U2954 ( .A(b[0]), .B(a[32]), .Z(n2590) );
  XNOR U2955 ( .A(b[1]), .B(n2590), .Z(n2592) );
  NANDN U2956 ( .A(b[0]), .B(a[31]), .Z(n2591) );
  NAND U2957 ( .A(n2592), .B(n2591), .Z(n2757) );
  XNOR U2958 ( .A(n2756), .B(n2757), .Z(n2744) );
  NANDN U2959 ( .A(n32996), .B(n2593), .Z(n2595) );
  XOR U2960 ( .A(b[21]), .B(a[12]), .Z(n2785) );
  NANDN U2961 ( .A(n33271), .B(n2785), .Z(n2594) );
  AND U2962 ( .A(n2595), .B(n2594), .Z(n2828) );
  NANDN U2963 ( .A(n2596), .B(n32023), .Z(n2598) );
  XOR U2964 ( .A(b[15]), .B(a[18]), .Z(n2815) );
  NANDN U2965 ( .A(n31925), .B(n2815), .Z(n2597) );
  AND U2966 ( .A(n2598), .B(n2597), .Z(n2827) );
  NANDN U2967 ( .A(n31055), .B(n2599), .Z(n2601) );
  XOR U2968 ( .A(b[13]), .B(a[20]), .Z(n2800) );
  NANDN U2969 ( .A(n31293), .B(n2800), .Z(n2600) );
  NAND U2970 ( .A(n2601), .B(n2600), .Z(n2826) );
  XOR U2971 ( .A(n2827), .B(n2826), .Z(n2829) );
  XOR U2972 ( .A(n2828), .B(n2829), .Z(n2743) );
  XOR U2973 ( .A(n2744), .B(n2743), .Z(n2746) );
  NANDN U2974 ( .A(n2603), .B(n2602), .Z(n2607) );
  OR U2975 ( .A(n2605), .B(n2604), .Z(n2606) );
  NAND U2976 ( .A(n2607), .B(n2606), .Z(n2745) );
  XOR U2977 ( .A(n2746), .B(n2745), .Z(n2733) );
  NANDN U2978 ( .A(n2609), .B(n2608), .Z(n2613) );
  NANDN U2979 ( .A(n2611), .B(n2610), .Z(n2612) );
  AND U2980 ( .A(n2613), .B(n2612), .Z(n2732) );
  NANDN U2981 ( .A(n2615), .B(n2614), .Z(n2619) );
  OR U2982 ( .A(n2617), .B(n2616), .Z(n2618) );
  AND U2983 ( .A(n2619), .B(n2618), .Z(n2731) );
  XOR U2984 ( .A(n2732), .B(n2731), .Z(n2734) );
  XNOR U2985 ( .A(n2733), .B(n2734), .Z(n2737) );
  XOR U2986 ( .A(n2738), .B(n2737), .Z(n2740) );
  XOR U2987 ( .A(n2739), .B(n2740), .Z(n2715) );
  NANDN U2988 ( .A(n2621), .B(n2620), .Z(n2625) );
  OR U2989 ( .A(n2623), .B(n2622), .Z(n2624) );
  AND U2990 ( .A(n2625), .B(n2624), .Z(n2841) );
  NANDN U2991 ( .A(n33875), .B(n2626), .Z(n2628) );
  XOR U2992 ( .A(b[25]), .B(a[8]), .Z(n2782) );
  NANDN U2993 ( .A(n33994), .B(n2782), .Z(n2627) );
  AND U2994 ( .A(n2628), .B(n2627), .Z(n2834) );
  NANDN U2995 ( .A(n34223), .B(n2629), .Z(n2631) );
  XOR U2996 ( .A(b[27]), .B(a[6]), .Z(n2809) );
  NANDN U2997 ( .A(n34458), .B(n2809), .Z(n2630) );
  AND U2998 ( .A(n2631), .B(n2630), .Z(n2833) );
  NANDN U2999 ( .A(n2632), .B(n31059), .Z(n2634) );
  XOR U3000 ( .A(b[11]), .B(a[22]), .Z(n2797) );
  NANDN U3001 ( .A(n30891), .B(n2797), .Z(n2633) );
  NAND U3002 ( .A(n2634), .B(n2633), .Z(n2832) );
  XOR U3003 ( .A(n2833), .B(n2832), .Z(n2835) );
  XOR U3004 ( .A(n2834), .B(n2835), .Z(n2720) );
  NANDN U3005 ( .A(n29499), .B(n2635), .Z(n2637) );
  XOR U3006 ( .A(b[7]), .B(a[26]), .Z(n2806) );
  NANDN U3007 ( .A(n29735), .B(n2806), .Z(n2636) );
  AND U3008 ( .A(n2637), .B(n2636), .Z(n2762) );
  NANDN U3009 ( .A(n28889), .B(n2638), .Z(n2640) );
  XOR U3010 ( .A(b[5]), .B(a[28]), .Z(n2803) );
  NANDN U3011 ( .A(n29138), .B(n2803), .Z(n2639) );
  AND U3012 ( .A(n2640), .B(n2639), .Z(n2761) );
  NANDN U3013 ( .A(n32483), .B(n2641), .Z(n2643) );
  XNOR U3014 ( .A(b[19]), .B(a[14]), .Z(n2820) );
  NANDN U3015 ( .A(n2820), .B(n33001), .Z(n2642) );
  NAND U3016 ( .A(n2643), .B(n2642), .Z(n2760) );
  XOR U3017 ( .A(n2761), .B(n2760), .Z(n2763) );
  XNOR U3018 ( .A(n2762), .B(n2763), .Z(n2719) );
  XNOR U3019 ( .A(n2720), .B(n2719), .Z(n2722) );
  NANDN U3020 ( .A(n2645), .B(n2644), .Z(n2649) );
  OR U3021 ( .A(n2647), .B(n2646), .Z(n2648) );
  AND U3022 ( .A(n2649), .B(n2648), .Z(n2721) );
  XOR U3023 ( .A(n2722), .B(n2721), .Z(n2839) );
  NANDN U3024 ( .A(n2651), .B(n2650), .Z(n2655) );
  NANDN U3025 ( .A(n2653), .B(n2652), .Z(n2654) );
  AND U3026 ( .A(n2655), .B(n2654), .Z(n2728) );
  NANDN U3027 ( .A(n209), .B(n2656), .Z(n2658) );
  XOR U3028 ( .A(b[3]), .B(a[30]), .Z(n2812) );
  NANDN U3029 ( .A(n28941), .B(n2812), .Z(n2657) );
  AND U3030 ( .A(n2658), .B(n2657), .Z(n2789) );
  NANDN U3031 ( .A(n32013), .B(n2659), .Z(n2661) );
  XOR U3032 ( .A(b[17]), .B(a[16]), .Z(n2769) );
  NANDN U3033 ( .A(n32292), .B(n2769), .Z(n2660) );
  NAND U3034 ( .A(n2661), .B(n2660), .Z(n2788) );
  XNOR U3035 ( .A(n2789), .B(n2788), .Z(n2790) );
  OR U3036 ( .A(n2663), .B(n2662), .Z(n2791) );
  XNOR U3037 ( .A(n2790), .B(n2791), .Z(n2725) );
  NANDN U3038 ( .A(n210), .B(n2664), .Z(n2666) );
  XOR U3039 ( .A(b[9]), .B(a[24]), .Z(n2794) );
  NANDN U3040 ( .A(n30267), .B(n2794), .Z(n2665) );
  AND U3041 ( .A(n2666), .B(n2665), .Z(n2752) );
  ANDN U3042 ( .B(n2667), .A(n35310), .Z(n35309) );
  IV U3043 ( .A(n35309), .Z(n34909) );
  NANDN U3044 ( .A(n34909), .B(n2668), .Z(n2670) );
  XOR U3045 ( .A(b[31]), .B(a[2]), .Z(n2772) );
  NANDN U3046 ( .A(n35145), .B(n2772), .Z(n2669) );
  AND U3047 ( .A(n2670), .B(n2669), .Z(n2750) );
  NANDN U3048 ( .A(n33866), .B(n2671), .Z(n2673) );
  XOR U3049 ( .A(b[23]), .B(a[10]), .Z(n2779) );
  NANDN U3050 ( .A(n33644), .B(n2779), .Z(n2672) );
  NAND U3051 ( .A(n2673), .B(n2672), .Z(n2749) );
  XNOR U3052 ( .A(n2750), .B(n2749), .Z(n2751) );
  XOR U3053 ( .A(n2752), .B(n2751), .Z(n2726) );
  XNOR U3054 ( .A(n2725), .B(n2726), .Z(n2727) );
  XNOR U3055 ( .A(n2728), .B(n2727), .Z(n2838) );
  XNOR U3056 ( .A(n2839), .B(n2838), .Z(n2840) );
  XOR U3057 ( .A(n2841), .B(n2840), .Z(n2714) );
  NANDN U3058 ( .A(n2675), .B(n2674), .Z(n2679) );
  NANDN U3059 ( .A(n2677), .B(n2676), .Z(n2678) );
  AND U3060 ( .A(n2679), .B(n2678), .Z(n2713) );
  XOR U3061 ( .A(n2714), .B(n2713), .Z(n2716) );
  XOR U3062 ( .A(n2715), .B(n2716), .Z(n2710) );
  NANDN U3063 ( .A(n2681), .B(n2680), .Z(n2685) );
  NANDN U3064 ( .A(n2683), .B(n2682), .Z(n2684) );
  AND U3065 ( .A(n2685), .B(n2684), .Z(n2708) );
  NANDN U3066 ( .A(n2687), .B(n2686), .Z(n2691) );
  NANDN U3067 ( .A(n2689), .B(n2688), .Z(n2690) );
  NAND U3068 ( .A(n2691), .B(n2690), .Z(n2707) );
  XNOR U3069 ( .A(n2708), .B(n2707), .Z(n2709) );
  XOR U3070 ( .A(n2710), .B(n2709), .Z(n2845) );
  XOR U3071 ( .A(n2844), .B(n2845), .Z(n2847) );
  XOR U3072 ( .A(n2846), .B(n2847), .Z(n2702) );
  NANDN U3073 ( .A(n2693), .B(n2692), .Z(n2697) );
  NANDN U3074 ( .A(n2695), .B(n2694), .Z(n2696) );
  NAND U3075 ( .A(n2697), .B(n2696), .Z(n2701) );
  XNOR U3076 ( .A(n2702), .B(n2701), .Z(n2703) );
  XNOR U3077 ( .A(n2704), .B(n2703), .Z(n2700) );
  XNOR U3078 ( .A(sreg[96]), .B(n2700), .Z(n2698) );
  XOR U3079 ( .A(n2699), .B(n2698), .Z(c[96]) );
  NANDN U3080 ( .A(n2702), .B(n2701), .Z(n2706) );
  NANDN U3081 ( .A(n2704), .B(n2703), .Z(n2705) );
  AND U3082 ( .A(n2706), .B(n2705), .Z(n2858) );
  NANDN U3083 ( .A(n2708), .B(n2707), .Z(n2712) );
  NANDN U3084 ( .A(n2710), .B(n2709), .Z(n2711) );
  AND U3085 ( .A(n2712), .B(n2711), .Z(n3001) );
  NANDN U3086 ( .A(n2714), .B(n2713), .Z(n2718) );
  OR U3087 ( .A(n2716), .B(n2715), .Z(n2717) );
  AND U3088 ( .A(n2718), .B(n2717), .Z(n2863) );
  NANDN U3089 ( .A(n2720), .B(n2719), .Z(n2724) );
  NAND U3090 ( .A(n2722), .B(n2721), .Z(n2723) );
  AND U3091 ( .A(n2724), .B(n2723), .Z(n2944) );
  NANDN U3092 ( .A(n2726), .B(n2725), .Z(n2730) );
  NANDN U3093 ( .A(n2728), .B(n2727), .Z(n2729) );
  AND U3094 ( .A(n2730), .B(n2729), .Z(n2943) );
  XNOR U3095 ( .A(n2944), .B(n2943), .Z(n2945) );
  NANDN U3096 ( .A(n2732), .B(n2731), .Z(n2736) );
  NANDN U3097 ( .A(n2734), .B(n2733), .Z(n2735) );
  NAND U3098 ( .A(n2736), .B(n2735), .Z(n2946) );
  XNOR U3099 ( .A(n2945), .B(n2946), .Z(n2861) );
  NANDN U3100 ( .A(n2738), .B(n2737), .Z(n2742) );
  OR U3101 ( .A(n2740), .B(n2739), .Z(n2741) );
  NAND U3102 ( .A(n2742), .B(n2741), .Z(n2862) );
  XOR U3103 ( .A(n2861), .B(n2862), .Z(n2864) );
  XOR U3104 ( .A(n2863), .B(n2864), .Z(n3000) );
  NAND U3105 ( .A(n2744), .B(n2743), .Z(n2748) );
  NAND U3106 ( .A(n2746), .B(n2745), .Z(n2747) );
  AND U3107 ( .A(n2748), .B(n2747), .Z(n2993) );
  NANDN U3108 ( .A(n2750), .B(n2749), .Z(n2754) );
  NANDN U3109 ( .A(n2752), .B(n2751), .Z(n2753) );
  AND U3110 ( .A(n2754), .B(n2753), .Z(n2950) );
  NANDN U3111 ( .A(n2755), .B(n2819), .Z(n2759) );
  NANDN U3112 ( .A(n2757), .B(n2756), .Z(n2758) );
  NAND U3113 ( .A(n2759), .B(n2758), .Z(n2949) );
  XNOR U3114 ( .A(n2950), .B(n2949), .Z(n2952) );
  NANDN U3115 ( .A(n2761), .B(n2760), .Z(n2765) );
  OR U3116 ( .A(n2763), .B(n2762), .Z(n2764) );
  AND U3117 ( .A(n2765), .B(n2764), .Z(n2882) );
  NAND U3118 ( .A(b[0]), .B(a[33]), .Z(n2766) );
  XNOR U3119 ( .A(b[1]), .B(n2766), .Z(n2768) );
  NANDN U3120 ( .A(b[0]), .B(a[32]), .Z(n2767) );
  NAND U3121 ( .A(n2768), .B(n2767), .Z(n2988) );
  NANDN U3122 ( .A(n32013), .B(n2769), .Z(n2771) );
  XOR U3123 ( .A(b[17]), .B(a[17]), .Z(n2912) );
  NANDN U3124 ( .A(n32292), .B(n2912), .Z(n2770) );
  NAND U3125 ( .A(n2771), .B(n2770), .Z(n2987) );
  XNOR U3126 ( .A(n2988), .B(n2987), .Z(n2989) );
  NANDN U3127 ( .A(n34909), .B(n2772), .Z(n2774) );
  XOR U3128 ( .A(b[31]), .B(a[3]), .Z(n2961) );
  NANDN U3129 ( .A(n35145), .B(n2961), .Z(n2773) );
  AND U3130 ( .A(n2774), .B(n2773), .Z(n2973) );
  XOR U3131 ( .A(b[33]), .B(b[32]), .Z(n2918) );
  XOR U3132 ( .A(b[33]), .B(a[0]), .Z(n2775) );
  NAND U3133 ( .A(n2918), .B(n2775), .Z(n2776) );
  OR U3134 ( .A(n2776), .B(n35655), .Z(n2778) );
  XOR U3135 ( .A(b[33]), .B(a[1]), .Z(n2919) );
  NAND U3136 ( .A(n35655), .B(n2919), .Z(n2777) );
  NAND U3137 ( .A(n2778), .B(n2777), .Z(n2974) );
  XOR U3138 ( .A(n2973), .B(n2974), .Z(n2990) );
  XNOR U3139 ( .A(n2989), .B(n2990), .Z(n2879) );
  NANDN U3140 ( .A(n33866), .B(n2779), .Z(n2781) );
  XOR U3141 ( .A(b[23]), .B(a[11]), .Z(n2897) );
  NANDN U3142 ( .A(n33644), .B(n2897), .Z(n2780) );
  AND U3143 ( .A(n2781), .B(n2780), .Z(n2928) );
  NANDN U3144 ( .A(n33875), .B(n2782), .Z(n2784) );
  XOR U3145 ( .A(b[25]), .B(a[9]), .Z(n2885) );
  NANDN U3146 ( .A(n33994), .B(n2885), .Z(n2783) );
  AND U3147 ( .A(n2784), .B(n2783), .Z(n2926) );
  NANDN U3148 ( .A(n32996), .B(n2785), .Z(n2787) );
  XOR U3149 ( .A(b[21]), .B(a[13]), .Z(n2915) );
  NANDN U3150 ( .A(n33271), .B(n2915), .Z(n2786) );
  NAND U3151 ( .A(n2787), .B(n2786), .Z(n2925) );
  XNOR U3152 ( .A(n2926), .B(n2925), .Z(n2927) );
  XOR U3153 ( .A(n2928), .B(n2927), .Z(n2880) );
  XNOR U3154 ( .A(n2879), .B(n2880), .Z(n2881) );
  XNOR U3155 ( .A(n2882), .B(n2881), .Z(n2951) );
  XOR U3156 ( .A(n2952), .B(n2951), .Z(n2870) );
  NANDN U3157 ( .A(n2789), .B(n2788), .Z(n2793) );
  NANDN U3158 ( .A(n2791), .B(n2790), .Z(n2792) );
  AND U3159 ( .A(n2793), .B(n2792), .Z(n2867) );
  NAND U3160 ( .A(n30627), .B(n2794), .Z(n2796) );
  XNOR U3161 ( .A(b[9]), .B(a[25]), .Z(n2891) );
  NANDN U3162 ( .A(n2891), .B(n30628), .Z(n2795) );
  NAND U3163 ( .A(n2796), .B(n2795), .Z(n2937) );
  NANDN U3164 ( .A(n30482), .B(n2797), .Z(n2799) );
  XOR U3165 ( .A(b[11]), .B(a[23]), .Z(n2900) );
  NANDN U3166 ( .A(n30891), .B(n2900), .Z(n2798) );
  AND U3167 ( .A(n2799), .B(n2798), .Z(n2978) );
  NANDN U3168 ( .A(n31055), .B(n2800), .Z(n2802) );
  XOR U3169 ( .A(b[13]), .B(a[21]), .Z(n2894) );
  NANDN U3170 ( .A(n31293), .B(n2894), .Z(n2801) );
  AND U3171 ( .A(n2802), .B(n2801), .Z(n2976) );
  NANDN U3172 ( .A(n28889), .B(n2803), .Z(n2805) );
  XOR U3173 ( .A(b[5]), .B(a[29]), .Z(n2922) );
  NANDN U3174 ( .A(n29138), .B(n2922), .Z(n2804) );
  NAND U3175 ( .A(n2805), .B(n2804), .Z(n2975) );
  XNOR U3176 ( .A(n2976), .B(n2975), .Z(n2977) );
  XNOR U3177 ( .A(n2978), .B(n2977), .Z(n2938) );
  XOR U3178 ( .A(n2937), .B(n2938), .Z(n2940) );
  NANDN U3179 ( .A(n29499), .B(n2806), .Z(n2808) );
  XOR U3180 ( .A(b[7]), .B(a[27]), .Z(n2906) );
  NANDN U3181 ( .A(n29735), .B(n2906), .Z(n2807) );
  NAND U3182 ( .A(n2808), .B(n2807), .Z(n2939) );
  XOR U3183 ( .A(n2940), .B(n2939), .Z(n2876) );
  NANDN U3184 ( .A(n34223), .B(n2809), .Z(n2811) );
  XOR U3185 ( .A(b[27]), .B(a[7]), .Z(n2888) );
  NANDN U3186 ( .A(n34458), .B(n2888), .Z(n2810) );
  AND U3187 ( .A(n2811), .B(n2810), .Z(n2983) );
  NANDN U3188 ( .A(n209), .B(n2812), .Z(n2814) );
  XOR U3189 ( .A(b[3]), .B(a[31]), .Z(n2967) );
  NANDN U3190 ( .A(n28941), .B(n2967), .Z(n2813) );
  AND U3191 ( .A(n2814), .B(n2813), .Z(n2982) );
  NANDN U3192 ( .A(n31536), .B(n2815), .Z(n2817) );
  XOR U3193 ( .A(b[15]), .B(a[19]), .Z(n2903) );
  NANDN U3194 ( .A(n31925), .B(n2903), .Z(n2816) );
  NAND U3195 ( .A(n2817), .B(n2816), .Z(n2981) );
  XOR U3196 ( .A(n2982), .B(n2981), .Z(n2984) );
  XOR U3197 ( .A(n2983), .B(n2984), .Z(n2874) );
  NAND U3198 ( .A(b[31]), .B(b[32]), .Z(n2818) );
  AND U3199 ( .A(b[33]), .B(n2818), .Z(n35961) );
  ANDN U3200 ( .B(n35961), .A(n2819), .Z(n2932) );
  NANDN U3201 ( .A(n2820), .B(n33000), .Z(n2822) );
  XNOR U3202 ( .A(b[19]), .B(a[15]), .Z(n2970) );
  NANDN U3203 ( .A(n2970), .B(n33001), .Z(n2821) );
  NAND U3204 ( .A(n2822), .B(n2821), .Z(n2931) );
  XOR U3205 ( .A(n2932), .B(n2931), .Z(n2934) );
  NANDN U3206 ( .A(n34634), .B(n2823), .Z(n2825) );
  XOR U3207 ( .A(b[29]), .B(a[5]), .Z(n2909) );
  NANDN U3208 ( .A(n34722), .B(n2909), .Z(n2824) );
  NAND U3209 ( .A(n2825), .B(n2824), .Z(n2933) );
  XNOR U3210 ( .A(n2934), .B(n2933), .Z(n2873) );
  XNOR U3211 ( .A(n2874), .B(n2873), .Z(n2875) );
  XNOR U3212 ( .A(n2876), .B(n2875), .Z(n2957) );
  NANDN U3213 ( .A(n2827), .B(n2826), .Z(n2831) );
  OR U3214 ( .A(n2829), .B(n2828), .Z(n2830) );
  AND U3215 ( .A(n2831), .B(n2830), .Z(n2955) );
  NANDN U3216 ( .A(n2833), .B(n2832), .Z(n2837) );
  OR U3217 ( .A(n2835), .B(n2834), .Z(n2836) );
  NAND U3218 ( .A(n2837), .B(n2836), .Z(n2956) );
  XOR U3219 ( .A(n2955), .B(n2956), .Z(n2958) );
  XOR U3220 ( .A(n2957), .B(n2958), .Z(n2868) );
  XNOR U3221 ( .A(n2867), .B(n2868), .Z(n2869) );
  XOR U3222 ( .A(n2870), .B(n2869), .Z(n2994) );
  XNOR U3223 ( .A(n2993), .B(n2994), .Z(n2996) );
  NANDN U3224 ( .A(n2839), .B(n2838), .Z(n2843) );
  NAND U3225 ( .A(n2841), .B(n2840), .Z(n2842) );
  AND U3226 ( .A(n2843), .B(n2842), .Z(n2995) );
  XNOR U3227 ( .A(n2996), .B(n2995), .Z(n2999) );
  XOR U3228 ( .A(n3000), .B(n2999), .Z(n3002) );
  XOR U3229 ( .A(n3001), .B(n3002), .Z(n2856) );
  NANDN U3230 ( .A(n2845), .B(n2844), .Z(n2849) );
  OR U3231 ( .A(n2847), .B(n2846), .Z(n2848) );
  AND U3232 ( .A(n2849), .B(n2848), .Z(n2855) );
  XNOR U3233 ( .A(n2856), .B(n2855), .Z(n2857) );
  XNOR U3234 ( .A(n2858), .B(n2857), .Z(n2850) );
  XNOR U3235 ( .A(sreg[97]), .B(n2850), .Z(n2851) );
  XNOR U3236 ( .A(n2852), .B(n2851), .Z(c[97]) );
  NANDN U3237 ( .A(sreg[97]), .B(n2850), .Z(n2854) );
  NAND U3238 ( .A(n2852), .B(n2851), .Z(n2853) );
  NAND U3239 ( .A(n2854), .B(n2853), .Z(n3165) );
  XNOR U3240 ( .A(sreg[98]), .B(n3165), .Z(n3167) );
  NANDN U3241 ( .A(n2856), .B(n2855), .Z(n2860) );
  NANDN U3242 ( .A(n2858), .B(n2857), .Z(n2859) );
  AND U3243 ( .A(n2860), .B(n2859), .Z(n3008) );
  NANDN U3244 ( .A(n2862), .B(n2861), .Z(n2866) );
  OR U3245 ( .A(n2864), .B(n2863), .Z(n2865) );
  AND U3246 ( .A(n2866), .B(n2865), .Z(n3162) );
  NANDN U3247 ( .A(n2868), .B(n2867), .Z(n2872) );
  NANDN U3248 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3249 ( .A(n2872), .B(n2871), .Z(n3155) );
  NANDN U3250 ( .A(n2874), .B(n2873), .Z(n2878) );
  NANDN U3251 ( .A(n2876), .B(n2875), .Z(n2877) );
  AND U3252 ( .A(n2878), .B(n2877), .Z(n3014) );
  NANDN U3253 ( .A(n2880), .B(n2879), .Z(n2884) );
  NANDN U3254 ( .A(n2882), .B(n2881), .Z(n2883) );
  AND U3255 ( .A(n2884), .B(n2883), .Z(n3012) );
  NANDN U3256 ( .A(n33875), .B(n2885), .Z(n2887) );
  XOR U3257 ( .A(b[25]), .B(a[10]), .Z(n3059) );
  NANDN U3258 ( .A(n33994), .B(n3059), .Z(n2886) );
  AND U3259 ( .A(n2887), .B(n2886), .Z(n3079) );
  NANDN U3260 ( .A(n34223), .B(n2888), .Z(n2890) );
  XOR U3261 ( .A(b[27]), .B(a[8]), .Z(n3062) );
  NANDN U3262 ( .A(n34458), .B(n3062), .Z(n2889) );
  AND U3263 ( .A(n2890), .B(n2889), .Z(n3078) );
  NANDN U3264 ( .A(n2891), .B(n30627), .Z(n2893) );
  XOR U3265 ( .A(b[9]), .B(a[26]), .Z(n3065) );
  NANDN U3266 ( .A(n30267), .B(n3065), .Z(n2892) );
  NAND U3267 ( .A(n2893), .B(n2892), .Z(n3077) );
  XOR U3268 ( .A(n3078), .B(n3077), .Z(n3080) );
  XOR U3269 ( .A(n3079), .B(n3080), .Z(n3091) );
  NANDN U3270 ( .A(n31055), .B(n2894), .Z(n2896) );
  XOR U3271 ( .A(b[13]), .B(a[22]), .Z(n3129) );
  NANDN U3272 ( .A(n31293), .B(n3129), .Z(n2895) );
  AND U3273 ( .A(n2896), .B(n2895), .Z(n3049) );
  NANDN U3274 ( .A(n33866), .B(n2897), .Z(n2899) );
  XOR U3275 ( .A(b[23]), .B(a[12]), .Z(n3074) );
  NANDN U3276 ( .A(n33644), .B(n3074), .Z(n2898) );
  AND U3277 ( .A(n2899), .B(n2898), .Z(n3048) );
  NANDN U3278 ( .A(n30482), .B(n2900), .Z(n2902) );
  XOR U3279 ( .A(b[11]), .B(a[24]), .Z(n3132) );
  NANDN U3280 ( .A(n30891), .B(n3132), .Z(n2901) );
  NAND U3281 ( .A(n2902), .B(n2901), .Z(n3047) );
  XOR U3282 ( .A(n3048), .B(n3047), .Z(n3050) );
  XOR U3283 ( .A(n3049), .B(n3050), .Z(n3090) );
  NAND U3284 ( .A(n32023), .B(n2903), .Z(n2905) );
  XNOR U3285 ( .A(b[15]), .B(a[20]), .Z(n3126) );
  NANDN U3286 ( .A(n3126), .B(n32024), .Z(n2904) );
  AND U3287 ( .A(n2905), .B(n2904), .Z(n3089) );
  XOR U3288 ( .A(n3090), .B(n3089), .Z(n3092) );
  XNOR U3289 ( .A(n3091), .B(n3092), .Z(n3011) );
  XNOR U3290 ( .A(n3012), .B(n3011), .Z(n3013) );
  XOR U3291 ( .A(n3014), .B(n3013), .Z(n3154) );
  NANDN U3292 ( .A(n29499), .B(n2906), .Z(n2908) );
  XOR U3293 ( .A(b[7]), .B(a[28]), .Z(n3068) );
  NANDN U3294 ( .A(n29735), .B(n3068), .Z(n2907) );
  AND U3295 ( .A(n2908), .B(n2907), .Z(n3102) );
  NANDN U3296 ( .A(n34634), .B(n2909), .Z(n2911) );
  XOR U3297 ( .A(b[29]), .B(a[6]), .Z(n3071) );
  NANDN U3298 ( .A(n34722), .B(n3071), .Z(n2910) );
  AND U3299 ( .A(n2911), .B(n2910), .Z(n3101) );
  NANDN U3300 ( .A(n32013), .B(n2912), .Z(n2914) );
  XOR U3301 ( .A(b[17]), .B(a[18]), .Z(n3035) );
  NANDN U3302 ( .A(n32292), .B(n3035), .Z(n2913) );
  NAND U3303 ( .A(n2914), .B(n2913), .Z(n3100) );
  XOR U3304 ( .A(n3101), .B(n3100), .Z(n3103) );
  XOR U3305 ( .A(n3102), .B(n3103), .Z(n3018) );
  NAND U3306 ( .A(n33413), .B(n2915), .Z(n2917) );
  XNOR U3307 ( .A(b[21]), .B(a[14]), .Z(n3044) );
  NANDN U3308 ( .A(n3044), .B(n33414), .Z(n2916) );
  NAND U3309 ( .A(n2917), .B(n2916), .Z(n3054) );
  ANDN U3310 ( .B(n2918), .A(n35655), .Z(n35654) );
  IV U3311 ( .A(n35654), .Z(n35260) );
  NANDN U3312 ( .A(n35260), .B(n2919), .Z(n2921) );
  XOR U3313 ( .A(b[33]), .B(a[2]), .Z(n3112) );
  NANDN U3314 ( .A(n35456), .B(n3112), .Z(n2920) );
  NAND U3315 ( .A(n2921), .B(n2920), .Z(n3053) );
  XOR U3316 ( .A(n3054), .B(n3053), .Z(n3056) );
  NANDN U3317 ( .A(n28889), .B(n2922), .Z(n2924) );
  XOR U3318 ( .A(b[5]), .B(a[30]), .Z(n3038) );
  NANDN U3319 ( .A(n29138), .B(n3038), .Z(n2923) );
  NAND U3320 ( .A(n2924), .B(n2923), .Z(n3055) );
  XNOR U3321 ( .A(n3056), .B(n3055), .Z(n3017) );
  XNOR U3322 ( .A(n3018), .B(n3017), .Z(n3019) );
  NANDN U3323 ( .A(n2926), .B(n2925), .Z(n2930) );
  NANDN U3324 ( .A(n2928), .B(n2927), .Z(n2929) );
  NAND U3325 ( .A(n2930), .B(n2929), .Z(n3020) );
  XNOR U3326 ( .A(n3019), .B(n3020), .Z(n3135) );
  NAND U3327 ( .A(n2932), .B(n2931), .Z(n2936) );
  NAND U3328 ( .A(n2934), .B(n2933), .Z(n2935) );
  NAND U3329 ( .A(n2936), .B(n2935), .Z(n3136) );
  XNOR U3330 ( .A(n3135), .B(n3136), .Z(n3137) );
  NAND U3331 ( .A(n2938), .B(n2937), .Z(n2942) );
  NAND U3332 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3333 ( .A(n2942), .B(n2941), .Z(n3138) );
  XNOR U3334 ( .A(n3137), .B(n3138), .Z(n3153) );
  XOR U3335 ( .A(n3154), .B(n3153), .Z(n3156) );
  XOR U3336 ( .A(n3155), .B(n3156), .Z(n3149) );
  NANDN U3337 ( .A(n2944), .B(n2943), .Z(n2948) );
  NANDN U3338 ( .A(n2946), .B(n2945), .Z(n2947) );
  AND U3339 ( .A(n2948), .B(n2947), .Z(n3147) );
  NANDN U3340 ( .A(n2950), .B(n2949), .Z(n2954) );
  NAND U3341 ( .A(n2952), .B(n2951), .Z(n2953) );
  AND U3342 ( .A(n2954), .B(n2953), .Z(n3144) );
  NANDN U3343 ( .A(n2956), .B(n2955), .Z(n2960) );
  NANDN U3344 ( .A(n2958), .B(n2957), .Z(n2959) );
  AND U3345 ( .A(n2960), .B(n2959), .Z(n3141) );
  XOR U3346 ( .A(b[34]), .B(b[33]), .Z(n35929) );
  IV U3347 ( .A(n35929), .Z(n35801) );
  ANDN U3348 ( .B(a[0]), .A(n35801), .Z(n3122) );
  NANDN U3349 ( .A(n34909), .B(n2961), .Z(n2963) );
  XOR U3350 ( .A(b[31]), .B(a[4]), .Z(n3029) );
  NANDN U3351 ( .A(n35145), .B(n3029), .Z(n2962) );
  AND U3352 ( .A(n2963), .B(n2962), .Z(n3095) );
  XOR U3353 ( .A(n3122), .B(n3095), .Z(n3096) );
  NAND U3354 ( .A(b[0]), .B(a[34]), .Z(n2964) );
  XNOR U3355 ( .A(b[1]), .B(n2964), .Z(n2966) );
  NANDN U3356 ( .A(b[0]), .B(a[33]), .Z(n2965) );
  NAND U3357 ( .A(n2966), .B(n2965), .Z(n3097) );
  XOR U3358 ( .A(n3096), .B(n3097), .Z(n3024) );
  NANDN U3359 ( .A(n209), .B(n2967), .Z(n2969) );
  XOR U3360 ( .A(b[3]), .B(a[32]), .Z(n3041) );
  NANDN U3361 ( .A(n28941), .B(n3041), .Z(n2968) );
  AND U3362 ( .A(n2969), .B(n2968), .Z(n3107) );
  NANDN U3363 ( .A(n2970), .B(n33000), .Z(n2972) );
  XOR U3364 ( .A(b[19]), .B(a[16]), .Z(n3123) );
  NANDN U3365 ( .A(n32823), .B(n3123), .Z(n2971) );
  NAND U3366 ( .A(n2972), .B(n2971), .Z(n3106) );
  XNOR U3367 ( .A(n3107), .B(n3106), .Z(n3109) );
  ANDN U3368 ( .B(n2974), .A(n2973), .Z(n3108) );
  XNOR U3369 ( .A(n3109), .B(n3108), .Z(n3023) );
  XNOR U3370 ( .A(n3024), .B(n3023), .Z(n3026) );
  NANDN U3371 ( .A(n2976), .B(n2975), .Z(n2980) );
  NANDN U3372 ( .A(n2978), .B(n2977), .Z(n2979) );
  AND U3373 ( .A(n2980), .B(n2979), .Z(n3025) );
  XOR U3374 ( .A(n3026), .B(n3025), .Z(n3086) );
  NANDN U3375 ( .A(n2982), .B(n2981), .Z(n2986) );
  OR U3376 ( .A(n2984), .B(n2983), .Z(n2985) );
  AND U3377 ( .A(n2986), .B(n2985), .Z(n3084) );
  NANDN U3378 ( .A(n2988), .B(n2987), .Z(n2992) );
  NANDN U3379 ( .A(n2990), .B(n2989), .Z(n2991) );
  NAND U3380 ( .A(n2992), .B(n2991), .Z(n3083) );
  XNOR U3381 ( .A(n3084), .B(n3083), .Z(n3085) );
  XOR U3382 ( .A(n3086), .B(n3085), .Z(n3142) );
  XNOR U3383 ( .A(n3141), .B(n3142), .Z(n3143) );
  XOR U3384 ( .A(n3144), .B(n3143), .Z(n3148) );
  XOR U3385 ( .A(n3147), .B(n3148), .Z(n3150) );
  XOR U3386 ( .A(n3149), .B(n3150), .Z(n3160) );
  NANDN U3387 ( .A(n2994), .B(n2993), .Z(n2998) );
  NAND U3388 ( .A(n2996), .B(n2995), .Z(n2997) );
  NAND U3389 ( .A(n2998), .B(n2997), .Z(n3159) );
  XNOR U3390 ( .A(n3160), .B(n3159), .Z(n3161) );
  XNOR U3391 ( .A(n3162), .B(n3161), .Z(n3005) );
  NANDN U3392 ( .A(n3000), .B(n2999), .Z(n3004) );
  OR U3393 ( .A(n3002), .B(n3001), .Z(n3003) );
  NAND U3394 ( .A(n3004), .B(n3003), .Z(n3006) );
  XNOR U3395 ( .A(n3005), .B(n3006), .Z(n3007) );
  XNOR U3396 ( .A(n3008), .B(n3007), .Z(n3166) );
  XNOR U3397 ( .A(n3167), .B(n3166), .Z(c[98]) );
  NANDN U3398 ( .A(n3006), .B(n3005), .Z(n3010) );
  NANDN U3399 ( .A(n3008), .B(n3007), .Z(n3009) );
  AND U3400 ( .A(n3010), .B(n3009), .Z(n3175) );
  NANDN U3401 ( .A(n3012), .B(n3011), .Z(n3016) );
  NAND U3402 ( .A(n3014), .B(n3013), .Z(n3015) );
  AND U3403 ( .A(n3016), .B(n3015), .Z(n3187) );
  NANDN U3404 ( .A(n3018), .B(n3017), .Z(n3022) );
  NANDN U3405 ( .A(n3020), .B(n3019), .Z(n3021) );
  AND U3406 ( .A(n3022), .B(n3021), .Z(n3192) );
  NANDN U3407 ( .A(n3024), .B(n3023), .Z(n3028) );
  NAND U3408 ( .A(n3026), .B(n3025), .Z(n3027) );
  NAND U3409 ( .A(n3028), .B(n3027), .Z(n3191) );
  XNOR U3410 ( .A(n3192), .B(n3191), .Z(n3194) );
  NANDN U3411 ( .A(n34909), .B(n3029), .Z(n3031) );
  XOR U3412 ( .A(b[31]), .B(a[5]), .Z(n3251) );
  NANDN U3413 ( .A(n35145), .B(n3251), .Z(n3030) );
  AND U3414 ( .A(n3031), .B(n3030), .Z(n3283) );
  NAND U3415 ( .A(b[0]), .B(a[35]), .Z(n3032) );
  XNOR U3416 ( .A(b[1]), .B(n3032), .Z(n3034) );
  NANDN U3417 ( .A(b[0]), .B(a[34]), .Z(n3033) );
  NAND U3418 ( .A(n3034), .B(n3033), .Z(n3282) );
  NANDN U3419 ( .A(n32013), .B(n3035), .Z(n3037) );
  XOR U3420 ( .A(b[17]), .B(a[19]), .Z(n3206) );
  NANDN U3421 ( .A(n32292), .B(n3206), .Z(n3036) );
  NAND U3422 ( .A(n3037), .B(n3036), .Z(n3281) );
  XOR U3423 ( .A(n3282), .B(n3281), .Z(n3284) );
  XOR U3424 ( .A(n3283), .B(n3284), .Z(n3258) );
  NANDN U3425 ( .A(n28889), .B(n3038), .Z(n3040) );
  XOR U3426 ( .A(b[5]), .B(a[31]), .Z(n3218) );
  NANDN U3427 ( .A(n29138), .B(n3218), .Z(n3039) );
  AND U3428 ( .A(n3040), .B(n3039), .Z(n3289) );
  NANDN U3429 ( .A(n209), .B(n3041), .Z(n3043) );
  XOR U3430 ( .A(b[3]), .B(a[33]), .Z(n3245) );
  NANDN U3431 ( .A(n28941), .B(n3245), .Z(n3042) );
  AND U3432 ( .A(n3043), .B(n3042), .Z(n3288) );
  NANDN U3433 ( .A(n3044), .B(n33413), .Z(n3046) );
  XOR U3434 ( .A(b[21]), .B(a[15]), .Z(n3242) );
  NANDN U3435 ( .A(n33271), .B(n3242), .Z(n3045) );
  NAND U3436 ( .A(n3046), .B(n3045), .Z(n3287) );
  XOR U3437 ( .A(n3288), .B(n3287), .Z(n3290) );
  XNOR U3438 ( .A(n3289), .B(n3290), .Z(n3257) );
  XNOR U3439 ( .A(n3258), .B(n3257), .Z(n3259) );
  NANDN U3440 ( .A(n3048), .B(n3047), .Z(n3052) );
  OR U3441 ( .A(n3050), .B(n3049), .Z(n3051) );
  NAND U3442 ( .A(n3052), .B(n3051), .Z(n3260) );
  XNOR U3443 ( .A(n3259), .B(n3260), .Z(n3321) );
  NAND U3444 ( .A(n3054), .B(n3053), .Z(n3058) );
  NAND U3445 ( .A(n3056), .B(n3055), .Z(n3057) );
  AND U3446 ( .A(n3058), .B(n3057), .Z(n3320) );
  XOR U3447 ( .A(n3321), .B(n3320), .Z(n3323) );
  NANDN U3448 ( .A(n33875), .B(n3059), .Z(n3061) );
  XOR U3449 ( .A(b[25]), .B(a[11]), .Z(n3299) );
  NANDN U3450 ( .A(n33994), .B(n3299), .Z(n3060) );
  AND U3451 ( .A(n3061), .B(n3060), .Z(n3236) );
  NANDN U3452 ( .A(n34223), .B(n3062), .Z(n3064) );
  XOR U3453 ( .A(b[27]), .B(a[9]), .Z(n3302) );
  NANDN U3454 ( .A(n34458), .B(n3302), .Z(n3063) );
  AND U3455 ( .A(n3064), .B(n3063), .Z(n3235) );
  NANDN U3456 ( .A(n210), .B(n3065), .Z(n3067) );
  XOR U3457 ( .A(b[9]), .B(a[27]), .Z(n3209) );
  NANDN U3458 ( .A(n30267), .B(n3209), .Z(n3066) );
  NAND U3459 ( .A(n3067), .B(n3066), .Z(n3234) );
  XOR U3460 ( .A(n3235), .B(n3234), .Z(n3237) );
  XOR U3461 ( .A(n3236), .B(n3237), .Z(n3264) );
  NANDN U3462 ( .A(n29499), .B(n3068), .Z(n3070) );
  XOR U3463 ( .A(b[7]), .B(a[29]), .Z(n3305) );
  NANDN U3464 ( .A(n29735), .B(n3305), .Z(n3069) );
  AND U3465 ( .A(n3070), .B(n3069), .Z(n3230) );
  NANDN U3466 ( .A(n34634), .B(n3071), .Z(n3073) );
  XOR U3467 ( .A(b[29]), .B(a[7]), .Z(n3248) );
  NANDN U3468 ( .A(n34722), .B(n3248), .Z(n3072) );
  AND U3469 ( .A(n3073), .B(n3072), .Z(n3229) );
  NANDN U3470 ( .A(n33866), .B(n3074), .Z(n3076) );
  XOR U3471 ( .A(b[23]), .B(a[13]), .Z(n3225) );
  NANDN U3472 ( .A(n33644), .B(n3225), .Z(n3075) );
  NAND U3473 ( .A(n3076), .B(n3075), .Z(n3228) );
  XOR U3474 ( .A(n3229), .B(n3228), .Z(n3231) );
  XNOR U3475 ( .A(n3230), .B(n3231), .Z(n3263) );
  XNOR U3476 ( .A(n3264), .B(n3263), .Z(n3266) );
  NANDN U3477 ( .A(n3078), .B(n3077), .Z(n3082) );
  OR U3478 ( .A(n3080), .B(n3079), .Z(n3081) );
  AND U3479 ( .A(n3082), .B(n3081), .Z(n3265) );
  XOR U3480 ( .A(n3266), .B(n3265), .Z(n3322) );
  XOR U3481 ( .A(n3323), .B(n3322), .Z(n3193) );
  XOR U3482 ( .A(n3194), .B(n3193), .Z(n3186) );
  NANDN U3483 ( .A(n3084), .B(n3083), .Z(n3088) );
  NANDN U3484 ( .A(n3086), .B(n3085), .Z(n3087) );
  AND U3485 ( .A(n3088), .B(n3087), .Z(n3317) );
  NANDN U3486 ( .A(n3090), .B(n3089), .Z(n3094) );
  OR U3487 ( .A(n3092), .B(n3091), .Z(n3093) );
  AND U3488 ( .A(n3094), .B(n3093), .Z(n3314) );
  NANDN U3489 ( .A(n3095), .B(n3122), .Z(n3099) );
  OR U3490 ( .A(n3097), .B(n3096), .Z(n3098) );
  AND U3491 ( .A(n3099), .B(n3098), .Z(n3270) );
  NANDN U3492 ( .A(n3101), .B(n3100), .Z(n3105) );
  OR U3493 ( .A(n3103), .B(n3102), .Z(n3104) );
  NAND U3494 ( .A(n3105), .B(n3104), .Z(n3269) );
  XNOR U3495 ( .A(n3270), .B(n3269), .Z(n3271) );
  NANDN U3496 ( .A(n3107), .B(n3106), .Z(n3111) );
  NAND U3497 ( .A(n3109), .B(n3108), .Z(n3110) );
  AND U3498 ( .A(n3111), .B(n3110), .Z(n3311) );
  NANDN U3499 ( .A(n35260), .B(n3112), .Z(n3114) );
  XOR U3500 ( .A(b[33]), .B(a[3]), .Z(n3296) );
  NANDN U3501 ( .A(n35456), .B(n3296), .Z(n3113) );
  AND U3502 ( .A(n3114), .B(n3113), .Z(n3240) );
  XOR U3503 ( .A(b[35]), .B(a[1]), .Z(n3222) );
  NANDN U3504 ( .A(n35801), .B(n3222), .Z(n3121) );
  ANDN U3505 ( .B(b[34]), .A(b[35]), .Z(n3115) );
  NAND U3506 ( .A(n3115), .B(a[0]), .Z(n3118) );
  NAND U3507 ( .A(b[33]), .B(b[34]), .Z(n3116) );
  AND U3508 ( .A(b[35]), .B(n3116), .Z(n36182) );
  NANDN U3509 ( .A(a[0]), .B(n36182), .Z(n3117) );
  NAND U3510 ( .A(n3118), .B(n3117), .Z(n3119) );
  NAND U3511 ( .A(n35801), .B(n3119), .Z(n3120) );
  AND U3512 ( .A(n3121), .B(n3120), .Z(n3241) );
  XOR U3513 ( .A(n3240), .B(n3241), .Z(n3214) );
  ANDN U3514 ( .B(n36182), .A(n3122), .Z(n3213) );
  NAND U3515 ( .A(n33000), .B(n3123), .Z(n3125) );
  XNOR U3516 ( .A(b[19]), .B(a[17]), .Z(n3254) );
  NANDN U3517 ( .A(n3254), .B(n33001), .Z(n3124) );
  AND U3518 ( .A(n3125), .B(n3124), .Z(n3212) );
  XOR U3519 ( .A(n3213), .B(n3212), .Z(n3215) );
  XOR U3520 ( .A(n3214), .B(n3215), .Z(n3309) );
  NANDN U3521 ( .A(n3126), .B(n32023), .Z(n3128) );
  XOR U3522 ( .A(b[15]), .B(a[21]), .Z(n3203) );
  NANDN U3523 ( .A(n31925), .B(n3203), .Z(n3127) );
  AND U3524 ( .A(n3128), .B(n3127), .Z(n3278) );
  NANDN U3525 ( .A(n31055), .B(n3129), .Z(n3131) );
  XOR U3526 ( .A(b[13]), .B(a[23]), .Z(n3200) );
  NANDN U3527 ( .A(n31293), .B(n3200), .Z(n3130) );
  AND U3528 ( .A(n3131), .B(n3130), .Z(n3276) );
  NANDN U3529 ( .A(n30482), .B(n3132), .Z(n3134) );
  XOR U3530 ( .A(b[11]), .B(a[25]), .Z(n3197) );
  NANDN U3531 ( .A(n30891), .B(n3197), .Z(n3133) );
  NAND U3532 ( .A(n3134), .B(n3133), .Z(n3275) );
  XNOR U3533 ( .A(n3276), .B(n3275), .Z(n3277) );
  XNOR U3534 ( .A(n3278), .B(n3277), .Z(n3308) );
  XNOR U3535 ( .A(n3309), .B(n3308), .Z(n3310) );
  XOR U3536 ( .A(n3311), .B(n3310), .Z(n3272) );
  XOR U3537 ( .A(n3271), .B(n3272), .Z(n3315) );
  XNOR U3538 ( .A(n3314), .B(n3315), .Z(n3316) );
  XNOR U3539 ( .A(n3317), .B(n3316), .Z(n3185) );
  XOR U3540 ( .A(n3186), .B(n3185), .Z(n3188) );
  XOR U3541 ( .A(n3187), .B(n3188), .Z(n3181) );
  NANDN U3542 ( .A(n3136), .B(n3135), .Z(n3140) );
  NANDN U3543 ( .A(n3138), .B(n3137), .Z(n3139) );
  AND U3544 ( .A(n3140), .B(n3139), .Z(n3180) );
  NANDN U3545 ( .A(n3142), .B(n3141), .Z(n3146) );
  NANDN U3546 ( .A(n3144), .B(n3143), .Z(n3145) );
  AND U3547 ( .A(n3146), .B(n3145), .Z(n3179) );
  XOR U3548 ( .A(n3180), .B(n3179), .Z(n3182) );
  XOR U3549 ( .A(n3181), .B(n3182), .Z(n3328) );
  NANDN U3550 ( .A(n3148), .B(n3147), .Z(n3152) );
  OR U3551 ( .A(n3150), .B(n3149), .Z(n3151) );
  AND U3552 ( .A(n3152), .B(n3151), .Z(n3327) );
  NANDN U3553 ( .A(n3154), .B(n3153), .Z(n3158) );
  OR U3554 ( .A(n3156), .B(n3155), .Z(n3157) );
  AND U3555 ( .A(n3158), .B(n3157), .Z(n3326) );
  XOR U3556 ( .A(n3327), .B(n3326), .Z(n3329) );
  XOR U3557 ( .A(n3328), .B(n3329), .Z(n3174) );
  NANDN U3558 ( .A(n3160), .B(n3159), .Z(n3164) );
  NANDN U3559 ( .A(n3162), .B(n3161), .Z(n3163) );
  NAND U3560 ( .A(n3164), .B(n3163), .Z(n3173) );
  XOR U3561 ( .A(n3174), .B(n3173), .Z(n3176) );
  XOR U3562 ( .A(n3175), .B(n3176), .Z(n3171) );
  NANDN U3563 ( .A(sreg[98]), .B(n3165), .Z(n3169) );
  NAND U3564 ( .A(n3167), .B(n3166), .Z(n3168) );
  AND U3565 ( .A(n3169), .B(n3168), .Z(n3172) );
  XNOR U3566 ( .A(sreg[99]), .B(n3172), .Z(n3170) );
  XOR U3567 ( .A(n3171), .B(n3170), .Z(c[99]) );
  XOR U3568 ( .A(sreg[100]), .B(n3499), .Z(n3501) );
  NANDN U3569 ( .A(n3174), .B(n3173), .Z(n3178) );
  OR U3570 ( .A(n3176), .B(n3175), .Z(n3177) );
  AND U3571 ( .A(n3178), .B(n3177), .Z(n3335) );
  NANDN U3572 ( .A(n3180), .B(n3179), .Z(n3184) );
  OR U3573 ( .A(n3182), .B(n3181), .Z(n3183) );
  AND U3574 ( .A(n3184), .B(n3183), .Z(n3496) );
  NANDN U3575 ( .A(n3186), .B(n3185), .Z(n3190) );
  OR U3576 ( .A(n3188), .B(n3187), .Z(n3189) );
  AND U3577 ( .A(n3190), .B(n3189), .Z(n3494) );
  NANDN U3578 ( .A(n3192), .B(n3191), .Z(n3196) );
  NAND U3579 ( .A(n3194), .B(n3193), .Z(n3195) );
  AND U3580 ( .A(n3196), .B(n3195), .Z(n3489) );
  NANDN U3581 ( .A(n30482), .B(n3197), .Z(n3199) );
  XOR U3582 ( .A(b[11]), .B(a[26]), .Z(n3380) );
  NANDN U3583 ( .A(n30891), .B(n3380), .Z(n3198) );
  AND U3584 ( .A(n3199), .B(n3198), .Z(n3357) );
  NANDN U3585 ( .A(n31055), .B(n3200), .Z(n3202) );
  XOR U3586 ( .A(b[13]), .B(a[24]), .Z(n3389) );
  NANDN U3587 ( .A(n31293), .B(n3389), .Z(n3201) );
  NAND U3588 ( .A(n3202), .B(n3201), .Z(n3356) );
  XNOR U3589 ( .A(n3357), .B(n3356), .Z(n3359) );
  NANDN U3590 ( .A(n31536), .B(n3203), .Z(n3205) );
  XOR U3591 ( .A(b[15]), .B(a[22]), .Z(n3392) );
  NANDN U3592 ( .A(n31925), .B(n3392), .Z(n3204) );
  AND U3593 ( .A(n3205), .B(n3204), .Z(n3478) );
  NANDN U3594 ( .A(n32013), .B(n3206), .Z(n3208) );
  XOR U3595 ( .A(b[17]), .B(a[20]), .Z(n3407) );
  NANDN U3596 ( .A(n32292), .B(n3407), .Z(n3207) );
  AND U3597 ( .A(n3208), .B(n3207), .Z(n3476) );
  NANDN U3598 ( .A(n210), .B(n3209), .Z(n3211) );
  XOR U3599 ( .A(b[9]), .B(a[28]), .Z(n3395) );
  NANDN U3600 ( .A(n30267), .B(n3395), .Z(n3210) );
  NAND U3601 ( .A(n3211), .B(n3210), .Z(n3475) );
  XNOR U3602 ( .A(n3476), .B(n3475), .Z(n3477) );
  XNOR U3603 ( .A(n3478), .B(n3477), .Z(n3358) );
  XOR U3604 ( .A(n3359), .B(n3358), .Z(n3439) );
  NANDN U3605 ( .A(n3213), .B(n3212), .Z(n3217) );
  OR U3606 ( .A(n3215), .B(n3214), .Z(n3216) );
  AND U3607 ( .A(n3217), .B(n3216), .Z(n3438) );
  NANDN U3608 ( .A(n28889), .B(n3218), .Z(n3220) );
  XOR U3609 ( .A(b[5]), .B(a[32]), .Z(n3463) );
  NANDN U3610 ( .A(n29138), .B(n3463), .Z(n3219) );
  AND U3611 ( .A(n3220), .B(n3219), .Z(n3370) );
  XOR U3612 ( .A(b[34]), .B(b[35]), .Z(n3221) );
  ANDN U3613 ( .B(n3221), .A(n35929), .Z(n35928) );
  IV U3614 ( .A(n35928), .Z(n35611) );
  NANDN U3615 ( .A(n35611), .B(n3222), .Z(n3224) );
  XOR U3616 ( .A(b[35]), .B(a[2]), .Z(n3448) );
  NANDN U3617 ( .A(n35801), .B(n3448), .Z(n3223) );
  AND U3618 ( .A(n3224), .B(n3223), .Z(n3369) );
  NANDN U3619 ( .A(n33866), .B(n3225), .Z(n3227) );
  XOR U3620 ( .A(b[23]), .B(a[14]), .Z(n3466) );
  NANDN U3621 ( .A(n33644), .B(n3466), .Z(n3226) );
  NAND U3622 ( .A(n3227), .B(n3226), .Z(n3368) );
  XOR U3623 ( .A(n3369), .B(n3368), .Z(n3371) );
  XNOR U3624 ( .A(n3370), .B(n3371), .Z(n3437) );
  XOR U3625 ( .A(n3438), .B(n3437), .Z(n3440) );
  XOR U3626 ( .A(n3439), .B(n3440), .Z(n3433) );
  NANDN U3627 ( .A(n3229), .B(n3228), .Z(n3233) );
  OR U3628 ( .A(n3231), .B(n3230), .Z(n3232) );
  AND U3629 ( .A(n3233), .B(n3232), .Z(n3432) );
  NANDN U3630 ( .A(n3235), .B(n3234), .Z(n3239) );
  OR U3631 ( .A(n3237), .B(n3236), .Z(n3238) );
  AND U3632 ( .A(n3239), .B(n3238), .Z(n3422) );
  NOR U3633 ( .A(n3241), .B(n3240), .Z(n3471) );
  NAND U3634 ( .A(n33413), .B(n3242), .Z(n3244) );
  XNOR U3635 ( .A(b[21]), .B(a[16]), .Z(n3383) );
  NANDN U3636 ( .A(n3383), .B(n33414), .Z(n3243) );
  AND U3637 ( .A(n3244), .B(n3243), .Z(n3469) );
  NAND U3638 ( .A(n9942), .B(n3245), .Z(n3247) );
  XNOR U3639 ( .A(b[3]), .B(a[34]), .Z(n3404) );
  NANDN U3640 ( .A(n3404), .B(n9653), .Z(n3246) );
  NAND U3641 ( .A(n3247), .B(n3246), .Z(n3470) );
  XOR U3642 ( .A(n3469), .B(n3470), .Z(n3472) );
  XOR U3643 ( .A(n3471), .B(n3472), .Z(n3420) );
  NANDN U3644 ( .A(n34634), .B(n3248), .Z(n3250) );
  XOR U3645 ( .A(b[29]), .B(a[8]), .Z(n3374) );
  NANDN U3646 ( .A(n34722), .B(n3374), .Z(n3249) );
  AND U3647 ( .A(n3250), .B(n3249), .Z(n3365) );
  NANDN U3648 ( .A(n34909), .B(n3251), .Z(n3253) );
  XOR U3649 ( .A(b[31]), .B(a[6]), .Z(n3377) );
  NANDN U3650 ( .A(n35145), .B(n3377), .Z(n3252) );
  AND U3651 ( .A(n3253), .B(n3252), .Z(n3363) );
  NANDN U3652 ( .A(n3254), .B(n33000), .Z(n3256) );
  XOR U3653 ( .A(b[19]), .B(a[18]), .Z(n3457) );
  NANDN U3654 ( .A(n32823), .B(n3457), .Z(n3255) );
  NAND U3655 ( .A(n3256), .B(n3255), .Z(n3362) );
  XNOR U3656 ( .A(n3363), .B(n3362), .Z(n3364) );
  XNOR U3657 ( .A(n3365), .B(n3364), .Z(n3419) );
  XNOR U3658 ( .A(n3420), .B(n3419), .Z(n3421) );
  XNOR U3659 ( .A(n3422), .B(n3421), .Z(n3431) );
  XOR U3660 ( .A(n3432), .B(n3431), .Z(n3434) );
  XOR U3661 ( .A(n3433), .B(n3434), .Z(n3353) );
  NANDN U3662 ( .A(n3258), .B(n3257), .Z(n3262) );
  NANDN U3663 ( .A(n3260), .B(n3259), .Z(n3261) );
  AND U3664 ( .A(n3262), .B(n3261), .Z(n3351) );
  NANDN U3665 ( .A(n3264), .B(n3263), .Z(n3268) );
  NAND U3666 ( .A(n3266), .B(n3265), .Z(n3267) );
  NAND U3667 ( .A(n3268), .B(n3267), .Z(n3350) );
  XNOR U3668 ( .A(n3351), .B(n3350), .Z(n3352) );
  XNOR U3669 ( .A(n3353), .B(n3352), .Z(n3487) );
  NANDN U3670 ( .A(n3270), .B(n3269), .Z(n3274) );
  NANDN U3671 ( .A(n3272), .B(n3271), .Z(n3273) );
  AND U3672 ( .A(n3274), .B(n3273), .Z(n3346) );
  NANDN U3673 ( .A(n3276), .B(n3275), .Z(n3280) );
  NANDN U3674 ( .A(n3278), .B(n3277), .Z(n3279) );
  AND U3675 ( .A(n3280), .B(n3279), .Z(n3482) );
  NANDN U3676 ( .A(n3282), .B(n3281), .Z(n3286) );
  OR U3677 ( .A(n3284), .B(n3283), .Z(n3285) );
  NAND U3678 ( .A(n3286), .B(n3285), .Z(n3481) );
  XNOR U3679 ( .A(n3482), .B(n3481), .Z(n3484) );
  NANDN U3680 ( .A(n3288), .B(n3287), .Z(n3292) );
  OR U3681 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U3682 ( .A(n3292), .B(n3291), .Z(n3427) );
  NAND U3683 ( .A(b[0]), .B(a[36]), .Z(n3293) );
  XNOR U3684 ( .A(b[1]), .B(n3293), .Z(n3295) );
  NANDN U3685 ( .A(b[0]), .B(a[35]), .Z(n3294) );
  NAND U3686 ( .A(n3295), .B(n3294), .Z(n3445) );
  XOR U3687 ( .A(b[36]), .B(b[35]), .Z(n36239) );
  IV U3688 ( .A(n36239), .Z(n36047) );
  ANDN U3689 ( .B(a[0]), .A(n36047), .Z(n3456) );
  NANDN U3690 ( .A(n35260), .B(n3296), .Z(n3298) );
  XOR U3691 ( .A(b[33]), .B(a[4]), .Z(n3398) );
  NANDN U3692 ( .A(n35456), .B(n3398), .Z(n3297) );
  AND U3693 ( .A(n3298), .B(n3297), .Z(n3443) );
  XNOR U3694 ( .A(n3456), .B(n3443), .Z(n3444) );
  XNOR U3695 ( .A(n3445), .B(n3444), .Z(n3426) );
  NANDN U3696 ( .A(n33875), .B(n3299), .Z(n3301) );
  XOR U3697 ( .A(b[25]), .B(a[12]), .Z(n3386) );
  NANDN U3698 ( .A(n33994), .B(n3386), .Z(n3300) );
  AND U3699 ( .A(n3301), .B(n3300), .Z(n3415) );
  NANDN U3700 ( .A(n34223), .B(n3302), .Z(n3304) );
  XOR U3701 ( .A(b[27]), .B(a[10]), .Z(n3401) );
  NANDN U3702 ( .A(n34458), .B(n3401), .Z(n3303) );
  AND U3703 ( .A(n3304), .B(n3303), .Z(n3414) );
  NANDN U3704 ( .A(n29499), .B(n3305), .Z(n3307) );
  XOR U3705 ( .A(b[7]), .B(a[30]), .Z(n3460) );
  NANDN U3706 ( .A(n29735), .B(n3460), .Z(n3306) );
  NAND U3707 ( .A(n3307), .B(n3306), .Z(n3413) );
  XOR U3708 ( .A(n3414), .B(n3413), .Z(n3416) );
  XOR U3709 ( .A(n3415), .B(n3416), .Z(n3425) );
  XOR U3710 ( .A(n3426), .B(n3425), .Z(n3428) );
  XOR U3711 ( .A(n3427), .B(n3428), .Z(n3483) );
  XOR U3712 ( .A(n3484), .B(n3483), .Z(n3345) );
  NANDN U3713 ( .A(n3309), .B(n3308), .Z(n3313) );
  NANDN U3714 ( .A(n3311), .B(n3310), .Z(n3312) );
  AND U3715 ( .A(n3313), .B(n3312), .Z(n3344) );
  XOR U3716 ( .A(n3345), .B(n3344), .Z(n3347) );
  XOR U3717 ( .A(n3346), .B(n3347), .Z(n3488) );
  XOR U3718 ( .A(n3487), .B(n3488), .Z(n3490) );
  XOR U3719 ( .A(n3489), .B(n3490), .Z(n3341) );
  NANDN U3720 ( .A(n3315), .B(n3314), .Z(n3319) );
  NANDN U3721 ( .A(n3317), .B(n3316), .Z(n3318) );
  AND U3722 ( .A(n3319), .B(n3318), .Z(n3339) );
  NAND U3723 ( .A(n3321), .B(n3320), .Z(n3325) );
  NAND U3724 ( .A(n3323), .B(n3322), .Z(n3324) );
  AND U3725 ( .A(n3325), .B(n3324), .Z(n3338) );
  XNOR U3726 ( .A(n3339), .B(n3338), .Z(n3340) );
  XNOR U3727 ( .A(n3341), .B(n3340), .Z(n3493) );
  XNOR U3728 ( .A(n3494), .B(n3493), .Z(n3495) );
  XOR U3729 ( .A(n3496), .B(n3495), .Z(n3333) );
  NANDN U3730 ( .A(n3327), .B(n3326), .Z(n3331) );
  OR U3731 ( .A(n3329), .B(n3328), .Z(n3330) );
  AND U3732 ( .A(n3331), .B(n3330), .Z(n3332) );
  XNOR U3733 ( .A(n3333), .B(n3332), .Z(n3334) );
  XNOR U3734 ( .A(n3335), .B(n3334), .Z(n3500) );
  XNOR U3735 ( .A(n3501), .B(n3500), .Z(c[100]) );
  NANDN U3736 ( .A(n3333), .B(n3332), .Z(n3337) );
  NANDN U3737 ( .A(n3335), .B(n3334), .Z(n3336) );
  AND U3738 ( .A(n3337), .B(n3336), .Z(n3512) );
  NANDN U3739 ( .A(n3339), .B(n3338), .Z(n3343) );
  NANDN U3740 ( .A(n3341), .B(n3340), .Z(n3342) );
  AND U3741 ( .A(n3343), .B(n3342), .Z(n3673) );
  NANDN U3742 ( .A(n3345), .B(n3344), .Z(n3349) );
  NANDN U3743 ( .A(n3347), .B(n3346), .Z(n3348) );
  AND U3744 ( .A(n3349), .B(n3348), .Z(n3666) );
  NANDN U3745 ( .A(n3351), .B(n3350), .Z(n3355) );
  NANDN U3746 ( .A(n3353), .B(n3352), .Z(n3354) );
  NAND U3747 ( .A(n3355), .B(n3354), .Z(n3665) );
  XNOR U3748 ( .A(n3666), .B(n3665), .Z(n3668) );
  NANDN U3749 ( .A(n3357), .B(n3356), .Z(n3361) );
  NAND U3750 ( .A(n3359), .B(n3358), .Z(n3360) );
  AND U3751 ( .A(n3361), .B(n3360), .Z(n3598) );
  NANDN U3752 ( .A(n3363), .B(n3362), .Z(n3367) );
  NANDN U3753 ( .A(n3365), .B(n3364), .Z(n3366) );
  AND U3754 ( .A(n3367), .B(n3366), .Z(n3597) );
  NANDN U3755 ( .A(n3369), .B(n3368), .Z(n3373) );
  OR U3756 ( .A(n3371), .B(n3370), .Z(n3372) );
  NAND U3757 ( .A(n3373), .B(n3372), .Z(n3596) );
  XOR U3758 ( .A(n3597), .B(n3596), .Z(n3599) );
  XOR U3759 ( .A(n3598), .B(n3599), .Z(n3592) );
  NANDN U3760 ( .A(n34634), .B(n3374), .Z(n3376) );
  XOR U3761 ( .A(b[29]), .B(a[9]), .Z(n3557) );
  NANDN U3762 ( .A(n34722), .B(n3557), .Z(n3375) );
  AND U3763 ( .A(n3376), .B(n3375), .Z(n3637) );
  NANDN U3764 ( .A(n34909), .B(n3377), .Z(n3379) );
  XOR U3765 ( .A(b[31]), .B(a[7]), .Z(n3614) );
  NANDN U3766 ( .A(n35145), .B(n3614), .Z(n3378) );
  AND U3767 ( .A(n3379), .B(n3378), .Z(n3636) );
  NANDN U3768 ( .A(n30482), .B(n3380), .Z(n3382) );
  XOR U3769 ( .A(b[11]), .B(a[27]), .Z(n3545) );
  NANDN U3770 ( .A(n30891), .B(n3545), .Z(n3381) );
  NAND U3771 ( .A(n3382), .B(n3381), .Z(n3635) );
  XOR U3772 ( .A(n3636), .B(n3635), .Z(n3638) );
  XOR U3773 ( .A(n3637), .B(n3638), .Z(n3632) );
  NANDN U3774 ( .A(n3383), .B(n33413), .Z(n3385) );
  XOR U3775 ( .A(b[21]), .B(a[17]), .Z(n3647) );
  NANDN U3776 ( .A(n33271), .B(n3647), .Z(n3384) );
  AND U3777 ( .A(n3385), .B(n3384), .Z(n3529) );
  NANDN U3778 ( .A(n33875), .B(n3386), .Z(n3388) );
  XOR U3779 ( .A(b[25]), .B(a[13]), .Z(n3548) );
  NANDN U3780 ( .A(n33994), .B(n3548), .Z(n3387) );
  AND U3781 ( .A(n3388), .B(n3387), .Z(n3528) );
  NANDN U3782 ( .A(n31055), .B(n3389), .Z(n3391) );
  XOR U3783 ( .A(b[13]), .B(a[25]), .Z(n3542) );
  NANDN U3784 ( .A(n31293), .B(n3542), .Z(n3390) );
  NAND U3785 ( .A(n3391), .B(n3390), .Z(n3527) );
  XOR U3786 ( .A(n3528), .B(n3527), .Z(n3530) );
  XOR U3787 ( .A(n3529), .B(n3530), .Z(n3630) );
  NAND U3788 ( .A(n32023), .B(n3392), .Z(n3394) );
  XNOR U3789 ( .A(b[15]), .B(a[23]), .Z(n3650) );
  NANDN U3790 ( .A(n3650), .B(n32024), .Z(n3393) );
  AND U3791 ( .A(n3394), .B(n3393), .Z(n3629) );
  XNOR U3792 ( .A(n3630), .B(n3629), .Z(n3631) );
  XNOR U3793 ( .A(n3632), .B(n3631), .Z(n3590) );
  NANDN U3794 ( .A(n210), .B(n3395), .Z(n3397) );
  XOR U3795 ( .A(b[9]), .B(a[29]), .Z(n3539) );
  NANDN U3796 ( .A(n30267), .B(n3539), .Z(n3396) );
  AND U3797 ( .A(n3397), .B(n3396), .Z(n3568) );
  NANDN U3798 ( .A(n35260), .B(n3398), .Z(n3400) );
  XOR U3799 ( .A(b[33]), .B(a[5]), .Z(n3617) );
  NANDN U3800 ( .A(n35456), .B(n3617), .Z(n3399) );
  AND U3801 ( .A(n3400), .B(n3399), .Z(n3567) );
  NANDN U3802 ( .A(n34223), .B(n3401), .Z(n3403) );
  XOR U3803 ( .A(b[27]), .B(a[11]), .Z(n3551) );
  NANDN U3804 ( .A(n34458), .B(n3551), .Z(n3402) );
  NAND U3805 ( .A(n3403), .B(n3402), .Z(n3566) );
  XOR U3806 ( .A(n3567), .B(n3566), .Z(n3569) );
  XOR U3807 ( .A(n3568), .B(n3569), .Z(n3579) );
  NANDN U3808 ( .A(n3404), .B(n9942), .Z(n3406) );
  XOR U3809 ( .A(b[3]), .B(a[35]), .Z(n3560) );
  NANDN U3810 ( .A(n28941), .B(n3560), .Z(n3405) );
  AND U3811 ( .A(n3406), .B(n3405), .Z(n3574) );
  NANDN U3812 ( .A(n32013), .B(n3407), .Z(n3409) );
  XOR U3813 ( .A(b[17]), .B(a[21]), .Z(n3563) );
  NANDN U3814 ( .A(n32292), .B(n3563), .Z(n3408) );
  NAND U3815 ( .A(n3409), .B(n3408), .Z(n3572) );
  NAND U3816 ( .A(b[0]), .B(a[37]), .Z(n3410) );
  XNOR U3817 ( .A(b[1]), .B(n3410), .Z(n3412) );
  NANDN U3818 ( .A(b[0]), .B(a[36]), .Z(n3411) );
  NAND U3819 ( .A(n3412), .B(n3411), .Z(n3573) );
  XOR U3820 ( .A(n3572), .B(n3573), .Z(n3575) );
  XNOR U3821 ( .A(n3574), .B(n3575), .Z(n3578) );
  XNOR U3822 ( .A(n3579), .B(n3578), .Z(n3580) );
  NANDN U3823 ( .A(n3414), .B(n3413), .Z(n3418) );
  OR U3824 ( .A(n3416), .B(n3415), .Z(n3417) );
  NAND U3825 ( .A(n3418), .B(n3417), .Z(n3581) );
  XOR U3826 ( .A(n3580), .B(n3581), .Z(n3591) );
  XOR U3827 ( .A(n3590), .B(n3591), .Z(n3593) );
  XOR U3828 ( .A(n3592), .B(n3593), .Z(n3517) );
  NANDN U3829 ( .A(n3420), .B(n3419), .Z(n3424) );
  NANDN U3830 ( .A(n3422), .B(n3421), .Z(n3423) );
  AND U3831 ( .A(n3424), .B(n3423), .Z(n3516) );
  NAND U3832 ( .A(n3426), .B(n3425), .Z(n3430) );
  NAND U3833 ( .A(n3428), .B(n3427), .Z(n3429) );
  NAND U3834 ( .A(n3430), .B(n3429), .Z(n3515) );
  XOR U3835 ( .A(n3516), .B(n3515), .Z(n3518) );
  XOR U3836 ( .A(n3517), .B(n3518), .Z(n3660) );
  NANDN U3837 ( .A(n3432), .B(n3431), .Z(n3436) );
  OR U3838 ( .A(n3434), .B(n3433), .Z(n3435) );
  AND U3839 ( .A(n3436), .B(n3435), .Z(n3659) );
  XNOR U3840 ( .A(n3660), .B(n3659), .Z(n3661) );
  NANDN U3841 ( .A(n3438), .B(n3437), .Z(n3442) );
  OR U3842 ( .A(n3440), .B(n3439), .Z(n3441) );
  AND U3843 ( .A(n3442), .B(n3441), .Z(n3524) );
  NANDN U3844 ( .A(n3443), .B(n3456), .Z(n3447) );
  NANDN U3845 ( .A(n3445), .B(n3444), .Z(n3446) );
  AND U3846 ( .A(n3447), .B(n3446), .Z(n3586) );
  NANDN U3847 ( .A(n35611), .B(n3448), .Z(n3450) );
  XOR U3848 ( .A(b[35]), .B(a[3]), .Z(n3536) );
  NANDN U3849 ( .A(n35801), .B(n3536), .Z(n3449) );
  AND U3850 ( .A(n3450), .B(n3449), .Z(n3641) );
  XOR U3851 ( .A(b[37]), .B(b[36]), .Z(n3643) );
  XOR U3852 ( .A(b[37]), .B(a[0]), .Z(n3451) );
  NAND U3853 ( .A(n3643), .B(n3451), .Z(n3452) );
  OR U3854 ( .A(n3452), .B(n36239), .Z(n3454) );
  XOR U3855 ( .A(b[37]), .B(a[1]), .Z(n3644) );
  NAND U3856 ( .A(n36239), .B(n3644), .Z(n3453) );
  AND U3857 ( .A(n3454), .B(n3453), .Z(n3642) );
  XOR U3858 ( .A(n3641), .B(n3642), .Z(n3610) );
  NAND U3859 ( .A(b[35]), .B(b[36]), .Z(n3455) );
  NAND U3860 ( .A(b[37]), .B(n3455), .Z(n36327) );
  NOR U3861 ( .A(n36327), .B(n3456), .Z(n3609) );
  NAND U3862 ( .A(n33000), .B(n3457), .Z(n3459) );
  XNOR U3863 ( .A(b[19]), .B(a[19]), .Z(n3620) );
  NANDN U3864 ( .A(n3620), .B(n33001), .Z(n3458) );
  AND U3865 ( .A(n3459), .B(n3458), .Z(n3608) );
  XOR U3866 ( .A(n3609), .B(n3608), .Z(n3611) );
  XOR U3867 ( .A(n3610), .B(n3611), .Z(n3585) );
  NANDN U3868 ( .A(n29499), .B(n3460), .Z(n3462) );
  XOR U3869 ( .A(b[7]), .B(a[31]), .Z(n3656) );
  NANDN U3870 ( .A(n29735), .B(n3656), .Z(n3461) );
  AND U3871 ( .A(n3462), .B(n3461), .Z(n3626) );
  NANDN U3872 ( .A(n28889), .B(n3463), .Z(n3465) );
  XOR U3873 ( .A(b[5]), .B(a[33]), .Z(n3554) );
  NANDN U3874 ( .A(n29138), .B(n3554), .Z(n3464) );
  AND U3875 ( .A(n3465), .B(n3464), .Z(n3624) );
  NANDN U3876 ( .A(n33866), .B(n3466), .Z(n3468) );
  XOR U3877 ( .A(b[23]), .B(a[15]), .Z(n3653) );
  NANDN U3878 ( .A(n33644), .B(n3653), .Z(n3467) );
  NAND U3879 ( .A(n3468), .B(n3467), .Z(n3623) );
  XNOR U3880 ( .A(n3624), .B(n3623), .Z(n3625) );
  XNOR U3881 ( .A(n3626), .B(n3625), .Z(n3584) );
  XOR U3882 ( .A(n3585), .B(n3584), .Z(n3587) );
  XOR U3883 ( .A(n3586), .B(n3587), .Z(n3605) );
  NANDN U3884 ( .A(n3470), .B(n3469), .Z(n3474) );
  OR U3885 ( .A(n3472), .B(n3471), .Z(n3473) );
  AND U3886 ( .A(n3474), .B(n3473), .Z(n3603) );
  NANDN U3887 ( .A(n3476), .B(n3475), .Z(n3480) );
  NANDN U3888 ( .A(n3478), .B(n3477), .Z(n3479) );
  AND U3889 ( .A(n3480), .B(n3479), .Z(n3602) );
  XNOR U3890 ( .A(n3603), .B(n3602), .Z(n3604) );
  XNOR U3891 ( .A(n3605), .B(n3604), .Z(n3521) );
  NANDN U3892 ( .A(n3482), .B(n3481), .Z(n3486) );
  NAND U3893 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U3894 ( .A(n3486), .B(n3485), .Z(n3522) );
  XNOR U3895 ( .A(n3521), .B(n3522), .Z(n3523) );
  XOR U3896 ( .A(n3524), .B(n3523), .Z(n3662) );
  XNOR U3897 ( .A(n3661), .B(n3662), .Z(n3667) );
  XOR U3898 ( .A(n3668), .B(n3667), .Z(n3672) );
  NANDN U3899 ( .A(n3488), .B(n3487), .Z(n3492) );
  OR U3900 ( .A(n3490), .B(n3489), .Z(n3491) );
  AND U3901 ( .A(n3492), .B(n3491), .Z(n3671) );
  XOR U3902 ( .A(n3672), .B(n3671), .Z(n3674) );
  XOR U3903 ( .A(n3673), .B(n3674), .Z(n3510) );
  NANDN U3904 ( .A(n3494), .B(n3493), .Z(n3498) );
  NAND U3905 ( .A(n3496), .B(n3495), .Z(n3497) );
  AND U3906 ( .A(n3498), .B(n3497), .Z(n3509) );
  XNOR U3907 ( .A(n3510), .B(n3509), .Z(n3511) );
  XNOR U3908 ( .A(n3512), .B(n3511), .Z(n3504) );
  XNOR U3909 ( .A(sreg[101]), .B(n3504), .Z(n3506) );
  OR U3910 ( .A(sreg[100]), .B(n3499), .Z(n3503) );
  NAND U3911 ( .A(n3501), .B(n3500), .Z(n3502) );
  NAND U3912 ( .A(n3503), .B(n3502), .Z(n3505) );
  XNOR U3913 ( .A(n3506), .B(n3505), .Z(c[101]) );
  NANDN U3914 ( .A(sreg[101]), .B(n3504), .Z(n3508) );
  NAND U3915 ( .A(n3506), .B(n3505), .Z(n3507) );
  AND U3916 ( .A(n3508), .B(n3507), .Z(n3678) );
  NANDN U3917 ( .A(n3510), .B(n3509), .Z(n3514) );
  NANDN U3918 ( .A(n3512), .B(n3511), .Z(n3513) );
  AND U3919 ( .A(n3514), .B(n3513), .Z(n3683) );
  NANDN U3920 ( .A(n3516), .B(n3515), .Z(n3520) );
  OR U3921 ( .A(n3518), .B(n3517), .Z(n3519) );
  AND U3922 ( .A(n3520), .B(n3519), .Z(n3851) );
  NANDN U3923 ( .A(n3522), .B(n3521), .Z(n3526) );
  NANDN U3924 ( .A(n3524), .B(n3523), .Z(n3525) );
  AND U3925 ( .A(n3526), .B(n3525), .Z(n3850) );
  XNOR U3926 ( .A(n3851), .B(n3850), .Z(n3853) );
  NANDN U3927 ( .A(n3528), .B(n3527), .Z(n3532) );
  OR U3928 ( .A(n3530), .B(n3529), .Z(n3531) );
  AND U3929 ( .A(n3532), .B(n3531), .Z(n3828) );
  NAND U3930 ( .A(b[0]), .B(a[38]), .Z(n3533) );
  XNOR U3931 ( .A(b[1]), .B(n3533), .Z(n3535) );
  NANDN U3932 ( .A(b[0]), .B(a[37]), .Z(n3534) );
  NAND U3933 ( .A(n3535), .B(n3534), .Z(n3823) );
  XOR U3934 ( .A(b[38]), .B(b[37]), .Z(n36491) );
  IV U3935 ( .A(n36491), .Z(n36347) );
  ANDN U3936 ( .B(a[0]), .A(n36347), .Z(n3820) );
  NANDN U3937 ( .A(n35611), .B(n3536), .Z(n3538) );
  XOR U3938 ( .A(b[35]), .B(a[4]), .Z(n3740) );
  NANDN U3939 ( .A(n35801), .B(n3740), .Z(n3537) );
  AND U3940 ( .A(n3538), .B(n3537), .Z(n3821) );
  XNOR U3941 ( .A(n3820), .B(n3821), .Z(n3822) );
  XNOR U3942 ( .A(n3823), .B(n3822), .Z(n3826) );
  NANDN U3943 ( .A(n210), .B(n3539), .Z(n3541) );
  XOR U3944 ( .A(b[9]), .B(a[30]), .Z(n3810) );
  NANDN U3945 ( .A(n30267), .B(n3810), .Z(n3540) );
  AND U3946 ( .A(n3541), .B(n3540), .Z(n3795) );
  NANDN U3947 ( .A(n31055), .B(n3542), .Z(n3544) );
  XOR U3948 ( .A(b[13]), .B(a[26]), .Z(n3801) );
  NANDN U3949 ( .A(n31293), .B(n3801), .Z(n3543) );
  AND U3950 ( .A(n3544), .B(n3543), .Z(n3793) );
  NANDN U3951 ( .A(n30482), .B(n3545), .Z(n3547) );
  XOR U3952 ( .A(b[11]), .B(a[28]), .Z(n3804) );
  NANDN U3953 ( .A(n30891), .B(n3804), .Z(n3546) );
  NAND U3954 ( .A(n3547), .B(n3546), .Z(n3792) );
  XNOR U3955 ( .A(n3793), .B(n3792), .Z(n3794) );
  XOR U3956 ( .A(n3795), .B(n3794), .Z(n3827) );
  XOR U3957 ( .A(n3826), .B(n3827), .Z(n3829) );
  XOR U3958 ( .A(n3828), .B(n3829), .Z(n3701) );
  NANDN U3959 ( .A(n33875), .B(n3548), .Z(n3550) );
  XOR U3960 ( .A(b[25]), .B(a[14]), .Z(n3743) );
  NANDN U3961 ( .A(n33994), .B(n3743), .Z(n3549) );
  AND U3962 ( .A(n3550), .B(n3549), .Z(n3754) );
  NANDN U3963 ( .A(n34223), .B(n3551), .Z(n3553) );
  XOR U3964 ( .A(b[27]), .B(a[12]), .Z(n3777) );
  NANDN U3965 ( .A(n34458), .B(n3777), .Z(n3552) );
  AND U3966 ( .A(n3553), .B(n3552), .Z(n3753) );
  NANDN U3967 ( .A(n28889), .B(n3554), .Z(n3556) );
  XOR U3968 ( .A(b[5]), .B(a[34]), .Z(n3731) );
  NANDN U3969 ( .A(n29138), .B(n3731), .Z(n3555) );
  NAND U3970 ( .A(n3556), .B(n3555), .Z(n3752) );
  XOR U3971 ( .A(n3753), .B(n3752), .Z(n3755) );
  XOR U3972 ( .A(n3754), .B(n3755), .Z(n3839) );
  NANDN U3973 ( .A(n34634), .B(n3557), .Z(n3559) );
  XOR U3974 ( .A(b[29]), .B(a[10]), .Z(n3780) );
  NANDN U3975 ( .A(n34722), .B(n3780), .Z(n3558) );
  AND U3976 ( .A(n3559), .B(n3558), .Z(n3760) );
  NANDN U3977 ( .A(n209), .B(n3560), .Z(n3562) );
  XOR U3978 ( .A(b[3]), .B(a[36]), .Z(n3813) );
  NANDN U3979 ( .A(n28941), .B(n3813), .Z(n3561) );
  AND U3980 ( .A(n3562), .B(n3561), .Z(n3759) );
  NANDN U3981 ( .A(n32013), .B(n3563), .Z(n3565) );
  XOR U3982 ( .A(b[17]), .B(a[22]), .Z(n3734) );
  NANDN U3983 ( .A(n32292), .B(n3734), .Z(n3564) );
  NAND U3984 ( .A(n3565), .B(n3564), .Z(n3758) );
  XOR U3985 ( .A(n3759), .B(n3758), .Z(n3761) );
  XNOR U3986 ( .A(n3760), .B(n3761), .Z(n3838) );
  XNOR U3987 ( .A(n3839), .B(n3838), .Z(n3840) );
  NANDN U3988 ( .A(n3567), .B(n3566), .Z(n3571) );
  OR U3989 ( .A(n3569), .B(n3568), .Z(n3570) );
  NAND U3990 ( .A(n3571), .B(n3570), .Z(n3841) );
  XNOR U3991 ( .A(n3840), .B(n3841), .Z(n3698) );
  NANDN U3992 ( .A(n3573), .B(n3572), .Z(n3577) );
  OR U3993 ( .A(n3575), .B(n3574), .Z(n3576) );
  NAND U3994 ( .A(n3577), .B(n3576), .Z(n3699) );
  XNOR U3995 ( .A(n3698), .B(n3699), .Z(n3700) );
  XNOR U3996 ( .A(n3701), .B(n3700), .Z(n3695) );
  NANDN U3997 ( .A(n3579), .B(n3578), .Z(n3583) );
  NANDN U3998 ( .A(n3581), .B(n3580), .Z(n3582) );
  AND U3999 ( .A(n3583), .B(n3582), .Z(n3693) );
  NANDN U4000 ( .A(n3585), .B(n3584), .Z(n3589) );
  OR U4001 ( .A(n3587), .B(n3586), .Z(n3588) );
  AND U4002 ( .A(n3589), .B(n3588), .Z(n3692) );
  XNOR U4003 ( .A(n3693), .B(n3692), .Z(n3694) );
  XOR U4004 ( .A(n3695), .B(n3694), .Z(n3845) );
  NANDN U4005 ( .A(n3591), .B(n3590), .Z(n3595) );
  OR U4006 ( .A(n3593), .B(n3592), .Z(n3594) );
  AND U4007 ( .A(n3595), .B(n3594), .Z(n3844) );
  XNOR U4008 ( .A(n3845), .B(n3844), .Z(n3846) );
  NANDN U4009 ( .A(n3597), .B(n3596), .Z(n3601) );
  OR U4010 ( .A(n3599), .B(n3598), .Z(n3600) );
  AND U4011 ( .A(n3601), .B(n3600), .Z(n3711) );
  NANDN U4012 ( .A(n3603), .B(n3602), .Z(n3607) );
  NANDN U4013 ( .A(n3605), .B(n3604), .Z(n3606) );
  AND U4014 ( .A(n3607), .B(n3606), .Z(n3710) );
  XNOR U4015 ( .A(n3711), .B(n3710), .Z(n3712) );
  NANDN U4016 ( .A(n3609), .B(n3608), .Z(n3613) );
  OR U4017 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U4018 ( .A(n3613), .B(n3612), .Z(n3717) );
  NANDN U4019 ( .A(n34909), .B(n3614), .Z(n3616) );
  XOR U4020 ( .A(b[31]), .B(a[8]), .Z(n3728) );
  NANDN U4021 ( .A(n35145), .B(n3728), .Z(n3615) );
  AND U4022 ( .A(n3616), .B(n3615), .Z(n3748) );
  NANDN U4023 ( .A(n35260), .B(n3617), .Z(n3619) );
  XOR U4024 ( .A(b[33]), .B(a[6]), .Z(n3737) );
  NANDN U4025 ( .A(n35456), .B(n3737), .Z(n3618) );
  AND U4026 ( .A(n3619), .B(n3618), .Z(n3747) );
  NANDN U4027 ( .A(n3620), .B(n33000), .Z(n3622) );
  XOR U4028 ( .A(b[19]), .B(a[20]), .Z(n3807) );
  NANDN U4029 ( .A(n32823), .B(n3807), .Z(n3621) );
  NAND U4030 ( .A(n3622), .B(n3621), .Z(n3746) );
  XOR U4031 ( .A(n3747), .B(n3746), .Z(n3749) );
  XNOR U4032 ( .A(n3748), .B(n3749), .Z(n3716) );
  XNOR U4033 ( .A(n3717), .B(n3716), .Z(n3719) );
  NANDN U4034 ( .A(n3624), .B(n3623), .Z(n3628) );
  NANDN U4035 ( .A(n3626), .B(n3625), .Z(n3627) );
  AND U4036 ( .A(n3628), .B(n3627), .Z(n3718) );
  XOR U4037 ( .A(n3719), .B(n3718), .Z(n3707) );
  NANDN U4038 ( .A(n3630), .B(n3629), .Z(n3634) );
  NANDN U4039 ( .A(n3632), .B(n3631), .Z(n3633) );
  AND U4040 ( .A(n3634), .B(n3633), .Z(n3704) );
  NANDN U4041 ( .A(n3636), .B(n3635), .Z(n3640) );
  OR U4042 ( .A(n3638), .B(n3637), .Z(n3639) );
  AND U4043 ( .A(n3640), .B(n3639), .Z(n3835) );
  NOR U4044 ( .A(n3642), .B(n3641), .Z(n3788) );
  ANDN U4045 ( .B(n3643), .A(n36239), .Z(n36238) );
  NAND U4046 ( .A(n36238), .B(n3644), .Z(n3646) );
  XNOR U4047 ( .A(b[37]), .B(a[2]), .Z(n3768) );
  NANDN U4048 ( .A(n3768), .B(n36239), .Z(n3645) );
  AND U4049 ( .A(n3646), .B(n3645), .Z(n3786) );
  NAND U4050 ( .A(n33413), .B(n3647), .Z(n3649) );
  XNOR U4051 ( .A(b[21]), .B(a[18]), .Z(n3774) );
  NANDN U4052 ( .A(n3774), .B(n33414), .Z(n3648) );
  NAND U4053 ( .A(n3649), .B(n3648), .Z(n3787) );
  XOR U4054 ( .A(n3786), .B(n3787), .Z(n3789) );
  XOR U4055 ( .A(n3788), .B(n3789), .Z(n3833) );
  NANDN U4056 ( .A(n3650), .B(n32023), .Z(n3652) );
  XOR U4057 ( .A(b[15]), .B(a[24]), .Z(n3798) );
  NANDN U4058 ( .A(n31925), .B(n3798), .Z(n3651) );
  AND U4059 ( .A(n3652), .B(n3651), .Z(n3725) );
  NANDN U4060 ( .A(n33866), .B(n3653), .Z(n3655) );
  XOR U4061 ( .A(b[23]), .B(a[16]), .Z(n3816) );
  NANDN U4062 ( .A(n33644), .B(n3816), .Z(n3654) );
  AND U4063 ( .A(n3655), .B(n3654), .Z(n3723) );
  NANDN U4064 ( .A(n29499), .B(n3656), .Z(n3658) );
  XOR U4065 ( .A(b[7]), .B(a[32]), .Z(n3783) );
  NANDN U4066 ( .A(n29735), .B(n3783), .Z(n3657) );
  NAND U4067 ( .A(n3658), .B(n3657), .Z(n3722) );
  XNOR U4068 ( .A(n3723), .B(n3722), .Z(n3724) );
  XNOR U4069 ( .A(n3725), .B(n3724), .Z(n3832) );
  XNOR U4070 ( .A(n3833), .B(n3832), .Z(n3834) );
  XOR U4071 ( .A(n3835), .B(n3834), .Z(n3705) );
  XNOR U4072 ( .A(n3704), .B(n3705), .Z(n3706) );
  XOR U4073 ( .A(n3707), .B(n3706), .Z(n3713) );
  XOR U4074 ( .A(n3712), .B(n3713), .Z(n3847) );
  XNOR U4075 ( .A(n3846), .B(n3847), .Z(n3852) );
  XOR U4076 ( .A(n3853), .B(n3852), .Z(n3689) );
  NANDN U4077 ( .A(n3660), .B(n3659), .Z(n3664) );
  NANDN U4078 ( .A(n3662), .B(n3661), .Z(n3663) );
  AND U4079 ( .A(n3664), .B(n3663), .Z(n3687) );
  NANDN U4080 ( .A(n3666), .B(n3665), .Z(n3670) );
  NAND U4081 ( .A(n3668), .B(n3667), .Z(n3669) );
  NAND U4082 ( .A(n3670), .B(n3669), .Z(n3686) );
  XNOR U4083 ( .A(n3687), .B(n3686), .Z(n3688) );
  XNOR U4084 ( .A(n3689), .B(n3688), .Z(n3680) );
  NANDN U4085 ( .A(n3672), .B(n3671), .Z(n3676) );
  OR U4086 ( .A(n3674), .B(n3673), .Z(n3675) );
  NAND U4087 ( .A(n3676), .B(n3675), .Z(n3681) );
  XNOR U4088 ( .A(n3680), .B(n3681), .Z(n3682) );
  XNOR U4089 ( .A(n3683), .B(n3682), .Z(n3679) );
  XNOR U4090 ( .A(sreg[102]), .B(n3679), .Z(n3677) );
  XOR U4091 ( .A(n3678), .B(n3677), .Z(c[102]) );
  NANDN U4092 ( .A(n3681), .B(n3680), .Z(n3685) );
  NANDN U4093 ( .A(n3683), .B(n3682), .Z(n3684) );
  AND U4094 ( .A(n3685), .B(n3684), .Z(n3859) );
  NANDN U4095 ( .A(n3687), .B(n3686), .Z(n3691) );
  NANDN U4096 ( .A(n3689), .B(n3688), .Z(n3690) );
  AND U4097 ( .A(n3691), .B(n3690), .Z(n3857) );
  NANDN U4098 ( .A(n3693), .B(n3692), .Z(n3697) );
  NAND U4099 ( .A(n3695), .B(n3694), .Z(n3696) );
  AND U4100 ( .A(n3697), .B(n3696), .Z(n3870) );
  NANDN U4101 ( .A(n3699), .B(n3698), .Z(n3703) );
  NANDN U4102 ( .A(n3701), .B(n3700), .Z(n3702) );
  AND U4103 ( .A(n3703), .B(n3702), .Z(n3869) );
  NANDN U4104 ( .A(n3705), .B(n3704), .Z(n3709) );
  NANDN U4105 ( .A(n3707), .B(n3706), .Z(n3708) );
  AND U4106 ( .A(n3709), .B(n3708), .Z(n3868) );
  XOR U4107 ( .A(n3869), .B(n3868), .Z(n3871) );
  XOR U4108 ( .A(n3870), .B(n3871), .Z(n3864) );
  NANDN U4109 ( .A(n3711), .B(n3710), .Z(n3715) );
  NANDN U4110 ( .A(n3713), .B(n3712), .Z(n3714) );
  AND U4111 ( .A(n3715), .B(n3714), .Z(n3863) );
  NANDN U4112 ( .A(n3717), .B(n3716), .Z(n3721) );
  NAND U4113 ( .A(n3719), .B(n3718), .Z(n3720) );
  AND U4114 ( .A(n3721), .B(n3720), .Z(n3882) );
  NANDN U4115 ( .A(n3723), .B(n3722), .Z(n3727) );
  NANDN U4116 ( .A(n3725), .B(n3724), .Z(n3726) );
  AND U4117 ( .A(n3727), .B(n3726), .Z(n3895) );
  NANDN U4118 ( .A(n34909), .B(n3728), .Z(n3730) );
  XOR U4119 ( .A(b[31]), .B(a[9]), .Z(n3999) );
  NANDN U4120 ( .A(n35145), .B(n3999), .Z(n3729) );
  AND U4121 ( .A(n3730), .B(n3729), .Z(n4018) );
  NANDN U4122 ( .A(n28889), .B(n3731), .Z(n3733) );
  XOR U4123 ( .A(b[5]), .B(a[35]), .Z(n4009) );
  NANDN U4124 ( .A(n29138), .B(n4009), .Z(n3732) );
  AND U4125 ( .A(n3733), .B(n3732), .Z(n4016) );
  NANDN U4126 ( .A(n32013), .B(n3734), .Z(n3736) );
  XOR U4127 ( .A(b[17]), .B(a[23]), .Z(n3972) );
  NANDN U4128 ( .A(n32292), .B(n3972), .Z(n3735) );
  NAND U4129 ( .A(n3736), .B(n3735), .Z(n4015) );
  XNOR U4130 ( .A(n4016), .B(n4015), .Z(n4017) );
  XOR U4131 ( .A(n4018), .B(n4017), .Z(n3893) );
  NANDN U4132 ( .A(n35260), .B(n3737), .Z(n3739) );
  XOR U4133 ( .A(b[33]), .B(a[7]), .Z(n4002) );
  NANDN U4134 ( .A(n35456), .B(n4002), .Z(n3738) );
  AND U4135 ( .A(n3739), .B(n3738), .Z(n3986) );
  NANDN U4136 ( .A(n35611), .B(n3740), .Z(n3742) );
  XOR U4137 ( .A(b[35]), .B(a[5]), .Z(n3951) );
  NANDN U4138 ( .A(n35801), .B(n3951), .Z(n3741) );
  AND U4139 ( .A(n3742), .B(n3741), .Z(n3985) );
  NANDN U4140 ( .A(n33875), .B(n3743), .Z(n3745) );
  XOR U4141 ( .A(b[25]), .B(a[15]), .Z(n4012) );
  NANDN U4142 ( .A(n33994), .B(n4012), .Z(n3744) );
  NAND U4143 ( .A(n3745), .B(n3744), .Z(n3984) );
  XOR U4144 ( .A(n3985), .B(n3984), .Z(n3987) );
  XNOR U4145 ( .A(n3986), .B(n3987), .Z(n3892) );
  XOR U4146 ( .A(n3893), .B(n3892), .Z(n3894) );
  XOR U4147 ( .A(n3895), .B(n3894), .Z(n3932) );
  NANDN U4148 ( .A(n3747), .B(n3746), .Z(n3751) );
  OR U4149 ( .A(n3749), .B(n3748), .Z(n3750) );
  AND U4150 ( .A(n3751), .B(n3750), .Z(n3931) );
  NANDN U4151 ( .A(n3753), .B(n3752), .Z(n3757) );
  OR U4152 ( .A(n3755), .B(n3754), .Z(n3756) );
  NAND U4153 ( .A(n3757), .B(n3756), .Z(n3930) );
  XOR U4154 ( .A(n3931), .B(n3930), .Z(n3933) );
  XOR U4155 ( .A(n3932), .B(n3933), .Z(n3881) );
  NANDN U4156 ( .A(n3759), .B(n3758), .Z(n3763) );
  OR U4157 ( .A(n3761), .B(n3760), .Z(n3762) );
  NAND U4158 ( .A(n3763), .B(n3762), .Z(n3900) );
  XOR U4159 ( .A(b[39]), .B(b[38]), .Z(n4005) );
  XOR U4160 ( .A(b[39]), .B(a[0]), .Z(n3764) );
  NAND U4161 ( .A(n4005), .B(n3764), .Z(n3765) );
  OR U4162 ( .A(n3765), .B(n36491), .Z(n3767) );
  XOR U4163 ( .A(b[39]), .B(a[1]), .Z(n4006) );
  NAND U4164 ( .A(n36491), .B(n4006), .Z(n3766) );
  AND U4165 ( .A(n3767), .B(n3766), .Z(n3923) );
  NANDN U4166 ( .A(n3768), .B(n36238), .Z(n3770) );
  XOR U4167 ( .A(b[37]), .B(a[3]), .Z(n3913) );
  NANDN U4168 ( .A(n36047), .B(n3913), .Z(n3769) );
  AND U4169 ( .A(n3770), .B(n3769), .Z(n3922) );
  XOR U4170 ( .A(n3923), .B(n3922), .Z(n3945) );
  NAND U4171 ( .A(b[0]), .B(a[39]), .Z(n3771) );
  XNOR U4172 ( .A(b[1]), .B(n3771), .Z(n3773) );
  NANDN U4173 ( .A(b[0]), .B(a[38]), .Z(n3772) );
  NAND U4174 ( .A(n3773), .B(n3772), .Z(n3942) );
  NANDN U4175 ( .A(n3774), .B(n33413), .Z(n3776) );
  XNOR U4176 ( .A(b[21]), .B(a[19]), .Z(n3954) );
  NANDN U4177 ( .A(n3954), .B(n33414), .Z(n3775) );
  NAND U4178 ( .A(n3776), .B(n3775), .Z(n3943) );
  XNOR U4179 ( .A(n3942), .B(n3943), .Z(n3944) );
  XOR U4180 ( .A(n3945), .B(n3944), .Z(n3898) );
  NANDN U4181 ( .A(n34223), .B(n3777), .Z(n3779) );
  XOR U4182 ( .A(b[27]), .B(a[13]), .Z(n3966) );
  NANDN U4183 ( .A(n34458), .B(n3966), .Z(n3778) );
  AND U4184 ( .A(n3779), .B(n3778), .Z(n3906) );
  NANDN U4185 ( .A(n34634), .B(n3780), .Z(n3782) );
  XOR U4186 ( .A(b[29]), .B(a[11]), .Z(n3996) );
  NANDN U4187 ( .A(n34722), .B(n3996), .Z(n3781) );
  AND U4188 ( .A(n3782), .B(n3781), .Z(n3905) );
  NANDN U4189 ( .A(n29499), .B(n3783), .Z(n3785) );
  XOR U4190 ( .A(b[7]), .B(a[33]), .Z(n3948) );
  NANDN U4191 ( .A(n29735), .B(n3948), .Z(n3784) );
  NAND U4192 ( .A(n3785), .B(n3784), .Z(n3904) );
  XOR U4193 ( .A(n3905), .B(n3904), .Z(n3907) );
  XOR U4194 ( .A(n3906), .B(n3907), .Z(n3899) );
  XNOR U4195 ( .A(n3898), .B(n3899), .Z(n3901) );
  NANDN U4196 ( .A(n3787), .B(n3786), .Z(n3791) );
  OR U4197 ( .A(n3789), .B(n3788), .Z(n3790) );
  AND U4198 ( .A(n3791), .B(n3790), .Z(n3925) );
  NANDN U4199 ( .A(n3793), .B(n3792), .Z(n3797) );
  NANDN U4200 ( .A(n3795), .B(n3794), .Z(n3796) );
  AND U4201 ( .A(n3797), .B(n3796), .Z(n3924) );
  XNOR U4202 ( .A(n3925), .B(n3924), .Z(n3926) );
  XOR U4203 ( .A(n3927), .B(n3926), .Z(n3880) );
  XOR U4204 ( .A(n3881), .B(n3880), .Z(n3883) );
  XOR U4205 ( .A(n3882), .B(n3883), .Z(n3877) );
  NANDN U4206 ( .A(n31536), .B(n3798), .Z(n3800) );
  XOR U4207 ( .A(b[15]), .B(a[25]), .Z(n3981) );
  NANDN U4208 ( .A(n31925), .B(n3981), .Z(n3799) );
  AND U4209 ( .A(n3800), .B(n3799), .Z(n4022) );
  NANDN U4210 ( .A(n31055), .B(n3801), .Z(n3803) );
  XOR U4211 ( .A(b[13]), .B(a[27]), .Z(n3975) );
  NANDN U4212 ( .A(n31293), .B(n3975), .Z(n3802) );
  NAND U4213 ( .A(n3803), .B(n3802), .Z(n4021) );
  XNOR U4214 ( .A(n4022), .B(n4021), .Z(n4024) );
  NANDN U4215 ( .A(n30482), .B(n3804), .Z(n3806) );
  XOR U4216 ( .A(b[11]), .B(a[29]), .Z(n3978) );
  NANDN U4217 ( .A(n30891), .B(n3978), .Z(n3805) );
  AND U4218 ( .A(n3806), .B(n3805), .Z(n3960) );
  NANDN U4219 ( .A(n32483), .B(n3807), .Z(n3809) );
  XOR U4220 ( .A(b[19]), .B(a[21]), .Z(n3963) );
  NANDN U4221 ( .A(n32823), .B(n3963), .Z(n3808) );
  AND U4222 ( .A(n3809), .B(n3808), .Z(n3958) );
  NANDN U4223 ( .A(n210), .B(n3810), .Z(n3812) );
  XOR U4224 ( .A(b[9]), .B(a[31]), .Z(n3969) );
  NANDN U4225 ( .A(n30267), .B(n3969), .Z(n3811) );
  NAND U4226 ( .A(n3812), .B(n3811), .Z(n3957) );
  XNOR U4227 ( .A(n3958), .B(n3957), .Z(n3959) );
  XNOR U4228 ( .A(n3960), .B(n3959), .Z(n4023) );
  XOR U4229 ( .A(n4024), .B(n4023), .Z(n3939) );
  NANDN U4230 ( .A(n209), .B(n3813), .Z(n3815) );
  XOR U4231 ( .A(b[3]), .B(a[37]), .Z(n3916) );
  NANDN U4232 ( .A(n28941), .B(n3916), .Z(n3814) );
  AND U4233 ( .A(n3815), .B(n3814), .Z(n3992) );
  NANDN U4234 ( .A(n33866), .B(n3816), .Z(n3818) );
  XOR U4235 ( .A(b[23]), .B(a[17]), .Z(n3919) );
  NANDN U4236 ( .A(n33644), .B(n3919), .Z(n3817) );
  AND U4237 ( .A(n3818), .B(n3817), .Z(n3991) );
  NAND U4238 ( .A(b[37]), .B(b[38]), .Z(n3819) );
  AND U4239 ( .A(b[39]), .B(n3819), .Z(n36728) );
  ANDN U4240 ( .B(n36728), .A(n3820), .Z(n3990) );
  XOR U4241 ( .A(n3991), .B(n3990), .Z(n3993) );
  XOR U4242 ( .A(n3992), .B(n3993), .Z(n3937) );
  NANDN U4243 ( .A(n3821), .B(n3820), .Z(n3825) );
  NANDN U4244 ( .A(n3823), .B(n3822), .Z(n3824) );
  AND U4245 ( .A(n3825), .B(n3824), .Z(n3936) );
  XNOR U4246 ( .A(n3937), .B(n3936), .Z(n3938) );
  XNOR U4247 ( .A(n3939), .B(n3938), .Z(n3886) );
  NANDN U4248 ( .A(n3827), .B(n3826), .Z(n3831) );
  OR U4249 ( .A(n3829), .B(n3828), .Z(n3830) );
  NAND U4250 ( .A(n3831), .B(n3830), .Z(n3887) );
  XNOR U4251 ( .A(n3886), .B(n3887), .Z(n3889) );
  NANDN U4252 ( .A(n3833), .B(n3832), .Z(n3837) );
  NANDN U4253 ( .A(n3835), .B(n3834), .Z(n3836) );
  AND U4254 ( .A(n3837), .B(n3836), .Z(n3888) );
  XOR U4255 ( .A(n3889), .B(n3888), .Z(n3875) );
  NANDN U4256 ( .A(n3839), .B(n3838), .Z(n3843) );
  NANDN U4257 ( .A(n3841), .B(n3840), .Z(n3842) );
  AND U4258 ( .A(n3843), .B(n3842), .Z(n3874) );
  XNOR U4259 ( .A(n3875), .B(n3874), .Z(n3876) );
  XNOR U4260 ( .A(n3877), .B(n3876), .Z(n3862) );
  XOR U4261 ( .A(n3863), .B(n3862), .Z(n3865) );
  XOR U4262 ( .A(n3864), .B(n3865), .Z(n4028) );
  NANDN U4263 ( .A(n3845), .B(n3844), .Z(n3849) );
  NANDN U4264 ( .A(n3847), .B(n3846), .Z(n3848) );
  AND U4265 ( .A(n3849), .B(n3848), .Z(n4027) );
  XNOR U4266 ( .A(n4028), .B(n4027), .Z(n4029) );
  NANDN U4267 ( .A(n3851), .B(n3850), .Z(n3855) );
  NAND U4268 ( .A(n3853), .B(n3852), .Z(n3854) );
  NAND U4269 ( .A(n3855), .B(n3854), .Z(n4030) );
  XNOR U4270 ( .A(n4029), .B(n4030), .Z(n3856) );
  XNOR U4271 ( .A(n3857), .B(n3856), .Z(n3858) );
  XNOR U4272 ( .A(n3859), .B(n3858), .Z(n4033) );
  XNOR U4273 ( .A(sreg[103]), .B(n4033), .Z(n4034) );
  XNOR U4274 ( .A(n4035), .B(n4034), .Z(c[103]) );
  NANDN U4275 ( .A(n3857), .B(n3856), .Z(n3861) );
  NANDN U4276 ( .A(n3859), .B(n3858), .Z(n3860) );
  AND U4277 ( .A(n3861), .B(n3860), .Z(n4041) );
  NANDN U4278 ( .A(n3863), .B(n3862), .Z(n3867) );
  OR U4279 ( .A(n3865), .B(n3864), .Z(n3866) );
  AND U4280 ( .A(n3867), .B(n3866), .Z(n4216) );
  NANDN U4281 ( .A(n3869), .B(n3868), .Z(n3873) );
  OR U4282 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U4283 ( .A(n3873), .B(n3872), .Z(n4215) );
  XNOR U4284 ( .A(n4216), .B(n4215), .Z(n4218) );
  NANDN U4285 ( .A(n3875), .B(n3874), .Z(n3879) );
  NANDN U4286 ( .A(n3877), .B(n3876), .Z(n3878) );
  AND U4287 ( .A(n3879), .B(n3878), .Z(n4210) );
  NANDN U4288 ( .A(n3881), .B(n3880), .Z(n3885) );
  OR U4289 ( .A(n3883), .B(n3882), .Z(n3884) );
  AND U4290 ( .A(n3885), .B(n3884), .Z(n4209) );
  XNOR U4291 ( .A(n4210), .B(n4209), .Z(n4211) );
  NANDN U4292 ( .A(n3887), .B(n3886), .Z(n3891) );
  NAND U4293 ( .A(n3889), .B(n3888), .Z(n3890) );
  AND U4294 ( .A(n3891), .B(n3890), .Z(n4205) );
  NAND U4295 ( .A(n3893), .B(n3892), .Z(n3897) );
  NAND U4296 ( .A(n3895), .B(n3894), .Z(n3896) );
  NAND U4297 ( .A(n3897), .B(n3896), .Z(n4047) );
  NAND U4298 ( .A(n3899), .B(n3898), .Z(n3903) );
  NANDN U4299 ( .A(n3901), .B(n3900), .Z(n3902) );
  AND U4300 ( .A(n3903), .B(n3902), .Z(n4046) );
  NANDN U4301 ( .A(n3905), .B(n3904), .Z(n3909) );
  OR U4302 ( .A(n3907), .B(n3906), .Z(n3908) );
  AND U4303 ( .A(n3909), .B(n3908), .Z(n4194) );
  NAND U4304 ( .A(b[0]), .B(a[40]), .Z(n3910) );
  XNOR U4305 ( .A(b[1]), .B(n3910), .Z(n3912) );
  NANDN U4306 ( .A(b[0]), .B(a[39]), .Z(n3911) );
  NAND U4307 ( .A(n3912), .B(n3911), .Z(n4068) );
  XOR U4308 ( .A(b[39]), .B(b[40]), .Z(n36733) );
  IV U4309 ( .A(n36733), .Z(n36594) );
  ANDN U4310 ( .B(a[0]), .A(n36594), .Z(n4169) );
  IV U4311 ( .A(n36238), .Z(n35936) );
  NANDN U4312 ( .A(n35936), .B(n3913), .Z(n3915) );
  XOR U4313 ( .A(b[37]), .B(a[4]), .Z(n4162) );
  NANDN U4314 ( .A(n36047), .B(n4162), .Z(n3914) );
  AND U4315 ( .A(n3915), .B(n3914), .Z(n4066) );
  XOR U4316 ( .A(n4169), .B(n4066), .Z(n4067) );
  XOR U4317 ( .A(n4068), .B(n4067), .Z(n4192) );
  NANDN U4318 ( .A(n209), .B(n3916), .Z(n3918) );
  XOR U4319 ( .A(b[3]), .B(a[38]), .Z(n4170) );
  NANDN U4320 ( .A(n28941), .B(n4170), .Z(n3917) );
  AND U4321 ( .A(n3918), .B(n3917), .Z(n4133) );
  NANDN U4322 ( .A(n33866), .B(n3919), .Z(n3921) );
  XOR U4323 ( .A(b[23]), .B(a[18]), .Z(n4165) );
  NANDN U4324 ( .A(n33644), .B(n4165), .Z(n3920) );
  NAND U4325 ( .A(n3921), .B(n3920), .Z(n4132) );
  XNOR U4326 ( .A(n4133), .B(n4132), .Z(n4135) );
  NOR U4327 ( .A(n3923), .B(n3922), .Z(n4134) );
  XNOR U4328 ( .A(n4135), .B(n4134), .Z(n4191) );
  XNOR U4329 ( .A(n4192), .B(n4191), .Z(n4193) );
  XOR U4330 ( .A(n4194), .B(n4193), .Z(n4045) );
  XOR U4331 ( .A(n4046), .B(n4045), .Z(n4048) );
  XOR U4332 ( .A(n4047), .B(n4048), .Z(n4092) );
  NANDN U4333 ( .A(n3925), .B(n3924), .Z(n3929) );
  NAND U4334 ( .A(n3927), .B(n3926), .Z(n3928) );
  AND U4335 ( .A(n3929), .B(n3928), .Z(n4090) );
  NANDN U4336 ( .A(n3931), .B(n3930), .Z(n3935) );
  OR U4337 ( .A(n3933), .B(n3932), .Z(n3934) );
  AND U4338 ( .A(n3935), .B(n3934), .Z(n4089) );
  XNOR U4339 ( .A(n4090), .B(n4089), .Z(n4091) );
  XOR U4340 ( .A(n4092), .B(n4091), .Z(n4204) );
  NANDN U4341 ( .A(n3937), .B(n3936), .Z(n3941) );
  NANDN U4342 ( .A(n3939), .B(n3938), .Z(n3940) );
  AND U4343 ( .A(n3941), .B(n3940), .Z(n4084) );
  NANDN U4344 ( .A(n3943), .B(n3942), .Z(n3947) );
  NANDN U4345 ( .A(n3945), .B(n3944), .Z(n3946) );
  AND U4346 ( .A(n3947), .B(n3946), .Z(n4186) );
  NANDN U4347 ( .A(n29499), .B(n3948), .Z(n3950) );
  XOR U4348 ( .A(b[7]), .B(a[34]), .Z(n4144) );
  NANDN U4349 ( .A(n29735), .B(n4144), .Z(n3949) );
  AND U4350 ( .A(n3950), .B(n3949), .Z(n4158) );
  NANDN U4351 ( .A(n35611), .B(n3951), .Z(n3953) );
  XOR U4352 ( .A(b[35]), .B(a[6]), .Z(n4173) );
  NANDN U4353 ( .A(n35801), .B(n4173), .Z(n3952) );
  AND U4354 ( .A(n3953), .B(n3952), .Z(n4157) );
  NANDN U4355 ( .A(n3954), .B(n33413), .Z(n3956) );
  XOR U4356 ( .A(b[21]), .B(a[20]), .Z(n4107) );
  NANDN U4357 ( .A(n33271), .B(n4107), .Z(n3955) );
  NAND U4358 ( .A(n3956), .B(n3955), .Z(n4156) );
  XOR U4359 ( .A(n4157), .B(n4156), .Z(n4159) );
  XNOR U4360 ( .A(n4158), .B(n4159), .Z(n4185) );
  XNOR U4361 ( .A(n4186), .B(n4185), .Z(n4187) );
  NANDN U4362 ( .A(n3958), .B(n3957), .Z(n3962) );
  NANDN U4363 ( .A(n3960), .B(n3959), .Z(n3961) );
  NAND U4364 ( .A(n3962), .B(n3961), .Z(n4188) );
  XNOR U4365 ( .A(n4187), .B(n4188), .Z(n4083) );
  XNOR U4366 ( .A(n4084), .B(n4083), .Z(n4086) );
  NANDN U4367 ( .A(n32483), .B(n3963), .Z(n3965) );
  XOR U4368 ( .A(b[19]), .B(a[22]), .Z(n4176) );
  NANDN U4369 ( .A(n32823), .B(n4176), .Z(n3964) );
  AND U4370 ( .A(n3965), .B(n3964), .Z(n4103) );
  NANDN U4371 ( .A(n34223), .B(n3966), .Z(n3968) );
  XOR U4372 ( .A(b[27]), .B(a[14]), .Z(n4141) );
  NANDN U4373 ( .A(n34458), .B(n4141), .Z(n3967) );
  AND U4374 ( .A(n3968), .B(n3967), .Z(n4102) );
  NANDN U4375 ( .A(n210), .B(n3969), .Z(n3971) );
  XOR U4376 ( .A(b[9]), .B(a[32]), .Z(n4117) );
  NANDN U4377 ( .A(n30267), .B(n4117), .Z(n3970) );
  NAND U4378 ( .A(n3971), .B(n3970), .Z(n4101) );
  XOR U4379 ( .A(n4102), .B(n4101), .Z(n4104) );
  XOR U4380 ( .A(n4103), .B(n4104), .Z(n4053) );
  NANDN U4381 ( .A(n32013), .B(n3972), .Z(n3974) );
  XOR U4382 ( .A(b[17]), .B(a[24]), .Z(n4138) );
  NANDN U4383 ( .A(n32292), .B(n4138), .Z(n3973) );
  AND U4384 ( .A(n3974), .B(n3973), .Z(n4073) );
  NANDN U4385 ( .A(n31055), .B(n3975), .Z(n3977) );
  XOR U4386 ( .A(b[13]), .B(a[28]), .Z(n4120) );
  NANDN U4387 ( .A(n31293), .B(n4120), .Z(n3976) );
  AND U4388 ( .A(n3977), .B(n3976), .Z(n4072) );
  NANDN U4389 ( .A(n30482), .B(n3978), .Z(n3980) );
  XOR U4390 ( .A(b[11]), .B(a[30]), .Z(n4123) );
  NANDN U4391 ( .A(n30891), .B(n4123), .Z(n3979) );
  NAND U4392 ( .A(n3980), .B(n3979), .Z(n4071) );
  XOR U4393 ( .A(n4072), .B(n4071), .Z(n4074) );
  XOR U4394 ( .A(n4073), .B(n4074), .Z(n4052) );
  NAND U4395 ( .A(n32023), .B(n3981), .Z(n3983) );
  XNOR U4396 ( .A(b[15]), .B(a[26]), .Z(n4063) );
  NANDN U4397 ( .A(n4063), .B(n32024), .Z(n3982) );
  AND U4398 ( .A(n3983), .B(n3982), .Z(n4051) );
  XOR U4399 ( .A(n4052), .B(n4051), .Z(n4054) );
  XOR U4400 ( .A(n4053), .B(n4054), .Z(n4079) );
  NANDN U4401 ( .A(n3985), .B(n3984), .Z(n3989) );
  OR U4402 ( .A(n3987), .B(n3986), .Z(n3988) );
  AND U4403 ( .A(n3989), .B(n3988), .Z(n4078) );
  NANDN U4404 ( .A(n3991), .B(n3990), .Z(n3995) );
  OR U4405 ( .A(n3993), .B(n3992), .Z(n3994) );
  NAND U4406 ( .A(n3995), .B(n3994), .Z(n4077) );
  XOR U4407 ( .A(n4078), .B(n4077), .Z(n4080) );
  XOR U4408 ( .A(n4079), .B(n4080), .Z(n4098) );
  NANDN U4409 ( .A(n34634), .B(n3996), .Z(n3998) );
  XOR U4410 ( .A(b[29]), .B(a[12]), .Z(n4057) );
  NANDN U4411 ( .A(n34722), .B(n4057), .Z(n3997) );
  AND U4412 ( .A(n3998), .B(n3997), .Z(n4181) );
  NANDN U4413 ( .A(n34909), .B(n3999), .Z(n4001) );
  XOR U4414 ( .A(b[31]), .B(a[10]), .Z(n4060) );
  NANDN U4415 ( .A(n35145), .B(n4060), .Z(n4000) );
  AND U4416 ( .A(n4001), .B(n4000), .Z(n4180) );
  NANDN U4417 ( .A(n35260), .B(n4002), .Z(n4004) );
  XOR U4418 ( .A(b[33]), .B(a[8]), .Z(n4147) );
  NANDN U4419 ( .A(n35456), .B(n4147), .Z(n4003) );
  NAND U4420 ( .A(n4004), .B(n4003), .Z(n4179) );
  XOR U4421 ( .A(n4180), .B(n4179), .Z(n4182) );
  XOR U4422 ( .A(n4181), .B(n4182), .Z(n4198) );
  ANDN U4423 ( .B(n4005), .A(n36491), .Z(n36490) );
  IV U4424 ( .A(n36490), .Z(n36210) );
  NANDN U4425 ( .A(n36210), .B(n4006), .Z(n4008) );
  XOR U4426 ( .A(b[39]), .B(a[2]), .Z(n4110) );
  NANDN U4427 ( .A(n36347), .B(n4110), .Z(n4007) );
  AND U4428 ( .A(n4008), .B(n4007), .Z(n4128) );
  NANDN U4429 ( .A(n28889), .B(n4009), .Z(n4011) );
  XOR U4430 ( .A(b[5]), .B(a[36]), .Z(n4150) );
  NANDN U4431 ( .A(n29138), .B(n4150), .Z(n4010) );
  AND U4432 ( .A(n4011), .B(n4010), .Z(n4127) );
  NANDN U4433 ( .A(n33875), .B(n4012), .Z(n4014) );
  XOR U4434 ( .A(b[25]), .B(a[16]), .Z(n4153) );
  NANDN U4435 ( .A(n33994), .B(n4153), .Z(n4013) );
  NAND U4436 ( .A(n4014), .B(n4013), .Z(n4126) );
  XOR U4437 ( .A(n4127), .B(n4126), .Z(n4129) );
  XNOR U4438 ( .A(n4128), .B(n4129), .Z(n4197) );
  XNOR U4439 ( .A(n4198), .B(n4197), .Z(n4199) );
  NANDN U4440 ( .A(n4016), .B(n4015), .Z(n4020) );
  NANDN U4441 ( .A(n4018), .B(n4017), .Z(n4019) );
  NAND U4442 ( .A(n4020), .B(n4019), .Z(n4200) );
  XNOR U4443 ( .A(n4199), .B(n4200), .Z(n4095) );
  NANDN U4444 ( .A(n4022), .B(n4021), .Z(n4026) );
  NAND U4445 ( .A(n4024), .B(n4023), .Z(n4025) );
  NAND U4446 ( .A(n4026), .B(n4025), .Z(n4096) );
  XNOR U4447 ( .A(n4095), .B(n4096), .Z(n4097) );
  XNOR U4448 ( .A(n4098), .B(n4097), .Z(n4085) );
  XNOR U4449 ( .A(n4086), .B(n4085), .Z(n4203) );
  XOR U4450 ( .A(n4204), .B(n4203), .Z(n4206) );
  XOR U4451 ( .A(n4205), .B(n4206), .Z(n4212) );
  XNOR U4452 ( .A(n4211), .B(n4212), .Z(n4217) );
  XOR U4453 ( .A(n4218), .B(n4217), .Z(n4040) );
  NANDN U4454 ( .A(n4028), .B(n4027), .Z(n4032) );
  NANDN U4455 ( .A(n4030), .B(n4029), .Z(n4031) );
  NAND U4456 ( .A(n4032), .B(n4031), .Z(n4039) );
  XOR U4457 ( .A(n4040), .B(n4039), .Z(n4042) );
  XNOR U4458 ( .A(n4041), .B(n4042), .Z(n4222) );
  NANDN U4459 ( .A(sreg[103]), .B(n4033), .Z(n4037) );
  NAND U4460 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U4461 ( .A(n4037), .B(n4036), .Z(n4221) );
  XOR U4462 ( .A(sreg[104]), .B(n4221), .Z(n4038) );
  XNOR U4463 ( .A(n4222), .B(n4038), .Z(c[104]) );
  NANDN U4464 ( .A(n4040), .B(n4039), .Z(n4044) );
  OR U4465 ( .A(n4042), .B(n4041), .Z(n4043) );
  AND U4466 ( .A(n4044), .B(n4043), .Z(n4228) );
  NAND U4467 ( .A(n4046), .B(n4045), .Z(n4050) );
  NAND U4468 ( .A(n4048), .B(n4047), .Z(n4049) );
  AND U4469 ( .A(n4050), .B(n4049), .Z(n4239) );
  NANDN U4470 ( .A(n4052), .B(n4051), .Z(n4056) );
  OR U4471 ( .A(n4054), .B(n4053), .Z(n4055) );
  AND U4472 ( .A(n4056), .B(n4055), .Z(n4251) );
  NANDN U4473 ( .A(n34634), .B(n4057), .Z(n4059) );
  XOR U4474 ( .A(b[29]), .B(a[13]), .Z(n4328) );
  NANDN U4475 ( .A(n34722), .B(n4328), .Z(n4058) );
  AND U4476 ( .A(n4059), .B(n4058), .Z(n4276) );
  NANDN U4477 ( .A(n34909), .B(n4060), .Z(n4062) );
  XOR U4478 ( .A(b[31]), .B(a[11]), .Z(n4316) );
  NANDN U4479 ( .A(n35145), .B(n4316), .Z(n4061) );
  AND U4480 ( .A(n4062), .B(n4061), .Z(n4275) );
  NANDN U4481 ( .A(n4063), .B(n32023), .Z(n4065) );
  XOR U4482 ( .A(b[15]), .B(a[27]), .Z(n4319) );
  NANDN U4483 ( .A(n31925), .B(n4319), .Z(n4064) );
  NAND U4484 ( .A(n4065), .B(n4064), .Z(n4274) );
  XOR U4485 ( .A(n4275), .B(n4274), .Z(n4277) );
  XOR U4486 ( .A(n4276), .B(n4277), .Z(n4257) );
  NANDN U4487 ( .A(n4066), .B(n4169), .Z(n4070) );
  OR U4488 ( .A(n4068), .B(n4067), .Z(n4069) );
  AND U4489 ( .A(n4070), .B(n4069), .Z(n4256) );
  XNOR U4490 ( .A(n4257), .B(n4256), .Z(n4258) );
  NANDN U4491 ( .A(n4072), .B(n4071), .Z(n4076) );
  OR U4492 ( .A(n4074), .B(n4073), .Z(n4075) );
  NAND U4493 ( .A(n4076), .B(n4075), .Z(n4259) );
  XNOR U4494 ( .A(n4258), .B(n4259), .Z(n4250) );
  XNOR U4495 ( .A(n4251), .B(n4250), .Z(n4252) );
  NANDN U4496 ( .A(n4078), .B(n4077), .Z(n4082) );
  OR U4497 ( .A(n4080), .B(n4079), .Z(n4081) );
  NAND U4498 ( .A(n4082), .B(n4081), .Z(n4253) );
  XOR U4499 ( .A(n4252), .B(n4253), .Z(n4238) );
  XOR U4500 ( .A(n4239), .B(n4238), .Z(n4241) );
  NANDN U4501 ( .A(n4084), .B(n4083), .Z(n4088) );
  NAND U4502 ( .A(n4086), .B(n4085), .Z(n4087) );
  AND U4503 ( .A(n4088), .B(n4087), .Z(n4240) );
  XOR U4504 ( .A(n4241), .B(n4240), .Z(n4235) );
  NANDN U4505 ( .A(n4090), .B(n4089), .Z(n4094) );
  NAND U4506 ( .A(n4092), .B(n4091), .Z(n4093) );
  AND U4507 ( .A(n4094), .B(n4093), .Z(n4232) );
  NANDN U4508 ( .A(n4096), .B(n4095), .Z(n4100) );
  NANDN U4509 ( .A(n4098), .B(n4097), .Z(n4099) );
  AND U4510 ( .A(n4100), .B(n4099), .Z(n4303) );
  NANDN U4511 ( .A(n4102), .B(n4101), .Z(n4106) );
  OR U4512 ( .A(n4104), .B(n4103), .Z(n4105) );
  AND U4513 ( .A(n4106), .B(n4105), .Z(n4298) );
  NANDN U4514 ( .A(n32996), .B(n4107), .Z(n4109) );
  XOR U4515 ( .A(b[21]), .B(a[21]), .Z(n4307) );
  NANDN U4516 ( .A(n33271), .B(n4307), .Z(n4108) );
  AND U4517 ( .A(n4109), .B(n4108), .Z(n4347) );
  XNOR U4518 ( .A(n4347), .B(n4346), .Z(n4348) );
  NANDN U4519 ( .A(n36210), .B(n4110), .Z(n4112) );
  XOR U4520 ( .A(b[39]), .B(a[3]), .Z(n4283) );
  NANDN U4521 ( .A(n36347), .B(n4283), .Z(n4111) );
  AND U4522 ( .A(n4112), .B(n4111), .Z(n4364) );
  XOR U4523 ( .A(b[41]), .B(b[40]), .Z(n4369) );
  XOR U4524 ( .A(b[41]), .B(a[0]), .Z(n4113) );
  NAND U4525 ( .A(n4369), .B(n4113), .Z(n4114) );
  OR U4526 ( .A(n4114), .B(n36733), .Z(n4116) );
  XOR U4527 ( .A(b[41]), .B(a[1]), .Z(n4370) );
  NAND U4528 ( .A(n36733), .B(n4370), .Z(n4115) );
  NAND U4529 ( .A(n4116), .B(n4115), .Z(n4365) );
  XOR U4530 ( .A(n4364), .B(n4365), .Z(n4349) );
  XNOR U4531 ( .A(n4348), .B(n4349), .Z(n4295) );
  NANDN U4532 ( .A(n210), .B(n4117), .Z(n4119) );
  XOR U4533 ( .A(b[9]), .B(a[33]), .Z(n4325) );
  NANDN U4534 ( .A(n30267), .B(n4325), .Z(n4118) );
  AND U4535 ( .A(n4119), .B(n4118), .Z(n4343) );
  NANDN U4536 ( .A(n31055), .B(n4120), .Z(n4122) );
  XOR U4537 ( .A(b[13]), .B(a[29]), .Z(n4292) );
  NANDN U4538 ( .A(n31293), .B(n4292), .Z(n4121) );
  AND U4539 ( .A(n4122), .B(n4121), .Z(n4341) );
  NANDN U4540 ( .A(n30482), .B(n4123), .Z(n4125) );
  XOR U4541 ( .A(b[11]), .B(a[31]), .Z(n4322) );
  NANDN U4542 ( .A(n30891), .B(n4322), .Z(n4124) );
  NAND U4543 ( .A(n4125), .B(n4124), .Z(n4340) );
  XNOR U4544 ( .A(n4341), .B(n4340), .Z(n4342) );
  XOR U4545 ( .A(n4343), .B(n4342), .Z(n4296) );
  XNOR U4546 ( .A(n4295), .B(n4296), .Z(n4297) );
  XNOR U4547 ( .A(n4298), .B(n4297), .Z(n4397) );
  NANDN U4548 ( .A(n4127), .B(n4126), .Z(n4131) );
  OR U4549 ( .A(n4129), .B(n4128), .Z(n4130) );
  AND U4550 ( .A(n4131), .B(n4130), .Z(n4395) );
  NANDN U4551 ( .A(n4133), .B(n4132), .Z(n4137) );
  NAND U4552 ( .A(n4135), .B(n4134), .Z(n4136) );
  NAND U4553 ( .A(n4137), .B(n4136), .Z(n4394) );
  XNOR U4554 ( .A(n4395), .B(n4394), .Z(n4396) );
  XOR U4555 ( .A(n4397), .B(n4396), .Z(n4402) );
  NANDN U4556 ( .A(n32013), .B(n4138), .Z(n4140) );
  XOR U4557 ( .A(b[17]), .B(a[25]), .Z(n4313) );
  NANDN U4558 ( .A(n32292), .B(n4313), .Z(n4139) );
  AND U4559 ( .A(n4140), .B(n4139), .Z(n4354) );
  NANDN U4560 ( .A(n34223), .B(n4141), .Z(n4143) );
  XOR U4561 ( .A(b[27]), .B(a[15]), .Z(n4337) );
  NANDN U4562 ( .A(n34458), .B(n4337), .Z(n4142) );
  AND U4563 ( .A(n4143), .B(n4142), .Z(n4353) );
  NANDN U4564 ( .A(n29499), .B(n4144), .Z(n4146) );
  XOR U4565 ( .A(b[7]), .B(a[35]), .Z(n4331) );
  NANDN U4566 ( .A(n29735), .B(n4331), .Z(n4145) );
  NAND U4567 ( .A(n4146), .B(n4145), .Z(n4352) );
  XOR U4568 ( .A(n4353), .B(n4352), .Z(n4355) );
  XOR U4569 ( .A(n4354), .B(n4355), .Z(n4389) );
  NANDN U4570 ( .A(n35260), .B(n4147), .Z(n4149) );
  XOR U4571 ( .A(b[33]), .B(a[9]), .Z(n4286) );
  NANDN U4572 ( .A(n35456), .B(n4286), .Z(n4148) );
  AND U4573 ( .A(n4149), .B(n4148), .Z(n4378) );
  NANDN U4574 ( .A(n28889), .B(n4150), .Z(n4152) );
  XOR U4575 ( .A(b[5]), .B(a[37]), .Z(n4366) );
  NANDN U4576 ( .A(n29138), .B(n4366), .Z(n4151) );
  AND U4577 ( .A(n4152), .B(n4151), .Z(n4377) );
  NANDN U4578 ( .A(n33875), .B(n4153), .Z(n4155) );
  XOR U4579 ( .A(b[25]), .B(a[17]), .Z(n4373) );
  NANDN U4580 ( .A(n33994), .B(n4373), .Z(n4154) );
  NAND U4581 ( .A(n4155), .B(n4154), .Z(n4376) );
  XOR U4582 ( .A(n4377), .B(n4376), .Z(n4379) );
  XNOR U4583 ( .A(n4378), .B(n4379), .Z(n4388) );
  XNOR U4584 ( .A(n4389), .B(n4388), .Z(n4390) );
  NANDN U4585 ( .A(n4157), .B(n4156), .Z(n4161) );
  OR U4586 ( .A(n4159), .B(n4158), .Z(n4160) );
  NAND U4587 ( .A(n4161), .B(n4160), .Z(n4391) );
  XNOR U4588 ( .A(n4390), .B(n4391), .Z(n4400) );
  NANDN U4589 ( .A(n35936), .B(n4162), .Z(n4164) );
  XOR U4590 ( .A(b[37]), .B(a[5]), .Z(n4334) );
  NANDN U4591 ( .A(n36047), .B(n4334), .Z(n4163) );
  AND U4592 ( .A(n4164), .B(n4163), .Z(n4270) );
  NANDN U4593 ( .A(n33866), .B(n4165), .Z(n4167) );
  XOR U4594 ( .A(b[23]), .B(a[19]), .Z(n4361) );
  NANDN U4595 ( .A(n33644), .B(n4361), .Z(n4166) );
  AND U4596 ( .A(n4167), .B(n4166), .Z(n4269) );
  NAND U4597 ( .A(b[39]), .B(b[40]), .Z(n4168) );
  AND U4598 ( .A(b[41]), .B(n4168), .Z(n36943) );
  ANDN U4599 ( .B(n36943), .A(n4169), .Z(n4268) );
  XOR U4600 ( .A(n4269), .B(n4268), .Z(n4271) );
  XOR U4601 ( .A(n4270), .B(n4271), .Z(n4383) );
  NANDN U4602 ( .A(n209), .B(n4170), .Z(n4172) );
  XOR U4603 ( .A(b[3]), .B(a[39]), .Z(n4358) );
  NANDN U4604 ( .A(n28941), .B(n4358), .Z(n4171) );
  AND U4605 ( .A(n4172), .B(n4171), .Z(n4264) );
  NANDN U4606 ( .A(n35611), .B(n4173), .Z(n4175) );
  XOR U4607 ( .A(b[35]), .B(a[7]), .Z(n4289) );
  NANDN U4608 ( .A(n35801), .B(n4289), .Z(n4174) );
  AND U4609 ( .A(n4175), .B(n4174), .Z(n4263) );
  NANDN U4610 ( .A(n32483), .B(n4176), .Z(n4178) );
  XOR U4611 ( .A(b[19]), .B(a[23]), .Z(n4310) );
  NANDN U4612 ( .A(n32823), .B(n4310), .Z(n4177) );
  NAND U4613 ( .A(n4178), .B(n4177), .Z(n4262) );
  XOR U4614 ( .A(n4263), .B(n4262), .Z(n4265) );
  XNOR U4615 ( .A(n4264), .B(n4265), .Z(n4382) );
  XNOR U4616 ( .A(n4383), .B(n4382), .Z(n4384) );
  NANDN U4617 ( .A(n4180), .B(n4179), .Z(n4184) );
  OR U4618 ( .A(n4182), .B(n4181), .Z(n4183) );
  NAND U4619 ( .A(n4184), .B(n4183), .Z(n4385) );
  XOR U4620 ( .A(n4384), .B(n4385), .Z(n4401) );
  XOR U4621 ( .A(n4400), .B(n4401), .Z(n4403) );
  XOR U4622 ( .A(n4402), .B(n4403), .Z(n4302) );
  NANDN U4623 ( .A(n4186), .B(n4185), .Z(n4190) );
  NANDN U4624 ( .A(n4188), .B(n4187), .Z(n4189) );
  AND U4625 ( .A(n4190), .B(n4189), .Z(n4246) );
  NANDN U4626 ( .A(n4192), .B(n4191), .Z(n4196) );
  NAND U4627 ( .A(n4194), .B(n4193), .Z(n4195) );
  AND U4628 ( .A(n4196), .B(n4195), .Z(n4245) );
  NANDN U4629 ( .A(n4198), .B(n4197), .Z(n4202) );
  NANDN U4630 ( .A(n4200), .B(n4199), .Z(n4201) );
  NAND U4631 ( .A(n4202), .B(n4201), .Z(n4244) );
  XOR U4632 ( .A(n4245), .B(n4244), .Z(n4247) );
  XNOR U4633 ( .A(n4246), .B(n4247), .Z(n4301) );
  XOR U4634 ( .A(n4302), .B(n4301), .Z(n4304) );
  XOR U4635 ( .A(n4303), .B(n4304), .Z(n4233) );
  XNOR U4636 ( .A(n4232), .B(n4233), .Z(n4234) );
  XOR U4637 ( .A(n4235), .B(n4234), .Z(n4407) );
  NANDN U4638 ( .A(n4204), .B(n4203), .Z(n4208) );
  NANDN U4639 ( .A(n4206), .B(n4205), .Z(n4207) );
  AND U4640 ( .A(n4208), .B(n4207), .Z(n4406) );
  XNOR U4641 ( .A(n4407), .B(n4406), .Z(n4408) );
  NANDN U4642 ( .A(n4210), .B(n4209), .Z(n4214) );
  NANDN U4643 ( .A(n4212), .B(n4211), .Z(n4213) );
  NAND U4644 ( .A(n4214), .B(n4213), .Z(n4409) );
  XNOR U4645 ( .A(n4408), .B(n4409), .Z(n4226) );
  NANDN U4646 ( .A(n4216), .B(n4215), .Z(n4220) );
  NAND U4647 ( .A(n4218), .B(n4217), .Z(n4219) );
  NAND U4648 ( .A(n4220), .B(n4219), .Z(n4227) );
  XOR U4649 ( .A(n4226), .B(n4227), .Z(n4229) );
  XOR U4650 ( .A(n4228), .B(n4229), .Z(n4224) );
  XNOR U4651 ( .A(sreg[105]), .B(n4225), .Z(n4223) );
  XOR U4652 ( .A(n4224), .B(n4223), .Z(c[105]) );
  XOR U4653 ( .A(sreg[106]), .B(n4604), .Z(n4606) );
  NANDN U4654 ( .A(n4227), .B(n4226), .Z(n4231) );
  OR U4655 ( .A(n4229), .B(n4228), .Z(n4230) );
  AND U4656 ( .A(n4231), .B(n4230), .Z(n4415) );
  NANDN U4657 ( .A(n4233), .B(n4232), .Z(n4237) );
  NAND U4658 ( .A(n4235), .B(n4234), .Z(n4236) );
  AND U4659 ( .A(n4237), .B(n4236), .Z(n4599) );
  NAND U4660 ( .A(n4239), .B(n4238), .Z(n4243) );
  NAND U4661 ( .A(n4241), .B(n4240), .Z(n4242) );
  NAND U4662 ( .A(n4243), .B(n4242), .Z(n4598) );
  XNOR U4663 ( .A(n4599), .B(n4598), .Z(n4601) );
  NANDN U4664 ( .A(n4245), .B(n4244), .Z(n4249) );
  OR U4665 ( .A(n4247), .B(n4246), .Z(n4248) );
  AND U4666 ( .A(n4249), .B(n4248), .Z(n4594) );
  NANDN U4667 ( .A(n4251), .B(n4250), .Z(n4255) );
  NANDN U4668 ( .A(n4253), .B(n4252), .Z(n4254) );
  AND U4669 ( .A(n4255), .B(n4254), .Z(n4593) );
  NANDN U4670 ( .A(n4257), .B(n4256), .Z(n4261) );
  NANDN U4671 ( .A(n4259), .B(n4258), .Z(n4260) );
  AND U4672 ( .A(n4261), .B(n4260), .Z(n4513) );
  NANDN U4673 ( .A(n4263), .B(n4262), .Z(n4267) );
  OR U4674 ( .A(n4265), .B(n4264), .Z(n4266) );
  AND U4675 ( .A(n4267), .B(n4266), .Z(n4523) );
  NANDN U4676 ( .A(n4269), .B(n4268), .Z(n4273) );
  OR U4677 ( .A(n4271), .B(n4270), .Z(n4272) );
  NAND U4678 ( .A(n4273), .B(n4272), .Z(n4522) );
  XNOR U4679 ( .A(n4523), .B(n4522), .Z(n4525) );
  NANDN U4680 ( .A(n4275), .B(n4274), .Z(n4279) );
  OR U4681 ( .A(n4277), .B(n4276), .Z(n4278) );
  AND U4682 ( .A(n4279), .B(n4278), .Z(n4547) );
  NAND U4683 ( .A(b[0]), .B(a[42]), .Z(n4280) );
  XNOR U4684 ( .A(b[1]), .B(n4280), .Z(n4282) );
  NANDN U4685 ( .A(b[0]), .B(a[41]), .Z(n4281) );
  NAND U4686 ( .A(n4282), .B(n4281), .Z(n4459) );
  XOR U4687 ( .A(b[42]), .B(b[41]), .Z(n36963) );
  IV U4688 ( .A(n36963), .Z(n36891) );
  ANDN U4689 ( .B(a[0]), .A(n36891), .Z(n4484) );
  NANDN U4690 ( .A(n36210), .B(n4283), .Z(n4285) );
  XOR U4691 ( .A(b[39]), .B(a[4]), .Z(n4583) );
  NANDN U4692 ( .A(n36347), .B(n4583), .Z(n4284) );
  AND U4693 ( .A(n4285), .B(n4284), .Z(n4457) );
  XNOR U4694 ( .A(n4484), .B(n4457), .Z(n4458) );
  XNOR U4695 ( .A(n4459), .B(n4458), .Z(n4544) );
  NANDN U4696 ( .A(n35260), .B(n4286), .Z(n4288) );
  XOR U4697 ( .A(b[33]), .B(a[10]), .Z(n4430) );
  NANDN U4698 ( .A(n35456), .B(n4430), .Z(n4287) );
  AND U4699 ( .A(n4288), .B(n4287), .Z(n4497) );
  NANDN U4700 ( .A(n35611), .B(n4289), .Z(n4291) );
  XOR U4701 ( .A(b[35]), .B(a[8]), .Z(n4433) );
  NANDN U4702 ( .A(n35801), .B(n4433), .Z(n4290) );
  AND U4703 ( .A(n4291), .B(n4290), .Z(n4495) );
  NANDN U4704 ( .A(n31055), .B(n4292), .Z(n4294) );
  XOR U4705 ( .A(b[13]), .B(a[30]), .Z(n4580) );
  NANDN U4706 ( .A(n31293), .B(n4580), .Z(n4293) );
  NAND U4707 ( .A(n4294), .B(n4293), .Z(n4494) );
  XNOR U4708 ( .A(n4495), .B(n4494), .Z(n4496) );
  XOR U4709 ( .A(n4497), .B(n4496), .Z(n4545) );
  XNOR U4710 ( .A(n4544), .B(n4545), .Z(n4546) );
  XNOR U4711 ( .A(n4547), .B(n4546), .Z(n4524) );
  XOR U4712 ( .A(n4525), .B(n4524), .Z(n4511) );
  NANDN U4713 ( .A(n4296), .B(n4295), .Z(n4300) );
  NANDN U4714 ( .A(n4298), .B(n4297), .Z(n4299) );
  AND U4715 ( .A(n4300), .B(n4299), .Z(n4510) );
  XNOR U4716 ( .A(n4511), .B(n4510), .Z(n4512) );
  XNOR U4717 ( .A(n4513), .B(n4512), .Z(n4592) );
  XOR U4718 ( .A(n4593), .B(n4592), .Z(n4595) );
  XOR U4719 ( .A(n4594), .B(n4595), .Z(n4421) );
  NANDN U4720 ( .A(n4302), .B(n4301), .Z(n4306) );
  NANDN U4721 ( .A(n4304), .B(n4303), .Z(n4305) );
  AND U4722 ( .A(n4306), .B(n4305), .Z(n4419) );
  NANDN U4723 ( .A(n32996), .B(n4307), .Z(n4309) );
  XOR U4724 ( .A(b[21]), .B(a[22]), .Z(n4462) );
  NANDN U4725 ( .A(n33271), .B(n4462), .Z(n4308) );
  AND U4726 ( .A(n4309), .B(n4308), .Z(n4557) );
  NANDN U4727 ( .A(n32483), .B(n4310), .Z(n4312) );
  XOR U4728 ( .A(b[19]), .B(a[24]), .Z(n4442) );
  NANDN U4729 ( .A(n32823), .B(n4442), .Z(n4311) );
  NAND U4730 ( .A(n4312), .B(n4311), .Z(n4556) );
  XNOR U4731 ( .A(n4557), .B(n4556), .Z(n4559) );
  NANDN U4732 ( .A(n32013), .B(n4313), .Z(n4315) );
  XOR U4733 ( .A(b[17]), .B(a[26]), .Z(n4445) );
  NANDN U4734 ( .A(n32292), .B(n4445), .Z(n4314) );
  AND U4735 ( .A(n4315), .B(n4314), .Z(n4454) );
  NANDN U4736 ( .A(n34909), .B(n4316), .Z(n4318) );
  XOR U4737 ( .A(b[31]), .B(a[12]), .Z(n4439) );
  NANDN U4738 ( .A(n35145), .B(n4439), .Z(n4317) );
  AND U4739 ( .A(n4318), .B(n4317), .Z(n4452) );
  NANDN U4740 ( .A(n31536), .B(n4319), .Z(n4321) );
  XOR U4741 ( .A(b[15]), .B(a[28]), .Z(n4436) );
  NANDN U4742 ( .A(n31925), .B(n4436), .Z(n4320) );
  NAND U4743 ( .A(n4321), .B(n4320), .Z(n4451) );
  XNOR U4744 ( .A(n4452), .B(n4451), .Z(n4453) );
  XNOR U4745 ( .A(n4454), .B(n4453), .Z(n4558) );
  XOR U4746 ( .A(n4559), .B(n4558), .Z(n4553) );
  NANDN U4747 ( .A(n30482), .B(n4322), .Z(n4324) );
  XOR U4748 ( .A(b[11]), .B(a[32]), .Z(n4568) );
  NANDN U4749 ( .A(n30891), .B(n4568), .Z(n4323) );
  AND U4750 ( .A(n4324), .B(n4323), .Z(n4588) );
  NANDN U4751 ( .A(n210), .B(n4325), .Z(n4327) );
  XOR U4752 ( .A(b[9]), .B(a[34]), .Z(n4571) );
  NANDN U4753 ( .A(n30267), .B(n4571), .Z(n4326) );
  AND U4754 ( .A(n4327), .B(n4326), .Z(n4587) );
  NANDN U4755 ( .A(n34634), .B(n4328), .Z(n4330) );
  XOR U4756 ( .A(b[29]), .B(a[14]), .Z(n4574) );
  NANDN U4757 ( .A(n34722), .B(n4574), .Z(n4329) );
  NAND U4758 ( .A(n4330), .B(n4329), .Z(n4586) );
  XOR U4759 ( .A(n4587), .B(n4586), .Z(n4589) );
  XOR U4760 ( .A(n4588), .B(n4589), .Z(n4551) );
  NANDN U4761 ( .A(n29499), .B(n4331), .Z(n4333) );
  XOR U4762 ( .A(b[7]), .B(a[36]), .Z(n4485) );
  NANDN U4763 ( .A(n29735), .B(n4485), .Z(n4332) );
  AND U4764 ( .A(n4333), .B(n4332), .Z(n4502) );
  NANDN U4765 ( .A(n35936), .B(n4334), .Z(n4336) );
  XOR U4766 ( .A(b[37]), .B(a[6]), .Z(n4577) );
  NANDN U4767 ( .A(n36047), .B(n4577), .Z(n4335) );
  AND U4768 ( .A(n4336), .B(n4335), .Z(n4501) );
  NANDN U4769 ( .A(n34223), .B(n4337), .Z(n4339) );
  XOR U4770 ( .A(b[27]), .B(a[16]), .Z(n4491) );
  NANDN U4771 ( .A(n34458), .B(n4491), .Z(n4338) );
  NAND U4772 ( .A(n4339), .B(n4338), .Z(n4500) );
  XOR U4773 ( .A(n4501), .B(n4500), .Z(n4503) );
  XNOR U4774 ( .A(n4502), .B(n4503), .Z(n4550) );
  XNOR U4775 ( .A(n4551), .B(n4550), .Z(n4552) );
  XOR U4776 ( .A(n4553), .B(n4552), .Z(n4530) );
  NANDN U4777 ( .A(n4341), .B(n4340), .Z(n4345) );
  NANDN U4778 ( .A(n4343), .B(n4342), .Z(n4344) );
  NAND U4779 ( .A(n4345), .B(n4344), .Z(n4529) );
  NANDN U4780 ( .A(n4347), .B(n4346), .Z(n4351) );
  NANDN U4781 ( .A(n4349), .B(n4348), .Z(n4350) );
  NAND U4782 ( .A(n4351), .B(n4350), .Z(n4528) );
  XOR U4783 ( .A(n4529), .B(n4528), .Z(n4531) );
  XNOR U4784 ( .A(n4530), .B(n4531), .Z(n4543) );
  NANDN U4785 ( .A(n4353), .B(n4352), .Z(n4357) );
  OR U4786 ( .A(n4355), .B(n4354), .Z(n4356) );
  NAND U4787 ( .A(n4357), .B(n4356), .Z(n4536) );
  NANDN U4788 ( .A(n209), .B(n4358), .Z(n4360) );
  XOR U4789 ( .A(b[3]), .B(a[40]), .Z(n4478) );
  NANDN U4790 ( .A(n28941), .B(n4478), .Z(n4359) );
  AND U4791 ( .A(n4360), .B(n4359), .Z(n4507) );
  NANDN U4792 ( .A(n33866), .B(n4361), .Z(n4363) );
  XOR U4793 ( .A(b[23]), .B(a[20]), .Z(n4448) );
  NANDN U4794 ( .A(n33644), .B(n4448), .Z(n4362) );
  NAND U4795 ( .A(n4363), .B(n4362), .Z(n4506) );
  XNOR U4796 ( .A(n4507), .B(n4506), .Z(n4509) );
  ANDN U4797 ( .B(n4365), .A(n4364), .Z(n4508) );
  XOR U4798 ( .A(n4509), .B(n4508), .Z(n4535) );
  NANDN U4799 ( .A(n28889), .B(n4366), .Z(n4368) );
  XOR U4800 ( .A(b[5]), .B(a[38]), .Z(n4488) );
  NANDN U4801 ( .A(n29138), .B(n4488), .Z(n4367) );
  AND U4802 ( .A(n4368), .B(n4367), .Z(n4565) );
  ANDN U4803 ( .B(n4369), .A(n36733), .Z(n36735) );
  IV U4804 ( .A(n36735), .Z(n36480) );
  NANDN U4805 ( .A(n36480), .B(n4370), .Z(n4372) );
  XOR U4806 ( .A(b[41]), .B(a[2]), .Z(n4468) );
  NANDN U4807 ( .A(n36594), .B(n4468), .Z(n4371) );
  AND U4808 ( .A(n4372), .B(n4371), .Z(n4563) );
  NANDN U4809 ( .A(n33875), .B(n4373), .Z(n4375) );
  XOR U4810 ( .A(b[25]), .B(a[18]), .Z(n4481) );
  NANDN U4811 ( .A(n33994), .B(n4481), .Z(n4374) );
  NAND U4812 ( .A(n4375), .B(n4374), .Z(n4562) );
  XNOR U4813 ( .A(n4563), .B(n4562), .Z(n4564) );
  XNOR U4814 ( .A(n4565), .B(n4564), .Z(n4534) );
  XOR U4815 ( .A(n4535), .B(n4534), .Z(n4537) );
  XNOR U4816 ( .A(n4536), .B(n4537), .Z(n4540) );
  NANDN U4817 ( .A(n4377), .B(n4376), .Z(n4381) );
  OR U4818 ( .A(n4379), .B(n4378), .Z(n4380) );
  AND U4819 ( .A(n4381), .B(n4380), .Z(n4541) );
  XOR U4820 ( .A(n4540), .B(n4541), .Z(n4542) );
  XNOR U4821 ( .A(n4543), .B(n4542), .Z(n4517) );
  NANDN U4822 ( .A(n4383), .B(n4382), .Z(n4387) );
  NANDN U4823 ( .A(n4385), .B(n4384), .Z(n4386) );
  AND U4824 ( .A(n4387), .B(n4386), .Z(n4425) );
  NANDN U4825 ( .A(n4389), .B(n4388), .Z(n4393) );
  NANDN U4826 ( .A(n4391), .B(n4390), .Z(n4392) );
  NAND U4827 ( .A(n4393), .B(n4392), .Z(n4424) );
  XNOR U4828 ( .A(n4425), .B(n4424), .Z(n4427) );
  NANDN U4829 ( .A(n4395), .B(n4394), .Z(n4399) );
  NAND U4830 ( .A(n4397), .B(n4396), .Z(n4398) );
  AND U4831 ( .A(n4399), .B(n4398), .Z(n4426) );
  XNOR U4832 ( .A(n4427), .B(n4426), .Z(n4516) );
  XOR U4833 ( .A(n4517), .B(n4516), .Z(n4518) );
  NANDN U4834 ( .A(n4401), .B(n4400), .Z(n4405) );
  OR U4835 ( .A(n4403), .B(n4402), .Z(n4404) );
  NAND U4836 ( .A(n4405), .B(n4404), .Z(n4519) );
  XNOR U4837 ( .A(n4518), .B(n4519), .Z(n4418) );
  XNOR U4838 ( .A(n4419), .B(n4418), .Z(n4420) );
  XNOR U4839 ( .A(n4421), .B(n4420), .Z(n4600) );
  XOR U4840 ( .A(n4601), .B(n4600), .Z(n4413) );
  NANDN U4841 ( .A(n4407), .B(n4406), .Z(n4411) );
  NANDN U4842 ( .A(n4409), .B(n4408), .Z(n4410) );
  NAND U4843 ( .A(n4411), .B(n4410), .Z(n4412) );
  XNOR U4844 ( .A(n4413), .B(n4412), .Z(n4414) );
  XNOR U4845 ( .A(n4415), .B(n4414), .Z(n4605) );
  XNOR U4846 ( .A(n4606), .B(n4605), .Z(c[106]) );
  NANDN U4847 ( .A(n4413), .B(n4412), .Z(n4417) );
  NANDN U4848 ( .A(n4415), .B(n4414), .Z(n4416) );
  AND U4849 ( .A(n4417), .B(n4416), .Z(n4617) );
  NANDN U4850 ( .A(n4419), .B(n4418), .Z(n4423) );
  NANDN U4851 ( .A(n4421), .B(n4420), .Z(n4422) );
  AND U4852 ( .A(n4423), .B(n4422), .Z(n4803) );
  NANDN U4853 ( .A(n4425), .B(n4424), .Z(n4429) );
  NAND U4854 ( .A(n4427), .B(n4426), .Z(n4428) );
  AND U4855 ( .A(n4429), .B(n4428), .Z(n4627) );
  NANDN U4856 ( .A(n35260), .B(n4430), .Z(n4432) );
  XOR U4857 ( .A(b[33]), .B(a[11]), .Z(n4725) );
  NANDN U4858 ( .A(n35456), .B(n4725), .Z(n4431) );
  AND U4859 ( .A(n4432), .B(n4431), .Z(n4767) );
  NANDN U4860 ( .A(n35611), .B(n4433), .Z(n4435) );
  XOR U4861 ( .A(b[35]), .B(a[9]), .Z(n4728) );
  NANDN U4862 ( .A(n35801), .B(n4728), .Z(n4434) );
  AND U4863 ( .A(n4435), .B(n4434), .Z(n4766) );
  NANDN U4864 ( .A(n31536), .B(n4436), .Z(n4438) );
  XOR U4865 ( .A(b[15]), .B(a[29]), .Z(n4698) );
  NANDN U4866 ( .A(n31925), .B(n4698), .Z(n4437) );
  NAND U4867 ( .A(n4438), .B(n4437), .Z(n4765) );
  XOR U4868 ( .A(n4766), .B(n4765), .Z(n4768) );
  XOR U4869 ( .A(n4767), .B(n4768), .Z(n4656) );
  NANDN U4870 ( .A(n34909), .B(n4439), .Z(n4441) );
  XOR U4871 ( .A(b[31]), .B(a[13]), .Z(n4749) );
  NANDN U4872 ( .A(n35145), .B(n4749), .Z(n4440) );
  AND U4873 ( .A(n4441), .B(n4440), .Z(n4712) );
  NANDN U4874 ( .A(n32483), .B(n4442), .Z(n4444) );
  XOR U4875 ( .A(b[19]), .B(a[25]), .Z(n4695) );
  NANDN U4876 ( .A(n32823), .B(n4695), .Z(n4443) );
  AND U4877 ( .A(n4444), .B(n4443), .Z(n4711) );
  NANDN U4878 ( .A(n32013), .B(n4445), .Z(n4447) );
  XOR U4879 ( .A(b[17]), .B(a[27]), .Z(n4701) );
  NANDN U4880 ( .A(n32292), .B(n4701), .Z(n4446) );
  NAND U4881 ( .A(n4447), .B(n4446), .Z(n4710) );
  XOR U4882 ( .A(n4711), .B(n4710), .Z(n4713) );
  XOR U4883 ( .A(n4712), .B(n4713), .Z(n4655) );
  NAND U4884 ( .A(n33492), .B(n4448), .Z(n4450) );
  XNOR U4885 ( .A(b[23]), .B(a[21]), .Z(n4669) );
  NANDN U4886 ( .A(n4669), .B(n33868), .Z(n4449) );
  AND U4887 ( .A(n4450), .B(n4449), .Z(n4654) );
  XOR U4888 ( .A(n4655), .B(n4654), .Z(n4657) );
  XOR U4889 ( .A(n4656), .B(n4657), .Z(n4784) );
  NANDN U4890 ( .A(n4452), .B(n4451), .Z(n4456) );
  NANDN U4891 ( .A(n4454), .B(n4453), .Z(n4455) );
  AND U4892 ( .A(n4456), .B(n4455), .Z(n4645) );
  NANDN U4893 ( .A(n4457), .B(n4484), .Z(n4461) );
  NANDN U4894 ( .A(n4459), .B(n4458), .Z(n4460) );
  AND U4895 ( .A(n4461), .B(n4460), .Z(n4643) );
  NANDN U4896 ( .A(n32996), .B(n4462), .Z(n4464) );
  XOR U4897 ( .A(b[21]), .B(a[23]), .Z(n4746) );
  NANDN U4898 ( .A(n33271), .B(n4746), .Z(n4463) );
  NAND U4899 ( .A(n4464), .B(n4463), .Z(n4689) );
  NAND U4900 ( .A(b[0]), .B(a[43]), .Z(n4465) );
  XNOR U4901 ( .A(b[1]), .B(n4465), .Z(n4467) );
  NANDN U4902 ( .A(b[0]), .B(a[42]), .Z(n4466) );
  NAND U4903 ( .A(n4467), .B(n4466), .Z(n4690) );
  XNOR U4904 ( .A(n4689), .B(n4690), .Z(n4691) );
  NANDN U4905 ( .A(n36480), .B(n4468), .Z(n4470) );
  XOR U4906 ( .A(b[41]), .B(a[3]), .Z(n4707) );
  NANDN U4907 ( .A(n36594), .B(n4707), .Z(n4469) );
  AND U4908 ( .A(n4470), .B(n4469), .Z(n4672) );
  XOR U4909 ( .A(b[43]), .B(a[1]), .Z(n4759) );
  NANDN U4910 ( .A(n36891), .B(n4759), .Z(n4477) );
  ANDN U4911 ( .B(b[42]), .A(b[43]), .Z(n4471) );
  NAND U4912 ( .A(n4471), .B(a[0]), .Z(n4474) );
  NAND U4913 ( .A(b[41]), .B(b[42]), .Z(n4472) );
  NAND U4914 ( .A(b[43]), .B(n4472), .Z(n37090) );
  OR U4915 ( .A(a[0]), .B(n37090), .Z(n4473) );
  NAND U4916 ( .A(n4474), .B(n4473), .Z(n4475) );
  NAND U4917 ( .A(n36891), .B(n4475), .Z(n4476) );
  NAND U4918 ( .A(n4477), .B(n4476), .Z(n4673) );
  XOR U4919 ( .A(n4672), .B(n4673), .Z(n4692) );
  XNOR U4920 ( .A(n4691), .B(n4692), .Z(n4642) );
  XNOR U4921 ( .A(n4643), .B(n4642), .Z(n4644) );
  XNOR U4922 ( .A(n4645), .B(n4644), .Z(n4783) );
  XNOR U4923 ( .A(n4784), .B(n4783), .Z(n4786) );
  NANDN U4924 ( .A(n209), .B(n4478), .Z(n4480) );
  XOR U4925 ( .A(b[3]), .B(a[41]), .Z(n4666) );
  NANDN U4926 ( .A(n28941), .B(n4666), .Z(n4479) );
  AND U4927 ( .A(n4480), .B(n4479), .Z(n4741) );
  NANDN U4928 ( .A(n33875), .B(n4481), .Z(n4483) );
  XOR U4929 ( .A(b[25]), .B(a[19]), .Z(n4722) );
  NANDN U4930 ( .A(n33994), .B(n4722), .Z(n4482) );
  NAND U4931 ( .A(n4483), .B(n4482), .Z(n4740) );
  XNOR U4932 ( .A(n4741), .B(n4740), .Z(n4743) );
  IV U4933 ( .A(n37090), .Z(n37180) );
  ANDN U4934 ( .B(n37180), .A(n4484), .Z(n4742) );
  XOR U4935 ( .A(n4743), .B(n4742), .Z(n4778) );
  NANDN U4936 ( .A(n29499), .B(n4485), .Z(n4487) );
  XOR U4937 ( .A(b[7]), .B(a[37]), .Z(n4677) );
  NANDN U4938 ( .A(n29735), .B(n4677), .Z(n4486) );
  AND U4939 ( .A(n4487), .B(n4486), .Z(n4685) );
  NANDN U4940 ( .A(n28889), .B(n4488), .Z(n4490) );
  XOR U4941 ( .A(b[5]), .B(a[39]), .Z(n4755) );
  NANDN U4942 ( .A(n29138), .B(n4755), .Z(n4489) );
  AND U4943 ( .A(n4490), .B(n4489), .Z(n4684) );
  NANDN U4944 ( .A(n34223), .B(n4491), .Z(n4493) );
  XOR U4945 ( .A(b[27]), .B(a[17]), .Z(n4762) );
  NANDN U4946 ( .A(n34458), .B(n4762), .Z(n4492) );
  NAND U4947 ( .A(n4493), .B(n4492), .Z(n4683) );
  XOR U4948 ( .A(n4684), .B(n4683), .Z(n4686) );
  XNOR U4949 ( .A(n4685), .B(n4686), .Z(n4777) );
  XNOR U4950 ( .A(n4778), .B(n4777), .Z(n4780) );
  NANDN U4951 ( .A(n4495), .B(n4494), .Z(n4499) );
  NANDN U4952 ( .A(n4497), .B(n4496), .Z(n4498) );
  AND U4953 ( .A(n4499), .B(n4498), .Z(n4779) );
  XOR U4954 ( .A(n4780), .B(n4779), .Z(n4639) );
  NANDN U4955 ( .A(n4501), .B(n4500), .Z(n4505) );
  OR U4956 ( .A(n4503), .B(n4502), .Z(n4504) );
  AND U4957 ( .A(n4505), .B(n4504), .Z(n4637) );
  XNOR U4958 ( .A(n4637), .B(n4636), .Z(n4638) );
  XNOR U4959 ( .A(n4639), .B(n4638), .Z(n4785) );
  XOR U4960 ( .A(n4786), .B(n4785), .Z(n4625) );
  NANDN U4961 ( .A(n4511), .B(n4510), .Z(n4515) );
  NANDN U4962 ( .A(n4513), .B(n4512), .Z(n4514) );
  NAND U4963 ( .A(n4515), .B(n4514), .Z(n4624) );
  XNOR U4964 ( .A(n4625), .B(n4624), .Z(n4626) );
  XNOR U4965 ( .A(n4627), .B(n4626), .Z(n4623) );
  NAND U4966 ( .A(n4517), .B(n4516), .Z(n4521) );
  NANDN U4967 ( .A(n4519), .B(n4518), .Z(n4520) );
  AND U4968 ( .A(n4521), .B(n4520), .Z(n4621) );
  NANDN U4969 ( .A(n4523), .B(n4522), .Z(n4527) );
  NAND U4970 ( .A(n4525), .B(n4524), .Z(n4526) );
  NAND U4971 ( .A(n4527), .B(n4526), .Z(n4791) );
  NAND U4972 ( .A(n4529), .B(n4528), .Z(n4533) );
  NAND U4973 ( .A(n4531), .B(n4530), .Z(n4532) );
  NAND U4974 ( .A(n4533), .B(n4532), .Z(n4790) );
  NAND U4975 ( .A(n4535), .B(n4534), .Z(n4539) );
  NAND U4976 ( .A(n4537), .B(n4536), .Z(n4538) );
  NAND U4977 ( .A(n4539), .B(n4538), .Z(n4789) );
  XOR U4978 ( .A(n4790), .B(n4789), .Z(n4792) );
  XNOR U4979 ( .A(n4791), .B(n4792), .Z(n4798) );
  NANDN U4980 ( .A(n4545), .B(n4544), .Z(n4549) );
  NANDN U4981 ( .A(n4547), .B(n4546), .Z(n4548) );
  AND U4982 ( .A(n4549), .B(n4548), .Z(n4649) );
  NANDN U4983 ( .A(n4551), .B(n4550), .Z(n4555) );
  NANDN U4984 ( .A(n4553), .B(n4552), .Z(n4554) );
  AND U4985 ( .A(n4555), .B(n4554), .Z(n4648) );
  XNOR U4986 ( .A(n4649), .B(n4648), .Z(n4651) );
  NANDN U4987 ( .A(n4557), .B(n4556), .Z(n4561) );
  NAND U4988 ( .A(n4559), .B(n4558), .Z(n4560) );
  AND U4989 ( .A(n4561), .B(n4560), .Z(n4633) );
  NANDN U4990 ( .A(n4563), .B(n4562), .Z(n4567) );
  NANDN U4991 ( .A(n4565), .B(n4564), .Z(n4566) );
  AND U4992 ( .A(n4567), .B(n4566), .Z(n4631) );
  NANDN U4993 ( .A(n30482), .B(n4568), .Z(n4570) );
  XOR U4994 ( .A(b[11]), .B(a[33]), .Z(n4731) );
  NANDN U4995 ( .A(n30891), .B(n4731), .Z(n4569) );
  AND U4996 ( .A(n4570), .B(n4569), .Z(n4736) );
  NANDN U4997 ( .A(n210), .B(n4571), .Z(n4573) );
  XOR U4998 ( .A(b[9]), .B(a[35]), .Z(n4716) );
  NANDN U4999 ( .A(n30267), .B(n4716), .Z(n4572) );
  AND U5000 ( .A(n4573), .B(n4572), .Z(n4735) );
  NANDN U5001 ( .A(n34634), .B(n4574), .Z(n4576) );
  XOR U5002 ( .A(b[29]), .B(a[15]), .Z(n4680) );
  NANDN U5003 ( .A(n34722), .B(n4680), .Z(n4575) );
  NAND U5004 ( .A(n4576), .B(n4575), .Z(n4734) );
  XOR U5005 ( .A(n4735), .B(n4734), .Z(n4737) );
  XOR U5006 ( .A(n4736), .B(n4737), .Z(n4772) );
  NANDN U5007 ( .A(n35936), .B(n4577), .Z(n4579) );
  XOR U5008 ( .A(b[37]), .B(a[7]), .Z(n4719) );
  NANDN U5009 ( .A(n36047), .B(n4719), .Z(n4578) );
  AND U5010 ( .A(n4579), .B(n4578), .Z(n4662) );
  NANDN U5011 ( .A(n31055), .B(n4580), .Z(n4582) );
  XOR U5012 ( .A(b[13]), .B(a[31]), .Z(n4752) );
  NANDN U5013 ( .A(n31293), .B(n4752), .Z(n4581) );
  AND U5014 ( .A(n4582), .B(n4581), .Z(n4661) );
  NANDN U5015 ( .A(n36210), .B(n4583), .Z(n4585) );
  XOR U5016 ( .A(b[39]), .B(a[5]), .Z(n4674) );
  NANDN U5017 ( .A(n36347), .B(n4674), .Z(n4584) );
  NAND U5018 ( .A(n4585), .B(n4584), .Z(n4660) );
  XOR U5019 ( .A(n4661), .B(n4660), .Z(n4663) );
  XNOR U5020 ( .A(n4662), .B(n4663), .Z(n4771) );
  XNOR U5021 ( .A(n4772), .B(n4771), .Z(n4774) );
  NANDN U5022 ( .A(n4587), .B(n4586), .Z(n4591) );
  OR U5023 ( .A(n4589), .B(n4588), .Z(n4590) );
  AND U5024 ( .A(n4591), .B(n4590), .Z(n4773) );
  XNOR U5025 ( .A(n4774), .B(n4773), .Z(n4630) );
  XNOR U5026 ( .A(n4631), .B(n4630), .Z(n4632) );
  XNOR U5027 ( .A(n4633), .B(n4632), .Z(n4650) );
  XNOR U5028 ( .A(n4651), .B(n4650), .Z(n4795) );
  XNOR U5029 ( .A(n4796), .B(n4795), .Z(n4797) );
  XOR U5030 ( .A(n4798), .B(n4797), .Z(n4620) );
  XOR U5031 ( .A(n4621), .B(n4620), .Z(n4622) );
  XOR U5032 ( .A(n4623), .B(n4622), .Z(n4802) );
  NANDN U5033 ( .A(n4593), .B(n4592), .Z(n4597) );
  OR U5034 ( .A(n4595), .B(n4594), .Z(n4596) );
  AND U5035 ( .A(n4597), .B(n4596), .Z(n4801) );
  XOR U5036 ( .A(n4802), .B(n4801), .Z(n4804) );
  XOR U5037 ( .A(n4803), .B(n4804), .Z(n4615) );
  NANDN U5038 ( .A(n4599), .B(n4598), .Z(n4603) );
  NAND U5039 ( .A(n4601), .B(n4600), .Z(n4602) );
  AND U5040 ( .A(n4603), .B(n4602), .Z(n4614) );
  XNOR U5041 ( .A(n4615), .B(n4614), .Z(n4616) );
  XNOR U5042 ( .A(n4617), .B(n4616), .Z(n4609) );
  XNOR U5043 ( .A(sreg[107]), .B(n4609), .Z(n4611) );
  OR U5044 ( .A(sreg[106]), .B(n4604), .Z(n4608) );
  NAND U5045 ( .A(n4606), .B(n4605), .Z(n4607) );
  NAND U5046 ( .A(n4608), .B(n4607), .Z(n4610) );
  XNOR U5047 ( .A(n4611), .B(n4610), .Z(c[107]) );
  NANDN U5048 ( .A(sreg[107]), .B(n4609), .Z(n4613) );
  NAND U5049 ( .A(n4611), .B(n4610), .Z(n4612) );
  AND U5050 ( .A(n4613), .B(n4612), .Z(n4808) );
  NANDN U5051 ( .A(n4615), .B(n4614), .Z(n4619) );
  NANDN U5052 ( .A(n4617), .B(n4616), .Z(n4618) );
  AND U5053 ( .A(n4619), .B(n4618), .Z(n4813) );
  NANDN U5054 ( .A(n4625), .B(n4624), .Z(n4629) );
  NANDN U5055 ( .A(n4627), .B(n4626), .Z(n4628) );
  AND U5056 ( .A(n4629), .B(n4628), .Z(n5003) );
  NANDN U5057 ( .A(n4631), .B(n4630), .Z(n4635) );
  NANDN U5058 ( .A(n4633), .B(n4632), .Z(n4634) );
  AND U5059 ( .A(n4635), .B(n4634), .Z(n4993) );
  NANDN U5060 ( .A(n4637), .B(n4636), .Z(n4641) );
  NANDN U5061 ( .A(n4639), .B(n4638), .Z(n4640) );
  AND U5062 ( .A(n4641), .B(n4640), .Z(n4992) );
  NANDN U5063 ( .A(n4643), .B(n4642), .Z(n4647) );
  NANDN U5064 ( .A(n4645), .B(n4644), .Z(n4646) );
  NAND U5065 ( .A(n4647), .B(n4646), .Z(n4991) );
  XOR U5066 ( .A(n4992), .B(n4991), .Z(n4994) );
  XOR U5067 ( .A(n4993), .B(n4994), .Z(n4998) );
  NANDN U5068 ( .A(n4649), .B(n4648), .Z(n4653) );
  NAND U5069 ( .A(n4651), .B(n4650), .Z(n4652) );
  AND U5070 ( .A(n4653), .B(n4652), .Z(n4997) );
  XNOR U5071 ( .A(n4998), .B(n4997), .Z(n5000) );
  NANDN U5072 ( .A(n4655), .B(n4654), .Z(n4659) );
  OR U5073 ( .A(n4657), .B(n4656), .Z(n4658) );
  AND U5074 ( .A(n4659), .B(n4658), .Z(n4822) );
  NANDN U5075 ( .A(n4661), .B(n4660), .Z(n4665) );
  OR U5076 ( .A(n4663), .B(n4662), .Z(n4664) );
  AND U5077 ( .A(n4665), .B(n4664), .Z(n4976) );
  NANDN U5078 ( .A(n209), .B(n4666), .Z(n4668) );
  XOR U5079 ( .A(b[3]), .B(a[42]), .Z(n4882) );
  NANDN U5080 ( .A(n28941), .B(n4882), .Z(n4667) );
  AND U5081 ( .A(n4668), .B(n4667), .Z(n4841) );
  NANDN U5082 ( .A(n4669), .B(n33492), .Z(n4671) );
  XOR U5083 ( .A(b[23]), .B(a[22]), .Z(n4860) );
  NANDN U5084 ( .A(n33644), .B(n4860), .Z(n4670) );
  NAND U5085 ( .A(n4671), .B(n4670), .Z(n4840) );
  XNOR U5086 ( .A(n4841), .B(n4840), .Z(n4843) );
  ANDN U5087 ( .B(n4673), .A(n4672), .Z(n4842) );
  XOR U5088 ( .A(n4843), .B(n4842), .Z(n4973) );
  NANDN U5089 ( .A(n36210), .B(n4674), .Z(n4676) );
  XOR U5090 ( .A(b[39]), .B(a[6]), .Z(n4885) );
  NANDN U5091 ( .A(n36347), .B(n4885), .Z(n4675) );
  AND U5092 ( .A(n4676), .B(n4675), .Z(n4915) );
  NANDN U5093 ( .A(n29499), .B(n4677), .Z(n4679) );
  XOR U5094 ( .A(b[7]), .B(a[38]), .Z(n4891) );
  NANDN U5095 ( .A(n29735), .B(n4891), .Z(n4678) );
  AND U5096 ( .A(n4679), .B(n4678), .Z(n4913) );
  NANDN U5097 ( .A(n34634), .B(n4680), .Z(n4682) );
  XOR U5098 ( .A(b[29]), .B(a[16]), .Z(n4921) );
  NANDN U5099 ( .A(n34722), .B(n4921), .Z(n4681) );
  NAND U5100 ( .A(n4682), .B(n4681), .Z(n4912) );
  XNOR U5101 ( .A(n4913), .B(n4912), .Z(n4914) );
  XOR U5102 ( .A(n4915), .B(n4914), .Z(n4974) );
  XNOR U5103 ( .A(n4973), .B(n4974), .Z(n4975) );
  XOR U5104 ( .A(n4976), .B(n4975), .Z(n4823) );
  XNOR U5105 ( .A(n4822), .B(n4823), .Z(n4825) );
  NANDN U5106 ( .A(n4684), .B(n4683), .Z(n4688) );
  OR U5107 ( .A(n4686), .B(n4685), .Z(n4687) );
  AND U5108 ( .A(n4688), .B(n4687), .Z(n4879) );
  NANDN U5109 ( .A(n4690), .B(n4689), .Z(n4694) );
  NANDN U5110 ( .A(n4692), .B(n4691), .Z(n4693) );
  NAND U5111 ( .A(n4694), .B(n4693), .Z(n4878) );
  XNOR U5112 ( .A(n4879), .B(n4878), .Z(n4881) );
  NANDN U5113 ( .A(n32483), .B(n4695), .Z(n4697) );
  XOR U5114 ( .A(b[19]), .B(a[26]), .Z(n4918) );
  NANDN U5115 ( .A(n32823), .B(n4918), .Z(n4696) );
  AND U5116 ( .A(n4697), .B(n4696), .Z(n4958) );
  NANDN U5117 ( .A(n31536), .B(n4698), .Z(n4700) );
  XOR U5118 ( .A(b[15]), .B(a[30]), .Z(n4930) );
  NANDN U5119 ( .A(n31925), .B(n4930), .Z(n4699) );
  AND U5120 ( .A(n4700), .B(n4699), .Z(n4956) );
  NANDN U5121 ( .A(n32013), .B(n4701), .Z(n4703) );
  XOR U5122 ( .A(b[17]), .B(a[28]), .Z(n4924) );
  NANDN U5123 ( .A(n32292), .B(n4924), .Z(n4702) );
  NAND U5124 ( .A(n4703), .B(n4702), .Z(n4955) );
  XNOR U5125 ( .A(n4956), .B(n4955), .Z(n4957) );
  XNOR U5126 ( .A(n4958), .B(n4957), .Z(n4968) );
  NAND U5127 ( .A(b[0]), .B(a[44]), .Z(n4704) );
  XNOR U5128 ( .A(b[1]), .B(n4704), .Z(n4706) );
  NANDN U5129 ( .A(b[0]), .B(a[43]), .Z(n4705) );
  NAND U5130 ( .A(n4706), .B(n4705), .Z(n4952) );
  XOR U5131 ( .A(b[43]), .B(b[44]), .Z(n37200) );
  IV U5132 ( .A(n37200), .Z(n37083) );
  ANDN U5133 ( .B(a[0]), .A(n37083), .Z(n4949) );
  NANDN U5134 ( .A(n36480), .B(n4707), .Z(n4709) );
  XOR U5135 ( .A(b[41]), .B(a[4]), .Z(n4942) );
  NANDN U5136 ( .A(n36594), .B(n4942), .Z(n4708) );
  AND U5137 ( .A(n4709), .B(n4708), .Z(n4950) );
  XOR U5138 ( .A(n4949), .B(n4950), .Z(n4951) );
  XOR U5139 ( .A(n4952), .B(n4951), .Z(n4967) );
  XOR U5140 ( .A(n4968), .B(n4967), .Z(n4970) );
  NANDN U5141 ( .A(n4711), .B(n4710), .Z(n4715) );
  OR U5142 ( .A(n4713), .B(n4712), .Z(n4714) );
  NAND U5143 ( .A(n4715), .B(n4714), .Z(n4969) );
  XOR U5144 ( .A(n4970), .B(n4969), .Z(n4880) );
  XOR U5145 ( .A(n4881), .B(n4880), .Z(n4824) );
  XOR U5146 ( .A(n4825), .B(n4824), .Z(n4986) );
  NANDN U5147 ( .A(n210), .B(n4716), .Z(n4718) );
  XOR U5148 ( .A(b[9]), .B(a[36]), .Z(n4936) );
  NANDN U5149 ( .A(n30267), .B(n4936), .Z(n4717) );
  AND U5150 ( .A(n4718), .B(n4717), .Z(n4908) );
  NANDN U5151 ( .A(n35936), .B(n4719), .Z(n4721) );
  XOR U5152 ( .A(b[37]), .B(a[8]), .Z(n4866) );
  NANDN U5153 ( .A(n36047), .B(n4866), .Z(n4720) );
  AND U5154 ( .A(n4721), .B(n4720), .Z(n4907) );
  NANDN U5155 ( .A(n33875), .B(n4722), .Z(n4724) );
  XOR U5156 ( .A(b[25]), .B(a[20]), .Z(n4945) );
  NANDN U5157 ( .A(n33994), .B(n4945), .Z(n4723) );
  NAND U5158 ( .A(n4724), .B(n4723), .Z(n4906) );
  XOR U5159 ( .A(n4907), .B(n4906), .Z(n4909) );
  XOR U5160 ( .A(n4908), .B(n4909), .Z(n4962) );
  NANDN U5161 ( .A(n35260), .B(n4725), .Z(n4727) );
  XOR U5162 ( .A(b[33]), .B(a[12]), .Z(n4927) );
  NANDN U5163 ( .A(n35456), .B(n4927), .Z(n4726) );
  AND U5164 ( .A(n4727), .B(n4726), .Z(n4836) );
  NANDN U5165 ( .A(n35611), .B(n4728), .Z(n4730) );
  XOR U5166 ( .A(b[35]), .B(a[10]), .Z(n4863) );
  NANDN U5167 ( .A(n35801), .B(n4863), .Z(n4729) );
  AND U5168 ( .A(n4730), .B(n4729), .Z(n4835) );
  NANDN U5169 ( .A(n30482), .B(n4731), .Z(n4733) );
  XOR U5170 ( .A(b[11]), .B(a[34]), .Z(n4933) );
  NANDN U5171 ( .A(n30891), .B(n4933), .Z(n4732) );
  NAND U5172 ( .A(n4733), .B(n4732), .Z(n4834) );
  XOR U5173 ( .A(n4835), .B(n4834), .Z(n4837) );
  XNOR U5174 ( .A(n4836), .B(n4837), .Z(n4961) );
  XNOR U5175 ( .A(n4962), .B(n4961), .Z(n4963) );
  NANDN U5176 ( .A(n4735), .B(n4734), .Z(n4739) );
  OR U5177 ( .A(n4737), .B(n4736), .Z(n4738) );
  NAND U5178 ( .A(n4739), .B(n4738), .Z(n4964) );
  XNOR U5179 ( .A(n4963), .B(n4964), .Z(n4828) );
  NANDN U5180 ( .A(n4741), .B(n4740), .Z(n4745) );
  NAND U5181 ( .A(n4743), .B(n4742), .Z(n4744) );
  NAND U5182 ( .A(n4745), .B(n4744), .Z(n4829) );
  XNOR U5183 ( .A(n4828), .B(n4829), .Z(n4830) );
  NANDN U5184 ( .A(n32996), .B(n4746), .Z(n4748) );
  XOR U5185 ( .A(b[21]), .B(a[24]), .Z(n4897) );
  NANDN U5186 ( .A(n33271), .B(n4897), .Z(n4747) );
  AND U5187 ( .A(n4748), .B(n4747), .Z(n4902) );
  NANDN U5188 ( .A(n34909), .B(n4749), .Z(n4751) );
  XOR U5189 ( .A(b[31]), .B(a[14]), .Z(n4939) );
  NANDN U5190 ( .A(n35145), .B(n4939), .Z(n4750) );
  AND U5191 ( .A(n4751), .B(n4750), .Z(n4901) );
  NANDN U5192 ( .A(n31055), .B(n4752), .Z(n4754) );
  XOR U5193 ( .A(b[13]), .B(a[32]), .Z(n4869) );
  NANDN U5194 ( .A(n31293), .B(n4869), .Z(n4753) );
  NAND U5195 ( .A(n4754), .B(n4753), .Z(n4900) );
  XOR U5196 ( .A(n4901), .B(n4900), .Z(n4903) );
  XOR U5197 ( .A(n4902), .B(n4903), .Z(n4873) );
  NANDN U5198 ( .A(n28889), .B(n4755), .Z(n4757) );
  XOR U5199 ( .A(b[5]), .B(a[40]), .Z(n4894) );
  NANDN U5200 ( .A(n29138), .B(n4894), .Z(n4756) );
  AND U5201 ( .A(n4757), .B(n4756), .Z(n4846) );
  XOR U5202 ( .A(b[42]), .B(b[43]), .Z(n4758) );
  ANDN U5203 ( .B(n4758), .A(n36963), .Z(n36962) );
  IV U5204 ( .A(n36962), .Z(n36742) );
  NANDN U5205 ( .A(n36742), .B(n4759), .Z(n4761) );
  XOR U5206 ( .A(b[43]), .B(a[2]), .Z(n4850) );
  NANDN U5207 ( .A(n36891), .B(n4850), .Z(n4760) );
  AND U5208 ( .A(n4761), .B(n4760), .Z(n4845) );
  NANDN U5209 ( .A(n34223), .B(n4762), .Z(n4764) );
  XOR U5210 ( .A(b[27]), .B(a[18]), .Z(n4888) );
  NANDN U5211 ( .A(n34458), .B(n4888), .Z(n4763) );
  NAND U5212 ( .A(n4764), .B(n4763), .Z(n4844) );
  XOR U5213 ( .A(n4845), .B(n4844), .Z(n4847) );
  XNOR U5214 ( .A(n4846), .B(n4847), .Z(n4872) );
  XNOR U5215 ( .A(n4873), .B(n4872), .Z(n4874) );
  NANDN U5216 ( .A(n4766), .B(n4765), .Z(n4770) );
  OR U5217 ( .A(n4768), .B(n4767), .Z(n4769) );
  NAND U5218 ( .A(n4770), .B(n4769), .Z(n4875) );
  XOR U5219 ( .A(n4874), .B(n4875), .Z(n4831) );
  XNOR U5220 ( .A(n4830), .B(n4831), .Z(n4981) );
  NANDN U5221 ( .A(n4772), .B(n4771), .Z(n4776) );
  NAND U5222 ( .A(n4774), .B(n4773), .Z(n4775) );
  AND U5223 ( .A(n4776), .B(n4775), .Z(n4980) );
  NANDN U5224 ( .A(n4778), .B(n4777), .Z(n4782) );
  NAND U5225 ( .A(n4780), .B(n4779), .Z(n4781) );
  NAND U5226 ( .A(n4782), .B(n4781), .Z(n4979) );
  XOR U5227 ( .A(n4980), .B(n4979), .Z(n4982) );
  XNOR U5228 ( .A(n4981), .B(n4982), .Z(n4985) );
  XNOR U5229 ( .A(n4986), .B(n4985), .Z(n4987) );
  NANDN U5230 ( .A(n4784), .B(n4783), .Z(n4788) );
  NAND U5231 ( .A(n4786), .B(n4785), .Z(n4787) );
  NAND U5232 ( .A(n4788), .B(n4787), .Z(n4988) );
  XNOR U5233 ( .A(n4987), .B(n4988), .Z(n4999) );
  XOR U5234 ( .A(n5000), .B(n4999), .Z(n4819) );
  NAND U5235 ( .A(n4790), .B(n4789), .Z(n4794) );
  NAND U5236 ( .A(n4792), .B(n4791), .Z(n4793) );
  AND U5237 ( .A(n4794), .B(n4793), .Z(n4817) );
  NANDN U5238 ( .A(n4796), .B(n4795), .Z(n4800) );
  NAND U5239 ( .A(n4798), .B(n4797), .Z(n4799) );
  AND U5240 ( .A(n4800), .B(n4799), .Z(n4816) );
  XNOR U5241 ( .A(n4817), .B(n4816), .Z(n4818) );
  XOR U5242 ( .A(n4819), .B(n4818), .Z(n5004) );
  XNOR U5243 ( .A(n5003), .B(n5004), .Z(n5005) );
  XOR U5244 ( .A(n5006), .B(n5005), .Z(n4811) );
  NANDN U5245 ( .A(n4802), .B(n4801), .Z(n4806) );
  OR U5246 ( .A(n4804), .B(n4803), .Z(n4805) );
  AND U5247 ( .A(n4806), .B(n4805), .Z(n4810) );
  XNOR U5248 ( .A(n4811), .B(n4810), .Z(n4812) );
  XNOR U5249 ( .A(n4813), .B(n4812), .Z(n4809) );
  XNOR U5250 ( .A(sreg[108]), .B(n4809), .Z(n4807) );
  XOR U5251 ( .A(n4808), .B(n4807), .Z(c[108]) );
  NANDN U5252 ( .A(n4811), .B(n4810), .Z(n4815) );
  NANDN U5253 ( .A(n4813), .B(n4812), .Z(n4814) );
  AND U5254 ( .A(n4815), .B(n4814), .Z(n5017) );
  NANDN U5255 ( .A(n4817), .B(n4816), .Z(n4821) );
  NANDN U5256 ( .A(n4819), .B(n4818), .Z(n4820) );
  AND U5257 ( .A(n4821), .B(n4820), .Z(n5212) );
  NANDN U5258 ( .A(n4823), .B(n4822), .Z(n4827) );
  NAND U5259 ( .A(n4825), .B(n4824), .Z(n4826) );
  AND U5260 ( .A(n4827), .B(n4826), .Z(n5035) );
  NANDN U5261 ( .A(n4829), .B(n4828), .Z(n4833) );
  NANDN U5262 ( .A(n4831), .B(n4830), .Z(n4832) );
  AND U5263 ( .A(n4833), .B(n4832), .Z(n5033) );
  NANDN U5264 ( .A(n4835), .B(n4834), .Z(n4839) );
  OR U5265 ( .A(n4837), .B(n4836), .Z(n4838) );
  AND U5266 ( .A(n4839), .B(n4838), .Z(n5051) );
  XNOR U5267 ( .A(n5051), .B(n5050), .Z(n5053) );
  NANDN U5268 ( .A(n4845), .B(n4844), .Z(n4849) );
  OR U5269 ( .A(n4847), .B(n4846), .Z(n4848) );
  AND U5270 ( .A(n4849), .B(n4848), .Z(n5191) );
  NANDN U5271 ( .A(n36742), .B(n4850), .Z(n4852) );
  XOR U5272 ( .A(b[43]), .B(a[3]), .Z(n5095) );
  NANDN U5273 ( .A(n36891), .B(n5095), .Z(n4851) );
  AND U5274 ( .A(n4852), .B(n4851), .Z(n5134) );
  XOR U5275 ( .A(b[45]), .B(b[44]), .Z(n5136) );
  XOR U5276 ( .A(b[45]), .B(a[0]), .Z(n4853) );
  NAND U5277 ( .A(n5136), .B(n4853), .Z(n4854) );
  OR U5278 ( .A(n4854), .B(n37200), .Z(n4856) );
  XNOR U5279 ( .A(b[45]), .B(a[1]), .Z(n5137) );
  NANDN U5280 ( .A(n5137), .B(n37200), .Z(n4855) );
  NAND U5281 ( .A(n4856), .B(n4855), .Z(n5135) );
  XOR U5282 ( .A(n5134), .B(n5135), .Z(n5154) );
  NAND U5283 ( .A(b[0]), .B(a[45]), .Z(n4857) );
  XNOR U5284 ( .A(b[1]), .B(n4857), .Z(n4859) );
  NANDN U5285 ( .A(b[0]), .B(a[44]), .Z(n4858) );
  NAND U5286 ( .A(n4859), .B(n4858), .Z(n5153) );
  NAND U5287 ( .A(n33492), .B(n4860), .Z(n4862) );
  XNOR U5288 ( .A(b[23]), .B(a[23]), .Z(n5179) );
  NANDN U5289 ( .A(n5179), .B(n33868), .Z(n4861) );
  AND U5290 ( .A(n4862), .B(n4861), .Z(n5152) );
  XOR U5291 ( .A(n5153), .B(n5152), .Z(n5155) );
  XNOR U5292 ( .A(n5154), .B(n5155), .Z(n5188) );
  NANDN U5293 ( .A(n35611), .B(n4863), .Z(n4865) );
  XOR U5294 ( .A(b[35]), .B(a[11]), .Z(n5164) );
  NANDN U5295 ( .A(n35801), .B(n5164), .Z(n4864) );
  AND U5296 ( .A(n4865), .B(n4864), .Z(n5185) );
  NANDN U5297 ( .A(n35936), .B(n4866), .Z(n4868) );
  XOR U5298 ( .A(b[37]), .B(a[9]), .Z(n5167) );
  NANDN U5299 ( .A(n36047), .B(n5167), .Z(n4867) );
  AND U5300 ( .A(n4868), .B(n4867), .Z(n5183) );
  NANDN U5301 ( .A(n31055), .B(n4869), .Z(n4871) );
  XOR U5302 ( .A(b[13]), .B(a[33]), .Z(n5062) );
  NANDN U5303 ( .A(n31293), .B(n5062), .Z(n4870) );
  NAND U5304 ( .A(n4871), .B(n4870), .Z(n5182) );
  XNOR U5305 ( .A(n5183), .B(n5182), .Z(n5184) );
  XNOR U5306 ( .A(n5185), .B(n5184), .Z(n5189) );
  XOR U5307 ( .A(n5188), .B(n5189), .Z(n5190) );
  XNOR U5308 ( .A(n5191), .B(n5190), .Z(n5052) );
  XOR U5309 ( .A(n5053), .B(n5052), .Z(n5045) );
  NANDN U5310 ( .A(n4873), .B(n4872), .Z(n4877) );
  NANDN U5311 ( .A(n4875), .B(n4874), .Z(n4876) );
  NAND U5312 ( .A(n4877), .B(n4876), .Z(n5044) );
  XNOR U5313 ( .A(n5045), .B(n5044), .Z(n5046) );
  XNOR U5314 ( .A(n5046), .B(n5047), .Z(n5032) );
  XNOR U5315 ( .A(n5033), .B(n5032), .Z(n5034) );
  XOR U5316 ( .A(n5035), .B(n5034), .Z(n5206) );
  NANDN U5317 ( .A(n209), .B(n4882), .Z(n4884) );
  XOR U5318 ( .A(b[3]), .B(a[43]), .Z(n5173) );
  NANDN U5319 ( .A(n28941), .B(n5173), .Z(n4883) );
  AND U5320 ( .A(n4884), .B(n4883), .Z(n5079) );
  NANDN U5321 ( .A(n36210), .B(n4885), .Z(n4887) );
  XOR U5322 ( .A(b[39]), .B(a[7]), .Z(n5143) );
  NANDN U5323 ( .A(n36347), .B(n5143), .Z(n4886) );
  AND U5324 ( .A(n4887), .B(n4886), .Z(n5078) );
  NANDN U5325 ( .A(n34223), .B(n4888), .Z(n4890) );
  XOR U5326 ( .A(b[27]), .B(a[19]), .Z(n5149) );
  NANDN U5327 ( .A(n34458), .B(n5149), .Z(n4889) );
  NAND U5328 ( .A(n4890), .B(n4889), .Z(n5077) );
  XOR U5329 ( .A(n5078), .B(n5077), .Z(n5080) );
  XOR U5330 ( .A(n5079), .B(n5080), .Z(n5123) );
  NANDN U5331 ( .A(n29499), .B(n4891), .Z(n4893) );
  XOR U5332 ( .A(b[7]), .B(a[39]), .Z(n5104) );
  NANDN U5333 ( .A(n29735), .B(n5104), .Z(n4892) );
  AND U5334 ( .A(n4893), .B(n4892), .Z(n5160) );
  NANDN U5335 ( .A(n28889), .B(n4894), .Z(n4896) );
  XOR U5336 ( .A(b[5]), .B(a[41]), .Z(n5146) );
  NANDN U5337 ( .A(n29138), .B(n5146), .Z(n4895) );
  AND U5338 ( .A(n4896), .B(n4895), .Z(n5159) );
  NANDN U5339 ( .A(n32996), .B(n4897), .Z(n4899) );
  XOR U5340 ( .A(b[21]), .B(a[25]), .Z(n5074) );
  NANDN U5341 ( .A(n33271), .B(n5074), .Z(n4898) );
  NAND U5342 ( .A(n4899), .B(n4898), .Z(n5158) );
  XOR U5343 ( .A(n5159), .B(n5158), .Z(n5161) );
  XNOR U5344 ( .A(n5160), .B(n5161), .Z(n5122) );
  XNOR U5345 ( .A(n5123), .B(n5122), .Z(n5125) );
  NANDN U5346 ( .A(n4901), .B(n4900), .Z(n4905) );
  OR U5347 ( .A(n4903), .B(n4902), .Z(n4904) );
  AND U5348 ( .A(n4905), .B(n4904), .Z(n5124) );
  XOR U5349 ( .A(n5125), .B(n5124), .Z(n5195) );
  NANDN U5350 ( .A(n4907), .B(n4906), .Z(n4911) );
  OR U5351 ( .A(n4909), .B(n4908), .Z(n4910) );
  AND U5352 ( .A(n4911), .B(n4910), .Z(n5193) );
  NANDN U5353 ( .A(n4913), .B(n4912), .Z(n4917) );
  NANDN U5354 ( .A(n4915), .B(n4914), .Z(n4916) );
  NAND U5355 ( .A(n4917), .B(n4916), .Z(n5192) );
  XNOR U5356 ( .A(n5193), .B(n5192), .Z(n5194) );
  XNOR U5357 ( .A(n5195), .B(n5194), .Z(n5038) );
  NANDN U5358 ( .A(n32483), .B(n4918), .Z(n4920) );
  XOR U5359 ( .A(b[19]), .B(a[27]), .Z(n5071) );
  NANDN U5360 ( .A(n32823), .B(n5071), .Z(n4919) );
  AND U5361 ( .A(n4920), .B(n4919), .Z(n5112) );
  NANDN U5362 ( .A(n34634), .B(n4921), .Z(n4923) );
  XOR U5363 ( .A(b[29]), .B(a[17]), .Z(n5107) );
  NANDN U5364 ( .A(n34722), .B(n5107), .Z(n4922) );
  AND U5365 ( .A(n4923), .B(n4922), .Z(n5111) );
  NANDN U5366 ( .A(n32013), .B(n4924), .Z(n4926) );
  XOR U5367 ( .A(b[17]), .B(a[29]), .Z(n5065) );
  NANDN U5368 ( .A(n32292), .B(n5065), .Z(n4925) );
  AND U5369 ( .A(n4926), .B(n4925), .Z(n5131) );
  NANDN U5370 ( .A(n35260), .B(n4927), .Z(n4929) );
  XOR U5371 ( .A(b[33]), .B(a[13]), .Z(n5059) );
  NANDN U5372 ( .A(n35456), .B(n5059), .Z(n4928) );
  AND U5373 ( .A(n4929), .B(n4928), .Z(n5129) );
  NANDN U5374 ( .A(n31536), .B(n4930), .Z(n4932) );
  XOR U5375 ( .A(b[15]), .B(a[31]), .Z(n5068) );
  NANDN U5376 ( .A(n31925), .B(n5068), .Z(n4931) );
  NAND U5377 ( .A(n4932), .B(n4931), .Z(n5128) );
  XNOR U5378 ( .A(n5129), .B(n5128), .Z(n5130) );
  XNOR U5379 ( .A(n5131), .B(n5130), .Z(n5110) );
  XOR U5380 ( .A(n5111), .B(n5110), .Z(n5113) );
  XOR U5381 ( .A(n5112), .B(n5113), .Z(n5118) );
  NANDN U5382 ( .A(n30482), .B(n4933), .Z(n4935) );
  XOR U5383 ( .A(b[11]), .B(a[35]), .Z(n5170) );
  NANDN U5384 ( .A(n30891), .B(n5170), .Z(n4934) );
  AND U5385 ( .A(n4935), .B(n4934), .Z(n5091) );
  NANDN U5386 ( .A(n210), .B(n4936), .Z(n4938) );
  XOR U5387 ( .A(b[9]), .B(a[37]), .Z(n5101) );
  NANDN U5388 ( .A(n30267), .B(n5101), .Z(n4937) );
  AND U5389 ( .A(n4938), .B(n4937), .Z(n5090) );
  NANDN U5390 ( .A(n34909), .B(n4939), .Z(n4941) );
  XOR U5391 ( .A(b[31]), .B(a[15]), .Z(n5056) );
  NANDN U5392 ( .A(n35145), .B(n5056), .Z(n4940) );
  NAND U5393 ( .A(n4941), .B(n4940), .Z(n5089) );
  XOR U5394 ( .A(n5090), .B(n5089), .Z(n5092) );
  XOR U5395 ( .A(n5091), .B(n5092), .Z(n5117) );
  NANDN U5396 ( .A(n36480), .B(n4942), .Z(n4944) );
  XOR U5397 ( .A(b[41]), .B(a[5]), .Z(n5176) );
  NANDN U5398 ( .A(n36594), .B(n5176), .Z(n4943) );
  AND U5399 ( .A(n4944), .B(n4943), .Z(n5085) );
  NANDN U5400 ( .A(n33875), .B(n4945), .Z(n4947) );
  XOR U5401 ( .A(b[25]), .B(a[21]), .Z(n5140) );
  NANDN U5402 ( .A(n33994), .B(n5140), .Z(n4946) );
  AND U5403 ( .A(n4947), .B(n4946), .Z(n5084) );
  NAND U5404 ( .A(b[43]), .B(b[44]), .Z(n4948) );
  AND U5405 ( .A(b[45]), .B(n4948), .Z(n37336) );
  ANDN U5406 ( .B(n37336), .A(n4949), .Z(n5083) );
  XOR U5407 ( .A(n5084), .B(n5083), .Z(n5086) );
  XNOR U5408 ( .A(n5085), .B(n5086), .Z(n5116) );
  XOR U5409 ( .A(n5117), .B(n5116), .Z(n5119) );
  XOR U5410 ( .A(n5118), .B(n5119), .Z(n5201) );
  NANDN U5411 ( .A(n4950), .B(n4949), .Z(n4954) );
  OR U5412 ( .A(n4952), .B(n4951), .Z(n4953) );
  AND U5413 ( .A(n4954), .B(n4953), .Z(n5199) );
  NANDN U5414 ( .A(n4956), .B(n4955), .Z(n4960) );
  NANDN U5415 ( .A(n4958), .B(n4957), .Z(n4959) );
  NAND U5416 ( .A(n4960), .B(n4959), .Z(n5198) );
  XNOR U5417 ( .A(n5199), .B(n5198), .Z(n5200) );
  XOR U5418 ( .A(n5201), .B(n5200), .Z(n5039) );
  XNOR U5419 ( .A(n5038), .B(n5039), .Z(n5041) );
  NANDN U5420 ( .A(n4962), .B(n4961), .Z(n4966) );
  NANDN U5421 ( .A(n4964), .B(n4963), .Z(n4965) );
  AND U5422 ( .A(n4966), .B(n4965), .Z(n5040) );
  XOR U5423 ( .A(n5041), .B(n5040), .Z(n5028) );
  NAND U5424 ( .A(n4968), .B(n4967), .Z(n4972) );
  NAND U5425 ( .A(n4970), .B(n4969), .Z(n4971) );
  AND U5426 ( .A(n4972), .B(n4971), .Z(n5026) );
  NANDN U5427 ( .A(n4974), .B(n4973), .Z(n4978) );
  NANDN U5428 ( .A(n4976), .B(n4975), .Z(n4977) );
  NAND U5429 ( .A(n4978), .B(n4977), .Z(n5027) );
  XOR U5430 ( .A(n5026), .B(n5027), .Z(n5029) );
  XOR U5431 ( .A(n5028), .B(n5029), .Z(n5205) );
  NANDN U5432 ( .A(n4980), .B(n4979), .Z(n4984) );
  NANDN U5433 ( .A(n4982), .B(n4981), .Z(n4983) );
  AND U5434 ( .A(n4984), .B(n4983), .Z(n5204) );
  XOR U5435 ( .A(n5205), .B(n5204), .Z(n5207) );
  XOR U5436 ( .A(n5206), .B(n5207), .Z(n5022) );
  NANDN U5437 ( .A(n4986), .B(n4985), .Z(n4990) );
  NANDN U5438 ( .A(n4988), .B(n4987), .Z(n4989) );
  AND U5439 ( .A(n4990), .B(n4989), .Z(n5021) );
  NANDN U5440 ( .A(n4992), .B(n4991), .Z(n4996) );
  OR U5441 ( .A(n4994), .B(n4993), .Z(n4995) );
  AND U5442 ( .A(n4996), .B(n4995), .Z(n5020) );
  XOR U5443 ( .A(n5021), .B(n5020), .Z(n5023) );
  XOR U5444 ( .A(n5022), .B(n5023), .Z(n5211) );
  NANDN U5445 ( .A(n4998), .B(n4997), .Z(n5002) );
  NAND U5446 ( .A(n5000), .B(n4999), .Z(n5001) );
  AND U5447 ( .A(n5002), .B(n5001), .Z(n5210) );
  XOR U5448 ( .A(n5211), .B(n5210), .Z(n5213) );
  XOR U5449 ( .A(n5212), .B(n5213), .Z(n5015) );
  NANDN U5450 ( .A(n5004), .B(n5003), .Z(n5008) );
  NAND U5451 ( .A(n5006), .B(n5005), .Z(n5007) );
  AND U5452 ( .A(n5008), .B(n5007), .Z(n5014) );
  XNOR U5453 ( .A(n5015), .B(n5014), .Z(n5016) );
  XNOR U5454 ( .A(n5017), .B(n5016), .Z(n5009) );
  XNOR U5455 ( .A(sreg[109]), .B(n5009), .Z(n5010) );
  XNOR U5456 ( .A(n5011), .B(n5010), .Z(c[109]) );
  NANDN U5457 ( .A(sreg[109]), .B(n5009), .Z(n5013) );
  NAND U5458 ( .A(n5011), .B(n5010), .Z(n5012) );
  NAND U5459 ( .A(n5013), .B(n5012), .Z(n5216) );
  XNOR U5460 ( .A(sreg[110]), .B(n5216), .Z(n5218) );
  NANDN U5461 ( .A(n5015), .B(n5014), .Z(n5019) );
  NANDN U5462 ( .A(n5017), .B(n5016), .Z(n5018) );
  AND U5463 ( .A(n5019), .B(n5018), .Z(n5224) );
  NANDN U5464 ( .A(n5021), .B(n5020), .Z(n5025) );
  OR U5465 ( .A(n5023), .B(n5022), .Z(n5024) );
  AND U5466 ( .A(n5025), .B(n5024), .Z(n5430) );
  NANDN U5467 ( .A(n5027), .B(n5026), .Z(n5031) );
  OR U5468 ( .A(n5029), .B(n5028), .Z(n5030) );
  AND U5469 ( .A(n5031), .B(n5030), .Z(n5227) );
  NANDN U5470 ( .A(n5033), .B(n5032), .Z(n5037) );
  NAND U5471 ( .A(n5035), .B(n5034), .Z(n5036) );
  NAND U5472 ( .A(n5037), .B(n5036), .Z(n5228) );
  XNOR U5473 ( .A(n5227), .B(n5228), .Z(n5230) );
  NANDN U5474 ( .A(n5039), .B(n5038), .Z(n5043) );
  NAND U5475 ( .A(n5041), .B(n5040), .Z(n5042) );
  AND U5476 ( .A(n5043), .B(n5042), .Z(n5234) );
  NANDN U5477 ( .A(n5045), .B(n5044), .Z(n5049) );
  NANDN U5478 ( .A(n5047), .B(n5046), .Z(n5048) );
  AND U5479 ( .A(n5049), .B(n5048), .Z(n5233) );
  XNOR U5480 ( .A(n5234), .B(n5233), .Z(n5235) );
  NANDN U5481 ( .A(n5051), .B(n5050), .Z(n5055) );
  NAND U5482 ( .A(n5053), .B(n5052), .Z(n5054) );
  AND U5483 ( .A(n5055), .B(n5054), .Z(n5246) );
  NANDN U5484 ( .A(n34909), .B(n5056), .Z(n5058) );
  XOR U5485 ( .A(b[31]), .B(a[16]), .Z(n5317) );
  NANDN U5486 ( .A(n35145), .B(n5317), .Z(n5057) );
  AND U5487 ( .A(n5058), .B(n5057), .Z(n5293) );
  NANDN U5488 ( .A(n35260), .B(n5059), .Z(n5061) );
  XOR U5489 ( .A(b[33]), .B(a[14]), .Z(n5382) );
  NANDN U5490 ( .A(n35456), .B(n5382), .Z(n5060) );
  AND U5491 ( .A(n5061), .B(n5060), .Z(n5292) );
  NANDN U5492 ( .A(n31055), .B(n5062), .Z(n5064) );
  XOR U5493 ( .A(b[13]), .B(a[34]), .Z(n5352) );
  NANDN U5494 ( .A(n31293), .B(n5352), .Z(n5063) );
  NAND U5495 ( .A(n5064), .B(n5063), .Z(n5291) );
  XOR U5496 ( .A(n5292), .B(n5291), .Z(n5294) );
  XOR U5497 ( .A(n5293), .B(n5294), .Z(n5405) );
  NANDN U5498 ( .A(n32013), .B(n5065), .Z(n5067) );
  XOR U5499 ( .A(b[17]), .B(a[30]), .Z(n5288) );
  NANDN U5500 ( .A(n32292), .B(n5288), .Z(n5066) );
  AND U5501 ( .A(n5067), .B(n5066), .Z(n5310) );
  NANDN U5502 ( .A(n31536), .B(n5068), .Z(n5070) );
  XOR U5503 ( .A(b[15]), .B(a[32]), .Z(n5373) );
  NANDN U5504 ( .A(n31925), .B(n5373), .Z(n5069) );
  AND U5505 ( .A(n5070), .B(n5069), .Z(n5309) );
  NANDN U5506 ( .A(n32483), .B(n5071), .Z(n5073) );
  XOR U5507 ( .A(b[19]), .B(a[28]), .Z(n5285) );
  NANDN U5508 ( .A(n32823), .B(n5285), .Z(n5072) );
  NAND U5509 ( .A(n5073), .B(n5072), .Z(n5308) );
  XOR U5510 ( .A(n5309), .B(n5308), .Z(n5311) );
  XOR U5511 ( .A(n5310), .B(n5311), .Z(n5404) );
  NAND U5512 ( .A(n33413), .B(n5074), .Z(n5076) );
  XNOR U5513 ( .A(b[21]), .B(a[26]), .Z(n5282) );
  NANDN U5514 ( .A(n5282), .B(n33414), .Z(n5075) );
  AND U5515 ( .A(n5076), .B(n5075), .Z(n5403) );
  XOR U5516 ( .A(n5404), .B(n5403), .Z(n5406) );
  XOR U5517 ( .A(n5405), .B(n5406), .Z(n5411) );
  NANDN U5518 ( .A(n5078), .B(n5077), .Z(n5082) );
  OR U5519 ( .A(n5080), .B(n5079), .Z(n5081) );
  AND U5520 ( .A(n5082), .B(n5081), .Z(n5410) );
  NANDN U5521 ( .A(n5084), .B(n5083), .Z(n5088) );
  OR U5522 ( .A(n5086), .B(n5085), .Z(n5087) );
  NAND U5523 ( .A(n5088), .B(n5087), .Z(n5409) );
  XOR U5524 ( .A(n5410), .B(n5409), .Z(n5412) );
  XOR U5525 ( .A(n5411), .B(n5412), .Z(n5417) );
  NANDN U5526 ( .A(n5090), .B(n5089), .Z(n5094) );
  OR U5527 ( .A(n5092), .B(n5091), .Z(n5093) );
  AND U5528 ( .A(n5094), .B(n5093), .Z(n5265) );
  XOR U5529 ( .A(b[45]), .B(b[46]), .Z(n37341) );
  IV U5530 ( .A(n37341), .Z(n37172) );
  ANDN U5531 ( .B(a[0]), .A(n37172), .Z(n5321) );
  NANDN U5532 ( .A(n36742), .B(n5095), .Z(n5097) );
  XOR U5533 ( .A(b[43]), .B(a[4]), .Z(n5376) );
  NANDN U5534 ( .A(n36891), .B(n5376), .Z(n5096) );
  AND U5535 ( .A(n5097), .B(n5096), .Z(n5303) );
  XNOR U5536 ( .A(n5321), .B(n5303), .Z(n5304) );
  NAND U5537 ( .A(b[0]), .B(a[46]), .Z(n5098) );
  XNOR U5538 ( .A(b[1]), .B(n5098), .Z(n5100) );
  NANDN U5539 ( .A(b[0]), .B(a[45]), .Z(n5099) );
  NAND U5540 ( .A(n5100), .B(n5099), .Z(n5305) );
  XOR U5541 ( .A(n5304), .B(n5305), .Z(n5264) );
  NANDN U5542 ( .A(n210), .B(n5101), .Z(n5103) );
  XOR U5543 ( .A(b[9]), .B(a[38]), .Z(n5379) );
  NANDN U5544 ( .A(n30267), .B(n5379), .Z(n5102) );
  AND U5545 ( .A(n5103), .B(n5102), .Z(n5334) );
  NANDN U5546 ( .A(n29499), .B(n5104), .Z(n5106) );
  XOR U5547 ( .A(b[7]), .B(a[40]), .Z(n5314) );
  NANDN U5548 ( .A(n29735), .B(n5314), .Z(n5105) );
  AND U5549 ( .A(n5106), .B(n5105), .Z(n5332) );
  NANDN U5550 ( .A(n34634), .B(n5107), .Z(n5109) );
  XOR U5551 ( .A(b[29]), .B(a[18]), .Z(n5328) );
  NANDN U5552 ( .A(n34722), .B(n5328), .Z(n5108) );
  NAND U5553 ( .A(n5109), .B(n5108), .Z(n5331) );
  XNOR U5554 ( .A(n5332), .B(n5331), .Z(n5333) );
  XOR U5555 ( .A(n5334), .B(n5333), .Z(n5263) );
  XNOR U5556 ( .A(n5264), .B(n5263), .Z(n5266) );
  NANDN U5557 ( .A(n5111), .B(n5110), .Z(n5115) );
  OR U5558 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U5559 ( .A(n5115), .B(n5114), .Z(n5416) );
  XOR U5560 ( .A(n5415), .B(n5416), .Z(n5418) );
  XOR U5561 ( .A(n5417), .B(n5418), .Z(n5254) );
  NANDN U5562 ( .A(n5117), .B(n5116), .Z(n5121) );
  OR U5563 ( .A(n5119), .B(n5118), .Z(n5120) );
  AND U5564 ( .A(n5121), .B(n5120), .Z(n5251) );
  NANDN U5565 ( .A(n5123), .B(n5122), .Z(n5127) );
  NAND U5566 ( .A(n5125), .B(n5124), .Z(n5126) );
  NAND U5567 ( .A(n5127), .B(n5126), .Z(n5252) );
  XNOR U5568 ( .A(n5251), .B(n5252), .Z(n5253) );
  XNOR U5569 ( .A(n5254), .B(n5253), .Z(n5245) );
  XNOR U5570 ( .A(n5246), .B(n5245), .Z(n5247) );
  NANDN U5571 ( .A(n5129), .B(n5128), .Z(n5133) );
  NANDN U5572 ( .A(n5131), .B(n5130), .Z(n5132) );
  AND U5573 ( .A(n5133), .B(n5132), .Z(n5358) );
  ANDN U5574 ( .B(n5135), .A(n5134), .Z(n5400) );
  ANDN U5575 ( .B(n5136), .A(n37200), .Z(n37202) );
  NANDN U5576 ( .A(n5137), .B(n37202), .Z(n5139) );
  XNOR U5577 ( .A(b[45]), .B(a[2]), .Z(n5275) );
  NANDN U5578 ( .A(n5275), .B(n37200), .Z(n5138) );
  AND U5579 ( .A(n5139), .B(n5138), .Z(n5398) );
  NAND U5580 ( .A(n34297), .B(n5140), .Z(n5142) );
  XNOR U5581 ( .A(b[25]), .B(a[22]), .Z(n5272) );
  NANDN U5582 ( .A(n5272), .B(n34298), .Z(n5141) );
  AND U5583 ( .A(n5142), .B(n5141), .Z(n5397) );
  XOR U5584 ( .A(n5398), .B(n5397), .Z(n5399) );
  NANDN U5585 ( .A(n36210), .B(n5143), .Z(n5145) );
  XOR U5586 ( .A(b[39]), .B(a[8]), .Z(n5349) );
  NANDN U5587 ( .A(n36347), .B(n5349), .Z(n5144) );
  AND U5588 ( .A(n5145), .B(n5144), .Z(n5300) );
  NANDN U5589 ( .A(n28889), .B(n5146), .Z(n5148) );
  XOR U5590 ( .A(b[5]), .B(a[42]), .Z(n5337) );
  NANDN U5591 ( .A(n29138), .B(n5337), .Z(n5147) );
  AND U5592 ( .A(n5148), .B(n5147), .Z(n5298) );
  NANDN U5593 ( .A(n34223), .B(n5149), .Z(n5151) );
  XOR U5594 ( .A(b[27]), .B(a[20]), .Z(n5343) );
  NANDN U5595 ( .A(n34458), .B(n5343), .Z(n5150) );
  NAND U5596 ( .A(n5151), .B(n5150), .Z(n5297) );
  XNOR U5597 ( .A(n5298), .B(n5297), .Z(n5299) );
  XNOR U5598 ( .A(n5300), .B(n5299), .Z(n5355) );
  XOR U5599 ( .A(n5356), .B(n5355), .Z(n5357) );
  XOR U5600 ( .A(n5358), .B(n5357), .Z(n5259) );
  NAND U5601 ( .A(n5153), .B(n5152), .Z(n5157) );
  NAND U5602 ( .A(n5155), .B(n5154), .Z(n5156) );
  NAND U5603 ( .A(n5157), .B(n5156), .Z(n5257) );
  NANDN U5604 ( .A(n5159), .B(n5158), .Z(n5163) );
  OR U5605 ( .A(n5161), .B(n5160), .Z(n5162) );
  AND U5606 ( .A(n5163), .B(n5162), .Z(n5258) );
  XOR U5607 ( .A(n5257), .B(n5258), .Z(n5260) );
  XOR U5608 ( .A(n5259), .B(n5260), .Z(n5424) );
  NAND U5609 ( .A(n35928), .B(n5164), .Z(n5166) );
  XNOR U5610 ( .A(b[35]), .B(a[12]), .Z(n5370) );
  NANDN U5611 ( .A(n5370), .B(n35929), .Z(n5165) );
  NAND U5612 ( .A(n5166), .B(n5165), .Z(n5387) );
  NAND U5613 ( .A(n36238), .B(n5167), .Z(n5169) );
  XNOR U5614 ( .A(b[37]), .B(a[10]), .Z(n5346) );
  NANDN U5615 ( .A(n5346), .B(n36239), .Z(n5168) );
  NAND U5616 ( .A(n5169), .B(n5168), .Z(n5386) );
  NAND U5617 ( .A(n31059), .B(n5170), .Z(n5172) );
  XNOR U5618 ( .A(b[11]), .B(a[36]), .Z(n5322) );
  NANDN U5619 ( .A(n5322), .B(n31060), .Z(n5171) );
  NAND U5620 ( .A(n5172), .B(n5171), .Z(n5385) );
  XNOR U5621 ( .A(n5386), .B(n5385), .Z(n5388) );
  NAND U5622 ( .A(n9942), .B(n5173), .Z(n5175) );
  XNOR U5623 ( .A(b[3]), .B(a[44]), .Z(n5340) );
  NANDN U5624 ( .A(n5340), .B(n9653), .Z(n5174) );
  NAND U5625 ( .A(n5175), .B(n5174), .Z(n5393) );
  NAND U5626 ( .A(n36735), .B(n5176), .Z(n5178) );
  XNOR U5627 ( .A(b[41]), .B(a[6]), .Z(n5325) );
  NANDN U5628 ( .A(n5325), .B(n36733), .Z(n5177) );
  NAND U5629 ( .A(n5178), .B(n5177), .Z(n5392) );
  NANDN U5630 ( .A(n5179), .B(n33492), .Z(n5181) );
  XNOR U5631 ( .A(b[23]), .B(a[24]), .Z(n5367) );
  NANDN U5632 ( .A(n5367), .B(n33868), .Z(n5180) );
  NAND U5633 ( .A(n5181), .B(n5180), .Z(n5391) );
  XNOR U5634 ( .A(n5392), .B(n5391), .Z(n5394) );
  XOR U5635 ( .A(n5393), .B(n5394), .Z(n5361) );
  XOR U5636 ( .A(n5362), .B(n5361), .Z(n5363) );
  NANDN U5637 ( .A(n5183), .B(n5182), .Z(n5187) );
  NANDN U5638 ( .A(n5185), .B(n5184), .Z(n5186) );
  NAND U5639 ( .A(n5187), .B(n5186), .Z(n5364) );
  XNOR U5640 ( .A(n5363), .B(n5364), .Z(n5421) );
  XNOR U5641 ( .A(n5421), .B(n5422), .Z(n5423) );
  XOR U5642 ( .A(n5424), .B(n5423), .Z(n5242) );
  NANDN U5643 ( .A(n5193), .B(n5192), .Z(n5197) );
  NANDN U5644 ( .A(n5195), .B(n5194), .Z(n5196) );
  AND U5645 ( .A(n5197), .B(n5196), .Z(n5240) );
  NANDN U5646 ( .A(n5199), .B(n5198), .Z(n5203) );
  NANDN U5647 ( .A(n5201), .B(n5200), .Z(n5202) );
  NAND U5648 ( .A(n5203), .B(n5202), .Z(n5239) );
  XNOR U5649 ( .A(n5240), .B(n5239), .Z(n5241) );
  XOR U5650 ( .A(n5242), .B(n5241), .Z(n5248) );
  XOR U5651 ( .A(n5247), .B(n5248), .Z(n5236) );
  XNOR U5652 ( .A(n5235), .B(n5236), .Z(n5229) );
  XOR U5653 ( .A(n5230), .B(n5229), .Z(n5428) );
  NANDN U5654 ( .A(n5205), .B(n5204), .Z(n5209) );
  OR U5655 ( .A(n5207), .B(n5206), .Z(n5208) );
  AND U5656 ( .A(n5209), .B(n5208), .Z(n5427) );
  XNOR U5657 ( .A(n5428), .B(n5427), .Z(n5429) );
  XNOR U5658 ( .A(n5430), .B(n5429), .Z(n5221) );
  NANDN U5659 ( .A(n5211), .B(n5210), .Z(n5215) );
  OR U5660 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U5661 ( .A(n5215), .B(n5214), .Z(n5222) );
  XNOR U5662 ( .A(n5221), .B(n5222), .Z(n5223) );
  XNOR U5663 ( .A(n5224), .B(n5223), .Z(n5217) );
  XNOR U5664 ( .A(n5218), .B(n5217), .Z(c[110]) );
  NANDN U5665 ( .A(sreg[110]), .B(n5216), .Z(n5220) );
  NAND U5666 ( .A(n5218), .B(n5217), .Z(n5219) );
  AND U5667 ( .A(n5220), .B(n5219), .Z(n5435) );
  NANDN U5668 ( .A(n5222), .B(n5221), .Z(n5226) );
  NANDN U5669 ( .A(n5224), .B(n5223), .Z(n5225) );
  AND U5670 ( .A(n5226), .B(n5225), .Z(n5440) );
  NANDN U5671 ( .A(n5228), .B(n5227), .Z(n5232) );
  NAND U5672 ( .A(n5230), .B(n5229), .Z(n5231) );
  AND U5673 ( .A(n5232), .B(n5231), .Z(n5641) );
  NANDN U5674 ( .A(n5234), .B(n5233), .Z(n5238) );
  NANDN U5675 ( .A(n5236), .B(n5235), .Z(n5237) );
  AND U5676 ( .A(n5238), .B(n5237), .Z(n5640) );
  NANDN U5677 ( .A(n5240), .B(n5239), .Z(n5244) );
  NANDN U5678 ( .A(n5242), .B(n5241), .Z(n5243) );
  AND U5679 ( .A(n5244), .B(n5243), .Z(n5634) );
  NANDN U5680 ( .A(n5246), .B(n5245), .Z(n5250) );
  NANDN U5681 ( .A(n5248), .B(n5247), .Z(n5249) );
  NAND U5682 ( .A(n5250), .B(n5249), .Z(n5633) );
  XNOR U5683 ( .A(n5634), .B(n5633), .Z(n5635) );
  NANDN U5684 ( .A(n5252), .B(n5251), .Z(n5256) );
  NANDN U5685 ( .A(n5254), .B(n5253), .Z(n5255) );
  AND U5686 ( .A(n5256), .B(n5255), .Z(n5618) );
  NAND U5687 ( .A(n5258), .B(n5257), .Z(n5262) );
  NAND U5688 ( .A(n5260), .B(n5259), .Z(n5261) );
  AND U5689 ( .A(n5262), .B(n5261), .Z(n5629) );
  NAND U5690 ( .A(n5264), .B(n5263), .Z(n5268) );
  NANDN U5691 ( .A(n5266), .B(n5265), .Z(n5267) );
  NAND U5692 ( .A(n5268), .B(n5267), .Z(n5630) );
  XNOR U5693 ( .A(n5629), .B(n5630), .Z(n5632) );
  NAND U5694 ( .A(b[0]), .B(a[47]), .Z(n5269) );
  XNOR U5695 ( .A(b[1]), .B(n5269), .Z(n5271) );
  NANDN U5696 ( .A(b[0]), .B(a[46]), .Z(n5270) );
  NAND U5697 ( .A(n5271), .B(n5270), .Z(n5473) );
  NANDN U5698 ( .A(n5272), .B(n34297), .Z(n5274) );
  XOR U5699 ( .A(b[25]), .B(a[23]), .Z(n5535) );
  NANDN U5700 ( .A(n33994), .B(n5535), .Z(n5273) );
  NAND U5701 ( .A(n5274), .B(n5273), .Z(n5472) );
  XNOR U5702 ( .A(n5473), .B(n5472), .Z(n5474) );
  NANDN U5703 ( .A(n5275), .B(n37202), .Z(n5277) );
  XOR U5704 ( .A(b[45]), .B(a[3]), .Z(n5569) );
  NANDN U5705 ( .A(n37083), .B(n5569), .Z(n5276) );
  AND U5706 ( .A(n5277), .B(n5276), .Z(n5520) );
  XOR U5707 ( .A(b[47]), .B(b[46]), .Z(n5531) );
  XOR U5708 ( .A(b[47]), .B(a[0]), .Z(n5278) );
  NAND U5709 ( .A(n5531), .B(n5278), .Z(n5279) );
  OR U5710 ( .A(n5279), .B(n37341), .Z(n5281) );
  XOR U5711 ( .A(b[47]), .B(a[1]), .Z(n5532) );
  NAND U5712 ( .A(n37341), .B(n5532), .Z(n5280) );
  NAND U5713 ( .A(n5281), .B(n5280), .Z(n5521) );
  XOR U5714 ( .A(n5520), .B(n5521), .Z(n5475) );
  XNOR U5715 ( .A(n5474), .B(n5475), .Z(n5582) );
  NANDN U5716 ( .A(n5282), .B(n33413), .Z(n5284) );
  XOR U5717 ( .A(b[21]), .B(a[27]), .Z(n5451) );
  NANDN U5718 ( .A(n33271), .B(n5451), .Z(n5283) );
  AND U5719 ( .A(n5284), .B(n5283), .Z(n5504) );
  NANDN U5720 ( .A(n32483), .B(n5285), .Z(n5287) );
  XOR U5721 ( .A(b[19]), .B(a[29]), .Z(n5448) );
  NANDN U5722 ( .A(n32823), .B(n5448), .Z(n5286) );
  AND U5723 ( .A(n5287), .B(n5286), .Z(n5503) );
  NANDN U5724 ( .A(n32013), .B(n5288), .Z(n5290) );
  XOR U5725 ( .A(b[17]), .B(a[31]), .Z(n5460) );
  NANDN U5726 ( .A(n32292), .B(n5460), .Z(n5289) );
  NAND U5727 ( .A(n5290), .B(n5289), .Z(n5502) );
  XOR U5728 ( .A(n5503), .B(n5502), .Z(n5505) );
  XOR U5729 ( .A(n5504), .B(n5505), .Z(n5581) );
  XOR U5730 ( .A(n5582), .B(n5581), .Z(n5584) );
  NANDN U5731 ( .A(n5292), .B(n5291), .Z(n5296) );
  OR U5732 ( .A(n5294), .B(n5293), .Z(n5295) );
  NAND U5733 ( .A(n5296), .B(n5295), .Z(n5583) );
  XOR U5734 ( .A(n5584), .B(n5583), .Z(n5596) );
  NANDN U5735 ( .A(n5298), .B(n5297), .Z(n5302) );
  NANDN U5736 ( .A(n5300), .B(n5299), .Z(n5301) );
  NAND U5737 ( .A(n5302), .B(n5301), .Z(n5594) );
  NANDN U5738 ( .A(n5303), .B(n5321), .Z(n5307) );
  NANDN U5739 ( .A(n5305), .B(n5304), .Z(n5306) );
  NAND U5740 ( .A(n5307), .B(n5306), .Z(n5593) );
  XOR U5741 ( .A(n5594), .B(n5593), .Z(n5595) );
  XOR U5742 ( .A(n5596), .B(n5595), .Z(n5541) );
  NANDN U5743 ( .A(n5309), .B(n5308), .Z(n5313) );
  OR U5744 ( .A(n5311), .B(n5310), .Z(n5312) );
  AND U5745 ( .A(n5313), .B(n5312), .Z(n5601) );
  NANDN U5746 ( .A(n29499), .B(n5314), .Z(n5316) );
  XOR U5747 ( .A(b[7]), .B(a[41]), .Z(n5466) );
  NANDN U5748 ( .A(n29735), .B(n5466), .Z(n5315) );
  AND U5749 ( .A(n5316), .B(n5315), .Z(n5557) );
  NANDN U5750 ( .A(n34909), .B(n5317), .Z(n5319) );
  XOR U5751 ( .A(b[31]), .B(a[17]), .Z(n5469) );
  NANDN U5752 ( .A(n35145), .B(n5469), .Z(n5318) );
  AND U5753 ( .A(n5319), .B(n5318), .Z(n5555) );
  NAND U5754 ( .A(b[45]), .B(b[46]), .Z(n5320) );
  AND U5755 ( .A(b[47]), .B(n5320), .Z(n37553) );
  ANDN U5756 ( .B(n37553), .A(n5321), .Z(n5554) );
  XNOR U5757 ( .A(n5555), .B(n5554), .Z(n5556) );
  XOR U5758 ( .A(n5557), .B(n5556), .Z(n5600) );
  NANDN U5759 ( .A(n5322), .B(n31059), .Z(n5324) );
  XOR U5760 ( .A(b[11]), .B(a[37]), .Z(n5487) );
  NANDN U5761 ( .A(n30891), .B(n5487), .Z(n5323) );
  AND U5762 ( .A(n5324), .B(n5323), .Z(n5517) );
  NANDN U5763 ( .A(n5325), .B(n36735), .Z(n5327) );
  XOR U5764 ( .A(b[41]), .B(a[7]), .Z(n5481) );
  NANDN U5765 ( .A(n36594), .B(n5481), .Z(n5326) );
  AND U5766 ( .A(n5327), .B(n5326), .Z(n5515) );
  NANDN U5767 ( .A(n34634), .B(n5328), .Z(n5330) );
  XOR U5768 ( .A(b[29]), .B(a[19]), .Z(n5457) );
  NANDN U5769 ( .A(n34722), .B(n5457), .Z(n5329) );
  NAND U5770 ( .A(n5330), .B(n5329), .Z(n5514) );
  XNOR U5771 ( .A(n5515), .B(n5514), .Z(n5516) );
  XOR U5772 ( .A(n5517), .B(n5516), .Z(n5599) );
  XNOR U5773 ( .A(n5600), .B(n5599), .Z(n5602) );
  NANDN U5774 ( .A(n5332), .B(n5331), .Z(n5336) );
  NANDN U5775 ( .A(n5334), .B(n5333), .Z(n5335) );
  AND U5776 ( .A(n5336), .B(n5335), .Z(n5613) );
  NANDN U5777 ( .A(n28889), .B(n5337), .Z(n5339) );
  XOR U5778 ( .A(b[5]), .B(a[43]), .Z(n5528) );
  NANDN U5779 ( .A(n29138), .B(n5528), .Z(n5338) );
  AND U5780 ( .A(n5339), .B(n5338), .Z(n5511) );
  NANDN U5781 ( .A(n5340), .B(n9942), .Z(n5342) );
  XOR U5782 ( .A(b[3]), .B(a[45]), .Z(n5522) );
  NANDN U5783 ( .A(n28941), .B(n5522), .Z(n5341) );
  AND U5784 ( .A(n5342), .B(n5341), .Z(n5509) );
  NANDN U5785 ( .A(n34223), .B(n5343), .Z(n5345) );
  XOR U5786 ( .A(b[27]), .B(a[21]), .Z(n5525) );
  NANDN U5787 ( .A(n34458), .B(n5525), .Z(n5344) );
  NAND U5788 ( .A(n5345), .B(n5344), .Z(n5508) );
  XNOR U5789 ( .A(n5509), .B(n5508), .Z(n5510) );
  XOR U5790 ( .A(n5511), .B(n5510), .Z(n5612) );
  NANDN U5791 ( .A(n5346), .B(n36238), .Z(n5348) );
  XOR U5792 ( .A(b[37]), .B(a[11]), .Z(n5575) );
  NANDN U5793 ( .A(n36047), .B(n5575), .Z(n5347) );
  AND U5794 ( .A(n5348), .B(n5347), .Z(n5563) );
  NANDN U5795 ( .A(n36210), .B(n5349), .Z(n5351) );
  XOR U5796 ( .A(b[39]), .B(a[9]), .Z(n5478) );
  NANDN U5797 ( .A(n36347), .B(n5478), .Z(n5350) );
  AND U5798 ( .A(n5351), .B(n5350), .Z(n5561) );
  NANDN U5799 ( .A(n31055), .B(n5352), .Z(n5354) );
  XOR U5800 ( .A(b[13]), .B(a[35]), .Z(n5484) );
  NANDN U5801 ( .A(n31293), .B(n5484), .Z(n5353) );
  NAND U5802 ( .A(n5354), .B(n5353), .Z(n5560) );
  XNOR U5803 ( .A(n5561), .B(n5560), .Z(n5562) );
  XOR U5804 ( .A(n5563), .B(n5562), .Z(n5611) );
  XNOR U5805 ( .A(n5612), .B(n5611), .Z(n5614) );
  XOR U5806 ( .A(n5539), .B(n5538), .Z(n5540) );
  XOR U5807 ( .A(n5541), .B(n5540), .Z(n5446) );
  NAND U5808 ( .A(n5356), .B(n5355), .Z(n5360) );
  NANDN U5809 ( .A(n5358), .B(n5357), .Z(n5359) );
  AND U5810 ( .A(n5360), .B(n5359), .Z(n5445) );
  NAND U5811 ( .A(n5362), .B(n5361), .Z(n5366) );
  NANDN U5812 ( .A(n5364), .B(n5363), .Z(n5365) );
  AND U5813 ( .A(n5366), .B(n5365), .Z(n5444) );
  XNOR U5814 ( .A(n5445), .B(n5444), .Z(n5447) );
  XOR U5815 ( .A(n5446), .B(n5447), .Z(n5631) );
  XOR U5816 ( .A(n5632), .B(n5631), .Z(n5617) );
  XNOR U5817 ( .A(n5618), .B(n5617), .Z(n5619) );
  NANDN U5818 ( .A(n5367), .B(n33492), .Z(n5369) );
  XOR U5819 ( .A(b[23]), .B(a[25]), .Z(n5454) );
  NANDN U5820 ( .A(n33644), .B(n5454), .Z(n5368) );
  AND U5821 ( .A(n5369), .B(n5368), .Z(n5499) );
  NANDN U5822 ( .A(n5370), .B(n35928), .Z(n5372) );
  XOR U5823 ( .A(b[35]), .B(a[13]), .Z(n5572) );
  NANDN U5824 ( .A(n35801), .B(n5572), .Z(n5371) );
  AND U5825 ( .A(n5372), .B(n5371), .Z(n5497) );
  NANDN U5826 ( .A(n31536), .B(n5373), .Z(n5375) );
  XOR U5827 ( .A(b[15]), .B(a[33]), .Z(n5578) );
  NANDN U5828 ( .A(n31925), .B(n5578), .Z(n5374) );
  NAND U5829 ( .A(n5375), .B(n5374), .Z(n5496) );
  XNOR U5830 ( .A(n5497), .B(n5496), .Z(n5498) );
  XOR U5831 ( .A(n5499), .B(n5498), .Z(n5606) );
  NANDN U5832 ( .A(n36742), .B(n5376), .Z(n5378) );
  XOR U5833 ( .A(b[43]), .B(a[5]), .Z(n5490) );
  NANDN U5834 ( .A(n36891), .B(n5490), .Z(n5377) );
  AND U5835 ( .A(n5378), .B(n5377), .Z(n5550) );
  NANDN U5836 ( .A(n210), .B(n5379), .Z(n5381) );
  XOR U5837 ( .A(b[9]), .B(a[39]), .Z(n5463) );
  NANDN U5838 ( .A(n30267), .B(n5463), .Z(n5380) );
  AND U5839 ( .A(n5381), .B(n5380), .Z(n5549) );
  NANDN U5840 ( .A(n35260), .B(n5382), .Z(n5384) );
  XOR U5841 ( .A(b[33]), .B(a[15]), .Z(n5493) );
  NANDN U5842 ( .A(n35456), .B(n5493), .Z(n5383) );
  NAND U5843 ( .A(n5384), .B(n5383), .Z(n5548) );
  XOR U5844 ( .A(n5549), .B(n5548), .Z(n5551) );
  XNOR U5845 ( .A(n5550), .B(n5551), .Z(n5605) );
  XOR U5846 ( .A(n5606), .B(n5605), .Z(n5608) );
  NAND U5847 ( .A(n5386), .B(n5385), .Z(n5390) );
  NANDN U5848 ( .A(n5388), .B(n5387), .Z(n5389) );
  AND U5849 ( .A(n5390), .B(n5389), .Z(n5607) );
  XOR U5850 ( .A(n5608), .B(n5607), .Z(n5589) );
  NAND U5851 ( .A(n5392), .B(n5391), .Z(n5396) );
  NANDN U5852 ( .A(n5394), .B(n5393), .Z(n5395) );
  AND U5853 ( .A(n5396), .B(n5395), .Z(n5588) );
  NAND U5854 ( .A(n5398), .B(n5397), .Z(n5402) );
  NANDN U5855 ( .A(n5400), .B(n5399), .Z(n5401) );
  AND U5856 ( .A(n5402), .B(n5401), .Z(n5587) );
  XOR U5857 ( .A(n5588), .B(n5587), .Z(n5590) );
  XOR U5858 ( .A(n5589), .B(n5590), .Z(n5543) );
  NANDN U5859 ( .A(n5404), .B(n5403), .Z(n5408) );
  OR U5860 ( .A(n5406), .B(n5405), .Z(n5407) );
  NAND U5861 ( .A(n5408), .B(n5407), .Z(n5542) );
  XNOR U5862 ( .A(n5543), .B(n5542), .Z(n5545) );
  NANDN U5863 ( .A(n5410), .B(n5409), .Z(n5414) );
  OR U5864 ( .A(n5412), .B(n5411), .Z(n5413) );
  AND U5865 ( .A(n5414), .B(n5413), .Z(n5544) );
  XOR U5866 ( .A(n5545), .B(n5544), .Z(n5624) );
  NANDN U5867 ( .A(n5416), .B(n5415), .Z(n5420) );
  OR U5868 ( .A(n5418), .B(n5417), .Z(n5419) );
  AND U5869 ( .A(n5420), .B(n5419), .Z(n5623) );
  XNOR U5870 ( .A(n5624), .B(n5623), .Z(n5625) );
  NANDN U5871 ( .A(n5422), .B(n5421), .Z(n5426) );
  NAND U5872 ( .A(n5424), .B(n5423), .Z(n5425) );
  NAND U5873 ( .A(n5426), .B(n5425), .Z(n5626) );
  XOR U5874 ( .A(n5625), .B(n5626), .Z(n5620) );
  XOR U5875 ( .A(n5619), .B(n5620), .Z(n5636) );
  XNOR U5876 ( .A(n5635), .B(n5636), .Z(n5639) );
  XOR U5877 ( .A(n5640), .B(n5639), .Z(n5642) );
  XOR U5878 ( .A(n5641), .B(n5642), .Z(n5439) );
  NANDN U5879 ( .A(n5428), .B(n5427), .Z(n5432) );
  NANDN U5880 ( .A(n5430), .B(n5429), .Z(n5431) );
  NAND U5881 ( .A(n5432), .B(n5431), .Z(n5438) );
  XOR U5882 ( .A(n5439), .B(n5438), .Z(n5441) );
  XOR U5883 ( .A(n5440), .B(n5441), .Z(n5433) );
  XNOR U5884 ( .A(n5433), .B(sreg[111]), .Z(n5434) );
  XOR U5885 ( .A(n5435), .B(n5434), .Z(c[111]) );
  NANDN U5886 ( .A(n5433), .B(sreg[111]), .Z(n5437) );
  NAND U5887 ( .A(n5435), .B(n5434), .Z(n5436) );
  AND U5888 ( .A(n5437), .B(n5436), .Z(n5869) );
  XNOR U5889 ( .A(sreg[112]), .B(n5869), .Z(n5871) );
  NANDN U5890 ( .A(n5439), .B(n5438), .Z(n5443) );
  OR U5891 ( .A(n5441), .B(n5440), .Z(n5442) );
  AND U5892 ( .A(n5443), .B(n5442), .Z(n5648) );
  NANDN U5893 ( .A(n32483), .B(n5448), .Z(n5450) );
  XOR U5894 ( .A(b[19]), .B(a[30]), .Z(n5690) );
  NANDN U5895 ( .A(n32823), .B(n5690), .Z(n5449) );
  AND U5896 ( .A(n5450), .B(n5449), .Z(n5840) );
  NANDN U5897 ( .A(n32996), .B(n5451), .Z(n5453) );
  XOR U5898 ( .A(b[21]), .B(a[28]), .Z(n5696) );
  NANDN U5899 ( .A(n33271), .B(n5696), .Z(n5452) );
  NAND U5900 ( .A(n5453), .B(n5452), .Z(n5839) );
  XNOR U5901 ( .A(n5840), .B(n5839), .Z(n5842) );
  NANDN U5902 ( .A(n33866), .B(n5454), .Z(n5456) );
  XOR U5903 ( .A(b[23]), .B(a[26]), .Z(n5751) );
  NANDN U5904 ( .A(n33644), .B(n5751), .Z(n5455) );
  AND U5905 ( .A(n5456), .B(n5455), .Z(n5848) );
  NANDN U5906 ( .A(n34634), .B(n5457), .Z(n5459) );
  XOR U5907 ( .A(b[29]), .B(a[20]), .Z(n5693) );
  NANDN U5908 ( .A(n34722), .B(n5693), .Z(n5458) );
  AND U5909 ( .A(n5459), .B(n5458), .Z(n5846) );
  NANDN U5910 ( .A(n32013), .B(n5460), .Z(n5462) );
  XOR U5911 ( .A(b[17]), .B(a[32]), .Z(n5699) );
  NANDN U5912 ( .A(n32292), .B(n5699), .Z(n5461) );
  NAND U5913 ( .A(n5462), .B(n5461), .Z(n5845) );
  XNOR U5914 ( .A(n5846), .B(n5845), .Z(n5847) );
  XNOR U5915 ( .A(n5848), .B(n5847), .Z(n5841) );
  XOR U5916 ( .A(n5842), .B(n5841), .Z(n5716) );
  NANDN U5917 ( .A(n210), .B(n5463), .Z(n5465) );
  XOR U5918 ( .A(b[9]), .B(a[40]), .Z(n5797) );
  NANDN U5919 ( .A(n30267), .B(n5797), .Z(n5464) );
  AND U5920 ( .A(n5465), .B(n5464), .Z(n5704) );
  NANDN U5921 ( .A(n29499), .B(n5466), .Z(n5468) );
  XOR U5922 ( .A(b[7]), .B(a[42]), .Z(n5821) );
  NANDN U5923 ( .A(n29735), .B(n5821), .Z(n5467) );
  AND U5924 ( .A(n5468), .B(n5467), .Z(n5703) );
  NANDN U5925 ( .A(n34909), .B(n5469), .Z(n5471) );
  XOR U5926 ( .A(b[31]), .B(a[18]), .Z(n5824) );
  NANDN U5927 ( .A(n35145), .B(n5824), .Z(n5470) );
  NAND U5928 ( .A(n5471), .B(n5470), .Z(n5702) );
  XOR U5929 ( .A(n5703), .B(n5702), .Z(n5705) );
  XOR U5930 ( .A(n5704), .B(n5705), .Z(n5715) );
  NANDN U5931 ( .A(n5473), .B(n5472), .Z(n5477) );
  NANDN U5932 ( .A(n5475), .B(n5474), .Z(n5476) );
  AND U5933 ( .A(n5477), .B(n5476), .Z(n5714) );
  XOR U5934 ( .A(n5715), .B(n5714), .Z(n5717) );
  XOR U5935 ( .A(n5716), .B(n5717), .Z(n5728) );
  NANDN U5936 ( .A(n36210), .B(n5478), .Z(n5480) );
  XOR U5937 ( .A(b[39]), .B(a[10]), .Z(n5809) );
  NANDN U5938 ( .A(n36347), .B(n5809), .Z(n5479) );
  AND U5939 ( .A(n5480), .B(n5479), .Z(n5756) );
  NANDN U5940 ( .A(n36480), .B(n5481), .Z(n5483) );
  XOR U5941 ( .A(b[41]), .B(a[8]), .Z(n5812) );
  NANDN U5942 ( .A(n36594), .B(n5812), .Z(n5482) );
  AND U5943 ( .A(n5483), .B(n5482), .Z(n5755) );
  NANDN U5944 ( .A(n31055), .B(n5484), .Z(n5486) );
  XOR U5945 ( .A(b[13]), .B(a[36]), .Z(n5815) );
  NANDN U5946 ( .A(n31293), .B(n5815), .Z(n5485) );
  NAND U5947 ( .A(n5486), .B(n5485), .Z(n5754) );
  XOR U5948 ( .A(n5755), .B(n5754), .Z(n5757) );
  XOR U5949 ( .A(n5756), .B(n5757), .Z(n5733) );
  NANDN U5950 ( .A(n30482), .B(n5487), .Z(n5489) );
  XOR U5951 ( .A(b[11]), .B(a[38]), .Z(n5794) );
  NANDN U5952 ( .A(n30891), .B(n5794), .Z(n5488) );
  AND U5953 ( .A(n5489), .B(n5488), .Z(n5710) );
  NANDN U5954 ( .A(n36742), .B(n5490), .Z(n5492) );
  XOR U5955 ( .A(b[43]), .B(a[6]), .Z(n5818) );
  NANDN U5956 ( .A(n36891), .B(n5818), .Z(n5491) );
  AND U5957 ( .A(n5492), .B(n5491), .Z(n5709) );
  NANDN U5958 ( .A(n35260), .B(n5493), .Z(n5495) );
  XOR U5959 ( .A(b[33]), .B(a[16]), .Z(n5800) );
  NANDN U5960 ( .A(n35456), .B(n5800), .Z(n5494) );
  NAND U5961 ( .A(n5495), .B(n5494), .Z(n5708) );
  XOR U5962 ( .A(n5709), .B(n5708), .Z(n5711) );
  XNOR U5963 ( .A(n5710), .B(n5711), .Z(n5732) );
  XNOR U5964 ( .A(n5733), .B(n5732), .Z(n5735) );
  NANDN U5965 ( .A(n5497), .B(n5496), .Z(n5501) );
  NANDN U5966 ( .A(n5499), .B(n5498), .Z(n5500) );
  AND U5967 ( .A(n5501), .B(n5500), .Z(n5734) );
  XOR U5968 ( .A(n5735), .B(n5734), .Z(n5769) );
  NANDN U5969 ( .A(n5503), .B(n5502), .Z(n5507) );
  OR U5970 ( .A(n5505), .B(n5504), .Z(n5506) );
  AND U5971 ( .A(n5507), .B(n5506), .Z(n5767) );
  NANDN U5972 ( .A(n5509), .B(n5508), .Z(n5513) );
  NANDN U5973 ( .A(n5511), .B(n5510), .Z(n5512) );
  NAND U5974 ( .A(n5513), .B(n5512), .Z(n5766) );
  XNOR U5975 ( .A(n5767), .B(n5766), .Z(n5768) );
  XNOR U5976 ( .A(n5769), .B(n5768), .Z(n5726) );
  NANDN U5977 ( .A(n5515), .B(n5514), .Z(n5519) );
  NANDN U5978 ( .A(n5517), .B(n5516), .Z(n5518) );
  AND U5979 ( .A(n5519), .B(n5518), .Z(n5836) );
  ANDN U5980 ( .B(n5521), .A(n5520), .Z(n5853) );
  NAND U5981 ( .A(n9942), .B(n5522), .Z(n5524) );
  XNOR U5982 ( .A(b[3]), .B(a[46]), .Z(n5748) );
  NANDN U5983 ( .A(n5748), .B(n9653), .Z(n5523) );
  AND U5984 ( .A(n5524), .B(n5523), .Z(n5851) );
  NAND U5985 ( .A(n34647), .B(n5525), .Z(n5527) );
  XNOR U5986 ( .A(b[27]), .B(a[22]), .Z(n5741) );
  NANDN U5987 ( .A(n5741), .B(n34648), .Z(n5526) );
  NAND U5988 ( .A(n5527), .B(n5526), .Z(n5852) );
  XOR U5989 ( .A(n5851), .B(n5852), .Z(n5854) );
  XOR U5990 ( .A(n5853), .B(n5854), .Z(n5834) );
  NANDN U5991 ( .A(n28889), .B(n5528), .Z(n5530) );
  XOR U5992 ( .A(b[5]), .B(a[44]), .Z(n5745) );
  NANDN U5993 ( .A(n29138), .B(n5745), .Z(n5529) );
  AND U5994 ( .A(n5530), .B(n5529), .Z(n5806) );
  ANDN U5995 ( .B(n5531), .A(n37341), .Z(n37294) );
  NANDN U5996 ( .A(n211), .B(n5532), .Z(n5534) );
  XOR U5997 ( .A(b[47]), .B(a[2]), .Z(n5784) );
  NANDN U5998 ( .A(n37172), .B(n5784), .Z(n5533) );
  AND U5999 ( .A(n5534), .B(n5533), .Z(n5804) );
  NANDN U6000 ( .A(n33875), .B(n5535), .Z(n5537) );
  XOR U6001 ( .A(b[25]), .B(a[24]), .Z(n5781) );
  NANDN U6002 ( .A(n33994), .B(n5781), .Z(n5536) );
  NAND U6003 ( .A(n5537), .B(n5536), .Z(n5803) );
  XNOR U6004 ( .A(n5804), .B(n5803), .Z(n5805) );
  XNOR U6005 ( .A(n5806), .B(n5805), .Z(n5833) );
  XNOR U6006 ( .A(n5834), .B(n5833), .Z(n5835) );
  XOR U6007 ( .A(n5836), .B(n5835), .Z(n5727) );
  XOR U6008 ( .A(n5726), .B(n5727), .Z(n5729) );
  XOR U6009 ( .A(n5728), .B(n5729), .Z(n5858) );
  XNOR U6010 ( .A(n5858), .B(n5857), .Z(n5859) );
  XOR U6011 ( .A(n5860), .B(n5859), .Z(n5659) );
  NANDN U6012 ( .A(n5543), .B(n5542), .Z(n5547) );
  NAND U6013 ( .A(n5545), .B(n5544), .Z(n5546) );
  AND U6014 ( .A(n5547), .B(n5546), .Z(n5657) );
  NANDN U6015 ( .A(n5549), .B(n5548), .Z(n5553) );
  OR U6016 ( .A(n5551), .B(n5550), .Z(n5552) );
  AND U6017 ( .A(n5553), .B(n5552), .Z(n5721) );
  NANDN U6018 ( .A(n5555), .B(n5554), .Z(n5559) );
  NANDN U6019 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U6020 ( .A(n5559), .B(n5558), .Z(n5720) );
  XNOR U6021 ( .A(n5721), .B(n5720), .Z(n5723) );
  NANDN U6022 ( .A(n5561), .B(n5560), .Z(n5565) );
  NANDN U6023 ( .A(n5563), .B(n5562), .Z(n5564) );
  AND U6024 ( .A(n5565), .B(n5564), .Z(n5763) );
  NAND U6025 ( .A(b[0]), .B(a[48]), .Z(n5566) );
  XNOR U6026 ( .A(b[1]), .B(n5566), .Z(n5568) );
  NANDN U6027 ( .A(b[0]), .B(a[47]), .Z(n5567) );
  NAND U6028 ( .A(n5568), .B(n5567), .Z(n5775) );
  XOR U6029 ( .A(b[48]), .B(b[47]), .Z(n37537) );
  IV U6030 ( .A(n37537), .Z(n37432) );
  ANDN U6031 ( .B(a[0]), .A(n37432), .Z(n5772) );
  IV U6032 ( .A(n37202), .Z(n36991) );
  NANDN U6033 ( .A(n36991), .B(n5569), .Z(n5571) );
  XOR U6034 ( .A(b[45]), .B(a[4]), .Z(n5738) );
  NANDN U6035 ( .A(n37083), .B(n5738), .Z(n5570) );
  AND U6036 ( .A(n5571), .B(n5570), .Z(n5773) );
  XNOR U6037 ( .A(n5772), .B(n5773), .Z(n5774) );
  XNOR U6038 ( .A(n5775), .B(n5774), .Z(n5760) );
  NANDN U6039 ( .A(n35611), .B(n5572), .Z(n5574) );
  XOR U6040 ( .A(b[35]), .B(a[14]), .Z(n5681) );
  NANDN U6041 ( .A(n35801), .B(n5681), .Z(n5573) );
  AND U6042 ( .A(n5574), .B(n5573), .Z(n5830) );
  NANDN U6043 ( .A(n35936), .B(n5575), .Z(n5577) );
  XOR U6044 ( .A(b[37]), .B(a[12]), .Z(n5684) );
  NANDN U6045 ( .A(n36047), .B(n5684), .Z(n5576) );
  AND U6046 ( .A(n5577), .B(n5576), .Z(n5828) );
  NANDN U6047 ( .A(n31536), .B(n5578), .Z(n5580) );
  XOR U6048 ( .A(b[15]), .B(a[34]), .Z(n5687) );
  NANDN U6049 ( .A(n31925), .B(n5687), .Z(n5579) );
  NAND U6050 ( .A(n5580), .B(n5579), .Z(n5827) );
  XNOR U6051 ( .A(n5828), .B(n5827), .Z(n5829) );
  XOR U6052 ( .A(n5830), .B(n5829), .Z(n5761) );
  XNOR U6053 ( .A(n5760), .B(n5761), .Z(n5762) );
  XNOR U6054 ( .A(n5763), .B(n5762), .Z(n5722) );
  XOR U6055 ( .A(n5723), .B(n5722), .Z(n5664) );
  NAND U6056 ( .A(n5582), .B(n5581), .Z(n5586) );
  NAND U6057 ( .A(n5584), .B(n5583), .Z(n5585) );
  AND U6058 ( .A(n5586), .B(n5585), .Z(n5663) );
  XNOR U6059 ( .A(n5664), .B(n5663), .Z(n5666) );
  NANDN U6060 ( .A(n5588), .B(n5587), .Z(n5592) );
  OR U6061 ( .A(n5590), .B(n5589), .Z(n5591) );
  AND U6062 ( .A(n5592), .B(n5591), .Z(n5665) );
  XOR U6063 ( .A(n5666), .B(n5665), .Z(n5678) );
  NAND U6064 ( .A(n5594), .B(n5593), .Z(n5598) );
  NAND U6065 ( .A(n5596), .B(n5595), .Z(n5597) );
  AND U6066 ( .A(n5598), .B(n5597), .Z(n5672) );
  NAND U6067 ( .A(n5600), .B(n5599), .Z(n5604) );
  NANDN U6068 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U6069 ( .A(n5604), .B(n5603), .Z(n5669) );
  NAND U6070 ( .A(n5606), .B(n5605), .Z(n5610) );
  NAND U6071 ( .A(n5608), .B(n5607), .Z(n5609) );
  NAND U6072 ( .A(n5610), .B(n5609), .Z(n5670) );
  XNOR U6073 ( .A(n5669), .B(n5670), .Z(n5671) );
  XNOR U6074 ( .A(n5672), .B(n5671), .Z(n5675) );
  NAND U6075 ( .A(n5612), .B(n5611), .Z(n5616) );
  NANDN U6076 ( .A(n5614), .B(n5613), .Z(n5615) );
  NAND U6077 ( .A(n5616), .B(n5615), .Z(n5676) );
  XNOR U6078 ( .A(n5675), .B(n5676), .Z(n5677) );
  XOR U6079 ( .A(n5678), .B(n5677), .Z(n5658) );
  XOR U6080 ( .A(n5657), .B(n5658), .Z(n5660) );
  XOR U6081 ( .A(n5659), .B(n5660), .Z(n5864) );
  NANDN U6082 ( .A(n5618), .B(n5617), .Z(n5622) );
  NANDN U6083 ( .A(n5620), .B(n5619), .Z(n5621) );
  AND U6084 ( .A(n5622), .B(n5621), .Z(n5653) );
  NANDN U6085 ( .A(n5624), .B(n5623), .Z(n5628) );
  NANDN U6086 ( .A(n5626), .B(n5625), .Z(n5627) );
  AND U6087 ( .A(n5628), .B(n5627), .Z(n5652) );
  XOR U6088 ( .A(n5652), .B(n5651), .Z(n5654) );
  XNOR U6089 ( .A(n5653), .B(n5654), .Z(n5863) );
  XNOR U6090 ( .A(n5864), .B(n5863), .Z(n5865) );
  NANDN U6091 ( .A(n5634), .B(n5633), .Z(n5638) );
  NANDN U6092 ( .A(n5636), .B(n5635), .Z(n5637) );
  NAND U6093 ( .A(n5638), .B(n5637), .Z(n5866) );
  XNOR U6094 ( .A(n5865), .B(n5866), .Z(n5645) );
  NANDN U6095 ( .A(n5640), .B(n5639), .Z(n5644) );
  OR U6096 ( .A(n5642), .B(n5641), .Z(n5643) );
  NAND U6097 ( .A(n5644), .B(n5643), .Z(n5646) );
  XNOR U6098 ( .A(n5645), .B(n5646), .Z(n5647) );
  XNOR U6099 ( .A(n5648), .B(n5647), .Z(n5870) );
  XNOR U6100 ( .A(n5871), .B(n5870), .Z(c[112]) );
  NANDN U6101 ( .A(n5646), .B(n5645), .Z(n5650) );
  NANDN U6102 ( .A(n5648), .B(n5647), .Z(n5649) );
  AND U6103 ( .A(n5650), .B(n5649), .Z(n5882) );
  NANDN U6104 ( .A(n5652), .B(n5651), .Z(n5656) );
  OR U6105 ( .A(n5654), .B(n5653), .Z(n5655) );
  AND U6106 ( .A(n5656), .B(n5655), .Z(n6097) );
  NANDN U6107 ( .A(n5658), .B(n5657), .Z(n5662) );
  OR U6108 ( .A(n5660), .B(n5659), .Z(n5661) );
  AND U6109 ( .A(n5662), .B(n5661), .Z(n6096) );
  NANDN U6110 ( .A(n5664), .B(n5663), .Z(n5668) );
  NAND U6111 ( .A(n5666), .B(n5665), .Z(n5667) );
  AND U6112 ( .A(n5668), .B(n5667), .Z(n5892) );
  NANDN U6113 ( .A(n5670), .B(n5669), .Z(n5674) );
  NANDN U6114 ( .A(n5672), .B(n5671), .Z(n5673) );
  NAND U6115 ( .A(n5674), .B(n5673), .Z(n5891) );
  XOR U6116 ( .A(n5892), .B(n5891), .Z(n5894) );
  NANDN U6117 ( .A(n5676), .B(n5675), .Z(n5680) );
  NANDN U6118 ( .A(n5678), .B(n5677), .Z(n5679) );
  NAND U6119 ( .A(n5680), .B(n5679), .Z(n5893) );
  XOR U6120 ( .A(n5894), .B(n5893), .Z(n5887) );
  NANDN U6121 ( .A(n35611), .B(n5681), .Z(n5683) );
  XOR U6122 ( .A(b[35]), .B(a[15]), .Z(n6035) );
  NANDN U6123 ( .A(n35801), .B(n6035), .Z(n5682) );
  AND U6124 ( .A(n5683), .B(n5682), .Z(n5987) );
  NANDN U6125 ( .A(n35936), .B(n5684), .Z(n5686) );
  XOR U6126 ( .A(b[37]), .B(a[13]), .Z(n5933) );
  NANDN U6127 ( .A(n36047), .B(n5933), .Z(n5685) );
  AND U6128 ( .A(n5686), .B(n5685), .Z(n5986) );
  NANDN U6129 ( .A(n31536), .B(n5687), .Z(n5689) );
  XOR U6130 ( .A(b[15]), .B(a[35]), .Z(n6026) );
  NANDN U6131 ( .A(n31925), .B(n6026), .Z(n5688) );
  NAND U6132 ( .A(n5689), .B(n5688), .Z(n5985) );
  XOR U6133 ( .A(n5986), .B(n5985), .Z(n5988) );
  XOR U6134 ( .A(n5987), .B(n5988), .Z(n5957) );
  NANDN U6135 ( .A(n32483), .B(n5690), .Z(n5692) );
  XOR U6136 ( .A(b[19]), .B(a[31]), .Z(n6000) );
  NANDN U6137 ( .A(n32823), .B(n6000), .Z(n5691) );
  AND U6138 ( .A(n5692), .B(n5691), .Z(n6008) );
  NANDN U6139 ( .A(n34634), .B(n5693), .Z(n5695) );
  XOR U6140 ( .A(b[29]), .B(a[21]), .Z(n5915) );
  NANDN U6141 ( .A(n34722), .B(n5915), .Z(n5694) );
  AND U6142 ( .A(n5695), .B(n5694), .Z(n6007) );
  NANDN U6143 ( .A(n32996), .B(n5696), .Z(n5698) );
  XOR U6144 ( .A(b[21]), .B(a[29]), .Z(n6003) );
  NANDN U6145 ( .A(n33271), .B(n6003), .Z(n5697) );
  NAND U6146 ( .A(n5698), .B(n5697), .Z(n6006) );
  XOR U6147 ( .A(n6007), .B(n6006), .Z(n6009) );
  XOR U6148 ( .A(n6008), .B(n6009), .Z(n5956) );
  NAND U6149 ( .A(n32544), .B(n5699), .Z(n5701) );
  XNOR U6150 ( .A(b[17]), .B(a[33]), .Z(n5997) );
  NANDN U6151 ( .A(n5997), .B(n32545), .Z(n5700) );
  AND U6152 ( .A(n5701), .B(n5700), .Z(n5955) );
  XOR U6153 ( .A(n5956), .B(n5955), .Z(n5958) );
  XOR U6154 ( .A(n5957), .B(n5958), .Z(n6085) );
  NANDN U6155 ( .A(n5703), .B(n5702), .Z(n5707) );
  OR U6156 ( .A(n5705), .B(n5704), .Z(n5706) );
  AND U6157 ( .A(n5707), .B(n5706), .Z(n6084) );
  NANDN U6158 ( .A(n5709), .B(n5708), .Z(n5713) );
  OR U6159 ( .A(n5711), .B(n5710), .Z(n5712) );
  NAND U6160 ( .A(n5713), .B(n5712), .Z(n6083) );
  XOR U6161 ( .A(n6084), .B(n6083), .Z(n6086) );
  XOR U6162 ( .A(n6085), .B(n6086), .Z(n6090) );
  NANDN U6163 ( .A(n5715), .B(n5714), .Z(n5719) );
  OR U6164 ( .A(n5717), .B(n5716), .Z(n5718) );
  NAND U6165 ( .A(n5719), .B(n5718), .Z(n6089) );
  XNOR U6166 ( .A(n6090), .B(n6089), .Z(n6092) );
  NANDN U6167 ( .A(n5721), .B(n5720), .Z(n5725) );
  NAND U6168 ( .A(n5723), .B(n5722), .Z(n5724) );
  AND U6169 ( .A(n5725), .B(n5724), .Z(n6091) );
  XOR U6170 ( .A(n6092), .B(n6091), .Z(n5904) );
  NANDN U6171 ( .A(n5727), .B(n5726), .Z(n5731) );
  OR U6172 ( .A(n5729), .B(n5728), .Z(n5730) );
  NAND U6173 ( .A(n5731), .B(n5730), .Z(n5903) );
  XNOR U6174 ( .A(n5904), .B(n5903), .Z(n5905) );
  NANDN U6175 ( .A(n5733), .B(n5732), .Z(n5737) );
  NAND U6176 ( .A(n5735), .B(n5734), .Z(n5736) );
  AND U6177 ( .A(n5737), .B(n5736), .Z(n5963) );
  NANDN U6178 ( .A(n36991), .B(n5738), .Z(n5740) );
  XOR U6179 ( .A(b[45]), .B(a[5]), .Z(n6029) );
  NANDN U6180 ( .A(n37083), .B(n6029), .Z(n5739) );
  AND U6181 ( .A(n5740), .B(n5739), .Z(n5981) );
  NANDN U6182 ( .A(n5741), .B(n34647), .Z(n5743) );
  XOR U6183 ( .A(b[27]), .B(a[23]), .Z(n6015) );
  NANDN U6184 ( .A(n34458), .B(n6015), .Z(n5742) );
  AND U6185 ( .A(n5743), .B(n5742), .Z(n5980) );
  NAND U6186 ( .A(b[47]), .B(b[48]), .Z(n5744) );
  NAND U6187 ( .A(b[49]), .B(n5744), .Z(n5788) );
  IV U6188 ( .A(n5788), .Z(n37724) );
  ANDN U6189 ( .B(n37724), .A(n5772), .Z(n5979) );
  XOR U6190 ( .A(n5980), .B(n5979), .Z(n5982) );
  XOR U6191 ( .A(n5981), .B(n5982), .Z(n6072) );
  NANDN U6192 ( .A(n28889), .B(n5745), .Z(n5747) );
  XOR U6193 ( .A(b[5]), .B(a[45]), .Z(n5912) );
  NANDN U6194 ( .A(n29138), .B(n5912), .Z(n5746) );
  AND U6195 ( .A(n5747), .B(n5746), .Z(n5975) );
  NANDN U6196 ( .A(n5748), .B(n9942), .Z(n5750) );
  XOR U6197 ( .A(b[3]), .B(a[47]), .Z(n6012) );
  NANDN U6198 ( .A(n28941), .B(n6012), .Z(n5749) );
  AND U6199 ( .A(n5750), .B(n5749), .Z(n5974) );
  NANDN U6200 ( .A(n33866), .B(n5751), .Z(n5753) );
  XOR U6201 ( .A(b[23]), .B(a[27]), .Z(n6020) );
  NANDN U6202 ( .A(n33644), .B(n6020), .Z(n5752) );
  NAND U6203 ( .A(n5753), .B(n5752), .Z(n5973) );
  XOR U6204 ( .A(n5974), .B(n5973), .Z(n5976) );
  XNOR U6205 ( .A(n5975), .B(n5976), .Z(n6071) );
  XNOR U6206 ( .A(n6072), .B(n6071), .Z(n6073) );
  NANDN U6207 ( .A(n5755), .B(n5754), .Z(n5759) );
  OR U6208 ( .A(n5757), .B(n5756), .Z(n5758) );
  NAND U6209 ( .A(n5759), .B(n5758), .Z(n6074) );
  XNOR U6210 ( .A(n6073), .B(n6074), .Z(n5961) );
  NANDN U6211 ( .A(n5761), .B(n5760), .Z(n5765) );
  NANDN U6212 ( .A(n5763), .B(n5762), .Z(n5764) );
  NAND U6213 ( .A(n5765), .B(n5764), .Z(n5962) );
  XOR U6214 ( .A(n5961), .B(n5962), .Z(n5964) );
  XOR U6215 ( .A(n5963), .B(n5964), .Z(n5900) );
  NANDN U6216 ( .A(n5767), .B(n5766), .Z(n5771) );
  NANDN U6217 ( .A(n5769), .B(n5768), .Z(n5770) );
  AND U6218 ( .A(n5771), .B(n5770), .Z(n5898) );
  NANDN U6219 ( .A(n5773), .B(n5772), .Z(n5777) );
  NANDN U6220 ( .A(n5775), .B(n5774), .Z(n5776) );
  AND U6221 ( .A(n5777), .B(n5776), .Z(n6055) );
  NAND U6222 ( .A(b[0]), .B(a[49]), .Z(n5778) );
  XNOR U6223 ( .A(b[1]), .B(n5778), .Z(n5780) );
  NANDN U6224 ( .A(b[0]), .B(a[48]), .Z(n5779) );
  NAND U6225 ( .A(n5780), .B(n5779), .Z(n5919) );
  NANDN U6226 ( .A(n33875), .B(n5781), .Z(n5783) );
  XOR U6227 ( .A(b[25]), .B(a[25]), .Z(n6023) );
  NANDN U6228 ( .A(n33994), .B(n6023), .Z(n5782) );
  NAND U6229 ( .A(n5783), .B(n5782), .Z(n5918) );
  XNOR U6230 ( .A(n5919), .B(n5918), .Z(n5920) );
  NANDN U6231 ( .A(n211), .B(n5784), .Z(n5786) );
  XOR U6232 ( .A(b[47]), .B(a[3]), .Z(n5991) );
  NANDN U6233 ( .A(n37172), .B(n5991), .Z(n5785) );
  AND U6234 ( .A(n5786), .B(n5785), .Z(n6018) );
  XOR U6235 ( .A(b[49]), .B(a[1]), .Z(n5940) );
  NANDN U6236 ( .A(n37432), .B(n5940), .Z(n5793) );
  ANDN U6237 ( .B(b[48]), .A(b[49]), .Z(n5787) );
  NAND U6238 ( .A(n5787), .B(a[0]), .Z(n5790) );
  OR U6239 ( .A(a[0]), .B(n5788), .Z(n5789) );
  NAND U6240 ( .A(n5790), .B(n5789), .Z(n5791) );
  NAND U6241 ( .A(n37432), .B(n5791), .Z(n5792) );
  NAND U6242 ( .A(n5793), .B(n5792), .Z(n6019) );
  XOR U6243 ( .A(n6018), .B(n6019), .Z(n5921) );
  XNOR U6244 ( .A(n5920), .B(n5921), .Z(n6053) );
  NANDN U6245 ( .A(n30482), .B(n5794), .Z(n5796) );
  XOR U6246 ( .A(b[11]), .B(a[39]), .Z(n6032) );
  NANDN U6247 ( .A(n30891), .B(n6032), .Z(n5795) );
  AND U6248 ( .A(n5796), .B(n5795), .Z(n6050) );
  NANDN U6249 ( .A(n210), .B(n5797), .Z(n5799) );
  XOR U6250 ( .A(b[9]), .B(a[41]), .Z(n5943) );
  NANDN U6251 ( .A(n30267), .B(n5943), .Z(n5798) );
  AND U6252 ( .A(n5799), .B(n5798), .Z(n6048) );
  NANDN U6253 ( .A(n35260), .B(n5800), .Z(n5802) );
  XOR U6254 ( .A(b[33]), .B(a[17]), .Z(n5946) );
  NANDN U6255 ( .A(n35456), .B(n5946), .Z(n5801) );
  NAND U6256 ( .A(n5802), .B(n5801), .Z(n6047) );
  XNOR U6257 ( .A(n6048), .B(n6047), .Z(n6049) );
  XOR U6258 ( .A(n6050), .B(n6049), .Z(n6054) );
  XOR U6259 ( .A(n6053), .B(n6054), .Z(n6056) );
  XOR U6260 ( .A(n6055), .B(n6056), .Z(n6066) );
  NANDN U6261 ( .A(n5804), .B(n5803), .Z(n5808) );
  NANDN U6262 ( .A(n5806), .B(n5805), .Z(n5807) );
  AND U6263 ( .A(n5808), .B(n5807), .Z(n6065) );
  XNOR U6264 ( .A(n6066), .B(n6065), .Z(n6068) );
  NANDN U6265 ( .A(n36210), .B(n5809), .Z(n5811) );
  XOR U6266 ( .A(b[39]), .B(a[11]), .Z(n6038) );
  NANDN U6267 ( .A(n36347), .B(n6038), .Z(n5810) );
  AND U6268 ( .A(n5811), .B(n5810), .Z(n5951) );
  NANDN U6269 ( .A(n36480), .B(n5812), .Z(n5814) );
  XOR U6270 ( .A(b[41]), .B(a[9]), .Z(n6041) );
  NANDN U6271 ( .A(n36594), .B(n6041), .Z(n5813) );
  AND U6272 ( .A(n5814), .B(n5813), .Z(n5950) );
  NANDN U6273 ( .A(n31055), .B(n5815), .Z(n5817) );
  XOR U6274 ( .A(b[13]), .B(a[37]), .Z(n5936) );
  NANDN U6275 ( .A(n31293), .B(n5936), .Z(n5816) );
  NAND U6276 ( .A(n5817), .B(n5816), .Z(n5949) );
  XOR U6277 ( .A(n5950), .B(n5949), .Z(n5952) );
  XOR U6278 ( .A(n5951), .B(n5952), .Z(n6060) );
  NANDN U6279 ( .A(n36742), .B(n5818), .Z(n5820) );
  XOR U6280 ( .A(b[43]), .B(a[7]), .Z(n6044) );
  NANDN U6281 ( .A(n36891), .B(n6044), .Z(n5819) );
  AND U6282 ( .A(n5820), .B(n5819), .Z(n5926) );
  NANDN U6283 ( .A(n29499), .B(n5821), .Z(n5823) );
  XOR U6284 ( .A(b[7]), .B(a[43]), .Z(n5909) );
  NANDN U6285 ( .A(n29735), .B(n5909), .Z(n5822) );
  AND U6286 ( .A(n5823), .B(n5822), .Z(n5925) );
  NANDN U6287 ( .A(n34909), .B(n5824), .Z(n5826) );
  XOR U6288 ( .A(b[31]), .B(a[19]), .Z(n5930) );
  NANDN U6289 ( .A(n35145), .B(n5930), .Z(n5825) );
  NAND U6290 ( .A(n5826), .B(n5825), .Z(n5924) );
  XOR U6291 ( .A(n5925), .B(n5924), .Z(n5927) );
  XNOR U6292 ( .A(n5926), .B(n5927), .Z(n6059) );
  XNOR U6293 ( .A(n6060), .B(n6059), .Z(n6061) );
  NANDN U6294 ( .A(n5828), .B(n5827), .Z(n5832) );
  NANDN U6295 ( .A(n5830), .B(n5829), .Z(n5831) );
  NAND U6296 ( .A(n5832), .B(n5831), .Z(n6062) );
  XNOR U6297 ( .A(n6061), .B(n6062), .Z(n6067) );
  XOR U6298 ( .A(n6068), .B(n6067), .Z(n5970) );
  NANDN U6299 ( .A(n5834), .B(n5833), .Z(n5838) );
  NANDN U6300 ( .A(n5836), .B(n5835), .Z(n5837) );
  AND U6301 ( .A(n5838), .B(n5837), .Z(n5968) );
  NANDN U6302 ( .A(n5840), .B(n5839), .Z(n5844) );
  NAND U6303 ( .A(n5842), .B(n5841), .Z(n5843) );
  AND U6304 ( .A(n5844), .B(n5843), .Z(n6080) );
  NANDN U6305 ( .A(n5846), .B(n5845), .Z(n5850) );
  NANDN U6306 ( .A(n5848), .B(n5847), .Z(n5849) );
  AND U6307 ( .A(n5850), .B(n5849), .Z(n6078) );
  NANDN U6308 ( .A(n5852), .B(n5851), .Z(n5856) );
  OR U6309 ( .A(n5854), .B(n5853), .Z(n5855) );
  AND U6310 ( .A(n5856), .B(n5855), .Z(n6077) );
  XNOR U6311 ( .A(n6078), .B(n6077), .Z(n6079) );
  XNOR U6312 ( .A(n6080), .B(n6079), .Z(n5967) );
  XNOR U6313 ( .A(n5968), .B(n5967), .Z(n5969) );
  XNOR U6314 ( .A(n5970), .B(n5969), .Z(n5897) );
  XNOR U6315 ( .A(n5898), .B(n5897), .Z(n5899) );
  XOR U6316 ( .A(n5900), .B(n5899), .Z(n5906) );
  XNOR U6317 ( .A(n5905), .B(n5906), .Z(n5885) );
  NANDN U6318 ( .A(n5858), .B(n5857), .Z(n5862) );
  NAND U6319 ( .A(n5860), .B(n5859), .Z(n5861) );
  NAND U6320 ( .A(n5862), .B(n5861), .Z(n5886) );
  XOR U6321 ( .A(n5885), .B(n5886), .Z(n5888) );
  XNOR U6322 ( .A(n5887), .B(n5888), .Z(n6095) );
  XOR U6323 ( .A(n6096), .B(n6095), .Z(n6098) );
  XOR U6324 ( .A(n6097), .B(n6098), .Z(n5880) );
  NANDN U6325 ( .A(n5864), .B(n5863), .Z(n5868) );
  NANDN U6326 ( .A(n5866), .B(n5865), .Z(n5867) );
  NAND U6327 ( .A(n5868), .B(n5867), .Z(n5879) );
  XNOR U6328 ( .A(n5880), .B(n5879), .Z(n5881) );
  XNOR U6329 ( .A(n5882), .B(n5881), .Z(n5874) );
  XNOR U6330 ( .A(sreg[113]), .B(n5874), .Z(n5876) );
  NANDN U6331 ( .A(sreg[112]), .B(n5869), .Z(n5873) );
  NAND U6332 ( .A(n5871), .B(n5870), .Z(n5872) );
  NAND U6333 ( .A(n5873), .B(n5872), .Z(n5875) );
  XNOR U6334 ( .A(n5876), .B(n5875), .Z(c[113]) );
  NANDN U6335 ( .A(sreg[113]), .B(n5874), .Z(n5878) );
  NAND U6336 ( .A(n5876), .B(n5875), .Z(n5877) );
  NAND U6337 ( .A(n5878), .B(n5877), .Z(n6329) );
  XNOR U6338 ( .A(sreg[114]), .B(n6329), .Z(n6331) );
  NANDN U6339 ( .A(n5880), .B(n5879), .Z(n5884) );
  NANDN U6340 ( .A(n5882), .B(n5881), .Z(n5883) );
  AND U6341 ( .A(n5884), .B(n5883), .Z(n6104) );
  NANDN U6342 ( .A(n5886), .B(n5885), .Z(n5890) );
  NANDN U6343 ( .A(n5888), .B(n5887), .Z(n5889) );
  AND U6344 ( .A(n5890), .B(n5889), .Z(n6324) );
  NAND U6345 ( .A(n5892), .B(n5891), .Z(n5896) );
  NAND U6346 ( .A(n5894), .B(n5893), .Z(n5895) );
  NAND U6347 ( .A(n5896), .B(n5895), .Z(n6323) );
  XNOR U6348 ( .A(n6324), .B(n6323), .Z(n6326) );
  NANDN U6349 ( .A(n5898), .B(n5897), .Z(n5902) );
  NANDN U6350 ( .A(n5900), .B(n5899), .Z(n5901) );
  AND U6351 ( .A(n5902), .B(n5901), .Z(n6318) );
  NANDN U6352 ( .A(n5904), .B(n5903), .Z(n5908) );
  NANDN U6353 ( .A(n5906), .B(n5905), .Z(n5907) );
  NAND U6354 ( .A(n5908), .B(n5907), .Z(n6317) );
  XNOR U6355 ( .A(n6318), .B(n6317), .Z(n6319) );
  NANDN U6356 ( .A(n29499), .B(n5909), .Z(n5911) );
  XOR U6357 ( .A(b[7]), .B(a[44]), .Z(n6206) );
  NANDN U6358 ( .A(n29735), .B(n6206), .Z(n5910) );
  AND U6359 ( .A(n5911), .B(n5910), .Z(n6229) );
  NANDN U6360 ( .A(n28889), .B(n5912), .Z(n5914) );
  XOR U6361 ( .A(b[5]), .B(a[46]), .Z(n6146) );
  NANDN U6362 ( .A(n29138), .B(n6146), .Z(n5913) );
  AND U6363 ( .A(n5914), .B(n5913), .Z(n6228) );
  NANDN U6364 ( .A(n34634), .B(n5915), .Z(n5917) );
  XOR U6365 ( .A(b[29]), .B(a[22]), .Z(n6143) );
  NANDN U6366 ( .A(n34722), .B(n6143), .Z(n5916) );
  NAND U6367 ( .A(n5917), .B(n5916), .Z(n6227) );
  XOR U6368 ( .A(n6228), .B(n6227), .Z(n6230) );
  XOR U6369 ( .A(n6229), .B(n6230), .Z(n6288) );
  NANDN U6370 ( .A(n5919), .B(n5918), .Z(n5923) );
  NANDN U6371 ( .A(n5921), .B(n5920), .Z(n5922) );
  AND U6372 ( .A(n5923), .B(n5922), .Z(n6287) );
  XNOR U6373 ( .A(n6288), .B(n6287), .Z(n6290) );
  NANDN U6374 ( .A(n5925), .B(n5924), .Z(n5929) );
  OR U6375 ( .A(n5927), .B(n5926), .Z(n5928) );
  AND U6376 ( .A(n5929), .B(n5928), .Z(n6289) );
  XOR U6377 ( .A(n6290), .B(n6289), .Z(n6127) );
  NANDN U6378 ( .A(n34909), .B(n5930), .Z(n5932) );
  XOR U6379 ( .A(b[31]), .B(a[20]), .Z(n6188) );
  NANDN U6380 ( .A(n35145), .B(n6188), .Z(n5931) );
  AND U6381 ( .A(n5932), .B(n5931), .Z(n6157) );
  NANDN U6382 ( .A(n35936), .B(n5933), .Z(n5935) );
  XOR U6383 ( .A(b[37]), .B(a[14]), .Z(n6197) );
  NANDN U6384 ( .A(n36047), .B(n6197), .Z(n5934) );
  AND U6385 ( .A(n5935), .B(n5934), .Z(n6156) );
  NANDN U6386 ( .A(n31055), .B(n5936), .Z(n5938) );
  XOR U6387 ( .A(b[13]), .B(a[38]), .Z(n6266) );
  NANDN U6388 ( .A(n31293), .B(n6266), .Z(n5937) );
  NAND U6389 ( .A(n5938), .B(n5937), .Z(n6155) );
  XOR U6390 ( .A(n6156), .B(n6155), .Z(n6158) );
  XOR U6391 ( .A(n6157), .B(n6158), .Z(n6300) );
  XOR U6392 ( .A(b[48]), .B(b[49]), .Z(n5939) );
  ANDN U6393 ( .B(n5939), .A(n37537), .Z(n37536) );
  NANDN U6394 ( .A(n212), .B(n5940), .Z(n5942) );
  XOR U6395 ( .A(b[49]), .B(a[2]), .Z(n6177) );
  NANDN U6396 ( .A(n37432), .B(n6177), .Z(n5941) );
  AND U6397 ( .A(n5942), .B(n5941), .Z(n6133) );
  NANDN U6398 ( .A(n210), .B(n5943), .Z(n5945) );
  XOR U6399 ( .A(b[9]), .B(a[42]), .Z(n6194) );
  NANDN U6400 ( .A(n30267), .B(n6194), .Z(n5944) );
  AND U6401 ( .A(n5945), .B(n5944), .Z(n6132) );
  NANDN U6402 ( .A(n35260), .B(n5946), .Z(n5948) );
  XOR U6403 ( .A(b[33]), .B(a[18]), .Z(n6212) );
  NANDN U6404 ( .A(n35456), .B(n6212), .Z(n5947) );
  NAND U6405 ( .A(n5948), .B(n5947), .Z(n6131) );
  XOR U6406 ( .A(n6132), .B(n6131), .Z(n6134) );
  XNOR U6407 ( .A(n6133), .B(n6134), .Z(n6299) );
  XNOR U6408 ( .A(n6300), .B(n6299), .Z(n6302) );
  NANDN U6409 ( .A(n5950), .B(n5949), .Z(n5954) );
  OR U6410 ( .A(n5952), .B(n5951), .Z(n5953) );
  AND U6411 ( .A(n5954), .B(n5953), .Z(n6301) );
  XOR U6412 ( .A(n6302), .B(n6301), .Z(n6126) );
  NANDN U6413 ( .A(n5956), .B(n5955), .Z(n5960) );
  OR U6414 ( .A(n5958), .B(n5957), .Z(n5959) );
  AND U6415 ( .A(n5960), .B(n5959), .Z(n6125) );
  XOR U6416 ( .A(n6126), .B(n6125), .Z(n6128) );
  XOR U6417 ( .A(n6127), .B(n6128), .Z(n6108) );
  NANDN U6418 ( .A(n5962), .B(n5961), .Z(n5966) );
  OR U6419 ( .A(n5964), .B(n5963), .Z(n5965) );
  NAND U6420 ( .A(n5966), .B(n5965), .Z(n6107) );
  XNOR U6421 ( .A(n6108), .B(n6107), .Z(n6110) );
  NANDN U6422 ( .A(n5968), .B(n5967), .Z(n5972) );
  NANDN U6423 ( .A(n5970), .B(n5969), .Z(n5971) );
  AND U6424 ( .A(n5972), .B(n5971), .Z(n6109) );
  XOR U6425 ( .A(n6110), .B(n6109), .Z(n6314) );
  NANDN U6426 ( .A(n5974), .B(n5973), .Z(n5978) );
  OR U6427 ( .A(n5976), .B(n5975), .Z(n5977) );
  AND U6428 ( .A(n5978), .B(n5977), .Z(n6240) );
  NANDN U6429 ( .A(n5980), .B(n5979), .Z(n5984) );
  OR U6430 ( .A(n5982), .B(n5981), .Z(n5983) );
  NAND U6431 ( .A(n5984), .B(n5983), .Z(n6239) );
  XNOR U6432 ( .A(n6240), .B(n6239), .Z(n6242) );
  NANDN U6433 ( .A(n5986), .B(n5985), .Z(n5990) );
  OR U6434 ( .A(n5988), .B(n5987), .Z(n5989) );
  AND U6435 ( .A(n5990), .B(n5989), .Z(n6278) );
  XOR U6436 ( .A(b[50]), .B(b[49]), .Z(n37734) );
  IV U6437 ( .A(n37734), .Z(n37605) );
  ANDN U6438 ( .B(a[0]), .A(n37605), .Z(n6245) );
  NANDN U6439 ( .A(n211), .B(n5991), .Z(n5993) );
  XOR U6440 ( .A(b[47]), .B(a[4]), .Z(n6251) );
  NANDN U6441 ( .A(n37172), .B(n6251), .Z(n5992) );
  AND U6442 ( .A(n5993), .B(n5992), .Z(n6246) );
  XNOR U6443 ( .A(n6245), .B(n6246), .Z(n6247) );
  NAND U6444 ( .A(b[0]), .B(a[50]), .Z(n5994) );
  XNOR U6445 ( .A(b[1]), .B(n5994), .Z(n5996) );
  NANDN U6446 ( .A(b[0]), .B(a[49]), .Z(n5995) );
  NAND U6447 ( .A(n5996), .B(n5995), .Z(n6248) );
  XNOR U6448 ( .A(n6247), .B(n6248), .Z(n6275) );
  NANDN U6449 ( .A(n5997), .B(n32544), .Z(n5999) );
  XOR U6450 ( .A(b[17]), .B(a[34]), .Z(n6260) );
  NANDN U6451 ( .A(n32292), .B(n6260), .Z(n5998) );
  AND U6452 ( .A(n5999), .B(n5998), .Z(n6164) );
  NANDN U6453 ( .A(n32483), .B(n6000), .Z(n6002) );
  XOR U6454 ( .A(b[19]), .B(a[32]), .Z(n6203) );
  NANDN U6455 ( .A(n32823), .B(n6203), .Z(n6001) );
  AND U6456 ( .A(n6002), .B(n6001), .Z(n6162) );
  NANDN U6457 ( .A(n32996), .B(n6003), .Z(n6005) );
  XOR U6458 ( .A(b[21]), .B(a[30]), .Z(n6269) );
  NANDN U6459 ( .A(n33271), .B(n6269), .Z(n6004) );
  NAND U6460 ( .A(n6005), .B(n6004), .Z(n6161) );
  XNOR U6461 ( .A(n6162), .B(n6161), .Z(n6163) );
  XOR U6462 ( .A(n6164), .B(n6163), .Z(n6276) );
  XNOR U6463 ( .A(n6275), .B(n6276), .Z(n6277) );
  XNOR U6464 ( .A(n6278), .B(n6277), .Z(n6241) );
  XOR U6465 ( .A(n6242), .B(n6241), .Z(n6307) );
  NANDN U6466 ( .A(n6007), .B(n6006), .Z(n6011) );
  OR U6467 ( .A(n6009), .B(n6008), .Z(n6010) );
  AND U6468 ( .A(n6011), .B(n6010), .Z(n6235) );
  NANDN U6469 ( .A(n209), .B(n6012), .Z(n6014) );
  XOR U6470 ( .A(b[3]), .B(a[48]), .Z(n6149) );
  NANDN U6471 ( .A(n28941), .B(n6149), .Z(n6013) );
  AND U6472 ( .A(n6014), .B(n6013), .Z(n6168) );
  NANDN U6473 ( .A(n34223), .B(n6015), .Z(n6017) );
  XOR U6474 ( .A(b[27]), .B(a[24]), .Z(n6185) );
  NANDN U6475 ( .A(n34458), .B(n6185), .Z(n6016) );
  NAND U6476 ( .A(n6017), .B(n6016), .Z(n6167) );
  XNOR U6477 ( .A(n6168), .B(n6167), .Z(n6170) );
  ANDN U6478 ( .B(n6019), .A(n6018), .Z(n6169) );
  XOR U6479 ( .A(n6170), .B(n6169), .Z(n6233) );
  NANDN U6480 ( .A(n33866), .B(n6020), .Z(n6022) );
  XOR U6481 ( .A(b[23]), .B(a[28]), .Z(n6152) );
  NANDN U6482 ( .A(n33644), .B(n6152), .Z(n6021) );
  AND U6483 ( .A(n6022), .B(n6021), .Z(n6218) );
  NANDN U6484 ( .A(n33875), .B(n6023), .Z(n6025) );
  XOR U6485 ( .A(b[25]), .B(a[26]), .Z(n6257) );
  NANDN U6486 ( .A(n33994), .B(n6257), .Z(n6024) );
  AND U6487 ( .A(n6025), .B(n6024), .Z(n6216) );
  NANDN U6488 ( .A(n31536), .B(n6026), .Z(n6028) );
  XOR U6489 ( .A(b[15]), .B(a[36]), .Z(n6263) );
  NANDN U6490 ( .A(n31925), .B(n6263), .Z(n6027) );
  NAND U6491 ( .A(n6028), .B(n6027), .Z(n6215) );
  XNOR U6492 ( .A(n6216), .B(n6215), .Z(n6217) );
  XOR U6493 ( .A(n6218), .B(n6217), .Z(n6234) );
  XOR U6494 ( .A(n6233), .B(n6234), .Z(n6236) );
  XOR U6495 ( .A(n6235), .B(n6236), .Z(n6306) );
  NANDN U6496 ( .A(n36991), .B(n6029), .Z(n6031) );
  XOR U6497 ( .A(b[45]), .B(a[6]), .Z(n6140) );
  NANDN U6498 ( .A(n37083), .B(n6140), .Z(n6030) );
  AND U6499 ( .A(n6031), .B(n6030), .Z(n6223) );
  NANDN U6500 ( .A(n30482), .B(n6032), .Z(n6034) );
  XOR U6501 ( .A(b[11]), .B(a[40]), .Z(n6272) );
  NANDN U6502 ( .A(n30891), .B(n6272), .Z(n6033) );
  AND U6503 ( .A(n6034), .B(n6033), .Z(n6222) );
  NANDN U6504 ( .A(n35611), .B(n6035), .Z(n6037) );
  XOR U6505 ( .A(b[35]), .B(a[16]), .Z(n6191) );
  NANDN U6506 ( .A(n35801), .B(n6191), .Z(n6036) );
  NAND U6507 ( .A(n6037), .B(n6036), .Z(n6221) );
  XOR U6508 ( .A(n6222), .B(n6221), .Z(n6224) );
  XOR U6509 ( .A(n6223), .B(n6224), .Z(n6294) );
  NANDN U6510 ( .A(n36210), .B(n6038), .Z(n6040) );
  XOR U6511 ( .A(b[39]), .B(a[12]), .Z(n6200) );
  NANDN U6512 ( .A(n36347), .B(n6200), .Z(n6039) );
  AND U6513 ( .A(n6040), .B(n6039), .Z(n6173) );
  NANDN U6514 ( .A(n36480), .B(n6041), .Z(n6043) );
  XOR U6515 ( .A(b[41]), .B(a[10]), .Z(n6209) );
  NANDN U6516 ( .A(n36594), .B(n6209), .Z(n6042) );
  AND U6517 ( .A(n6043), .B(n6042), .Z(n6172) );
  NANDN U6518 ( .A(n36742), .B(n6044), .Z(n6046) );
  XOR U6519 ( .A(b[43]), .B(a[8]), .Z(n6137) );
  NANDN U6520 ( .A(n36891), .B(n6137), .Z(n6045) );
  NAND U6521 ( .A(n6046), .B(n6045), .Z(n6171) );
  XOR U6522 ( .A(n6172), .B(n6171), .Z(n6174) );
  XNOR U6523 ( .A(n6173), .B(n6174), .Z(n6293) );
  XNOR U6524 ( .A(n6294), .B(n6293), .Z(n6295) );
  NANDN U6525 ( .A(n6048), .B(n6047), .Z(n6052) );
  NANDN U6526 ( .A(n6050), .B(n6049), .Z(n6051) );
  NAND U6527 ( .A(n6052), .B(n6051), .Z(n6296) );
  XNOR U6528 ( .A(n6295), .B(n6296), .Z(n6305) );
  XOR U6529 ( .A(n6306), .B(n6305), .Z(n6308) );
  XOR U6530 ( .A(n6307), .B(n6308), .Z(n6283) );
  NANDN U6531 ( .A(n6054), .B(n6053), .Z(n6058) );
  OR U6532 ( .A(n6056), .B(n6055), .Z(n6057) );
  AND U6533 ( .A(n6058), .B(n6057), .Z(n6282) );
  NANDN U6534 ( .A(n6060), .B(n6059), .Z(n6064) );
  NANDN U6535 ( .A(n6062), .B(n6061), .Z(n6063) );
  AND U6536 ( .A(n6064), .B(n6063), .Z(n6281) );
  XOR U6537 ( .A(n6282), .B(n6281), .Z(n6284) );
  XOR U6538 ( .A(n6283), .B(n6284), .Z(n6120) );
  NANDN U6539 ( .A(n6066), .B(n6065), .Z(n6070) );
  NAND U6540 ( .A(n6068), .B(n6067), .Z(n6069) );
  NAND U6541 ( .A(n6070), .B(n6069), .Z(n6119) );
  XNOR U6542 ( .A(n6120), .B(n6119), .Z(n6122) );
  NANDN U6543 ( .A(n6072), .B(n6071), .Z(n6076) );
  NANDN U6544 ( .A(n6074), .B(n6073), .Z(n6075) );
  NAND U6545 ( .A(n6076), .B(n6075), .Z(n6113) );
  NANDN U6546 ( .A(n6078), .B(n6077), .Z(n6082) );
  NANDN U6547 ( .A(n6080), .B(n6079), .Z(n6081) );
  AND U6548 ( .A(n6082), .B(n6081), .Z(n6114) );
  XOR U6549 ( .A(n6113), .B(n6114), .Z(n6116) );
  NANDN U6550 ( .A(n6084), .B(n6083), .Z(n6088) );
  OR U6551 ( .A(n6086), .B(n6085), .Z(n6087) );
  AND U6552 ( .A(n6088), .B(n6087), .Z(n6115) );
  XOR U6553 ( .A(n6116), .B(n6115), .Z(n6121) );
  XOR U6554 ( .A(n6122), .B(n6121), .Z(n6312) );
  NANDN U6555 ( .A(n6090), .B(n6089), .Z(n6094) );
  NAND U6556 ( .A(n6092), .B(n6091), .Z(n6093) );
  AND U6557 ( .A(n6094), .B(n6093), .Z(n6311) );
  XNOR U6558 ( .A(n6312), .B(n6311), .Z(n6313) );
  XOR U6559 ( .A(n6314), .B(n6313), .Z(n6320) );
  XNOR U6560 ( .A(n6319), .B(n6320), .Z(n6325) );
  XOR U6561 ( .A(n6326), .B(n6325), .Z(n6102) );
  NANDN U6562 ( .A(n6096), .B(n6095), .Z(n6100) );
  OR U6563 ( .A(n6098), .B(n6097), .Z(n6099) );
  AND U6564 ( .A(n6100), .B(n6099), .Z(n6101) );
  XNOR U6565 ( .A(n6102), .B(n6101), .Z(n6103) );
  XNOR U6566 ( .A(n6104), .B(n6103), .Z(n6330) );
  XNOR U6567 ( .A(n6331), .B(n6330), .Z(c[114]) );
  NANDN U6568 ( .A(n6102), .B(n6101), .Z(n6106) );
  NANDN U6569 ( .A(n6104), .B(n6103), .Z(n6105) );
  AND U6570 ( .A(n6106), .B(n6105), .Z(n6342) );
  NANDN U6571 ( .A(n6108), .B(n6107), .Z(n6112) );
  NAND U6572 ( .A(n6110), .B(n6109), .Z(n6111) );
  AND U6573 ( .A(n6112), .B(n6111), .Z(n6562) );
  NAND U6574 ( .A(n6114), .B(n6113), .Z(n6118) );
  NAND U6575 ( .A(n6116), .B(n6115), .Z(n6117) );
  NAND U6576 ( .A(n6118), .B(n6117), .Z(n6563) );
  XNOR U6577 ( .A(n6562), .B(n6563), .Z(n6565) );
  NANDN U6578 ( .A(n6120), .B(n6119), .Z(n6124) );
  NAND U6579 ( .A(n6122), .B(n6121), .Z(n6123) );
  AND U6580 ( .A(n6124), .B(n6123), .Z(n6558) );
  NANDN U6581 ( .A(n6126), .B(n6125), .Z(n6130) );
  OR U6582 ( .A(n6128), .B(n6127), .Z(n6129) );
  AND U6583 ( .A(n6130), .B(n6129), .Z(n6354) );
  NANDN U6584 ( .A(n6132), .B(n6131), .Z(n6136) );
  OR U6585 ( .A(n6134), .B(n6133), .Z(n6135) );
  AND U6586 ( .A(n6136), .B(n6135), .Z(n6459) );
  NAND U6587 ( .A(n36962), .B(n6137), .Z(n6139) );
  XNOR U6588 ( .A(b[43]), .B(a[9]), .Z(n6476) );
  NANDN U6589 ( .A(n6476), .B(n36963), .Z(n6138) );
  NAND U6590 ( .A(n6139), .B(n6138), .Z(n6399) );
  NAND U6591 ( .A(n37202), .B(n6140), .Z(n6142) );
  XNOR U6592 ( .A(b[45]), .B(a[7]), .Z(n6505) );
  NANDN U6593 ( .A(n6505), .B(n37200), .Z(n6141) );
  NAND U6594 ( .A(n6142), .B(n6141), .Z(n6398) );
  NAND U6595 ( .A(n35001), .B(n6143), .Z(n6145) );
  XNOR U6596 ( .A(b[29]), .B(a[23]), .Z(n6500) );
  NANDN U6597 ( .A(n6500), .B(n35002), .Z(n6144) );
  NAND U6598 ( .A(n6145), .B(n6144), .Z(n6397) );
  XOR U6599 ( .A(n6398), .B(n6397), .Z(n6400) );
  XNOR U6600 ( .A(n6399), .B(n6400), .Z(n6410) );
  NANDN U6601 ( .A(n28889), .B(n6146), .Z(n6148) );
  XOR U6602 ( .A(b[5]), .B(a[47]), .Z(n6387) );
  NANDN U6603 ( .A(n29138), .B(n6387), .Z(n6147) );
  AND U6604 ( .A(n6148), .B(n6147), .Z(n6438) );
  NANDN U6605 ( .A(n209), .B(n6149), .Z(n6151) );
  XOR U6606 ( .A(b[3]), .B(a[49]), .Z(n6497) );
  NANDN U6607 ( .A(n28941), .B(n6497), .Z(n6150) );
  AND U6608 ( .A(n6151), .B(n6150), .Z(n6437) );
  NANDN U6609 ( .A(n33866), .B(n6152), .Z(n6154) );
  XOR U6610 ( .A(b[23]), .B(a[29]), .Z(n6424) );
  NANDN U6611 ( .A(n33644), .B(n6424), .Z(n6153) );
  NAND U6612 ( .A(n6154), .B(n6153), .Z(n6436) );
  XOR U6613 ( .A(n6437), .B(n6436), .Z(n6439) );
  XNOR U6614 ( .A(n6438), .B(n6439), .Z(n6409) );
  XOR U6615 ( .A(n6410), .B(n6409), .Z(n6412) );
  NANDN U6616 ( .A(n6156), .B(n6155), .Z(n6160) );
  OR U6617 ( .A(n6158), .B(n6157), .Z(n6159) );
  AND U6618 ( .A(n6160), .B(n6159), .Z(n6411) );
  XNOR U6619 ( .A(n6412), .B(n6411), .Z(n6458) );
  XNOR U6620 ( .A(n6459), .B(n6458), .Z(n6461) );
  NANDN U6621 ( .A(n6162), .B(n6161), .Z(n6166) );
  NANDN U6622 ( .A(n6164), .B(n6163), .Z(n6165) );
  AND U6623 ( .A(n6166), .B(n6165), .Z(n6449) );
  XNOR U6624 ( .A(n6449), .B(n6448), .Z(n6451) );
  NANDN U6625 ( .A(n6172), .B(n6171), .Z(n6176) );
  OR U6626 ( .A(n6174), .B(n6173), .Z(n6175) );
  NAND U6627 ( .A(n6176), .B(n6175), .Z(n6365) );
  NANDN U6628 ( .A(n212), .B(n6177), .Z(n6179) );
  XOR U6629 ( .A(b[49]), .B(a[3]), .Z(n6384) );
  NANDN U6630 ( .A(n37432), .B(n6384), .Z(n6178) );
  AND U6631 ( .A(n6179), .B(n6178), .Z(n6503) );
  XOR U6632 ( .A(b[51]), .B(b[50]), .Z(n6390) );
  XOR U6633 ( .A(b[51]), .B(a[0]), .Z(n6180) );
  NAND U6634 ( .A(n6390), .B(n6180), .Z(n6181) );
  OR U6635 ( .A(n6181), .B(n37734), .Z(n6183) );
  XOR U6636 ( .A(b[51]), .B(a[1]), .Z(n6391) );
  NAND U6637 ( .A(n37734), .B(n6391), .Z(n6182) );
  AND U6638 ( .A(n6183), .B(n6182), .Z(n6504) );
  XOR U6639 ( .A(n6503), .B(n6504), .Z(n6473) );
  NAND U6640 ( .A(b[49]), .B(b[50]), .Z(n6184) );
  NAND U6641 ( .A(b[51]), .B(n6184), .Z(n37831) );
  NOR U6642 ( .A(n37831), .B(n6245), .Z(n6471) );
  NAND U6643 ( .A(n34647), .B(n6185), .Z(n6187) );
  XNOR U6644 ( .A(b[27]), .B(a[25]), .Z(n6511) );
  NANDN U6645 ( .A(n6511), .B(n34648), .Z(n6186) );
  AND U6646 ( .A(n6187), .B(n6186), .Z(n6470) );
  XNOR U6647 ( .A(n6471), .B(n6470), .Z(n6472) );
  XOR U6648 ( .A(n6473), .B(n6472), .Z(n6363) );
  NANDN U6649 ( .A(n34909), .B(n6188), .Z(n6190) );
  XOR U6650 ( .A(b[31]), .B(a[21]), .Z(n6394) );
  NANDN U6651 ( .A(n35145), .B(n6394), .Z(n6189) );
  AND U6652 ( .A(n6190), .B(n6189), .Z(n6488) );
  NANDN U6653 ( .A(n35611), .B(n6191), .Z(n6193) );
  XOR U6654 ( .A(b[35]), .B(a[17]), .Z(n6418) );
  NANDN U6655 ( .A(n35801), .B(n6418), .Z(n6192) );
  AND U6656 ( .A(n6193), .B(n6192), .Z(n6486) );
  NANDN U6657 ( .A(n210), .B(n6194), .Z(n6196) );
  XOR U6658 ( .A(b[9]), .B(a[43]), .Z(n6532) );
  NANDN U6659 ( .A(n30267), .B(n6532), .Z(n6195) );
  NAND U6660 ( .A(n6196), .B(n6195), .Z(n6485) );
  XNOR U6661 ( .A(n6486), .B(n6485), .Z(n6487) );
  XNOR U6662 ( .A(n6488), .B(n6487), .Z(n6364) );
  XOR U6663 ( .A(n6363), .B(n6364), .Z(n6366) );
  XOR U6664 ( .A(n6365), .B(n6366), .Z(n6450) );
  XOR U6665 ( .A(n6451), .B(n6450), .Z(n6460) );
  XOR U6666 ( .A(n6461), .B(n6460), .Z(n6546) );
  NANDN U6667 ( .A(n35936), .B(n6197), .Z(n6199) );
  XOR U6668 ( .A(b[37]), .B(a[15]), .Z(n6520) );
  NANDN U6669 ( .A(n36047), .B(n6520), .Z(n6198) );
  AND U6670 ( .A(n6199), .B(n6198), .Z(n6516) );
  NANDN U6671 ( .A(n36210), .B(n6200), .Z(n6202) );
  XOR U6672 ( .A(b[39]), .B(a[13]), .Z(n6535) );
  NANDN U6673 ( .A(n36347), .B(n6535), .Z(n6201) );
  AND U6674 ( .A(n6202), .B(n6201), .Z(n6515) );
  NANDN U6675 ( .A(n32483), .B(n6203), .Z(n6205) );
  XOR U6676 ( .A(b[19]), .B(a[33]), .Z(n6433) );
  NANDN U6677 ( .A(n32823), .B(n6433), .Z(n6204) );
  NAND U6678 ( .A(n6205), .B(n6204), .Z(n6514) );
  XOR U6679 ( .A(n6515), .B(n6514), .Z(n6517) );
  XOR U6680 ( .A(n6516), .B(n6517), .Z(n6358) );
  NANDN U6681 ( .A(n29499), .B(n6206), .Z(n6208) );
  XOR U6682 ( .A(b[7]), .B(a[45]), .Z(n6479) );
  NANDN U6683 ( .A(n29735), .B(n6479), .Z(n6207) );
  AND U6684 ( .A(n6208), .B(n6207), .Z(n6493) );
  NANDN U6685 ( .A(n36480), .B(n6209), .Z(n6211) );
  XOR U6686 ( .A(b[41]), .B(a[11]), .Z(n6523) );
  NANDN U6687 ( .A(n36594), .B(n6523), .Z(n6210) );
  AND U6688 ( .A(n6211), .B(n6210), .Z(n6492) );
  NANDN U6689 ( .A(n35260), .B(n6212), .Z(n6214) );
  XOR U6690 ( .A(b[33]), .B(a[19]), .Z(n6415) );
  NANDN U6691 ( .A(n35456), .B(n6415), .Z(n6213) );
  NAND U6692 ( .A(n6214), .B(n6213), .Z(n6491) );
  XOR U6693 ( .A(n6492), .B(n6491), .Z(n6494) );
  XNOR U6694 ( .A(n6493), .B(n6494), .Z(n6357) );
  XNOR U6695 ( .A(n6358), .B(n6357), .Z(n6360) );
  NANDN U6696 ( .A(n6216), .B(n6215), .Z(n6220) );
  NANDN U6697 ( .A(n6218), .B(n6217), .Z(n6219) );
  AND U6698 ( .A(n6220), .B(n6219), .Z(n6359) );
  XOR U6699 ( .A(n6360), .B(n6359), .Z(n6371) );
  NANDN U6700 ( .A(n6222), .B(n6221), .Z(n6226) );
  OR U6701 ( .A(n6224), .B(n6223), .Z(n6225) );
  AND U6702 ( .A(n6226), .B(n6225), .Z(n6370) );
  NANDN U6703 ( .A(n6228), .B(n6227), .Z(n6232) );
  OR U6704 ( .A(n6230), .B(n6229), .Z(n6231) );
  NAND U6705 ( .A(n6232), .B(n6231), .Z(n6369) );
  XOR U6706 ( .A(n6370), .B(n6369), .Z(n6372) );
  XOR U6707 ( .A(n6371), .B(n6372), .Z(n6545) );
  NANDN U6708 ( .A(n6234), .B(n6233), .Z(n6238) );
  OR U6709 ( .A(n6236), .B(n6235), .Z(n6237) );
  AND U6710 ( .A(n6238), .B(n6237), .Z(n6544) );
  XOR U6711 ( .A(n6545), .B(n6544), .Z(n6547) );
  XOR U6712 ( .A(n6546), .B(n6547), .Z(n6352) );
  NANDN U6713 ( .A(n6240), .B(n6239), .Z(n6244) );
  NAND U6714 ( .A(n6242), .B(n6241), .Z(n6243) );
  AND U6715 ( .A(n6244), .B(n6243), .Z(n6455) );
  NANDN U6716 ( .A(n6246), .B(n6245), .Z(n6250) );
  NANDN U6717 ( .A(n6248), .B(n6247), .Z(n6249) );
  AND U6718 ( .A(n6250), .B(n6249), .Z(n6465) );
  NANDN U6719 ( .A(n211), .B(n6251), .Z(n6253) );
  XOR U6720 ( .A(b[47]), .B(a[5]), .Z(n6508) );
  NANDN U6721 ( .A(n37172), .B(n6508), .Z(n6252) );
  AND U6722 ( .A(n6253), .B(n6252), .Z(n6445) );
  NAND U6723 ( .A(b[0]), .B(a[51]), .Z(n6254) );
  XNOR U6724 ( .A(b[1]), .B(n6254), .Z(n6256) );
  NANDN U6725 ( .A(b[0]), .B(a[50]), .Z(n6255) );
  NAND U6726 ( .A(n6256), .B(n6255), .Z(n6443) );
  NANDN U6727 ( .A(n33875), .B(n6257), .Z(n6259) );
  XOR U6728 ( .A(b[25]), .B(a[27]), .Z(n6482) );
  NANDN U6729 ( .A(n33994), .B(n6482), .Z(n6258) );
  NAND U6730 ( .A(n6259), .B(n6258), .Z(n6442) );
  XNOR U6731 ( .A(n6443), .B(n6442), .Z(n6444) );
  XNOR U6732 ( .A(n6445), .B(n6444), .Z(n6464) );
  XNOR U6733 ( .A(n6465), .B(n6464), .Z(n6467) );
  NANDN U6734 ( .A(n32013), .B(n6260), .Z(n6262) );
  XOR U6735 ( .A(b[17]), .B(a[35]), .Z(n6427) );
  NANDN U6736 ( .A(n32292), .B(n6427), .Z(n6261) );
  AND U6737 ( .A(n6262), .B(n6261), .Z(n6406) );
  NANDN U6738 ( .A(n31536), .B(n6263), .Z(n6265) );
  XOR U6739 ( .A(b[15]), .B(a[37]), .Z(n6421) );
  NANDN U6740 ( .A(n31925), .B(n6421), .Z(n6264) );
  AND U6741 ( .A(n6265), .B(n6264), .Z(n6404) );
  NANDN U6742 ( .A(n31055), .B(n6266), .Z(n6268) );
  XOR U6743 ( .A(b[13]), .B(a[39]), .Z(n6526) );
  NANDN U6744 ( .A(n31293), .B(n6526), .Z(n6267) );
  AND U6745 ( .A(n6268), .B(n6267), .Z(n6378) );
  NANDN U6746 ( .A(n32996), .B(n6269), .Z(n6271) );
  XOR U6747 ( .A(b[21]), .B(a[31]), .Z(n6430) );
  NANDN U6748 ( .A(n33271), .B(n6430), .Z(n6270) );
  AND U6749 ( .A(n6271), .B(n6270), .Z(n6376) );
  NANDN U6750 ( .A(n30482), .B(n6272), .Z(n6274) );
  XOR U6751 ( .A(b[11]), .B(a[41]), .Z(n6529) );
  NANDN U6752 ( .A(n30891), .B(n6529), .Z(n6273) );
  NAND U6753 ( .A(n6274), .B(n6273), .Z(n6375) );
  XNOR U6754 ( .A(n6376), .B(n6375), .Z(n6377) );
  XNOR U6755 ( .A(n6378), .B(n6377), .Z(n6403) );
  XNOR U6756 ( .A(n6404), .B(n6403), .Z(n6405) );
  XNOR U6757 ( .A(n6406), .B(n6405), .Z(n6466) );
  XOR U6758 ( .A(n6467), .B(n6466), .Z(n6453) );
  NANDN U6759 ( .A(n6276), .B(n6275), .Z(n6280) );
  NANDN U6760 ( .A(n6278), .B(n6277), .Z(n6279) );
  AND U6761 ( .A(n6280), .B(n6279), .Z(n6452) );
  XNOR U6762 ( .A(n6453), .B(n6452), .Z(n6454) );
  XNOR U6763 ( .A(n6455), .B(n6454), .Z(n6351) );
  XNOR U6764 ( .A(n6352), .B(n6351), .Z(n6353) );
  XNOR U6765 ( .A(n6354), .B(n6353), .Z(n6556) );
  NANDN U6766 ( .A(n6282), .B(n6281), .Z(n6286) );
  OR U6767 ( .A(n6284), .B(n6283), .Z(n6285) );
  AND U6768 ( .A(n6286), .B(n6285), .Z(n6541) );
  NANDN U6769 ( .A(n6288), .B(n6287), .Z(n6292) );
  NAND U6770 ( .A(n6290), .B(n6289), .Z(n6291) );
  AND U6771 ( .A(n6292), .B(n6291), .Z(n6552) );
  NANDN U6772 ( .A(n6294), .B(n6293), .Z(n6298) );
  NANDN U6773 ( .A(n6296), .B(n6295), .Z(n6297) );
  AND U6774 ( .A(n6298), .B(n6297), .Z(n6551) );
  NANDN U6775 ( .A(n6300), .B(n6299), .Z(n6304) );
  NAND U6776 ( .A(n6302), .B(n6301), .Z(n6303) );
  NAND U6777 ( .A(n6304), .B(n6303), .Z(n6550) );
  XOR U6778 ( .A(n6551), .B(n6550), .Z(n6553) );
  XOR U6779 ( .A(n6552), .B(n6553), .Z(n6539) );
  NANDN U6780 ( .A(n6306), .B(n6305), .Z(n6310) );
  OR U6781 ( .A(n6308), .B(n6307), .Z(n6309) );
  AND U6782 ( .A(n6310), .B(n6309), .Z(n6538) );
  XNOR U6783 ( .A(n6539), .B(n6538), .Z(n6540) );
  XOR U6784 ( .A(n6541), .B(n6540), .Z(n6557) );
  XOR U6785 ( .A(n6556), .B(n6557), .Z(n6559) );
  XNOR U6786 ( .A(n6558), .B(n6559), .Z(n6564) );
  XOR U6787 ( .A(n6565), .B(n6564), .Z(n6346) );
  NANDN U6788 ( .A(n6312), .B(n6311), .Z(n6316) );
  NANDN U6789 ( .A(n6314), .B(n6313), .Z(n6315) );
  AND U6790 ( .A(n6316), .B(n6315), .Z(n6345) );
  XNOR U6791 ( .A(n6346), .B(n6345), .Z(n6347) );
  NANDN U6792 ( .A(n6318), .B(n6317), .Z(n6322) );
  NANDN U6793 ( .A(n6320), .B(n6319), .Z(n6321) );
  NAND U6794 ( .A(n6322), .B(n6321), .Z(n6348) );
  XNOR U6795 ( .A(n6347), .B(n6348), .Z(n6339) );
  NANDN U6796 ( .A(n6324), .B(n6323), .Z(n6328) );
  NAND U6797 ( .A(n6326), .B(n6325), .Z(n6327) );
  NAND U6798 ( .A(n6328), .B(n6327), .Z(n6340) );
  XNOR U6799 ( .A(n6339), .B(n6340), .Z(n6341) );
  XNOR U6800 ( .A(n6342), .B(n6341), .Z(n6334) );
  XNOR U6801 ( .A(sreg[115]), .B(n6334), .Z(n6336) );
  NANDN U6802 ( .A(sreg[114]), .B(n6329), .Z(n6333) );
  NAND U6803 ( .A(n6331), .B(n6330), .Z(n6332) );
  NAND U6804 ( .A(n6333), .B(n6332), .Z(n6335) );
  XNOR U6805 ( .A(n6336), .B(n6335), .Z(c[115]) );
  NANDN U6806 ( .A(sreg[115]), .B(n6334), .Z(n6338) );
  NAND U6807 ( .A(n6336), .B(n6335), .Z(n6337) );
  NAND U6808 ( .A(n6338), .B(n6337), .Z(n6568) );
  XNOR U6809 ( .A(sreg[116]), .B(n6568), .Z(n6570) );
  NANDN U6810 ( .A(n6340), .B(n6339), .Z(n6344) );
  NANDN U6811 ( .A(n6342), .B(n6341), .Z(n6343) );
  AND U6812 ( .A(n6344), .B(n6343), .Z(n6575) );
  NANDN U6813 ( .A(n6346), .B(n6345), .Z(n6350) );
  NANDN U6814 ( .A(n6348), .B(n6347), .Z(n6349) );
  AND U6815 ( .A(n6350), .B(n6349), .Z(n6574) );
  NANDN U6816 ( .A(n6352), .B(n6351), .Z(n6356) );
  NANDN U6817 ( .A(n6354), .B(n6353), .Z(n6355) );
  AND U6818 ( .A(n6356), .B(n6355), .Z(n6801) );
  NANDN U6819 ( .A(n6358), .B(n6357), .Z(n6362) );
  NAND U6820 ( .A(n6360), .B(n6359), .Z(n6361) );
  AND U6821 ( .A(n6362), .B(n6361), .Z(n6580) );
  NAND U6822 ( .A(n6364), .B(n6363), .Z(n6368) );
  NAND U6823 ( .A(n6366), .B(n6365), .Z(n6367) );
  AND U6824 ( .A(n6368), .B(n6367), .Z(n6579) );
  XNOR U6825 ( .A(n6580), .B(n6579), .Z(n6581) );
  NANDN U6826 ( .A(n6370), .B(n6369), .Z(n6374) );
  OR U6827 ( .A(n6372), .B(n6371), .Z(n6373) );
  NAND U6828 ( .A(n6374), .B(n6373), .Z(n6582) );
  XNOR U6829 ( .A(n6581), .B(n6582), .Z(n6791) );
  NANDN U6830 ( .A(n6376), .B(n6375), .Z(n6380) );
  NANDN U6831 ( .A(n6378), .B(n6377), .Z(n6379) );
  AND U6832 ( .A(n6380), .B(n6379), .Z(n6673) );
  NAND U6833 ( .A(b[0]), .B(a[52]), .Z(n6381) );
  XNOR U6834 ( .A(b[1]), .B(n6381), .Z(n6383) );
  NANDN U6835 ( .A(b[0]), .B(a[51]), .Z(n6382) );
  NAND U6836 ( .A(n6383), .B(n6382), .Z(n6596) );
  XOR U6837 ( .A(b[52]), .B(b[51]), .Z(n37850) );
  IV U6838 ( .A(n37850), .Z(n37778) );
  ANDN U6839 ( .B(a[0]), .A(n37778), .Z(n6723) );
  NANDN U6840 ( .A(n212), .B(n6384), .Z(n6386) );
  XOR U6841 ( .A(b[49]), .B(a[4]), .Z(n6689) );
  NANDN U6842 ( .A(n37432), .B(n6689), .Z(n6385) );
  AND U6843 ( .A(n6386), .B(n6385), .Z(n6594) );
  XNOR U6844 ( .A(n6723), .B(n6594), .Z(n6595) );
  XNOR U6845 ( .A(n6596), .B(n6595), .Z(n6671) );
  NANDN U6846 ( .A(n28889), .B(n6387), .Z(n6389) );
  XOR U6847 ( .A(b[5]), .B(a[48]), .Z(n6588) );
  NANDN U6848 ( .A(n29138), .B(n6588), .Z(n6388) );
  AND U6849 ( .A(n6389), .B(n6388), .Z(n6743) );
  ANDN U6850 ( .B(n6390), .A(n37734), .Z(n37733) );
  IV U6851 ( .A(n37733), .Z(n37526) );
  NANDN U6852 ( .A(n37526), .B(n6391), .Z(n6393) );
  XOR U6853 ( .A(b[51]), .B(a[2]), .Z(n6724) );
  NANDN U6854 ( .A(n37605), .B(n6724), .Z(n6392) );
  AND U6855 ( .A(n6393), .B(n6392), .Z(n6741) );
  NANDN U6856 ( .A(n34909), .B(n6394), .Z(n6396) );
  XOR U6857 ( .A(b[31]), .B(a[22]), .Z(n6761) );
  NANDN U6858 ( .A(n35145), .B(n6761), .Z(n6395) );
  NAND U6859 ( .A(n6396), .B(n6395), .Z(n6740) );
  XNOR U6860 ( .A(n6741), .B(n6740), .Z(n6742) );
  XOR U6861 ( .A(n6743), .B(n6742), .Z(n6672) );
  XOR U6862 ( .A(n6671), .B(n6672), .Z(n6674) );
  XOR U6863 ( .A(n6673), .B(n6674), .Z(n6638) );
  NAND U6864 ( .A(n6398), .B(n6397), .Z(n6402) );
  NAND U6865 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U6866 ( .A(n6402), .B(n6401), .Z(n6635) );
  NANDN U6867 ( .A(n6404), .B(n6403), .Z(n6408) );
  NANDN U6868 ( .A(n6406), .B(n6405), .Z(n6407) );
  NAND U6869 ( .A(n6408), .B(n6407), .Z(n6636) );
  XNOR U6870 ( .A(n6635), .B(n6636), .Z(n6637) );
  XNOR U6871 ( .A(n6638), .B(n6637), .Z(n6788) );
  NAND U6872 ( .A(n6410), .B(n6409), .Z(n6414) );
  NAND U6873 ( .A(n6412), .B(n6411), .Z(n6413) );
  AND U6874 ( .A(n6414), .B(n6413), .Z(n6648) );
  NANDN U6875 ( .A(n35260), .B(n6415), .Z(n6417) );
  XOR U6876 ( .A(b[33]), .B(a[20]), .Z(n6617) );
  NANDN U6877 ( .A(n35456), .B(n6617), .Z(n6416) );
  AND U6878 ( .A(n6417), .B(n6416), .Z(n6715) );
  NANDN U6879 ( .A(n35611), .B(n6418), .Z(n6420) );
  XOR U6880 ( .A(b[35]), .B(a[18]), .Z(n6585) );
  NANDN U6881 ( .A(n35801), .B(n6585), .Z(n6419) );
  AND U6882 ( .A(n6420), .B(n6419), .Z(n6714) );
  NANDN U6883 ( .A(n31536), .B(n6421), .Z(n6423) );
  XOR U6884 ( .A(b[15]), .B(a[38]), .Z(n6737) );
  NANDN U6885 ( .A(n31925), .B(n6737), .Z(n6422) );
  NAND U6886 ( .A(n6423), .B(n6422), .Z(n6713) );
  XOR U6887 ( .A(n6714), .B(n6713), .Z(n6716) );
  XOR U6888 ( .A(n6715), .B(n6716), .Z(n6631) );
  NANDN U6889 ( .A(n33866), .B(n6424), .Z(n6426) );
  XOR U6890 ( .A(b[23]), .B(a[30]), .Z(n6752) );
  NANDN U6891 ( .A(n33644), .B(n6752), .Z(n6425) );
  AND U6892 ( .A(n6426), .B(n6425), .Z(n6697) );
  NANDN U6893 ( .A(n32013), .B(n6427), .Z(n6429) );
  XOR U6894 ( .A(b[17]), .B(a[36]), .Z(n6605) );
  NANDN U6895 ( .A(n32292), .B(n6605), .Z(n6428) );
  AND U6896 ( .A(n6429), .B(n6428), .Z(n6696) );
  NANDN U6897 ( .A(n32996), .B(n6430), .Z(n6432) );
  XOR U6898 ( .A(b[21]), .B(a[32]), .Z(n6614) );
  NANDN U6899 ( .A(n33271), .B(n6614), .Z(n6431) );
  NAND U6900 ( .A(n6432), .B(n6431), .Z(n6695) );
  XOR U6901 ( .A(n6696), .B(n6695), .Z(n6698) );
  XOR U6902 ( .A(n6697), .B(n6698), .Z(n6630) );
  NAND U6903 ( .A(n33000), .B(n6433), .Z(n6435) );
  XNOR U6904 ( .A(b[19]), .B(a[34]), .Z(n6608) );
  NANDN U6905 ( .A(n6608), .B(n33001), .Z(n6434) );
  AND U6906 ( .A(n6435), .B(n6434), .Z(n6629) );
  XOR U6907 ( .A(n6630), .B(n6629), .Z(n6632) );
  XOR U6908 ( .A(n6631), .B(n6632), .Z(n6655) );
  NANDN U6909 ( .A(n6437), .B(n6436), .Z(n6441) );
  OR U6910 ( .A(n6439), .B(n6438), .Z(n6440) );
  AND U6911 ( .A(n6441), .B(n6440), .Z(n6654) );
  NANDN U6912 ( .A(n6443), .B(n6442), .Z(n6447) );
  NANDN U6913 ( .A(n6445), .B(n6444), .Z(n6446) );
  NAND U6914 ( .A(n6447), .B(n6446), .Z(n6653) );
  XOR U6915 ( .A(n6654), .B(n6653), .Z(n6656) );
  XNOR U6916 ( .A(n6655), .B(n6656), .Z(n6647) );
  XNOR U6917 ( .A(n6648), .B(n6647), .Z(n6649) );
  XOR U6918 ( .A(n6649), .B(n6650), .Z(n6789) );
  XNOR U6919 ( .A(n6788), .B(n6789), .Z(n6790) );
  XOR U6920 ( .A(n6791), .B(n6790), .Z(n6785) );
  NANDN U6921 ( .A(n6453), .B(n6452), .Z(n6457) );
  NAND U6922 ( .A(n6455), .B(n6454), .Z(n6456) );
  AND U6923 ( .A(n6457), .B(n6456), .Z(n6782) );
  NANDN U6924 ( .A(n6459), .B(n6458), .Z(n6463) );
  NAND U6925 ( .A(n6461), .B(n6460), .Z(n6462) );
  AND U6926 ( .A(n6463), .B(n6462), .Z(n6779) );
  NANDN U6927 ( .A(n6465), .B(n6464), .Z(n6469) );
  NAND U6928 ( .A(n6467), .B(n6466), .Z(n6468) );
  AND U6929 ( .A(n6469), .B(n6468), .Z(n6777) );
  NANDN U6930 ( .A(n6471), .B(n6470), .Z(n6475) );
  NANDN U6931 ( .A(n6473), .B(n6472), .Z(n6474) );
  AND U6932 ( .A(n6475), .B(n6474), .Z(n6771) );
  NANDN U6933 ( .A(n6476), .B(n36962), .Z(n6478) );
  XOR U6934 ( .A(b[43]), .B(a[10]), .Z(n6680) );
  NANDN U6935 ( .A(n36891), .B(n6680), .Z(n6477) );
  AND U6936 ( .A(n6478), .B(n6477), .Z(n6766) );
  NANDN U6937 ( .A(n29499), .B(n6479), .Z(n6481) );
  XOR U6938 ( .A(b[7]), .B(a[46]), .Z(n6620) );
  NANDN U6939 ( .A(n29735), .B(n6620), .Z(n6480) );
  AND U6940 ( .A(n6481), .B(n6480), .Z(n6765) );
  NANDN U6941 ( .A(n33875), .B(n6482), .Z(n6484) );
  XOR U6942 ( .A(b[25]), .B(a[28]), .Z(n6692) );
  NANDN U6943 ( .A(n33994), .B(n6692), .Z(n6483) );
  NAND U6944 ( .A(n6484), .B(n6483), .Z(n6764) );
  XOR U6945 ( .A(n6765), .B(n6764), .Z(n6767) );
  XNOR U6946 ( .A(n6766), .B(n6767), .Z(n6770) );
  XNOR U6947 ( .A(n6771), .B(n6770), .Z(n6773) );
  NANDN U6948 ( .A(n6486), .B(n6485), .Z(n6490) );
  NANDN U6949 ( .A(n6488), .B(n6487), .Z(n6489) );
  AND U6950 ( .A(n6490), .B(n6489), .Z(n6772) );
  XOR U6951 ( .A(n6773), .B(n6772), .Z(n6644) );
  NANDN U6952 ( .A(n6492), .B(n6491), .Z(n6496) );
  OR U6953 ( .A(n6494), .B(n6493), .Z(n6495) );
  AND U6954 ( .A(n6496), .B(n6495), .Z(n6662) );
  NANDN U6955 ( .A(n209), .B(n6497), .Z(n6499) );
  XOR U6956 ( .A(b[3]), .B(a[50]), .Z(n6677) );
  NANDN U6957 ( .A(n28941), .B(n6677), .Z(n6498) );
  AND U6958 ( .A(n6499), .B(n6498), .Z(n6708) );
  NANDN U6959 ( .A(n6500), .B(n35001), .Z(n6502) );
  XOR U6960 ( .A(b[29]), .B(a[24]), .Z(n6683) );
  NANDN U6961 ( .A(n34722), .B(n6683), .Z(n6501) );
  NAND U6962 ( .A(n6502), .B(n6501), .Z(n6707) );
  XNOR U6963 ( .A(n6708), .B(n6707), .Z(n6710) );
  NOR U6964 ( .A(n6504), .B(n6503), .Z(n6709) );
  XOR U6965 ( .A(n6710), .B(n6709), .Z(n6660) );
  NANDN U6966 ( .A(n6505), .B(n37202), .Z(n6507) );
  XOR U6967 ( .A(b[45]), .B(a[8]), .Z(n6749) );
  NANDN U6968 ( .A(n37083), .B(n6749), .Z(n6506) );
  AND U6969 ( .A(n6507), .B(n6506), .Z(n6703) );
  NANDN U6970 ( .A(n211), .B(n6508), .Z(n6510) );
  XOR U6971 ( .A(b[47]), .B(a[6]), .Z(n6686) );
  NANDN U6972 ( .A(n37172), .B(n6686), .Z(n6509) );
  AND U6973 ( .A(n6510), .B(n6509), .Z(n6702) );
  NANDN U6974 ( .A(n6511), .B(n34647), .Z(n6513) );
  XOR U6975 ( .A(b[27]), .B(a[26]), .Z(n6719) );
  NANDN U6976 ( .A(n34458), .B(n6719), .Z(n6512) );
  NAND U6977 ( .A(n6513), .B(n6512), .Z(n6701) );
  XOR U6978 ( .A(n6702), .B(n6701), .Z(n6704) );
  XNOR U6979 ( .A(n6703), .B(n6704), .Z(n6659) );
  XNOR U6980 ( .A(n6660), .B(n6659), .Z(n6661) );
  XOR U6981 ( .A(n6662), .B(n6661), .Z(n6642) );
  NANDN U6982 ( .A(n6515), .B(n6514), .Z(n6519) );
  OR U6983 ( .A(n6517), .B(n6516), .Z(n6518) );
  AND U6984 ( .A(n6519), .B(n6518), .Z(n6668) );
  NANDN U6985 ( .A(n35936), .B(n6520), .Z(n6522) );
  XOR U6986 ( .A(b[37]), .B(a[16]), .Z(n6591) );
  NANDN U6987 ( .A(n36047), .B(n6591), .Z(n6521) );
  AND U6988 ( .A(n6522), .B(n6521), .Z(n6601) );
  NANDN U6989 ( .A(n36480), .B(n6523), .Z(n6525) );
  XOR U6990 ( .A(b[41]), .B(a[12]), .Z(n6758) );
  NANDN U6991 ( .A(n36594), .B(n6758), .Z(n6524) );
  AND U6992 ( .A(n6525), .B(n6524), .Z(n6600) );
  NANDN U6993 ( .A(n31055), .B(n6526), .Z(n6528) );
  XOR U6994 ( .A(b[13]), .B(a[40]), .Z(n6734) );
  NANDN U6995 ( .A(n31293), .B(n6734), .Z(n6527) );
  NAND U6996 ( .A(n6528), .B(n6527), .Z(n6599) );
  XOR U6997 ( .A(n6600), .B(n6599), .Z(n6602) );
  XOR U6998 ( .A(n6601), .B(n6602), .Z(n6666) );
  NANDN U6999 ( .A(n30482), .B(n6529), .Z(n6531) );
  XOR U7000 ( .A(b[11]), .B(a[42]), .Z(n6731) );
  NANDN U7001 ( .A(n30891), .B(n6731), .Z(n6530) );
  AND U7002 ( .A(n6531), .B(n6530), .Z(n6625) );
  NANDN U7003 ( .A(n210), .B(n6532), .Z(n6534) );
  XOR U7004 ( .A(b[9]), .B(a[44]), .Z(n6611) );
  NANDN U7005 ( .A(n30267), .B(n6611), .Z(n6533) );
  AND U7006 ( .A(n6534), .B(n6533), .Z(n6624) );
  NANDN U7007 ( .A(n36210), .B(n6535), .Z(n6537) );
  XOR U7008 ( .A(b[39]), .B(a[14]), .Z(n6755) );
  NANDN U7009 ( .A(n36347), .B(n6755), .Z(n6536) );
  NAND U7010 ( .A(n6537), .B(n6536), .Z(n6623) );
  XOR U7011 ( .A(n6624), .B(n6623), .Z(n6626) );
  XNOR U7012 ( .A(n6625), .B(n6626), .Z(n6665) );
  XNOR U7013 ( .A(n6666), .B(n6665), .Z(n6667) );
  XNOR U7014 ( .A(n6668), .B(n6667), .Z(n6641) );
  XNOR U7015 ( .A(n6642), .B(n6641), .Z(n6643) );
  XNOR U7016 ( .A(n6644), .B(n6643), .Z(n6776) );
  XNOR U7017 ( .A(n6777), .B(n6776), .Z(n6778) );
  XOR U7018 ( .A(n6779), .B(n6778), .Z(n6783) );
  XNOR U7019 ( .A(n6782), .B(n6783), .Z(n6784) );
  XNOR U7020 ( .A(n6785), .B(n6784), .Z(n6800) );
  XNOR U7021 ( .A(n6801), .B(n6800), .Z(n6803) );
  NANDN U7022 ( .A(n6539), .B(n6538), .Z(n6543) );
  NANDN U7023 ( .A(n6541), .B(n6540), .Z(n6542) );
  AND U7024 ( .A(n6543), .B(n6542), .Z(n6797) );
  NANDN U7025 ( .A(n6545), .B(n6544), .Z(n6549) );
  OR U7026 ( .A(n6547), .B(n6546), .Z(n6548) );
  AND U7027 ( .A(n6549), .B(n6548), .Z(n6794) );
  NANDN U7028 ( .A(n6551), .B(n6550), .Z(n6555) );
  OR U7029 ( .A(n6553), .B(n6552), .Z(n6554) );
  NAND U7030 ( .A(n6555), .B(n6554), .Z(n6795) );
  XNOR U7031 ( .A(n6794), .B(n6795), .Z(n6796) );
  XNOR U7032 ( .A(n6797), .B(n6796), .Z(n6802) );
  XOR U7033 ( .A(n6803), .B(n6802), .Z(n6807) );
  NANDN U7034 ( .A(n6557), .B(n6556), .Z(n6561) );
  NANDN U7035 ( .A(n6559), .B(n6558), .Z(n6560) );
  AND U7036 ( .A(n6561), .B(n6560), .Z(n6806) );
  XNOR U7037 ( .A(n6807), .B(n6806), .Z(n6808) );
  NANDN U7038 ( .A(n6563), .B(n6562), .Z(n6567) );
  NAND U7039 ( .A(n6565), .B(n6564), .Z(n6566) );
  NAND U7040 ( .A(n6567), .B(n6566), .Z(n6809) );
  XNOR U7041 ( .A(n6808), .B(n6809), .Z(n6573) );
  XOR U7042 ( .A(n6574), .B(n6573), .Z(n6576) );
  XNOR U7043 ( .A(n6575), .B(n6576), .Z(n6569) );
  XOR U7044 ( .A(n6570), .B(n6569), .Z(c[116]) );
  NANDN U7045 ( .A(n6568), .B(sreg[116]), .Z(n6572) );
  NAND U7046 ( .A(n6570), .B(n6569), .Z(n6571) );
  AND U7047 ( .A(n6572), .B(n6571), .Z(n6814) );
  NANDN U7048 ( .A(n6574), .B(n6573), .Z(n6578) );
  OR U7049 ( .A(n6576), .B(n6575), .Z(n6577) );
  AND U7050 ( .A(n6578), .B(n6577), .Z(n6820) );
  NANDN U7051 ( .A(n6580), .B(n6579), .Z(n6584) );
  NANDN U7052 ( .A(n6582), .B(n6581), .Z(n6583) );
  NAND U7053 ( .A(n6584), .B(n6583), .Z(n7039) );
  NANDN U7054 ( .A(n35611), .B(n6585), .Z(n6587) );
  XOR U7055 ( .A(b[35]), .B(a[19]), .Z(n7022) );
  NANDN U7056 ( .A(n35801), .B(n7022), .Z(n6586) );
  AND U7057 ( .A(n6587), .B(n6586), .Z(n6986) );
  NANDN U7058 ( .A(n28889), .B(n6588), .Z(n6590) );
  XOR U7059 ( .A(b[5]), .B(a[49]), .Z(n6938) );
  NANDN U7060 ( .A(n29138), .B(n6938), .Z(n6589) );
  AND U7061 ( .A(n6590), .B(n6589), .Z(n6985) );
  NANDN U7062 ( .A(n35936), .B(n6591), .Z(n6593) );
  XOR U7063 ( .A(b[37]), .B(a[17]), .Z(n6887) );
  NANDN U7064 ( .A(n36047), .B(n6887), .Z(n6592) );
  NAND U7065 ( .A(n6593), .B(n6592), .Z(n6984) );
  XOR U7066 ( .A(n6985), .B(n6984), .Z(n6987) );
  XOR U7067 ( .A(n6986), .B(n6987), .Z(n6858) );
  NANDN U7068 ( .A(n6594), .B(n6723), .Z(n6598) );
  NANDN U7069 ( .A(n6596), .B(n6595), .Z(n6597) );
  AND U7070 ( .A(n6598), .B(n6597), .Z(n6857) );
  XNOR U7071 ( .A(n6858), .B(n6857), .Z(n6860) );
  NANDN U7072 ( .A(n6600), .B(n6599), .Z(n6604) );
  OR U7073 ( .A(n6602), .B(n6601), .Z(n6603) );
  AND U7074 ( .A(n6604), .B(n6603), .Z(n6859) );
  XOR U7075 ( .A(n6860), .B(n6859), .Z(n6911) );
  NANDN U7076 ( .A(n32013), .B(n6605), .Z(n6607) );
  XOR U7077 ( .A(b[17]), .B(a[37]), .Z(n6972) );
  NANDN U7078 ( .A(n32292), .B(n6972), .Z(n6606) );
  AND U7079 ( .A(n6607), .B(n6606), .Z(n6962) );
  NANDN U7080 ( .A(n6608), .B(n33000), .Z(n6610) );
  XOR U7081 ( .A(b[19]), .B(a[35]), .Z(n6893) );
  NANDN U7082 ( .A(n32823), .B(n6893), .Z(n6609) );
  AND U7083 ( .A(n6610), .B(n6609), .Z(n6961) );
  NANDN U7084 ( .A(n210), .B(n6611), .Z(n6613) );
  XOR U7085 ( .A(b[9]), .B(a[45]), .Z(n7019) );
  NANDN U7086 ( .A(n30267), .B(n7019), .Z(n6612) );
  NAND U7087 ( .A(n6613), .B(n6612), .Z(n6960) );
  XOR U7088 ( .A(n6961), .B(n6960), .Z(n6963) );
  XOR U7089 ( .A(n6962), .B(n6963), .Z(n6897) );
  NANDN U7090 ( .A(n32996), .B(n6614), .Z(n6616) );
  XOR U7091 ( .A(b[21]), .B(a[33]), .Z(n6932) );
  NANDN U7092 ( .A(n33271), .B(n6932), .Z(n6615) );
  AND U7093 ( .A(n6616), .B(n6615), .Z(n6877) );
  NANDN U7094 ( .A(n35260), .B(n6617), .Z(n6619) );
  XOR U7095 ( .A(b[33]), .B(a[21]), .Z(n6929) );
  NANDN U7096 ( .A(n35456), .B(n6929), .Z(n6618) );
  AND U7097 ( .A(n6619), .B(n6618), .Z(n6876) );
  NANDN U7098 ( .A(n29499), .B(n6620), .Z(n6622) );
  XOR U7099 ( .A(b[7]), .B(a[47]), .Z(n6935) );
  NANDN U7100 ( .A(n29735), .B(n6935), .Z(n6621) );
  NAND U7101 ( .A(n6622), .B(n6621), .Z(n6875) );
  XOR U7102 ( .A(n6876), .B(n6875), .Z(n6878) );
  XNOR U7103 ( .A(n6877), .B(n6878), .Z(n6896) );
  XNOR U7104 ( .A(n6897), .B(n6896), .Z(n6899) );
  NANDN U7105 ( .A(n6624), .B(n6623), .Z(n6628) );
  OR U7106 ( .A(n6626), .B(n6625), .Z(n6627) );
  AND U7107 ( .A(n6628), .B(n6627), .Z(n6898) );
  XOR U7108 ( .A(n6899), .B(n6898), .Z(n6909) );
  NANDN U7109 ( .A(n6630), .B(n6629), .Z(n6634) );
  OR U7110 ( .A(n6632), .B(n6631), .Z(n6633) );
  AND U7111 ( .A(n6634), .B(n6633), .Z(n6908) );
  XNOR U7112 ( .A(n6909), .B(n6908), .Z(n6910) );
  XOR U7113 ( .A(n6911), .B(n6910), .Z(n7038) );
  NANDN U7114 ( .A(n6636), .B(n6635), .Z(n6640) );
  NANDN U7115 ( .A(n6638), .B(n6637), .Z(n6639) );
  NAND U7116 ( .A(n6640), .B(n6639), .Z(n7037) );
  XOR U7117 ( .A(n7038), .B(n7037), .Z(n7040) );
  XNOR U7118 ( .A(n7039), .B(n7040), .Z(n7045) );
  NANDN U7119 ( .A(n6642), .B(n6641), .Z(n6646) );
  NANDN U7120 ( .A(n6644), .B(n6643), .Z(n6645) );
  AND U7121 ( .A(n6646), .B(n6645), .Z(n7044) );
  NANDN U7122 ( .A(n6648), .B(n6647), .Z(n6652) );
  NANDN U7123 ( .A(n6650), .B(n6649), .Z(n6651) );
  AND U7124 ( .A(n6652), .B(n6651), .Z(n7043) );
  XOR U7125 ( .A(n7044), .B(n7043), .Z(n7046) );
  XOR U7126 ( .A(n7045), .B(n7046), .Z(n7033) );
  NANDN U7127 ( .A(n6654), .B(n6653), .Z(n6658) );
  OR U7128 ( .A(n6656), .B(n6655), .Z(n6657) );
  AND U7129 ( .A(n6658), .B(n6657), .Z(n6835) );
  NANDN U7130 ( .A(n6660), .B(n6659), .Z(n6664) );
  NAND U7131 ( .A(n6662), .B(n6661), .Z(n6663) );
  AND U7132 ( .A(n6664), .B(n6663), .Z(n6834) );
  NANDN U7133 ( .A(n6666), .B(n6665), .Z(n6670) );
  NAND U7134 ( .A(n6668), .B(n6667), .Z(n6669) );
  NAND U7135 ( .A(n6670), .B(n6669), .Z(n6833) );
  XOR U7136 ( .A(n6834), .B(n6833), .Z(n6836) );
  XNOR U7137 ( .A(n6835), .B(n6836), .Z(n7027) );
  NANDN U7138 ( .A(n6672), .B(n6671), .Z(n6676) );
  OR U7139 ( .A(n6674), .B(n6673), .Z(n6675) );
  AND U7140 ( .A(n6676), .B(n6675), .Z(n6828) );
  NANDN U7141 ( .A(n209), .B(n6677), .Z(n6679) );
  XOR U7142 ( .A(b[3]), .B(a[51]), .Z(n7010) );
  NANDN U7143 ( .A(n28941), .B(n7010), .Z(n6678) );
  AND U7144 ( .A(n6679), .B(n6678), .Z(n6871) );
  NANDN U7145 ( .A(n36742), .B(n6680), .Z(n6682) );
  XOR U7146 ( .A(b[43]), .B(a[11]), .Z(n6890) );
  NANDN U7147 ( .A(n36891), .B(n6890), .Z(n6681) );
  AND U7148 ( .A(n6682), .B(n6681), .Z(n6870) );
  NANDN U7149 ( .A(n34634), .B(n6683), .Z(n6685) );
  XOR U7150 ( .A(b[29]), .B(a[25]), .Z(n7013) );
  NANDN U7151 ( .A(n34722), .B(n7013), .Z(n6684) );
  NAND U7152 ( .A(n6685), .B(n6684), .Z(n6869) );
  XOR U7153 ( .A(n6870), .B(n6869), .Z(n6872) );
  XOR U7154 ( .A(n6871), .B(n6872), .Z(n6840) );
  NANDN U7155 ( .A(n211), .B(n6686), .Z(n6688) );
  XOR U7156 ( .A(b[47]), .B(a[7]), .Z(n6969) );
  NANDN U7157 ( .A(n37172), .B(n6969), .Z(n6687) );
  AND U7158 ( .A(n6688), .B(n6687), .Z(n6992) );
  NANDN U7159 ( .A(n212), .B(n6689), .Z(n6691) );
  XOR U7160 ( .A(b[49]), .B(a[5]), .Z(n6978) );
  NANDN U7161 ( .A(n37432), .B(n6978), .Z(n6690) );
  AND U7162 ( .A(n6691), .B(n6690), .Z(n6991) );
  NANDN U7163 ( .A(n33875), .B(n6692), .Z(n6694) );
  XOR U7164 ( .A(b[25]), .B(a[29]), .Z(n6923) );
  NANDN U7165 ( .A(n33994), .B(n6923), .Z(n6693) );
  NAND U7166 ( .A(n6694), .B(n6693), .Z(n6990) );
  XOR U7167 ( .A(n6991), .B(n6990), .Z(n6993) );
  XNOR U7168 ( .A(n6992), .B(n6993), .Z(n6839) );
  XNOR U7169 ( .A(n6840), .B(n6839), .Z(n6842) );
  NANDN U7170 ( .A(n6696), .B(n6695), .Z(n6700) );
  OR U7171 ( .A(n6698), .B(n6697), .Z(n6699) );
  AND U7172 ( .A(n6700), .B(n6699), .Z(n6841) );
  XOR U7173 ( .A(n6842), .B(n6841), .Z(n6854) );
  NANDN U7174 ( .A(n6702), .B(n6701), .Z(n6706) );
  OR U7175 ( .A(n6704), .B(n6703), .Z(n6705) );
  AND U7176 ( .A(n6706), .B(n6705), .Z(n6852) );
  NANDN U7177 ( .A(n6708), .B(n6707), .Z(n6712) );
  NAND U7178 ( .A(n6710), .B(n6709), .Z(n6711) );
  NAND U7179 ( .A(n6712), .B(n6711), .Z(n6851) );
  XNOR U7180 ( .A(n6852), .B(n6851), .Z(n6853) );
  XNOR U7181 ( .A(n6854), .B(n6853), .Z(n6827) );
  XNOR U7182 ( .A(n6828), .B(n6827), .Z(n6830) );
  NANDN U7183 ( .A(n6714), .B(n6713), .Z(n6718) );
  OR U7184 ( .A(n6716), .B(n6715), .Z(n6717) );
  AND U7185 ( .A(n6718), .B(n6717), .Z(n6848) );
  NANDN U7186 ( .A(n34223), .B(n6719), .Z(n6721) );
  XOR U7187 ( .A(b[27]), .B(a[27]), .Z(n6920) );
  NANDN U7188 ( .A(n34458), .B(n6920), .Z(n6720) );
  AND U7189 ( .A(n6721), .B(n6720), .Z(n6955) );
  NAND U7190 ( .A(b[51]), .B(b[52]), .Z(n6722) );
  NAND U7191 ( .A(b[53]), .B(n6722), .Z(n37964) );
  NOR U7192 ( .A(n37964), .B(n6723), .Z(n6954) );
  XNOR U7193 ( .A(n6955), .B(n6954), .Z(n6956) );
  NANDN U7194 ( .A(n37526), .B(n6724), .Z(n6726) );
  XOR U7195 ( .A(b[51]), .B(a[3]), .Z(n6881) );
  NANDN U7196 ( .A(n37605), .B(n6881), .Z(n6725) );
  AND U7197 ( .A(n6726), .B(n6725), .Z(n7008) );
  XOR U7198 ( .A(b[53]), .B(b[52]), .Z(n6947) );
  XOR U7199 ( .A(b[53]), .B(a[0]), .Z(n6727) );
  NAND U7200 ( .A(n6947), .B(n6727), .Z(n6728) );
  OR U7201 ( .A(n6728), .B(n37850), .Z(n6730) );
  XOR U7202 ( .A(b[53]), .B(a[1]), .Z(n6948) );
  NAND U7203 ( .A(n37850), .B(n6948), .Z(n6729) );
  NAND U7204 ( .A(n6730), .B(n6729), .Z(n7009) );
  XOR U7205 ( .A(n7008), .B(n7009), .Z(n6957) );
  XNOR U7206 ( .A(n6956), .B(n6957), .Z(n6845) );
  NANDN U7207 ( .A(n30482), .B(n6731), .Z(n6733) );
  XOR U7208 ( .A(b[11]), .B(a[43]), .Z(n7016) );
  NANDN U7209 ( .A(n30891), .B(n7016), .Z(n6732) );
  AND U7210 ( .A(n6733), .B(n6732), .Z(n7005) );
  NANDN U7211 ( .A(n31055), .B(n6734), .Z(n6736) );
  XOR U7212 ( .A(b[13]), .B(a[41]), .Z(n6944) );
  NANDN U7213 ( .A(n31293), .B(n6944), .Z(n6735) );
  AND U7214 ( .A(n6736), .B(n6735), .Z(n7003) );
  NANDN U7215 ( .A(n31536), .B(n6737), .Z(n6739) );
  XOR U7216 ( .A(b[15]), .B(a[39]), .Z(n6975) );
  NANDN U7217 ( .A(n31925), .B(n6975), .Z(n6738) );
  NAND U7218 ( .A(n6739), .B(n6738), .Z(n7002) );
  XNOR U7219 ( .A(n7003), .B(n7002), .Z(n7004) );
  XOR U7220 ( .A(n7005), .B(n7004), .Z(n6846) );
  XNOR U7221 ( .A(n6845), .B(n6846), .Z(n6847) );
  XNOR U7222 ( .A(n6848), .B(n6847), .Z(n6916) );
  NANDN U7223 ( .A(n6741), .B(n6740), .Z(n6745) );
  NANDN U7224 ( .A(n6743), .B(n6742), .Z(n6744) );
  AND U7225 ( .A(n6745), .B(n6744), .Z(n6915) );
  NAND U7226 ( .A(b[0]), .B(a[53]), .Z(n6746) );
  XNOR U7227 ( .A(b[1]), .B(n6746), .Z(n6748) );
  NANDN U7228 ( .A(b[0]), .B(a[52]), .Z(n6747) );
  NAND U7229 ( .A(n6748), .B(n6747), .Z(n6866) );
  NANDN U7230 ( .A(n36991), .B(n6749), .Z(n6751) );
  XOR U7231 ( .A(b[45]), .B(a[9]), .Z(n6966) );
  NANDN U7232 ( .A(n37083), .B(n6966), .Z(n6750) );
  AND U7233 ( .A(n6751), .B(n6750), .Z(n6864) );
  NANDN U7234 ( .A(n33866), .B(n6752), .Z(n6754) );
  XOR U7235 ( .A(b[23]), .B(a[31]), .Z(n6926) );
  NANDN U7236 ( .A(n33644), .B(n6926), .Z(n6753) );
  NAND U7237 ( .A(n6754), .B(n6753), .Z(n6863) );
  XOR U7238 ( .A(n6864), .B(n6863), .Z(n6865) );
  XOR U7239 ( .A(n6866), .B(n6865), .Z(n6903) );
  NANDN U7240 ( .A(n36210), .B(n6755), .Z(n6757) );
  XOR U7241 ( .A(b[39]), .B(a[15]), .Z(n6951) );
  NANDN U7242 ( .A(n36347), .B(n6951), .Z(n6756) );
  AND U7243 ( .A(n6757), .B(n6756), .Z(n6998) );
  NANDN U7244 ( .A(n36480), .B(n6758), .Z(n6760) );
  XOR U7245 ( .A(b[41]), .B(a[13]), .Z(n6981) );
  NANDN U7246 ( .A(n36594), .B(n6981), .Z(n6759) );
  AND U7247 ( .A(n6760), .B(n6759), .Z(n6997) );
  NANDN U7248 ( .A(n34909), .B(n6761), .Z(n6763) );
  XOR U7249 ( .A(b[31]), .B(a[23]), .Z(n6941) );
  NANDN U7250 ( .A(n35145), .B(n6941), .Z(n6762) );
  NAND U7251 ( .A(n6763), .B(n6762), .Z(n6996) );
  XOR U7252 ( .A(n6997), .B(n6996), .Z(n6999) );
  XNOR U7253 ( .A(n6998), .B(n6999), .Z(n6902) );
  XNOR U7254 ( .A(n6903), .B(n6902), .Z(n6905) );
  NANDN U7255 ( .A(n6765), .B(n6764), .Z(n6769) );
  OR U7256 ( .A(n6767), .B(n6766), .Z(n6768) );
  AND U7257 ( .A(n6769), .B(n6768), .Z(n6904) );
  XNOR U7258 ( .A(n6905), .B(n6904), .Z(n6914) );
  XOR U7259 ( .A(n6915), .B(n6914), .Z(n6917) );
  XNOR U7260 ( .A(n6916), .B(n6917), .Z(n6829) );
  XOR U7261 ( .A(n6830), .B(n6829), .Z(n7026) );
  NANDN U7262 ( .A(n6771), .B(n6770), .Z(n6775) );
  NAND U7263 ( .A(n6773), .B(n6772), .Z(n6774) );
  NAND U7264 ( .A(n6775), .B(n6774), .Z(n7025) );
  XOR U7265 ( .A(n7026), .B(n7025), .Z(n7028) );
  XNOR U7266 ( .A(n7027), .B(n7028), .Z(n7031) );
  NANDN U7267 ( .A(n6777), .B(n6776), .Z(n6781) );
  NANDN U7268 ( .A(n6779), .B(n6778), .Z(n6780) );
  NAND U7269 ( .A(n6781), .B(n6780), .Z(n7032) );
  XOR U7270 ( .A(n7031), .B(n7032), .Z(n7034) );
  XOR U7271 ( .A(n7033), .B(n7034), .Z(n6825) );
  NANDN U7272 ( .A(n6783), .B(n6782), .Z(n6787) );
  NANDN U7273 ( .A(n6785), .B(n6784), .Z(n6786) );
  AND U7274 ( .A(n6787), .B(n6786), .Z(n6824) );
  NANDN U7275 ( .A(n6789), .B(n6788), .Z(n6793) );
  NAND U7276 ( .A(n6791), .B(n6790), .Z(n6792) );
  AND U7277 ( .A(n6793), .B(n6792), .Z(n6823) );
  XNOR U7278 ( .A(n6824), .B(n6823), .Z(n6826) );
  XOR U7279 ( .A(n6825), .B(n6826), .Z(n7052) );
  NANDN U7280 ( .A(n6795), .B(n6794), .Z(n6799) );
  NANDN U7281 ( .A(n6797), .B(n6796), .Z(n6798) );
  AND U7282 ( .A(n6799), .B(n6798), .Z(n7050) );
  NANDN U7283 ( .A(n6801), .B(n6800), .Z(n6805) );
  NAND U7284 ( .A(n6803), .B(n6802), .Z(n6804) );
  NAND U7285 ( .A(n6805), .B(n6804), .Z(n7049) );
  XNOR U7286 ( .A(n7050), .B(n7049), .Z(n7051) );
  XOR U7287 ( .A(n7052), .B(n7051), .Z(n6818) );
  NANDN U7288 ( .A(n6807), .B(n6806), .Z(n6811) );
  NANDN U7289 ( .A(n6809), .B(n6808), .Z(n6810) );
  NAND U7290 ( .A(n6811), .B(n6810), .Z(n6817) );
  XNOR U7291 ( .A(n6818), .B(n6817), .Z(n6819) );
  XNOR U7292 ( .A(n6820), .B(n6819), .Z(n6812) );
  XNOR U7293 ( .A(sreg[117]), .B(n6812), .Z(n6813) );
  XNOR U7294 ( .A(n6814), .B(n6813), .Z(c[117]) );
  NANDN U7295 ( .A(sreg[117]), .B(n6812), .Z(n6816) );
  NAND U7296 ( .A(n6814), .B(n6813), .Z(n6815) );
  NAND U7297 ( .A(n6816), .B(n6815), .Z(n7055) );
  XNOR U7298 ( .A(sreg[118]), .B(n7055), .Z(n7057) );
  NANDN U7299 ( .A(n6818), .B(n6817), .Z(n6822) );
  NANDN U7300 ( .A(n6820), .B(n6819), .Z(n6821) );
  AND U7301 ( .A(n6822), .B(n6821), .Z(n7063) );
  NANDN U7302 ( .A(n6828), .B(n6827), .Z(n6832) );
  NAND U7303 ( .A(n6830), .B(n6829), .Z(n6831) );
  AND U7304 ( .A(n6832), .B(n6831), .Z(n7158) );
  NANDN U7305 ( .A(n6834), .B(n6833), .Z(n6838) );
  NANDN U7306 ( .A(n6836), .B(n6835), .Z(n6837) );
  AND U7307 ( .A(n6838), .B(n6837), .Z(n7157) );
  XNOR U7308 ( .A(n7158), .B(n7157), .Z(n7160) );
  NANDN U7309 ( .A(n6840), .B(n6839), .Z(n6844) );
  NAND U7310 ( .A(n6842), .B(n6841), .Z(n6843) );
  AND U7311 ( .A(n6844), .B(n6843), .Z(n7293) );
  NANDN U7312 ( .A(n6846), .B(n6845), .Z(n6850) );
  NANDN U7313 ( .A(n6848), .B(n6847), .Z(n6849) );
  AND U7314 ( .A(n6850), .B(n6849), .Z(n7292) );
  XNOR U7315 ( .A(n7293), .B(n7292), .Z(n7295) );
  NANDN U7316 ( .A(n6852), .B(n6851), .Z(n6856) );
  NANDN U7317 ( .A(n6854), .B(n6853), .Z(n6855) );
  AND U7318 ( .A(n6856), .B(n6855), .Z(n7294) );
  XOR U7319 ( .A(n7295), .B(n7294), .Z(n7154) );
  NANDN U7320 ( .A(n6858), .B(n6857), .Z(n6862) );
  NAND U7321 ( .A(n6860), .B(n6859), .Z(n6861) );
  AND U7322 ( .A(n6862), .B(n6861), .Z(n7300) );
  NANDN U7323 ( .A(n6864), .B(n6863), .Z(n6868) );
  OR U7324 ( .A(n6866), .B(n6865), .Z(n6867) );
  AND U7325 ( .A(n6868), .B(n6867), .Z(n7170) );
  NANDN U7326 ( .A(n6870), .B(n6869), .Z(n6874) );
  OR U7327 ( .A(n6872), .B(n6871), .Z(n6873) );
  NAND U7328 ( .A(n6874), .B(n6873), .Z(n7169) );
  XNOR U7329 ( .A(n7170), .B(n7169), .Z(n7172) );
  NANDN U7330 ( .A(n6876), .B(n6875), .Z(n6880) );
  OR U7331 ( .A(n6878), .B(n6877), .Z(n6879) );
  AND U7332 ( .A(n6880), .B(n6879), .Z(n7136) );
  XOR U7333 ( .A(b[54]), .B(b[53]), .Z(n37985) );
  IV U7334 ( .A(n37985), .Z(n37911) );
  ANDN U7335 ( .B(a[0]), .A(n37911), .Z(n7103) );
  NANDN U7336 ( .A(n37526), .B(n6881), .Z(n6883) );
  XOR U7337 ( .A(b[51]), .B(a[4]), .Z(n7256) );
  NANDN U7338 ( .A(n37605), .B(n7256), .Z(n6882) );
  AND U7339 ( .A(n6883), .B(n6882), .Z(n7104) );
  XNOR U7340 ( .A(n7103), .B(n7104), .Z(n7105) );
  NAND U7341 ( .A(b[0]), .B(a[54]), .Z(n6884) );
  XNOR U7342 ( .A(b[1]), .B(n6884), .Z(n6886) );
  NANDN U7343 ( .A(b[0]), .B(a[53]), .Z(n6885) );
  NAND U7344 ( .A(n6886), .B(n6885), .Z(n7106) );
  XNOR U7345 ( .A(n7105), .B(n7106), .Z(n7133) );
  NANDN U7346 ( .A(n35936), .B(n6887), .Z(n6889) );
  XOR U7347 ( .A(b[37]), .B(a[18]), .Z(n7226) );
  NANDN U7348 ( .A(n36047), .B(n7226), .Z(n6888) );
  AND U7349 ( .A(n6889), .B(n6888), .Z(n7130) );
  NANDN U7350 ( .A(n36742), .B(n6890), .Z(n6892) );
  XOR U7351 ( .A(b[43]), .B(a[12]), .Z(n7220) );
  NANDN U7352 ( .A(n36891), .B(n7220), .Z(n6891) );
  AND U7353 ( .A(n6892), .B(n6891), .Z(n7128) );
  NANDN U7354 ( .A(n32483), .B(n6893), .Z(n6895) );
  XOR U7355 ( .A(b[19]), .B(a[36]), .Z(n7271) );
  NANDN U7356 ( .A(n32823), .B(n7271), .Z(n6894) );
  NAND U7357 ( .A(n6895), .B(n6894), .Z(n7127) );
  XNOR U7358 ( .A(n7128), .B(n7127), .Z(n7129) );
  XOR U7359 ( .A(n7130), .B(n7129), .Z(n7134) );
  XNOR U7360 ( .A(n7133), .B(n7134), .Z(n7135) );
  XNOR U7361 ( .A(n7136), .B(n7135), .Z(n7171) );
  XOR U7362 ( .A(n7172), .B(n7171), .Z(n7299) );
  NANDN U7363 ( .A(n6897), .B(n6896), .Z(n6901) );
  NAND U7364 ( .A(n6899), .B(n6898), .Z(n6900) );
  NAND U7365 ( .A(n6901), .B(n6900), .Z(n7298) );
  XOR U7366 ( .A(n7299), .B(n7298), .Z(n7301) );
  XOR U7367 ( .A(n7300), .B(n7301), .Z(n7152) );
  NANDN U7368 ( .A(n6903), .B(n6902), .Z(n6907) );
  NAND U7369 ( .A(n6905), .B(n6904), .Z(n6906) );
  AND U7370 ( .A(n6907), .B(n6906), .Z(n7151) );
  XNOR U7371 ( .A(n7152), .B(n7151), .Z(n7153) );
  XNOR U7372 ( .A(n7154), .B(n7153), .Z(n7159) );
  XOR U7373 ( .A(n7160), .B(n7159), .Z(n7306) );
  NANDN U7374 ( .A(n6909), .B(n6908), .Z(n6913) );
  NANDN U7375 ( .A(n6911), .B(n6910), .Z(n6912) );
  AND U7376 ( .A(n6913), .B(n6912), .Z(n7080) );
  NANDN U7377 ( .A(n6915), .B(n6914), .Z(n6919) );
  NANDN U7378 ( .A(n6917), .B(n6916), .Z(n6918) );
  AND U7379 ( .A(n6919), .B(n6918), .Z(n7079) );
  NANDN U7380 ( .A(n34223), .B(n6920), .Z(n6922) );
  XOR U7381 ( .A(b[27]), .B(a[28]), .Z(n7115) );
  NANDN U7382 ( .A(n34458), .B(n7115), .Z(n6921) );
  AND U7383 ( .A(n6922), .B(n6921), .Z(n7189) );
  NANDN U7384 ( .A(n33875), .B(n6923), .Z(n6925) );
  XOR U7385 ( .A(b[25]), .B(a[30]), .Z(n7235) );
  NANDN U7386 ( .A(n33994), .B(n7235), .Z(n6924) );
  AND U7387 ( .A(n6925), .B(n6924), .Z(n7188) );
  NANDN U7388 ( .A(n33866), .B(n6926), .Z(n6928) );
  XOR U7389 ( .A(b[23]), .B(a[32]), .Z(n7229) );
  NANDN U7390 ( .A(n33644), .B(n7229), .Z(n6927) );
  AND U7391 ( .A(n6928), .B(n6927), .Z(n7087) );
  NANDN U7392 ( .A(n35260), .B(n6929), .Z(n6931) );
  XOR U7393 ( .A(b[33]), .B(a[22]), .Z(n7262) );
  NANDN U7394 ( .A(n35456), .B(n7262), .Z(n6930) );
  AND U7395 ( .A(n6931), .B(n6930), .Z(n7085) );
  NANDN U7396 ( .A(n32996), .B(n6932), .Z(n6934) );
  XOR U7397 ( .A(b[21]), .B(a[34]), .Z(n7223) );
  NANDN U7398 ( .A(n33271), .B(n7223), .Z(n6933) );
  NAND U7399 ( .A(n6934), .B(n6933), .Z(n7084) );
  XNOR U7400 ( .A(n7085), .B(n7084), .Z(n7086) );
  XNOR U7401 ( .A(n7087), .B(n7086), .Z(n7187) );
  XOR U7402 ( .A(n7188), .B(n7187), .Z(n7190) );
  XOR U7403 ( .A(n7189), .B(n7190), .Z(n7178) );
  NANDN U7404 ( .A(n29499), .B(n6935), .Z(n6937) );
  XOR U7405 ( .A(b[7]), .B(a[48]), .Z(n7196) );
  NANDN U7406 ( .A(n29735), .B(n7196), .Z(n6936) );
  AND U7407 ( .A(n6937), .B(n6936), .Z(n7246) );
  NANDN U7408 ( .A(n28889), .B(n6938), .Z(n6940) );
  XOR U7409 ( .A(b[5]), .B(a[50]), .Z(n7259) );
  NANDN U7410 ( .A(n29138), .B(n7259), .Z(n6939) );
  AND U7411 ( .A(n6940), .B(n6939), .Z(n7245) );
  NANDN U7412 ( .A(n34909), .B(n6941), .Z(n6943) );
  XOR U7413 ( .A(b[31]), .B(a[24]), .Z(n7232) );
  NANDN U7414 ( .A(n35145), .B(n7232), .Z(n6942) );
  NAND U7415 ( .A(n6943), .B(n6942), .Z(n7244) );
  XOR U7416 ( .A(n7245), .B(n7244), .Z(n7247) );
  XOR U7417 ( .A(n7246), .B(n7247), .Z(n7176) );
  NANDN U7418 ( .A(n31055), .B(n6944), .Z(n6946) );
  XOR U7419 ( .A(b[13]), .B(a[42]), .Z(n7118) );
  NANDN U7420 ( .A(n31293), .B(n7118), .Z(n6945) );
  AND U7421 ( .A(n6946), .B(n6945), .Z(n7282) );
  ANDN U7422 ( .B(n6947), .A(n37850), .Z(n37849) );
  IV U7423 ( .A(n37849), .Z(n37705) );
  NANDN U7424 ( .A(n37705), .B(n6948), .Z(n6950) );
  XOR U7425 ( .A(b[53]), .B(a[2]), .Z(n7090) );
  NANDN U7426 ( .A(n37778), .B(n7090), .Z(n6949) );
  AND U7427 ( .A(n6950), .B(n6949), .Z(n7281) );
  NANDN U7428 ( .A(n36210), .B(n6951), .Z(n6953) );
  XOR U7429 ( .A(b[39]), .B(a[16]), .Z(n7124) );
  NANDN U7430 ( .A(n36347), .B(n7124), .Z(n6952) );
  NAND U7431 ( .A(n6953), .B(n6952), .Z(n7280) );
  XOR U7432 ( .A(n7281), .B(n7280), .Z(n7283) );
  XNOR U7433 ( .A(n7282), .B(n7283), .Z(n7175) );
  XNOR U7434 ( .A(n7176), .B(n7175), .Z(n7177) );
  XNOR U7435 ( .A(n7178), .B(n7177), .Z(n7148) );
  NANDN U7436 ( .A(n6955), .B(n6954), .Z(n6959) );
  NANDN U7437 ( .A(n6957), .B(n6956), .Z(n6958) );
  AND U7438 ( .A(n6959), .B(n6958), .Z(n7145) );
  NANDN U7439 ( .A(n6961), .B(n6960), .Z(n6965) );
  OR U7440 ( .A(n6963), .B(n6962), .Z(n6964) );
  NAND U7441 ( .A(n6965), .B(n6964), .Z(n7146) );
  XNOR U7442 ( .A(n7145), .B(n7146), .Z(n7147) );
  XOR U7443 ( .A(n7148), .B(n7147), .Z(n7166) );
  NANDN U7444 ( .A(n36991), .B(n6966), .Z(n6968) );
  XOR U7445 ( .A(b[45]), .B(a[10]), .Z(n7265) );
  NANDN U7446 ( .A(n37083), .B(n7265), .Z(n6967) );
  AND U7447 ( .A(n6968), .B(n6967), .Z(n7276) );
  NANDN U7448 ( .A(n211), .B(n6969), .Z(n6971) );
  XOR U7449 ( .A(b[47]), .B(a[8]), .Z(n7268) );
  NANDN U7450 ( .A(n37172), .B(n7268), .Z(n6970) );
  AND U7451 ( .A(n6971), .B(n6970), .Z(n7275) );
  NANDN U7452 ( .A(n32013), .B(n6972), .Z(n6974) );
  XOR U7453 ( .A(b[17]), .B(a[38]), .Z(n7202) );
  NANDN U7454 ( .A(n32292), .B(n7202), .Z(n6973) );
  NAND U7455 ( .A(n6974), .B(n6973), .Z(n7274) );
  XOR U7456 ( .A(n7275), .B(n7274), .Z(n7277) );
  XOR U7457 ( .A(n7276), .B(n7277), .Z(n7182) );
  NANDN U7458 ( .A(n31536), .B(n6975), .Z(n6977) );
  XOR U7459 ( .A(b[15]), .B(a[40]), .Z(n7205) );
  NANDN U7460 ( .A(n31925), .B(n7205), .Z(n6976) );
  AND U7461 ( .A(n6977), .B(n6976), .Z(n7213) );
  NANDN U7462 ( .A(n212), .B(n6978), .Z(n6980) );
  XOR U7463 ( .A(b[49]), .B(a[6]), .Z(n7208) );
  NANDN U7464 ( .A(n37432), .B(n7208), .Z(n6979) );
  AND U7465 ( .A(n6980), .B(n6979), .Z(n7212) );
  NANDN U7466 ( .A(n36480), .B(n6981), .Z(n6983) );
  XOR U7467 ( .A(b[41]), .B(a[14]), .Z(n7217) );
  NANDN U7468 ( .A(n36594), .B(n7217), .Z(n6982) );
  NAND U7469 ( .A(n6983), .B(n6982), .Z(n7211) );
  XOR U7470 ( .A(n7212), .B(n7211), .Z(n7214) );
  XNOR U7471 ( .A(n7213), .B(n7214), .Z(n7181) );
  XNOR U7472 ( .A(n7182), .B(n7181), .Z(n7184) );
  NANDN U7473 ( .A(n6985), .B(n6984), .Z(n6989) );
  OR U7474 ( .A(n6987), .B(n6986), .Z(n6988) );
  AND U7475 ( .A(n6989), .B(n6988), .Z(n7183) );
  XOR U7476 ( .A(n7184), .B(n7183), .Z(n7164) );
  NANDN U7477 ( .A(n6991), .B(n6990), .Z(n6995) );
  OR U7478 ( .A(n6993), .B(n6992), .Z(n6994) );
  AND U7479 ( .A(n6995), .B(n6994), .Z(n7140) );
  NANDN U7480 ( .A(n6997), .B(n6996), .Z(n7001) );
  OR U7481 ( .A(n6999), .B(n6998), .Z(n7000) );
  NAND U7482 ( .A(n7001), .B(n7000), .Z(n7139) );
  XNOR U7483 ( .A(n7140), .B(n7139), .Z(n7141) );
  NANDN U7484 ( .A(n7003), .B(n7002), .Z(n7007) );
  NANDN U7485 ( .A(n7005), .B(n7004), .Z(n7006) );
  AND U7486 ( .A(n7007), .B(n7006), .Z(n7253) );
  ANDN U7487 ( .B(n7009), .A(n7008), .Z(n7288) );
  NAND U7488 ( .A(n9942), .B(n7010), .Z(n7012) );
  XNOR U7489 ( .A(b[3]), .B(a[52]), .Z(n7109) );
  NANDN U7490 ( .A(n7109), .B(n9653), .Z(n7011) );
  AND U7491 ( .A(n7012), .B(n7011), .Z(n7286) );
  NAND U7492 ( .A(n35001), .B(n7013), .Z(n7015) );
  XNOR U7493 ( .A(b[29]), .B(a[26]), .Z(n7100) );
  NANDN U7494 ( .A(n7100), .B(n35002), .Z(n7014) );
  NAND U7495 ( .A(n7015), .B(n7014), .Z(n7287) );
  XOR U7496 ( .A(n7286), .B(n7287), .Z(n7289) );
  XOR U7497 ( .A(n7288), .B(n7289), .Z(n7251) );
  NANDN U7498 ( .A(n30482), .B(n7016), .Z(n7018) );
  XOR U7499 ( .A(b[11]), .B(a[44]), .Z(n7121) );
  NANDN U7500 ( .A(n30891), .B(n7121), .Z(n7017) );
  AND U7501 ( .A(n7018), .B(n7017), .Z(n7241) );
  NANDN U7502 ( .A(n210), .B(n7019), .Z(n7021) );
  XOR U7503 ( .A(b[9]), .B(a[46]), .Z(n7193) );
  NANDN U7504 ( .A(n30267), .B(n7193), .Z(n7020) );
  AND U7505 ( .A(n7021), .B(n7020), .Z(n7239) );
  NANDN U7506 ( .A(n35611), .B(n7022), .Z(n7024) );
  XOR U7507 ( .A(b[35]), .B(a[20]), .Z(n7199) );
  NANDN U7508 ( .A(n35801), .B(n7199), .Z(n7023) );
  NAND U7509 ( .A(n7024), .B(n7023), .Z(n7238) );
  XNOR U7510 ( .A(n7239), .B(n7238), .Z(n7240) );
  XNOR U7511 ( .A(n7241), .B(n7240), .Z(n7250) );
  XNOR U7512 ( .A(n7251), .B(n7250), .Z(n7252) );
  XOR U7513 ( .A(n7253), .B(n7252), .Z(n7142) );
  XNOR U7514 ( .A(n7141), .B(n7142), .Z(n7163) );
  XNOR U7515 ( .A(n7164), .B(n7163), .Z(n7165) );
  XNOR U7516 ( .A(n7166), .B(n7165), .Z(n7078) );
  XOR U7517 ( .A(n7079), .B(n7078), .Z(n7081) );
  XOR U7518 ( .A(n7080), .B(n7081), .Z(n7305) );
  NANDN U7519 ( .A(n7026), .B(n7025), .Z(n7030) );
  NANDN U7520 ( .A(n7028), .B(n7027), .Z(n7029) );
  NAND U7521 ( .A(n7030), .B(n7029), .Z(n7304) );
  XOR U7522 ( .A(n7305), .B(n7304), .Z(n7307) );
  XOR U7523 ( .A(n7306), .B(n7307), .Z(n7067) );
  NANDN U7524 ( .A(n7032), .B(n7031), .Z(n7036) );
  NANDN U7525 ( .A(n7034), .B(n7033), .Z(n7035) );
  AND U7526 ( .A(n7036), .B(n7035), .Z(n7074) );
  NAND U7527 ( .A(n7038), .B(n7037), .Z(n7042) );
  NAND U7528 ( .A(n7040), .B(n7039), .Z(n7041) );
  AND U7529 ( .A(n7042), .B(n7041), .Z(n7073) );
  NANDN U7530 ( .A(n7044), .B(n7043), .Z(n7048) );
  NANDN U7531 ( .A(n7046), .B(n7045), .Z(n7047) );
  AND U7532 ( .A(n7048), .B(n7047), .Z(n7072) );
  XOR U7533 ( .A(n7073), .B(n7072), .Z(n7075) );
  XNOR U7534 ( .A(n7074), .B(n7075), .Z(n7066) );
  XOR U7535 ( .A(n7067), .B(n7066), .Z(n7069) );
  XOR U7536 ( .A(n7068), .B(n7069), .Z(n7061) );
  NANDN U7537 ( .A(n7050), .B(n7049), .Z(n7054) );
  NAND U7538 ( .A(n7052), .B(n7051), .Z(n7053) );
  AND U7539 ( .A(n7054), .B(n7053), .Z(n7060) );
  XNOR U7540 ( .A(n7061), .B(n7060), .Z(n7062) );
  XNOR U7541 ( .A(n7063), .B(n7062), .Z(n7056) );
  XNOR U7542 ( .A(n7057), .B(n7056), .Z(c[118]) );
  NANDN U7543 ( .A(sreg[118]), .B(n7055), .Z(n7059) );
  NAND U7544 ( .A(n7057), .B(n7056), .Z(n7058) );
  AND U7545 ( .A(n7059), .B(n7058), .Z(n7312) );
  NANDN U7546 ( .A(n7061), .B(n7060), .Z(n7065) );
  NANDN U7547 ( .A(n7063), .B(n7062), .Z(n7064) );
  AND U7548 ( .A(n7065), .B(n7064), .Z(n7317) );
  NANDN U7549 ( .A(n7067), .B(n7066), .Z(n7071) );
  OR U7550 ( .A(n7069), .B(n7068), .Z(n7070) );
  AND U7551 ( .A(n7071), .B(n7070), .Z(n7315) );
  NANDN U7552 ( .A(n7073), .B(n7072), .Z(n7077) );
  OR U7553 ( .A(n7075), .B(n7074), .Z(n7076) );
  AND U7554 ( .A(n7077), .B(n7076), .Z(n7324) );
  NANDN U7555 ( .A(n7079), .B(n7078), .Z(n7083) );
  OR U7556 ( .A(n7081), .B(n7080), .Z(n7082) );
  AND U7557 ( .A(n7083), .B(n7082), .Z(n7555) );
  NANDN U7558 ( .A(n7085), .B(n7084), .Z(n7089) );
  NANDN U7559 ( .A(n7087), .B(n7086), .Z(n7088) );
  AND U7560 ( .A(n7089), .B(n7088), .Z(n7347) );
  NANDN U7561 ( .A(n37705), .B(n7090), .Z(n7092) );
  XOR U7562 ( .A(b[53]), .B(a[3]), .Z(n7408) );
  NANDN U7563 ( .A(n37778), .B(n7408), .Z(n7091) );
  AND U7564 ( .A(n7092), .B(n7091), .Z(n7456) );
  XNOR U7565 ( .A(b[55]), .B(a[1]), .Z(n7459) );
  NANDN U7566 ( .A(n7459), .B(n37985), .Z(n7099) );
  ANDN U7567 ( .B(b[54]), .A(b[55]), .Z(n7093) );
  NAND U7568 ( .A(n7093), .B(a[0]), .Z(n7096) );
  NAND U7569 ( .A(b[53]), .B(b[54]), .Z(n7094) );
  NAND U7570 ( .A(b[55]), .B(n7094), .Z(n38038) );
  OR U7571 ( .A(a[0]), .B(n38038), .Z(n7095) );
  NAND U7572 ( .A(n7096), .B(n7095), .Z(n7097) );
  NAND U7573 ( .A(n37911), .B(n7097), .Z(n7098) );
  AND U7574 ( .A(n7099), .B(n7098), .Z(n7457) );
  XOR U7575 ( .A(n7456), .B(n7457), .Z(n7395) );
  NOR U7576 ( .A(n38038), .B(n7103), .Z(n7394) );
  NANDN U7577 ( .A(n7100), .B(n35001), .Z(n7102) );
  XNOR U7578 ( .A(b[29]), .B(a[27]), .Z(n7513) );
  NANDN U7579 ( .A(n7513), .B(n35002), .Z(n7101) );
  AND U7580 ( .A(n7102), .B(n7101), .Z(n7393) );
  XOR U7581 ( .A(n7394), .B(n7393), .Z(n7396) );
  XOR U7582 ( .A(n7395), .B(n7396), .Z(n7346) );
  NANDN U7583 ( .A(n7104), .B(n7103), .Z(n7108) );
  NANDN U7584 ( .A(n7106), .B(n7105), .Z(n7107) );
  NAND U7585 ( .A(n7108), .B(n7107), .Z(n7345) );
  XOR U7586 ( .A(n7346), .B(n7345), .Z(n7348) );
  XOR U7587 ( .A(n7347), .B(n7348), .Z(n7422) );
  NANDN U7588 ( .A(n7109), .B(n9942), .Z(n7111) );
  XOR U7589 ( .A(b[3]), .B(a[53]), .Z(n7507) );
  NANDN U7590 ( .A(n28941), .B(n7507), .Z(n7110) );
  AND U7591 ( .A(n7111), .B(n7110), .Z(n7446) );
  NAND U7592 ( .A(b[0]), .B(a[55]), .Z(n7112) );
  XNOR U7593 ( .A(b[1]), .B(n7112), .Z(n7114) );
  NANDN U7594 ( .A(b[0]), .B(a[54]), .Z(n7113) );
  NAND U7595 ( .A(n7114), .B(n7113), .Z(n7445) );
  NANDN U7596 ( .A(n34223), .B(n7115), .Z(n7117) );
  XOR U7597 ( .A(b[27]), .B(a[29]), .Z(n7489) );
  NANDN U7598 ( .A(n34458), .B(n7489), .Z(n7116) );
  NAND U7599 ( .A(n7117), .B(n7116), .Z(n7444) );
  XOR U7600 ( .A(n7445), .B(n7444), .Z(n7447) );
  XOR U7601 ( .A(n7446), .B(n7447), .Z(n7529) );
  NANDN U7602 ( .A(n31055), .B(n7118), .Z(n7120) );
  XOR U7603 ( .A(b[13]), .B(a[43]), .Z(n7375) );
  NANDN U7604 ( .A(n31293), .B(n7375), .Z(n7119) );
  AND U7605 ( .A(n7120), .B(n7119), .Z(n7494) );
  NANDN U7606 ( .A(n30482), .B(n7121), .Z(n7123) );
  XOR U7607 ( .A(b[11]), .B(a[45]), .Z(n7480) );
  NANDN U7608 ( .A(n30891), .B(n7480), .Z(n7122) );
  AND U7609 ( .A(n7123), .B(n7122), .Z(n7493) );
  NANDN U7610 ( .A(n36210), .B(n7124), .Z(n7126) );
  XOR U7611 ( .A(b[39]), .B(a[17]), .Z(n7372) );
  NANDN U7612 ( .A(n36347), .B(n7372), .Z(n7125) );
  NAND U7613 ( .A(n7126), .B(n7125), .Z(n7492) );
  XOR U7614 ( .A(n7493), .B(n7492), .Z(n7495) );
  XNOR U7615 ( .A(n7494), .B(n7495), .Z(n7528) );
  XNOR U7616 ( .A(n7529), .B(n7528), .Z(n7530) );
  NANDN U7617 ( .A(n7128), .B(n7127), .Z(n7132) );
  NANDN U7618 ( .A(n7130), .B(n7129), .Z(n7131) );
  NAND U7619 ( .A(n7132), .B(n7131), .Z(n7531) );
  XNOR U7620 ( .A(n7530), .B(n7531), .Z(n7420) );
  NANDN U7621 ( .A(n7134), .B(n7133), .Z(n7138) );
  NANDN U7622 ( .A(n7136), .B(n7135), .Z(n7137) );
  NAND U7623 ( .A(n7138), .B(n7137), .Z(n7421) );
  XOR U7624 ( .A(n7420), .B(n7421), .Z(n7423) );
  XOR U7625 ( .A(n7422), .B(n7423), .Z(n7536) );
  NANDN U7626 ( .A(n7140), .B(n7139), .Z(n7144) );
  NANDN U7627 ( .A(n7142), .B(n7141), .Z(n7143) );
  AND U7628 ( .A(n7144), .B(n7143), .Z(n7535) );
  NANDN U7629 ( .A(n7146), .B(n7145), .Z(n7150) );
  NAND U7630 ( .A(n7148), .B(n7147), .Z(n7149) );
  AND U7631 ( .A(n7150), .B(n7149), .Z(n7534) );
  XOR U7632 ( .A(n7535), .B(n7534), .Z(n7537) );
  XOR U7633 ( .A(n7536), .B(n7537), .Z(n7553) );
  NANDN U7634 ( .A(n7152), .B(n7151), .Z(n7156) );
  NANDN U7635 ( .A(n7154), .B(n7153), .Z(n7155) );
  AND U7636 ( .A(n7156), .B(n7155), .Z(n7552) );
  XNOR U7637 ( .A(n7553), .B(n7552), .Z(n7554) );
  XOR U7638 ( .A(n7555), .B(n7554), .Z(n7560) );
  NANDN U7639 ( .A(n7158), .B(n7157), .Z(n7162) );
  NAND U7640 ( .A(n7160), .B(n7159), .Z(n7161) );
  AND U7641 ( .A(n7162), .B(n7161), .Z(n7559) );
  NANDN U7642 ( .A(n7164), .B(n7163), .Z(n7168) );
  NANDN U7643 ( .A(n7166), .B(n7165), .Z(n7167) );
  AND U7644 ( .A(n7168), .B(n7167), .Z(n7336) );
  NANDN U7645 ( .A(n7170), .B(n7169), .Z(n7174) );
  NAND U7646 ( .A(n7172), .B(n7171), .Z(n7173) );
  AND U7647 ( .A(n7174), .B(n7173), .Z(n7542) );
  NANDN U7648 ( .A(n7176), .B(n7175), .Z(n7180) );
  NANDN U7649 ( .A(n7178), .B(n7177), .Z(n7179) );
  AND U7650 ( .A(n7180), .B(n7179), .Z(n7540) );
  NANDN U7651 ( .A(n7182), .B(n7181), .Z(n7186) );
  NAND U7652 ( .A(n7184), .B(n7183), .Z(n7185) );
  NAND U7653 ( .A(n7186), .B(n7185), .Z(n7541) );
  XOR U7654 ( .A(n7540), .B(n7541), .Z(n7543) );
  XOR U7655 ( .A(n7542), .B(n7543), .Z(n7334) );
  NANDN U7656 ( .A(n7188), .B(n7187), .Z(n7192) );
  OR U7657 ( .A(n7190), .B(n7189), .Z(n7191) );
  AND U7658 ( .A(n7192), .B(n7191), .Z(n7427) );
  NANDN U7659 ( .A(n210), .B(n7193), .Z(n7195) );
  XOR U7660 ( .A(b[9]), .B(a[47]), .Z(n7378) );
  NANDN U7661 ( .A(n30267), .B(n7378), .Z(n7194) );
  AND U7662 ( .A(n7195), .B(n7194), .Z(n7389) );
  NANDN U7663 ( .A(n29499), .B(n7196), .Z(n7198) );
  XOR U7664 ( .A(b[7]), .B(a[49]), .Z(n7486) );
  NANDN U7665 ( .A(n29735), .B(n7486), .Z(n7197) );
  AND U7666 ( .A(n7198), .B(n7197), .Z(n7388) );
  NANDN U7667 ( .A(n35611), .B(n7199), .Z(n7201) );
  XOR U7668 ( .A(b[35]), .B(a[21]), .Z(n7384) );
  NANDN U7669 ( .A(n35801), .B(n7384), .Z(n7200) );
  NAND U7670 ( .A(n7201), .B(n7200), .Z(n7387) );
  XOR U7671 ( .A(n7388), .B(n7387), .Z(n7390) );
  XOR U7672 ( .A(n7389), .B(n7390), .Z(n7352) );
  NANDN U7673 ( .A(n32013), .B(n7202), .Z(n7204) );
  XOR U7674 ( .A(b[17]), .B(a[39]), .Z(n7414) );
  NANDN U7675 ( .A(n32292), .B(n7414), .Z(n7203) );
  AND U7676 ( .A(n7204), .B(n7203), .Z(n7518) );
  NANDN U7677 ( .A(n31536), .B(n7205), .Z(n7207) );
  XOR U7678 ( .A(b[15]), .B(a[41]), .Z(n7471) );
  NANDN U7679 ( .A(n31925), .B(n7471), .Z(n7206) );
  AND U7680 ( .A(n7207), .B(n7206), .Z(n7517) );
  NANDN U7681 ( .A(n212), .B(n7208), .Z(n7210) );
  XOR U7682 ( .A(b[49]), .B(a[7]), .Z(n7501) );
  NANDN U7683 ( .A(n37432), .B(n7501), .Z(n7209) );
  NAND U7684 ( .A(n7210), .B(n7209), .Z(n7516) );
  XOR U7685 ( .A(n7517), .B(n7516), .Z(n7519) );
  XNOR U7686 ( .A(n7518), .B(n7519), .Z(n7351) );
  XNOR U7687 ( .A(n7352), .B(n7351), .Z(n7354) );
  NANDN U7688 ( .A(n7212), .B(n7211), .Z(n7216) );
  OR U7689 ( .A(n7214), .B(n7213), .Z(n7215) );
  AND U7690 ( .A(n7216), .B(n7215), .Z(n7353) );
  XNOR U7691 ( .A(n7354), .B(n7353), .Z(n7426) );
  XNOR U7692 ( .A(n7427), .B(n7426), .Z(n7428) );
  NANDN U7693 ( .A(n36480), .B(n7217), .Z(n7219) );
  XOR U7694 ( .A(b[41]), .B(a[15]), .Z(n7474) );
  NANDN U7695 ( .A(n36594), .B(n7474), .Z(n7218) );
  AND U7696 ( .A(n7219), .B(n7218), .Z(n7401) );
  NANDN U7697 ( .A(n36742), .B(n7220), .Z(n7222) );
  XOR U7698 ( .A(b[43]), .B(a[13]), .Z(n7477) );
  NANDN U7699 ( .A(n36891), .B(n7477), .Z(n7221) );
  AND U7700 ( .A(n7222), .B(n7221), .Z(n7400) );
  NANDN U7701 ( .A(n32996), .B(n7223), .Z(n7225) );
  XOR U7702 ( .A(b[21]), .B(a[35]), .Z(n7417) );
  NANDN U7703 ( .A(n33271), .B(n7417), .Z(n7224) );
  NAND U7704 ( .A(n7225), .B(n7224), .Z(n7399) );
  XOR U7705 ( .A(n7400), .B(n7399), .Z(n7402) );
  XOR U7706 ( .A(n7401), .B(n7402), .Z(n7359) );
  NANDN U7707 ( .A(n35936), .B(n7226), .Z(n7228) );
  XOR U7708 ( .A(b[37]), .B(a[19]), .Z(n7369) );
  NANDN U7709 ( .A(n36047), .B(n7369), .Z(n7227) );
  AND U7710 ( .A(n7228), .B(n7227), .Z(n7452) );
  NANDN U7711 ( .A(n33866), .B(n7229), .Z(n7231) );
  XOR U7712 ( .A(b[23]), .B(a[33]), .Z(n7465) );
  NANDN U7713 ( .A(n33644), .B(n7465), .Z(n7230) );
  AND U7714 ( .A(n7231), .B(n7230), .Z(n7451) );
  NANDN U7715 ( .A(n34909), .B(n7232), .Z(n7234) );
  XOR U7716 ( .A(b[31]), .B(a[25]), .Z(n7462) );
  NANDN U7717 ( .A(n35145), .B(n7462), .Z(n7233) );
  NAND U7718 ( .A(n7234), .B(n7233), .Z(n7450) );
  XOR U7719 ( .A(n7451), .B(n7450), .Z(n7453) );
  XOR U7720 ( .A(n7452), .B(n7453), .Z(n7358) );
  NAND U7721 ( .A(n34297), .B(n7235), .Z(n7237) );
  XNOR U7722 ( .A(b[25]), .B(a[31]), .Z(n7468) );
  NANDN U7723 ( .A(n7468), .B(n34298), .Z(n7236) );
  AND U7724 ( .A(n7237), .B(n7236), .Z(n7357) );
  XOR U7725 ( .A(n7358), .B(n7357), .Z(n7360) );
  XOR U7726 ( .A(n7359), .B(n7360), .Z(n7342) );
  NANDN U7727 ( .A(n7239), .B(n7238), .Z(n7243) );
  NANDN U7728 ( .A(n7241), .B(n7240), .Z(n7242) );
  AND U7729 ( .A(n7243), .B(n7242), .Z(n7340) );
  NANDN U7730 ( .A(n7245), .B(n7244), .Z(n7249) );
  OR U7731 ( .A(n7247), .B(n7246), .Z(n7248) );
  NAND U7732 ( .A(n7249), .B(n7248), .Z(n7339) );
  XNOR U7733 ( .A(n7340), .B(n7339), .Z(n7341) );
  XOR U7734 ( .A(n7342), .B(n7341), .Z(n7429) );
  XNOR U7735 ( .A(n7428), .B(n7429), .Z(n7549) );
  NANDN U7736 ( .A(n7251), .B(n7250), .Z(n7255) );
  NANDN U7737 ( .A(n7253), .B(n7252), .Z(n7254) );
  AND U7738 ( .A(n7255), .B(n7254), .Z(n7547) );
  NANDN U7739 ( .A(n37526), .B(n7256), .Z(n7258) );
  XOR U7740 ( .A(b[51]), .B(a[5]), .Z(n7510) );
  NANDN U7741 ( .A(n37605), .B(n7510), .Z(n7257) );
  AND U7742 ( .A(n7258), .B(n7257), .Z(n7440) );
  NANDN U7743 ( .A(n28889), .B(n7259), .Z(n7261) );
  XOR U7744 ( .A(b[5]), .B(a[51]), .Z(n7498) );
  NANDN U7745 ( .A(n29138), .B(n7498), .Z(n7260) );
  AND U7746 ( .A(n7261), .B(n7260), .Z(n7439) );
  NANDN U7747 ( .A(n35260), .B(n7262), .Z(n7264) );
  XOR U7748 ( .A(b[33]), .B(a[23]), .Z(n7504) );
  NANDN U7749 ( .A(n35456), .B(n7504), .Z(n7263) );
  NAND U7750 ( .A(n7264), .B(n7263), .Z(n7438) );
  XOR U7751 ( .A(n7439), .B(n7438), .Z(n7441) );
  XOR U7752 ( .A(n7440), .B(n7441), .Z(n7523) );
  NANDN U7753 ( .A(n36991), .B(n7265), .Z(n7267) );
  XOR U7754 ( .A(b[45]), .B(a[11]), .Z(n7381) );
  NANDN U7755 ( .A(n37083), .B(n7381), .Z(n7266) );
  AND U7756 ( .A(n7267), .B(n7266), .Z(n7365) );
  NANDN U7757 ( .A(n211), .B(n7268), .Z(n7270) );
  XOR U7758 ( .A(b[47]), .B(a[9]), .Z(n7483) );
  NANDN U7759 ( .A(n37172), .B(n7483), .Z(n7269) );
  AND U7760 ( .A(n7270), .B(n7269), .Z(n7364) );
  NANDN U7761 ( .A(n32483), .B(n7271), .Z(n7273) );
  XOR U7762 ( .A(b[19]), .B(a[37]), .Z(n7411) );
  NANDN U7763 ( .A(n32823), .B(n7411), .Z(n7272) );
  NAND U7764 ( .A(n7273), .B(n7272), .Z(n7363) );
  XOR U7765 ( .A(n7364), .B(n7363), .Z(n7366) );
  XNOR U7766 ( .A(n7365), .B(n7366), .Z(n7522) );
  XNOR U7767 ( .A(n7523), .B(n7522), .Z(n7525) );
  NANDN U7768 ( .A(n7275), .B(n7274), .Z(n7279) );
  OR U7769 ( .A(n7277), .B(n7276), .Z(n7278) );
  AND U7770 ( .A(n7279), .B(n7278), .Z(n7524) );
  XOR U7771 ( .A(n7525), .B(n7524), .Z(n7435) );
  NANDN U7772 ( .A(n7281), .B(n7280), .Z(n7285) );
  OR U7773 ( .A(n7283), .B(n7282), .Z(n7284) );
  AND U7774 ( .A(n7285), .B(n7284), .Z(n7433) );
  NANDN U7775 ( .A(n7287), .B(n7286), .Z(n7291) );
  OR U7776 ( .A(n7289), .B(n7288), .Z(n7290) );
  AND U7777 ( .A(n7291), .B(n7290), .Z(n7432) );
  XNOR U7778 ( .A(n7433), .B(n7432), .Z(n7434) );
  XNOR U7779 ( .A(n7435), .B(n7434), .Z(n7546) );
  XNOR U7780 ( .A(n7547), .B(n7546), .Z(n7548) );
  XNOR U7781 ( .A(n7549), .B(n7548), .Z(n7333) );
  XNOR U7782 ( .A(n7334), .B(n7333), .Z(n7335) );
  XOR U7783 ( .A(n7336), .B(n7335), .Z(n7330) );
  NANDN U7784 ( .A(n7293), .B(n7292), .Z(n7297) );
  NAND U7785 ( .A(n7295), .B(n7294), .Z(n7296) );
  AND U7786 ( .A(n7297), .B(n7296), .Z(n7327) );
  NANDN U7787 ( .A(n7299), .B(n7298), .Z(n7303) );
  OR U7788 ( .A(n7301), .B(n7300), .Z(n7302) );
  NAND U7789 ( .A(n7303), .B(n7302), .Z(n7328) );
  XNOR U7790 ( .A(n7327), .B(n7328), .Z(n7329) );
  XNOR U7791 ( .A(n7330), .B(n7329), .Z(n7558) );
  XOR U7792 ( .A(n7559), .B(n7558), .Z(n7561) );
  XOR U7793 ( .A(n7560), .B(n7561), .Z(n7322) );
  NANDN U7794 ( .A(n7305), .B(n7304), .Z(n7309) );
  OR U7795 ( .A(n7307), .B(n7306), .Z(n7308) );
  NAND U7796 ( .A(n7309), .B(n7308), .Z(n7321) );
  XNOR U7797 ( .A(n7322), .B(n7321), .Z(n7323) );
  XOR U7798 ( .A(n7324), .B(n7323), .Z(n7316) );
  XOR U7799 ( .A(n7315), .B(n7316), .Z(n7318) );
  XOR U7800 ( .A(n7317), .B(n7318), .Z(n7310) );
  XNOR U7801 ( .A(n7310), .B(sreg[119]), .Z(n7311) );
  XOR U7802 ( .A(n7312), .B(n7311), .Z(c[119]) );
  NANDN U7803 ( .A(n7310), .B(sreg[119]), .Z(n7314) );
  NAND U7804 ( .A(n7312), .B(n7311), .Z(n7313) );
  AND U7805 ( .A(n7314), .B(n7313), .Z(n7821) );
  XNOR U7806 ( .A(sreg[120]), .B(n7821), .Z(n7823) );
  NANDN U7807 ( .A(n7316), .B(n7315), .Z(n7320) );
  OR U7808 ( .A(n7318), .B(n7317), .Z(n7319) );
  AND U7809 ( .A(n7320), .B(n7319), .Z(n7567) );
  NANDN U7810 ( .A(n7322), .B(n7321), .Z(n7326) );
  NANDN U7811 ( .A(n7324), .B(n7323), .Z(n7325) );
  AND U7812 ( .A(n7326), .B(n7325), .Z(n7565) );
  NANDN U7813 ( .A(n7328), .B(n7327), .Z(n7332) );
  NANDN U7814 ( .A(n7330), .B(n7329), .Z(n7331) );
  AND U7815 ( .A(n7332), .B(n7331), .Z(n7816) );
  NANDN U7816 ( .A(n7334), .B(n7333), .Z(n7338) );
  NAND U7817 ( .A(n7336), .B(n7335), .Z(n7337) );
  AND U7818 ( .A(n7338), .B(n7337), .Z(n7815) );
  XNOR U7819 ( .A(n7816), .B(n7815), .Z(n7818) );
  NANDN U7820 ( .A(n7340), .B(n7339), .Z(n7344) );
  NANDN U7821 ( .A(n7342), .B(n7341), .Z(n7343) );
  AND U7822 ( .A(n7344), .B(n7343), .Z(n7584) );
  NANDN U7823 ( .A(n7346), .B(n7345), .Z(n7350) );
  OR U7824 ( .A(n7348), .B(n7347), .Z(n7349) );
  AND U7825 ( .A(n7350), .B(n7349), .Z(n7583) );
  NANDN U7826 ( .A(n7352), .B(n7351), .Z(n7356) );
  NAND U7827 ( .A(n7354), .B(n7353), .Z(n7355) );
  AND U7828 ( .A(n7356), .B(n7355), .Z(n7582) );
  XOR U7829 ( .A(n7583), .B(n7582), .Z(n7585) );
  XOR U7830 ( .A(n7584), .B(n7585), .Z(n7664) );
  NANDN U7831 ( .A(n7358), .B(n7357), .Z(n7362) );
  OR U7832 ( .A(n7360), .B(n7359), .Z(n7361) );
  AND U7833 ( .A(n7362), .B(n7361), .Z(n7597) );
  NANDN U7834 ( .A(n7364), .B(n7363), .Z(n7368) );
  OR U7835 ( .A(n7366), .B(n7365), .Z(n7367) );
  AND U7836 ( .A(n7368), .B(n7367), .Z(n7695) );
  NANDN U7837 ( .A(n35936), .B(n7369), .Z(n7371) );
  XOR U7838 ( .A(b[37]), .B(a[20]), .Z(n7735) );
  NANDN U7839 ( .A(n36047), .B(n7735), .Z(n7370) );
  AND U7840 ( .A(n7371), .B(n7370), .Z(n7770) );
  NANDN U7841 ( .A(n36210), .B(n7372), .Z(n7374) );
  XOR U7842 ( .A(b[39]), .B(a[18]), .Z(n7642) );
  NANDN U7843 ( .A(n36347), .B(n7642), .Z(n7373) );
  AND U7844 ( .A(n7374), .B(n7373), .Z(n7768) );
  NANDN U7845 ( .A(n31055), .B(n7375), .Z(n7377) );
  XOR U7846 ( .A(b[13]), .B(a[44]), .Z(n7636) );
  NANDN U7847 ( .A(n31293), .B(n7636), .Z(n7376) );
  NAND U7848 ( .A(n7377), .B(n7376), .Z(n7767) );
  XNOR U7849 ( .A(n7768), .B(n7767), .Z(n7769) );
  XOR U7850 ( .A(n7770), .B(n7769), .Z(n7693) );
  NANDN U7851 ( .A(n210), .B(n7378), .Z(n7380) );
  XOR U7852 ( .A(b[9]), .B(a[48]), .Z(n7750) );
  NANDN U7853 ( .A(n30267), .B(n7750), .Z(n7379) );
  AND U7854 ( .A(n7380), .B(n7379), .Z(n7799) );
  NANDN U7855 ( .A(n36991), .B(n7381), .Z(n7383) );
  XOR U7856 ( .A(b[45]), .B(a[12]), .Z(n7782) );
  NANDN U7857 ( .A(n37083), .B(n7782), .Z(n7382) );
  AND U7858 ( .A(n7383), .B(n7382), .Z(n7798) );
  NANDN U7859 ( .A(n35611), .B(n7384), .Z(n7386) );
  XOR U7860 ( .A(b[35]), .B(a[22]), .Z(n7756) );
  NANDN U7861 ( .A(n35801), .B(n7756), .Z(n7385) );
  NAND U7862 ( .A(n7386), .B(n7385), .Z(n7797) );
  XOR U7863 ( .A(n7798), .B(n7797), .Z(n7800) );
  XNOR U7864 ( .A(n7799), .B(n7800), .Z(n7692) );
  XOR U7865 ( .A(n7693), .B(n7692), .Z(n7694) );
  XOR U7866 ( .A(n7695), .B(n7694), .Z(n7595) );
  NANDN U7867 ( .A(n7388), .B(n7387), .Z(n7392) );
  OR U7868 ( .A(n7390), .B(n7389), .Z(n7391) );
  AND U7869 ( .A(n7392), .B(n7391), .Z(n7601) );
  NANDN U7870 ( .A(n7394), .B(n7393), .Z(n7398) );
  OR U7871 ( .A(n7396), .B(n7395), .Z(n7397) );
  AND U7872 ( .A(n7398), .B(n7397), .Z(n7600) );
  XNOR U7873 ( .A(n7601), .B(n7600), .Z(n7602) );
  NANDN U7874 ( .A(n7400), .B(n7399), .Z(n7404) );
  OR U7875 ( .A(n7402), .B(n7401), .Z(n7403) );
  AND U7876 ( .A(n7404), .B(n7403), .Z(n7609) );
  NAND U7877 ( .A(b[0]), .B(a[56]), .Z(n7405) );
  XNOR U7878 ( .A(b[1]), .B(n7405), .Z(n7407) );
  NANDN U7879 ( .A(b[0]), .B(a[55]), .Z(n7406) );
  NAND U7880 ( .A(n7407), .B(n7406), .Z(n7653) );
  XOR U7881 ( .A(b[56]), .B(b[55]), .Z(n38077) );
  IV U7882 ( .A(n38077), .Z(n38031) );
  ANDN U7883 ( .B(a[0]), .A(n38031), .Z(n7766) );
  NANDN U7884 ( .A(n37705), .B(n7408), .Z(n7410) );
  XOR U7885 ( .A(b[53]), .B(a[4]), .Z(n7779) );
  NANDN U7886 ( .A(n37778), .B(n7779), .Z(n7409) );
  AND U7887 ( .A(n7410), .B(n7409), .Z(n7651) );
  XNOR U7888 ( .A(n7766), .B(n7651), .Z(n7652) );
  XNOR U7889 ( .A(n7653), .B(n7652), .Z(n7606) );
  NANDN U7890 ( .A(n32483), .B(n7411), .Z(n7413) );
  XOR U7891 ( .A(b[19]), .B(a[38]), .Z(n7618) );
  NANDN U7892 ( .A(n32823), .B(n7618), .Z(n7412) );
  AND U7893 ( .A(n7413), .B(n7412), .Z(n7648) );
  NANDN U7894 ( .A(n32013), .B(n7414), .Z(n7416) );
  XOR U7895 ( .A(b[17]), .B(a[40]), .Z(n7741) );
  NANDN U7896 ( .A(n32292), .B(n7741), .Z(n7415) );
  AND U7897 ( .A(n7416), .B(n7415), .Z(n7646) );
  NANDN U7898 ( .A(n32996), .B(n7417), .Z(n7419) );
  XOR U7899 ( .A(b[21]), .B(a[36]), .Z(n7612) );
  NANDN U7900 ( .A(n33271), .B(n7612), .Z(n7418) );
  NAND U7901 ( .A(n7419), .B(n7418), .Z(n7645) );
  XNOR U7902 ( .A(n7646), .B(n7645), .Z(n7647) );
  XOR U7903 ( .A(n7648), .B(n7647), .Z(n7607) );
  XNOR U7904 ( .A(n7606), .B(n7607), .Z(n7608) );
  XOR U7905 ( .A(n7609), .B(n7608), .Z(n7603) );
  XNOR U7906 ( .A(n7602), .B(n7603), .Z(n7594) );
  XNOR U7907 ( .A(n7595), .B(n7594), .Z(n7596) );
  XOR U7908 ( .A(n7597), .B(n7596), .Z(n7663) );
  NANDN U7909 ( .A(n7421), .B(n7420), .Z(n7425) );
  OR U7910 ( .A(n7423), .B(n7422), .Z(n7424) );
  NAND U7911 ( .A(n7425), .B(n7424), .Z(n7662) );
  XOR U7912 ( .A(n7663), .B(n7662), .Z(n7665) );
  XOR U7913 ( .A(n7664), .B(n7665), .Z(n7810) );
  NANDN U7914 ( .A(n7427), .B(n7426), .Z(n7431) );
  NANDN U7915 ( .A(n7429), .B(n7428), .Z(n7430) );
  AND U7916 ( .A(n7431), .B(n7430), .Z(n7671) );
  NANDN U7917 ( .A(n7433), .B(n7432), .Z(n7437) );
  NANDN U7918 ( .A(n7435), .B(n7434), .Z(n7436) );
  AND U7919 ( .A(n7437), .B(n7436), .Z(n7669) );
  NANDN U7920 ( .A(n7439), .B(n7438), .Z(n7443) );
  OR U7921 ( .A(n7441), .B(n7440), .Z(n7442) );
  AND U7922 ( .A(n7443), .B(n7442), .Z(n7687) );
  NANDN U7923 ( .A(n7445), .B(n7444), .Z(n7449) );
  OR U7924 ( .A(n7447), .B(n7446), .Z(n7448) );
  NAND U7925 ( .A(n7449), .B(n7448), .Z(n7686) );
  XNOR U7926 ( .A(n7687), .B(n7686), .Z(n7689) );
  NANDN U7927 ( .A(n7451), .B(n7450), .Z(n7455) );
  OR U7928 ( .A(n7453), .B(n7452), .Z(n7454) );
  NAND U7929 ( .A(n7455), .B(n7454), .Z(n7700) );
  OR U7930 ( .A(n7457), .B(n7456), .Z(n7806) );
  XOR U7931 ( .A(b[54]), .B(b[55]), .Z(n7458) );
  ANDN U7932 ( .B(n7458), .A(n37985), .Z(n37984) );
  NANDN U7933 ( .A(n7459), .B(n37984), .Z(n7461) );
  XNOR U7934 ( .A(b[55]), .B(a[2]), .Z(n7722) );
  NANDN U7935 ( .A(n7722), .B(n37985), .Z(n7460) );
  AND U7936 ( .A(n7461), .B(n7460), .Z(n7804) );
  NANDN U7937 ( .A(n34909), .B(n7462), .Z(n7464) );
  XOR U7938 ( .A(b[31]), .B(a[26]), .Z(n7732) );
  NANDN U7939 ( .A(n35145), .B(n7732), .Z(n7463) );
  AND U7940 ( .A(n7464), .B(n7463), .Z(n7803) );
  XOR U7941 ( .A(n7804), .B(n7803), .Z(n7805) );
  XNOR U7942 ( .A(n7806), .B(n7805), .Z(n7699) );
  NANDN U7943 ( .A(n33866), .B(n7465), .Z(n7467) );
  XOR U7944 ( .A(b[23]), .B(a[34]), .Z(n7624) );
  NANDN U7945 ( .A(n33644), .B(n7624), .Z(n7466) );
  AND U7946 ( .A(n7467), .B(n7466), .Z(n7794) );
  NANDN U7947 ( .A(n7468), .B(n34297), .Z(n7470) );
  XOR U7948 ( .A(b[25]), .B(a[32]), .Z(n7615) );
  NANDN U7949 ( .A(n33994), .B(n7615), .Z(n7469) );
  AND U7950 ( .A(n7470), .B(n7469), .Z(n7792) );
  NANDN U7951 ( .A(n31536), .B(n7471), .Z(n7473) );
  XOR U7952 ( .A(b[15]), .B(a[42]), .Z(n7788) );
  NANDN U7953 ( .A(n31925), .B(n7788), .Z(n7472) );
  NAND U7954 ( .A(n7473), .B(n7472), .Z(n7791) );
  XNOR U7955 ( .A(n7792), .B(n7791), .Z(n7793) );
  XNOR U7956 ( .A(n7794), .B(n7793), .Z(n7698) );
  XOR U7957 ( .A(n7699), .B(n7698), .Z(n7701) );
  XOR U7958 ( .A(n7700), .B(n7701), .Z(n7688) );
  XOR U7959 ( .A(n7689), .B(n7688), .Z(n7658) );
  NANDN U7960 ( .A(n36480), .B(n7474), .Z(n7476) );
  XOR U7961 ( .A(b[41]), .B(a[16]), .Z(n7738) );
  NANDN U7962 ( .A(n36594), .B(n7738), .Z(n7475) );
  AND U7963 ( .A(n7476), .B(n7475), .Z(n7718) );
  NANDN U7964 ( .A(n36742), .B(n7477), .Z(n7479) );
  XOR U7965 ( .A(b[43]), .B(a[14]), .Z(n7633) );
  NANDN U7966 ( .A(n36891), .B(n7633), .Z(n7478) );
  AND U7967 ( .A(n7479), .B(n7478), .Z(n7717) );
  NANDN U7968 ( .A(n30482), .B(n7480), .Z(n7482) );
  XOR U7969 ( .A(b[11]), .B(a[46]), .Z(n7639) );
  NANDN U7970 ( .A(n30891), .B(n7639), .Z(n7481) );
  NAND U7971 ( .A(n7482), .B(n7481), .Z(n7716) );
  XOR U7972 ( .A(n7717), .B(n7716), .Z(n7719) );
  XOR U7973 ( .A(n7718), .B(n7719), .Z(n7675) );
  NANDN U7974 ( .A(n211), .B(n7483), .Z(n7485) );
  XOR U7975 ( .A(b[47]), .B(a[10]), .Z(n7785) );
  NANDN U7976 ( .A(n37172), .B(n7785), .Z(n7484) );
  AND U7977 ( .A(n7485), .B(n7484), .Z(n7706) );
  NANDN U7978 ( .A(n29499), .B(n7486), .Z(n7488) );
  XOR U7979 ( .A(b[7]), .B(a[50]), .Z(n7753) );
  NANDN U7980 ( .A(n29735), .B(n7753), .Z(n7487) );
  AND U7981 ( .A(n7488), .B(n7487), .Z(n7705) );
  NANDN U7982 ( .A(n34223), .B(n7489), .Z(n7491) );
  XOR U7983 ( .A(b[27]), .B(a[30]), .Z(n7621) );
  NANDN U7984 ( .A(n34458), .B(n7621), .Z(n7490) );
  NAND U7985 ( .A(n7491), .B(n7490), .Z(n7704) );
  XOR U7986 ( .A(n7705), .B(n7704), .Z(n7707) );
  XNOR U7987 ( .A(n7706), .B(n7707), .Z(n7674) );
  XNOR U7988 ( .A(n7675), .B(n7674), .Z(n7676) );
  NANDN U7989 ( .A(n7493), .B(n7492), .Z(n7497) );
  OR U7990 ( .A(n7495), .B(n7494), .Z(n7496) );
  NAND U7991 ( .A(n7497), .B(n7496), .Z(n7677) );
  XNOR U7992 ( .A(n7676), .B(n7677), .Z(n7656) );
  NAND U7993 ( .A(n29551), .B(n7498), .Z(n7500) );
  XNOR U7994 ( .A(b[5]), .B(a[52]), .Z(n7776) );
  NANDN U7995 ( .A(n7776), .B(n29552), .Z(n7499) );
  NAND U7996 ( .A(n7500), .B(n7499), .Z(n7746) );
  NAND U7997 ( .A(n37536), .B(n7501), .Z(n7503) );
  XNOR U7998 ( .A(b[49]), .B(a[8]), .Z(n7627) );
  NANDN U7999 ( .A(n7627), .B(n37537), .Z(n7502) );
  NAND U8000 ( .A(n7503), .B(n7502), .Z(n7745) );
  NAND U8001 ( .A(n35654), .B(n7504), .Z(n7506) );
  XNOR U8002 ( .A(b[33]), .B(a[24]), .Z(n7762) );
  NANDN U8003 ( .A(n7762), .B(n35655), .Z(n7505) );
  NAND U8004 ( .A(n7506), .B(n7505), .Z(n7744) );
  XOR U8005 ( .A(n7745), .B(n7744), .Z(n7747) );
  XNOR U8006 ( .A(n7746), .B(n7747), .Z(n7681) );
  NANDN U8007 ( .A(n209), .B(n7507), .Z(n7509) );
  XOR U8008 ( .A(b[3]), .B(a[54]), .Z(n7759) );
  NANDN U8009 ( .A(n28941), .B(n7759), .Z(n7508) );
  AND U8010 ( .A(n7509), .B(n7508), .Z(n7712) );
  NANDN U8011 ( .A(n37526), .B(n7510), .Z(n7512) );
  XOR U8012 ( .A(b[51]), .B(a[6]), .Z(n7630) );
  NANDN U8013 ( .A(n37605), .B(n7630), .Z(n7511) );
  AND U8014 ( .A(n7512), .B(n7511), .Z(n7711) );
  NANDN U8015 ( .A(n7513), .B(n35001), .Z(n7515) );
  XOR U8016 ( .A(b[29]), .B(a[28]), .Z(n7773) );
  NANDN U8017 ( .A(n34722), .B(n7773), .Z(n7514) );
  NAND U8018 ( .A(n7515), .B(n7514), .Z(n7710) );
  XOR U8019 ( .A(n7711), .B(n7710), .Z(n7713) );
  XNOR U8020 ( .A(n7712), .B(n7713), .Z(n7680) );
  XOR U8021 ( .A(n7681), .B(n7680), .Z(n7682) );
  NANDN U8022 ( .A(n7517), .B(n7516), .Z(n7521) );
  OR U8023 ( .A(n7519), .B(n7518), .Z(n7520) );
  NAND U8024 ( .A(n7521), .B(n7520), .Z(n7683) );
  XOR U8025 ( .A(n7682), .B(n7683), .Z(n7657) );
  XOR U8026 ( .A(n7656), .B(n7657), .Z(n7659) );
  XOR U8027 ( .A(n7658), .B(n7659), .Z(n7591) );
  NANDN U8028 ( .A(n7523), .B(n7522), .Z(n7527) );
  NAND U8029 ( .A(n7525), .B(n7524), .Z(n7526) );
  AND U8030 ( .A(n7527), .B(n7526), .Z(n7588) );
  NANDN U8031 ( .A(n7529), .B(n7528), .Z(n7533) );
  NANDN U8032 ( .A(n7531), .B(n7530), .Z(n7532) );
  NAND U8033 ( .A(n7533), .B(n7532), .Z(n7589) );
  XNOR U8034 ( .A(n7588), .B(n7589), .Z(n7590) );
  XNOR U8035 ( .A(n7591), .B(n7590), .Z(n7668) );
  XNOR U8036 ( .A(n7669), .B(n7668), .Z(n7670) );
  XNOR U8037 ( .A(n7671), .B(n7670), .Z(n7809) );
  XNOR U8038 ( .A(n7810), .B(n7809), .Z(n7811) );
  NANDN U8039 ( .A(n7535), .B(n7534), .Z(n7539) );
  OR U8040 ( .A(n7537), .B(n7536), .Z(n7538) );
  AND U8041 ( .A(n7539), .B(n7538), .Z(n7579) );
  NANDN U8042 ( .A(n7541), .B(n7540), .Z(n7545) );
  OR U8043 ( .A(n7543), .B(n7542), .Z(n7544) );
  AND U8044 ( .A(n7545), .B(n7544), .Z(n7577) );
  NANDN U8045 ( .A(n7547), .B(n7546), .Z(n7551) );
  NAND U8046 ( .A(n7549), .B(n7548), .Z(n7550) );
  NAND U8047 ( .A(n7551), .B(n7550), .Z(n7576) );
  XNOR U8048 ( .A(n7577), .B(n7576), .Z(n7578) );
  XOR U8049 ( .A(n7579), .B(n7578), .Z(n7812) );
  XNOR U8050 ( .A(n7811), .B(n7812), .Z(n7817) );
  XOR U8051 ( .A(n7818), .B(n7817), .Z(n7571) );
  NANDN U8052 ( .A(n7553), .B(n7552), .Z(n7557) );
  NAND U8053 ( .A(n7555), .B(n7554), .Z(n7556) );
  NAND U8054 ( .A(n7557), .B(n7556), .Z(n7570) );
  XNOR U8055 ( .A(n7571), .B(n7570), .Z(n7572) );
  NANDN U8056 ( .A(n7559), .B(n7558), .Z(n7563) );
  OR U8057 ( .A(n7561), .B(n7560), .Z(n7562) );
  NAND U8058 ( .A(n7563), .B(n7562), .Z(n7573) );
  XNOR U8059 ( .A(n7572), .B(n7573), .Z(n7564) );
  XNOR U8060 ( .A(n7565), .B(n7564), .Z(n7566) );
  XNOR U8061 ( .A(n7567), .B(n7566), .Z(n7822) );
  XNOR U8062 ( .A(n7823), .B(n7822), .Z(c[120]) );
  NANDN U8063 ( .A(n7565), .B(n7564), .Z(n7569) );
  NANDN U8064 ( .A(n7567), .B(n7566), .Z(n7568) );
  AND U8065 ( .A(n7569), .B(n7568), .Z(n7834) );
  NANDN U8066 ( .A(n7571), .B(n7570), .Z(n7575) );
  NANDN U8067 ( .A(n7573), .B(n7572), .Z(n7574) );
  AND U8068 ( .A(n7575), .B(n7574), .Z(n7832) );
  NANDN U8069 ( .A(n7577), .B(n7576), .Z(n7581) );
  NANDN U8070 ( .A(n7579), .B(n7578), .Z(n7580) );
  AND U8071 ( .A(n7581), .B(n7580), .Z(n7844) );
  NANDN U8072 ( .A(n7583), .B(n7582), .Z(n7587) );
  OR U8073 ( .A(n7585), .B(n7584), .Z(n7586) );
  AND U8074 ( .A(n7587), .B(n7586), .Z(n8072) );
  NANDN U8075 ( .A(n7589), .B(n7588), .Z(n7593) );
  NANDN U8076 ( .A(n7591), .B(n7590), .Z(n7592) );
  AND U8077 ( .A(n7593), .B(n7592), .Z(n8070) );
  NANDN U8078 ( .A(n7595), .B(n7594), .Z(n7599) );
  NAND U8079 ( .A(n7597), .B(n7596), .Z(n7598) );
  AND U8080 ( .A(n7599), .B(n7598), .Z(n7852) );
  NANDN U8081 ( .A(n7601), .B(n7600), .Z(n7605) );
  NANDN U8082 ( .A(n7603), .B(n7602), .Z(n7604) );
  AND U8083 ( .A(n7605), .B(n7604), .Z(n7995) );
  NANDN U8084 ( .A(n7607), .B(n7606), .Z(n7611) );
  NANDN U8085 ( .A(n7609), .B(n7608), .Z(n7610) );
  AND U8086 ( .A(n7611), .B(n7610), .Z(n7993) );
  NAND U8087 ( .A(n33413), .B(n7612), .Z(n7614) );
  XNOR U8088 ( .A(b[21]), .B(a[37]), .Z(n7974) );
  NANDN U8089 ( .A(n7974), .B(n33414), .Z(n7613) );
  NAND U8090 ( .A(n7614), .B(n7613), .Z(n8030) );
  NANDN U8091 ( .A(n33875), .B(n7615), .Z(n7617) );
  XOR U8092 ( .A(b[25]), .B(a[33]), .Z(n7968) );
  NANDN U8093 ( .A(n33994), .B(n7968), .Z(n7616) );
  NAND U8094 ( .A(n7617), .B(n7616), .Z(n8029) );
  XOR U8095 ( .A(n8030), .B(n8029), .Z(n8032) );
  NANDN U8096 ( .A(n32483), .B(n7618), .Z(n7620) );
  XOR U8097 ( .A(b[19]), .B(a[39]), .Z(n7965) );
  NANDN U8098 ( .A(n32823), .B(n7965), .Z(n7619) );
  AND U8099 ( .A(n7620), .B(n7619), .Z(n7908) );
  NANDN U8100 ( .A(n34223), .B(n7621), .Z(n7623) );
  XOR U8101 ( .A(b[27]), .B(a[31]), .Z(n7977) );
  NANDN U8102 ( .A(n34458), .B(n7977), .Z(n7622) );
  AND U8103 ( .A(n7623), .B(n7622), .Z(n7906) );
  NANDN U8104 ( .A(n33866), .B(n7624), .Z(n7626) );
  XOR U8105 ( .A(b[23]), .B(a[35]), .Z(n7971) );
  NANDN U8106 ( .A(n33644), .B(n7971), .Z(n7625) );
  NAND U8107 ( .A(n7626), .B(n7625), .Z(n7905) );
  XNOR U8108 ( .A(n7906), .B(n7905), .Z(n7907) );
  XNOR U8109 ( .A(n7908), .B(n7907), .Z(n8031) );
  XOR U8110 ( .A(n8032), .B(n8031), .Z(n8037) );
  NANDN U8111 ( .A(n7627), .B(n37536), .Z(n7629) );
  XOR U8112 ( .A(b[49]), .B(a[9]), .Z(n7923) );
  NANDN U8113 ( .A(n37432), .B(n7923), .Z(n7628) );
  AND U8114 ( .A(n7629), .B(n7628), .Z(n7931) );
  NANDN U8115 ( .A(n37526), .B(n7630), .Z(n7632) );
  XOR U8116 ( .A(b[51]), .B(a[7]), .Z(n7911) );
  NANDN U8117 ( .A(n37605), .B(n7911), .Z(n7631) );
  AND U8118 ( .A(n7632), .B(n7631), .Z(n7930) );
  NANDN U8119 ( .A(n36742), .B(n7633), .Z(n7635) );
  XOR U8120 ( .A(b[43]), .B(a[15]), .Z(n7887) );
  NANDN U8121 ( .A(n36891), .B(n7887), .Z(n7634) );
  NAND U8122 ( .A(n7635), .B(n7634), .Z(n7929) );
  XOR U8123 ( .A(n7930), .B(n7929), .Z(n7932) );
  XOR U8124 ( .A(n7931), .B(n7932), .Z(n8036) );
  NANDN U8125 ( .A(n31055), .B(n7636), .Z(n7638) );
  XOR U8126 ( .A(b[13]), .B(a[45]), .Z(n7914) );
  NANDN U8127 ( .A(n31293), .B(n7914), .Z(n7637) );
  AND U8128 ( .A(n7638), .B(n7637), .Z(n7877) );
  NANDN U8129 ( .A(n30482), .B(n7639), .Z(n7641) );
  XOR U8130 ( .A(b[11]), .B(a[47]), .Z(n8008) );
  NANDN U8131 ( .A(n30891), .B(n8008), .Z(n7640) );
  AND U8132 ( .A(n7641), .B(n7640), .Z(n7876) );
  NANDN U8133 ( .A(n36210), .B(n7642), .Z(n7644) );
  XOR U8134 ( .A(b[39]), .B(a[19]), .Z(n7962) );
  NANDN U8135 ( .A(n36347), .B(n7962), .Z(n7643) );
  NAND U8136 ( .A(n7644), .B(n7643), .Z(n7875) );
  XOR U8137 ( .A(n7876), .B(n7875), .Z(n7878) );
  XNOR U8138 ( .A(n7877), .B(n7878), .Z(n8035) );
  XOR U8139 ( .A(n8036), .B(n8035), .Z(n8038) );
  XOR U8140 ( .A(n8037), .B(n8038), .Z(n7938) );
  NANDN U8141 ( .A(n7646), .B(n7645), .Z(n7650) );
  NANDN U8142 ( .A(n7648), .B(n7647), .Z(n7649) );
  AND U8143 ( .A(n7650), .B(n7649), .Z(n7936) );
  NANDN U8144 ( .A(n7651), .B(n7766), .Z(n7655) );
  NANDN U8145 ( .A(n7653), .B(n7652), .Z(n7654) );
  NAND U8146 ( .A(n7655), .B(n7654), .Z(n7935) );
  XNOR U8147 ( .A(n7936), .B(n7935), .Z(n7937) );
  XNOR U8148 ( .A(n7938), .B(n7937), .Z(n7992) );
  XNOR U8149 ( .A(n7993), .B(n7992), .Z(n7994) );
  XNOR U8150 ( .A(n7995), .B(n7994), .Z(n7849) );
  NANDN U8151 ( .A(n7657), .B(n7656), .Z(n7661) );
  OR U8152 ( .A(n7659), .B(n7658), .Z(n7660) );
  NAND U8153 ( .A(n7661), .B(n7660), .Z(n7850) );
  XNOR U8154 ( .A(n7849), .B(n7850), .Z(n7851) );
  XNOR U8155 ( .A(n7852), .B(n7851), .Z(n8069) );
  XNOR U8156 ( .A(n8070), .B(n8069), .Z(n8071) );
  XNOR U8157 ( .A(n8072), .B(n8071), .Z(n7843) );
  XNOR U8158 ( .A(n7844), .B(n7843), .Z(n7846) );
  NANDN U8159 ( .A(n7663), .B(n7662), .Z(n7667) );
  OR U8160 ( .A(n7665), .B(n7664), .Z(n7666) );
  AND U8161 ( .A(n7667), .B(n7666), .Z(n7839) );
  NANDN U8162 ( .A(n7669), .B(n7668), .Z(n7673) );
  NANDN U8163 ( .A(n7671), .B(n7670), .Z(n7672) );
  AND U8164 ( .A(n7673), .B(n7672), .Z(n7838) );
  NANDN U8165 ( .A(n7675), .B(n7674), .Z(n7679) );
  NANDN U8166 ( .A(n7677), .B(n7676), .Z(n7678) );
  AND U8167 ( .A(n7679), .B(n7678), .Z(n8064) );
  NAND U8168 ( .A(n7681), .B(n7680), .Z(n7685) );
  NANDN U8169 ( .A(n7683), .B(n7682), .Z(n7684) );
  NAND U8170 ( .A(n7685), .B(n7684), .Z(n8063) );
  XNOR U8171 ( .A(n8064), .B(n8063), .Z(n8066) );
  NANDN U8172 ( .A(n7687), .B(n7686), .Z(n7691) );
  NAND U8173 ( .A(n7689), .B(n7688), .Z(n7690) );
  AND U8174 ( .A(n7691), .B(n7690), .Z(n8065) );
  XOR U8175 ( .A(n8066), .B(n8065), .Z(n8076) );
  NAND U8176 ( .A(n7693), .B(n7692), .Z(n7697) );
  NAND U8177 ( .A(n7695), .B(n7694), .Z(n7696) );
  AND U8178 ( .A(n7697), .B(n7696), .Z(n8075) );
  XNOR U8179 ( .A(n8076), .B(n8075), .Z(n8078) );
  NAND U8180 ( .A(n7699), .B(n7698), .Z(n7703) );
  NAND U8181 ( .A(n7701), .B(n7700), .Z(n7702) );
  AND U8182 ( .A(n7703), .B(n7702), .Z(n8060) );
  NANDN U8183 ( .A(n7705), .B(n7704), .Z(n7709) );
  OR U8184 ( .A(n7707), .B(n7706), .Z(n7708) );
  AND U8185 ( .A(n7709), .B(n7708), .Z(n7948) );
  NANDN U8186 ( .A(n7711), .B(n7710), .Z(n7715) );
  OR U8187 ( .A(n7713), .B(n7712), .Z(n7714) );
  NAND U8188 ( .A(n7715), .B(n7714), .Z(n7947) );
  XNOR U8189 ( .A(n7948), .B(n7947), .Z(n7949) );
  NANDN U8190 ( .A(n7717), .B(n7716), .Z(n7721) );
  OR U8191 ( .A(n7719), .B(n7718), .Z(n7720) );
  AND U8192 ( .A(n7721), .B(n7720), .Z(n7956) );
  NANDN U8193 ( .A(n7722), .B(n37984), .Z(n7724) );
  XOR U8194 ( .A(b[55]), .B(a[3]), .Z(n7858) );
  NANDN U8195 ( .A(n37911), .B(n7858), .Z(n7723) );
  AND U8196 ( .A(n7724), .B(n7723), .Z(n7867) );
  XOR U8197 ( .A(b[57]), .B(b[56]), .Z(n8001) );
  XOR U8198 ( .A(b[57]), .B(a[0]), .Z(n7725) );
  NAND U8199 ( .A(n8001), .B(n7725), .Z(n7726) );
  OR U8200 ( .A(n7726), .B(n38077), .Z(n7728) );
  XOR U8201 ( .A(b[57]), .B(a[1]), .Z(n8002) );
  NAND U8202 ( .A(n38077), .B(n8002), .Z(n7727) );
  AND U8203 ( .A(n7728), .B(n7727), .Z(n7868) );
  XOR U8204 ( .A(n7867), .B(n7868), .Z(n7883) );
  NAND U8205 ( .A(b[0]), .B(a[57]), .Z(n7729) );
  XNOR U8206 ( .A(b[1]), .B(n7729), .Z(n7731) );
  NANDN U8207 ( .A(b[0]), .B(a[56]), .Z(n7730) );
  NAND U8208 ( .A(n7731), .B(n7730), .Z(n7881) );
  NAND U8209 ( .A(n35309), .B(n7732), .Z(n7734) );
  XNOR U8210 ( .A(b[31]), .B(a[27]), .Z(n7864) );
  NANDN U8211 ( .A(n7864), .B(n35310), .Z(n7733) );
  NAND U8212 ( .A(n7734), .B(n7733), .Z(n7882) );
  XOR U8213 ( .A(n7881), .B(n7882), .Z(n7884) );
  XOR U8214 ( .A(n7883), .B(n7884), .Z(n7954) );
  NANDN U8215 ( .A(n35936), .B(n7735), .Z(n7737) );
  XOR U8216 ( .A(b[37]), .B(a[21]), .Z(n8005) );
  NANDN U8217 ( .A(n36047), .B(n8005), .Z(n7736) );
  AND U8218 ( .A(n7737), .B(n7736), .Z(n7872) );
  NANDN U8219 ( .A(n36480), .B(n7738), .Z(n7740) );
  XOR U8220 ( .A(b[41]), .B(a[17]), .Z(n7917) );
  NANDN U8221 ( .A(n36594), .B(n7917), .Z(n7739) );
  AND U8222 ( .A(n7740), .B(n7739), .Z(n7870) );
  NANDN U8223 ( .A(n32013), .B(n7741), .Z(n7743) );
  XOR U8224 ( .A(b[17]), .B(a[41]), .Z(n7893) );
  NANDN U8225 ( .A(n32292), .B(n7893), .Z(n7742) );
  NAND U8226 ( .A(n7743), .B(n7742), .Z(n7869) );
  XNOR U8227 ( .A(n7870), .B(n7869), .Z(n7871) );
  XNOR U8228 ( .A(n7872), .B(n7871), .Z(n7953) );
  XNOR U8229 ( .A(n7954), .B(n7953), .Z(n7955) );
  XOR U8230 ( .A(n7956), .B(n7955), .Z(n7950) );
  XNOR U8231 ( .A(n7949), .B(n7950), .Z(n8059) );
  XNOR U8232 ( .A(n8060), .B(n8059), .Z(n8062) );
  NAND U8233 ( .A(n7745), .B(n7744), .Z(n7749) );
  NAND U8234 ( .A(n7747), .B(n7746), .Z(n7748) );
  NAND U8235 ( .A(n7749), .B(n7748), .Z(n8054) );
  NANDN U8236 ( .A(n210), .B(n7750), .Z(n7752) );
  XOR U8237 ( .A(b[9]), .B(a[49]), .Z(n8011) );
  NANDN U8238 ( .A(n30267), .B(n8011), .Z(n7751) );
  AND U8239 ( .A(n7752), .B(n7751), .Z(n7982) );
  NANDN U8240 ( .A(n29499), .B(n7753), .Z(n7755) );
  XOR U8241 ( .A(b[7]), .B(a[51]), .Z(n7896) );
  NANDN U8242 ( .A(n29735), .B(n7896), .Z(n7754) );
  AND U8243 ( .A(n7755), .B(n7754), .Z(n7981) );
  NANDN U8244 ( .A(n35611), .B(n7756), .Z(n7758) );
  XOR U8245 ( .A(b[35]), .B(a[23]), .Z(n8014) );
  NANDN U8246 ( .A(n35801), .B(n8014), .Z(n7757) );
  NAND U8247 ( .A(n7758), .B(n7757), .Z(n7980) );
  XOR U8248 ( .A(n7981), .B(n7980), .Z(n7983) );
  XOR U8249 ( .A(n7982), .B(n7983), .Z(n7942) );
  NANDN U8250 ( .A(n209), .B(n7759), .Z(n7761) );
  XOR U8251 ( .A(b[3]), .B(a[55]), .Z(n7861) );
  NANDN U8252 ( .A(n28941), .B(n7861), .Z(n7760) );
  AND U8253 ( .A(n7761), .B(n7760), .Z(n7988) );
  NANDN U8254 ( .A(n7762), .B(n35654), .Z(n7764) );
  XOR U8255 ( .A(b[33]), .B(a[25]), .Z(n7902) );
  NANDN U8256 ( .A(n35456), .B(n7902), .Z(n7763) );
  AND U8257 ( .A(n7764), .B(n7763), .Z(n7987) );
  NAND U8258 ( .A(b[55]), .B(b[56]), .Z(n7765) );
  AND U8259 ( .A(b[57]), .B(n7765), .Z(n38167) );
  ANDN U8260 ( .B(n38167), .A(n7766), .Z(n7986) );
  XOR U8261 ( .A(n7987), .B(n7986), .Z(n7989) );
  XNOR U8262 ( .A(n7988), .B(n7989), .Z(n7941) );
  XNOR U8263 ( .A(n7942), .B(n7941), .Z(n7944) );
  NANDN U8264 ( .A(n7768), .B(n7767), .Z(n7772) );
  NANDN U8265 ( .A(n7770), .B(n7769), .Z(n7771) );
  AND U8266 ( .A(n7772), .B(n7771), .Z(n7943) );
  XNOR U8267 ( .A(n7944), .B(n7943), .Z(n8053) );
  XOR U8268 ( .A(n8054), .B(n8053), .Z(n8055) );
  NAND U8269 ( .A(n35001), .B(n7773), .Z(n7775) );
  XNOR U8270 ( .A(b[29]), .B(a[29]), .Z(n7959) );
  NANDN U8271 ( .A(n7959), .B(n35002), .Z(n7774) );
  NAND U8272 ( .A(n7775), .B(n7774), .Z(n8024) );
  NANDN U8273 ( .A(n7776), .B(n29551), .Z(n7778) );
  XOR U8274 ( .A(b[5]), .B(a[53]), .Z(n7899) );
  NANDN U8275 ( .A(n29138), .B(n7899), .Z(n7777) );
  NAND U8276 ( .A(n7778), .B(n7777), .Z(n8023) );
  XOR U8277 ( .A(n8024), .B(n8023), .Z(n8026) );
  NANDN U8278 ( .A(n37705), .B(n7779), .Z(n7781) );
  XOR U8279 ( .A(b[53]), .B(a[5]), .Z(n7998) );
  NANDN U8280 ( .A(n37778), .B(n7998), .Z(n7780) );
  NAND U8281 ( .A(n7781), .B(n7780), .Z(n8025) );
  XOR U8282 ( .A(n8026), .B(n8025), .Z(n8042) );
  NANDN U8283 ( .A(n36991), .B(n7782), .Z(n7784) );
  XOR U8284 ( .A(b[45]), .B(a[13]), .Z(n7890) );
  NANDN U8285 ( .A(n37083), .B(n7890), .Z(n7783) );
  AND U8286 ( .A(n7784), .B(n7783), .Z(n8019) );
  NANDN U8287 ( .A(n211), .B(n7785), .Z(n7787) );
  XOR U8288 ( .A(b[47]), .B(a[11]), .Z(n7920) );
  NANDN U8289 ( .A(n37172), .B(n7920), .Z(n7786) );
  AND U8290 ( .A(n7787), .B(n7786), .Z(n8018) );
  NANDN U8291 ( .A(n31536), .B(n7788), .Z(n7790) );
  XOR U8292 ( .A(b[15]), .B(a[43]), .Z(n7926) );
  NANDN U8293 ( .A(n31925), .B(n7926), .Z(n7789) );
  NAND U8294 ( .A(n7790), .B(n7789), .Z(n8017) );
  XOR U8295 ( .A(n8018), .B(n8017), .Z(n8020) );
  XNOR U8296 ( .A(n8019), .B(n8020), .Z(n8041) );
  XNOR U8297 ( .A(n8042), .B(n8041), .Z(n8043) );
  NANDN U8298 ( .A(n7792), .B(n7791), .Z(n7796) );
  NANDN U8299 ( .A(n7794), .B(n7793), .Z(n7795) );
  NAND U8300 ( .A(n7796), .B(n7795), .Z(n8044) );
  XOR U8301 ( .A(n8043), .B(n8044), .Z(n8049) );
  NANDN U8302 ( .A(n7798), .B(n7797), .Z(n7802) );
  OR U8303 ( .A(n7800), .B(n7799), .Z(n7801) );
  NAND U8304 ( .A(n7802), .B(n7801), .Z(n8047) );
  NAND U8305 ( .A(n7804), .B(n7803), .Z(n7808) );
  NAND U8306 ( .A(n7806), .B(n7805), .Z(n7807) );
  AND U8307 ( .A(n7808), .B(n7807), .Z(n8048) );
  XOR U8308 ( .A(n8047), .B(n8048), .Z(n8050) );
  XNOR U8309 ( .A(n8049), .B(n8050), .Z(n8056) );
  XNOR U8310 ( .A(n8055), .B(n8056), .Z(n8061) );
  XOR U8311 ( .A(n8062), .B(n8061), .Z(n8077) );
  XOR U8312 ( .A(n8078), .B(n8077), .Z(n7837) );
  XOR U8313 ( .A(n7838), .B(n7837), .Z(n7840) );
  XNOR U8314 ( .A(n7839), .B(n7840), .Z(n7845) );
  XOR U8315 ( .A(n7846), .B(n7845), .Z(n8080) );
  NANDN U8316 ( .A(n7810), .B(n7809), .Z(n7814) );
  NANDN U8317 ( .A(n7812), .B(n7811), .Z(n7813) );
  AND U8318 ( .A(n7814), .B(n7813), .Z(n8079) );
  XNOR U8319 ( .A(n8080), .B(n8079), .Z(n8081) );
  NANDN U8320 ( .A(n7816), .B(n7815), .Z(n7820) );
  NAND U8321 ( .A(n7818), .B(n7817), .Z(n7819) );
  NAND U8322 ( .A(n7820), .B(n7819), .Z(n8082) );
  XNOR U8323 ( .A(n8081), .B(n8082), .Z(n7831) );
  XNOR U8324 ( .A(n7832), .B(n7831), .Z(n7833) );
  XNOR U8325 ( .A(n7834), .B(n7833), .Z(n7826) );
  XNOR U8326 ( .A(sreg[121]), .B(n7826), .Z(n7828) );
  NANDN U8327 ( .A(sreg[120]), .B(n7821), .Z(n7825) );
  NAND U8328 ( .A(n7823), .B(n7822), .Z(n7824) );
  NAND U8329 ( .A(n7825), .B(n7824), .Z(n7827) );
  XNOR U8330 ( .A(n7828), .B(n7827), .Z(c[121]) );
  NANDN U8331 ( .A(sreg[121]), .B(n7826), .Z(n7830) );
  NAND U8332 ( .A(n7828), .B(n7827), .Z(n7829) );
  NAND U8333 ( .A(n7830), .B(n7829), .Z(n8352) );
  XNOR U8334 ( .A(sreg[122]), .B(n8352), .Z(n8354) );
  NANDN U8335 ( .A(n7832), .B(n7831), .Z(n7836) );
  NANDN U8336 ( .A(n7834), .B(n7833), .Z(n7835) );
  AND U8337 ( .A(n7836), .B(n7835), .Z(n8088) );
  NANDN U8338 ( .A(n7838), .B(n7837), .Z(n7842) );
  NANDN U8339 ( .A(n7840), .B(n7839), .Z(n7841) );
  AND U8340 ( .A(n7842), .B(n7841), .Z(n8347) );
  NANDN U8341 ( .A(n7844), .B(n7843), .Z(n7848) );
  NAND U8342 ( .A(n7846), .B(n7845), .Z(n7847) );
  NAND U8343 ( .A(n7848), .B(n7847), .Z(n8346) );
  XNOR U8344 ( .A(n8347), .B(n8346), .Z(n8349) );
  NANDN U8345 ( .A(n7850), .B(n7849), .Z(n7854) );
  NANDN U8346 ( .A(n7852), .B(n7851), .Z(n7853) );
  AND U8347 ( .A(n7854), .B(n7853), .Z(n8094) );
  NAND U8348 ( .A(b[0]), .B(a[58]), .Z(n7855) );
  XNOR U8349 ( .A(b[1]), .B(n7855), .Z(n7857) );
  NANDN U8350 ( .A(b[0]), .B(a[57]), .Z(n7856) );
  NAND U8351 ( .A(n7857), .B(n7856), .Z(n8123) );
  XOR U8352 ( .A(b[58]), .B(b[57]), .Z(n38175) );
  IV U8353 ( .A(n38175), .Z(n38130) );
  ANDN U8354 ( .B(a[0]), .A(n38130), .Z(n8141) );
  IV U8355 ( .A(n37984), .Z(n37857) );
  NANDN U8356 ( .A(n37857), .B(n7858), .Z(n7860) );
  XOR U8357 ( .A(b[55]), .B(a[4]), .Z(n8202) );
  NANDN U8358 ( .A(n37911), .B(n8202), .Z(n7859) );
  AND U8359 ( .A(n7860), .B(n7859), .Z(n8121) );
  XOR U8360 ( .A(n8141), .B(n8121), .Z(n8122) );
  XOR U8361 ( .A(n8123), .B(n8122), .Z(n8245) );
  NANDN U8362 ( .A(n209), .B(n7861), .Z(n7863) );
  XOR U8363 ( .A(b[3]), .B(a[56]), .Z(n8265) );
  NANDN U8364 ( .A(n28941), .B(n8265), .Z(n7862) );
  AND U8365 ( .A(n7863), .B(n7862), .Z(n8287) );
  NANDN U8366 ( .A(n7864), .B(n35309), .Z(n7866) );
  XOR U8367 ( .A(b[31]), .B(a[28]), .Z(n8142) );
  NANDN U8368 ( .A(n35145), .B(n8142), .Z(n7865) );
  NAND U8369 ( .A(n7866), .B(n7865), .Z(n8286) );
  XNOR U8370 ( .A(n8287), .B(n8286), .Z(n8289) );
  NOR U8371 ( .A(n7868), .B(n7867), .Z(n8288) );
  XNOR U8372 ( .A(n8289), .B(n8288), .Z(n8244) );
  XNOR U8373 ( .A(n8245), .B(n8244), .Z(n8247) );
  NANDN U8374 ( .A(n7870), .B(n7869), .Z(n7874) );
  NANDN U8375 ( .A(n7872), .B(n7871), .Z(n7873) );
  AND U8376 ( .A(n7874), .B(n7873), .Z(n8246) );
  XOR U8377 ( .A(n8247), .B(n8246), .Z(n8306) );
  NANDN U8378 ( .A(n7876), .B(n7875), .Z(n7880) );
  OR U8379 ( .A(n7878), .B(n7877), .Z(n7879) );
  AND U8380 ( .A(n7880), .B(n7879), .Z(n8305) );
  NANDN U8381 ( .A(n7882), .B(n7881), .Z(n7886) );
  OR U8382 ( .A(n7884), .B(n7883), .Z(n7885) );
  AND U8383 ( .A(n7886), .B(n7885), .Z(n8304) );
  XOR U8384 ( .A(n8305), .B(n8304), .Z(n8307) );
  XOR U8385 ( .A(n8306), .B(n8307), .Z(n8330) );
  NANDN U8386 ( .A(n36742), .B(n7887), .Z(n7889) );
  XOR U8387 ( .A(b[43]), .B(a[16]), .Z(n8226) );
  NANDN U8388 ( .A(n36891), .B(n8226), .Z(n7888) );
  AND U8389 ( .A(n7889), .B(n7888), .Z(n8186) );
  NANDN U8390 ( .A(n36991), .B(n7890), .Z(n7892) );
  XOR U8391 ( .A(b[45]), .B(a[14]), .Z(n8214) );
  NANDN U8392 ( .A(n37083), .B(n8214), .Z(n7891) );
  AND U8393 ( .A(n7892), .B(n7891), .Z(n8185) );
  NANDN U8394 ( .A(n32013), .B(n7893), .Z(n7895) );
  XOR U8395 ( .A(b[17]), .B(a[42]), .Z(n8148) );
  NANDN U8396 ( .A(n32292), .B(n8148), .Z(n7894) );
  NAND U8397 ( .A(n7895), .B(n7894), .Z(n8184) );
  XOR U8398 ( .A(n8185), .B(n8184), .Z(n8187) );
  XOR U8399 ( .A(n8186), .B(n8187), .Z(n8293) );
  NANDN U8400 ( .A(n29499), .B(n7896), .Z(n7898) );
  XOR U8401 ( .A(b[7]), .B(a[52]), .Z(n8166) );
  NANDN U8402 ( .A(n29735), .B(n8166), .Z(n7897) );
  AND U8403 ( .A(n7898), .B(n7897), .Z(n8210) );
  NANDN U8404 ( .A(n28889), .B(n7899), .Z(n7901) );
  XOR U8405 ( .A(b[5]), .B(a[54]), .Z(n8223) );
  NANDN U8406 ( .A(n29138), .B(n8223), .Z(n7900) );
  AND U8407 ( .A(n7901), .B(n7900), .Z(n8209) );
  NANDN U8408 ( .A(n35260), .B(n7902), .Z(n7904) );
  XOR U8409 ( .A(b[33]), .B(a[26]), .Z(n8271) );
  NANDN U8410 ( .A(n35456), .B(n8271), .Z(n7903) );
  NAND U8411 ( .A(n7904), .B(n7903), .Z(n8208) );
  XOR U8412 ( .A(n8209), .B(n8208), .Z(n8211) );
  XNOR U8413 ( .A(n8210), .B(n8211), .Z(n8292) );
  XNOR U8414 ( .A(n8293), .B(n8292), .Z(n8294) );
  NANDN U8415 ( .A(n7906), .B(n7905), .Z(n7910) );
  NANDN U8416 ( .A(n7908), .B(n7907), .Z(n7909) );
  NAND U8417 ( .A(n7910), .B(n7909), .Z(n8295) );
  XNOR U8418 ( .A(n8294), .B(n8295), .Z(n8328) );
  NANDN U8419 ( .A(n37526), .B(n7911), .Z(n7913) );
  XOR U8420 ( .A(b[51]), .B(a[8]), .Z(n8193) );
  NANDN U8421 ( .A(n37605), .B(n8193), .Z(n7912) );
  AND U8422 ( .A(n7913), .B(n7912), .Z(n8180) );
  NANDN U8423 ( .A(n31055), .B(n7914), .Z(n7916) );
  XOR U8424 ( .A(b[13]), .B(a[46]), .Z(n8259) );
  NANDN U8425 ( .A(n31293), .B(n8259), .Z(n7915) );
  AND U8426 ( .A(n7916), .B(n7915), .Z(n8179) );
  NANDN U8427 ( .A(n36480), .B(n7917), .Z(n7919) );
  XOR U8428 ( .A(b[41]), .B(a[18]), .Z(n8163) );
  NANDN U8429 ( .A(n36594), .B(n8163), .Z(n7918) );
  NAND U8430 ( .A(n7919), .B(n7918), .Z(n8178) );
  XOR U8431 ( .A(n8179), .B(n8178), .Z(n8181) );
  XOR U8432 ( .A(n8180), .B(n8181), .Z(n8311) );
  NANDN U8433 ( .A(n211), .B(n7920), .Z(n7922) );
  XOR U8434 ( .A(b[47]), .B(a[12]), .Z(n8217) );
  NANDN U8435 ( .A(n37172), .B(n8217), .Z(n7921) );
  AND U8436 ( .A(n7922), .B(n7921), .Z(n8234) );
  NANDN U8437 ( .A(n212), .B(n7923), .Z(n7925) );
  XOR U8438 ( .A(b[49]), .B(a[10]), .Z(n8268) );
  NANDN U8439 ( .A(n37432), .B(n8268), .Z(n7924) );
  AND U8440 ( .A(n7925), .B(n7924), .Z(n8233) );
  NANDN U8441 ( .A(n31536), .B(n7926), .Z(n7928) );
  XOR U8442 ( .A(b[15]), .B(a[44]), .Z(n8151) );
  NANDN U8443 ( .A(n31925), .B(n8151), .Z(n7927) );
  NAND U8444 ( .A(n7928), .B(n7927), .Z(n8232) );
  XOR U8445 ( .A(n8233), .B(n8232), .Z(n8235) );
  XNOR U8446 ( .A(n8234), .B(n8235), .Z(n8310) );
  XNOR U8447 ( .A(n8311), .B(n8310), .Z(n8312) );
  NANDN U8448 ( .A(n7930), .B(n7929), .Z(n7934) );
  OR U8449 ( .A(n7932), .B(n7931), .Z(n7933) );
  NAND U8450 ( .A(n7934), .B(n7933), .Z(n8313) );
  XOR U8451 ( .A(n8312), .B(n8313), .Z(n8329) );
  XOR U8452 ( .A(n8328), .B(n8329), .Z(n8331) );
  XOR U8453 ( .A(n8330), .B(n8331), .Z(n8252) );
  NANDN U8454 ( .A(n7936), .B(n7935), .Z(n7940) );
  NANDN U8455 ( .A(n7938), .B(n7937), .Z(n7939) );
  AND U8456 ( .A(n7940), .B(n7939), .Z(n8251) );
  NANDN U8457 ( .A(n7942), .B(n7941), .Z(n7946) );
  NAND U8458 ( .A(n7944), .B(n7943), .Z(n7945) );
  AND U8459 ( .A(n7946), .B(n7945), .Z(n8250) );
  XOR U8460 ( .A(n8251), .B(n8250), .Z(n8253) );
  XOR U8461 ( .A(n8252), .B(n8253), .Z(n8099) );
  NANDN U8462 ( .A(n7948), .B(n7947), .Z(n7952) );
  NANDN U8463 ( .A(n7950), .B(n7949), .Z(n7951) );
  AND U8464 ( .A(n7952), .B(n7951), .Z(n8318) );
  NANDN U8465 ( .A(n7954), .B(n7953), .Z(n7958) );
  NANDN U8466 ( .A(n7956), .B(n7955), .Z(n7957) );
  AND U8467 ( .A(n7958), .B(n7957), .Z(n8317) );
  NANDN U8468 ( .A(n7959), .B(n35001), .Z(n7961) );
  XOR U8469 ( .A(b[29]), .B(a[30]), .Z(n8205) );
  NANDN U8470 ( .A(n34722), .B(n8205), .Z(n7960) );
  AND U8471 ( .A(n7961), .B(n7960), .Z(n8128) );
  NANDN U8472 ( .A(n36210), .B(n7962), .Z(n7964) );
  XOR U8473 ( .A(b[39]), .B(a[20]), .Z(n8160) );
  NANDN U8474 ( .A(n36347), .B(n8160), .Z(n7963) );
  AND U8475 ( .A(n7964), .B(n7963), .Z(n8127) );
  NANDN U8476 ( .A(n32483), .B(n7965), .Z(n7967) );
  XOR U8477 ( .A(b[19]), .B(a[40]), .Z(n8145) );
  NANDN U8478 ( .A(n32823), .B(n8145), .Z(n7966) );
  NAND U8479 ( .A(n7967), .B(n7966), .Z(n8126) );
  XOR U8480 ( .A(n8127), .B(n8126), .Z(n8129) );
  XOR U8481 ( .A(n8128), .B(n8129), .Z(n8156) );
  NANDN U8482 ( .A(n33875), .B(n7968), .Z(n7970) );
  XOR U8483 ( .A(b[25]), .B(a[34]), .Z(n8220) );
  NANDN U8484 ( .A(n33994), .B(n8220), .Z(n7969) );
  AND U8485 ( .A(n7970), .B(n7969), .Z(n8276) );
  NANDN U8486 ( .A(n33866), .B(n7971), .Z(n7973) );
  XOR U8487 ( .A(b[23]), .B(a[36]), .Z(n8169) );
  NANDN U8488 ( .A(n33644), .B(n8169), .Z(n7972) );
  AND U8489 ( .A(n7973), .B(n7972), .Z(n8275) );
  NANDN U8490 ( .A(n7974), .B(n33413), .Z(n7976) );
  XOR U8491 ( .A(b[21]), .B(a[38]), .Z(n8256) );
  NANDN U8492 ( .A(n33271), .B(n8256), .Z(n7975) );
  NAND U8493 ( .A(n7976), .B(n7975), .Z(n8274) );
  XOR U8494 ( .A(n8275), .B(n8274), .Z(n8277) );
  XOR U8495 ( .A(n8276), .B(n8277), .Z(n8155) );
  NAND U8496 ( .A(n34647), .B(n7977), .Z(n7979) );
  XNOR U8497 ( .A(b[27]), .B(a[32]), .Z(n8196) );
  NANDN U8498 ( .A(n8196), .B(n34648), .Z(n7978) );
  AND U8499 ( .A(n7979), .B(n7978), .Z(n8154) );
  XOR U8500 ( .A(n8155), .B(n8154), .Z(n8157) );
  XOR U8501 ( .A(n8156), .B(n8157), .Z(n8301) );
  NANDN U8502 ( .A(n7981), .B(n7980), .Z(n7985) );
  OR U8503 ( .A(n7983), .B(n7982), .Z(n7984) );
  AND U8504 ( .A(n7985), .B(n7984), .Z(n8299) );
  NANDN U8505 ( .A(n7987), .B(n7986), .Z(n7991) );
  OR U8506 ( .A(n7989), .B(n7988), .Z(n7990) );
  NAND U8507 ( .A(n7991), .B(n7990), .Z(n8298) );
  XNOR U8508 ( .A(n8299), .B(n8298), .Z(n8300) );
  XNOR U8509 ( .A(n8301), .B(n8300), .Z(n8316) );
  XOR U8510 ( .A(n8317), .B(n8316), .Z(n8319) );
  XOR U8511 ( .A(n8318), .B(n8319), .Z(n8098) );
  NANDN U8512 ( .A(n7993), .B(n7992), .Z(n7997) );
  NANDN U8513 ( .A(n7995), .B(n7994), .Z(n7996) );
  AND U8514 ( .A(n7997), .B(n7996), .Z(n8097) );
  XOR U8515 ( .A(n8098), .B(n8097), .Z(n8100) );
  XOR U8516 ( .A(n8099), .B(n8100), .Z(n8092) );
  NANDN U8517 ( .A(n37705), .B(n7998), .Z(n8000) );
  XOR U8518 ( .A(b[53]), .B(a[6]), .Z(n8199) );
  NANDN U8519 ( .A(n37778), .B(n8199), .Z(n7999) );
  AND U8520 ( .A(n8000), .B(n7999), .Z(n8282) );
  ANDN U8521 ( .B(n8001), .A(n38077), .Z(n38076) );
  IV U8522 ( .A(n38076), .Z(n37974) );
  NANDN U8523 ( .A(n37974), .B(n8002), .Z(n8004) );
  XOR U8524 ( .A(b[57]), .B(a[2]), .Z(n8137) );
  NANDN U8525 ( .A(n38031), .B(n8137), .Z(n8003) );
  AND U8526 ( .A(n8004), .B(n8003), .Z(n8281) );
  NANDN U8527 ( .A(n35936), .B(n8005), .Z(n8007) );
  XOR U8528 ( .A(b[37]), .B(a[22]), .Z(n8172) );
  NANDN U8529 ( .A(n36047), .B(n8172), .Z(n8006) );
  NAND U8530 ( .A(n8007), .B(n8006), .Z(n8280) );
  XOR U8531 ( .A(n8281), .B(n8280), .Z(n8283) );
  XOR U8532 ( .A(n8282), .B(n8283), .Z(n8239) );
  NANDN U8533 ( .A(n30482), .B(n8008), .Z(n8010) );
  XOR U8534 ( .A(b[11]), .B(a[48]), .Z(n8262) );
  NANDN U8535 ( .A(n30891), .B(n8262), .Z(n8009) );
  AND U8536 ( .A(n8010), .B(n8009), .Z(n8117) );
  NANDN U8537 ( .A(n210), .B(n8011), .Z(n8013) );
  XOR U8538 ( .A(b[9]), .B(a[50]), .Z(n8175) );
  NANDN U8539 ( .A(n30267), .B(n8175), .Z(n8012) );
  AND U8540 ( .A(n8013), .B(n8012), .Z(n8116) );
  NANDN U8541 ( .A(n35611), .B(n8014), .Z(n8016) );
  XOR U8542 ( .A(b[35]), .B(a[24]), .Z(n8229) );
  NANDN U8543 ( .A(n35801), .B(n8229), .Z(n8015) );
  NAND U8544 ( .A(n8016), .B(n8015), .Z(n8115) );
  XOR U8545 ( .A(n8116), .B(n8115), .Z(n8118) );
  XNOR U8546 ( .A(n8117), .B(n8118), .Z(n8238) );
  XNOR U8547 ( .A(n8239), .B(n8238), .Z(n8240) );
  NANDN U8548 ( .A(n8018), .B(n8017), .Z(n8022) );
  OR U8549 ( .A(n8020), .B(n8019), .Z(n8021) );
  NAND U8550 ( .A(n8022), .B(n8021), .Z(n8241) );
  XOR U8551 ( .A(n8240), .B(n8241), .Z(n8323) );
  NAND U8552 ( .A(n8024), .B(n8023), .Z(n8028) );
  NAND U8553 ( .A(n8026), .B(n8025), .Z(n8027) );
  NAND U8554 ( .A(n8028), .B(n8027), .Z(n8322) );
  XOR U8555 ( .A(n8323), .B(n8322), .Z(n8325) );
  NAND U8556 ( .A(n8030), .B(n8029), .Z(n8034) );
  NAND U8557 ( .A(n8032), .B(n8031), .Z(n8033) );
  NAND U8558 ( .A(n8034), .B(n8033), .Z(n8324) );
  XOR U8559 ( .A(n8325), .B(n8324), .Z(n8112) );
  NANDN U8560 ( .A(n8036), .B(n8035), .Z(n8040) );
  OR U8561 ( .A(n8038), .B(n8037), .Z(n8039) );
  AND U8562 ( .A(n8040), .B(n8039), .Z(n8110) );
  NANDN U8563 ( .A(n8042), .B(n8041), .Z(n8046) );
  NANDN U8564 ( .A(n8044), .B(n8043), .Z(n8045) );
  NAND U8565 ( .A(n8046), .B(n8045), .Z(n8109) );
  XNOR U8566 ( .A(n8110), .B(n8109), .Z(n8111) );
  XNOR U8567 ( .A(n8112), .B(n8111), .Z(n8104) );
  NAND U8568 ( .A(n8048), .B(n8047), .Z(n8052) );
  NAND U8569 ( .A(n8050), .B(n8049), .Z(n8051) );
  AND U8570 ( .A(n8052), .B(n8051), .Z(n8103) );
  XOR U8571 ( .A(n8104), .B(n8103), .Z(n8106) );
  NAND U8572 ( .A(n8054), .B(n8053), .Z(n8058) );
  NANDN U8573 ( .A(n8056), .B(n8055), .Z(n8057) );
  AND U8574 ( .A(n8058), .B(n8057), .Z(n8105) );
  XOR U8575 ( .A(n8106), .B(n8105), .Z(n8337) );
  NANDN U8576 ( .A(n8064), .B(n8063), .Z(n8068) );
  NAND U8577 ( .A(n8066), .B(n8065), .Z(n8067) );
  AND U8578 ( .A(n8068), .B(n8067), .Z(n8334) );
  XNOR U8579 ( .A(n8335), .B(n8334), .Z(n8336) );
  XNOR U8580 ( .A(n8337), .B(n8336), .Z(n8091) );
  XNOR U8581 ( .A(n8092), .B(n8091), .Z(n8093) );
  XNOR U8582 ( .A(n8094), .B(n8093), .Z(n8342) );
  NANDN U8583 ( .A(n8070), .B(n8069), .Z(n8074) );
  NANDN U8584 ( .A(n8072), .B(n8071), .Z(n8073) );
  AND U8585 ( .A(n8074), .B(n8073), .Z(n8341) );
  XOR U8586 ( .A(n8341), .B(n8340), .Z(n8343) );
  XNOR U8587 ( .A(n8342), .B(n8343), .Z(n8348) );
  XOR U8588 ( .A(n8349), .B(n8348), .Z(n8086) );
  NANDN U8589 ( .A(n8080), .B(n8079), .Z(n8084) );
  NANDN U8590 ( .A(n8082), .B(n8081), .Z(n8083) );
  NAND U8591 ( .A(n8084), .B(n8083), .Z(n8085) );
  XNOR U8592 ( .A(n8086), .B(n8085), .Z(n8087) );
  XNOR U8593 ( .A(n8088), .B(n8087), .Z(n8353) );
  XNOR U8594 ( .A(n8354), .B(n8353), .Z(c[122]) );
  NANDN U8595 ( .A(n8086), .B(n8085), .Z(n8090) );
  NANDN U8596 ( .A(n8088), .B(n8087), .Z(n8089) );
  AND U8597 ( .A(n8090), .B(n8089), .Z(n8365) );
  NANDN U8598 ( .A(n8092), .B(n8091), .Z(n8096) );
  NANDN U8599 ( .A(n8094), .B(n8093), .Z(n8095) );
  AND U8600 ( .A(n8096), .B(n8095), .Z(n8623) );
  NANDN U8601 ( .A(n8098), .B(n8097), .Z(n8102) );
  OR U8602 ( .A(n8100), .B(n8099), .Z(n8101) );
  AND U8603 ( .A(n8102), .B(n8101), .Z(n8614) );
  NAND U8604 ( .A(n8104), .B(n8103), .Z(n8108) );
  NAND U8605 ( .A(n8106), .B(n8105), .Z(n8107) );
  AND U8606 ( .A(n8108), .B(n8107), .Z(n8612) );
  NANDN U8607 ( .A(n8110), .B(n8109), .Z(n8114) );
  NANDN U8608 ( .A(n8112), .B(n8111), .Z(n8113) );
  AND U8609 ( .A(n8114), .B(n8113), .Z(n8371) );
  NANDN U8610 ( .A(n8116), .B(n8115), .Z(n8120) );
  OR U8611 ( .A(n8118), .B(n8117), .Z(n8119) );
  AND U8612 ( .A(n8120), .B(n8119), .Z(n8546) );
  NANDN U8613 ( .A(n8121), .B(n8141), .Z(n8125) );
  OR U8614 ( .A(n8123), .B(n8122), .Z(n8124) );
  NAND U8615 ( .A(n8125), .B(n8124), .Z(n8545) );
  XNOR U8616 ( .A(n8546), .B(n8545), .Z(n8548) );
  NANDN U8617 ( .A(n8127), .B(n8126), .Z(n8131) );
  OR U8618 ( .A(n8129), .B(n8128), .Z(n8130) );
  AND U8619 ( .A(n8131), .B(n8130), .Z(n8419) );
  XOR U8620 ( .A(b[59]), .B(a[0]), .Z(n8134) );
  XOR U8621 ( .A(b[59]), .B(b[57]), .Z(n8132) );
  XOR U8622 ( .A(b[59]), .B(b[58]), .Z(n8577) );
  AND U8623 ( .A(n8132), .B(n8577), .Z(n8133) );
  NAND U8624 ( .A(n8134), .B(n8133), .Z(n8136) );
  XOR U8625 ( .A(b[59]), .B(a[1]), .Z(n8578) );
  NANDN U8626 ( .A(n38130), .B(n8578), .Z(n8135) );
  AND U8627 ( .A(n8136), .B(n8135), .Z(n8576) );
  NANDN U8628 ( .A(n37974), .B(n8137), .Z(n8139) );
  XOR U8629 ( .A(b[57]), .B(a[3]), .Z(n8491) );
  NANDN U8630 ( .A(n38031), .B(n8491), .Z(n8138) );
  AND U8631 ( .A(n8139), .B(n8138), .Z(n8575) );
  XOR U8632 ( .A(n8576), .B(n8575), .Z(n8403) );
  NAND U8633 ( .A(b[57]), .B(b[58]), .Z(n8140) );
  NAND U8634 ( .A(b[59]), .B(n8140), .Z(n38210) );
  NOR U8635 ( .A(n38210), .B(n8141), .Z(n8402) );
  NAND U8636 ( .A(n35309), .B(n8142), .Z(n8144) );
  XNOR U8637 ( .A(b[31]), .B(a[29]), .Z(n8413) );
  NANDN U8638 ( .A(n8413), .B(n35310), .Z(n8143) );
  AND U8639 ( .A(n8144), .B(n8143), .Z(n8401) );
  XOR U8640 ( .A(n8402), .B(n8401), .Z(n8404) );
  XOR U8641 ( .A(n8403), .B(n8404), .Z(n8417) );
  NANDN U8642 ( .A(n32483), .B(n8145), .Z(n8147) );
  XOR U8643 ( .A(b[19]), .B(a[41]), .Z(n8389) );
  NANDN U8644 ( .A(n32823), .B(n8389), .Z(n8146) );
  AND U8645 ( .A(n8147), .B(n8146), .Z(n8524) );
  NANDN U8646 ( .A(n32013), .B(n8148), .Z(n8150) );
  XOR U8647 ( .A(b[17]), .B(a[43]), .Z(n8500) );
  NANDN U8648 ( .A(n32292), .B(n8500), .Z(n8149) );
  AND U8649 ( .A(n8150), .B(n8149), .Z(n8522) );
  NANDN U8650 ( .A(n31536), .B(n8151), .Z(n8153) );
  XOR U8651 ( .A(b[15]), .B(a[45]), .Z(n8509) );
  NANDN U8652 ( .A(n31925), .B(n8509), .Z(n8152) );
  NAND U8653 ( .A(n8153), .B(n8152), .Z(n8521) );
  XNOR U8654 ( .A(n8522), .B(n8521), .Z(n8523) );
  XNOR U8655 ( .A(n8524), .B(n8523), .Z(n8416) );
  XNOR U8656 ( .A(n8417), .B(n8416), .Z(n8418) );
  XNOR U8657 ( .A(n8419), .B(n8418), .Z(n8547) );
  XOR U8658 ( .A(n8548), .B(n8547), .Z(n8376) );
  NANDN U8659 ( .A(n8155), .B(n8154), .Z(n8159) );
  OR U8660 ( .A(n8157), .B(n8156), .Z(n8158) );
  AND U8661 ( .A(n8159), .B(n8158), .Z(n8375) );
  NANDN U8662 ( .A(n36210), .B(n8160), .Z(n8162) );
  XOR U8663 ( .A(b[39]), .B(a[21]), .Z(n8455) );
  NANDN U8664 ( .A(n36347), .B(n8455), .Z(n8161) );
  AND U8665 ( .A(n8162), .B(n8161), .Z(n8460) );
  NANDN U8666 ( .A(n36480), .B(n8163), .Z(n8165) );
  XOR U8667 ( .A(b[41]), .B(a[19]), .Z(n8497) );
  NANDN U8668 ( .A(n36594), .B(n8497), .Z(n8164) );
  AND U8669 ( .A(n8165), .B(n8164), .Z(n8459) );
  NANDN U8670 ( .A(n29499), .B(n8166), .Z(n8168) );
  XOR U8671 ( .A(b[7]), .B(a[53]), .Z(n8443) );
  NANDN U8672 ( .A(n29735), .B(n8443), .Z(n8167) );
  NAND U8673 ( .A(n8168), .B(n8167), .Z(n8458) );
  XOR U8674 ( .A(n8459), .B(n8458), .Z(n8461) );
  XOR U8675 ( .A(n8460), .B(n8461), .Z(n8540) );
  NANDN U8676 ( .A(n33866), .B(n8169), .Z(n8171) );
  XOR U8677 ( .A(b[23]), .B(a[37]), .Z(n8398) );
  NANDN U8678 ( .A(n33644), .B(n8398), .Z(n8170) );
  AND U8679 ( .A(n8171), .B(n8170), .Z(n8484) );
  NANDN U8680 ( .A(n35936), .B(n8172), .Z(n8174) );
  XOR U8681 ( .A(b[37]), .B(a[23]), .Z(n8446) );
  NANDN U8682 ( .A(n36047), .B(n8446), .Z(n8173) );
  AND U8683 ( .A(n8174), .B(n8173), .Z(n8483) );
  NANDN U8684 ( .A(n210), .B(n8175), .Z(n8177) );
  XOR U8685 ( .A(b[9]), .B(a[51]), .Z(n8440) );
  NANDN U8686 ( .A(n30267), .B(n8440), .Z(n8176) );
  NAND U8687 ( .A(n8177), .B(n8176), .Z(n8482) );
  XOR U8688 ( .A(n8483), .B(n8482), .Z(n8485) );
  XNOR U8689 ( .A(n8484), .B(n8485), .Z(n8539) );
  XNOR U8690 ( .A(n8540), .B(n8539), .Z(n8541) );
  NANDN U8691 ( .A(n8179), .B(n8178), .Z(n8183) );
  OR U8692 ( .A(n8181), .B(n8180), .Z(n8182) );
  NAND U8693 ( .A(n8183), .B(n8182), .Z(n8542) );
  XNOR U8694 ( .A(n8541), .B(n8542), .Z(n8374) );
  XOR U8695 ( .A(n8375), .B(n8374), .Z(n8377) );
  XOR U8696 ( .A(n8376), .B(n8377), .Z(n8369) );
  NANDN U8697 ( .A(n8185), .B(n8184), .Z(n8189) );
  OR U8698 ( .A(n8187), .B(n8186), .Z(n8188) );
  AND U8699 ( .A(n8189), .B(n8188), .Z(n8535) );
  NAND U8700 ( .A(b[0]), .B(a[59]), .Z(n8190) );
  XNOR U8701 ( .A(b[1]), .B(n8190), .Z(n8192) );
  NANDN U8702 ( .A(b[0]), .B(a[58]), .Z(n8191) );
  NAND U8703 ( .A(n8192), .B(n8191), .Z(n8566) );
  NANDN U8704 ( .A(n37526), .B(n8193), .Z(n8195) );
  XOR U8705 ( .A(b[51]), .B(a[9]), .Z(n8590) );
  NANDN U8706 ( .A(n37605), .B(n8590), .Z(n8194) );
  AND U8707 ( .A(n8195), .B(n8194), .Z(n8564) );
  NANDN U8708 ( .A(n8196), .B(n34647), .Z(n8198) );
  XOR U8709 ( .A(b[27]), .B(a[33]), .Z(n8395) );
  NANDN U8710 ( .A(n34458), .B(n8395), .Z(n8197) );
  NAND U8711 ( .A(n8198), .B(n8197), .Z(n8563) );
  XNOR U8712 ( .A(n8564), .B(n8563), .Z(n8565) );
  XNOR U8713 ( .A(n8566), .B(n8565), .Z(n8533) );
  NANDN U8714 ( .A(n37705), .B(n8199), .Z(n8201) );
  XOR U8715 ( .A(b[53]), .B(a[7]), .Z(n8512) );
  NANDN U8716 ( .A(n37778), .B(n8512), .Z(n8200) );
  AND U8717 ( .A(n8201), .B(n8200), .Z(n8473) );
  NANDN U8718 ( .A(n37857), .B(n8202), .Z(n8204) );
  XOR U8719 ( .A(b[55]), .B(a[5]), .Z(n8410) );
  NANDN U8720 ( .A(n37911), .B(n8410), .Z(n8203) );
  AND U8721 ( .A(n8204), .B(n8203), .Z(n8471) );
  NANDN U8722 ( .A(n34634), .B(n8205), .Z(n8207) );
  XOR U8723 ( .A(b[29]), .B(a[31]), .Z(n8494) );
  NANDN U8724 ( .A(n34722), .B(n8494), .Z(n8206) );
  NAND U8725 ( .A(n8207), .B(n8206), .Z(n8470) );
  XNOR U8726 ( .A(n8471), .B(n8470), .Z(n8472) );
  XOR U8727 ( .A(n8473), .B(n8472), .Z(n8534) );
  XOR U8728 ( .A(n8533), .B(n8534), .Z(n8536) );
  XOR U8729 ( .A(n8535), .B(n8536), .Z(n8594) );
  NANDN U8730 ( .A(n8209), .B(n8208), .Z(n8213) );
  OR U8731 ( .A(n8211), .B(n8210), .Z(n8212) );
  AND U8732 ( .A(n8213), .B(n8212), .Z(n8593) );
  XNOR U8733 ( .A(n8594), .B(n8593), .Z(n8595) );
  NANDN U8734 ( .A(n36991), .B(n8214), .Z(n8216) );
  XOR U8735 ( .A(b[45]), .B(a[15]), .Z(n8506) );
  NANDN U8736 ( .A(n37083), .B(n8506), .Z(n8215) );
  AND U8737 ( .A(n8216), .B(n8215), .Z(n8559) );
  NANDN U8738 ( .A(n211), .B(n8217), .Z(n8219) );
  XOR U8739 ( .A(b[47]), .B(a[13]), .Z(n8584) );
  NANDN U8740 ( .A(n37172), .B(n8584), .Z(n8218) );
  AND U8741 ( .A(n8219), .B(n8218), .Z(n8558) );
  NANDN U8742 ( .A(n33875), .B(n8220), .Z(n8222) );
  XOR U8743 ( .A(b[25]), .B(a[35]), .Z(n8392) );
  NANDN U8744 ( .A(n33994), .B(n8392), .Z(n8221) );
  NAND U8745 ( .A(n8222), .B(n8221), .Z(n8557) );
  XOR U8746 ( .A(n8558), .B(n8557), .Z(n8560) );
  XOR U8747 ( .A(n8559), .B(n8560), .Z(n8477) );
  NANDN U8748 ( .A(n28889), .B(n8223), .Z(n8225) );
  XOR U8749 ( .A(b[5]), .B(a[55]), .Z(n8515) );
  NANDN U8750 ( .A(n29138), .B(n8515), .Z(n8224) );
  AND U8751 ( .A(n8225), .B(n8224), .Z(n8571) );
  NANDN U8752 ( .A(n36742), .B(n8226), .Z(n8228) );
  XOR U8753 ( .A(b[43]), .B(a[17]), .Z(n8503) );
  NANDN U8754 ( .A(n36891), .B(n8503), .Z(n8227) );
  AND U8755 ( .A(n8228), .B(n8227), .Z(n8570) );
  NANDN U8756 ( .A(n35611), .B(n8229), .Z(n8231) );
  XOR U8757 ( .A(b[35]), .B(a[25]), .Z(n8518) );
  NANDN U8758 ( .A(n35801), .B(n8518), .Z(n8230) );
  NAND U8759 ( .A(n8231), .B(n8230), .Z(n8569) );
  XOR U8760 ( .A(n8570), .B(n8569), .Z(n8572) );
  XNOR U8761 ( .A(n8571), .B(n8572), .Z(n8476) );
  XNOR U8762 ( .A(n8477), .B(n8476), .Z(n8478) );
  NANDN U8763 ( .A(n8233), .B(n8232), .Z(n8237) );
  OR U8764 ( .A(n8235), .B(n8234), .Z(n8236) );
  NAND U8765 ( .A(n8237), .B(n8236), .Z(n8479) );
  XOR U8766 ( .A(n8478), .B(n8479), .Z(n8596) );
  XNOR U8767 ( .A(n8595), .B(n8596), .Z(n8383) );
  NANDN U8768 ( .A(n8239), .B(n8238), .Z(n8243) );
  NANDN U8769 ( .A(n8241), .B(n8240), .Z(n8242) );
  AND U8770 ( .A(n8243), .B(n8242), .Z(n8381) );
  NANDN U8771 ( .A(n8245), .B(n8244), .Z(n8249) );
  NAND U8772 ( .A(n8247), .B(n8246), .Z(n8248) );
  NAND U8773 ( .A(n8249), .B(n8248), .Z(n8380) );
  XNOR U8774 ( .A(n8381), .B(n8380), .Z(n8382) );
  XNOR U8775 ( .A(n8383), .B(n8382), .Z(n8368) );
  XNOR U8776 ( .A(n8369), .B(n8368), .Z(n8370) );
  XOR U8777 ( .A(n8371), .B(n8370), .Z(n8611) );
  XOR U8778 ( .A(n8612), .B(n8611), .Z(n8613) );
  XOR U8779 ( .A(n8614), .B(n8613), .Z(n8620) );
  NANDN U8780 ( .A(n8251), .B(n8250), .Z(n8255) );
  OR U8781 ( .A(n8253), .B(n8252), .Z(n8254) );
  AND U8782 ( .A(n8255), .B(n8254), .Z(n8607) );
  NANDN U8783 ( .A(n32996), .B(n8256), .Z(n8258) );
  XOR U8784 ( .A(b[21]), .B(a[39]), .Z(n8386) );
  NANDN U8785 ( .A(n33271), .B(n8386), .Z(n8257) );
  AND U8786 ( .A(n8258), .B(n8257), .Z(n8467) );
  NANDN U8787 ( .A(n31055), .B(n8259), .Z(n8261) );
  XOR U8788 ( .A(b[13]), .B(a[47]), .Z(n8449) );
  NANDN U8789 ( .A(n31293), .B(n8449), .Z(n8260) );
  AND U8790 ( .A(n8261), .B(n8260), .Z(n8465) );
  NANDN U8791 ( .A(n30482), .B(n8262), .Z(n8264) );
  XOR U8792 ( .A(b[11]), .B(a[49]), .Z(n8452) );
  NANDN U8793 ( .A(n30891), .B(n8452), .Z(n8263) );
  NAND U8794 ( .A(n8264), .B(n8263), .Z(n8464) );
  XNOR U8795 ( .A(n8465), .B(n8464), .Z(n8466) );
  XOR U8796 ( .A(n8467), .B(n8466), .Z(n8552) );
  NANDN U8797 ( .A(n209), .B(n8265), .Z(n8267) );
  XOR U8798 ( .A(b[3]), .B(a[57]), .Z(n8407) );
  NANDN U8799 ( .A(n28941), .B(n8407), .Z(n8266) );
  AND U8800 ( .A(n8267), .B(n8266), .Z(n8529) );
  NANDN U8801 ( .A(n212), .B(n8268), .Z(n8270) );
  XOR U8802 ( .A(b[49]), .B(a[11]), .Z(n8587) );
  NANDN U8803 ( .A(n37432), .B(n8587), .Z(n8269) );
  AND U8804 ( .A(n8270), .B(n8269), .Z(n8528) );
  NANDN U8805 ( .A(n35260), .B(n8271), .Z(n8273) );
  XOR U8806 ( .A(b[33]), .B(a[27]), .Z(n8581) );
  NANDN U8807 ( .A(n35456), .B(n8581), .Z(n8272) );
  NAND U8808 ( .A(n8273), .B(n8272), .Z(n8527) );
  XOR U8809 ( .A(n8528), .B(n8527), .Z(n8530) );
  XNOR U8810 ( .A(n8529), .B(n8530), .Z(n8551) );
  XOR U8811 ( .A(n8552), .B(n8551), .Z(n8554) );
  NANDN U8812 ( .A(n8275), .B(n8274), .Z(n8279) );
  OR U8813 ( .A(n8277), .B(n8276), .Z(n8278) );
  AND U8814 ( .A(n8279), .B(n8278), .Z(n8553) );
  XOR U8815 ( .A(n8554), .B(n8553), .Z(n8424) );
  NANDN U8816 ( .A(n8281), .B(n8280), .Z(n8285) );
  OR U8817 ( .A(n8283), .B(n8282), .Z(n8284) );
  AND U8818 ( .A(n8285), .B(n8284), .Z(n8423) );
  NANDN U8819 ( .A(n8287), .B(n8286), .Z(n8291) );
  NAND U8820 ( .A(n8289), .B(n8288), .Z(n8290) );
  NAND U8821 ( .A(n8291), .B(n8290), .Z(n8422) );
  XOR U8822 ( .A(n8423), .B(n8422), .Z(n8425) );
  XOR U8823 ( .A(n8424), .B(n8425), .Z(n8435) );
  NANDN U8824 ( .A(n8293), .B(n8292), .Z(n8297) );
  NANDN U8825 ( .A(n8295), .B(n8294), .Z(n8296) );
  NAND U8826 ( .A(n8297), .B(n8296), .Z(n8434) );
  XNOR U8827 ( .A(n8435), .B(n8434), .Z(n8437) );
  NANDN U8828 ( .A(n8299), .B(n8298), .Z(n8303) );
  NANDN U8829 ( .A(n8301), .B(n8300), .Z(n8302) );
  AND U8830 ( .A(n8303), .B(n8302), .Z(n8436) );
  XOR U8831 ( .A(n8437), .B(n8436), .Z(n8431) );
  NANDN U8832 ( .A(n8305), .B(n8304), .Z(n8309) );
  OR U8833 ( .A(n8307), .B(n8306), .Z(n8308) );
  AND U8834 ( .A(n8309), .B(n8308), .Z(n8429) );
  NANDN U8835 ( .A(n8311), .B(n8310), .Z(n8315) );
  NANDN U8836 ( .A(n8313), .B(n8312), .Z(n8314) );
  AND U8837 ( .A(n8315), .B(n8314), .Z(n8428) );
  XNOR U8838 ( .A(n8429), .B(n8428), .Z(n8430) );
  XNOR U8839 ( .A(n8431), .B(n8430), .Z(n8605) );
  NANDN U8840 ( .A(n8317), .B(n8316), .Z(n8321) );
  OR U8841 ( .A(n8319), .B(n8318), .Z(n8320) );
  AND U8842 ( .A(n8321), .B(n8320), .Z(n8602) );
  NAND U8843 ( .A(n8323), .B(n8322), .Z(n8327) );
  NAND U8844 ( .A(n8325), .B(n8324), .Z(n8326) );
  AND U8845 ( .A(n8327), .B(n8326), .Z(n8600) );
  NANDN U8846 ( .A(n8329), .B(n8328), .Z(n8333) );
  OR U8847 ( .A(n8331), .B(n8330), .Z(n8332) );
  AND U8848 ( .A(n8333), .B(n8332), .Z(n8599) );
  XNOR U8849 ( .A(n8600), .B(n8599), .Z(n8601) );
  XOR U8850 ( .A(n8602), .B(n8601), .Z(n8606) );
  XOR U8851 ( .A(n8605), .B(n8606), .Z(n8608) );
  XOR U8852 ( .A(n8607), .B(n8608), .Z(n8618) );
  NANDN U8853 ( .A(n8335), .B(n8334), .Z(n8339) );
  NANDN U8854 ( .A(n8337), .B(n8336), .Z(n8338) );
  AND U8855 ( .A(n8339), .B(n8338), .Z(n8617) );
  XNOR U8856 ( .A(n8618), .B(n8617), .Z(n8619) );
  XOR U8857 ( .A(n8620), .B(n8619), .Z(n8624) );
  XNOR U8858 ( .A(n8623), .B(n8624), .Z(n8625) );
  NANDN U8859 ( .A(n8341), .B(n8340), .Z(n8345) );
  NANDN U8860 ( .A(n8343), .B(n8342), .Z(n8344) );
  NAND U8861 ( .A(n8345), .B(n8344), .Z(n8626) );
  XNOR U8862 ( .A(n8625), .B(n8626), .Z(n8362) );
  NANDN U8863 ( .A(n8347), .B(n8346), .Z(n8351) );
  NAND U8864 ( .A(n8349), .B(n8348), .Z(n8350) );
  NAND U8865 ( .A(n8351), .B(n8350), .Z(n8363) );
  XNOR U8866 ( .A(n8362), .B(n8363), .Z(n8364) );
  XNOR U8867 ( .A(n8365), .B(n8364), .Z(n8357) );
  XNOR U8868 ( .A(sreg[123]), .B(n8357), .Z(n8359) );
  NANDN U8869 ( .A(sreg[122]), .B(n8352), .Z(n8356) );
  NAND U8870 ( .A(n8354), .B(n8353), .Z(n8355) );
  NAND U8871 ( .A(n8356), .B(n8355), .Z(n8358) );
  XNOR U8872 ( .A(n8359), .B(n8358), .Z(c[123]) );
  NANDN U8873 ( .A(sreg[123]), .B(n8357), .Z(n8361) );
  NAND U8874 ( .A(n8359), .B(n8358), .Z(n8360) );
  NAND U8875 ( .A(n8361), .B(n8360), .Z(n8904) );
  XNOR U8876 ( .A(sreg[124]), .B(n8904), .Z(n8906) );
  NANDN U8877 ( .A(n8363), .B(n8362), .Z(n8367) );
  NANDN U8878 ( .A(n8365), .B(n8364), .Z(n8366) );
  AND U8879 ( .A(n8367), .B(n8366), .Z(n8632) );
  NANDN U8880 ( .A(n8369), .B(n8368), .Z(n8373) );
  NAND U8881 ( .A(n8371), .B(n8370), .Z(n8372) );
  AND U8882 ( .A(n8373), .B(n8372), .Z(n8642) );
  NANDN U8883 ( .A(n8375), .B(n8374), .Z(n8379) );
  OR U8884 ( .A(n8377), .B(n8376), .Z(n8378) );
  AND U8885 ( .A(n8379), .B(n8378), .Z(n8655) );
  NANDN U8886 ( .A(n8381), .B(n8380), .Z(n8385) );
  NAND U8887 ( .A(n8383), .B(n8382), .Z(n8384) );
  AND U8888 ( .A(n8385), .B(n8384), .Z(n8654) );
  NANDN U8889 ( .A(n32996), .B(n8386), .Z(n8388) );
  XOR U8890 ( .A(b[21]), .B(a[40]), .Z(n8871) );
  NANDN U8891 ( .A(n33271), .B(n8871), .Z(n8387) );
  AND U8892 ( .A(n8388), .B(n8387), .Z(n8774) );
  NANDN U8893 ( .A(n32483), .B(n8389), .Z(n8391) );
  XOR U8894 ( .A(b[19]), .B(a[42]), .Z(n8868) );
  NANDN U8895 ( .A(n32823), .B(n8868), .Z(n8390) );
  NAND U8896 ( .A(n8391), .B(n8390), .Z(n8773) );
  XNOR U8897 ( .A(n8774), .B(n8773), .Z(n8776) );
  NANDN U8898 ( .A(n33875), .B(n8392), .Z(n8394) );
  XOR U8899 ( .A(b[25]), .B(a[36]), .Z(n8862) );
  NANDN U8900 ( .A(n33994), .B(n8862), .Z(n8393) );
  AND U8901 ( .A(n8394), .B(n8393), .Z(n8752) );
  NANDN U8902 ( .A(n34223), .B(n8395), .Z(n8397) );
  XOR U8903 ( .A(b[27]), .B(a[34]), .Z(n8746) );
  NANDN U8904 ( .A(n34458), .B(n8746), .Z(n8396) );
  AND U8905 ( .A(n8397), .B(n8396), .Z(n8750) );
  NANDN U8906 ( .A(n33866), .B(n8398), .Z(n8400) );
  XOR U8907 ( .A(b[23]), .B(a[38]), .Z(n8686) );
  NANDN U8908 ( .A(n33644), .B(n8686), .Z(n8399) );
  NAND U8909 ( .A(n8400), .B(n8399), .Z(n8749) );
  XNOR U8910 ( .A(n8750), .B(n8749), .Z(n8751) );
  XNOR U8911 ( .A(n8752), .B(n8751), .Z(n8775) );
  XOR U8912 ( .A(n8776), .B(n8775), .Z(n8826) );
  NANDN U8913 ( .A(n8402), .B(n8401), .Z(n8406) );
  OR U8914 ( .A(n8404), .B(n8403), .Z(n8405) );
  AND U8915 ( .A(n8406), .B(n8405), .Z(n8824) );
  NANDN U8916 ( .A(n209), .B(n8407), .Z(n8409) );
  XOR U8917 ( .A(b[3]), .B(a[58]), .Z(n8808) );
  NANDN U8918 ( .A(n28941), .B(n8808), .Z(n8408) );
  AND U8919 ( .A(n8409), .B(n8408), .Z(n8703) );
  NANDN U8920 ( .A(n37857), .B(n8410), .Z(n8412) );
  XOR U8921 ( .A(b[55]), .B(a[6]), .Z(n8671) );
  NANDN U8922 ( .A(n37911), .B(n8671), .Z(n8411) );
  AND U8923 ( .A(n8412), .B(n8411), .Z(n8702) );
  NANDN U8924 ( .A(n8413), .B(n35309), .Z(n8415) );
  XOR U8925 ( .A(b[31]), .B(a[30]), .Z(n8805) );
  NANDN U8926 ( .A(n35145), .B(n8805), .Z(n8414) );
  NAND U8927 ( .A(n8415), .B(n8414), .Z(n8701) );
  XOR U8928 ( .A(n8702), .B(n8701), .Z(n8704) );
  XNOR U8929 ( .A(n8703), .B(n8704), .Z(n8823) );
  XNOR U8930 ( .A(n8824), .B(n8823), .Z(n8825) );
  XNOR U8931 ( .A(n8826), .B(n8825), .Z(n8841) );
  NANDN U8932 ( .A(n8417), .B(n8416), .Z(n8421) );
  NANDN U8933 ( .A(n8419), .B(n8418), .Z(n8420) );
  NAND U8934 ( .A(n8421), .B(n8420), .Z(n8842) );
  XNOR U8935 ( .A(n8841), .B(n8842), .Z(n8843) );
  NANDN U8936 ( .A(n8423), .B(n8422), .Z(n8427) );
  OR U8937 ( .A(n8425), .B(n8424), .Z(n8426) );
  NAND U8938 ( .A(n8427), .B(n8426), .Z(n8844) );
  XNOR U8939 ( .A(n8843), .B(n8844), .Z(n8653) );
  XOR U8940 ( .A(n8654), .B(n8653), .Z(n8656) );
  XNOR U8941 ( .A(n8655), .B(n8656), .Z(n8641) );
  XNOR U8942 ( .A(n8642), .B(n8641), .Z(n8643) );
  NANDN U8943 ( .A(n8429), .B(n8428), .Z(n8433) );
  NANDN U8944 ( .A(n8431), .B(n8430), .Z(n8432) );
  AND U8945 ( .A(n8433), .B(n8432), .Z(n8650) );
  NANDN U8946 ( .A(n8435), .B(n8434), .Z(n8439) );
  NAND U8947 ( .A(n8437), .B(n8436), .Z(n8438) );
  AND U8948 ( .A(n8439), .B(n8438), .Z(n8647) );
  NANDN U8949 ( .A(n210), .B(n8440), .Z(n8442) );
  XOR U8950 ( .A(b[9]), .B(a[52]), .Z(n8734) );
  NANDN U8951 ( .A(n30267), .B(n8734), .Z(n8441) );
  AND U8952 ( .A(n8442), .B(n8441), .Z(n8876) );
  NANDN U8953 ( .A(n29499), .B(n8443), .Z(n8445) );
  XOR U8954 ( .A(b[7]), .B(a[54]), .Z(n8740) );
  NANDN U8955 ( .A(n29735), .B(n8740), .Z(n8444) );
  AND U8956 ( .A(n8445), .B(n8444), .Z(n8875) );
  NANDN U8957 ( .A(n35936), .B(n8446), .Z(n8448) );
  XOR U8958 ( .A(b[37]), .B(a[24]), .Z(n8865) );
  NANDN U8959 ( .A(n36047), .B(n8865), .Z(n8447) );
  NAND U8960 ( .A(n8448), .B(n8447), .Z(n8874) );
  XOR U8961 ( .A(n8875), .B(n8874), .Z(n8877) );
  XOR U8962 ( .A(n8876), .B(n8877), .Z(n8762) );
  NANDN U8963 ( .A(n31055), .B(n8449), .Z(n8451) );
  XOR U8964 ( .A(b[13]), .B(a[48]), .Z(n8713) );
  NANDN U8965 ( .A(n31293), .B(n8713), .Z(n8450) );
  AND U8966 ( .A(n8451), .B(n8450), .Z(n8781) );
  NANDN U8967 ( .A(n30482), .B(n8452), .Z(n8454) );
  XOR U8968 ( .A(b[11]), .B(a[50]), .Z(n8731) );
  NANDN U8969 ( .A(n30891), .B(n8731), .Z(n8453) );
  AND U8970 ( .A(n8454), .B(n8453), .Z(n8780) );
  NANDN U8971 ( .A(n36210), .B(n8455), .Z(n8457) );
  XOR U8972 ( .A(b[39]), .B(a[22]), .Z(n8737) );
  NANDN U8973 ( .A(n36347), .B(n8737), .Z(n8456) );
  NAND U8974 ( .A(n8457), .B(n8456), .Z(n8779) );
  XOR U8975 ( .A(n8780), .B(n8779), .Z(n8782) );
  XNOR U8976 ( .A(n8781), .B(n8782), .Z(n8761) );
  XNOR U8977 ( .A(n8762), .B(n8761), .Z(n8764) );
  NANDN U8978 ( .A(n8459), .B(n8458), .Z(n8463) );
  OR U8979 ( .A(n8461), .B(n8460), .Z(n8462) );
  AND U8980 ( .A(n8463), .B(n8462), .Z(n8763) );
  XOR U8981 ( .A(n8764), .B(n8763), .Z(n8831) );
  NANDN U8982 ( .A(n8465), .B(n8464), .Z(n8469) );
  NANDN U8983 ( .A(n8467), .B(n8466), .Z(n8468) );
  AND U8984 ( .A(n8469), .B(n8468), .Z(n8830) );
  NANDN U8985 ( .A(n8471), .B(n8470), .Z(n8475) );
  NANDN U8986 ( .A(n8473), .B(n8472), .Z(n8474) );
  NAND U8987 ( .A(n8475), .B(n8474), .Z(n8829) );
  XOR U8988 ( .A(n8830), .B(n8829), .Z(n8832) );
  XOR U8989 ( .A(n8831), .B(n8832), .Z(n8893) );
  NANDN U8990 ( .A(n8477), .B(n8476), .Z(n8481) );
  NANDN U8991 ( .A(n8479), .B(n8478), .Z(n8480) );
  NAND U8992 ( .A(n8481), .B(n8480), .Z(n8892) );
  XNOR U8993 ( .A(n8893), .B(n8892), .Z(n8895) );
  NANDN U8994 ( .A(n8483), .B(n8482), .Z(n8487) );
  OR U8995 ( .A(n8485), .B(n8484), .Z(n8486) );
  AND U8996 ( .A(n8487), .B(n8486), .Z(n8819) );
  AND U8997 ( .A(b[0]), .B(a[60]), .Z(n8488) );
  XOR U8998 ( .A(b[1]), .B(n8488), .Z(n8490) );
  NANDN U8999 ( .A(b[0]), .B(a[59]), .Z(n8489) );
  AND U9000 ( .A(n8490), .B(n8489), .Z(n8786) );
  XOR U9001 ( .A(b[59]), .B(b[60]), .Z(n37864) );
  IV U9002 ( .A(n37864), .Z(n38248) );
  ANDN U9003 ( .B(a[0]), .A(n38248), .Z(n8804) );
  NANDN U9004 ( .A(n37974), .B(n8491), .Z(n8493) );
  XOR U9005 ( .A(b[57]), .B(a[4]), .Z(n8674) );
  NANDN U9006 ( .A(n38031), .B(n8674), .Z(n8492) );
  AND U9007 ( .A(n8493), .B(n8492), .Z(n8785) );
  XOR U9008 ( .A(n8804), .B(n8785), .Z(n8787) );
  XNOR U9009 ( .A(n8786), .B(n8787), .Z(n8817) );
  NANDN U9010 ( .A(n34634), .B(n8494), .Z(n8496) );
  XOR U9011 ( .A(b[29]), .B(a[32]), .Z(n8814) );
  NANDN U9012 ( .A(n34722), .B(n8814), .Z(n8495) );
  AND U9013 ( .A(n8496), .B(n8495), .Z(n8728) );
  NANDN U9014 ( .A(n36480), .B(n8497), .Z(n8499) );
  XOR U9015 ( .A(b[41]), .B(a[20]), .Z(n8856) );
  NANDN U9016 ( .A(n36594), .B(n8856), .Z(n8498) );
  AND U9017 ( .A(n8499), .B(n8498), .Z(n8726) );
  NANDN U9018 ( .A(n32013), .B(n8500), .Z(n8502) );
  XOR U9019 ( .A(b[17]), .B(a[44]), .Z(n8853) );
  NANDN U9020 ( .A(n32292), .B(n8853), .Z(n8501) );
  NAND U9021 ( .A(n8502), .B(n8501), .Z(n8725) );
  XNOR U9022 ( .A(n8726), .B(n8725), .Z(n8727) );
  XOR U9023 ( .A(n8728), .B(n8727), .Z(n8818) );
  XOR U9024 ( .A(n8817), .B(n8818), .Z(n8820) );
  XOR U9025 ( .A(n8819), .B(n8820), .Z(n8770) );
  NANDN U9026 ( .A(n36742), .B(n8503), .Z(n8505) );
  XOR U9027 ( .A(b[43]), .B(a[18]), .Z(n8707) );
  NANDN U9028 ( .A(n36891), .B(n8707), .Z(n8504) );
  AND U9029 ( .A(n8505), .B(n8504), .Z(n8792) );
  NANDN U9030 ( .A(n36991), .B(n8506), .Z(n8508) );
  XOR U9031 ( .A(b[45]), .B(a[16]), .Z(n8710) );
  NANDN U9032 ( .A(n37083), .B(n8710), .Z(n8507) );
  AND U9033 ( .A(n8508), .B(n8507), .Z(n8791) );
  NANDN U9034 ( .A(n31536), .B(n8509), .Z(n8511) );
  XOR U9035 ( .A(b[15]), .B(a[46]), .Z(n8859) );
  NANDN U9036 ( .A(n31925), .B(n8859), .Z(n8510) );
  NAND U9037 ( .A(n8511), .B(n8510), .Z(n8790) );
  XOR U9038 ( .A(n8791), .B(n8790), .Z(n8793) );
  XOR U9039 ( .A(n8792), .B(n8793), .Z(n8887) );
  NANDN U9040 ( .A(n37705), .B(n8512), .Z(n8514) );
  XOR U9041 ( .A(b[53]), .B(a[8]), .Z(n8719) );
  NANDN U9042 ( .A(n37778), .B(n8719), .Z(n8513) );
  AND U9043 ( .A(n8514), .B(n8513), .Z(n8697) );
  NANDN U9044 ( .A(n28889), .B(n8515), .Z(n8517) );
  XOR U9045 ( .A(b[5]), .B(a[56]), .Z(n8743) );
  NANDN U9046 ( .A(n29138), .B(n8743), .Z(n8516) );
  AND U9047 ( .A(n8517), .B(n8516), .Z(n8696) );
  NANDN U9048 ( .A(n35611), .B(n8518), .Z(n8520) );
  XOR U9049 ( .A(b[35]), .B(a[26]), .Z(n8722) );
  NANDN U9050 ( .A(n35801), .B(n8722), .Z(n8519) );
  NAND U9051 ( .A(n8520), .B(n8519), .Z(n8695) );
  XOR U9052 ( .A(n8696), .B(n8695), .Z(n8698) );
  XNOR U9053 ( .A(n8697), .B(n8698), .Z(n8886) );
  XNOR U9054 ( .A(n8887), .B(n8886), .Z(n8888) );
  NANDN U9055 ( .A(n8522), .B(n8521), .Z(n8526) );
  NANDN U9056 ( .A(n8524), .B(n8523), .Z(n8525) );
  NAND U9057 ( .A(n8526), .B(n8525), .Z(n8889) );
  XNOR U9058 ( .A(n8888), .B(n8889), .Z(n8767) );
  NANDN U9059 ( .A(n8528), .B(n8527), .Z(n8532) );
  OR U9060 ( .A(n8530), .B(n8529), .Z(n8531) );
  NAND U9061 ( .A(n8532), .B(n8531), .Z(n8768) );
  XNOR U9062 ( .A(n8767), .B(n8768), .Z(n8769) );
  XNOR U9063 ( .A(n8770), .B(n8769), .Z(n8894) );
  XOR U9064 ( .A(n8895), .B(n8894), .Z(n8662) );
  NANDN U9065 ( .A(n8534), .B(n8533), .Z(n8538) );
  OR U9066 ( .A(n8536), .B(n8535), .Z(n8537) );
  AND U9067 ( .A(n8538), .B(n8537), .Z(n8660) );
  NANDN U9068 ( .A(n8540), .B(n8539), .Z(n8544) );
  NANDN U9069 ( .A(n8542), .B(n8541), .Z(n8543) );
  AND U9070 ( .A(n8544), .B(n8543), .Z(n8659) );
  XNOR U9071 ( .A(n8660), .B(n8659), .Z(n8661) );
  XNOR U9072 ( .A(n8662), .B(n8661), .Z(n8837) );
  NANDN U9073 ( .A(n8546), .B(n8545), .Z(n8550) );
  NAND U9074 ( .A(n8548), .B(n8547), .Z(n8549) );
  AND U9075 ( .A(n8550), .B(n8549), .Z(n8668) );
  NAND U9076 ( .A(n8552), .B(n8551), .Z(n8556) );
  NAND U9077 ( .A(n8554), .B(n8553), .Z(n8555) );
  AND U9078 ( .A(n8556), .B(n8555), .Z(n8666) );
  NANDN U9079 ( .A(n8558), .B(n8557), .Z(n8562) );
  OR U9080 ( .A(n8560), .B(n8559), .Z(n8561) );
  AND U9081 ( .A(n8562), .B(n8561), .Z(n8848) );
  NANDN U9082 ( .A(n8564), .B(n8563), .Z(n8568) );
  NANDN U9083 ( .A(n8566), .B(n8565), .Z(n8567) );
  NAND U9084 ( .A(n8568), .B(n8567), .Z(n8847) );
  XNOR U9085 ( .A(n8848), .B(n8847), .Z(n8850) );
  NANDN U9086 ( .A(n8570), .B(n8569), .Z(n8574) );
  OR U9087 ( .A(n8572), .B(n8571), .Z(n8573) );
  AND U9088 ( .A(n8574), .B(n8573), .Z(n8758) );
  NOR U9089 ( .A(n8576), .B(n8575), .Z(n8882) );
  ANDN U9090 ( .B(n8577), .A(n38175), .Z(n38174) );
  NAND U9091 ( .A(n38174), .B(n8578), .Z(n8580) );
  XNOR U9092 ( .A(b[59]), .B(a[2]), .Z(n8796) );
  NANDN U9093 ( .A(n8796), .B(n38175), .Z(n8579) );
  AND U9094 ( .A(n8580), .B(n8579), .Z(n8880) );
  NAND U9095 ( .A(n35654), .B(n8581), .Z(n8583) );
  XNOR U9096 ( .A(b[33]), .B(a[28]), .Z(n8677) );
  NANDN U9097 ( .A(n8677), .B(n35655), .Z(n8582) );
  NAND U9098 ( .A(n8583), .B(n8582), .Z(n8881) );
  XOR U9099 ( .A(n8880), .B(n8881), .Z(n8883) );
  XOR U9100 ( .A(n8882), .B(n8883), .Z(n8756) );
  NANDN U9101 ( .A(n211), .B(n8584), .Z(n8586) );
  XOR U9102 ( .A(b[47]), .B(a[14]), .Z(n8680) );
  NANDN U9103 ( .A(n37172), .B(n8680), .Z(n8585) );
  AND U9104 ( .A(n8586), .B(n8585), .Z(n8692) );
  NANDN U9105 ( .A(n212), .B(n8587), .Z(n8589) );
  XOR U9106 ( .A(b[49]), .B(a[12]), .Z(n8683) );
  NANDN U9107 ( .A(n37432), .B(n8683), .Z(n8588) );
  AND U9108 ( .A(n8589), .B(n8588), .Z(n8690) );
  NANDN U9109 ( .A(n37526), .B(n8590), .Z(n8592) );
  XOR U9110 ( .A(b[51]), .B(a[10]), .Z(n8716) );
  NANDN U9111 ( .A(n37605), .B(n8716), .Z(n8591) );
  NAND U9112 ( .A(n8592), .B(n8591), .Z(n8689) );
  XNOR U9113 ( .A(n8690), .B(n8689), .Z(n8691) );
  XNOR U9114 ( .A(n8692), .B(n8691), .Z(n8755) );
  XNOR U9115 ( .A(n8756), .B(n8755), .Z(n8757) );
  XNOR U9116 ( .A(n8758), .B(n8757), .Z(n8849) );
  XNOR U9117 ( .A(n8850), .B(n8849), .Z(n8665) );
  XNOR U9118 ( .A(n8666), .B(n8665), .Z(n8667) );
  XOR U9119 ( .A(n8668), .B(n8667), .Z(n8836) );
  NANDN U9120 ( .A(n8594), .B(n8593), .Z(n8598) );
  NANDN U9121 ( .A(n8596), .B(n8595), .Z(n8597) );
  AND U9122 ( .A(n8598), .B(n8597), .Z(n8835) );
  XOR U9123 ( .A(n8836), .B(n8835), .Z(n8838) );
  XOR U9124 ( .A(n8837), .B(n8838), .Z(n8648) );
  XNOR U9125 ( .A(n8647), .B(n8648), .Z(n8649) );
  XOR U9126 ( .A(n8650), .B(n8649), .Z(n8644) );
  XNOR U9127 ( .A(n8643), .B(n8644), .Z(n8637) );
  NANDN U9128 ( .A(n8600), .B(n8599), .Z(n8604) );
  NANDN U9129 ( .A(n8602), .B(n8601), .Z(n8603) );
  AND U9130 ( .A(n8604), .B(n8603), .Z(n8636) );
  NANDN U9131 ( .A(n8606), .B(n8605), .Z(n8610) );
  OR U9132 ( .A(n8608), .B(n8607), .Z(n8609) );
  NAND U9133 ( .A(n8610), .B(n8609), .Z(n8635) );
  XOR U9134 ( .A(n8636), .B(n8635), .Z(n8638) );
  XNOR U9135 ( .A(n8637), .B(n8638), .Z(n8901) );
  NAND U9136 ( .A(n8612), .B(n8611), .Z(n8616) );
  NAND U9137 ( .A(n8614), .B(n8613), .Z(n8615) );
  AND U9138 ( .A(n8616), .B(n8615), .Z(n8899) );
  NANDN U9139 ( .A(n8618), .B(n8617), .Z(n8622) );
  NANDN U9140 ( .A(n8620), .B(n8619), .Z(n8621) );
  AND U9141 ( .A(n8622), .B(n8621), .Z(n8898) );
  XNOR U9142 ( .A(n8899), .B(n8898), .Z(n8900) );
  XOR U9143 ( .A(n8901), .B(n8900), .Z(n8630) );
  NANDN U9144 ( .A(n8624), .B(n8623), .Z(n8628) );
  NANDN U9145 ( .A(n8626), .B(n8625), .Z(n8627) );
  NAND U9146 ( .A(n8628), .B(n8627), .Z(n8629) );
  XNOR U9147 ( .A(n8630), .B(n8629), .Z(n8631) );
  XNOR U9148 ( .A(n8632), .B(n8631), .Z(n8905) );
  XNOR U9149 ( .A(n8906), .B(n8905), .Z(c[124]) );
  NANDN U9150 ( .A(n8630), .B(n8629), .Z(n8634) );
  NANDN U9151 ( .A(n8632), .B(n8631), .Z(n8633) );
  AND U9152 ( .A(n8634), .B(n8633), .Z(n8917) );
  NANDN U9153 ( .A(n8636), .B(n8635), .Z(n8640) );
  NANDN U9154 ( .A(n8638), .B(n8637), .Z(n8639) );
  AND U9155 ( .A(n8640), .B(n8639), .Z(n8922) );
  NANDN U9156 ( .A(n8642), .B(n8641), .Z(n8646) );
  NANDN U9157 ( .A(n8644), .B(n8643), .Z(n8645) );
  AND U9158 ( .A(n8646), .B(n8645), .Z(n8921) );
  NANDN U9159 ( .A(n8648), .B(n8647), .Z(n8652) );
  NANDN U9160 ( .A(n8650), .B(n8649), .Z(n8651) );
  AND U9161 ( .A(n8652), .B(n8651), .Z(n9183) );
  NANDN U9162 ( .A(n8654), .B(n8653), .Z(n8658) );
  OR U9163 ( .A(n8656), .B(n8655), .Z(n8657) );
  AND U9164 ( .A(n8658), .B(n8657), .Z(n9182) );
  XNOR U9165 ( .A(n9183), .B(n9182), .Z(n9184) );
  NANDN U9166 ( .A(n8660), .B(n8659), .Z(n8664) );
  NANDN U9167 ( .A(n8662), .B(n8661), .Z(n8663) );
  AND U9168 ( .A(n8664), .B(n8663), .Z(n8929) );
  NANDN U9169 ( .A(n8666), .B(n8665), .Z(n8670) );
  NAND U9170 ( .A(n8668), .B(n8667), .Z(n8669) );
  AND U9171 ( .A(n8670), .B(n8669), .Z(n8927) );
  NANDN U9172 ( .A(n37857), .B(n8671), .Z(n8673) );
  XOR U9173 ( .A(b[55]), .B(a[7]), .Z(n9134) );
  NANDN U9174 ( .A(n37911), .B(n9134), .Z(n8672) );
  AND U9175 ( .A(n8673), .B(n8672), .Z(n9027) );
  NANDN U9176 ( .A(n37974), .B(n8674), .Z(n8676) );
  XOR U9177 ( .A(b[57]), .B(a[5]), .Z(n8989) );
  NANDN U9178 ( .A(n38031), .B(n8989), .Z(n8675) );
  AND U9179 ( .A(n8676), .B(n8675), .Z(n9026) );
  NANDN U9180 ( .A(n8677), .B(n35654), .Z(n8679) );
  XOR U9181 ( .A(b[33]), .B(a[29]), .Z(n8971) );
  NANDN U9182 ( .A(n35456), .B(n8971), .Z(n8678) );
  NAND U9183 ( .A(n8679), .B(n8678), .Z(n9025) );
  XOR U9184 ( .A(n9026), .B(n9025), .Z(n9028) );
  XOR U9185 ( .A(n9027), .B(n9028), .Z(n9095) );
  NANDN U9186 ( .A(n211), .B(n8680), .Z(n8682) );
  XOR U9187 ( .A(b[47]), .B(a[15]), .Z(n8998) );
  NANDN U9188 ( .A(n37172), .B(n8998), .Z(n8681) );
  AND U9189 ( .A(n8682), .B(n8681), .Z(n9009) );
  NANDN U9190 ( .A(n212), .B(n8683), .Z(n8685) );
  XOR U9191 ( .A(b[49]), .B(a[13]), .Z(n9001) );
  NANDN U9192 ( .A(n37432), .B(n9001), .Z(n8684) );
  AND U9193 ( .A(n8685), .B(n8684), .Z(n9008) );
  NANDN U9194 ( .A(n33866), .B(n8686), .Z(n8688) );
  XOR U9195 ( .A(b[23]), .B(a[39]), .Z(n8977) );
  NANDN U9196 ( .A(n33644), .B(n8977), .Z(n8687) );
  NAND U9197 ( .A(n8688), .B(n8687), .Z(n9007) );
  XOR U9198 ( .A(n9008), .B(n9007), .Z(n9010) );
  XNOR U9199 ( .A(n9009), .B(n9010), .Z(n9094) );
  XNOR U9200 ( .A(n9095), .B(n9094), .Z(n9097) );
  NANDN U9201 ( .A(n8690), .B(n8689), .Z(n8694) );
  NANDN U9202 ( .A(n8692), .B(n8691), .Z(n8693) );
  AND U9203 ( .A(n8694), .B(n8693), .Z(n9096) );
  XOR U9204 ( .A(n9097), .B(n9096), .Z(n9067) );
  NANDN U9205 ( .A(n8696), .B(n8695), .Z(n8700) );
  OR U9206 ( .A(n8698), .B(n8697), .Z(n8699) );
  AND U9207 ( .A(n8700), .B(n8699), .Z(n9065) );
  NANDN U9208 ( .A(n8702), .B(n8701), .Z(n8706) );
  OR U9209 ( .A(n8704), .B(n8703), .Z(n8705) );
  NAND U9210 ( .A(n8706), .B(n8705), .Z(n9064) );
  XNOR U9211 ( .A(n9065), .B(n9064), .Z(n9066) );
  XOR U9212 ( .A(n9067), .B(n9066), .Z(n9084) );
  NANDN U9213 ( .A(n36742), .B(n8707), .Z(n8709) );
  XOR U9214 ( .A(b[43]), .B(a[19]), .Z(n9137) );
  NANDN U9215 ( .A(n36891), .B(n9137), .Z(n8708) );
  AND U9216 ( .A(n8709), .B(n8708), .Z(n9142) );
  NANDN U9217 ( .A(n36991), .B(n8710), .Z(n8712) );
  XOR U9218 ( .A(b[45]), .B(a[17]), .Z(n9125) );
  NANDN U9219 ( .A(n37083), .B(n9125), .Z(n8711) );
  AND U9220 ( .A(n8712), .B(n8711), .Z(n9141) );
  NANDN U9221 ( .A(n31055), .B(n8713), .Z(n8715) );
  XOR U9222 ( .A(b[13]), .B(a[49]), .Z(n9158) );
  NANDN U9223 ( .A(n31293), .B(n9158), .Z(n8714) );
  NAND U9224 ( .A(n8715), .B(n8714), .Z(n9140) );
  XOR U9225 ( .A(n9141), .B(n9140), .Z(n9143) );
  XOR U9226 ( .A(n9142), .B(n9143), .Z(n8955) );
  NANDN U9227 ( .A(n37526), .B(n8716), .Z(n8718) );
  XOR U9228 ( .A(b[51]), .B(a[11]), .Z(n9161) );
  NANDN U9229 ( .A(n37605), .B(n9161), .Z(n8717) );
  AND U9230 ( .A(n8718), .B(n8717), .Z(n9033) );
  NANDN U9231 ( .A(n37705), .B(n8719), .Z(n8721) );
  XOR U9232 ( .A(b[53]), .B(a[9]), .Z(n9131) );
  NANDN U9233 ( .A(n37778), .B(n9131), .Z(n8720) );
  AND U9234 ( .A(n8721), .B(n8720), .Z(n9032) );
  NANDN U9235 ( .A(n35611), .B(n8722), .Z(n8724) );
  XOR U9236 ( .A(b[35]), .B(a[27]), .Z(n9113) );
  NANDN U9237 ( .A(n35801), .B(n9113), .Z(n8723) );
  NAND U9238 ( .A(n8724), .B(n8723), .Z(n9031) );
  XOR U9239 ( .A(n9032), .B(n9031), .Z(n9034) );
  XNOR U9240 ( .A(n9033), .B(n9034), .Z(n8954) );
  XNOR U9241 ( .A(n8955), .B(n8954), .Z(n8956) );
  NANDN U9242 ( .A(n8726), .B(n8725), .Z(n8730) );
  NANDN U9243 ( .A(n8728), .B(n8727), .Z(n8729) );
  NAND U9244 ( .A(n8730), .B(n8729), .Z(n8957) );
  XNOR U9245 ( .A(n8956), .B(n8957), .Z(n9083) );
  NANDN U9246 ( .A(n30482), .B(n8731), .Z(n8733) );
  XOR U9247 ( .A(b[11]), .B(a[51]), .Z(n9146) );
  NANDN U9248 ( .A(n30891), .B(n9146), .Z(n8732) );
  AND U9249 ( .A(n8733), .B(n8732), .Z(n9166) );
  NANDN U9250 ( .A(n210), .B(n8734), .Z(n8736) );
  XOR U9251 ( .A(b[9]), .B(a[53]), .Z(n9149) );
  NANDN U9252 ( .A(n30267), .B(n9149), .Z(n8735) );
  AND U9253 ( .A(n8736), .B(n8735), .Z(n9165) );
  NANDN U9254 ( .A(n36210), .B(n8737), .Z(n8739) );
  XOR U9255 ( .A(b[39]), .B(a[23]), .Z(n9152) );
  NANDN U9256 ( .A(n36347), .B(n9152), .Z(n8738) );
  NAND U9257 ( .A(n8739), .B(n8738), .Z(n9164) );
  XOR U9258 ( .A(n9165), .B(n9164), .Z(n9167) );
  XOR U9259 ( .A(n9166), .B(n9167), .Z(n8949) );
  NANDN U9260 ( .A(n29499), .B(n8740), .Z(n8742) );
  XOR U9261 ( .A(b[7]), .B(a[55]), .Z(n8992) );
  NANDN U9262 ( .A(n29735), .B(n8992), .Z(n8741) );
  AND U9263 ( .A(n8742), .B(n8741), .Z(n9118) );
  NANDN U9264 ( .A(n28889), .B(n8743), .Z(n8745) );
  XOR U9265 ( .A(b[5]), .B(a[57]), .Z(n9110) );
  NANDN U9266 ( .A(n29138), .B(n9110), .Z(n8744) );
  AND U9267 ( .A(n8745), .B(n8744), .Z(n9117) );
  NANDN U9268 ( .A(n34223), .B(n8746), .Z(n8748) );
  XOR U9269 ( .A(b[27]), .B(a[35]), .Z(n9049) );
  NANDN U9270 ( .A(n34458), .B(n9049), .Z(n8747) );
  NAND U9271 ( .A(n8748), .B(n8747), .Z(n9116) );
  XOR U9272 ( .A(n9117), .B(n9116), .Z(n9119) );
  XNOR U9273 ( .A(n9118), .B(n9119), .Z(n8948) );
  XNOR U9274 ( .A(n8949), .B(n8948), .Z(n8950) );
  NANDN U9275 ( .A(n8750), .B(n8749), .Z(n8754) );
  NANDN U9276 ( .A(n8752), .B(n8751), .Z(n8753) );
  NAND U9277 ( .A(n8754), .B(n8753), .Z(n8951) );
  XNOR U9278 ( .A(n8950), .B(n8951), .Z(n9082) );
  XOR U9279 ( .A(n9083), .B(n9082), .Z(n9085) );
  XNOR U9280 ( .A(n9084), .B(n9085), .Z(n9015) );
  NANDN U9281 ( .A(n8756), .B(n8755), .Z(n8760) );
  NANDN U9282 ( .A(n8758), .B(n8757), .Z(n8759) );
  AND U9283 ( .A(n8760), .B(n8759), .Z(n9014) );
  NANDN U9284 ( .A(n8762), .B(n8761), .Z(n8766) );
  NAND U9285 ( .A(n8764), .B(n8763), .Z(n8765) );
  AND U9286 ( .A(n8766), .B(n8765), .Z(n9013) );
  XOR U9287 ( .A(n9014), .B(n9013), .Z(n9016) );
  XOR U9288 ( .A(n9015), .B(n9016), .Z(n8938) );
  NANDN U9289 ( .A(n8768), .B(n8767), .Z(n8772) );
  NANDN U9290 ( .A(n8770), .B(n8769), .Z(n8771) );
  NAND U9291 ( .A(n8772), .B(n8771), .Z(n8939) );
  XOR U9292 ( .A(n8938), .B(n8939), .Z(n8940) );
  NANDN U9293 ( .A(n8774), .B(n8773), .Z(n8778) );
  NAND U9294 ( .A(n8776), .B(n8775), .Z(n8777) );
  AND U9295 ( .A(n8778), .B(n8777), .Z(n9078) );
  NANDN U9296 ( .A(n8780), .B(n8779), .Z(n8784) );
  OR U9297 ( .A(n8782), .B(n8781), .Z(n8783) );
  AND U9298 ( .A(n8784), .B(n8783), .Z(n9077) );
  NANDN U9299 ( .A(n8785), .B(n8804), .Z(n8789) );
  NANDN U9300 ( .A(n8787), .B(n8786), .Z(n8788) );
  NAND U9301 ( .A(n8789), .B(n8788), .Z(n9076) );
  XOR U9302 ( .A(n9077), .B(n9076), .Z(n9079) );
  XOR U9303 ( .A(n9078), .B(n9079), .Z(n8945) );
  NANDN U9304 ( .A(n8791), .B(n8790), .Z(n8795) );
  OR U9305 ( .A(n8793), .B(n8792), .Z(n8794) );
  AND U9306 ( .A(n8795), .B(n8794), .Z(n9090) );
  NANDN U9307 ( .A(n8796), .B(n38174), .Z(n8798) );
  XOR U9308 ( .A(b[59]), .B(a[3]), .Z(n9046) );
  NANDN U9309 ( .A(n38130), .B(n9046), .Z(n8797) );
  AND U9310 ( .A(n8798), .B(n8797), .Z(n8966) );
  XOR U9311 ( .A(b[61]), .B(b[60]), .Z(n9106) );
  XOR U9312 ( .A(b[61]), .B(a[0]), .Z(n8799) );
  NAND U9313 ( .A(n9106), .B(n8799), .Z(n8800) );
  OR U9314 ( .A(n8800), .B(n37864), .Z(n8802) );
  XOR U9315 ( .A(b[61]), .B(a[1]), .Z(n9107) );
  NAND U9316 ( .A(n37864), .B(n9107), .Z(n8801) );
  AND U9317 ( .A(n8802), .B(n8801), .Z(n8967) );
  XOR U9318 ( .A(n8966), .B(n8967), .Z(n9102) );
  NAND U9319 ( .A(b[59]), .B(b[60]), .Z(n8803) );
  NAND U9320 ( .A(b[61]), .B(n8803), .Z(n38273) );
  NOR U9321 ( .A(n38273), .B(n8804), .Z(n9101) );
  NAND U9322 ( .A(n35309), .B(n8805), .Z(n8807) );
  XNOR U9323 ( .A(b[31]), .B(a[31]), .Z(n8974) );
  NANDN U9324 ( .A(n8974), .B(n35310), .Z(n8806) );
  AND U9325 ( .A(n8807), .B(n8806), .Z(n9100) );
  XOR U9326 ( .A(n9101), .B(n9100), .Z(n9103) );
  XOR U9327 ( .A(n9102), .B(n9103), .Z(n9089) );
  NAND U9328 ( .A(n9942), .B(n8808), .Z(n8810) );
  XNOR U9329 ( .A(b[3]), .B(a[59]), .Z(n8968) );
  NANDN U9330 ( .A(n8968), .B(n9653), .Z(n8809) );
  NAND U9331 ( .A(n8810), .B(n8809), .Z(n8985) );
  NAND U9332 ( .A(b[0]), .B(a[61]), .Z(n8811) );
  XNOR U9333 ( .A(b[1]), .B(n8811), .Z(n8813) );
  NANDN U9334 ( .A(b[0]), .B(a[60]), .Z(n8812) );
  NAND U9335 ( .A(n8813), .B(n8812), .Z(n8984) );
  NANDN U9336 ( .A(n34634), .B(n8814), .Z(n8816) );
  XOR U9337 ( .A(b[29]), .B(a[33]), .Z(n9052) );
  NANDN U9338 ( .A(n34722), .B(n9052), .Z(n8815) );
  NAND U9339 ( .A(n8816), .B(n8815), .Z(n8983) );
  XNOR U9340 ( .A(n8984), .B(n8983), .Z(n8986) );
  XOR U9341 ( .A(n8985), .B(n8986), .Z(n9088) );
  XOR U9342 ( .A(n9089), .B(n9088), .Z(n9091) );
  XOR U9343 ( .A(n9090), .B(n9091), .Z(n8943) );
  NANDN U9344 ( .A(n8818), .B(n8817), .Z(n8822) );
  OR U9345 ( .A(n8820), .B(n8819), .Z(n8821) );
  AND U9346 ( .A(n8822), .B(n8821), .Z(n8942) );
  XNOR U9347 ( .A(n8943), .B(n8942), .Z(n8944) );
  XNOR U9348 ( .A(n8945), .B(n8944), .Z(n9021) );
  NANDN U9349 ( .A(n8824), .B(n8823), .Z(n8828) );
  NANDN U9350 ( .A(n8826), .B(n8825), .Z(n8827) );
  AND U9351 ( .A(n8828), .B(n8827), .Z(n9020) );
  NANDN U9352 ( .A(n8830), .B(n8829), .Z(n8834) );
  OR U9353 ( .A(n8832), .B(n8831), .Z(n8833) );
  AND U9354 ( .A(n8834), .B(n8833), .Z(n9019) );
  XOR U9355 ( .A(n9020), .B(n9019), .Z(n9022) );
  XOR U9356 ( .A(n9021), .B(n9022), .Z(n8941) );
  XNOR U9357 ( .A(n8940), .B(n8941), .Z(n8926) );
  XNOR U9358 ( .A(n8927), .B(n8926), .Z(n8928) );
  XOR U9359 ( .A(n8929), .B(n8928), .Z(n9179) );
  NANDN U9360 ( .A(n8836), .B(n8835), .Z(n8840) );
  NANDN U9361 ( .A(n8838), .B(n8837), .Z(n8839) );
  AND U9362 ( .A(n8840), .B(n8839), .Z(n9177) );
  NANDN U9363 ( .A(n8842), .B(n8841), .Z(n8846) );
  NANDN U9364 ( .A(n8844), .B(n8843), .Z(n8845) );
  AND U9365 ( .A(n8846), .B(n8845), .Z(n8934) );
  NANDN U9366 ( .A(n8848), .B(n8847), .Z(n8852) );
  NAND U9367 ( .A(n8850), .B(n8849), .Z(n8851) );
  AND U9368 ( .A(n8852), .B(n8851), .Z(n9173) );
  NANDN U9369 ( .A(n32013), .B(n8853), .Z(n8855) );
  XOR U9370 ( .A(b[17]), .B(a[45]), .Z(n9004) );
  NANDN U9371 ( .A(n32292), .B(n9004), .Z(n8854) );
  AND U9372 ( .A(n8855), .B(n8854), .Z(n9039) );
  NANDN U9373 ( .A(n36480), .B(n8856), .Z(n8858) );
  XOR U9374 ( .A(b[41]), .B(a[21]), .Z(n9122) );
  NANDN U9375 ( .A(n36594), .B(n9122), .Z(n8857) );
  AND U9376 ( .A(n8858), .B(n8857), .Z(n9038) );
  NANDN U9377 ( .A(n31536), .B(n8859), .Z(n8861) );
  XOR U9378 ( .A(b[15]), .B(a[47]), .Z(n9155) );
  NANDN U9379 ( .A(n31925), .B(n9155), .Z(n8860) );
  NAND U9380 ( .A(n8861), .B(n8860), .Z(n9037) );
  XOR U9381 ( .A(n9038), .B(n9037), .Z(n9040) );
  XOR U9382 ( .A(n9039), .B(n9040), .Z(n9060) );
  NANDN U9383 ( .A(n33875), .B(n8862), .Z(n8864) );
  XOR U9384 ( .A(b[25]), .B(a[37]), .Z(n9055) );
  NANDN U9385 ( .A(n33994), .B(n9055), .Z(n8863) );
  AND U9386 ( .A(n8864), .B(n8863), .Z(n8962) );
  NANDN U9387 ( .A(n35936), .B(n8865), .Z(n8867) );
  XOR U9388 ( .A(b[37]), .B(a[25]), .Z(n8995) );
  NANDN U9389 ( .A(n36047), .B(n8995), .Z(n8866) );
  AND U9390 ( .A(n8867), .B(n8866), .Z(n8961) );
  NANDN U9391 ( .A(n32483), .B(n8868), .Z(n8870) );
  XOR U9392 ( .A(b[19]), .B(a[43]), .Z(n9128) );
  NANDN U9393 ( .A(n32823), .B(n9128), .Z(n8869) );
  NAND U9394 ( .A(n8870), .B(n8869), .Z(n8960) );
  XOR U9395 ( .A(n8961), .B(n8960), .Z(n8963) );
  XOR U9396 ( .A(n8962), .B(n8963), .Z(n9059) );
  NAND U9397 ( .A(n33413), .B(n8871), .Z(n8873) );
  XNOR U9398 ( .A(b[21]), .B(a[41]), .Z(n8980) );
  NANDN U9399 ( .A(n8980), .B(n33414), .Z(n8872) );
  AND U9400 ( .A(n8873), .B(n8872), .Z(n9058) );
  XOR U9401 ( .A(n9059), .B(n9058), .Z(n9061) );
  XOR U9402 ( .A(n9060), .B(n9061), .Z(n9072) );
  NANDN U9403 ( .A(n8875), .B(n8874), .Z(n8879) );
  OR U9404 ( .A(n8877), .B(n8876), .Z(n8878) );
  AND U9405 ( .A(n8879), .B(n8878), .Z(n9071) );
  NANDN U9406 ( .A(n8881), .B(n8880), .Z(n8885) );
  OR U9407 ( .A(n8883), .B(n8882), .Z(n8884) );
  AND U9408 ( .A(n8885), .B(n8884), .Z(n9070) );
  XOR U9409 ( .A(n9071), .B(n9070), .Z(n9073) );
  XOR U9410 ( .A(n9072), .B(n9073), .Z(n9171) );
  NANDN U9411 ( .A(n8887), .B(n8886), .Z(n8891) );
  NANDN U9412 ( .A(n8889), .B(n8888), .Z(n8890) );
  NAND U9413 ( .A(n8891), .B(n8890), .Z(n9170) );
  XNOR U9414 ( .A(n9171), .B(n9170), .Z(n9172) );
  XOR U9415 ( .A(n9173), .B(n9172), .Z(n8933) );
  NANDN U9416 ( .A(n8893), .B(n8892), .Z(n8897) );
  NAND U9417 ( .A(n8895), .B(n8894), .Z(n8896) );
  AND U9418 ( .A(n8897), .B(n8896), .Z(n8932) );
  XOR U9419 ( .A(n8933), .B(n8932), .Z(n8935) );
  XNOR U9420 ( .A(n8934), .B(n8935), .Z(n9176) );
  XNOR U9421 ( .A(n9177), .B(n9176), .Z(n9178) );
  XOR U9422 ( .A(n9179), .B(n9178), .Z(n9185) );
  XNOR U9423 ( .A(n9184), .B(n9185), .Z(n8920) );
  XOR U9424 ( .A(n8921), .B(n8920), .Z(n8923) );
  XOR U9425 ( .A(n8922), .B(n8923), .Z(n8915) );
  NANDN U9426 ( .A(n8899), .B(n8898), .Z(n8903) );
  NAND U9427 ( .A(n8901), .B(n8900), .Z(n8902) );
  AND U9428 ( .A(n8903), .B(n8902), .Z(n8914) );
  XNOR U9429 ( .A(n8915), .B(n8914), .Z(n8916) );
  XNOR U9430 ( .A(n8917), .B(n8916), .Z(n8909) );
  XNOR U9431 ( .A(sreg[125]), .B(n8909), .Z(n8911) );
  NANDN U9432 ( .A(sreg[124]), .B(n8904), .Z(n8908) );
  NAND U9433 ( .A(n8906), .B(n8905), .Z(n8907) );
  NAND U9434 ( .A(n8908), .B(n8907), .Z(n8910) );
  XNOR U9435 ( .A(n8911), .B(n8910), .Z(c[125]) );
  NANDN U9436 ( .A(sreg[125]), .B(n8909), .Z(n8913) );
  NAND U9437 ( .A(n8911), .B(n8910), .Z(n8912) );
  NAND U9438 ( .A(n8913), .B(n8912), .Z(n9466) );
  XNOR U9439 ( .A(sreg[126]), .B(n9466), .Z(n9468) );
  NANDN U9440 ( .A(n8915), .B(n8914), .Z(n8919) );
  NANDN U9441 ( .A(n8917), .B(n8916), .Z(n8918) );
  AND U9442 ( .A(n8919), .B(n8918), .Z(n9191) );
  NANDN U9443 ( .A(n8921), .B(n8920), .Z(n8925) );
  OR U9444 ( .A(n8923), .B(n8922), .Z(n8924) );
  AND U9445 ( .A(n8925), .B(n8924), .Z(n9188) );
  NANDN U9446 ( .A(n8927), .B(n8926), .Z(n8931) );
  NAND U9447 ( .A(n8929), .B(n8928), .Z(n8930) );
  AND U9448 ( .A(n8931), .B(n8930), .Z(n9201) );
  NANDN U9449 ( .A(n8933), .B(n8932), .Z(n8937) );
  NANDN U9450 ( .A(n8935), .B(n8934), .Z(n8936) );
  AND U9451 ( .A(n8937), .B(n8936), .Z(n9200) );
  XNOR U9452 ( .A(n9201), .B(n9200), .Z(n9202) );
  NANDN U9453 ( .A(n8943), .B(n8942), .Z(n8947) );
  NANDN U9454 ( .A(n8945), .B(n8944), .Z(n8946) );
  AND U9455 ( .A(n8947), .B(n8946), .Z(n9215) );
  NANDN U9456 ( .A(n8949), .B(n8948), .Z(n8953) );
  NANDN U9457 ( .A(n8951), .B(n8950), .Z(n8952) );
  AND U9458 ( .A(n8953), .B(n8952), .Z(n9442) );
  NANDN U9459 ( .A(n8955), .B(n8954), .Z(n8959) );
  NANDN U9460 ( .A(n8957), .B(n8956), .Z(n8958) );
  NAND U9461 ( .A(n8959), .B(n8958), .Z(n9443) );
  XNOR U9462 ( .A(n9442), .B(n9443), .Z(n9445) );
  NANDN U9463 ( .A(n8961), .B(n8960), .Z(n8965) );
  OR U9464 ( .A(n8963), .B(n8962), .Z(n8964) );
  AND U9465 ( .A(n8965), .B(n8964), .Z(n9421) );
  NOR U9466 ( .A(n8967), .B(n8966), .Z(n9342) );
  NANDN U9467 ( .A(n8968), .B(n9942), .Z(n8970) );
  XNOR U9468 ( .A(b[3]), .B(a[60]), .Z(n9254) );
  NANDN U9469 ( .A(n9254), .B(n9653), .Z(n8969) );
  AND U9470 ( .A(n8970), .B(n8969), .Z(n9340) );
  NAND U9471 ( .A(n35654), .B(n8971), .Z(n8973) );
  XNOR U9472 ( .A(b[33]), .B(a[30]), .Z(n9328) );
  NANDN U9473 ( .A(n9328), .B(n35655), .Z(n8972) );
  NAND U9474 ( .A(n8973), .B(n8972), .Z(n9341) );
  XOR U9475 ( .A(n9340), .B(n9341), .Z(n9343) );
  XOR U9476 ( .A(n9342), .B(n9343), .Z(n9419) );
  NANDN U9477 ( .A(n8974), .B(n35309), .Z(n8976) );
  XOR U9478 ( .A(b[31]), .B(a[32]), .Z(n9409) );
  NANDN U9479 ( .A(n35145), .B(n9409), .Z(n8975) );
  AND U9480 ( .A(n8976), .B(n8975), .Z(n9263) );
  NANDN U9481 ( .A(n33866), .B(n8977), .Z(n8979) );
  XOR U9482 ( .A(b[23]), .B(a[40]), .Z(n9257) );
  NANDN U9483 ( .A(n33644), .B(n9257), .Z(n8978) );
  AND U9484 ( .A(n8979), .B(n8978), .Z(n9261) );
  NANDN U9485 ( .A(n8980), .B(n33413), .Z(n8982) );
  XOR U9486 ( .A(b[21]), .B(a[42]), .Z(n9394) );
  NANDN U9487 ( .A(n33271), .B(n9394), .Z(n8981) );
  NAND U9488 ( .A(n8982), .B(n8981), .Z(n9260) );
  XNOR U9489 ( .A(n9261), .B(n9260), .Z(n9262) );
  XNOR U9490 ( .A(n9263), .B(n9262), .Z(n9418) );
  XNOR U9491 ( .A(n9419), .B(n9418), .Z(n9420) );
  XNOR U9492 ( .A(n9421), .B(n9420), .Z(n9462) );
  NANDN U9493 ( .A(n8984), .B(n8983), .Z(n8988) );
  NAND U9494 ( .A(n8986), .B(n8985), .Z(n8987) );
  AND U9495 ( .A(n8988), .B(n8987), .Z(n9461) );
  NANDN U9496 ( .A(n37974), .B(n8989), .Z(n8991) );
  XOR U9497 ( .A(b[57]), .B(a[6]), .Z(n9403) );
  NANDN U9498 ( .A(n38031), .B(n9403), .Z(n8990) );
  AND U9499 ( .A(n8991), .B(n8990), .Z(n9310) );
  NANDN U9500 ( .A(n29499), .B(n8992), .Z(n8994) );
  XOR U9501 ( .A(b[7]), .B(a[56]), .Z(n9290) );
  NANDN U9502 ( .A(n29735), .B(n9290), .Z(n8993) );
  AND U9503 ( .A(n8994), .B(n8993), .Z(n9309) );
  NANDN U9504 ( .A(n35936), .B(n8995), .Z(n8997) );
  XOR U9505 ( .A(b[37]), .B(a[26]), .Z(n9331) );
  NANDN U9506 ( .A(n36047), .B(n9331), .Z(n8996) );
  NAND U9507 ( .A(n8997), .B(n8996), .Z(n9308) );
  XOR U9508 ( .A(n9309), .B(n9308), .Z(n9311) );
  XOR U9509 ( .A(n9310), .B(n9311), .Z(n9437) );
  NANDN U9510 ( .A(n211), .B(n8998), .Z(n9000) );
  XOR U9511 ( .A(b[47]), .B(a[16]), .Z(n9227) );
  NANDN U9512 ( .A(n37172), .B(n9227), .Z(n8999) );
  AND U9513 ( .A(n9000), .B(n8999), .Z(n9316) );
  NANDN U9514 ( .A(n212), .B(n9001), .Z(n9003) );
  XOR U9515 ( .A(b[49]), .B(a[14]), .Z(n9230) );
  NANDN U9516 ( .A(n37432), .B(n9230), .Z(n9002) );
  AND U9517 ( .A(n9003), .B(n9002), .Z(n9315) );
  NANDN U9518 ( .A(n32013), .B(n9004), .Z(n9006) );
  XOR U9519 ( .A(b[17]), .B(a[46]), .Z(n9400) );
  NANDN U9520 ( .A(n32292), .B(n9400), .Z(n9005) );
  NAND U9521 ( .A(n9006), .B(n9005), .Z(n9314) );
  XOR U9522 ( .A(n9315), .B(n9314), .Z(n9317) );
  XNOR U9523 ( .A(n9316), .B(n9317), .Z(n9436) );
  XNOR U9524 ( .A(n9437), .B(n9436), .Z(n9439) );
  NANDN U9525 ( .A(n9008), .B(n9007), .Z(n9012) );
  OR U9526 ( .A(n9010), .B(n9009), .Z(n9011) );
  AND U9527 ( .A(n9012), .B(n9011), .Z(n9438) );
  XNOR U9528 ( .A(n9439), .B(n9438), .Z(n9460) );
  XOR U9529 ( .A(n9461), .B(n9460), .Z(n9463) );
  XNOR U9530 ( .A(n9462), .B(n9463), .Z(n9444) );
  XOR U9531 ( .A(n9445), .B(n9444), .Z(n9213) );
  NANDN U9532 ( .A(n9014), .B(n9013), .Z(n9018) );
  NANDN U9533 ( .A(n9016), .B(n9015), .Z(n9017) );
  AND U9534 ( .A(n9018), .B(n9017), .Z(n9212) );
  XNOR U9535 ( .A(n9213), .B(n9212), .Z(n9214) );
  XNOR U9536 ( .A(n9215), .B(n9214), .Z(n9206) );
  XNOR U9537 ( .A(n9207), .B(n9206), .Z(n9208) );
  NANDN U9538 ( .A(n9020), .B(n9019), .Z(n9024) );
  NANDN U9539 ( .A(n9022), .B(n9021), .Z(n9023) );
  AND U9540 ( .A(n9024), .B(n9023), .Z(n9377) );
  NANDN U9541 ( .A(n9026), .B(n9025), .Z(n9030) );
  OR U9542 ( .A(n9028), .B(n9027), .Z(n9029) );
  AND U9543 ( .A(n9030), .B(n9029), .Z(n9359) );
  NANDN U9544 ( .A(n9032), .B(n9031), .Z(n9036) );
  OR U9545 ( .A(n9034), .B(n9033), .Z(n9035) );
  NAND U9546 ( .A(n9036), .B(n9035), .Z(n9358) );
  XNOR U9547 ( .A(n9359), .B(n9358), .Z(n9361) );
  NANDN U9548 ( .A(n9038), .B(n9037), .Z(n9042) );
  OR U9549 ( .A(n9040), .B(n9039), .Z(n9041) );
  AND U9550 ( .A(n9042), .B(n9041), .Z(n9355) );
  NAND U9551 ( .A(b[0]), .B(a[62]), .Z(n9043) );
  XNOR U9552 ( .A(b[1]), .B(n9043), .Z(n9045) );
  NANDN U9553 ( .A(b[0]), .B(a[61]), .Z(n9044) );
  NAND U9554 ( .A(n9045), .B(n9044), .Z(n9415) );
  XOR U9555 ( .A(b[61]), .B(b[62]), .Z(n38264) );
  IV U9556 ( .A(n38264), .Z(n38279) );
  ANDN U9557 ( .B(a[0]), .A(n38279), .Z(n9412) );
  IV U9558 ( .A(n38174), .Z(n38090) );
  NANDN U9559 ( .A(n38090), .B(n9046), .Z(n9048) );
  XOR U9560 ( .A(b[59]), .B(a[4]), .Z(n9406) );
  NANDN U9561 ( .A(n38130), .B(n9406), .Z(n9047) );
  AND U9562 ( .A(n9048), .B(n9047), .Z(n9413) );
  XNOR U9563 ( .A(n9412), .B(n9413), .Z(n9414) );
  XNOR U9564 ( .A(n9415), .B(n9414), .Z(n9352) );
  NANDN U9565 ( .A(n34223), .B(n9049), .Z(n9051) );
  XOR U9566 ( .A(b[27]), .B(a[36]), .Z(n9233) );
  NANDN U9567 ( .A(n34458), .B(n9233), .Z(n9050) );
  AND U9568 ( .A(n9051), .B(n9050), .Z(n9349) );
  NANDN U9569 ( .A(n34634), .B(n9052), .Z(n9054) );
  XOR U9570 ( .A(b[29]), .B(a[34]), .Z(n9284) );
  NANDN U9571 ( .A(n34722), .B(n9284), .Z(n9053) );
  AND U9572 ( .A(n9054), .B(n9053), .Z(n9347) );
  NANDN U9573 ( .A(n33875), .B(n9055), .Z(n9057) );
  XOR U9574 ( .A(b[25]), .B(a[38]), .Z(n9397) );
  NANDN U9575 ( .A(n33994), .B(n9397), .Z(n9056) );
  NAND U9576 ( .A(n9057), .B(n9056), .Z(n9346) );
  XNOR U9577 ( .A(n9347), .B(n9346), .Z(n9348) );
  XOR U9578 ( .A(n9349), .B(n9348), .Z(n9353) );
  XNOR U9579 ( .A(n9352), .B(n9353), .Z(n9354) );
  XNOR U9580 ( .A(n9355), .B(n9354), .Z(n9360) );
  XOR U9581 ( .A(n9361), .B(n9360), .Z(n9449) );
  NANDN U9582 ( .A(n9059), .B(n9058), .Z(n9063) );
  OR U9583 ( .A(n9061), .B(n9060), .Z(n9062) );
  NAND U9584 ( .A(n9063), .B(n9062), .Z(n9448) );
  XNOR U9585 ( .A(n9449), .B(n9448), .Z(n9450) );
  NANDN U9586 ( .A(n9065), .B(n9064), .Z(n9069) );
  NANDN U9587 ( .A(n9067), .B(n9066), .Z(n9068) );
  NAND U9588 ( .A(n9069), .B(n9068), .Z(n9451) );
  XNOR U9589 ( .A(n9450), .B(n9451), .Z(n9371) );
  NANDN U9590 ( .A(n9071), .B(n9070), .Z(n9075) );
  OR U9591 ( .A(n9073), .B(n9072), .Z(n9074) );
  AND U9592 ( .A(n9075), .B(n9074), .Z(n9368) );
  NANDN U9593 ( .A(n9077), .B(n9076), .Z(n9081) );
  OR U9594 ( .A(n9079), .B(n9078), .Z(n9080) );
  NAND U9595 ( .A(n9081), .B(n9080), .Z(n9369) );
  XNOR U9596 ( .A(n9368), .B(n9369), .Z(n9370) );
  XOR U9597 ( .A(n9371), .B(n9370), .Z(n9381) );
  NAND U9598 ( .A(n9083), .B(n9082), .Z(n9087) );
  NAND U9599 ( .A(n9085), .B(n9084), .Z(n9086) );
  AND U9600 ( .A(n9087), .B(n9086), .Z(n9379) );
  NANDN U9601 ( .A(n9089), .B(n9088), .Z(n9093) );
  OR U9602 ( .A(n9091), .B(n9090), .Z(n9092) );
  AND U9603 ( .A(n9093), .B(n9092), .Z(n9365) );
  NANDN U9604 ( .A(n9095), .B(n9094), .Z(n9099) );
  NAND U9605 ( .A(n9097), .B(n9096), .Z(n9098) );
  AND U9606 ( .A(n9099), .B(n9098), .Z(n9364) );
  XNOR U9607 ( .A(n9365), .B(n9364), .Z(n9367) );
  NANDN U9608 ( .A(n9101), .B(n9100), .Z(n9105) );
  OR U9609 ( .A(n9103), .B(n9102), .Z(n9104) );
  AND U9610 ( .A(n9105), .B(n9104), .Z(n9383) );
  ANDN U9611 ( .B(n9106), .A(n37864), .Z(n37921) );
  IV U9612 ( .A(n37921), .Z(n38247) );
  NANDN U9613 ( .A(n38247), .B(n9107), .Z(n9109) );
  XOR U9614 ( .A(b[61]), .B(a[2]), .Z(n9320) );
  NANDN U9615 ( .A(n38248), .B(n9320), .Z(n9108) );
  AND U9616 ( .A(n9109), .B(n9108), .Z(n9274) );
  NANDN U9617 ( .A(n28889), .B(n9110), .Z(n9112) );
  XOR U9618 ( .A(b[5]), .B(a[58]), .Z(n9251) );
  NANDN U9619 ( .A(n29138), .B(n9251), .Z(n9111) );
  AND U9620 ( .A(n9112), .B(n9111), .Z(n9273) );
  NANDN U9621 ( .A(n35611), .B(n9113), .Z(n9115) );
  XOR U9622 ( .A(b[35]), .B(a[28]), .Z(n9224) );
  NANDN U9623 ( .A(n35801), .B(n9224), .Z(n9114) );
  NAND U9624 ( .A(n9115), .B(n9114), .Z(n9272) );
  XOR U9625 ( .A(n9273), .B(n9272), .Z(n9275) );
  XNOR U9626 ( .A(n9274), .B(n9275), .Z(n9382) );
  XNOR U9627 ( .A(n9383), .B(n9382), .Z(n9384) );
  NANDN U9628 ( .A(n9117), .B(n9116), .Z(n9121) );
  OR U9629 ( .A(n9119), .B(n9118), .Z(n9120) );
  NAND U9630 ( .A(n9121), .B(n9120), .Z(n9385) );
  XOR U9631 ( .A(n9384), .B(n9385), .Z(n9456) );
  NANDN U9632 ( .A(n36480), .B(n9122), .Z(n9124) );
  XOR U9633 ( .A(b[41]), .B(a[22]), .Z(n9242) );
  NANDN U9634 ( .A(n36594), .B(n9242), .Z(n9123) );
  AND U9635 ( .A(n9124), .B(n9123), .Z(n9238) );
  NANDN U9636 ( .A(n36991), .B(n9125), .Z(n9127) );
  XOR U9637 ( .A(b[45]), .B(a[18]), .Z(n9287) );
  NANDN U9638 ( .A(n37083), .B(n9287), .Z(n9126) );
  AND U9639 ( .A(n9127), .B(n9126), .Z(n9237) );
  NANDN U9640 ( .A(n32483), .B(n9128), .Z(n9130) );
  XOR U9641 ( .A(b[19]), .B(a[44]), .Z(n9293) );
  NANDN U9642 ( .A(n32823), .B(n9293), .Z(n9129) );
  NAND U9643 ( .A(n9130), .B(n9129), .Z(n9236) );
  XOR U9644 ( .A(n9237), .B(n9236), .Z(n9239) );
  XOR U9645 ( .A(n9238), .B(n9239), .Z(n9431) );
  NANDN U9646 ( .A(n37705), .B(n9131), .Z(n9133) );
  XOR U9647 ( .A(b[53]), .B(a[10]), .Z(n9221) );
  NANDN U9648 ( .A(n37778), .B(n9221), .Z(n9132) );
  AND U9649 ( .A(n9133), .B(n9132), .Z(n9268) );
  NANDN U9650 ( .A(n37857), .B(n9134), .Z(n9136) );
  XOR U9651 ( .A(b[55]), .B(a[8]), .Z(n9281) );
  NANDN U9652 ( .A(n37911), .B(n9281), .Z(n9135) );
  AND U9653 ( .A(n9136), .B(n9135), .Z(n9267) );
  NANDN U9654 ( .A(n36742), .B(n9137), .Z(n9139) );
  XOR U9655 ( .A(b[43]), .B(a[20]), .Z(n9245) );
  NANDN U9656 ( .A(n36891), .B(n9245), .Z(n9138) );
  NAND U9657 ( .A(n9139), .B(n9138), .Z(n9266) );
  XOR U9658 ( .A(n9267), .B(n9266), .Z(n9269) );
  XNOR U9659 ( .A(n9268), .B(n9269), .Z(n9430) );
  XNOR U9660 ( .A(n9431), .B(n9430), .Z(n9432) );
  NANDN U9661 ( .A(n9141), .B(n9140), .Z(n9145) );
  OR U9662 ( .A(n9143), .B(n9142), .Z(n9144) );
  NAND U9663 ( .A(n9145), .B(n9144), .Z(n9433) );
  XOR U9664 ( .A(n9432), .B(n9433), .Z(n9455) );
  NANDN U9665 ( .A(n30482), .B(n9146), .Z(n9148) );
  XOR U9666 ( .A(b[11]), .B(a[52]), .Z(n9337) );
  NANDN U9667 ( .A(n30891), .B(n9337), .Z(n9147) );
  AND U9668 ( .A(n9148), .B(n9147), .Z(n9304) );
  NANDN U9669 ( .A(n210), .B(n9149), .Z(n9151) );
  XOR U9670 ( .A(b[9]), .B(a[54]), .Z(n9248) );
  NANDN U9671 ( .A(n30267), .B(n9248), .Z(n9150) );
  AND U9672 ( .A(n9151), .B(n9150), .Z(n9303) );
  NANDN U9673 ( .A(n36210), .B(n9152), .Z(n9154) );
  XOR U9674 ( .A(b[39]), .B(a[24]), .Z(n9334) );
  NANDN U9675 ( .A(n36347), .B(n9334), .Z(n9153) );
  NAND U9676 ( .A(n9154), .B(n9153), .Z(n9302) );
  XOR U9677 ( .A(n9303), .B(n9302), .Z(n9305) );
  XOR U9678 ( .A(n9304), .B(n9305), .Z(n9425) );
  NANDN U9679 ( .A(n31536), .B(n9155), .Z(n9157) );
  XOR U9680 ( .A(b[15]), .B(a[48]), .Z(n9391) );
  NANDN U9681 ( .A(n31925), .B(n9391), .Z(n9156) );
  AND U9682 ( .A(n9157), .B(n9156), .Z(n9298) );
  NANDN U9683 ( .A(n31055), .B(n9158), .Z(n9160) );
  XOR U9684 ( .A(b[13]), .B(a[50]), .Z(n9388) );
  NANDN U9685 ( .A(n31293), .B(n9388), .Z(n9159) );
  AND U9686 ( .A(n9160), .B(n9159), .Z(n9297) );
  NANDN U9687 ( .A(n37526), .B(n9161), .Z(n9163) );
  XOR U9688 ( .A(b[51]), .B(a[12]), .Z(n9218) );
  NANDN U9689 ( .A(n37605), .B(n9218), .Z(n9162) );
  NAND U9690 ( .A(n9163), .B(n9162), .Z(n9296) );
  XOR U9691 ( .A(n9297), .B(n9296), .Z(n9299) );
  XNOR U9692 ( .A(n9298), .B(n9299), .Z(n9424) );
  XNOR U9693 ( .A(n9425), .B(n9424), .Z(n9427) );
  NANDN U9694 ( .A(n9165), .B(n9164), .Z(n9169) );
  OR U9695 ( .A(n9167), .B(n9166), .Z(n9168) );
  AND U9696 ( .A(n9169), .B(n9168), .Z(n9426) );
  XNOR U9697 ( .A(n9427), .B(n9426), .Z(n9454) );
  XOR U9698 ( .A(n9455), .B(n9454), .Z(n9457) );
  XOR U9699 ( .A(n9456), .B(n9457), .Z(n9366) );
  XOR U9700 ( .A(n9367), .B(n9366), .Z(n9378) );
  XOR U9701 ( .A(n9379), .B(n9378), .Z(n9380) );
  XOR U9702 ( .A(n9381), .B(n9380), .Z(n9374) );
  NANDN U9703 ( .A(n9171), .B(n9170), .Z(n9175) );
  NAND U9704 ( .A(n9173), .B(n9172), .Z(n9174) );
  NAND U9705 ( .A(n9175), .B(n9174), .Z(n9375) );
  XOR U9706 ( .A(n9374), .B(n9375), .Z(n9376) );
  XOR U9707 ( .A(n9377), .B(n9376), .Z(n9209) );
  XOR U9708 ( .A(n9208), .B(n9209), .Z(n9203) );
  XNOR U9709 ( .A(n9202), .B(n9203), .Z(n9194) );
  NANDN U9710 ( .A(n9177), .B(n9176), .Z(n9181) );
  NANDN U9711 ( .A(n9179), .B(n9178), .Z(n9180) );
  NAND U9712 ( .A(n9181), .B(n9180), .Z(n9195) );
  XNOR U9713 ( .A(n9194), .B(n9195), .Z(n9196) );
  NANDN U9714 ( .A(n9183), .B(n9182), .Z(n9187) );
  NANDN U9715 ( .A(n9185), .B(n9184), .Z(n9186) );
  NAND U9716 ( .A(n9187), .B(n9186), .Z(n9197) );
  XOR U9717 ( .A(n9196), .B(n9197), .Z(n9189) );
  XNOR U9718 ( .A(n9188), .B(n9189), .Z(n9190) );
  XNOR U9719 ( .A(n9191), .B(n9190), .Z(n9467) );
  XNOR U9720 ( .A(n9468), .B(n9467), .Z(c[126]) );
  NANDN U9721 ( .A(n9189), .B(n9188), .Z(n9193) );
  NANDN U9722 ( .A(n9191), .B(n9190), .Z(n9192) );
  AND U9723 ( .A(n9193), .B(n9192), .Z(n9479) );
  NANDN U9724 ( .A(n9195), .B(n9194), .Z(n9199) );
  NANDN U9725 ( .A(n9197), .B(n9196), .Z(n9198) );
  AND U9726 ( .A(n9199), .B(n9198), .Z(n9477) );
  NANDN U9727 ( .A(n9201), .B(n9200), .Z(n9205) );
  NANDN U9728 ( .A(n9203), .B(n9202), .Z(n9204) );
  AND U9729 ( .A(n9205), .B(n9204), .Z(n9758) );
  NANDN U9730 ( .A(n9207), .B(n9206), .Z(n9211) );
  NANDN U9731 ( .A(n9209), .B(n9208), .Z(n9210) );
  AND U9732 ( .A(n9211), .B(n9210), .Z(n9756) );
  NANDN U9733 ( .A(n9213), .B(n9212), .Z(n9217) );
  NANDN U9734 ( .A(n9215), .B(n9214), .Z(n9216) );
  AND U9735 ( .A(n9217), .B(n9216), .Z(n9497) );
  NANDN U9736 ( .A(n37526), .B(n9218), .Z(n9220) );
  XOR U9737 ( .A(b[51]), .B(a[13]), .Z(n9662) );
  NANDN U9738 ( .A(n37605), .B(n9662), .Z(n9219) );
  AND U9739 ( .A(n9220), .B(n9219), .Z(n9706) );
  NANDN U9740 ( .A(n37705), .B(n9221), .Z(n9223) );
  XOR U9741 ( .A(b[53]), .B(a[11]), .Z(n9578) );
  NANDN U9742 ( .A(n37778), .B(n9578), .Z(n9222) );
  AND U9743 ( .A(n9223), .B(n9222), .Z(n9705) );
  NANDN U9744 ( .A(n35611), .B(n9224), .Z(n9226) );
  XOR U9745 ( .A(b[35]), .B(a[29]), .Z(n9656) );
  NANDN U9746 ( .A(n35801), .B(n9656), .Z(n9225) );
  NAND U9747 ( .A(n9226), .B(n9225), .Z(n9704) );
  XOR U9748 ( .A(n9705), .B(n9704), .Z(n9707) );
  XOR U9749 ( .A(n9706), .B(n9707), .Z(n9639) );
  NANDN U9750 ( .A(n211), .B(n9227), .Z(n9229) );
  XOR U9751 ( .A(b[47]), .B(a[17]), .Z(n9659) );
  NANDN U9752 ( .A(n37172), .B(n9659), .Z(n9228) );
  AND U9753 ( .A(n9229), .B(n9228), .Z(n9565) );
  NANDN U9754 ( .A(n212), .B(n9230), .Z(n9232) );
  XOR U9755 ( .A(b[49]), .B(a[15]), .Z(n9590) );
  NANDN U9756 ( .A(n37432), .B(n9590), .Z(n9231) );
  AND U9757 ( .A(n9232), .B(n9231), .Z(n9564) );
  NANDN U9758 ( .A(n34223), .B(n9233), .Z(n9235) );
  XOR U9759 ( .A(b[27]), .B(a[37]), .Z(n9557) );
  NANDN U9760 ( .A(n34458), .B(n9557), .Z(n9234) );
  NAND U9761 ( .A(n9235), .B(n9234), .Z(n9563) );
  XOR U9762 ( .A(n9564), .B(n9563), .Z(n9566) );
  XNOR U9763 ( .A(n9565), .B(n9566), .Z(n9638) );
  XNOR U9764 ( .A(n9639), .B(n9638), .Z(n9641) );
  NANDN U9765 ( .A(n9237), .B(n9236), .Z(n9241) );
  OR U9766 ( .A(n9239), .B(n9238), .Z(n9240) );
  AND U9767 ( .A(n9241), .B(n9240), .Z(n9640) );
  XOR U9768 ( .A(n9641), .B(n9640), .Z(n9633) );
  NANDN U9769 ( .A(n36480), .B(n9242), .Z(n9244) );
  XOR U9770 ( .A(b[41]), .B(a[23]), .Z(n9683) );
  NANDN U9771 ( .A(n36594), .B(n9683), .Z(n9243) );
  AND U9772 ( .A(n9244), .B(n9243), .Z(n9595) );
  NANDN U9773 ( .A(n36742), .B(n9245), .Z(n9247) );
  XOR U9774 ( .A(b[43]), .B(a[21]), .Z(n9668) );
  NANDN U9775 ( .A(n36891), .B(n9668), .Z(n9246) );
  AND U9776 ( .A(n9247), .B(n9246), .Z(n9594) );
  NANDN U9777 ( .A(n210), .B(n9248), .Z(n9250) );
  XOR U9778 ( .A(b[9]), .B(a[55]), .Z(n9575) );
  NANDN U9779 ( .A(n30267), .B(n9575), .Z(n9249) );
  NAND U9780 ( .A(n9250), .B(n9249), .Z(n9593) );
  XOR U9781 ( .A(n9594), .B(n9593), .Z(n9596) );
  XOR U9782 ( .A(n9595), .B(n9596), .Z(n9693) );
  NANDN U9783 ( .A(n28889), .B(n9251), .Z(n9253) );
  XOR U9784 ( .A(b[5]), .B(a[59]), .Z(n9722) );
  NANDN U9785 ( .A(n29138), .B(n9722), .Z(n9252) );
  AND U9786 ( .A(n9253), .B(n9252), .Z(n9646) );
  NANDN U9787 ( .A(n9254), .B(n9942), .Z(n9256) );
  XOR U9788 ( .A(b[3]), .B(a[61]), .Z(n9652) );
  NANDN U9789 ( .A(n28941), .B(n9652), .Z(n9255) );
  AND U9790 ( .A(n9256), .B(n9255), .Z(n9645) );
  NANDN U9791 ( .A(n33866), .B(n9257), .Z(n9259) );
  XOR U9792 ( .A(b[23]), .B(a[41]), .Z(n9560) );
  NANDN U9793 ( .A(n33644), .B(n9560), .Z(n9258) );
  NAND U9794 ( .A(n9259), .B(n9258), .Z(n9644) );
  XOR U9795 ( .A(n9645), .B(n9644), .Z(n9647) );
  XNOR U9796 ( .A(n9646), .B(n9647), .Z(n9692) );
  XNOR U9797 ( .A(n9693), .B(n9692), .Z(n9695) );
  NANDN U9798 ( .A(n9261), .B(n9260), .Z(n9265) );
  NANDN U9799 ( .A(n9263), .B(n9262), .Z(n9264) );
  AND U9800 ( .A(n9265), .B(n9264), .Z(n9694) );
  XOR U9801 ( .A(n9695), .B(n9694), .Z(n9527) );
  NANDN U9802 ( .A(n9267), .B(n9266), .Z(n9271) );
  OR U9803 ( .A(n9269), .B(n9268), .Z(n9270) );
  AND U9804 ( .A(n9271), .B(n9270), .Z(n9525) );
  NANDN U9805 ( .A(n9273), .B(n9272), .Z(n9277) );
  OR U9806 ( .A(n9275), .B(n9274), .Z(n9276) );
  NAND U9807 ( .A(n9277), .B(n9276), .Z(n9524) );
  XNOR U9808 ( .A(n9525), .B(n9524), .Z(n9526) );
  XNOR U9809 ( .A(n9527), .B(n9526), .Z(n9632) );
  XNOR U9810 ( .A(n9633), .B(n9632), .Z(n9635) );
  NAND U9811 ( .A(b[0]), .B(a[63]), .Z(n9278) );
  XNOR U9812 ( .A(b[1]), .B(n9278), .Z(n9280) );
  NANDN U9813 ( .A(b[0]), .B(a[62]), .Z(n9279) );
  NAND U9814 ( .A(n9280), .B(n9279), .Z(n9701) );
  NANDN U9815 ( .A(n37857), .B(n9281), .Z(n9283) );
  XOR U9816 ( .A(b[55]), .B(a[9]), .Z(n9677) );
  NANDN U9817 ( .A(n37911), .B(n9677), .Z(n9282) );
  AND U9818 ( .A(n9283), .B(n9282), .Z(n9699) );
  NANDN U9819 ( .A(n34634), .B(n9284), .Z(n9286) );
  XOR U9820 ( .A(b[29]), .B(a[35]), .Z(n9554) );
  NANDN U9821 ( .A(n34722), .B(n9554), .Z(n9285) );
  NAND U9822 ( .A(n9286), .B(n9285), .Z(n9698) );
  XOR U9823 ( .A(n9699), .B(n9698), .Z(n9700) );
  XOR U9824 ( .A(n9701), .B(n9700), .Z(n9738) );
  NANDN U9825 ( .A(n36991), .B(n9287), .Z(n9289) );
  XOR U9826 ( .A(b[45]), .B(a[19]), .Z(n9671) );
  NANDN U9827 ( .A(n37083), .B(n9671), .Z(n9288) );
  AND U9828 ( .A(n9289), .B(n9288), .Z(n9622) );
  NANDN U9829 ( .A(n29499), .B(n9290), .Z(n9292) );
  XOR U9830 ( .A(b[7]), .B(a[57]), .Z(n9614) );
  NANDN U9831 ( .A(n29735), .B(n9614), .Z(n9291) );
  AND U9832 ( .A(n9292), .B(n9291), .Z(n9621) );
  NANDN U9833 ( .A(n32483), .B(n9293), .Z(n9295) );
  XOR U9834 ( .A(b[19]), .B(a[45]), .Z(n9548) );
  NANDN U9835 ( .A(n32823), .B(n9548), .Z(n9294) );
  NAND U9836 ( .A(n9295), .B(n9294), .Z(n9620) );
  XOR U9837 ( .A(n9621), .B(n9620), .Z(n9623) );
  XNOR U9838 ( .A(n9622), .B(n9623), .Z(n9737) );
  XNOR U9839 ( .A(n9738), .B(n9737), .Z(n9740) );
  NANDN U9840 ( .A(n9297), .B(n9296), .Z(n9301) );
  OR U9841 ( .A(n9299), .B(n9298), .Z(n9300) );
  AND U9842 ( .A(n9301), .B(n9300), .Z(n9739) );
  XOR U9843 ( .A(n9740), .B(n9739), .Z(n9734) );
  NANDN U9844 ( .A(n9303), .B(n9302), .Z(n9307) );
  OR U9845 ( .A(n9305), .B(n9304), .Z(n9306) );
  AND U9846 ( .A(n9307), .B(n9306), .Z(n9732) );
  NANDN U9847 ( .A(n9309), .B(n9308), .Z(n9313) );
  OR U9848 ( .A(n9311), .B(n9310), .Z(n9312) );
  NAND U9849 ( .A(n9313), .B(n9312), .Z(n9731) );
  XNOR U9850 ( .A(n9732), .B(n9731), .Z(n9733) );
  XNOR U9851 ( .A(n9734), .B(n9733), .Z(n9634) );
  XOR U9852 ( .A(n9635), .B(n9634), .Z(n9513) );
  NANDN U9853 ( .A(n9315), .B(n9314), .Z(n9319) );
  OR U9854 ( .A(n9317), .B(n9316), .Z(n9318) );
  AND U9855 ( .A(n9319), .B(n9318), .Z(n9538) );
  NANDN U9856 ( .A(n38247), .B(n9320), .Z(n9322) );
  XOR U9857 ( .A(b[61]), .B(a[3]), .Z(n9719) );
  NANDN U9858 ( .A(n38248), .B(n9719), .Z(n9321) );
  AND U9859 ( .A(n9322), .B(n9321), .Z(n9651) );
  XOR U9860 ( .A(b[62]), .B(b[63]), .Z(n9323) );
  ANDN U9861 ( .B(n9323), .A(n38264), .Z(n38262) );
  IV U9862 ( .A(n38262), .Z(n38278) );
  XOR U9863 ( .A(a[0]), .B(b[63]), .Z(n9324) );
  NANDN U9864 ( .A(n38278), .B(n9324), .Z(n9326) );
  XOR U9865 ( .A(b[63]), .B(a[1]), .Z(n9725) );
  ANDN U9866 ( .B(n9725), .A(n38279), .Z(n9325) );
  ANDN U9867 ( .B(n9326), .A(n9325), .Z(n9650) );
  XOR U9868 ( .A(n9651), .B(n9650), .Z(n9607) );
  NAND U9869 ( .A(b[61]), .B(b[62]), .Z(n38296) );
  ANDN U9870 ( .B(n38296), .A(n9412), .Z(n9327) );
  AND U9871 ( .A(b[63]), .B(n9327), .Z(n9606) );
  NANDN U9872 ( .A(n9328), .B(n35654), .Z(n9330) );
  XNOR U9873 ( .A(b[33]), .B(a[31]), .Z(n9545) );
  NANDN U9874 ( .A(n9545), .B(n35655), .Z(n9329) );
  AND U9875 ( .A(n9330), .B(n9329), .Z(n9605) );
  XOR U9876 ( .A(n9606), .B(n9605), .Z(n9608) );
  XOR U9877 ( .A(n9607), .B(n9608), .Z(n9537) );
  NANDN U9878 ( .A(n35936), .B(n9331), .Z(n9333) );
  XOR U9879 ( .A(b[37]), .B(a[27]), .Z(n9728) );
  NANDN U9880 ( .A(n36047), .B(n9728), .Z(n9332) );
  AND U9881 ( .A(n9333), .B(n9332), .Z(n9689) );
  NANDN U9882 ( .A(n36210), .B(n9334), .Z(n9336) );
  XOR U9883 ( .A(b[39]), .B(a[25]), .Z(n9617) );
  NANDN U9884 ( .A(n36347), .B(n9617), .Z(n9335) );
  AND U9885 ( .A(n9336), .B(n9335), .Z(n9687) );
  NANDN U9886 ( .A(n30482), .B(n9337), .Z(n9339) );
  XOR U9887 ( .A(b[11]), .B(a[53]), .Z(n9587) );
  NANDN U9888 ( .A(n30891), .B(n9587), .Z(n9338) );
  NAND U9889 ( .A(n9339), .B(n9338), .Z(n9686) );
  XNOR U9890 ( .A(n9687), .B(n9686), .Z(n9688) );
  XNOR U9891 ( .A(n9689), .B(n9688), .Z(n9536) );
  XOR U9892 ( .A(n9537), .B(n9536), .Z(n9539) );
  XOR U9893 ( .A(n9538), .B(n9539), .Z(n9746) );
  NANDN U9894 ( .A(n9341), .B(n9340), .Z(n9345) );
  OR U9895 ( .A(n9343), .B(n9342), .Z(n9344) );
  AND U9896 ( .A(n9345), .B(n9344), .Z(n9744) );
  NANDN U9897 ( .A(n9347), .B(n9346), .Z(n9351) );
  NANDN U9898 ( .A(n9349), .B(n9348), .Z(n9350) );
  AND U9899 ( .A(n9351), .B(n9350), .Z(n9743) );
  XNOR U9900 ( .A(n9744), .B(n9743), .Z(n9745) );
  XNOR U9901 ( .A(n9746), .B(n9745), .Z(n9626) );
  NANDN U9902 ( .A(n9353), .B(n9352), .Z(n9357) );
  NANDN U9903 ( .A(n9355), .B(n9354), .Z(n9356) );
  NAND U9904 ( .A(n9357), .B(n9356), .Z(n9627) );
  XNOR U9905 ( .A(n9626), .B(n9627), .Z(n9628) );
  NANDN U9906 ( .A(n9359), .B(n9358), .Z(n9363) );
  NAND U9907 ( .A(n9361), .B(n9360), .Z(n9362) );
  NAND U9908 ( .A(n9363), .B(n9362), .Z(n9629) );
  XNOR U9909 ( .A(n9628), .B(n9629), .Z(n9512) );
  XNOR U9910 ( .A(n9513), .B(n9512), .Z(n9515) );
  XOR U9911 ( .A(n9515), .B(n9514), .Z(n9495) );
  NANDN U9912 ( .A(n9369), .B(n9368), .Z(n9373) );
  NAND U9913 ( .A(n9371), .B(n9370), .Z(n9372) );
  AND U9914 ( .A(n9373), .B(n9372), .Z(n9494) );
  XNOR U9915 ( .A(n9495), .B(n9494), .Z(n9496) );
  XOR U9916 ( .A(n9497), .B(n9496), .Z(n9485) );
  NANDN U9917 ( .A(n9383), .B(n9382), .Z(n9387) );
  NANDN U9918 ( .A(n9385), .B(n9384), .Z(n9386) );
  AND U9919 ( .A(n9387), .B(n9386), .Z(n9521) );
  NANDN U9920 ( .A(n31055), .B(n9388), .Z(n9390) );
  XOR U9921 ( .A(b[13]), .B(a[51]), .Z(n9584) );
  NANDN U9922 ( .A(n31293), .B(n9584), .Z(n9389) );
  AND U9923 ( .A(n9390), .B(n9389), .Z(n9600) );
  NANDN U9924 ( .A(n31536), .B(n9391), .Z(n9393) );
  XOR U9925 ( .A(b[15]), .B(a[49]), .Z(n9665) );
  NANDN U9926 ( .A(n31925), .B(n9665), .Z(n9392) );
  NAND U9927 ( .A(n9393), .B(n9392), .Z(n9599) );
  XNOR U9928 ( .A(n9600), .B(n9599), .Z(n9602) );
  NANDN U9929 ( .A(n32996), .B(n9394), .Z(n9396) );
  XOR U9930 ( .A(b[21]), .B(a[43]), .Z(n9542) );
  NANDN U9931 ( .A(n33271), .B(n9542), .Z(n9395) );
  AND U9932 ( .A(n9396), .B(n9395), .Z(n9713) );
  NANDN U9933 ( .A(n33875), .B(n9397), .Z(n9399) );
  XOR U9934 ( .A(b[25]), .B(a[39]), .Z(n9551) );
  NANDN U9935 ( .A(n33994), .B(n9551), .Z(n9398) );
  AND U9936 ( .A(n9399), .B(n9398), .Z(n9711) );
  NANDN U9937 ( .A(n32013), .B(n9400), .Z(n9402) );
  XOR U9938 ( .A(b[17]), .B(a[47]), .Z(n9674) );
  NANDN U9939 ( .A(n32292), .B(n9674), .Z(n9401) );
  NAND U9940 ( .A(n9402), .B(n9401), .Z(n9710) );
  XNOR U9941 ( .A(n9711), .B(n9710), .Z(n9712) );
  XNOR U9942 ( .A(n9713), .B(n9712), .Z(n9601) );
  XOR U9943 ( .A(n9602), .B(n9601), .Z(n9533) );
  NANDN U9944 ( .A(n37974), .B(n9403), .Z(n9405) );
  XOR U9945 ( .A(b[57]), .B(a[7]), .Z(n9680) );
  NANDN U9946 ( .A(n38031), .B(n9680), .Z(n9404) );
  AND U9947 ( .A(n9405), .B(n9404), .Z(n9571) );
  NANDN U9948 ( .A(n38090), .B(n9406), .Z(n9408) );
  XOR U9949 ( .A(b[59]), .B(a[5]), .Z(n9611) );
  NANDN U9950 ( .A(n38130), .B(n9611), .Z(n9407) );
  AND U9951 ( .A(n9408), .B(n9407), .Z(n9570) );
  NANDN U9952 ( .A(n34909), .B(n9409), .Z(n9411) );
  XOR U9953 ( .A(b[31]), .B(a[33]), .Z(n9581) );
  NANDN U9954 ( .A(n35145), .B(n9581), .Z(n9410) );
  NAND U9955 ( .A(n9411), .B(n9410), .Z(n9569) );
  XOR U9956 ( .A(n9570), .B(n9569), .Z(n9572) );
  XOR U9957 ( .A(n9571), .B(n9572), .Z(n9531) );
  NANDN U9958 ( .A(n9413), .B(n9412), .Z(n9417) );
  NANDN U9959 ( .A(n9415), .B(n9414), .Z(n9416) );
  AND U9960 ( .A(n9417), .B(n9416), .Z(n9530) );
  XNOR U9961 ( .A(n9531), .B(n9530), .Z(n9532) );
  XNOR U9962 ( .A(n9533), .B(n9532), .Z(n9518) );
  NANDN U9963 ( .A(n9419), .B(n9418), .Z(n9423) );
  NANDN U9964 ( .A(n9421), .B(n9420), .Z(n9422) );
  NAND U9965 ( .A(n9423), .B(n9422), .Z(n9519) );
  XNOR U9966 ( .A(n9518), .B(n9519), .Z(n9520) );
  XNOR U9967 ( .A(n9521), .B(n9520), .Z(n9500) );
  NANDN U9968 ( .A(n9425), .B(n9424), .Z(n9429) );
  NAND U9969 ( .A(n9427), .B(n9426), .Z(n9428) );
  AND U9970 ( .A(n9429), .B(n9428), .Z(n9752) );
  NANDN U9971 ( .A(n9431), .B(n9430), .Z(n9435) );
  NANDN U9972 ( .A(n9433), .B(n9432), .Z(n9434) );
  AND U9973 ( .A(n9435), .B(n9434), .Z(n9750) );
  NANDN U9974 ( .A(n9437), .B(n9436), .Z(n9441) );
  NAND U9975 ( .A(n9439), .B(n9438), .Z(n9440) );
  NAND U9976 ( .A(n9441), .B(n9440), .Z(n9749) );
  XNOR U9977 ( .A(n9750), .B(n9749), .Z(n9751) );
  XOR U9978 ( .A(n9752), .B(n9751), .Z(n9501) );
  XNOR U9979 ( .A(n9500), .B(n9501), .Z(n9503) );
  NANDN U9980 ( .A(n9443), .B(n9442), .Z(n9447) );
  NAND U9981 ( .A(n9445), .B(n9444), .Z(n9446) );
  AND U9982 ( .A(n9447), .B(n9446), .Z(n9502) );
  XOR U9983 ( .A(n9503), .B(n9502), .Z(n9489) );
  NANDN U9984 ( .A(n9449), .B(n9448), .Z(n9453) );
  NANDN U9985 ( .A(n9451), .B(n9450), .Z(n9452) );
  AND U9986 ( .A(n9453), .B(n9452), .Z(n9508) );
  NAND U9987 ( .A(n9455), .B(n9454), .Z(n9459) );
  NAND U9988 ( .A(n9457), .B(n9456), .Z(n9458) );
  AND U9989 ( .A(n9459), .B(n9458), .Z(n9507) );
  NANDN U9990 ( .A(n9461), .B(n9460), .Z(n9465) );
  NANDN U9991 ( .A(n9463), .B(n9462), .Z(n9464) );
  NAND U9992 ( .A(n9465), .B(n9464), .Z(n9506) );
  XOR U9993 ( .A(n9507), .B(n9506), .Z(n9509) );
  XNOR U9994 ( .A(n9508), .B(n9509), .Z(n9488) );
  XOR U9995 ( .A(n9489), .B(n9488), .Z(n9491) );
  XNOR U9996 ( .A(n9490), .B(n9491), .Z(n9482) );
  XNOR U9997 ( .A(n9483), .B(n9482), .Z(n9484) );
  XNOR U9998 ( .A(n9485), .B(n9484), .Z(n9755) );
  XNOR U9999 ( .A(n9756), .B(n9755), .Z(n9757) );
  XNOR U10000 ( .A(n9758), .B(n9757), .Z(n9476) );
  XNOR U10001 ( .A(n9477), .B(n9476), .Z(n9478) );
  XNOR U10002 ( .A(n9479), .B(n9478), .Z(n9471) );
  XNOR U10003 ( .A(sreg[127]), .B(n9471), .Z(n9473) );
  NANDN U10004 ( .A(sreg[126]), .B(n9466), .Z(n9470) );
  NAND U10005 ( .A(n9468), .B(n9467), .Z(n9469) );
  NAND U10006 ( .A(n9470), .B(n9469), .Z(n9472) );
  XNOR U10007 ( .A(n9473), .B(n9472), .Z(c[127]) );
  NANDN U10008 ( .A(sreg[127]), .B(n9471), .Z(n9475) );
  NAND U10009 ( .A(n9473), .B(n9472), .Z(n9474) );
  NAND U10010 ( .A(n9475), .B(n9474), .Z(n10048) );
  XNOR U10011 ( .A(sreg[128]), .B(n10048), .Z(n10050) );
  NANDN U10012 ( .A(n9477), .B(n9476), .Z(n9481) );
  NANDN U10013 ( .A(n9479), .B(n9478), .Z(n9480) );
  AND U10014 ( .A(n9481), .B(n9480), .Z(n9764) );
  NANDN U10015 ( .A(n9483), .B(n9482), .Z(n9487) );
  NANDN U10016 ( .A(n9485), .B(n9484), .Z(n9486) );
  AND U10017 ( .A(n9487), .B(n9486), .Z(n10045) );
  NANDN U10018 ( .A(n9489), .B(n9488), .Z(n9493) );
  OR U10019 ( .A(n9491), .B(n9490), .Z(n9492) );
  AND U10020 ( .A(n9493), .B(n9492), .Z(n10043) );
  NANDN U10021 ( .A(n9495), .B(n9494), .Z(n9499) );
  NAND U10022 ( .A(n9497), .B(n9496), .Z(n9498) );
  AND U10023 ( .A(n9499), .B(n9498), .Z(n9770) );
  NANDN U10024 ( .A(n9501), .B(n9500), .Z(n9505) );
  NAND U10025 ( .A(n9503), .B(n9502), .Z(n9504) );
  AND U10026 ( .A(n9505), .B(n9504), .Z(n9805) );
  NANDN U10027 ( .A(n9507), .B(n9506), .Z(n9511) );
  NANDN U10028 ( .A(n9509), .B(n9508), .Z(n9510) );
  AND U10029 ( .A(n9511), .B(n9510), .Z(n9804) );
  NANDN U10030 ( .A(n9513), .B(n9512), .Z(n9517) );
  NAND U10031 ( .A(n9515), .B(n9514), .Z(n9516) );
  AND U10032 ( .A(n9517), .B(n9516), .Z(n9803) );
  XOR U10033 ( .A(n9804), .B(n9803), .Z(n9806) );
  XNOR U10034 ( .A(n9805), .B(n9806), .Z(n9767) );
  NANDN U10035 ( .A(n9519), .B(n9518), .Z(n9523) );
  NANDN U10036 ( .A(n9521), .B(n9520), .Z(n9522) );
  AND U10037 ( .A(n9523), .B(n9522), .Z(n9775) );
  NANDN U10038 ( .A(n9525), .B(n9524), .Z(n9529) );
  NANDN U10039 ( .A(n9527), .B(n9526), .Z(n9528) );
  AND U10040 ( .A(n9529), .B(n9528), .Z(n10025) );
  NANDN U10041 ( .A(n9531), .B(n9530), .Z(n9535) );
  NANDN U10042 ( .A(n9533), .B(n9532), .Z(n9534) );
  AND U10043 ( .A(n9535), .B(n9534), .Z(n10024) );
  XNOR U10044 ( .A(n10025), .B(n10024), .Z(n10027) );
  NANDN U10045 ( .A(n9537), .B(n9536), .Z(n9541) );
  OR U10046 ( .A(n9539), .B(n9538), .Z(n9540) );
  AND U10047 ( .A(n9541), .B(n9540), .Z(n9810) );
  NANDN U10048 ( .A(n32996), .B(n9542), .Z(n9544) );
  XOR U10049 ( .A(b[21]), .B(a[44]), .Z(n9909) );
  NANDN U10050 ( .A(n33271), .B(n9909), .Z(n9543) );
  AND U10051 ( .A(n9544), .B(n9543), .Z(n9927) );
  NANDN U10052 ( .A(n9545), .B(n35654), .Z(n9547) );
  XOR U10053 ( .A(b[33]), .B(a[32]), .Z(n9882) );
  NANDN U10054 ( .A(n35456), .B(n9882), .Z(n9546) );
  AND U10055 ( .A(n9547), .B(n9546), .Z(n9925) );
  NANDN U10056 ( .A(n32483), .B(n9548), .Z(n9550) );
  XOR U10057 ( .A(b[19]), .B(a[46]), .Z(n9915) );
  NANDN U10058 ( .A(n32823), .B(n9915), .Z(n9549) );
  NAND U10059 ( .A(n9550), .B(n9549), .Z(n9924) );
  XNOR U10060 ( .A(n9925), .B(n9924), .Z(n9926) );
  XOR U10061 ( .A(n9927), .B(n9926), .Z(n10020) );
  NANDN U10062 ( .A(n33875), .B(n9551), .Z(n9553) );
  XOR U10063 ( .A(b[25]), .B(a[40]), .Z(n9825) );
  NANDN U10064 ( .A(n33994), .B(n9825), .Z(n9552) );
  AND U10065 ( .A(n9553), .B(n9552), .Z(n9876) );
  NANDN U10066 ( .A(n34634), .B(n9554), .Z(n9556) );
  XOR U10067 ( .A(b[29]), .B(a[36]), .Z(n9933) );
  NANDN U10068 ( .A(n34722), .B(n9933), .Z(n9555) );
  AND U10069 ( .A(n9556), .B(n9555), .Z(n9874) );
  NANDN U10070 ( .A(n34223), .B(n9557), .Z(n9559) );
  XOR U10071 ( .A(b[27]), .B(a[38]), .Z(n9930) );
  NANDN U10072 ( .A(n34458), .B(n9930), .Z(n9558) );
  NAND U10073 ( .A(n9559), .B(n9558), .Z(n9873) );
  XNOR U10074 ( .A(n9874), .B(n9873), .Z(n9875) );
  XOR U10075 ( .A(n9876), .B(n9875), .Z(n10018) );
  NANDN U10076 ( .A(n33866), .B(n9560), .Z(n9562) );
  XOR U10077 ( .A(b[23]), .B(a[42]), .Z(n9912) );
  NANDN U10078 ( .A(n33644), .B(n9912), .Z(n9561) );
  AND U10079 ( .A(n9562), .B(n9561), .Z(n10019) );
  XNOR U10080 ( .A(n10018), .B(n10019), .Z(n10021) );
  NANDN U10081 ( .A(n9564), .B(n9563), .Z(n9568) );
  OR U10082 ( .A(n9566), .B(n9565), .Z(n9567) );
  AND U10083 ( .A(n9568), .B(n9567), .Z(n9814) );
  NANDN U10084 ( .A(n9570), .B(n9569), .Z(n9574) );
  OR U10085 ( .A(n9572), .B(n9571), .Z(n9573) );
  NAND U10086 ( .A(n9574), .B(n9573), .Z(n9813) );
  XNOR U10087 ( .A(n9814), .B(n9813), .Z(n9815) );
  XOR U10088 ( .A(n9816), .B(n9815), .Z(n9809) );
  XNOR U10089 ( .A(n9810), .B(n9809), .Z(n9812) );
  NANDN U10090 ( .A(n210), .B(n9575), .Z(n9577) );
  XOR U10091 ( .A(b[9]), .B(a[56]), .Z(n9997) );
  NANDN U10092 ( .A(n30267), .B(n9997), .Z(n9576) );
  AND U10093 ( .A(n9577), .B(n9576), .Z(n9951) );
  NANDN U10094 ( .A(n37705), .B(n9578), .Z(n9580) );
  XOR U10095 ( .A(b[53]), .B(a[12]), .Z(n9837) );
  NANDN U10096 ( .A(n37778), .B(n9837), .Z(n9579) );
  AND U10097 ( .A(n9580), .B(n9579), .Z(n9950) );
  NANDN U10098 ( .A(n34909), .B(n9581), .Z(n9583) );
  XOR U10099 ( .A(b[31]), .B(a[34]), .Z(n9918) );
  NANDN U10100 ( .A(n35145), .B(n9918), .Z(n9582) );
  NAND U10101 ( .A(n9583), .B(n9582), .Z(n9949) );
  XOR U10102 ( .A(n9950), .B(n9949), .Z(n9952) );
  XOR U10103 ( .A(n9951), .B(n9952), .Z(n9904) );
  NANDN U10104 ( .A(n31055), .B(n9584), .Z(n9586) );
  XOR U10105 ( .A(b[13]), .B(a[52]), .Z(n9936) );
  NANDN U10106 ( .A(n31293), .B(n9936), .Z(n9585) );
  AND U10107 ( .A(n9586), .B(n9585), .Z(n9990) );
  NANDN U10108 ( .A(n30482), .B(n9587), .Z(n9589) );
  XOR U10109 ( .A(b[11]), .B(a[54]), .Z(n10009) );
  NANDN U10110 ( .A(n30891), .B(n10009), .Z(n9588) );
  AND U10111 ( .A(n9589), .B(n9588), .Z(n9989) );
  NANDN U10112 ( .A(n212), .B(n9590), .Z(n9592) );
  XOR U10113 ( .A(b[49]), .B(a[16]), .Z(n10000) );
  NANDN U10114 ( .A(n37432), .B(n10000), .Z(n9591) );
  NAND U10115 ( .A(n9592), .B(n9591), .Z(n9988) );
  XOR U10116 ( .A(n9989), .B(n9988), .Z(n9991) );
  XNOR U10117 ( .A(n9990), .B(n9991), .Z(n9903) );
  XNOR U10118 ( .A(n9904), .B(n9903), .Z(n9905) );
  NANDN U10119 ( .A(n9594), .B(n9593), .Z(n9598) );
  OR U10120 ( .A(n9596), .B(n9595), .Z(n9597) );
  NAND U10121 ( .A(n9598), .B(n9597), .Z(n9906) );
  XOR U10122 ( .A(n9905), .B(n9906), .Z(n9786) );
  NANDN U10123 ( .A(n9600), .B(n9599), .Z(n9604) );
  NAND U10124 ( .A(n9602), .B(n9601), .Z(n9603) );
  NAND U10125 ( .A(n9604), .B(n9603), .Z(n9785) );
  XOR U10126 ( .A(n9786), .B(n9785), .Z(n9788) );
  NANDN U10127 ( .A(n9606), .B(n9605), .Z(n9610) );
  OR U10128 ( .A(n9608), .B(n9607), .Z(n9609) );
  AND U10129 ( .A(n9610), .B(n9609), .Z(n9956) );
  NANDN U10130 ( .A(n38090), .B(n9611), .Z(n9613) );
  XOR U10131 ( .A(b[59]), .B(a[6]), .Z(n9891) );
  NANDN U10132 ( .A(n38130), .B(n9891), .Z(n9612) );
  AND U10133 ( .A(n9613), .B(n9612), .Z(n9863) );
  NANDN U10134 ( .A(n29499), .B(n9614), .Z(n9616) );
  XOR U10135 ( .A(b[7]), .B(a[58]), .Z(n9973) );
  NANDN U10136 ( .A(n29735), .B(n9973), .Z(n9615) );
  AND U10137 ( .A(n9616), .B(n9615), .Z(n9862) );
  NANDN U10138 ( .A(n36210), .B(n9617), .Z(n9619) );
  XOR U10139 ( .A(b[39]), .B(a[26]), .Z(n9840) );
  NANDN U10140 ( .A(n36347), .B(n9840), .Z(n9618) );
  NAND U10141 ( .A(n9619), .B(n9618), .Z(n9861) );
  XOR U10142 ( .A(n9862), .B(n9861), .Z(n9864) );
  XNOR U10143 ( .A(n9863), .B(n9864), .Z(n9955) );
  XNOR U10144 ( .A(n9956), .B(n9955), .Z(n9957) );
  NANDN U10145 ( .A(n9621), .B(n9620), .Z(n9625) );
  OR U10146 ( .A(n9623), .B(n9622), .Z(n9624) );
  NAND U10147 ( .A(n9625), .B(n9624), .Z(n9958) );
  XOR U10148 ( .A(n9957), .B(n9958), .Z(n9787) );
  XOR U10149 ( .A(n9788), .B(n9787), .Z(n9811) );
  XOR U10150 ( .A(n9812), .B(n9811), .Z(n10026) );
  XOR U10151 ( .A(n10027), .B(n10026), .Z(n9774) );
  NANDN U10152 ( .A(n9627), .B(n9626), .Z(n9631) );
  NANDN U10153 ( .A(n9629), .B(n9628), .Z(n9630) );
  NAND U10154 ( .A(n9631), .B(n9630), .Z(n9773) );
  XOR U10155 ( .A(n9774), .B(n9773), .Z(n9776) );
  XOR U10156 ( .A(n9775), .B(n9776), .Z(n10039) );
  NANDN U10157 ( .A(n9633), .B(n9632), .Z(n9637) );
  NAND U10158 ( .A(n9635), .B(n9634), .Z(n9636) );
  AND U10159 ( .A(n9637), .B(n9636), .Z(n9800) );
  NANDN U10160 ( .A(n9639), .B(n9638), .Z(n9643) );
  NAND U10161 ( .A(n9641), .B(n9640), .Z(n9642) );
  AND U10162 ( .A(n9643), .B(n9642), .Z(n9793) );
  NANDN U10163 ( .A(n9645), .B(n9644), .Z(n9649) );
  OR U10164 ( .A(n9647), .B(n9646), .Z(n9648) );
  AND U10165 ( .A(n9649), .B(n9648), .Z(n9963) );
  NOR U10166 ( .A(n9651), .B(n9650), .Z(n9857) );
  NAND U10167 ( .A(n9942), .B(n9652), .Z(n9655) );
  XNOR U10168 ( .A(b[3]), .B(a[62]), .Z(n9943) );
  NANDN U10169 ( .A(n9943), .B(n9653), .Z(n9654) );
  AND U10170 ( .A(n9655), .B(n9654), .Z(n9855) );
  NAND U10171 ( .A(n35928), .B(n9656), .Z(n9658) );
  XNOR U10172 ( .A(b[35]), .B(a[30]), .Z(n9979) );
  NANDN U10173 ( .A(n9979), .B(n35929), .Z(n9657) );
  NAND U10174 ( .A(n9658), .B(n9657), .Z(n9856) );
  XOR U10175 ( .A(n9855), .B(n9856), .Z(n9858) );
  XOR U10176 ( .A(n9857), .B(n9858), .Z(n9962) );
  NANDN U10177 ( .A(n211), .B(n9659), .Z(n9661) );
  XOR U10178 ( .A(b[47]), .B(a[18]), .Z(n9994) );
  NANDN U10179 ( .A(n37172), .B(n9994), .Z(n9660) );
  AND U10180 ( .A(n9661), .B(n9660), .Z(n10015) );
  NANDN U10181 ( .A(n37526), .B(n9662), .Z(n9664) );
  XOR U10182 ( .A(b[51]), .B(a[14]), .Z(n9834) );
  NANDN U10183 ( .A(n37605), .B(n9834), .Z(n9663) );
  AND U10184 ( .A(n9664), .B(n9663), .Z(n10013) );
  NANDN U10185 ( .A(n31536), .B(n9665), .Z(n9667) );
  XOR U10186 ( .A(b[15]), .B(a[50]), .Z(n9831) );
  NANDN U10187 ( .A(n31925), .B(n9831), .Z(n9666) );
  NAND U10188 ( .A(n9667), .B(n9666), .Z(n10012) );
  XNOR U10189 ( .A(n10013), .B(n10012), .Z(n10014) );
  XNOR U10190 ( .A(n10015), .B(n10014), .Z(n9961) );
  XOR U10191 ( .A(n9962), .B(n9961), .Z(n9964) );
  XOR U10192 ( .A(n9963), .B(n9964), .Z(n9792) );
  NANDN U10193 ( .A(n36742), .B(n9668), .Z(n9670) );
  XOR U10194 ( .A(b[43]), .B(a[22]), .Z(n10003) );
  NANDN U10195 ( .A(n36891), .B(n10003), .Z(n9669) );
  AND U10196 ( .A(n9670), .B(n9669), .Z(n9845) );
  NANDN U10197 ( .A(n36991), .B(n9671), .Z(n9673) );
  XOR U10198 ( .A(b[45]), .B(a[20]), .Z(n10006) );
  NANDN U10199 ( .A(n37083), .B(n10006), .Z(n9672) );
  AND U10200 ( .A(n9673), .B(n9672), .Z(n9844) );
  NANDN U10201 ( .A(n32013), .B(n9674), .Z(n9676) );
  XOR U10202 ( .A(b[17]), .B(a[48]), .Z(n9828) );
  NANDN U10203 ( .A(n32292), .B(n9828), .Z(n9675) );
  NAND U10204 ( .A(n9676), .B(n9675), .Z(n9843) );
  XOR U10205 ( .A(n9844), .B(n9843), .Z(n9846) );
  XOR U10206 ( .A(n9845), .B(n9846), .Z(n9898) );
  NANDN U10207 ( .A(n37857), .B(n9677), .Z(n9679) );
  XOR U10208 ( .A(b[55]), .B(a[10]), .Z(n9976) );
  NANDN U10209 ( .A(n37911), .B(n9976), .Z(n9678) );
  AND U10210 ( .A(n9679), .B(n9678), .Z(n9851) );
  NANDN U10211 ( .A(n37974), .B(n9680), .Z(n9682) );
  XOR U10212 ( .A(b[57]), .B(a[8]), .Z(n9888) );
  NANDN U10213 ( .A(n38031), .B(n9888), .Z(n9681) );
  AND U10214 ( .A(n9682), .B(n9681), .Z(n9850) );
  NANDN U10215 ( .A(n36480), .B(n9683), .Z(n9685) );
  XOR U10216 ( .A(b[41]), .B(a[24]), .Z(n9894) );
  NANDN U10217 ( .A(n36594), .B(n9894), .Z(n9684) );
  NAND U10218 ( .A(n9685), .B(n9684), .Z(n9849) );
  XOR U10219 ( .A(n9850), .B(n9849), .Z(n9852) );
  XNOR U10220 ( .A(n9851), .B(n9852), .Z(n9897) );
  XNOR U10221 ( .A(n9898), .B(n9897), .Z(n9899) );
  NANDN U10222 ( .A(n9687), .B(n9686), .Z(n9691) );
  NANDN U10223 ( .A(n9689), .B(n9688), .Z(n9690) );
  NAND U10224 ( .A(n9691), .B(n9690), .Z(n9900) );
  XNOR U10225 ( .A(n9899), .B(n9900), .Z(n9791) );
  XOR U10226 ( .A(n9792), .B(n9791), .Z(n9794) );
  XOR U10227 ( .A(n9793), .B(n9794), .Z(n9781) );
  NANDN U10228 ( .A(n9693), .B(n9692), .Z(n9697) );
  NAND U10229 ( .A(n9695), .B(n9694), .Z(n9696) );
  AND U10230 ( .A(n9697), .B(n9696), .Z(n9779) );
  NANDN U10231 ( .A(n9699), .B(n9698), .Z(n9703) );
  OR U10232 ( .A(n9701), .B(n9700), .Z(n9702) );
  AND U10233 ( .A(n9703), .B(n9702), .Z(n9968) );
  NANDN U10234 ( .A(n9705), .B(n9704), .Z(n9709) );
  OR U10235 ( .A(n9707), .B(n9706), .Z(n9708) );
  NAND U10236 ( .A(n9709), .B(n9708), .Z(n9967) );
  XNOR U10237 ( .A(n9968), .B(n9967), .Z(n9969) );
  NANDN U10238 ( .A(n9711), .B(n9710), .Z(n9715) );
  NANDN U10239 ( .A(n9713), .B(n9712), .Z(n9714) );
  AND U10240 ( .A(n9715), .B(n9714), .Z(n9822) );
  NAND U10241 ( .A(b[0]), .B(a[64]), .Z(n9716) );
  XNOR U10242 ( .A(b[1]), .B(n9716), .Z(n9718) );
  NANDN U10243 ( .A(b[0]), .B(a[63]), .Z(n9717) );
  NAND U10244 ( .A(n9718), .B(n9717), .Z(n9985) );
  NANDN U10245 ( .A(n38247), .B(n9719), .Z(n9721) );
  XOR U10246 ( .A(b[61]), .B(a[4]), .Z(n9921) );
  NANDN U10247 ( .A(n38248), .B(n9921), .Z(n9720) );
  AND U10248 ( .A(n9721), .B(n9720), .Z(n9983) );
  AND U10249 ( .A(b[63]), .B(a[0]), .Z(n9982) );
  XNOR U10250 ( .A(n9983), .B(n9982), .Z(n9984) );
  XNOR U10251 ( .A(n9985), .B(n9984), .Z(n9819) );
  NANDN U10252 ( .A(n28889), .B(n9722), .Z(n9724) );
  XOR U10253 ( .A(b[5]), .B(a[60]), .Z(n9939) );
  NANDN U10254 ( .A(n29138), .B(n9939), .Z(n9723) );
  AND U10255 ( .A(n9724), .B(n9723), .Z(n9870) );
  NANDN U10256 ( .A(n38278), .B(n9725), .Z(n9727) );
  XOR U10257 ( .A(b[63]), .B(a[2]), .Z(n9879) );
  NANDN U10258 ( .A(n38279), .B(n9879), .Z(n9726) );
  AND U10259 ( .A(n9727), .B(n9726), .Z(n9868) );
  NANDN U10260 ( .A(n35936), .B(n9728), .Z(n9730) );
  XOR U10261 ( .A(b[37]), .B(a[28]), .Z(n9946) );
  NANDN U10262 ( .A(n36047), .B(n9946), .Z(n9729) );
  NAND U10263 ( .A(n9730), .B(n9729), .Z(n9867) );
  XNOR U10264 ( .A(n9868), .B(n9867), .Z(n9869) );
  XOR U10265 ( .A(n9870), .B(n9869), .Z(n9820) );
  XNOR U10266 ( .A(n9819), .B(n9820), .Z(n9821) );
  XOR U10267 ( .A(n9822), .B(n9821), .Z(n9970) );
  XOR U10268 ( .A(n9969), .B(n9970), .Z(n9780) );
  XOR U10269 ( .A(n9779), .B(n9780), .Z(n9782) );
  XOR U10270 ( .A(n9781), .B(n9782), .Z(n9798) );
  NANDN U10271 ( .A(n9732), .B(n9731), .Z(n9736) );
  NANDN U10272 ( .A(n9734), .B(n9733), .Z(n9735) );
  AND U10273 ( .A(n9736), .B(n9735), .Z(n10032) );
  NANDN U10274 ( .A(n9738), .B(n9737), .Z(n9742) );
  NAND U10275 ( .A(n9740), .B(n9739), .Z(n9741) );
  AND U10276 ( .A(n9742), .B(n9741), .Z(n10030) );
  NANDN U10277 ( .A(n9744), .B(n9743), .Z(n9748) );
  NANDN U10278 ( .A(n9746), .B(n9745), .Z(n9747) );
  NAND U10279 ( .A(n9748), .B(n9747), .Z(n10031) );
  XOR U10280 ( .A(n10030), .B(n10031), .Z(n10033) );
  XNOR U10281 ( .A(n10032), .B(n10033), .Z(n9797) );
  XNOR U10282 ( .A(n9798), .B(n9797), .Z(n9799) );
  XOR U10283 ( .A(n9800), .B(n9799), .Z(n10037) );
  NANDN U10284 ( .A(n9750), .B(n9749), .Z(n9754) );
  NANDN U10285 ( .A(n9752), .B(n9751), .Z(n9753) );
  AND U10286 ( .A(n9754), .B(n9753), .Z(n10036) );
  XNOR U10287 ( .A(n10037), .B(n10036), .Z(n10038) );
  XOR U10288 ( .A(n10039), .B(n10038), .Z(n9768) );
  XNOR U10289 ( .A(n9767), .B(n9768), .Z(n9769) );
  XNOR U10290 ( .A(n9770), .B(n9769), .Z(n10042) );
  XNOR U10291 ( .A(n10043), .B(n10042), .Z(n10044) );
  XOR U10292 ( .A(n10045), .B(n10044), .Z(n9762) );
  NANDN U10293 ( .A(n9756), .B(n9755), .Z(n9760) );
  NANDN U10294 ( .A(n9758), .B(n9757), .Z(n9759) );
  NAND U10295 ( .A(n9760), .B(n9759), .Z(n9761) );
  XNOR U10296 ( .A(n9762), .B(n9761), .Z(n9763) );
  XNOR U10297 ( .A(n9764), .B(n9763), .Z(n10049) );
  XNOR U10298 ( .A(n10050), .B(n10049), .Z(c[128]) );
  NANDN U10299 ( .A(n9762), .B(n9761), .Z(n9766) );
  NANDN U10300 ( .A(n9764), .B(n9763), .Z(n9765) );
  AND U10301 ( .A(n9766), .B(n9765), .Z(n10056) );
  NANDN U10302 ( .A(n9768), .B(n9767), .Z(n9772) );
  NANDN U10303 ( .A(n9770), .B(n9769), .Z(n9771) );
  AND U10304 ( .A(n9772), .B(n9771), .Z(n10334) );
  NANDN U10305 ( .A(n9774), .B(n9773), .Z(n9778) );
  OR U10306 ( .A(n9776), .B(n9775), .Z(n9777) );
  AND U10307 ( .A(n9778), .B(n9777), .Z(n10065) );
  NANDN U10308 ( .A(n9780), .B(n9779), .Z(n9784) );
  OR U10309 ( .A(n9782), .B(n9781), .Z(n9783) );
  AND U10310 ( .A(n9784), .B(n9783), .Z(n10317) );
  NAND U10311 ( .A(n9786), .B(n9785), .Z(n9790) );
  NAND U10312 ( .A(n9788), .B(n9787), .Z(n9789) );
  AND U10313 ( .A(n9790), .B(n9789), .Z(n10316) );
  NANDN U10314 ( .A(n9792), .B(n9791), .Z(n9796) );
  OR U10315 ( .A(n9794), .B(n9793), .Z(n9795) );
  AND U10316 ( .A(n9796), .B(n9795), .Z(n10315) );
  XOR U10317 ( .A(n10316), .B(n10315), .Z(n10318) );
  XOR U10318 ( .A(n10317), .B(n10318), .Z(n10064) );
  NANDN U10319 ( .A(n9798), .B(n9797), .Z(n9802) );
  NAND U10320 ( .A(n9800), .B(n9799), .Z(n9801) );
  NAND U10321 ( .A(n9802), .B(n9801), .Z(n10063) );
  XOR U10322 ( .A(n10064), .B(n10063), .Z(n10066) );
  XNOR U10323 ( .A(n10065), .B(n10066), .Z(n10333) );
  XNOR U10324 ( .A(n10334), .B(n10333), .Z(n10336) );
  NANDN U10325 ( .A(n9804), .B(n9803), .Z(n9808) );
  NANDN U10326 ( .A(n9806), .B(n9805), .Z(n9807) );
  AND U10327 ( .A(n9808), .B(n9807), .Z(n10062) );
  NANDN U10328 ( .A(n9814), .B(n9813), .Z(n9818) );
  NAND U10329 ( .A(n9816), .B(n9815), .Z(n9817) );
  AND U10330 ( .A(n9818), .B(n9817), .Z(n10305) );
  NANDN U10331 ( .A(n9820), .B(n9819), .Z(n9824) );
  NANDN U10332 ( .A(n9822), .B(n9821), .Z(n9823) );
  AND U10333 ( .A(n9824), .B(n9823), .Z(n10304) );
  NANDN U10334 ( .A(n33875), .B(n9825), .Z(n9827) );
  XOR U10335 ( .A(b[25]), .B(a[41]), .Z(n10132) );
  NANDN U10336 ( .A(n33994), .B(n10132), .Z(n9826) );
  AND U10337 ( .A(n9827), .B(n9826), .Z(n10257) );
  NANDN U10338 ( .A(n32013), .B(n9828), .Z(n9830) );
  XOR U10339 ( .A(b[17]), .B(a[49]), .Z(n10135) );
  NANDN U10340 ( .A(n32292), .B(n10135), .Z(n9829) );
  AND U10341 ( .A(n9830), .B(n9829), .Z(n10256) );
  NANDN U10342 ( .A(n31536), .B(n9831), .Z(n9833) );
  XOR U10343 ( .A(b[15]), .B(a[51]), .Z(n10138) );
  NANDN U10344 ( .A(n31925), .B(n10138), .Z(n9832) );
  NAND U10345 ( .A(n9833), .B(n9832), .Z(n10255) );
  XOR U10346 ( .A(n10256), .B(n10255), .Z(n10258) );
  XOR U10347 ( .A(n10257), .B(n10258), .Z(n10229) );
  NANDN U10348 ( .A(n37526), .B(n9834), .Z(n9836) );
  XOR U10349 ( .A(b[51]), .B(a[15]), .Z(n10141) );
  NANDN U10350 ( .A(n37605), .B(n10141), .Z(n9835) );
  AND U10351 ( .A(n9836), .B(n9835), .Z(n10281) );
  NANDN U10352 ( .A(n37705), .B(n9837), .Z(n9839) );
  XOR U10353 ( .A(b[53]), .B(a[13]), .Z(n10144) );
  NANDN U10354 ( .A(n37778), .B(n10144), .Z(n9838) );
  AND U10355 ( .A(n9839), .B(n9838), .Z(n10280) );
  NANDN U10356 ( .A(n36210), .B(n9840), .Z(n9842) );
  XOR U10357 ( .A(b[39]), .B(a[27]), .Z(n10147) );
  NANDN U10358 ( .A(n36347), .B(n10147), .Z(n9841) );
  NAND U10359 ( .A(n9842), .B(n9841), .Z(n10279) );
  XOR U10360 ( .A(n10280), .B(n10279), .Z(n10282) );
  XNOR U10361 ( .A(n10281), .B(n10282), .Z(n10228) );
  XNOR U10362 ( .A(n10229), .B(n10228), .Z(n10231) );
  NANDN U10363 ( .A(n9844), .B(n9843), .Z(n9848) );
  OR U10364 ( .A(n9846), .B(n9845), .Z(n9847) );
  AND U10365 ( .A(n9848), .B(n9847), .Z(n10230) );
  XOR U10366 ( .A(n10231), .B(n10230), .Z(n10123) );
  NANDN U10367 ( .A(n9850), .B(n9849), .Z(n9854) );
  OR U10368 ( .A(n9852), .B(n9851), .Z(n9853) );
  AND U10369 ( .A(n9854), .B(n9853), .Z(n10121) );
  NANDN U10370 ( .A(n9856), .B(n9855), .Z(n9860) );
  OR U10371 ( .A(n9858), .B(n9857), .Z(n9859) );
  AND U10372 ( .A(n9860), .B(n9859), .Z(n10120) );
  XNOR U10373 ( .A(n10121), .B(n10120), .Z(n10122) );
  XNOR U10374 ( .A(n10123), .B(n10122), .Z(n10303) );
  XOR U10375 ( .A(n10304), .B(n10303), .Z(n10306) );
  XOR U10376 ( .A(n10305), .B(n10306), .Z(n10292) );
  NANDN U10377 ( .A(n9862), .B(n9861), .Z(n9866) );
  OR U10378 ( .A(n9864), .B(n9863), .Z(n9865) );
  AND U10379 ( .A(n9866), .B(n9865), .Z(n10187) );
  NANDN U10380 ( .A(n9868), .B(n9867), .Z(n9872) );
  NANDN U10381 ( .A(n9870), .B(n9869), .Z(n9871) );
  NAND U10382 ( .A(n9872), .B(n9871), .Z(n10186) );
  XNOR U10383 ( .A(n10187), .B(n10186), .Z(n10189) );
  NANDN U10384 ( .A(n9874), .B(n9873), .Z(n9878) );
  NANDN U10385 ( .A(n9876), .B(n9875), .Z(n9877) );
  AND U10386 ( .A(n9878), .B(n9877), .Z(n10129) );
  NANDN U10387 ( .A(n38278), .B(n9879), .Z(n9881) );
  XOR U10388 ( .A(b[63]), .B(a[3]), .Z(n10210) );
  NANDN U10389 ( .A(n38279), .B(n10210), .Z(n9880) );
  AND U10390 ( .A(n9881), .B(n9880), .Z(n10163) );
  NANDN U10391 ( .A(n35260), .B(n9882), .Z(n9884) );
  XOR U10392 ( .A(b[33]), .B(a[33]), .Z(n10213) );
  NANDN U10393 ( .A(n35456), .B(n10213), .Z(n9883) );
  NAND U10394 ( .A(n9884), .B(n9883), .Z(n10162) );
  XNOR U10395 ( .A(n10163), .B(n10162), .Z(n10164) );
  NAND U10396 ( .A(b[0]), .B(a[65]), .Z(n9885) );
  XNOR U10397 ( .A(b[1]), .B(n9885), .Z(n9887) );
  NANDN U10398 ( .A(b[0]), .B(a[64]), .Z(n9886) );
  NAND U10399 ( .A(n9887), .B(n9886), .Z(n10165) );
  XNOR U10400 ( .A(n10164), .B(n10165), .Z(n10126) );
  NANDN U10401 ( .A(n37974), .B(n9888), .Z(n9890) );
  XOR U10402 ( .A(b[57]), .B(a[9]), .Z(n10219) );
  NANDN U10403 ( .A(n38031), .B(n10219), .Z(n9889) );
  AND U10404 ( .A(n9890), .B(n9889), .Z(n10195) );
  NANDN U10405 ( .A(n38090), .B(n9891), .Z(n9893) );
  XOR U10406 ( .A(b[59]), .B(a[7]), .Z(n10222) );
  NANDN U10407 ( .A(n38130), .B(n10222), .Z(n9892) );
  AND U10408 ( .A(n9893), .B(n9892), .Z(n10193) );
  NANDN U10409 ( .A(n36480), .B(n9894), .Z(n9896) );
  XOR U10410 ( .A(b[41]), .B(a[25]), .Z(n10225) );
  NANDN U10411 ( .A(n36594), .B(n10225), .Z(n9895) );
  NAND U10412 ( .A(n9896), .B(n9895), .Z(n10192) );
  XNOR U10413 ( .A(n10193), .B(n10192), .Z(n10194) );
  XOR U10414 ( .A(n10195), .B(n10194), .Z(n10127) );
  XNOR U10415 ( .A(n10126), .B(n10127), .Z(n10128) );
  XNOR U10416 ( .A(n10129), .B(n10128), .Z(n10188) );
  XOR U10417 ( .A(n10189), .B(n10188), .Z(n10169) );
  NANDN U10418 ( .A(n9898), .B(n9897), .Z(n9902) );
  NANDN U10419 ( .A(n9900), .B(n9899), .Z(n9901) );
  NAND U10420 ( .A(n9902), .B(n9901), .Z(n10168) );
  XNOR U10421 ( .A(n10169), .B(n10168), .Z(n10170) );
  NANDN U10422 ( .A(n9904), .B(n9903), .Z(n9908) );
  NANDN U10423 ( .A(n9906), .B(n9905), .Z(n9907) );
  AND U10424 ( .A(n9908), .B(n9907), .Z(n10288) );
  NANDN U10425 ( .A(n32996), .B(n9909), .Z(n9911) );
  XOR U10426 ( .A(b[21]), .B(a[45]), .Z(n10240) );
  NANDN U10427 ( .A(n33271), .B(n10240), .Z(n9910) );
  AND U10428 ( .A(n9911), .B(n9910), .Z(n10206) );
  NANDN U10429 ( .A(n33866), .B(n9912), .Z(n9914) );
  XOR U10430 ( .A(b[23]), .B(a[43]), .Z(n10243) );
  NANDN U10431 ( .A(n33644), .B(n10243), .Z(n9913) );
  AND U10432 ( .A(n9914), .B(n9913), .Z(n10205) );
  NANDN U10433 ( .A(n32483), .B(n9915), .Z(n9917) );
  XOR U10434 ( .A(b[19]), .B(a[47]), .Z(n10246) );
  NANDN U10435 ( .A(n32823), .B(n10246), .Z(n9916) );
  NAND U10436 ( .A(n9917), .B(n9916), .Z(n10204) );
  XOR U10437 ( .A(n10205), .B(n10204), .Z(n10207) );
  XOR U10438 ( .A(n10206), .B(n10207), .Z(n10091) );
  NANDN U10439 ( .A(n34909), .B(n9918), .Z(n9920) );
  XOR U10440 ( .A(b[31]), .B(a[35]), .Z(n10249) );
  NANDN U10441 ( .A(n35145), .B(n10249), .Z(n9919) );
  AND U10442 ( .A(n9920), .B(n9919), .Z(n10080) );
  NANDN U10443 ( .A(n38247), .B(n9921), .Z(n9923) );
  XOR U10444 ( .A(b[61]), .B(a[5]), .Z(n10252) );
  NANDN U10445 ( .A(n38248), .B(n10252), .Z(n9922) );
  AND U10446 ( .A(n9923), .B(n9922), .Z(n10079) );
  AND U10447 ( .A(b[63]), .B(a[1]), .Z(n10078) );
  XOR U10448 ( .A(n10079), .B(n10078), .Z(n10081) );
  XNOR U10449 ( .A(n10080), .B(n10081), .Z(n10090) );
  XNOR U10450 ( .A(n10091), .B(n10090), .Z(n10092) );
  NANDN U10451 ( .A(n9925), .B(n9924), .Z(n9929) );
  NANDN U10452 ( .A(n9927), .B(n9926), .Z(n9928) );
  NAND U10453 ( .A(n9929), .B(n9928), .Z(n10093) );
  XNOR U10454 ( .A(n10092), .B(n10093), .Z(n10285) );
  NANDN U10455 ( .A(n34223), .B(n9930), .Z(n9932) );
  XOR U10456 ( .A(b[27]), .B(a[39]), .Z(n10261) );
  NANDN U10457 ( .A(n34458), .B(n10261), .Z(n9931) );
  AND U10458 ( .A(n9932), .B(n9931), .Z(n10152) );
  NANDN U10459 ( .A(n34634), .B(n9933), .Z(n9935) );
  XOR U10460 ( .A(b[29]), .B(a[37]), .Z(n10264) );
  NANDN U10461 ( .A(n34722), .B(n10264), .Z(n9934) );
  AND U10462 ( .A(n9935), .B(n9934), .Z(n10151) );
  NANDN U10463 ( .A(n31055), .B(n9936), .Z(n9938) );
  XOR U10464 ( .A(b[13]), .B(a[53]), .Z(n10267) );
  NANDN U10465 ( .A(n31293), .B(n10267), .Z(n9937) );
  NAND U10466 ( .A(n9938), .B(n9937), .Z(n10150) );
  XOR U10467 ( .A(n10151), .B(n10150), .Z(n10153) );
  XOR U10468 ( .A(n10152), .B(n10153), .Z(n10181) );
  NANDN U10469 ( .A(n28889), .B(n9939), .Z(n9941) );
  XOR U10470 ( .A(b[5]), .B(a[61]), .Z(n10270) );
  NANDN U10471 ( .A(n29138), .B(n10270), .Z(n9940) );
  AND U10472 ( .A(n9941), .B(n9940), .Z(n10200) );
  NANDN U10473 ( .A(n9943), .B(n9942), .Z(n9945) );
  XOR U10474 ( .A(b[3]), .B(a[63]), .Z(n10273) );
  NANDN U10475 ( .A(n28941), .B(n10273), .Z(n9944) );
  AND U10476 ( .A(n9945), .B(n9944), .Z(n10199) );
  NANDN U10477 ( .A(n35936), .B(n9946), .Z(n9948) );
  XOR U10478 ( .A(b[37]), .B(a[29]), .Z(n10276) );
  NANDN U10479 ( .A(n36047), .B(n10276), .Z(n9947) );
  NAND U10480 ( .A(n9948), .B(n9947), .Z(n10198) );
  XOR U10481 ( .A(n10199), .B(n10198), .Z(n10201) );
  XNOR U10482 ( .A(n10200), .B(n10201), .Z(n10180) );
  XNOR U10483 ( .A(n10181), .B(n10180), .Z(n10182) );
  NANDN U10484 ( .A(n9950), .B(n9949), .Z(n9954) );
  OR U10485 ( .A(n9952), .B(n9951), .Z(n9953) );
  NAND U10486 ( .A(n9954), .B(n9953), .Z(n10183) );
  XOR U10487 ( .A(n10182), .B(n10183), .Z(n10286) );
  XNOR U10488 ( .A(n10285), .B(n10286), .Z(n10287) );
  XOR U10489 ( .A(n10288), .B(n10287), .Z(n10171) );
  XNOR U10490 ( .A(n10170), .B(n10171), .Z(n10291) );
  XOR U10491 ( .A(n10292), .B(n10291), .Z(n10294) );
  XOR U10492 ( .A(n10293), .B(n10294), .Z(n10323) );
  NANDN U10493 ( .A(n9956), .B(n9955), .Z(n9960) );
  NANDN U10494 ( .A(n9958), .B(n9957), .Z(n9959) );
  AND U10495 ( .A(n9960), .B(n9959), .Z(n10300) );
  NANDN U10496 ( .A(n9962), .B(n9961), .Z(n9966) );
  OR U10497 ( .A(n9964), .B(n9963), .Z(n9965) );
  AND U10498 ( .A(n9966), .B(n9965), .Z(n10297) );
  NANDN U10499 ( .A(n9968), .B(n9967), .Z(n9972) );
  NANDN U10500 ( .A(n9970), .B(n9969), .Z(n9971) );
  NAND U10501 ( .A(n9972), .B(n9971), .Z(n10298) );
  XNOR U10502 ( .A(n10297), .B(n10298), .Z(n10299) );
  XOR U10503 ( .A(n10300), .B(n10299), .Z(n10321) );
  NANDN U10504 ( .A(n29499), .B(n9973), .Z(n9975) );
  XOR U10505 ( .A(b[7]), .B(a[59]), .Z(n10069) );
  NANDN U10506 ( .A(n29735), .B(n10069), .Z(n9974) );
  AND U10507 ( .A(n9975), .B(n9974), .Z(n10158) );
  NANDN U10508 ( .A(n37857), .B(n9976), .Z(n9978) );
  XOR U10509 ( .A(b[55]), .B(a[11]), .Z(n10072) );
  NANDN U10510 ( .A(n37911), .B(n10072), .Z(n9977) );
  AND U10511 ( .A(n9978), .B(n9977), .Z(n10157) );
  NANDN U10512 ( .A(n9979), .B(n35928), .Z(n9981) );
  XOR U10513 ( .A(b[35]), .B(a[31]), .Z(n10075) );
  NANDN U10514 ( .A(n35801), .B(n10075), .Z(n9980) );
  NAND U10515 ( .A(n9981), .B(n9980), .Z(n10156) );
  XOR U10516 ( .A(n10157), .B(n10156), .Z(n10159) );
  XOR U10517 ( .A(n10158), .B(n10159), .Z(n10175) );
  NANDN U10518 ( .A(n9983), .B(n9982), .Z(n9987) );
  NANDN U10519 ( .A(n9985), .B(n9984), .Z(n9986) );
  AND U10520 ( .A(n9987), .B(n9986), .Z(n10174) );
  XNOR U10521 ( .A(n10175), .B(n10174), .Z(n10177) );
  NANDN U10522 ( .A(n9989), .B(n9988), .Z(n9993) );
  OR U10523 ( .A(n9991), .B(n9990), .Z(n9992) );
  AND U10524 ( .A(n9993), .B(n9992), .Z(n10176) );
  XOR U10525 ( .A(n10177), .B(n10176), .Z(n10311) );
  NANDN U10526 ( .A(n211), .B(n9994), .Z(n9996) );
  XOR U10527 ( .A(b[47]), .B(a[19]), .Z(n10096) );
  NANDN U10528 ( .A(n37172), .B(n10096), .Z(n9995) );
  AND U10529 ( .A(n9996), .B(n9995), .Z(n10086) );
  NANDN U10530 ( .A(n210), .B(n9997), .Z(n9999) );
  XOR U10531 ( .A(b[9]), .B(a[57]), .Z(n10099) );
  NANDN U10532 ( .A(n30267), .B(n10099), .Z(n9998) );
  AND U10533 ( .A(n9999), .B(n9998), .Z(n10085) );
  NANDN U10534 ( .A(n212), .B(n10000), .Z(n10002) );
  XOR U10535 ( .A(b[49]), .B(a[17]), .Z(n10102) );
  NANDN U10536 ( .A(n37432), .B(n10102), .Z(n10001) );
  NAND U10537 ( .A(n10002), .B(n10001), .Z(n10084) );
  XOR U10538 ( .A(n10085), .B(n10084), .Z(n10087) );
  XOR U10539 ( .A(n10086), .B(n10087), .Z(n10235) );
  NANDN U10540 ( .A(n36742), .B(n10003), .Z(n10005) );
  XOR U10541 ( .A(b[43]), .B(a[23]), .Z(n10105) );
  NANDN U10542 ( .A(n36891), .B(n10105), .Z(n10004) );
  AND U10543 ( .A(n10005), .B(n10004), .Z(n10116) );
  NANDN U10544 ( .A(n36991), .B(n10006), .Z(n10008) );
  XOR U10545 ( .A(b[45]), .B(a[21]), .Z(n10108) );
  NANDN U10546 ( .A(n37083), .B(n10108), .Z(n10007) );
  AND U10547 ( .A(n10008), .B(n10007), .Z(n10115) );
  NANDN U10548 ( .A(n30482), .B(n10009), .Z(n10011) );
  XOR U10549 ( .A(b[11]), .B(a[55]), .Z(n10111) );
  NANDN U10550 ( .A(n30891), .B(n10111), .Z(n10010) );
  NAND U10551 ( .A(n10011), .B(n10010), .Z(n10114) );
  XOR U10552 ( .A(n10115), .B(n10114), .Z(n10117) );
  XNOR U10553 ( .A(n10116), .B(n10117), .Z(n10234) );
  XNOR U10554 ( .A(n10235), .B(n10234), .Z(n10237) );
  NANDN U10555 ( .A(n10013), .B(n10012), .Z(n10017) );
  NANDN U10556 ( .A(n10015), .B(n10014), .Z(n10016) );
  AND U10557 ( .A(n10017), .B(n10016), .Z(n10236) );
  XOR U10558 ( .A(n10237), .B(n10236), .Z(n10310) );
  NAND U10559 ( .A(n10019), .B(n10018), .Z(n10023) );
  NANDN U10560 ( .A(n10021), .B(n10020), .Z(n10022) );
  AND U10561 ( .A(n10023), .B(n10022), .Z(n10309) );
  XOR U10562 ( .A(n10310), .B(n10309), .Z(n10312) );
  XOR U10563 ( .A(n10311), .B(n10312), .Z(n10322) );
  XOR U10564 ( .A(n10321), .B(n10322), .Z(n10324) );
  XNOR U10565 ( .A(n10323), .B(n10324), .Z(n10329) );
  NANDN U10566 ( .A(n10025), .B(n10024), .Z(n10029) );
  NAND U10567 ( .A(n10027), .B(n10026), .Z(n10028) );
  AND U10568 ( .A(n10029), .B(n10028), .Z(n10327) );
  NANDN U10569 ( .A(n10031), .B(n10030), .Z(n10035) );
  OR U10570 ( .A(n10033), .B(n10032), .Z(n10034) );
  NAND U10571 ( .A(n10035), .B(n10034), .Z(n10328) );
  XOR U10572 ( .A(n10327), .B(n10328), .Z(n10330) );
  XOR U10573 ( .A(n10329), .B(n10330), .Z(n10059) );
  NANDN U10574 ( .A(n10037), .B(n10036), .Z(n10041) );
  NANDN U10575 ( .A(n10039), .B(n10038), .Z(n10040) );
  NAND U10576 ( .A(n10041), .B(n10040), .Z(n10060) );
  XOR U10577 ( .A(n10059), .B(n10060), .Z(n10061) );
  XNOR U10578 ( .A(n10062), .B(n10061), .Z(n10335) );
  XOR U10579 ( .A(n10336), .B(n10335), .Z(n10054) );
  NANDN U10580 ( .A(n10043), .B(n10042), .Z(n10047) );
  NAND U10581 ( .A(n10045), .B(n10044), .Z(n10046) );
  AND U10582 ( .A(n10047), .B(n10046), .Z(n10053) );
  XNOR U10583 ( .A(n10054), .B(n10053), .Z(n10055) );
  XNOR U10584 ( .A(n10056), .B(n10055), .Z(n10339) );
  XNOR U10585 ( .A(sreg[129]), .B(n10339), .Z(n10341) );
  NANDN U10586 ( .A(sreg[128]), .B(n10048), .Z(n10052) );
  NAND U10587 ( .A(n10050), .B(n10049), .Z(n10051) );
  NAND U10588 ( .A(n10052), .B(n10051), .Z(n10340) );
  XNOR U10589 ( .A(n10341), .B(n10340), .Z(c[129]) );
  NANDN U10590 ( .A(n10054), .B(n10053), .Z(n10058) );
  NANDN U10591 ( .A(n10056), .B(n10055), .Z(n10057) );
  AND U10592 ( .A(n10058), .B(n10057), .Z(n10347) );
  NANDN U10593 ( .A(n10064), .B(n10063), .Z(n10068) );
  OR U10594 ( .A(n10066), .B(n10065), .Z(n10067) );
  AND U10595 ( .A(n10068), .B(n10067), .Z(n10626) );
  NANDN U10596 ( .A(n29499), .B(n10069), .Z(n10071) );
  XOR U10597 ( .A(b[7]), .B(a[60]), .Z(n10464) );
  NANDN U10598 ( .A(n29735), .B(n10464), .Z(n10070) );
  AND U10599 ( .A(n10071), .B(n10070), .Z(n10424) );
  NANDN U10600 ( .A(n37857), .B(n10072), .Z(n10074) );
  XOR U10601 ( .A(b[55]), .B(a[12]), .Z(n10467) );
  NANDN U10602 ( .A(n37911), .B(n10467), .Z(n10073) );
  AND U10603 ( .A(n10074), .B(n10073), .Z(n10423) );
  NANDN U10604 ( .A(n35611), .B(n10075), .Z(n10077) );
  XOR U10605 ( .A(b[35]), .B(a[32]), .Z(n10470) );
  NANDN U10606 ( .A(n35801), .B(n10470), .Z(n10076) );
  NAND U10607 ( .A(n10077), .B(n10076), .Z(n10422) );
  XOR U10608 ( .A(n10423), .B(n10422), .Z(n10425) );
  XOR U10609 ( .A(n10424), .B(n10425), .Z(n10486) );
  NANDN U10610 ( .A(n10079), .B(n10078), .Z(n10083) );
  OR U10611 ( .A(n10081), .B(n10080), .Z(n10082) );
  AND U10612 ( .A(n10083), .B(n10082), .Z(n10485) );
  XNOR U10613 ( .A(n10486), .B(n10485), .Z(n10487) );
  NANDN U10614 ( .A(n10085), .B(n10084), .Z(n10089) );
  OR U10615 ( .A(n10087), .B(n10086), .Z(n10088) );
  NAND U10616 ( .A(n10089), .B(n10088), .Z(n10488) );
  XNOR U10617 ( .A(n10487), .B(n10488), .Z(n10359) );
  NANDN U10618 ( .A(n10091), .B(n10090), .Z(n10095) );
  NANDN U10619 ( .A(n10093), .B(n10092), .Z(n10094) );
  AND U10620 ( .A(n10095), .B(n10094), .Z(n10357) );
  NANDN U10621 ( .A(n211), .B(n10096), .Z(n10098) );
  XOR U10622 ( .A(b[47]), .B(a[20]), .Z(n10440) );
  NANDN U10623 ( .A(n37172), .B(n10440), .Z(n10097) );
  AND U10624 ( .A(n10098), .B(n10097), .Z(n10481) );
  NANDN U10625 ( .A(n210), .B(n10099), .Z(n10101) );
  XOR U10626 ( .A(b[9]), .B(a[58]), .Z(n10443) );
  NANDN U10627 ( .A(n30267), .B(n10443), .Z(n10100) );
  AND U10628 ( .A(n10101), .B(n10100), .Z(n10480) );
  NANDN U10629 ( .A(n212), .B(n10102), .Z(n10104) );
  XOR U10630 ( .A(b[49]), .B(a[18]), .Z(n10446) );
  NANDN U10631 ( .A(n37432), .B(n10446), .Z(n10103) );
  NAND U10632 ( .A(n10104), .B(n10103), .Z(n10479) );
  XOR U10633 ( .A(n10480), .B(n10479), .Z(n10482) );
  XOR U10634 ( .A(n10481), .B(n10482), .Z(n10546) );
  NANDN U10635 ( .A(n36742), .B(n10105), .Z(n10107) );
  XOR U10636 ( .A(b[43]), .B(a[24]), .Z(n10449) );
  NANDN U10637 ( .A(n36891), .B(n10449), .Z(n10106) );
  AND U10638 ( .A(n10107), .B(n10106), .Z(n10460) );
  NANDN U10639 ( .A(n36991), .B(n10108), .Z(n10110) );
  XOR U10640 ( .A(b[45]), .B(a[22]), .Z(n10452) );
  NANDN U10641 ( .A(n37083), .B(n10452), .Z(n10109) );
  AND U10642 ( .A(n10110), .B(n10109), .Z(n10459) );
  NANDN U10643 ( .A(n30482), .B(n10111), .Z(n10113) );
  XOR U10644 ( .A(b[11]), .B(a[56]), .Z(n10455) );
  NANDN U10645 ( .A(n30891), .B(n10455), .Z(n10112) );
  NAND U10646 ( .A(n10113), .B(n10112), .Z(n10458) );
  XOR U10647 ( .A(n10459), .B(n10458), .Z(n10461) );
  XNOR U10648 ( .A(n10460), .B(n10461), .Z(n10545) );
  XNOR U10649 ( .A(n10546), .B(n10545), .Z(n10547) );
  NANDN U10650 ( .A(n10115), .B(n10114), .Z(n10119) );
  OR U10651 ( .A(n10117), .B(n10116), .Z(n10118) );
  NAND U10652 ( .A(n10119), .B(n10118), .Z(n10548) );
  XNOR U10653 ( .A(n10547), .B(n10548), .Z(n10356) );
  XNOR U10654 ( .A(n10357), .B(n10356), .Z(n10358) );
  XOR U10655 ( .A(n10359), .B(n10358), .Z(n10369) );
  NANDN U10656 ( .A(n10121), .B(n10120), .Z(n10125) );
  NANDN U10657 ( .A(n10123), .B(n10122), .Z(n10124) );
  AND U10658 ( .A(n10125), .B(n10124), .Z(n10365) );
  NANDN U10659 ( .A(n10127), .B(n10126), .Z(n10131) );
  NANDN U10660 ( .A(n10129), .B(n10128), .Z(n10130) );
  AND U10661 ( .A(n10131), .B(n10130), .Z(n10363) );
  NANDN U10662 ( .A(n33875), .B(n10132), .Z(n10134) );
  XOR U10663 ( .A(b[25]), .B(a[42]), .Z(n10398) );
  NANDN U10664 ( .A(n33994), .B(n10398), .Z(n10133) );
  AND U10665 ( .A(n10134), .B(n10133), .Z(n10568) );
  NANDN U10666 ( .A(n32013), .B(n10135), .Z(n10137) );
  XOR U10667 ( .A(b[17]), .B(a[50]), .Z(n10401) );
  NANDN U10668 ( .A(n32292), .B(n10401), .Z(n10136) );
  AND U10669 ( .A(n10137), .B(n10136), .Z(n10567) );
  NANDN U10670 ( .A(n31536), .B(n10138), .Z(n10140) );
  XOR U10671 ( .A(b[15]), .B(a[52]), .Z(n10404) );
  NANDN U10672 ( .A(n31925), .B(n10404), .Z(n10139) );
  NAND U10673 ( .A(n10140), .B(n10139), .Z(n10566) );
  XOR U10674 ( .A(n10567), .B(n10566), .Z(n10569) );
  XOR U10675 ( .A(n10568), .B(n10569), .Z(n10540) );
  NANDN U10676 ( .A(n37526), .B(n10141), .Z(n10143) );
  XOR U10677 ( .A(b[51]), .B(a[16]), .Z(n10407) );
  NANDN U10678 ( .A(n37605), .B(n10407), .Z(n10142) );
  AND U10679 ( .A(n10143), .B(n10142), .Z(n10592) );
  NANDN U10680 ( .A(n37705), .B(n10144), .Z(n10146) );
  XOR U10681 ( .A(b[53]), .B(a[14]), .Z(n10410) );
  NANDN U10682 ( .A(n37778), .B(n10410), .Z(n10145) );
  AND U10683 ( .A(n10146), .B(n10145), .Z(n10591) );
  NANDN U10684 ( .A(n36210), .B(n10147), .Z(n10149) );
  XOR U10685 ( .A(b[39]), .B(a[28]), .Z(n10413) );
  NANDN U10686 ( .A(n36347), .B(n10413), .Z(n10148) );
  NAND U10687 ( .A(n10149), .B(n10148), .Z(n10590) );
  XOR U10688 ( .A(n10591), .B(n10590), .Z(n10593) );
  XNOR U10689 ( .A(n10592), .B(n10593), .Z(n10539) );
  XNOR U10690 ( .A(n10540), .B(n10539), .Z(n10542) );
  NANDN U10691 ( .A(n10151), .B(n10150), .Z(n10155) );
  OR U10692 ( .A(n10153), .B(n10152), .Z(n10154) );
  AND U10693 ( .A(n10155), .B(n10154), .Z(n10541) );
  XOR U10694 ( .A(n10542), .B(n10541), .Z(n10389) );
  NANDN U10695 ( .A(n10157), .B(n10156), .Z(n10161) );
  OR U10696 ( .A(n10159), .B(n10158), .Z(n10160) );
  AND U10697 ( .A(n10161), .B(n10160), .Z(n10387) );
  NANDN U10698 ( .A(n10163), .B(n10162), .Z(n10167) );
  NANDN U10699 ( .A(n10165), .B(n10164), .Z(n10166) );
  NAND U10700 ( .A(n10167), .B(n10166), .Z(n10386) );
  XNOR U10701 ( .A(n10387), .B(n10386), .Z(n10388) );
  XNOR U10702 ( .A(n10389), .B(n10388), .Z(n10362) );
  XNOR U10703 ( .A(n10363), .B(n10362), .Z(n10364) );
  XNOR U10704 ( .A(n10365), .B(n10364), .Z(n10368) );
  XNOR U10705 ( .A(n10369), .B(n10368), .Z(n10370) );
  NANDN U10706 ( .A(n10169), .B(n10168), .Z(n10173) );
  NANDN U10707 ( .A(n10171), .B(n10170), .Z(n10172) );
  NAND U10708 ( .A(n10173), .B(n10172), .Z(n10371) );
  XNOR U10709 ( .A(n10370), .B(n10371), .Z(n10608) );
  NANDN U10710 ( .A(n10175), .B(n10174), .Z(n10179) );
  NAND U10711 ( .A(n10177), .B(n10176), .Z(n10178) );
  AND U10712 ( .A(n10179), .B(n10178), .Z(n10352) );
  NANDN U10713 ( .A(n10181), .B(n10180), .Z(n10185) );
  NANDN U10714 ( .A(n10183), .B(n10182), .Z(n10184) );
  AND U10715 ( .A(n10185), .B(n10184), .Z(n10351) );
  NANDN U10716 ( .A(n10187), .B(n10186), .Z(n10191) );
  NAND U10717 ( .A(n10189), .B(n10188), .Z(n10190) );
  AND U10718 ( .A(n10191), .B(n10190), .Z(n10350) );
  XOR U10719 ( .A(n10351), .B(n10350), .Z(n10353) );
  XOR U10720 ( .A(n10352), .B(n10353), .Z(n10377) );
  NANDN U10721 ( .A(n10193), .B(n10192), .Z(n10197) );
  NANDN U10722 ( .A(n10195), .B(n10194), .Z(n10196) );
  AND U10723 ( .A(n10197), .B(n10196), .Z(n10498) );
  NANDN U10724 ( .A(n10199), .B(n10198), .Z(n10203) );
  OR U10725 ( .A(n10201), .B(n10200), .Z(n10202) );
  NAND U10726 ( .A(n10203), .B(n10202), .Z(n10497) );
  XNOR U10727 ( .A(n10498), .B(n10497), .Z(n10500) );
  NANDN U10728 ( .A(n10205), .B(n10204), .Z(n10209) );
  OR U10729 ( .A(n10207), .B(n10206), .Z(n10208) );
  AND U10730 ( .A(n10209), .B(n10208), .Z(n10395) );
  NANDN U10731 ( .A(n38278), .B(n10210), .Z(n10212) );
  XOR U10732 ( .A(b[63]), .B(a[4]), .Z(n10524) );
  NANDN U10733 ( .A(n38279), .B(n10524), .Z(n10211) );
  AND U10734 ( .A(n10212), .B(n10211), .Z(n10429) );
  NANDN U10735 ( .A(n35260), .B(n10213), .Z(n10215) );
  XOR U10736 ( .A(b[33]), .B(a[34]), .Z(n10527) );
  NANDN U10737 ( .A(n35456), .B(n10527), .Z(n10214) );
  NAND U10738 ( .A(n10215), .B(n10214), .Z(n10428) );
  XNOR U10739 ( .A(n10429), .B(n10428), .Z(n10430) );
  NAND U10740 ( .A(b[0]), .B(a[66]), .Z(n10216) );
  XNOR U10741 ( .A(b[1]), .B(n10216), .Z(n10218) );
  NANDN U10742 ( .A(b[0]), .B(a[65]), .Z(n10217) );
  NAND U10743 ( .A(n10218), .B(n10217), .Z(n10431) );
  XNOR U10744 ( .A(n10430), .B(n10431), .Z(n10392) );
  NANDN U10745 ( .A(n37974), .B(n10219), .Z(n10221) );
  XOR U10746 ( .A(b[57]), .B(a[10]), .Z(n10530) );
  NANDN U10747 ( .A(n38031), .B(n10530), .Z(n10220) );
  AND U10748 ( .A(n10221), .B(n10220), .Z(n10506) );
  NANDN U10749 ( .A(n38090), .B(n10222), .Z(n10224) );
  XOR U10750 ( .A(b[59]), .B(a[8]), .Z(n10533) );
  NANDN U10751 ( .A(n38130), .B(n10533), .Z(n10223) );
  AND U10752 ( .A(n10224), .B(n10223), .Z(n10504) );
  NANDN U10753 ( .A(n36480), .B(n10225), .Z(n10227) );
  XOR U10754 ( .A(b[41]), .B(a[26]), .Z(n10536) );
  NANDN U10755 ( .A(n36594), .B(n10536), .Z(n10226) );
  NAND U10756 ( .A(n10227), .B(n10226), .Z(n10503) );
  XNOR U10757 ( .A(n10504), .B(n10503), .Z(n10505) );
  XOR U10758 ( .A(n10506), .B(n10505), .Z(n10393) );
  XNOR U10759 ( .A(n10392), .B(n10393), .Z(n10394) );
  XNOR U10760 ( .A(n10395), .B(n10394), .Z(n10499) );
  XOR U10761 ( .A(n10500), .B(n10499), .Z(n10381) );
  NANDN U10762 ( .A(n10229), .B(n10228), .Z(n10233) );
  NAND U10763 ( .A(n10231), .B(n10230), .Z(n10232) );
  NAND U10764 ( .A(n10233), .B(n10232), .Z(n10380) );
  XNOR U10765 ( .A(n10381), .B(n10380), .Z(n10383) );
  NANDN U10766 ( .A(n10235), .B(n10234), .Z(n10239) );
  NAND U10767 ( .A(n10237), .B(n10236), .Z(n10238) );
  AND U10768 ( .A(n10239), .B(n10238), .Z(n10599) );
  NANDN U10769 ( .A(n32996), .B(n10240), .Z(n10242) );
  XOR U10770 ( .A(b[21]), .B(a[46]), .Z(n10551) );
  NANDN U10771 ( .A(n33271), .B(n10551), .Z(n10241) );
  AND U10772 ( .A(n10242), .B(n10241), .Z(n10517) );
  NANDN U10773 ( .A(n33866), .B(n10243), .Z(n10245) );
  XOR U10774 ( .A(b[23]), .B(a[44]), .Z(n10554) );
  NANDN U10775 ( .A(n33644), .B(n10554), .Z(n10244) );
  AND U10776 ( .A(n10245), .B(n10244), .Z(n10516) );
  NANDN U10777 ( .A(n32483), .B(n10246), .Z(n10248) );
  XOR U10778 ( .A(b[19]), .B(a[48]), .Z(n10557) );
  NANDN U10779 ( .A(n32823), .B(n10557), .Z(n10247) );
  NAND U10780 ( .A(n10248), .B(n10247), .Z(n10515) );
  XOR U10781 ( .A(n10516), .B(n10515), .Z(n10518) );
  XOR U10782 ( .A(n10517), .B(n10518), .Z(n10435) );
  NANDN U10783 ( .A(n34909), .B(n10249), .Z(n10251) );
  XOR U10784 ( .A(b[31]), .B(a[36]), .Z(n10560) );
  NANDN U10785 ( .A(n35145), .B(n10560), .Z(n10250) );
  AND U10786 ( .A(n10251), .B(n10250), .Z(n10475) );
  NANDN U10787 ( .A(n38247), .B(n10252), .Z(n10254) );
  XOR U10788 ( .A(b[61]), .B(a[6]), .Z(n10563) );
  NANDN U10789 ( .A(n38248), .B(n10563), .Z(n10253) );
  AND U10790 ( .A(n10254), .B(n10253), .Z(n10474) );
  AND U10791 ( .A(b[63]), .B(a[2]), .Z(n10473) );
  XOR U10792 ( .A(n10474), .B(n10473), .Z(n10476) );
  XNOR U10793 ( .A(n10475), .B(n10476), .Z(n10434) );
  XNOR U10794 ( .A(n10435), .B(n10434), .Z(n10436) );
  NANDN U10795 ( .A(n10256), .B(n10255), .Z(n10260) );
  OR U10796 ( .A(n10258), .B(n10257), .Z(n10259) );
  NAND U10797 ( .A(n10260), .B(n10259), .Z(n10437) );
  XNOR U10798 ( .A(n10436), .B(n10437), .Z(n10596) );
  NANDN U10799 ( .A(n34223), .B(n10261), .Z(n10263) );
  XOR U10800 ( .A(b[27]), .B(a[40]), .Z(n10572) );
  NANDN U10801 ( .A(n34458), .B(n10572), .Z(n10262) );
  AND U10802 ( .A(n10263), .B(n10262), .Z(n10418) );
  NANDN U10803 ( .A(n34634), .B(n10264), .Z(n10266) );
  XOR U10804 ( .A(b[29]), .B(a[38]), .Z(n10575) );
  NANDN U10805 ( .A(n34722), .B(n10575), .Z(n10265) );
  AND U10806 ( .A(n10266), .B(n10265), .Z(n10417) );
  NANDN U10807 ( .A(n31055), .B(n10267), .Z(n10269) );
  XOR U10808 ( .A(b[13]), .B(a[54]), .Z(n10578) );
  NANDN U10809 ( .A(n31293), .B(n10578), .Z(n10268) );
  NAND U10810 ( .A(n10269), .B(n10268), .Z(n10416) );
  XOR U10811 ( .A(n10417), .B(n10416), .Z(n10419) );
  XOR U10812 ( .A(n10418), .B(n10419), .Z(n10492) );
  NANDN U10813 ( .A(n28889), .B(n10270), .Z(n10272) );
  XOR U10814 ( .A(b[5]), .B(a[62]), .Z(n10581) );
  NANDN U10815 ( .A(n29138), .B(n10581), .Z(n10271) );
  AND U10816 ( .A(n10272), .B(n10271), .Z(n10511) );
  NANDN U10817 ( .A(n209), .B(n10273), .Z(n10275) );
  XOR U10818 ( .A(b[3]), .B(a[64]), .Z(n10584) );
  NANDN U10819 ( .A(n28941), .B(n10584), .Z(n10274) );
  AND U10820 ( .A(n10275), .B(n10274), .Z(n10510) );
  NANDN U10821 ( .A(n35936), .B(n10276), .Z(n10278) );
  XOR U10822 ( .A(b[37]), .B(a[30]), .Z(n10587) );
  NANDN U10823 ( .A(n36047), .B(n10587), .Z(n10277) );
  NAND U10824 ( .A(n10278), .B(n10277), .Z(n10509) );
  XOR U10825 ( .A(n10510), .B(n10509), .Z(n10512) );
  XNOR U10826 ( .A(n10511), .B(n10512), .Z(n10491) );
  XNOR U10827 ( .A(n10492), .B(n10491), .Z(n10493) );
  NANDN U10828 ( .A(n10280), .B(n10279), .Z(n10284) );
  OR U10829 ( .A(n10282), .B(n10281), .Z(n10283) );
  NAND U10830 ( .A(n10284), .B(n10283), .Z(n10494) );
  XOR U10831 ( .A(n10493), .B(n10494), .Z(n10597) );
  XNOR U10832 ( .A(n10596), .B(n10597), .Z(n10598) );
  XNOR U10833 ( .A(n10599), .B(n10598), .Z(n10382) );
  XOR U10834 ( .A(n10383), .B(n10382), .Z(n10375) );
  NANDN U10835 ( .A(n10286), .B(n10285), .Z(n10290) );
  NANDN U10836 ( .A(n10288), .B(n10287), .Z(n10289) );
  AND U10837 ( .A(n10290), .B(n10289), .Z(n10374) );
  XNOR U10838 ( .A(n10375), .B(n10374), .Z(n10376) );
  XOR U10839 ( .A(n10377), .B(n10376), .Z(n10609) );
  XNOR U10840 ( .A(n10608), .B(n10609), .Z(n10611) );
  NANDN U10841 ( .A(n10292), .B(n10291), .Z(n10296) );
  NANDN U10842 ( .A(n10294), .B(n10293), .Z(n10295) );
  AND U10843 ( .A(n10296), .B(n10295), .Z(n10610) );
  XOR U10844 ( .A(n10611), .B(n10610), .Z(n10616) );
  NANDN U10845 ( .A(n10298), .B(n10297), .Z(n10302) );
  NANDN U10846 ( .A(n10300), .B(n10299), .Z(n10301) );
  AND U10847 ( .A(n10302), .B(n10301), .Z(n10605) );
  NANDN U10848 ( .A(n10304), .B(n10303), .Z(n10308) );
  OR U10849 ( .A(n10306), .B(n10305), .Z(n10307) );
  AND U10850 ( .A(n10308), .B(n10307), .Z(n10603) );
  NANDN U10851 ( .A(n10310), .B(n10309), .Z(n10314) );
  OR U10852 ( .A(n10312), .B(n10311), .Z(n10313) );
  NAND U10853 ( .A(n10314), .B(n10313), .Z(n10602) );
  XNOR U10854 ( .A(n10603), .B(n10602), .Z(n10604) );
  XOR U10855 ( .A(n10605), .B(n10604), .Z(n10615) );
  NANDN U10856 ( .A(n10316), .B(n10315), .Z(n10320) );
  OR U10857 ( .A(n10318), .B(n10317), .Z(n10319) );
  AND U10858 ( .A(n10320), .B(n10319), .Z(n10614) );
  XOR U10859 ( .A(n10615), .B(n10614), .Z(n10617) );
  XOR U10860 ( .A(n10616), .B(n10617), .Z(n10623) );
  NAND U10861 ( .A(n10322), .B(n10321), .Z(n10326) );
  NAND U10862 ( .A(n10324), .B(n10323), .Z(n10325) );
  AND U10863 ( .A(n10326), .B(n10325), .Z(n10621) );
  NANDN U10864 ( .A(n10328), .B(n10327), .Z(n10332) );
  NANDN U10865 ( .A(n10330), .B(n10329), .Z(n10331) );
  AND U10866 ( .A(n10332), .B(n10331), .Z(n10620) );
  XNOR U10867 ( .A(n10621), .B(n10620), .Z(n10622) );
  XOR U10868 ( .A(n10623), .B(n10622), .Z(n10627) );
  XOR U10869 ( .A(n10626), .B(n10627), .Z(n10629) );
  XOR U10870 ( .A(n10628), .B(n10629), .Z(n10345) );
  NANDN U10871 ( .A(n10334), .B(n10333), .Z(n10338) );
  NAND U10872 ( .A(n10336), .B(n10335), .Z(n10337) );
  AND U10873 ( .A(n10338), .B(n10337), .Z(n10344) );
  XNOR U10874 ( .A(n10345), .B(n10344), .Z(n10346) );
  XNOR U10875 ( .A(n10347), .B(n10346), .Z(n10632) );
  XNOR U10876 ( .A(sreg[130]), .B(n10632), .Z(n10634) );
  NANDN U10877 ( .A(sreg[129]), .B(n10339), .Z(n10343) );
  NAND U10878 ( .A(n10341), .B(n10340), .Z(n10342) );
  NAND U10879 ( .A(n10343), .B(n10342), .Z(n10633) );
  XNOR U10880 ( .A(n10634), .B(n10633), .Z(c[130]) );
  NANDN U10881 ( .A(n10345), .B(n10344), .Z(n10349) );
  NANDN U10882 ( .A(n10347), .B(n10346), .Z(n10348) );
  AND U10883 ( .A(n10349), .B(n10348), .Z(n10640) );
  NANDN U10884 ( .A(n10351), .B(n10350), .Z(n10355) );
  OR U10885 ( .A(n10353), .B(n10352), .Z(n10354) );
  AND U10886 ( .A(n10355), .B(n10354), .Z(n10909) );
  NANDN U10887 ( .A(n10357), .B(n10356), .Z(n10361) );
  NAND U10888 ( .A(n10359), .B(n10358), .Z(n10360) );
  AND U10889 ( .A(n10361), .B(n10360), .Z(n10908) );
  NANDN U10890 ( .A(n10363), .B(n10362), .Z(n10367) );
  NANDN U10891 ( .A(n10365), .B(n10364), .Z(n10366) );
  AND U10892 ( .A(n10367), .B(n10366), .Z(n10907) );
  XOR U10893 ( .A(n10908), .B(n10907), .Z(n10910) );
  XOR U10894 ( .A(n10909), .B(n10910), .Z(n10914) );
  NANDN U10895 ( .A(n10369), .B(n10368), .Z(n10373) );
  NANDN U10896 ( .A(n10371), .B(n10370), .Z(n10372) );
  NAND U10897 ( .A(n10373), .B(n10372), .Z(n10913) );
  XNOR U10898 ( .A(n10914), .B(n10913), .Z(n10915) );
  NANDN U10899 ( .A(n10375), .B(n10374), .Z(n10379) );
  NANDN U10900 ( .A(n10377), .B(n10376), .Z(n10378) );
  AND U10901 ( .A(n10379), .B(n10378), .Z(n10904) );
  NANDN U10902 ( .A(n10381), .B(n10380), .Z(n10385) );
  NAND U10903 ( .A(n10383), .B(n10382), .Z(n10384) );
  AND U10904 ( .A(n10385), .B(n10384), .Z(n10669) );
  NANDN U10905 ( .A(n10387), .B(n10386), .Z(n10391) );
  NANDN U10906 ( .A(n10389), .B(n10388), .Z(n10390) );
  AND U10907 ( .A(n10391), .B(n10390), .Z(n10663) );
  NANDN U10908 ( .A(n10393), .B(n10392), .Z(n10397) );
  NANDN U10909 ( .A(n10395), .B(n10394), .Z(n10396) );
  AND U10910 ( .A(n10397), .B(n10396), .Z(n10662) );
  NANDN U10911 ( .A(n33875), .B(n10398), .Z(n10400) );
  XOR U10912 ( .A(b[25]), .B(a[43]), .Z(n10742) );
  NANDN U10913 ( .A(n33994), .B(n10742), .Z(n10399) );
  AND U10914 ( .A(n10400), .B(n10399), .Z(n10867) );
  NANDN U10915 ( .A(n32013), .B(n10401), .Z(n10403) );
  XOR U10916 ( .A(b[17]), .B(a[51]), .Z(n10745) );
  NANDN U10917 ( .A(n32292), .B(n10745), .Z(n10402) );
  AND U10918 ( .A(n10403), .B(n10402), .Z(n10866) );
  NANDN U10919 ( .A(n31536), .B(n10404), .Z(n10406) );
  XOR U10920 ( .A(b[15]), .B(a[53]), .Z(n10748) );
  NANDN U10921 ( .A(n31925), .B(n10748), .Z(n10405) );
  NAND U10922 ( .A(n10406), .B(n10405), .Z(n10865) );
  XOR U10923 ( .A(n10866), .B(n10865), .Z(n10868) );
  XOR U10924 ( .A(n10867), .B(n10868), .Z(n10839) );
  NANDN U10925 ( .A(n37526), .B(n10407), .Z(n10409) );
  XOR U10926 ( .A(b[51]), .B(a[17]), .Z(n10751) );
  NANDN U10927 ( .A(n37605), .B(n10751), .Z(n10408) );
  AND U10928 ( .A(n10409), .B(n10408), .Z(n10891) );
  NANDN U10929 ( .A(n37705), .B(n10410), .Z(n10412) );
  XOR U10930 ( .A(b[53]), .B(a[15]), .Z(n10754) );
  NANDN U10931 ( .A(n37778), .B(n10754), .Z(n10411) );
  AND U10932 ( .A(n10412), .B(n10411), .Z(n10890) );
  NANDN U10933 ( .A(n36210), .B(n10413), .Z(n10415) );
  XOR U10934 ( .A(b[39]), .B(a[29]), .Z(n10757) );
  NANDN U10935 ( .A(n36347), .B(n10757), .Z(n10414) );
  NAND U10936 ( .A(n10415), .B(n10414), .Z(n10889) );
  XOR U10937 ( .A(n10890), .B(n10889), .Z(n10892) );
  XNOR U10938 ( .A(n10891), .B(n10892), .Z(n10838) );
  XNOR U10939 ( .A(n10839), .B(n10838), .Z(n10841) );
  NANDN U10940 ( .A(n10417), .B(n10416), .Z(n10421) );
  OR U10941 ( .A(n10419), .B(n10418), .Z(n10420) );
  AND U10942 ( .A(n10421), .B(n10420), .Z(n10840) );
  XOR U10943 ( .A(n10841), .B(n10840), .Z(n10733) );
  NANDN U10944 ( .A(n10423), .B(n10422), .Z(n10427) );
  OR U10945 ( .A(n10425), .B(n10424), .Z(n10426) );
  AND U10946 ( .A(n10427), .B(n10426), .Z(n10731) );
  NANDN U10947 ( .A(n10429), .B(n10428), .Z(n10433) );
  NANDN U10948 ( .A(n10431), .B(n10430), .Z(n10432) );
  NAND U10949 ( .A(n10433), .B(n10432), .Z(n10730) );
  XNOR U10950 ( .A(n10731), .B(n10730), .Z(n10732) );
  XNOR U10951 ( .A(n10733), .B(n10732), .Z(n10661) );
  XOR U10952 ( .A(n10662), .B(n10661), .Z(n10664) );
  XOR U10953 ( .A(n10663), .B(n10664), .Z(n10668) );
  NANDN U10954 ( .A(n10435), .B(n10434), .Z(n10439) );
  NANDN U10955 ( .A(n10437), .B(n10436), .Z(n10438) );
  AND U10956 ( .A(n10439), .B(n10438), .Z(n10656) );
  NANDN U10957 ( .A(n211), .B(n10440), .Z(n10442) );
  XOR U10958 ( .A(b[47]), .B(a[21]), .Z(n10706) );
  NANDN U10959 ( .A(n37172), .B(n10706), .Z(n10441) );
  AND U10960 ( .A(n10442), .B(n10441), .Z(n10696) );
  NANDN U10961 ( .A(n210), .B(n10443), .Z(n10445) );
  XOR U10962 ( .A(b[9]), .B(a[59]), .Z(n10709) );
  NANDN U10963 ( .A(n30267), .B(n10709), .Z(n10444) );
  AND U10964 ( .A(n10445), .B(n10444), .Z(n10695) );
  NANDN U10965 ( .A(n212), .B(n10446), .Z(n10448) );
  XOR U10966 ( .A(b[49]), .B(a[19]), .Z(n10712) );
  NANDN U10967 ( .A(n37432), .B(n10712), .Z(n10447) );
  NAND U10968 ( .A(n10448), .B(n10447), .Z(n10694) );
  XOR U10969 ( .A(n10695), .B(n10694), .Z(n10697) );
  XOR U10970 ( .A(n10696), .B(n10697), .Z(n10845) );
  NANDN U10971 ( .A(n36742), .B(n10449), .Z(n10451) );
  XOR U10972 ( .A(b[43]), .B(a[25]), .Z(n10715) );
  NANDN U10973 ( .A(n36891), .B(n10715), .Z(n10450) );
  AND U10974 ( .A(n10451), .B(n10450), .Z(n10726) );
  NANDN U10975 ( .A(n36991), .B(n10452), .Z(n10454) );
  XOR U10976 ( .A(b[45]), .B(a[23]), .Z(n10718) );
  NANDN U10977 ( .A(n37083), .B(n10718), .Z(n10453) );
  AND U10978 ( .A(n10454), .B(n10453), .Z(n10725) );
  NANDN U10979 ( .A(n30482), .B(n10455), .Z(n10457) );
  XOR U10980 ( .A(b[11]), .B(a[57]), .Z(n10721) );
  NANDN U10981 ( .A(n30891), .B(n10721), .Z(n10456) );
  NAND U10982 ( .A(n10457), .B(n10456), .Z(n10724) );
  XOR U10983 ( .A(n10725), .B(n10724), .Z(n10727) );
  XNOR U10984 ( .A(n10726), .B(n10727), .Z(n10844) );
  XNOR U10985 ( .A(n10845), .B(n10844), .Z(n10846) );
  NANDN U10986 ( .A(n10459), .B(n10458), .Z(n10463) );
  OR U10987 ( .A(n10461), .B(n10460), .Z(n10462) );
  NAND U10988 ( .A(n10463), .B(n10462), .Z(n10847) );
  XNOR U10989 ( .A(n10846), .B(n10847), .Z(n10655) );
  XNOR U10990 ( .A(n10656), .B(n10655), .Z(n10657) );
  NANDN U10991 ( .A(n29499), .B(n10464), .Z(n10466) );
  XOR U10992 ( .A(b[7]), .B(a[61]), .Z(n10679) );
  NANDN U10993 ( .A(n29735), .B(n10679), .Z(n10465) );
  AND U10994 ( .A(n10466), .B(n10465), .Z(n10768) );
  NANDN U10995 ( .A(n37857), .B(n10467), .Z(n10469) );
  XOR U10996 ( .A(b[55]), .B(a[13]), .Z(n10682) );
  NANDN U10997 ( .A(n37911), .B(n10682), .Z(n10468) );
  AND U10998 ( .A(n10469), .B(n10468), .Z(n10767) );
  NANDN U10999 ( .A(n35611), .B(n10470), .Z(n10472) );
  XOR U11000 ( .A(b[35]), .B(a[33]), .Z(n10685) );
  NANDN U11001 ( .A(n35801), .B(n10685), .Z(n10471) );
  NAND U11002 ( .A(n10472), .B(n10471), .Z(n10766) );
  XOR U11003 ( .A(n10767), .B(n10766), .Z(n10769) );
  XOR U11004 ( .A(n10768), .B(n10769), .Z(n10785) );
  NANDN U11005 ( .A(n10474), .B(n10473), .Z(n10478) );
  OR U11006 ( .A(n10476), .B(n10475), .Z(n10477) );
  AND U11007 ( .A(n10478), .B(n10477), .Z(n10784) );
  XNOR U11008 ( .A(n10785), .B(n10784), .Z(n10786) );
  NANDN U11009 ( .A(n10480), .B(n10479), .Z(n10484) );
  OR U11010 ( .A(n10482), .B(n10481), .Z(n10483) );
  NAND U11011 ( .A(n10484), .B(n10483), .Z(n10787) );
  XOR U11012 ( .A(n10786), .B(n10787), .Z(n10658) );
  XNOR U11013 ( .A(n10657), .B(n10658), .Z(n10667) );
  XOR U11014 ( .A(n10668), .B(n10667), .Z(n10670) );
  XOR U11015 ( .A(n10669), .B(n10670), .Z(n10902) );
  NANDN U11016 ( .A(n10486), .B(n10485), .Z(n10490) );
  NANDN U11017 ( .A(n10488), .B(n10487), .Z(n10489) );
  AND U11018 ( .A(n10490), .B(n10489), .Z(n10651) );
  NANDN U11019 ( .A(n10492), .B(n10491), .Z(n10496) );
  NANDN U11020 ( .A(n10494), .B(n10493), .Z(n10495) );
  AND U11021 ( .A(n10496), .B(n10495), .Z(n10650) );
  NANDN U11022 ( .A(n10498), .B(n10497), .Z(n10502) );
  NAND U11023 ( .A(n10500), .B(n10499), .Z(n10501) );
  AND U11024 ( .A(n10502), .B(n10501), .Z(n10649) );
  XOR U11025 ( .A(n10650), .B(n10649), .Z(n10652) );
  XOR U11026 ( .A(n10651), .B(n10652), .Z(n10676) );
  NANDN U11027 ( .A(n10504), .B(n10503), .Z(n10508) );
  NANDN U11028 ( .A(n10506), .B(n10505), .Z(n10507) );
  AND U11029 ( .A(n10508), .B(n10507), .Z(n10797) );
  NANDN U11030 ( .A(n10510), .B(n10509), .Z(n10514) );
  OR U11031 ( .A(n10512), .B(n10511), .Z(n10513) );
  NAND U11032 ( .A(n10514), .B(n10513), .Z(n10796) );
  XNOR U11033 ( .A(n10797), .B(n10796), .Z(n10799) );
  NANDN U11034 ( .A(n10516), .B(n10515), .Z(n10520) );
  OR U11035 ( .A(n10518), .B(n10517), .Z(n10519) );
  AND U11036 ( .A(n10520), .B(n10519), .Z(n10739) );
  NAND U11037 ( .A(b[0]), .B(a[67]), .Z(n10521) );
  XNOR U11038 ( .A(b[1]), .B(n10521), .Z(n10523) );
  NANDN U11039 ( .A(b[0]), .B(a[66]), .Z(n10522) );
  NAND U11040 ( .A(n10523), .B(n10522), .Z(n10775) );
  NANDN U11041 ( .A(n38278), .B(n10524), .Z(n10526) );
  XOR U11042 ( .A(b[63]), .B(a[5]), .Z(n10823) );
  NANDN U11043 ( .A(n38279), .B(n10823), .Z(n10525) );
  AND U11044 ( .A(n10526), .B(n10525), .Z(n10773) );
  NANDN U11045 ( .A(n35260), .B(n10527), .Z(n10529) );
  XOR U11046 ( .A(b[33]), .B(a[35]), .Z(n10826) );
  NANDN U11047 ( .A(n35456), .B(n10826), .Z(n10528) );
  NAND U11048 ( .A(n10529), .B(n10528), .Z(n10772) );
  XNOR U11049 ( .A(n10773), .B(n10772), .Z(n10774) );
  XNOR U11050 ( .A(n10775), .B(n10774), .Z(n10736) );
  NANDN U11051 ( .A(n37974), .B(n10530), .Z(n10532) );
  XOR U11052 ( .A(b[57]), .B(a[11]), .Z(n10829) );
  NANDN U11053 ( .A(n38031), .B(n10829), .Z(n10531) );
  AND U11054 ( .A(n10532), .B(n10531), .Z(n10805) );
  NANDN U11055 ( .A(n38090), .B(n10533), .Z(n10535) );
  XOR U11056 ( .A(b[59]), .B(a[9]), .Z(n10832) );
  NANDN U11057 ( .A(n38130), .B(n10832), .Z(n10534) );
  AND U11058 ( .A(n10535), .B(n10534), .Z(n10803) );
  NANDN U11059 ( .A(n36480), .B(n10536), .Z(n10538) );
  XOR U11060 ( .A(b[41]), .B(a[27]), .Z(n10835) );
  NANDN U11061 ( .A(n36594), .B(n10835), .Z(n10537) );
  NAND U11062 ( .A(n10538), .B(n10537), .Z(n10802) );
  XNOR U11063 ( .A(n10803), .B(n10802), .Z(n10804) );
  XOR U11064 ( .A(n10805), .B(n10804), .Z(n10737) );
  XNOR U11065 ( .A(n10736), .B(n10737), .Z(n10738) );
  XNOR U11066 ( .A(n10739), .B(n10738), .Z(n10798) );
  XOR U11067 ( .A(n10799), .B(n10798), .Z(n10779) );
  NANDN U11068 ( .A(n10540), .B(n10539), .Z(n10544) );
  NAND U11069 ( .A(n10542), .B(n10541), .Z(n10543) );
  NAND U11070 ( .A(n10544), .B(n10543), .Z(n10778) );
  XNOR U11071 ( .A(n10779), .B(n10778), .Z(n10781) );
  NANDN U11072 ( .A(n10546), .B(n10545), .Z(n10550) );
  NANDN U11073 ( .A(n10548), .B(n10547), .Z(n10549) );
  AND U11074 ( .A(n10550), .B(n10549), .Z(n10898) );
  NANDN U11075 ( .A(n32996), .B(n10551), .Z(n10553) );
  XOR U11076 ( .A(b[21]), .B(a[47]), .Z(n10850) );
  NANDN U11077 ( .A(n33271), .B(n10850), .Z(n10552) );
  AND U11078 ( .A(n10553), .B(n10552), .Z(n10816) );
  NANDN U11079 ( .A(n33866), .B(n10554), .Z(n10556) );
  XOR U11080 ( .A(b[23]), .B(a[45]), .Z(n10853) );
  NANDN U11081 ( .A(n33644), .B(n10853), .Z(n10555) );
  AND U11082 ( .A(n10556), .B(n10555), .Z(n10815) );
  NANDN U11083 ( .A(n32483), .B(n10557), .Z(n10559) );
  XOR U11084 ( .A(b[19]), .B(a[49]), .Z(n10856) );
  NANDN U11085 ( .A(n32823), .B(n10856), .Z(n10558) );
  NAND U11086 ( .A(n10559), .B(n10558), .Z(n10814) );
  XOR U11087 ( .A(n10815), .B(n10814), .Z(n10817) );
  XOR U11088 ( .A(n10816), .B(n10817), .Z(n10701) );
  NANDN U11089 ( .A(n34909), .B(n10560), .Z(n10562) );
  XOR U11090 ( .A(b[31]), .B(a[37]), .Z(n10859) );
  NANDN U11091 ( .A(n35145), .B(n10859), .Z(n10561) );
  AND U11092 ( .A(n10562), .B(n10561), .Z(n10690) );
  NANDN U11093 ( .A(n38247), .B(n10563), .Z(n10565) );
  XOR U11094 ( .A(b[61]), .B(a[7]), .Z(n10862) );
  NANDN U11095 ( .A(n38248), .B(n10862), .Z(n10564) );
  AND U11096 ( .A(n10565), .B(n10564), .Z(n10689) );
  AND U11097 ( .A(b[63]), .B(a[3]), .Z(n10688) );
  XOR U11098 ( .A(n10689), .B(n10688), .Z(n10691) );
  XNOR U11099 ( .A(n10690), .B(n10691), .Z(n10700) );
  XNOR U11100 ( .A(n10701), .B(n10700), .Z(n10702) );
  NANDN U11101 ( .A(n10567), .B(n10566), .Z(n10571) );
  OR U11102 ( .A(n10569), .B(n10568), .Z(n10570) );
  NAND U11103 ( .A(n10571), .B(n10570), .Z(n10703) );
  XNOR U11104 ( .A(n10702), .B(n10703), .Z(n10895) );
  NANDN U11105 ( .A(n34223), .B(n10572), .Z(n10574) );
  XOR U11106 ( .A(b[27]), .B(a[41]), .Z(n10871) );
  NANDN U11107 ( .A(n34458), .B(n10871), .Z(n10573) );
  AND U11108 ( .A(n10574), .B(n10573), .Z(n10762) );
  NANDN U11109 ( .A(n34634), .B(n10575), .Z(n10577) );
  XOR U11110 ( .A(b[29]), .B(a[39]), .Z(n10874) );
  NANDN U11111 ( .A(n34722), .B(n10874), .Z(n10576) );
  AND U11112 ( .A(n10577), .B(n10576), .Z(n10761) );
  NANDN U11113 ( .A(n31055), .B(n10578), .Z(n10580) );
  XOR U11114 ( .A(b[13]), .B(a[55]), .Z(n10877) );
  NANDN U11115 ( .A(n31293), .B(n10877), .Z(n10579) );
  NAND U11116 ( .A(n10580), .B(n10579), .Z(n10760) );
  XOR U11117 ( .A(n10761), .B(n10760), .Z(n10763) );
  XOR U11118 ( .A(n10762), .B(n10763), .Z(n10791) );
  NANDN U11119 ( .A(n28889), .B(n10581), .Z(n10583) );
  XOR U11120 ( .A(b[5]), .B(a[63]), .Z(n10880) );
  NANDN U11121 ( .A(n29138), .B(n10880), .Z(n10582) );
  AND U11122 ( .A(n10583), .B(n10582), .Z(n10810) );
  NANDN U11123 ( .A(n209), .B(n10584), .Z(n10586) );
  XOR U11124 ( .A(b[3]), .B(a[65]), .Z(n10883) );
  NANDN U11125 ( .A(n28941), .B(n10883), .Z(n10585) );
  AND U11126 ( .A(n10586), .B(n10585), .Z(n10809) );
  NANDN U11127 ( .A(n35936), .B(n10587), .Z(n10589) );
  XOR U11128 ( .A(b[37]), .B(a[31]), .Z(n10886) );
  NANDN U11129 ( .A(n36047), .B(n10886), .Z(n10588) );
  NAND U11130 ( .A(n10589), .B(n10588), .Z(n10808) );
  XOR U11131 ( .A(n10809), .B(n10808), .Z(n10811) );
  XNOR U11132 ( .A(n10810), .B(n10811), .Z(n10790) );
  XNOR U11133 ( .A(n10791), .B(n10790), .Z(n10792) );
  NANDN U11134 ( .A(n10591), .B(n10590), .Z(n10595) );
  OR U11135 ( .A(n10593), .B(n10592), .Z(n10594) );
  NAND U11136 ( .A(n10595), .B(n10594), .Z(n10793) );
  XOR U11137 ( .A(n10792), .B(n10793), .Z(n10896) );
  XNOR U11138 ( .A(n10895), .B(n10896), .Z(n10897) );
  XNOR U11139 ( .A(n10898), .B(n10897), .Z(n10780) );
  XOR U11140 ( .A(n10781), .B(n10780), .Z(n10674) );
  NANDN U11141 ( .A(n10597), .B(n10596), .Z(n10601) );
  NANDN U11142 ( .A(n10599), .B(n10598), .Z(n10600) );
  AND U11143 ( .A(n10601), .B(n10600), .Z(n10673) );
  XNOR U11144 ( .A(n10674), .B(n10673), .Z(n10675) );
  XNOR U11145 ( .A(n10676), .B(n10675), .Z(n10901) );
  XNOR U11146 ( .A(n10902), .B(n10901), .Z(n10903) );
  XOR U11147 ( .A(n10904), .B(n10903), .Z(n10916) );
  XNOR U11148 ( .A(n10915), .B(n10916), .Z(n10922) );
  NANDN U11149 ( .A(n10603), .B(n10602), .Z(n10607) );
  NAND U11150 ( .A(n10605), .B(n10604), .Z(n10606) );
  AND U11151 ( .A(n10607), .B(n10606), .Z(n10920) );
  NANDN U11152 ( .A(n10609), .B(n10608), .Z(n10613) );
  NAND U11153 ( .A(n10611), .B(n10610), .Z(n10612) );
  NAND U11154 ( .A(n10613), .B(n10612), .Z(n10919) );
  XNOR U11155 ( .A(n10920), .B(n10919), .Z(n10921) );
  XOR U11156 ( .A(n10922), .B(n10921), .Z(n10644) );
  NANDN U11157 ( .A(n10615), .B(n10614), .Z(n10619) );
  OR U11158 ( .A(n10617), .B(n10616), .Z(n10618) );
  NAND U11159 ( .A(n10619), .B(n10618), .Z(n10643) );
  XNOR U11160 ( .A(n10644), .B(n10643), .Z(n10645) );
  NANDN U11161 ( .A(n10621), .B(n10620), .Z(n10625) );
  NANDN U11162 ( .A(n10623), .B(n10622), .Z(n10624) );
  NAND U11163 ( .A(n10625), .B(n10624), .Z(n10646) );
  XNOR U11164 ( .A(n10645), .B(n10646), .Z(n10637) );
  NANDN U11165 ( .A(n10627), .B(n10626), .Z(n10631) );
  OR U11166 ( .A(n10629), .B(n10628), .Z(n10630) );
  NAND U11167 ( .A(n10631), .B(n10630), .Z(n10638) );
  XNOR U11168 ( .A(n10637), .B(n10638), .Z(n10639) );
  XNOR U11169 ( .A(n10640), .B(n10639), .Z(n10925) );
  XNOR U11170 ( .A(sreg[131]), .B(n10925), .Z(n10927) );
  NANDN U11171 ( .A(sreg[130]), .B(n10632), .Z(n10636) );
  NAND U11172 ( .A(n10634), .B(n10633), .Z(n10635) );
  NAND U11173 ( .A(n10636), .B(n10635), .Z(n10926) );
  XNOR U11174 ( .A(n10927), .B(n10926), .Z(c[131]) );
  NANDN U11175 ( .A(n10638), .B(n10637), .Z(n10642) );
  NANDN U11176 ( .A(n10640), .B(n10639), .Z(n10641) );
  AND U11177 ( .A(n10642), .B(n10641), .Z(n10933) );
  NANDN U11178 ( .A(n10644), .B(n10643), .Z(n10648) );
  NANDN U11179 ( .A(n10646), .B(n10645), .Z(n10647) );
  AND U11180 ( .A(n10648), .B(n10647), .Z(n10931) );
  NANDN U11181 ( .A(n10650), .B(n10649), .Z(n10654) );
  OR U11182 ( .A(n10652), .B(n10651), .Z(n10653) );
  AND U11183 ( .A(n10654), .B(n10653), .Z(n11208) );
  NANDN U11184 ( .A(n10656), .B(n10655), .Z(n10660) );
  NANDN U11185 ( .A(n10658), .B(n10657), .Z(n10659) );
  AND U11186 ( .A(n10660), .B(n10659), .Z(n11207) );
  NANDN U11187 ( .A(n10662), .B(n10661), .Z(n10666) );
  OR U11188 ( .A(n10664), .B(n10663), .Z(n10665) );
  AND U11189 ( .A(n10666), .B(n10665), .Z(n11206) );
  XOR U11190 ( .A(n11207), .B(n11206), .Z(n11209) );
  XOR U11191 ( .A(n11208), .B(n11209), .Z(n10943) );
  NANDN U11192 ( .A(n10668), .B(n10667), .Z(n10672) );
  OR U11193 ( .A(n10670), .B(n10669), .Z(n10671) );
  AND U11194 ( .A(n10672), .B(n10671), .Z(n10942) );
  XNOR U11195 ( .A(n10943), .B(n10942), .Z(n10944) );
  NANDN U11196 ( .A(n10674), .B(n10673), .Z(n10678) );
  NANDN U11197 ( .A(n10676), .B(n10675), .Z(n10677) );
  AND U11198 ( .A(n10678), .B(n10677), .Z(n11203) );
  NANDN U11199 ( .A(n29499), .B(n10679), .Z(n10681) );
  XOR U11200 ( .A(b[7]), .B(a[62]), .Z(n11062) );
  NANDN U11201 ( .A(n29735), .B(n11062), .Z(n10680) );
  AND U11202 ( .A(n10681), .B(n10680), .Z(n11022) );
  NANDN U11203 ( .A(n37857), .B(n10682), .Z(n10684) );
  XOR U11204 ( .A(b[55]), .B(a[14]), .Z(n11065) );
  NANDN U11205 ( .A(n37911), .B(n11065), .Z(n10683) );
  AND U11206 ( .A(n10684), .B(n10683), .Z(n11021) );
  NANDN U11207 ( .A(n35611), .B(n10685), .Z(n10687) );
  XOR U11208 ( .A(b[35]), .B(a[34]), .Z(n11068) );
  NANDN U11209 ( .A(n35801), .B(n11068), .Z(n10686) );
  NAND U11210 ( .A(n10687), .B(n10686), .Z(n11020) );
  XOR U11211 ( .A(n11021), .B(n11020), .Z(n11023) );
  XOR U11212 ( .A(n11022), .B(n11023), .Z(n11084) );
  NANDN U11213 ( .A(n10689), .B(n10688), .Z(n10693) );
  OR U11214 ( .A(n10691), .B(n10690), .Z(n10692) );
  AND U11215 ( .A(n10693), .B(n10692), .Z(n11083) );
  XNOR U11216 ( .A(n11084), .B(n11083), .Z(n11085) );
  NANDN U11217 ( .A(n10695), .B(n10694), .Z(n10699) );
  OR U11218 ( .A(n10697), .B(n10696), .Z(n10698) );
  NAND U11219 ( .A(n10699), .B(n10698), .Z(n11086) );
  XNOR U11220 ( .A(n11085), .B(n11086), .Z(n10963) );
  NANDN U11221 ( .A(n10701), .B(n10700), .Z(n10705) );
  NANDN U11222 ( .A(n10703), .B(n10702), .Z(n10704) );
  AND U11223 ( .A(n10705), .B(n10704), .Z(n10961) );
  NAND U11224 ( .A(n37294), .B(n10706), .Z(n10708) );
  XNOR U11225 ( .A(b[47]), .B(a[22]), .Z(n11038) );
  NANDN U11226 ( .A(n11038), .B(n37341), .Z(n10707) );
  NAND U11227 ( .A(n10708), .B(n10707), .Z(n11079) );
  NAND U11228 ( .A(n30627), .B(n10709), .Z(n10711) );
  XNOR U11229 ( .A(b[9]), .B(a[60]), .Z(n11041) );
  NANDN U11230 ( .A(n11041), .B(n30628), .Z(n10710) );
  NAND U11231 ( .A(n10711), .B(n10710), .Z(n11078) );
  NAND U11232 ( .A(n37536), .B(n10712), .Z(n10714) );
  XNOR U11233 ( .A(b[49]), .B(a[20]), .Z(n11044) );
  NANDN U11234 ( .A(n11044), .B(n37537), .Z(n10713) );
  NAND U11235 ( .A(n10714), .B(n10713), .Z(n11077) );
  XNOR U11236 ( .A(n11078), .B(n11077), .Z(n11080) );
  NANDN U11237 ( .A(n36742), .B(n10715), .Z(n10717) );
  XOR U11238 ( .A(b[43]), .B(a[26]), .Z(n11047) );
  NANDN U11239 ( .A(n36891), .B(n11047), .Z(n10716) );
  AND U11240 ( .A(n10717), .B(n10716), .Z(n11058) );
  NANDN U11241 ( .A(n36991), .B(n10718), .Z(n10720) );
  XOR U11242 ( .A(b[45]), .B(a[24]), .Z(n11050) );
  NANDN U11243 ( .A(n37083), .B(n11050), .Z(n10719) );
  AND U11244 ( .A(n10720), .B(n10719), .Z(n11057) );
  NANDN U11245 ( .A(n30482), .B(n10721), .Z(n10723) );
  XOR U11246 ( .A(b[11]), .B(a[58]), .Z(n11053) );
  NANDN U11247 ( .A(n30891), .B(n11053), .Z(n10722) );
  NAND U11248 ( .A(n10723), .B(n10722), .Z(n11056) );
  XOR U11249 ( .A(n11057), .B(n11056), .Z(n11059) );
  XNOR U11250 ( .A(n11058), .B(n11059), .Z(n11143) );
  XOR U11251 ( .A(n11144), .B(n11143), .Z(n11145) );
  NANDN U11252 ( .A(n10725), .B(n10724), .Z(n10729) );
  OR U11253 ( .A(n10727), .B(n10726), .Z(n10728) );
  NAND U11254 ( .A(n10729), .B(n10728), .Z(n11146) );
  XNOR U11255 ( .A(n11145), .B(n11146), .Z(n10960) );
  XNOR U11256 ( .A(n10961), .B(n10960), .Z(n10962) );
  XOR U11257 ( .A(n10963), .B(n10962), .Z(n10949) );
  NANDN U11258 ( .A(n10731), .B(n10730), .Z(n10735) );
  NANDN U11259 ( .A(n10733), .B(n10732), .Z(n10734) );
  AND U11260 ( .A(n10735), .B(n10734), .Z(n10969) );
  NANDN U11261 ( .A(n10737), .B(n10736), .Z(n10741) );
  NANDN U11262 ( .A(n10739), .B(n10738), .Z(n10740) );
  AND U11263 ( .A(n10741), .B(n10740), .Z(n10967) );
  NANDN U11264 ( .A(n33875), .B(n10742), .Z(n10744) );
  XOR U11265 ( .A(b[25]), .B(a[44]), .Z(n10996) );
  NANDN U11266 ( .A(n33994), .B(n10996), .Z(n10743) );
  AND U11267 ( .A(n10744), .B(n10743), .Z(n11151) );
  NANDN U11268 ( .A(n32013), .B(n10745), .Z(n10747) );
  XOR U11269 ( .A(b[17]), .B(a[52]), .Z(n10999) );
  NANDN U11270 ( .A(n32292), .B(n10999), .Z(n10746) );
  AND U11271 ( .A(n10747), .B(n10746), .Z(n11150) );
  NANDN U11272 ( .A(n31536), .B(n10748), .Z(n10750) );
  XOR U11273 ( .A(b[15]), .B(a[54]), .Z(n11002) );
  NANDN U11274 ( .A(n31925), .B(n11002), .Z(n10749) );
  NAND U11275 ( .A(n10750), .B(n10749), .Z(n11149) );
  XOR U11276 ( .A(n11150), .B(n11149), .Z(n11152) );
  XOR U11277 ( .A(n11151), .B(n11152), .Z(n11138) );
  NANDN U11278 ( .A(n37526), .B(n10751), .Z(n10753) );
  XOR U11279 ( .A(b[51]), .B(a[18]), .Z(n11005) );
  NANDN U11280 ( .A(n37605), .B(n11005), .Z(n10752) );
  AND U11281 ( .A(n10753), .B(n10752), .Z(n11172) );
  NANDN U11282 ( .A(n37705), .B(n10754), .Z(n10756) );
  XOR U11283 ( .A(b[53]), .B(a[16]), .Z(n11008) );
  NANDN U11284 ( .A(n37778), .B(n11008), .Z(n10755) );
  AND U11285 ( .A(n10756), .B(n10755), .Z(n11171) );
  NANDN U11286 ( .A(n36210), .B(n10757), .Z(n10759) );
  XOR U11287 ( .A(b[39]), .B(a[30]), .Z(n11011) );
  NANDN U11288 ( .A(n36347), .B(n11011), .Z(n10758) );
  NAND U11289 ( .A(n10759), .B(n10758), .Z(n11170) );
  XOR U11290 ( .A(n11171), .B(n11170), .Z(n11173) );
  XNOR U11291 ( .A(n11172), .B(n11173), .Z(n11137) );
  XNOR U11292 ( .A(n11138), .B(n11137), .Z(n11140) );
  NANDN U11293 ( .A(n10761), .B(n10760), .Z(n10765) );
  OR U11294 ( .A(n10763), .B(n10762), .Z(n10764) );
  AND U11295 ( .A(n10765), .B(n10764), .Z(n11139) );
  XOR U11296 ( .A(n11140), .B(n11139), .Z(n10987) );
  NANDN U11297 ( .A(n10767), .B(n10766), .Z(n10771) );
  OR U11298 ( .A(n10769), .B(n10768), .Z(n10770) );
  AND U11299 ( .A(n10771), .B(n10770), .Z(n10985) );
  NANDN U11300 ( .A(n10773), .B(n10772), .Z(n10777) );
  NANDN U11301 ( .A(n10775), .B(n10774), .Z(n10776) );
  NAND U11302 ( .A(n10777), .B(n10776), .Z(n10984) );
  XNOR U11303 ( .A(n10985), .B(n10984), .Z(n10986) );
  XNOR U11304 ( .A(n10987), .B(n10986), .Z(n10966) );
  XNOR U11305 ( .A(n10967), .B(n10966), .Z(n10968) );
  XNOR U11306 ( .A(n10969), .B(n10968), .Z(n10948) );
  XNOR U11307 ( .A(n10949), .B(n10948), .Z(n10950) );
  NANDN U11308 ( .A(n10779), .B(n10778), .Z(n10783) );
  NAND U11309 ( .A(n10781), .B(n10780), .Z(n10782) );
  NAND U11310 ( .A(n10783), .B(n10782), .Z(n10951) );
  XNOR U11311 ( .A(n10950), .B(n10951), .Z(n11200) );
  NANDN U11312 ( .A(n10785), .B(n10784), .Z(n10789) );
  NANDN U11313 ( .A(n10787), .B(n10786), .Z(n10788) );
  AND U11314 ( .A(n10789), .B(n10788), .Z(n10956) );
  NANDN U11315 ( .A(n10791), .B(n10790), .Z(n10795) );
  NANDN U11316 ( .A(n10793), .B(n10792), .Z(n10794) );
  AND U11317 ( .A(n10795), .B(n10794), .Z(n10955) );
  NANDN U11318 ( .A(n10797), .B(n10796), .Z(n10801) );
  NAND U11319 ( .A(n10799), .B(n10798), .Z(n10800) );
  AND U11320 ( .A(n10801), .B(n10800), .Z(n10954) );
  XOR U11321 ( .A(n10955), .B(n10954), .Z(n10957) );
  XOR U11322 ( .A(n10956), .B(n10957), .Z(n10975) );
  NANDN U11323 ( .A(n10803), .B(n10802), .Z(n10807) );
  NANDN U11324 ( .A(n10805), .B(n10804), .Z(n10806) );
  AND U11325 ( .A(n10807), .B(n10806), .Z(n11096) );
  NANDN U11326 ( .A(n10809), .B(n10808), .Z(n10813) );
  OR U11327 ( .A(n10811), .B(n10810), .Z(n10812) );
  NAND U11328 ( .A(n10813), .B(n10812), .Z(n11095) );
  XNOR U11329 ( .A(n11096), .B(n11095), .Z(n11098) );
  NANDN U11330 ( .A(n10815), .B(n10814), .Z(n10819) );
  OR U11331 ( .A(n10817), .B(n10816), .Z(n10818) );
  AND U11332 ( .A(n10819), .B(n10818), .Z(n10993) );
  NAND U11333 ( .A(b[0]), .B(a[68]), .Z(n10820) );
  XNOR U11334 ( .A(b[1]), .B(n10820), .Z(n10822) );
  NANDN U11335 ( .A(b[0]), .B(a[67]), .Z(n10821) );
  NAND U11336 ( .A(n10822), .B(n10821), .Z(n11029) );
  NANDN U11337 ( .A(n38278), .B(n10823), .Z(n10825) );
  XOR U11338 ( .A(b[63]), .B(a[6]), .Z(n11122) );
  NANDN U11339 ( .A(n38279), .B(n11122), .Z(n10824) );
  AND U11340 ( .A(n10825), .B(n10824), .Z(n11027) );
  NANDN U11341 ( .A(n35260), .B(n10826), .Z(n10828) );
  XOR U11342 ( .A(b[33]), .B(a[36]), .Z(n11125) );
  NANDN U11343 ( .A(n35456), .B(n11125), .Z(n10827) );
  NAND U11344 ( .A(n10828), .B(n10827), .Z(n11026) );
  XNOR U11345 ( .A(n11027), .B(n11026), .Z(n11028) );
  XNOR U11346 ( .A(n11029), .B(n11028), .Z(n10990) );
  NANDN U11347 ( .A(n37974), .B(n10829), .Z(n10831) );
  XOR U11348 ( .A(b[57]), .B(a[12]), .Z(n11128) );
  NANDN U11349 ( .A(n38031), .B(n11128), .Z(n10830) );
  AND U11350 ( .A(n10831), .B(n10830), .Z(n11104) );
  NANDN U11351 ( .A(n38090), .B(n10832), .Z(n10834) );
  XOR U11352 ( .A(b[59]), .B(a[10]), .Z(n11131) );
  NANDN U11353 ( .A(n38130), .B(n11131), .Z(n10833) );
  AND U11354 ( .A(n10834), .B(n10833), .Z(n11102) );
  NANDN U11355 ( .A(n36480), .B(n10835), .Z(n10837) );
  XOR U11356 ( .A(b[41]), .B(a[28]), .Z(n11134) );
  NANDN U11357 ( .A(n36594), .B(n11134), .Z(n10836) );
  NAND U11358 ( .A(n10837), .B(n10836), .Z(n11101) );
  XNOR U11359 ( .A(n11102), .B(n11101), .Z(n11103) );
  XOR U11360 ( .A(n11104), .B(n11103), .Z(n10991) );
  XNOR U11361 ( .A(n10990), .B(n10991), .Z(n10992) );
  XNOR U11362 ( .A(n10993), .B(n10992), .Z(n11097) );
  XOR U11363 ( .A(n11098), .B(n11097), .Z(n10979) );
  NANDN U11364 ( .A(n10839), .B(n10838), .Z(n10843) );
  NAND U11365 ( .A(n10841), .B(n10840), .Z(n10842) );
  NAND U11366 ( .A(n10843), .B(n10842), .Z(n10978) );
  XNOR U11367 ( .A(n10979), .B(n10978), .Z(n10981) );
  NANDN U11368 ( .A(n10845), .B(n10844), .Z(n10849) );
  NANDN U11369 ( .A(n10847), .B(n10846), .Z(n10848) );
  AND U11370 ( .A(n10849), .B(n10848), .Z(n11197) );
  NANDN U11371 ( .A(n32996), .B(n10850), .Z(n10852) );
  XOR U11372 ( .A(b[21]), .B(a[48]), .Z(n11155) );
  NANDN U11373 ( .A(n33271), .B(n11155), .Z(n10851) );
  AND U11374 ( .A(n10852), .B(n10851), .Z(n11115) );
  NANDN U11375 ( .A(n33866), .B(n10853), .Z(n10855) );
  XOR U11376 ( .A(b[23]), .B(a[46]), .Z(n11158) );
  NANDN U11377 ( .A(n33644), .B(n11158), .Z(n10854) );
  AND U11378 ( .A(n10855), .B(n10854), .Z(n11114) );
  NANDN U11379 ( .A(n32483), .B(n10856), .Z(n10858) );
  XOR U11380 ( .A(b[19]), .B(a[50]), .Z(n11161) );
  NANDN U11381 ( .A(n32823), .B(n11161), .Z(n10857) );
  NAND U11382 ( .A(n10858), .B(n10857), .Z(n11113) );
  XOR U11383 ( .A(n11114), .B(n11113), .Z(n11116) );
  XOR U11384 ( .A(n11115), .B(n11116), .Z(n11033) );
  NANDN U11385 ( .A(n34909), .B(n10859), .Z(n10861) );
  XOR U11386 ( .A(b[31]), .B(a[38]), .Z(n11164) );
  NANDN U11387 ( .A(n35145), .B(n11164), .Z(n10860) );
  AND U11388 ( .A(n10861), .B(n10860), .Z(n11073) );
  NANDN U11389 ( .A(n38247), .B(n10862), .Z(n10864) );
  XOR U11390 ( .A(b[61]), .B(a[8]), .Z(n11167) );
  NANDN U11391 ( .A(n38248), .B(n11167), .Z(n10863) );
  AND U11392 ( .A(n10864), .B(n10863), .Z(n11072) );
  AND U11393 ( .A(b[63]), .B(a[4]), .Z(n11071) );
  XOR U11394 ( .A(n11072), .B(n11071), .Z(n11074) );
  XNOR U11395 ( .A(n11073), .B(n11074), .Z(n11032) );
  XNOR U11396 ( .A(n11033), .B(n11032), .Z(n11034) );
  NANDN U11397 ( .A(n10866), .B(n10865), .Z(n10870) );
  OR U11398 ( .A(n10868), .B(n10867), .Z(n10869) );
  NAND U11399 ( .A(n10870), .B(n10869), .Z(n11035) );
  XNOR U11400 ( .A(n11034), .B(n11035), .Z(n11194) );
  NANDN U11401 ( .A(n34223), .B(n10871), .Z(n10873) );
  XOR U11402 ( .A(b[27]), .B(a[42]), .Z(n11176) );
  NANDN U11403 ( .A(n34458), .B(n11176), .Z(n10872) );
  AND U11404 ( .A(n10873), .B(n10872), .Z(n11016) );
  NANDN U11405 ( .A(n34634), .B(n10874), .Z(n10876) );
  XOR U11406 ( .A(b[29]), .B(a[40]), .Z(n11179) );
  NANDN U11407 ( .A(n34722), .B(n11179), .Z(n10875) );
  AND U11408 ( .A(n10876), .B(n10875), .Z(n11015) );
  NANDN U11409 ( .A(n31055), .B(n10877), .Z(n10879) );
  XOR U11410 ( .A(b[13]), .B(a[56]), .Z(n11182) );
  NANDN U11411 ( .A(n31293), .B(n11182), .Z(n10878) );
  NAND U11412 ( .A(n10879), .B(n10878), .Z(n11014) );
  XOR U11413 ( .A(n11015), .B(n11014), .Z(n11017) );
  XOR U11414 ( .A(n11016), .B(n11017), .Z(n11090) );
  NANDN U11415 ( .A(n28889), .B(n10880), .Z(n10882) );
  XOR U11416 ( .A(b[5]), .B(a[64]), .Z(n11185) );
  NANDN U11417 ( .A(n29138), .B(n11185), .Z(n10881) );
  AND U11418 ( .A(n10882), .B(n10881), .Z(n11109) );
  NANDN U11419 ( .A(n209), .B(n10883), .Z(n10885) );
  XOR U11420 ( .A(b[3]), .B(a[66]), .Z(n11188) );
  NANDN U11421 ( .A(n28941), .B(n11188), .Z(n10884) );
  AND U11422 ( .A(n10885), .B(n10884), .Z(n11108) );
  NANDN U11423 ( .A(n35936), .B(n10886), .Z(n10888) );
  XOR U11424 ( .A(b[37]), .B(a[32]), .Z(n11191) );
  NANDN U11425 ( .A(n36047), .B(n11191), .Z(n10887) );
  NAND U11426 ( .A(n10888), .B(n10887), .Z(n11107) );
  XOR U11427 ( .A(n11108), .B(n11107), .Z(n11110) );
  XNOR U11428 ( .A(n11109), .B(n11110), .Z(n11089) );
  XNOR U11429 ( .A(n11090), .B(n11089), .Z(n11091) );
  NANDN U11430 ( .A(n10890), .B(n10889), .Z(n10894) );
  OR U11431 ( .A(n10892), .B(n10891), .Z(n10893) );
  NAND U11432 ( .A(n10894), .B(n10893), .Z(n11092) );
  XOR U11433 ( .A(n11091), .B(n11092), .Z(n11195) );
  XNOR U11434 ( .A(n11194), .B(n11195), .Z(n11196) );
  XNOR U11435 ( .A(n11197), .B(n11196), .Z(n10980) );
  XOR U11436 ( .A(n10981), .B(n10980), .Z(n10973) );
  NANDN U11437 ( .A(n10896), .B(n10895), .Z(n10900) );
  NANDN U11438 ( .A(n10898), .B(n10897), .Z(n10899) );
  AND U11439 ( .A(n10900), .B(n10899), .Z(n10972) );
  XNOR U11440 ( .A(n10973), .B(n10972), .Z(n10974) );
  XOR U11441 ( .A(n10975), .B(n10974), .Z(n11201) );
  XNOR U11442 ( .A(n11200), .B(n11201), .Z(n11202) );
  XOR U11443 ( .A(n11203), .B(n11202), .Z(n10945) );
  XNOR U11444 ( .A(n10944), .B(n10945), .Z(n10939) );
  NANDN U11445 ( .A(n10902), .B(n10901), .Z(n10906) );
  NANDN U11446 ( .A(n10904), .B(n10903), .Z(n10905) );
  AND U11447 ( .A(n10906), .B(n10905), .Z(n10937) );
  NANDN U11448 ( .A(n10908), .B(n10907), .Z(n10912) );
  OR U11449 ( .A(n10910), .B(n10909), .Z(n10911) );
  AND U11450 ( .A(n10912), .B(n10911), .Z(n10936) );
  XNOR U11451 ( .A(n10937), .B(n10936), .Z(n10938) );
  XOR U11452 ( .A(n10939), .B(n10938), .Z(n11213) );
  NANDN U11453 ( .A(n10914), .B(n10913), .Z(n10918) );
  NANDN U11454 ( .A(n10916), .B(n10915), .Z(n10917) );
  AND U11455 ( .A(n10918), .B(n10917), .Z(n11212) );
  XNOR U11456 ( .A(n11213), .B(n11212), .Z(n11214) );
  NANDN U11457 ( .A(n10920), .B(n10919), .Z(n10924) );
  NAND U11458 ( .A(n10922), .B(n10921), .Z(n10923) );
  NAND U11459 ( .A(n10924), .B(n10923), .Z(n11215) );
  XNOR U11460 ( .A(n11214), .B(n11215), .Z(n10930) );
  XNOR U11461 ( .A(n10931), .B(n10930), .Z(n10932) );
  XNOR U11462 ( .A(n10933), .B(n10932), .Z(n11218) );
  XNOR U11463 ( .A(sreg[132]), .B(n11218), .Z(n11220) );
  NANDN U11464 ( .A(sreg[131]), .B(n10925), .Z(n10929) );
  NAND U11465 ( .A(n10927), .B(n10926), .Z(n10928) );
  NAND U11466 ( .A(n10929), .B(n10928), .Z(n11219) );
  XNOR U11467 ( .A(n11220), .B(n11219), .Z(c[132]) );
  NANDN U11468 ( .A(n10931), .B(n10930), .Z(n10935) );
  NANDN U11469 ( .A(n10933), .B(n10932), .Z(n10934) );
  AND U11470 ( .A(n10935), .B(n10934), .Z(n11226) );
  NANDN U11471 ( .A(n10937), .B(n10936), .Z(n10941) );
  NAND U11472 ( .A(n10939), .B(n10938), .Z(n10940) );
  AND U11473 ( .A(n10941), .B(n10940), .Z(n11231) );
  NANDN U11474 ( .A(n10943), .B(n10942), .Z(n10947) );
  NANDN U11475 ( .A(n10945), .B(n10944), .Z(n10946) );
  AND U11476 ( .A(n10947), .B(n10946), .Z(n11230) );
  NANDN U11477 ( .A(n10949), .B(n10948), .Z(n10953) );
  NANDN U11478 ( .A(n10951), .B(n10950), .Z(n10952) );
  AND U11479 ( .A(n10953), .B(n10952), .Z(n11498) );
  NANDN U11480 ( .A(n10955), .B(n10954), .Z(n10959) );
  OR U11481 ( .A(n10957), .B(n10956), .Z(n10958) );
  AND U11482 ( .A(n10959), .B(n10958), .Z(n11493) );
  NANDN U11483 ( .A(n10961), .B(n10960), .Z(n10965) );
  NAND U11484 ( .A(n10963), .B(n10962), .Z(n10964) );
  AND U11485 ( .A(n10965), .B(n10964), .Z(n11492) );
  NANDN U11486 ( .A(n10967), .B(n10966), .Z(n10971) );
  NANDN U11487 ( .A(n10969), .B(n10968), .Z(n10970) );
  AND U11488 ( .A(n10971), .B(n10970), .Z(n11491) );
  XOR U11489 ( .A(n11492), .B(n11491), .Z(n11494) );
  XNOR U11490 ( .A(n11493), .B(n11494), .Z(n11497) );
  XNOR U11491 ( .A(n11498), .B(n11497), .Z(n11499) );
  NANDN U11492 ( .A(n10973), .B(n10972), .Z(n10977) );
  NANDN U11493 ( .A(n10975), .B(n10974), .Z(n10976) );
  AND U11494 ( .A(n10977), .B(n10976), .Z(n11488) );
  NANDN U11495 ( .A(n10979), .B(n10978), .Z(n10983) );
  NAND U11496 ( .A(n10981), .B(n10980), .Z(n10982) );
  AND U11497 ( .A(n10983), .B(n10982), .Z(n11463) );
  NANDN U11498 ( .A(n10985), .B(n10984), .Z(n10989) );
  NANDN U11499 ( .A(n10987), .B(n10986), .Z(n10988) );
  AND U11500 ( .A(n10989), .B(n10988), .Z(n11481) );
  NANDN U11501 ( .A(n10991), .B(n10990), .Z(n10995) );
  NANDN U11502 ( .A(n10993), .B(n10992), .Z(n10994) );
  AND U11503 ( .A(n10995), .B(n10994), .Z(n11480) );
  NANDN U11504 ( .A(n33875), .B(n10996), .Z(n10998) );
  XOR U11505 ( .A(b[25]), .B(a[45]), .Z(n11259) );
  NANDN U11506 ( .A(n33994), .B(n11259), .Z(n10997) );
  AND U11507 ( .A(n10998), .B(n10997), .Z(n11429) );
  NANDN U11508 ( .A(n32013), .B(n10999), .Z(n11001) );
  XOR U11509 ( .A(b[17]), .B(a[53]), .Z(n11262) );
  NANDN U11510 ( .A(n32292), .B(n11262), .Z(n11000) );
  AND U11511 ( .A(n11001), .B(n11000), .Z(n11428) );
  NANDN U11512 ( .A(n31536), .B(n11002), .Z(n11004) );
  XOR U11513 ( .A(b[15]), .B(a[55]), .Z(n11265) );
  NANDN U11514 ( .A(n31925), .B(n11265), .Z(n11003) );
  NAND U11515 ( .A(n11004), .B(n11003), .Z(n11427) );
  XOR U11516 ( .A(n11428), .B(n11427), .Z(n11430) );
  XOR U11517 ( .A(n11429), .B(n11430), .Z(n11401) );
  NANDN U11518 ( .A(n37526), .B(n11005), .Z(n11007) );
  XOR U11519 ( .A(b[51]), .B(a[19]), .Z(n11268) );
  NANDN U11520 ( .A(n37605), .B(n11268), .Z(n11006) );
  AND U11521 ( .A(n11007), .B(n11006), .Z(n11453) );
  NANDN U11522 ( .A(n37705), .B(n11008), .Z(n11010) );
  XOR U11523 ( .A(b[53]), .B(a[17]), .Z(n11271) );
  NANDN U11524 ( .A(n37778), .B(n11271), .Z(n11009) );
  AND U11525 ( .A(n11010), .B(n11009), .Z(n11452) );
  NANDN U11526 ( .A(n36210), .B(n11011), .Z(n11013) );
  XOR U11527 ( .A(b[39]), .B(a[31]), .Z(n11274) );
  NANDN U11528 ( .A(n36347), .B(n11274), .Z(n11012) );
  NAND U11529 ( .A(n11013), .B(n11012), .Z(n11451) );
  XOR U11530 ( .A(n11452), .B(n11451), .Z(n11454) );
  XNOR U11531 ( .A(n11453), .B(n11454), .Z(n11400) );
  XNOR U11532 ( .A(n11401), .B(n11400), .Z(n11403) );
  NANDN U11533 ( .A(n11015), .B(n11014), .Z(n11019) );
  OR U11534 ( .A(n11017), .B(n11016), .Z(n11018) );
  AND U11535 ( .A(n11019), .B(n11018), .Z(n11402) );
  XOR U11536 ( .A(n11403), .B(n11402), .Z(n11250) );
  NANDN U11537 ( .A(n11021), .B(n11020), .Z(n11025) );
  OR U11538 ( .A(n11023), .B(n11022), .Z(n11024) );
  AND U11539 ( .A(n11025), .B(n11024), .Z(n11248) );
  NANDN U11540 ( .A(n11027), .B(n11026), .Z(n11031) );
  NANDN U11541 ( .A(n11029), .B(n11028), .Z(n11030) );
  NAND U11542 ( .A(n11031), .B(n11030), .Z(n11247) );
  XNOR U11543 ( .A(n11248), .B(n11247), .Z(n11249) );
  XNOR U11544 ( .A(n11250), .B(n11249), .Z(n11479) );
  XOR U11545 ( .A(n11480), .B(n11479), .Z(n11482) );
  XOR U11546 ( .A(n11481), .B(n11482), .Z(n11462) );
  NANDN U11547 ( .A(n11033), .B(n11032), .Z(n11037) );
  NANDN U11548 ( .A(n11035), .B(n11034), .Z(n11036) );
  AND U11549 ( .A(n11037), .B(n11036), .Z(n11474) );
  NANDN U11550 ( .A(n11038), .B(n37294), .Z(n11040) );
  XOR U11551 ( .A(b[47]), .B(a[23]), .Z(n11322) );
  NANDN U11552 ( .A(n37172), .B(n11322), .Z(n11039) );
  AND U11553 ( .A(n11040), .B(n11039), .Z(n11312) );
  NANDN U11554 ( .A(n11041), .B(n30627), .Z(n11043) );
  XOR U11555 ( .A(b[9]), .B(a[61]), .Z(n11325) );
  NANDN U11556 ( .A(n30267), .B(n11325), .Z(n11042) );
  AND U11557 ( .A(n11043), .B(n11042), .Z(n11311) );
  NANDN U11558 ( .A(n11044), .B(n37536), .Z(n11046) );
  XOR U11559 ( .A(b[49]), .B(a[21]), .Z(n11328) );
  NANDN U11560 ( .A(n37432), .B(n11328), .Z(n11045) );
  NAND U11561 ( .A(n11046), .B(n11045), .Z(n11310) );
  XOR U11562 ( .A(n11311), .B(n11310), .Z(n11313) );
  XOR U11563 ( .A(n11312), .B(n11313), .Z(n11407) );
  NANDN U11564 ( .A(n36742), .B(n11047), .Z(n11049) );
  XOR U11565 ( .A(b[43]), .B(a[27]), .Z(n11331) );
  NANDN U11566 ( .A(n36891), .B(n11331), .Z(n11048) );
  AND U11567 ( .A(n11049), .B(n11048), .Z(n11342) );
  NANDN U11568 ( .A(n36991), .B(n11050), .Z(n11052) );
  XOR U11569 ( .A(b[45]), .B(a[25]), .Z(n11334) );
  NANDN U11570 ( .A(n37083), .B(n11334), .Z(n11051) );
  AND U11571 ( .A(n11052), .B(n11051), .Z(n11341) );
  NANDN U11572 ( .A(n30482), .B(n11053), .Z(n11055) );
  XOR U11573 ( .A(b[11]), .B(a[59]), .Z(n11337) );
  NANDN U11574 ( .A(n30891), .B(n11337), .Z(n11054) );
  NAND U11575 ( .A(n11055), .B(n11054), .Z(n11340) );
  XOR U11576 ( .A(n11341), .B(n11340), .Z(n11343) );
  XNOR U11577 ( .A(n11342), .B(n11343), .Z(n11406) );
  XNOR U11578 ( .A(n11407), .B(n11406), .Z(n11408) );
  NANDN U11579 ( .A(n11057), .B(n11056), .Z(n11061) );
  OR U11580 ( .A(n11059), .B(n11058), .Z(n11060) );
  NAND U11581 ( .A(n11061), .B(n11060), .Z(n11409) );
  XNOR U11582 ( .A(n11408), .B(n11409), .Z(n11473) );
  XNOR U11583 ( .A(n11474), .B(n11473), .Z(n11475) );
  NANDN U11584 ( .A(n29499), .B(n11062), .Z(n11064) );
  XOR U11585 ( .A(b[7]), .B(a[63]), .Z(n11295) );
  NANDN U11586 ( .A(n29735), .B(n11295), .Z(n11063) );
  AND U11587 ( .A(n11064), .B(n11063), .Z(n11285) );
  NANDN U11588 ( .A(n37857), .B(n11065), .Z(n11067) );
  XOR U11589 ( .A(b[55]), .B(a[15]), .Z(n11298) );
  NANDN U11590 ( .A(n37911), .B(n11298), .Z(n11066) );
  AND U11591 ( .A(n11067), .B(n11066), .Z(n11284) );
  NANDN U11592 ( .A(n35611), .B(n11068), .Z(n11070) );
  XOR U11593 ( .A(b[35]), .B(a[35]), .Z(n11301) );
  NANDN U11594 ( .A(n35801), .B(n11301), .Z(n11069) );
  NAND U11595 ( .A(n11070), .B(n11069), .Z(n11283) );
  XOR U11596 ( .A(n11284), .B(n11283), .Z(n11286) );
  XOR U11597 ( .A(n11285), .B(n11286), .Z(n11359) );
  NANDN U11598 ( .A(n11072), .B(n11071), .Z(n11076) );
  OR U11599 ( .A(n11074), .B(n11073), .Z(n11075) );
  AND U11600 ( .A(n11076), .B(n11075), .Z(n11358) );
  XNOR U11601 ( .A(n11359), .B(n11358), .Z(n11360) );
  NAND U11602 ( .A(n11078), .B(n11077), .Z(n11082) );
  NANDN U11603 ( .A(n11080), .B(n11079), .Z(n11081) );
  NAND U11604 ( .A(n11082), .B(n11081), .Z(n11361) );
  XOR U11605 ( .A(n11360), .B(n11361), .Z(n11476) );
  XNOR U11606 ( .A(n11475), .B(n11476), .Z(n11461) );
  XOR U11607 ( .A(n11462), .B(n11461), .Z(n11464) );
  XOR U11608 ( .A(n11463), .B(n11464), .Z(n11486) );
  NANDN U11609 ( .A(n11084), .B(n11083), .Z(n11088) );
  NANDN U11610 ( .A(n11086), .B(n11085), .Z(n11087) );
  AND U11611 ( .A(n11088), .B(n11087), .Z(n11469) );
  NANDN U11612 ( .A(n11090), .B(n11089), .Z(n11094) );
  NANDN U11613 ( .A(n11092), .B(n11091), .Z(n11093) );
  AND U11614 ( .A(n11094), .B(n11093), .Z(n11468) );
  NANDN U11615 ( .A(n11096), .B(n11095), .Z(n11100) );
  NAND U11616 ( .A(n11098), .B(n11097), .Z(n11099) );
  AND U11617 ( .A(n11100), .B(n11099), .Z(n11467) );
  XOR U11618 ( .A(n11468), .B(n11467), .Z(n11470) );
  XOR U11619 ( .A(n11469), .B(n11470), .Z(n11238) );
  NANDN U11620 ( .A(n11102), .B(n11101), .Z(n11106) );
  NANDN U11621 ( .A(n11104), .B(n11103), .Z(n11105) );
  AND U11622 ( .A(n11106), .B(n11105), .Z(n11353) );
  NANDN U11623 ( .A(n11108), .B(n11107), .Z(n11112) );
  OR U11624 ( .A(n11110), .B(n11109), .Z(n11111) );
  NAND U11625 ( .A(n11112), .B(n11111), .Z(n11352) );
  XNOR U11626 ( .A(n11353), .B(n11352), .Z(n11355) );
  NANDN U11627 ( .A(n11114), .B(n11113), .Z(n11118) );
  OR U11628 ( .A(n11116), .B(n11115), .Z(n11117) );
  NAND U11629 ( .A(n11118), .B(n11117), .Z(n11255) );
  NAND U11630 ( .A(b[0]), .B(a[69]), .Z(n11119) );
  XNOR U11631 ( .A(b[1]), .B(n11119), .Z(n11121) );
  NANDN U11632 ( .A(b[0]), .B(a[68]), .Z(n11120) );
  NAND U11633 ( .A(n11121), .B(n11120), .Z(n11292) );
  NANDN U11634 ( .A(n38278), .B(n11122), .Z(n11124) );
  XOR U11635 ( .A(b[63]), .B(a[7]), .Z(n11385) );
  NANDN U11636 ( .A(n38279), .B(n11385), .Z(n11123) );
  AND U11637 ( .A(n11124), .B(n11123), .Z(n11290) );
  NANDN U11638 ( .A(n35260), .B(n11125), .Z(n11127) );
  XOR U11639 ( .A(b[33]), .B(a[37]), .Z(n11388) );
  NANDN U11640 ( .A(n35456), .B(n11388), .Z(n11126) );
  NAND U11641 ( .A(n11127), .B(n11126), .Z(n11289) );
  XNOR U11642 ( .A(n11290), .B(n11289), .Z(n11291) );
  XNOR U11643 ( .A(n11292), .B(n11291), .Z(n11254) );
  NANDN U11644 ( .A(n37974), .B(n11128), .Z(n11130) );
  XOR U11645 ( .A(b[57]), .B(a[13]), .Z(n11391) );
  NANDN U11646 ( .A(n38031), .B(n11391), .Z(n11129) );
  AND U11647 ( .A(n11130), .B(n11129), .Z(n11366) );
  NANDN U11648 ( .A(n38090), .B(n11131), .Z(n11133) );
  XOR U11649 ( .A(b[59]), .B(a[11]), .Z(n11394) );
  NANDN U11650 ( .A(n38130), .B(n11394), .Z(n11132) );
  AND U11651 ( .A(n11133), .B(n11132), .Z(n11365) );
  NANDN U11652 ( .A(n36480), .B(n11134), .Z(n11136) );
  XOR U11653 ( .A(b[41]), .B(a[29]), .Z(n11397) );
  NANDN U11654 ( .A(n36594), .B(n11397), .Z(n11135) );
  NAND U11655 ( .A(n11136), .B(n11135), .Z(n11364) );
  XOR U11656 ( .A(n11365), .B(n11364), .Z(n11367) );
  XOR U11657 ( .A(n11366), .B(n11367), .Z(n11253) );
  XOR U11658 ( .A(n11254), .B(n11253), .Z(n11256) );
  XOR U11659 ( .A(n11255), .B(n11256), .Z(n11354) );
  XOR U11660 ( .A(n11355), .B(n11354), .Z(n11242) );
  NANDN U11661 ( .A(n11138), .B(n11137), .Z(n11142) );
  NAND U11662 ( .A(n11140), .B(n11139), .Z(n11141) );
  NAND U11663 ( .A(n11142), .B(n11141), .Z(n11241) );
  XNOR U11664 ( .A(n11242), .B(n11241), .Z(n11244) );
  NAND U11665 ( .A(n11144), .B(n11143), .Z(n11148) );
  NANDN U11666 ( .A(n11146), .B(n11145), .Z(n11147) );
  AND U11667 ( .A(n11148), .B(n11147), .Z(n11460) );
  NANDN U11668 ( .A(n11150), .B(n11149), .Z(n11154) );
  OR U11669 ( .A(n11152), .B(n11151), .Z(n11153) );
  AND U11670 ( .A(n11154), .B(n11153), .Z(n11318) );
  NANDN U11671 ( .A(n32996), .B(n11155), .Z(n11157) );
  XOR U11672 ( .A(b[21]), .B(a[49]), .Z(n11412) );
  NANDN U11673 ( .A(n33271), .B(n11412), .Z(n11156) );
  AND U11674 ( .A(n11157), .B(n11156), .Z(n11379) );
  NANDN U11675 ( .A(n33866), .B(n11158), .Z(n11160) );
  XOR U11676 ( .A(b[23]), .B(a[47]), .Z(n11415) );
  NANDN U11677 ( .A(n33644), .B(n11415), .Z(n11159) );
  AND U11678 ( .A(n11160), .B(n11159), .Z(n11377) );
  NANDN U11679 ( .A(n32483), .B(n11161), .Z(n11163) );
  XOR U11680 ( .A(b[19]), .B(a[51]), .Z(n11418) );
  NANDN U11681 ( .A(n32823), .B(n11418), .Z(n11162) );
  NAND U11682 ( .A(n11163), .B(n11162), .Z(n11376) );
  XNOR U11683 ( .A(n11377), .B(n11376), .Z(n11378) );
  XOR U11684 ( .A(n11379), .B(n11378), .Z(n11317) );
  NANDN U11685 ( .A(n34909), .B(n11164), .Z(n11166) );
  XOR U11686 ( .A(b[31]), .B(a[39]), .Z(n11421) );
  NANDN U11687 ( .A(n35145), .B(n11421), .Z(n11165) );
  AND U11688 ( .A(n11166), .B(n11165), .Z(n11307) );
  NANDN U11689 ( .A(n38247), .B(n11167), .Z(n11169) );
  XOR U11690 ( .A(b[61]), .B(a[9]), .Z(n11424) );
  NANDN U11691 ( .A(n38248), .B(n11424), .Z(n11168) );
  AND U11692 ( .A(n11169), .B(n11168), .Z(n11305) );
  AND U11693 ( .A(b[63]), .B(a[5]), .Z(n11304) );
  XNOR U11694 ( .A(n11305), .B(n11304), .Z(n11306) );
  XOR U11695 ( .A(n11307), .B(n11306), .Z(n11316) );
  XNOR U11696 ( .A(n11317), .B(n11316), .Z(n11319) );
  NANDN U11697 ( .A(n11171), .B(n11170), .Z(n11175) );
  OR U11698 ( .A(n11173), .B(n11172), .Z(n11174) );
  AND U11699 ( .A(n11175), .B(n11174), .Z(n11348) );
  NANDN U11700 ( .A(n34223), .B(n11176), .Z(n11178) );
  XOR U11701 ( .A(b[27]), .B(a[43]), .Z(n11433) );
  NANDN U11702 ( .A(n34458), .B(n11433), .Z(n11177) );
  AND U11703 ( .A(n11178), .B(n11177), .Z(n11280) );
  NANDN U11704 ( .A(n34634), .B(n11179), .Z(n11181) );
  XOR U11705 ( .A(b[29]), .B(a[41]), .Z(n11436) );
  NANDN U11706 ( .A(n34722), .B(n11436), .Z(n11180) );
  AND U11707 ( .A(n11181), .B(n11180), .Z(n11278) );
  NANDN U11708 ( .A(n31055), .B(n11182), .Z(n11184) );
  XOR U11709 ( .A(b[13]), .B(a[57]), .Z(n11439) );
  NANDN U11710 ( .A(n31293), .B(n11439), .Z(n11183) );
  NAND U11711 ( .A(n11184), .B(n11183), .Z(n11277) );
  XNOR U11712 ( .A(n11278), .B(n11277), .Z(n11279) );
  XOR U11713 ( .A(n11280), .B(n11279), .Z(n11347) );
  NANDN U11714 ( .A(n28889), .B(n11185), .Z(n11187) );
  XOR U11715 ( .A(b[5]), .B(a[65]), .Z(n11442) );
  NANDN U11716 ( .A(n29138), .B(n11442), .Z(n11186) );
  AND U11717 ( .A(n11187), .B(n11186), .Z(n11373) );
  NANDN U11718 ( .A(n209), .B(n11188), .Z(n11190) );
  XOR U11719 ( .A(b[3]), .B(a[67]), .Z(n11445) );
  NANDN U11720 ( .A(n28941), .B(n11445), .Z(n11189) );
  AND U11721 ( .A(n11190), .B(n11189), .Z(n11371) );
  NANDN U11722 ( .A(n35936), .B(n11191), .Z(n11193) );
  XOR U11723 ( .A(b[37]), .B(a[33]), .Z(n11448) );
  NANDN U11724 ( .A(n36047), .B(n11448), .Z(n11192) );
  NAND U11725 ( .A(n11193), .B(n11192), .Z(n11370) );
  XNOR U11726 ( .A(n11371), .B(n11370), .Z(n11372) );
  XOR U11727 ( .A(n11373), .B(n11372), .Z(n11346) );
  XNOR U11728 ( .A(n11347), .B(n11346), .Z(n11349) );
  XOR U11729 ( .A(n11458), .B(n11457), .Z(n11459) );
  XNOR U11730 ( .A(n11460), .B(n11459), .Z(n11243) );
  XOR U11731 ( .A(n11244), .B(n11243), .Z(n11236) );
  NANDN U11732 ( .A(n11195), .B(n11194), .Z(n11199) );
  NANDN U11733 ( .A(n11197), .B(n11196), .Z(n11198) );
  AND U11734 ( .A(n11199), .B(n11198), .Z(n11235) );
  XNOR U11735 ( .A(n11236), .B(n11235), .Z(n11237) );
  XNOR U11736 ( .A(n11238), .B(n11237), .Z(n11485) );
  XNOR U11737 ( .A(n11486), .B(n11485), .Z(n11487) );
  XOR U11738 ( .A(n11488), .B(n11487), .Z(n11500) );
  XNOR U11739 ( .A(n11499), .B(n11500), .Z(n11505) );
  NANDN U11740 ( .A(n11201), .B(n11200), .Z(n11205) );
  NANDN U11741 ( .A(n11203), .B(n11202), .Z(n11204) );
  AND U11742 ( .A(n11205), .B(n11204), .Z(n11504) );
  NANDN U11743 ( .A(n11207), .B(n11206), .Z(n11211) );
  OR U11744 ( .A(n11209), .B(n11208), .Z(n11210) );
  AND U11745 ( .A(n11211), .B(n11210), .Z(n11503) );
  XOR U11746 ( .A(n11504), .B(n11503), .Z(n11506) );
  XNOR U11747 ( .A(n11505), .B(n11506), .Z(n11229) );
  XOR U11748 ( .A(n11230), .B(n11229), .Z(n11232) );
  XOR U11749 ( .A(n11231), .B(n11232), .Z(n11224) );
  NANDN U11750 ( .A(n11213), .B(n11212), .Z(n11217) );
  NANDN U11751 ( .A(n11215), .B(n11214), .Z(n11216) );
  NAND U11752 ( .A(n11217), .B(n11216), .Z(n11223) );
  XNOR U11753 ( .A(n11224), .B(n11223), .Z(n11225) );
  XNOR U11754 ( .A(n11226), .B(n11225), .Z(n11509) );
  XNOR U11755 ( .A(sreg[133]), .B(n11509), .Z(n11511) );
  NANDN U11756 ( .A(sreg[132]), .B(n11218), .Z(n11222) );
  NAND U11757 ( .A(n11220), .B(n11219), .Z(n11221) );
  NAND U11758 ( .A(n11222), .B(n11221), .Z(n11510) );
  XNOR U11759 ( .A(n11511), .B(n11510), .Z(c[133]) );
  NANDN U11760 ( .A(n11224), .B(n11223), .Z(n11228) );
  NANDN U11761 ( .A(n11226), .B(n11225), .Z(n11227) );
  AND U11762 ( .A(n11228), .B(n11227), .Z(n11517) );
  NANDN U11763 ( .A(n11230), .B(n11229), .Z(n11234) );
  OR U11764 ( .A(n11232), .B(n11231), .Z(n11233) );
  AND U11765 ( .A(n11234), .B(n11233), .Z(n11514) );
  NANDN U11766 ( .A(n11236), .B(n11235), .Z(n11240) );
  NANDN U11767 ( .A(n11238), .B(n11237), .Z(n11239) );
  AND U11768 ( .A(n11240), .B(n11239), .Z(n11534) );
  NANDN U11769 ( .A(n11242), .B(n11241), .Z(n11246) );
  NAND U11770 ( .A(n11244), .B(n11243), .Z(n11245) );
  AND U11771 ( .A(n11246), .B(n11245), .Z(n11546) );
  NANDN U11772 ( .A(n11248), .B(n11247), .Z(n11252) );
  NANDN U11773 ( .A(n11250), .B(n11249), .Z(n11251) );
  AND U11774 ( .A(n11252), .B(n11251), .Z(n11558) );
  NAND U11775 ( .A(n11254), .B(n11253), .Z(n11258) );
  NAND U11776 ( .A(n11256), .B(n11255), .Z(n11257) );
  AND U11777 ( .A(n11258), .B(n11257), .Z(n11557) );
  NANDN U11778 ( .A(n33875), .B(n11259), .Z(n11261) );
  XOR U11779 ( .A(b[25]), .B(a[46]), .Z(n11592) );
  NANDN U11780 ( .A(n33994), .B(n11592), .Z(n11260) );
  AND U11781 ( .A(n11261), .B(n11260), .Z(n11720) );
  NANDN U11782 ( .A(n32013), .B(n11262), .Z(n11264) );
  XOR U11783 ( .A(b[17]), .B(a[54]), .Z(n11595) );
  NANDN U11784 ( .A(n32292), .B(n11595), .Z(n11263) );
  AND U11785 ( .A(n11264), .B(n11263), .Z(n11719) );
  NANDN U11786 ( .A(n31536), .B(n11265), .Z(n11267) );
  XOR U11787 ( .A(b[15]), .B(a[56]), .Z(n11598) );
  NANDN U11788 ( .A(n31925), .B(n11598), .Z(n11266) );
  NAND U11789 ( .A(n11267), .B(n11266), .Z(n11718) );
  XOR U11790 ( .A(n11719), .B(n11718), .Z(n11721) );
  XOR U11791 ( .A(n11720), .B(n11721), .Z(n11785) );
  NANDN U11792 ( .A(n37526), .B(n11268), .Z(n11270) );
  XOR U11793 ( .A(b[51]), .B(a[20]), .Z(n11601) );
  NANDN U11794 ( .A(n37605), .B(n11601), .Z(n11269) );
  AND U11795 ( .A(n11270), .B(n11269), .Z(n11744) );
  NANDN U11796 ( .A(n37705), .B(n11271), .Z(n11273) );
  XOR U11797 ( .A(b[53]), .B(a[18]), .Z(n11604) );
  NANDN U11798 ( .A(n37778), .B(n11604), .Z(n11272) );
  AND U11799 ( .A(n11273), .B(n11272), .Z(n11743) );
  NANDN U11800 ( .A(n36210), .B(n11274), .Z(n11276) );
  XOR U11801 ( .A(b[39]), .B(a[32]), .Z(n11607) );
  NANDN U11802 ( .A(n36347), .B(n11607), .Z(n11275) );
  NAND U11803 ( .A(n11276), .B(n11275), .Z(n11742) );
  XOR U11804 ( .A(n11743), .B(n11742), .Z(n11745) );
  XNOR U11805 ( .A(n11744), .B(n11745), .Z(n11784) );
  XNOR U11806 ( .A(n11785), .B(n11784), .Z(n11787) );
  NANDN U11807 ( .A(n11278), .B(n11277), .Z(n11282) );
  NANDN U11808 ( .A(n11280), .B(n11279), .Z(n11281) );
  AND U11809 ( .A(n11282), .B(n11281), .Z(n11786) );
  XOR U11810 ( .A(n11787), .B(n11786), .Z(n11583) );
  NANDN U11811 ( .A(n11284), .B(n11283), .Z(n11288) );
  OR U11812 ( .A(n11286), .B(n11285), .Z(n11287) );
  AND U11813 ( .A(n11288), .B(n11287), .Z(n11581) );
  NANDN U11814 ( .A(n11290), .B(n11289), .Z(n11294) );
  NANDN U11815 ( .A(n11292), .B(n11291), .Z(n11293) );
  NAND U11816 ( .A(n11294), .B(n11293), .Z(n11580) );
  XNOR U11817 ( .A(n11581), .B(n11580), .Z(n11582) );
  XNOR U11818 ( .A(n11583), .B(n11582), .Z(n11556) );
  XOR U11819 ( .A(n11557), .B(n11556), .Z(n11559) );
  XOR U11820 ( .A(n11558), .B(n11559), .Z(n11545) );
  NANDN U11821 ( .A(n29499), .B(n11295), .Z(n11297) );
  XOR U11822 ( .A(b[7]), .B(a[64]), .Z(n11628) );
  NANDN U11823 ( .A(n29735), .B(n11628), .Z(n11296) );
  AND U11824 ( .A(n11297), .B(n11296), .Z(n11618) );
  NANDN U11825 ( .A(n37857), .B(n11298), .Z(n11300) );
  XOR U11826 ( .A(b[55]), .B(a[16]), .Z(n11631) );
  NANDN U11827 ( .A(n37911), .B(n11631), .Z(n11299) );
  AND U11828 ( .A(n11300), .B(n11299), .Z(n11617) );
  NANDN U11829 ( .A(n35611), .B(n11301), .Z(n11303) );
  XOR U11830 ( .A(b[35]), .B(a[36]), .Z(n11634) );
  NANDN U11831 ( .A(n35801), .B(n11634), .Z(n11302) );
  NAND U11832 ( .A(n11303), .B(n11302), .Z(n11616) );
  XOR U11833 ( .A(n11617), .B(n11616), .Z(n11619) );
  XOR U11834 ( .A(n11618), .B(n11619), .Z(n11680) );
  NANDN U11835 ( .A(n11305), .B(n11304), .Z(n11309) );
  NANDN U11836 ( .A(n11307), .B(n11306), .Z(n11308) );
  AND U11837 ( .A(n11309), .B(n11308), .Z(n11679) );
  XNOR U11838 ( .A(n11680), .B(n11679), .Z(n11681) );
  NANDN U11839 ( .A(n11311), .B(n11310), .Z(n11315) );
  OR U11840 ( .A(n11313), .B(n11312), .Z(n11314) );
  NAND U11841 ( .A(n11315), .B(n11314), .Z(n11682) );
  XNOR U11842 ( .A(n11681), .B(n11682), .Z(n11564) );
  NAND U11843 ( .A(n11317), .B(n11316), .Z(n11321) );
  NANDN U11844 ( .A(n11319), .B(n11318), .Z(n11320) );
  AND U11845 ( .A(n11321), .B(n11320), .Z(n11563) );
  NANDN U11846 ( .A(n211), .B(n11322), .Z(n11324) );
  XOR U11847 ( .A(b[47]), .B(a[24]), .Z(n11655) );
  NANDN U11848 ( .A(n37172), .B(n11655), .Z(n11323) );
  AND U11849 ( .A(n11324), .B(n11323), .Z(n11645) );
  NANDN U11850 ( .A(n210), .B(n11325), .Z(n11327) );
  XOR U11851 ( .A(b[9]), .B(a[62]), .Z(n11658) );
  NANDN U11852 ( .A(n30267), .B(n11658), .Z(n11326) );
  AND U11853 ( .A(n11327), .B(n11326), .Z(n11644) );
  NANDN U11854 ( .A(n212), .B(n11328), .Z(n11330) );
  XOR U11855 ( .A(b[49]), .B(a[22]), .Z(n11661) );
  NANDN U11856 ( .A(n37432), .B(n11661), .Z(n11329) );
  NAND U11857 ( .A(n11330), .B(n11329), .Z(n11643) );
  XOR U11858 ( .A(n11644), .B(n11643), .Z(n11646) );
  XOR U11859 ( .A(n11645), .B(n11646), .Z(n11698) );
  NANDN U11860 ( .A(n36742), .B(n11331), .Z(n11333) );
  XOR U11861 ( .A(b[43]), .B(a[28]), .Z(n11664) );
  NANDN U11862 ( .A(n36891), .B(n11664), .Z(n11332) );
  AND U11863 ( .A(n11333), .B(n11332), .Z(n11675) );
  NANDN U11864 ( .A(n36991), .B(n11334), .Z(n11336) );
  XOR U11865 ( .A(b[45]), .B(a[26]), .Z(n11667) );
  NANDN U11866 ( .A(n37083), .B(n11667), .Z(n11335) );
  AND U11867 ( .A(n11336), .B(n11335), .Z(n11674) );
  NANDN U11868 ( .A(n30482), .B(n11337), .Z(n11339) );
  XOR U11869 ( .A(b[11]), .B(a[60]), .Z(n11670) );
  NANDN U11870 ( .A(n30891), .B(n11670), .Z(n11338) );
  NAND U11871 ( .A(n11339), .B(n11338), .Z(n11673) );
  XOR U11872 ( .A(n11674), .B(n11673), .Z(n11676) );
  XNOR U11873 ( .A(n11675), .B(n11676), .Z(n11697) );
  XNOR U11874 ( .A(n11698), .B(n11697), .Z(n11699) );
  NANDN U11875 ( .A(n11341), .B(n11340), .Z(n11345) );
  OR U11876 ( .A(n11343), .B(n11342), .Z(n11344) );
  NAND U11877 ( .A(n11345), .B(n11344), .Z(n11700) );
  XNOR U11878 ( .A(n11699), .B(n11700), .Z(n11562) );
  XOR U11879 ( .A(n11563), .B(n11562), .Z(n11565) );
  XNOR U11880 ( .A(n11564), .B(n11565), .Z(n11544) );
  XOR U11881 ( .A(n11545), .B(n11544), .Z(n11547) );
  XOR U11882 ( .A(n11546), .B(n11547), .Z(n11533) );
  NAND U11883 ( .A(n11347), .B(n11346), .Z(n11351) );
  NANDN U11884 ( .A(n11349), .B(n11348), .Z(n11350) );
  NAND U11885 ( .A(n11351), .B(n11350), .Z(n11550) );
  NANDN U11886 ( .A(n11353), .B(n11352), .Z(n11357) );
  NAND U11887 ( .A(n11355), .B(n11354), .Z(n11356) );
  AND U11888 ( .A(n11357), .B(n11356), .Z(n11551) );
  XOR U11889 ( .A(n11550), .B(n11551), .Z(n11553) );
  NANDN U11890 ( .A(n11359), .B(n11358), .Z(n11363) );
  NANDN U11891 ( .A(n11361), .B(n11360), .Z(n11362) );
  NAND U11892 ( .A(n11363), .B(n11362), .Z(n11552) );
  XOR U11893 ( .A(n11553), .B(n11552), .Z(n11571) );
  NANDN U11894 ( .A(n11365), .B(n11364), .Z(n11369) );
  OR U11895 ( .A(n11367), .B(n11366), .Z(n11368) );
  AND U11896 ( .A(n11369), .B(n11368), .Z(n11692) );
  NANDN U11897 ( .A(n11371), .B(n11370), .Z(n11375) );
  NANDN U11898 ( .A(n11373), .B(n11372), .Z(n11374) );
  NAND U11899 ( .A(n11375), .B(n11374), .Z(n11691) );
  XNOR U11900 ( .A(n11692), .B(n11691), .Z(n11694) );
  NANDN U11901 ( .A(n11377), .B(n11376), .Z(n11381) );
  NANDN U11902 ( .A(n11379), .B(n11378), .Z(n11380) );
  AND U11903 ( .A(n11381), .B(n11380), .Z(n11589) );
  NAND U11904 ( .A(b[0]), .B(a[70]), .Z(n11382) );
  XNOR U11905 ( .A(b[1]), .B(n11382), .Z(n11384) );
  NANDN U11906 ( .A(b[0]), .B(a[69]), .Z(n11383) );
  NAND U11907 ( .A(n11384), .B(n11383), .Z(n11625) );
  NANDN U11908 ( .A(n38278), .B(n11385), .Z(n11387) );
  XOR U11909 ( .A(b[63]), .B(a[8]), .Z(n11769) );
  NANDN U11910 ( .A(n38279), .B(n11769), .Z(n11386) );
  AND U11911 ( .A(n11387), .B(n11386), .Z(n11623) );
  NANDN U11912 ( .A(n35260), .B(n11388), .Z(n11390) );
  XOR U11913 ( .A(b[33]), .B(a[38]), .Z(n11772) );
  NANDN U11914 ( .A(n35456), .B(n11772), .Z(n11389) );
  NAND U11915 ( .A(n11390), .B(n11389), .Z(n11622) );
  XNOR U11916 ( .A(n11623), .B(n11622), .Z(n11624) );
  XNOR U11917 ( .A(n11625), .B(n11624), .Z(n11586) );
  NANDN U11918 ( .A(n37974), .B(n11391), .Z(n11393) );
  XOR U11919 ( .A(b[57]), .B(a[14]), .Z(n11775) );
  NANDN U11920 ( .A(n38031), .B(n11775), .Z(n11392) );
  AND U11921 ( .A(n11393), .B(n11392), .Z(n11751) );
  NANDN U11922 ( .A(n38090), .B(n11394), .Z(n11396) );
  XOR U11923 ( .A(b[59]), .B(a[12]), .Z(n11778) );
  NANDN U11924 ( .A(n38130), .B(n11778), .Z(n11395) );
  AND U11925 ( .A(n11396), .B(n11395), .Z(n11749) );
  NANDN U11926 ( .A(n36480), .B(n11397), .Z(n11399) );
  XOR U11927 ( .A(b[41]), .B(a[30]), .Z(n11781) );
  NANDN U11928 ( .A(n36594), .B(n11781), .Z(n11398) );
  NAND U11929 ( .A(n11399), .B(n11398), .Z(n11748) );
  XNOR U11930 ( .A(n11749), .B(n11748), .Z(n11750) );
  XOR U11931 ( .A(n11751), .B(n11750), .Z(n11587) );
  XNOR U11932 ( .A(n11586), .B(n11587), .Z(n11588) );
  XNOR U11933 ( .A(n11589), .B(n11588), .Z(n11693) );
  XOR U11934 ( .A(n11694), .B(n11693), .Z(n11575) );
  NANDN U11935 ( .A(n11401), .B(n11400), .Z(n11405) );
  NAND U11936 ( .A(n11403), .B(n11402), .Z(n11404) );
  NAND U11937 ( .A(n11405), .B(n11404), .Z(n11574) );
  XNOR U11938 ( .A(n11575), .B(n11574), .Z(n11577) );
  NANDN U11939 ( .A(n11407), .B(n11406), .Z(n11411) );
  NANDN U11940 ( .A(n11409), .B(n11408), .Z(n11410) );
  AND U11941 ( .A(n11411), .B(n11410), .Z(n11793) );
  NANDN U11942 ( .A(n32996), .B(n11412), .Z(n11414) );
  XOR U11943 ( .A(b[21]), .B(a[50]), .Z(n11703) );
  NANDN U11944 ( .A(n33271), .B(n11703), .Z(n11413) );
  AND U11945 ( .A(n11414), .B(n11413), .Z(n11762) );
  NANDN U11946 ( .A(n33866), .B(n11415), .Z(n11417) );
  XOR U11947 ( .A(b[23]), .B(a[48]), .Z(n11706) );
  NANDN U11948 ( .A(n33644), .B(n11706), .Z(n11416) );
  AND U11949 ( .A(n11417), .B(n11416), .Z(n11761) );
  NANDN U11950 ( .A(n32483), .B(n11418), .Z(n11420) );
  XOR U11951 ( .A(b[19]), .B(a[52]), .Z(n11709) );
  NANDN U11952 ( .A(n32823), .B(n11709), .Z(n11419) );
  NAND U11953 ( .A(n11420), .B(n11419), .Z(n11760) );
  XOR U11954 ( .A(n11761), .B(n11760), .Z(n11763) );
  XOR U11955 ( .A(n11762), .B(n11763), .Z(n11650) );
  NANDN U11956 ( .A(n34909), .B(n11421), .Z(n11423) );
  XOR U11957 ( .A(b[31]), .B(a[40]), .Z(n11712) );
  NANDN U11958 ( .A(n35145), .B(n11712), .Z(n11422) );
  AND U11959 ( .A(n11423), .B(n11422), .Z(n11639) );
  NANDN U11960 ( .A(n38247), .B(n11424), .Z(n11426) );
  XOR U11961 ( .A(b[61]), .B(a[10]), .Z(n11715) );
  NANDN U11962 ( .A(n38248), .B(n11715), .Z(n11425) );
  AND U11963 ( .A(n11426), .B(n11425), .Z(n11638) );
  AND U11964 ( .A(b[63]), .B(a[6]), .Z(n11637) );
  XOR U11965 ( .A(n11638), .B(n11637), .Z(n11640) );
  XNOR U11966 ( .A(n11639), .B(n11640), .Z(n11649) );
  XNOR U11967 ( .A(n11650), .B(n11649), .Z(n11651) );
  NANDN U11968 ( .A(n11428), .B(n11427), .Z(n11432) );
  OR U11969 ( .A(n11430), .B(n11429), .Z(n11431) );
  NAND U11970 ( .A(n11432), .B(n11431), .Z(n11652) );
  XNOR U11971 ( .A(n11651), .B(n11652), .Z(n11790) );
  NANDN U11972 ( .A(n34223), .B(n11433), .Z(n11435) );
  XOR U11973 ( .A(b[27]), .B(a[44]), .Z(n11724) );
  NANDN U11974 ( .A(n34458), .B(n11724), .Z(n11434) );
  AND U11975 ( .A(n11435), .B(n11434), .Z(n11612) );
  NANDN U11976 ( .A(n34634), .B(n11436), .Z(n11438) );
  XOR U11977 ( .A(b[29]), .B(a[42]), .Z(n11727) );
  NANDN U11978 ( .A(n34722), .B(n11727), .Z(n11437) );
  AND U11979 ( .A(n11438), .B(n11437), .Z(n11611) );
  NANDN U11980 ( .A(n31055), .B(n11439), .Z(n11441) );
  XOR U11981 ( .A(b[13]), .B(a[58]), .Z(n11730) );
  NANDN U11982 ( .A(n31293), .B(n11730), .Z(n11440) );
  NAND U11983 ( .A(n11441), .B(n11440), .Z(n11610) );
  XOR U11984 ( .A(n11611), .B(n11610), .Z(n11613) );
  XOR U11985 ( .A(n11612), .B(n11613), .Z(n11686) );
  NANDN U11986 ( .A(n28889), .B(n11442), .Z(n11444) );
  XOR U11987 ( .A(b[5]), .B(a[66]), .Z(n11733) );
  NANDN U11988 ( .A(n29138), .B(n11733), .Z(n11443) );
  AND U11989 ( .A(n11444), .B(n11443), .Z(n11756) );
  NANDN U11990 ( .A(n209), .B(n11445), .Z(n11447) );
  XOR U11991 ( .A(b[3]), .B(a[68]), .Z(n11736) );
  NANDN U11992 ( .A(n28941), .B(n11736), .Z(n11446) );
  AND U11993 ( .A(n11447), .B(n11446), .Z(n11755) );
  NANDN U11994 ( .A(n35936), .B(n11448), .Z(n11450) );
  XOR U11995 ( .A(b[37]), .B(a[34]), .Z(n11739) );
  NANDN U11996 ( .A(n36047), .B(n11739), .Z(n11449) );
  NAND U11997 ( .A(n11450), .B(n11449), .Z(n11754) );
  XOR U11998 ( .A(n11755), .B(n11754), .Z(n11757) );
  XNOR U11999 ( .A(n11756), .B(n11757), .Z(n11685) );
  XNOR U12000 ( .A(n11686), .B(n11685), .Z(n11687) );
  NANDN U12001 ( .A(n11452), .B(n11451), .Z(n11456) );
  OR U12002 ( .A(n11454), .B(n11453), .Z(n11455) );
  NAND U12003 ( .A(n11456), .B(n11455), .Z(n11688) );
  XOR U12004 ( .A(n11687), .B(n11688), .Z(n11791) );
  XNOR U12005 ( .A(n11790), .B(n11791), .Z(n11792) );
  XNOR U12006 ( .A(n11793), .B(n11792), .Z(n11576) );
  XOR U12007 ( .A(n11577), .B(n11576), .Z(n11569) );
  XNOR U12008 ( .A(n11569), .B(n11568), .Z(n11570) );
  XNOR U12009 ( .A(n11571), .B(n11570), .Z(n11532) );
  XOR U12010 ( .A(n11533), .B(n11532), .Z(n11535) );
  XOR U12011 ( .A(n11534), .B(n11535), .Z(n11528) );
  NANDN U12012 ( .A(n11462), .B(n11461), .Z(n11466) );
  OR U12013 ( .A(n11464), .B(n11463), .Z(n11465) );
  AND U12014 ( .A(n11466), .B(n11465), .Z(n11527) );
  NANDN U12015 ( .A(n11468), .B(n11467), .Z(n11472) );
  OR U12016 ( .A(n11470), .B(n11469), .Z(n11471) );
  AND U12017 ( .A(n11472), .B(n11471), .Z(n11541) );
  NANDN U12018 ( .A(n11474), .B(n11473), .Z(n11478) );
  NANDN U12019 ( .A(n11476), .B(n11475), .Z(n11477) );
  AND U12020 ( .A(n11478), .B(n11477), .Z(n11539) );
  NANDN U12021 ( .A(n11480), .B(n11479), .Z(n11484) );
  OR U12022 ( .A(n11482), .B(n11481), .Z(n11483) );
  AND U12023 ( .A(n11484), .B(n11483), .Z(n11538) );
  XNOR U12024 ( .A(n11539), .B(n11538), .Z(n11540) );
  XNOR U12025 ( .A(n11541), .B(n11540), .Z(n11526) );
  XOR U12026 ( .A(n11527), .B(n11526), .Z(n11529) );
  XOR U12027 ( .A(n11528), .B(n11529), .Z(n11522) );
  NANDN U12028 ( .A(n11486), .B(n11485), .Z(n11490) );
  NANDN U12029 ( .A(n11488), .B(n11487), .Z(n11489) );
  AND U12030 ( .A(n11490), .B(n11489), .Z(n11521) );
  NANDN U12031 ( .A(n11492), .B(n11491), .Z(n11496) );
  OR U12032 ( .A(n11494), .B(n11493), .Z(n11495) );
  AND U12033 ( .A(n11496), .B(n11495), .Z(n11520) );
  XOR U12034 ( .A(n11521), .B(n11520), .Z(n11523) );
  XOR U12035 ( .A(n11522), .B(n11523), .Z(n11797) );
  NANDN U12036 ( .A(n11498), .B(n11497), .Z(n11502) );
  NANDN U12037 ( .A(n11500), .B(n11499), .Z(n11501) );
  AND U12038 ( .A(n11502), .B(n11501), .Z(n11796) );
  XNOR U12039 ( .A(n11797), .B(n11796), .Z(n11798) );
  NANDN U12040 ( .A(n11504), .B(n11503), .Z(n11508) );
  NANDN U12041 ( .A(n11506), .B(n11505), .Z(n11507) );
  NAND U12042 ( .A(n11508), .B(n11507), .Z(n11799) );
  XOR U12043 ( .A(n11798), .B(n11799), .Z(n11515) );
  XNOR U12044 ( .A(n11514), .B(n11515), .Z(n11516) );
  XNOR U12045 ( .A(n11517), .B(n11516), .Z(n11802) );
  XNOR U12046 ( .A(sreg[134]), .B(n11802), .Z(n11804) );
  NANDN U12047 ( .A(sreg[133]), .B(n11509), .Z(n11513) );
  NAND U12048 ( .A(n11511), .B(n11510), .Z(n11512) );
  NAND U12049 ( .A(n11513), .B(n11512), .Z(n11803) );
  XNOR U12050 ( .A(n11804), .B(n11803), .Z(c[134]) );
  NANDN U12051 ( .A(n11515), .B(n11514), .Z(n11519) );
  NANDN U12052 ( .A(n11517), .B(n11516), .Z(n11518) );
  AND U12053 ( .A(n11519), .B(n11518), .Z(n11810) );
  NANDN U12054 ( .A(n11521), .B(n11520), .Z(n11525) );
  OR U12055 ( .A(n11523), .B(n11522), .Z(n11524) );
  AND U12056 ( .A(n11525), .B(n11524), .Z(n11815) );
  NANDN U12057 ( .A(n11527), .B(n11526), .Z(n11531) );
  OR U12058 ( .A(n11529), .B(n11528), .Z(n11530) );
  AND U12059 ( .A(n11531), .B(n11530), .Z(n11813) );
  NANDN U12060 ( .A(n11533), .B(n11532), .Z(n11537) );
  OR U12061 ( .A(n11535), .B(n11534), .Z(n11536) );
  AND U12062 ( .A(n11537), .B(n11536), .Z(n12090) );
  NANDN U12063 ( .A(n11539), .B(n11538), .Z(n11543) );
  NANDN U12064 ( .A(n11541), .B(n11540), .Z(n11542) );
  AND U12065 ( .A(n11543), .B(n11542), .Z(n12089) );
  XNOR U12066 ( .A(n12090), .B(n12089), .Z(n12091) );
  NANDN U12067 ( .A(n11545), .B(n11544), .Z(n11549) );
  OR U12068 ( .A(n11547), .B(n11546), .Z(n11548) );
  AND U12069 ( .A(n11549), .B(n11548), .Z(n12083) );
  NAND U12070 ( .A(n11551), .B(n11550), .Z(n11555) );
  NAND U12071 ( .A(n11553), .B(n11552), .Z(n11554) );
  AND U12072 ( .A(n11555), .B(n11554), .Z(n11827) );
  NANDN U12073 ( .A(n11557), .B(n11556), .Z(n11561) );
  OR U12074 ( .A(n11559), .B(n11558), .Z(n11560) );
  AND U12075 ( .A(n11561), .B(n11560), .Z(n11826) );
  NANDN U12076 ( .A(n11563), .B(n11562), .Z(n11567) );
  NANDN U12077 ( .A(n11565), .B(n11564), .Z(n11566) );
  AND U12078 ( .A(n11567), .B(n11566), .Z(n11825) );
  XOR U12079 ( .A(n11826), .B(n11825), .Z(n11828) );
  XOR U12080 ( .A(n11827), .B(n11828), .Z(n12084) );
  XNOR U12081 ( .A(n12083), .B(n12084), .Z(n12085) );
  NANDN U12082 ( .A(n11569), .B(n11568), .Z(n11573) );
  NANDN U12083 ( .A(n11571), .B(n11570), .Z(n11572) );
  AND U12084 ( .A(n11573), .B(n11572), .Z(n11822) );
  NANDN U12085 ( .A(n11575), .B(n11574), .Z(n11579) );
  NAND U12086 ( .A(n11577), .B(n11576), .Z(n11578) );
  AND U12087 ( .A(n11579), .B(n11578), .Z(n11851) );
  NANDN U12088 ( .A(n11581), .B(n11580), .Z(n11585) );
  NANDN U12089 ( .A(n11583), .B(n11582), .Z(n11584) );
  AND U12090 ( .A(n11585), .B(n11584), .Z(n11845) );
  NANDN U12091 ( .A(n11587), .B(n11586), .Z(n11591) );
  NANDN U12092 ( .A(n11589), .B(n11588), .Z(n11590) );
  AND U12093 ( .A(n11591), .B(n11590), .Z(n11844) );
  NANDN U12094 ( .A(n33875), .B(n11592), .Z(n11594) );
  XOR U12095 ( .A(b[25]), .B(a[47]), .Z(n11924) );
  NANDN U12096 ( .A(n33994), .B(n11924), .Z(n11593) );
  AND U12097 ( .A(n11594), .B(n11593), .Z(n12049) );
  NANDN U12098 ( .A(n32013), .B(n11595), .Z(n11597) );
  XOR U12099 ( .A(b[17]), .B(a[55]), .Z(n11927) );
  NANDN U12100 ( .A(n32292), .B(n11927), .Z(n11596) );
  AND U12101 ( .A(n11597), .B(n11596), .Z(n12048) );
  NANDN U12102 ( .A(n31536), .B(n11598), .Z(n11600) );
  XOR U12103 ( .A(b[15]), .B(a[57]), .Z(n11930) );
  NANDN U12104 ( .A(n31925), .B(n11930), .Z(n11599) );
  NAND U12105 ( .A(n11600), .B(n11599), .Z(n12047) );
  XOR U12106 ( .A(n12048), .B(n12047), .Z(n12050) );
  XOR U12107 ( .A(n12049), .B(n12050), .Z(n12021) );
  NANDN U12108 ( .A(n37526), .B(n11601), .Z(n11603) );
  XOR U12109 ( .A(b[51]), .B(a[21]), .Z(n11933) );
  NANDN U12110 ( .A(n37605), .B(n11933), .Z(n11602) );
  AND U12111 ( .A(n11603), .B(n11602), .Z(n12073) );
  NANDN U12112 ( .A(n37705), .B(n11604), .Z(n11606) );
  XOR U12113 ( .A(b[53]), .B(a[19]), .Z(n11936) );
  NANDN U12114 ( .A(n37778), .B(n11936), .Z(n11605) );
  AND U12115 ( .A(n11606), .B(n11605), .Z(n12072) );
  NANDN U12116 ( .A(n36210), .B(n11607), .Z(n11609) );
  XOR U12117 ( .A(b[39]), .B(a[33]), .Z(n11939) );
  NANDN U12118 ( .A(n36347), .B(n11939), .Z(n11608) );
  NAND U12119 ( .A(n11609), .B(n11608), .Z(n12071) );
  XOR U12120 ( .A(n12072), .B(n12071), .Z(n12074) );
  XNOR U12121 ( .A(n12073), .B(n12074), .Z(n12020) );
  XNOR U12122 ( .A(n12021), .B(n12020), .Z(n12023) );
  NANDN U12123 ( .A(n11611), .B(n11610), .Z(n11615) );
  OR U12124 ( .A(n11613), .B(n11612), .Z(n11614) );
  AND U12125 ( .A(n11615), .B(n11614), .Z(n12022) );
  XOR U12126 ( .A(n12023), .B(n12022), .Z(n11915) );
  NANDN U12127 ( .A(n11617), .B(n11616), .Z(n11621) );
  OR U12128 ( .A(n11619), .B(n11618), .Z(n11620) );
  AND U12129 ( .A(n11621), .B(n11620), .Z(n11913) );
  NANDN U12130 ( .A(n11623), .B(n11622), .Z(n11627) );
  NANDN U12131 ( .A(n11625), .B(n11624), .Z(n11626) );
  NAND U12132 ( .A(n11627), .B(n11626), .Z(n11912) );
  XNOR U12133 ( .A(n11913), .B(n11912), .Z(n11914) );
  XNOR U12134 ( .A(n11915), .B(n11914), .Z(n11843) );
  XOR U12135 ( .A(n11844), .B(n11843), .Z(n11846) );
  XOR U12136 ( .A(n11845), .B(n11846), .Z(n11850) );
  NANDN U12137 ( .A(n29499), .B(n11628), .Z(n11630) );
  XOR U12138 ( .A(b[7]), .B(a[65]), .Z(n11861) );
  NANDN U12139 ( .A(n29735), .B(n11861), .Z(n11629) );
  AND U12140 ( .A(n11630), .B(n11629), .Z(n11950) );
  NANDN U12141 ( .A(n37857), .B(n11631), .Z(n11633) );
  XOR U12142 ( .A(b[55]), .B(a[17]), .Z(n11864) );
  NANDN U12143 ( .A(n37911), .B(n11864), .Z(n11632) );
  AND U12144 ( .A(n11633), .B(n11632), .Z(n11949) );
  NANDN U12145 ( .A(n35611), .B(n11634), .Z(n11636) );
  XOR U12146 ( .A(b[35]), .B(a[37]), .Z(n11867) );
  NANDN U12147 ( .A(n35801), .B(n11867), .Z(n11635) );
  NAND U12148 ( .A(n11636), .B(n11635), .Z(n11948) );
  XOR U12149 ( .A(n11949), .B(n11948), .Z(n11951) );
  XOR U12150 ( .A(n11950), .B(n11951), .Z(n11967) );
  NANDN U12151 ( .A(n11638), .B(n11637), .Z(n11642) );
  OR U12152 ( .A(n11640), .B(n11639), .Z(n11641) );
  AND U12153 ( .A(n11642), .B(n11641), .Z(n11966) );
  XNOR U12154 ( .A(n11967), .B(n11966), .Z(n11968) );
  NANDN U12155 ( .A(n11644), .B(n11643), .Z(n11648) );
  OR U12156 ( .A(n11646), .B(n11645), .Z(n11647) );
  NAND U12157 ( .A(n11648), .B(n11647), .Z(n11969) );
  XNOR U12158 ( .A(n11968), .B(n11969), .Z(n11839) );
  NANDN U12159 ( .A(n11650), .B(n11649), .Z(n11654) );
  NANDN U12160 ( .A(n11652), .B(n11651), .Z(n11653) );
  AND U12161 ( .A(n11654), .B(n11653), .Z(n11838) );
  NANDN U12162 ( .A(n211), .B(n11655), .Z(n11657) );
  XOR U12163 ( .A(b[47]), .B(a[25]), .Z(n11888) );
  NANDN U12164 ( .A(n37172), .B(n11888), .Z(n11656) );
  AND U12165 ( .A(n11657), .B(n11656), .Z(n11878) );
  NANDN U12166 ( .A(n210), .B(n11658), .Z(n11660) );
  XOR U12167 ( .A(b[9]), .B(a[63]), .Z(n11891) );
  NANDN U12168 ( .A(n30267), .B(n11891), .Z(n11659) );
  AND U12169 ( .A(n11660), .B(n11659), .Z(n11877) );
  NANDN U12170 ( .A(n212), .B(n11661), .Z(n11663) );
  XOR U12171 ( .A(b[49]), .B(a[23]), .Z(n11894) );
  NANDN U12172 ( .A(n37432), .B(n11894), .Z(n11662) );
  NAND U12173 ( .A(n11663), .B(n11662), .Z(n11876) );
  XOR U12174 ( .A(n11877), .B(n11876), .Z(n11879) );
  XOR U12175 ( .A(n11878), .B(n11879), .Z(n12027) );
  NANDN U12176 ( .A(n36742), .B(n11664), .Z(n11666) );
  XOR U12177 ( .A(b[43]), .B(a[29]), .Z(n11897) );
  NANDN U12178 ( .A(n36891), .B(n11897), .Z(n11665) );
  AND U12179 ( .A(n11666), .B(n11665), .Z(n11908) );
  NANDN U12180 ( .A(n36991), .B(n11667), .Z(n11669) );
  XOR U12181 ( .A(b[45]), .B(a[27]), .Z(n11900) );
  NANDN U12182 ( .A(n37083), .B(n11900), .Z(n11668) );
  AND U12183 ( .A(n11669), .B(n11668), .Z(n11907) );
  NANDN U12184 ( .A(n30482), .B(n11670), .Z(n11672) );
  XOR U12185 ( .A(b[11]), .B(a[61]), .Z(n11903) );
  NANDN U12186 ( .A(n30891), .B(n11903), .Z(n11671) );
  NAND U12187 ( .A(n11672), .B(n11671), .Z(n11906) );
  XOR U12188 ( .A(n11907), .B(n11906), .Z(n11909) );
  XNOR U12189 ( .A(n11908), .B(n11909), .Z(n12026) );
  XNOR U12190 ( .A(n12027), .B(n12026), .Z(n12028) );
  NANDN U12191 ( .A(n11674), .B(n11673), .Z(n11678) );
  OR U12192 ( .A(n11676), .B(n11675), .Z(n11677) );
  NAND U12193 ( .A(n11678), .B(n11677), .Z(n12029) );
  XNOR U12194 ( .A(n12028), .B(n12029), .Z(n11837) );
  XOR U12195 ( .A(n11838), .B(n11837), .Z(n11840) );
  XNOR U12196 ( .A(n11839), .B(n11840), .Z(n11849) );
  XOR U12197 ( .A(n11850), .B(n11849), .Z(n11852) );
  XOR U12198 ( .A(n11851), .B(n11852), .Z(n11820) );
  NANDN U12199 ( .A(n11680), .B(n11679), .Z(n11684) );
  NANDN U12200 ( .A(n11682), .B(n11681), .Z(n11683) );
  AND U12201 ( .A(n11684), .B(n11683), .Z(n11833) );
  NANDN U12202 ( .A(n11686), .B(n11685), .Z(n11690) );
  NANDN U12203 ( .A(n11688), .B(n11687), .Z(n11689) );
  AND U12204 ( .A(n11690), .B(n11689), .Z(n11832) );
  NANDN U12205 ( .A(n11692), .B(n11691), .Z(n11696) );
  NAND U12206 ( .A(n11694), .B(n11693), .Z(n11695) );
  AND U12207 ( .A(n11696), .B(n11695), .Z(n11831) );
  XOR U12208 ( .A(n11832), .B(n11831), .Z(n11834) );
  XOR U12209 ( .A(n11833), .B(n11834), .Z(n11858) );
  NANDN U12210 ( .A(n11698), .B(n11697), .Z(n11702) );
  NANDN U12211 ( .A(n11700), .B(n11699), .Z(n11701) );
  AND U12212 ( .A(n11702), .B(n11701), .Z(n12080) );
  NANDN U12213 ( .A(n32996), .B(n11703), .Z(n11705) );
  XOR U12214 ( .A(b[21]), .B(a[51]), .Z(n12032) );
  NANDN U12215 ( .A(n33271), .B(n12032), .Z(n11704) );
  AND U12216 ( .A(n11705), .B(n11704), .Z(n11998) );
  NANDN U12217 ( .A(n33866), .B(n11706), .Z(n11708) );
  XOR U12218 ( .A(b[23]), .B(a[49]), .Z(n12035) );
  NANDN U12219 ( .A(n33644), .B(n12035), .Z(n11707) );
  AND U12220 ( .A(n11708), .B(n11707), .Z(n11997) );
  NANDN U12221 ( .A(n32483), .B(n11709), .Z(n11711) );
  XOR U12222 ( .A(b[19]), .B(a[53]), .Z(n12038) );
  NANDN U12223 ( .A(n32823), .B(n12038), .Z(n11710) );
  NAND U12224 ( .A(n11711), .B(n11710), .Z(n11996) );
  XOR U12225 ( .A(n11997), .B(n11996), .Z(n11999) );
  XOR U12226 ( .A(n11998), .B(n11999), .Z(n11883) );
  NANDN U12227 ( .A(n34909), .B(n11712), .Z(n11714) );
  XOR U12228 ( .A(b[31]), .B(a[41]), .Z(n12041) );
  NANDN U12229 ( .A(n35145), .B(n12041), .Z(n11713) );
  AND U12230 ( .A(n11714), .B(n11713), .Z(n11872) );
  NANDN U12231 ( .A(n38247), .B(n11715), .Z(n11717) );
  XOR U12232 ( .A(b[61]), .B(a[11]), .Z(n12044) );
  NANDN U12233 ( .A(n38248), .B(n12044), .Z(n11716) );
  AND U12234 ( .A(n11717), .B(n11716), .Z(n11871) );
  AND U12235 ( .A(b[63]), .B(a[7]), .Z(n11870) );
  XOR U12236 ( .A(n11871), .B(n11870), .Z(n11873) );
  XNOR U12237 ( .A(n11872), .B(n11873), .Z(n11882) );
  XNOR U12238 ( .A(n11883), .B(n11882), .Z(n11884) );
  NANDN U12239 ( .A(n11719), .B(n11718), .Z(n11723) );
  OR U12240 ( .A(n11721), .B(n11720), .Z(n11722) );
  NAND U12241 ( .A(n11723), .B(n11722), .Z(n11885) );
  XNOR U12242 ( .A(n11884), .B(n11885), .Z(n12077) );
  NANDN U12243 ( .A(n34223), .B(n11724), .Z(n11726) );
  XOR U12244 ( .A(b[27]), .B(a[45]), .Z(n12053) );
  NANDN U12245 ( .A(n34458), .B(n12053), .Z(n11725) );
  AND U12246 ( .A(n11726), .B(n11725), .Z(n11944) );
  NANDN U12247 ( .A(n34634), .B(n11727), .Z(n11729) );
  XOR U12248 ( .A(b[29]), .B(a[43]), .Z(n12056) );
  NANDN U12249 ( .A(n34722), .B(n12056), .Z(n11728) );
  AND U12250 ( .A(n11729), .B(n11728), .Z(n11943) );
  NANDN U12251 ( .A(n31055), .B(n11730), .Z(n11732) );
  XOR U12252 ( .A(b[13]), .B(a[59]), .Z(n12059) );
  NANDN U12253 ( .A(n31293), .B(n12059), .Z(n11731) );
  NAND U12254 ( .A(n11732), .B(n11731), .Z(n11942) );
  XOR U12255 ( .A(n11943), .B(n11942), .Z(n11945) );
  XOR U12256 ( .A(n11944), .B(n11945), .Z(n11973) );
  NANDN U12257 ( .A(n28889), .B(n11733), .Z(n11735) );
  XOR U12258 ( .A(b[5]), .B(a[67]), .Z(n12062) );
  NANDN U12259 ( .A(n29138), .B(n12062), .Z(n11734) );
  AND U12260 ( .A(n11735), .B(n11734), .Z(n11992) );
  NANDN U12261 ( .A(n209), .B(n11736), .Z(n11738) );
  XOR U12262 ( .A(b[3]), .B(a[69]), .Z(n12065) );
  NANDN U12263 ( .A(n28941), .B(n12065), .Z(n11737) );
  AND U12264 ( .A(n11738), .B(n11737), .Z(n11991) );
  NANDN U12265 ( .A(n35936), .B(n11739), .Z(n11741) );
  XOR U12266 ( .A(b[37]), .B(a[35]), .Z(n12068) );
  NANDN U12267 ( .A(n36047), .B(n12068), .Z(n11740) );
  NAND U12268 ( .A(n11741), .B(n11740), .Z(n11990) );
  XOR U12269 ( .A(n11991), .B(n11990), .Z(n11993) );
  XNOR U12270 ( .A(n11992), .B(n11993), .Z(n11972) );
  XNOR U12271 ( .A(n11973), .B(n11972), .Z(n11974) );
  NANDN U12272 ( .A(n11743), .B(n11742), .Z(n11747) );
  OR U12273 ( .A(n11745), .B(n11744), .Z(n11746) );
  NAND U12274 ( .A(n11747), .B(n11746), .Z(n11975) );
  XOR U12275 ( .A(n11974), .B(n11975), .Z(n12078) );
  XNOR U12276 ( .A(n12077), .B(n12078), .Z(n12079) );
  XNOR U12277 ( .A(n12080), .B(n12079), .Z(n11963) );
  NANDN U12278 ( .A(n11749), .B(n11748), .Z(n11753) );
  NANDN U12279 ( .A(n11751), .B(n11750), .Z(n11752) );
  AND U12280 ( .A(n11753), .B(n11752), .Z(n11979) );
  NANDN U12281 ( .A(n11755), .B(n11754), .Z(n11759) );
  OR U12282 ( .A(n11757), .B(n11756), .Z(n11758) );
  NAND U12283 ( .A(n11759), .B(n11758), .Z(n11978) );
  XNOR U12284 ( .A(n11979), .B(n11978), .Z(n11981) );
  NANDN U12285 ( .A(n11761), .B(n11760), .Z(n11765) );
  OR U12286 ( .A(n11763), .B(n11762), .Z(n11764) );
  AND U12287 ( .A(n11765), .B(n11764), .Z(n11921) );
  NAND U12288 ( .A(b[0]), .B(a[71]), .Z(n11766) );
  XNOR U12289 ( .A(b[1]), .B(n11766), .Z(n11768) );
  NANDN U12290 ( .A(b[0]), .B(a[70]), .Z(n11767) );
  NAND U12291 ( .A(n11768), .B(n11767), .Z(n11957) );
  NANDN U12292 ( .A(n38278), .B(n11769), .Z(n11771) );
  XOR U12293 ( .A(b[63]), .B(a[9]), .Z(n12005) );
  NANDN U12294 ( .A(n38279), .B(n12005), .Z(n11770) );
  AND U12295 ( .A(n11771), .B(n11770), .Z(n11955) );
  NANDN U12296 ( .A(n35260), .B(n11772), .Z(n11774) );
  XOR U12297 ( .A(b[33]), .B(a[39]), .Z(n12008) );
  NANDN U12298 ( .A(n35456), .B(n12008), .Z(n11773) );
  NAND U12299 ( .A(n11774), .B(n11773), .Z(n11954) );
  XNOR U12300 ( .A(n11955), .B(n11954), .Z(n11956) );
  XNOR U12301 ( .A(n11957), .B(n11956), .Z(n11918) );
  NANDN U12302 ( .A(n37974), .B(n11775), .Z(n11777) );
  XOR U12303 ( .A(b[57]), .B(a[15]), .Z(n12011) );
  NANDN U12304 ( .A(n38031), .B(n12011), .Z(n11776) );
  AND U12305 ( .A(n11777), .B(n11776), .Z(n11987) );
  NANDN U12306 ( .A(n38090), .B(n11778), .Z(n11780) );
  XOR U12307 ( .A(b[59]), .B(a[13]), .Z(n12014) );
  NANDN U12308 ( .A(n38130), .B(n12014), .Z(n11779) );
  AND U12309 ( .A(n11780), .B(n11779), .Z(n11985) );
  NANDN U12310 ( .A(n36480), .B(n11781), .Z(n11783) );
  XOR U12311 ( .A(b[41]), .B(a[31]), .Z(n12017) );
  NANDN U12312 ( .A(n36594), .B(n12017), .Z(n11782) );
  NAND U12313 ( .A(n11783), .B(n11782), .Z(n11984) );
  XNOR U12314 ( .A(n11985), .B(n11984), .Z(n11986) );
  XOR U12315 ( .A(n11987), .B(n11986), .Z(n11919) );
  XNOR U12316 ( .A(n11918), .B(n11919), .Z(n11920) );
  XNOR U12317 ( .A(n11921), .B(n11920), .Z(n11980) );
  XOR U12318 ( .A(n11981), .B(n11980), .Z(n11961) );
  NANDN U12319 ( .A(n11785), .B(n11784), .Z(n11789) );
  NAND U12320 ( .A(n11787), .B(n11786), .Z(n11788) );
  NAND U12321 ( .A(n11789), .B(n11788), .Z(n11960) );
  XNOR U12322 ( .A(n11961), .B(n11960), .Z(n11962) );
  XOR U12323 ( .A(n11963), .B(n11962), .Z(n11856) );
  NANDN U12324 ( .A(n11791), .B(n11790), .Z(n11795) );
  NANDN U12325 ( .A(n11793), .B(n11792), .Z(n11794) );
  AND U12326 ( .A(n11795), .B(n11794), .Z(n11855) );
  XNOR U12327 ( .A(n11856), .B(n11855), .Z(n11857) );
  XNOR U12328 ( .A(n11858), .B(n11857), .Z(n11819) );
  XNOR U12329 ( .A(n11820), .B(n11819), .Z(n11821) );
  XOR U12330 ( .A(n11822), .B(n11821), .Z(n12086) );
  XOR U12331 ( .A(n12085), .B(n12086), .Z(n12092) );
  XOR U12332 ( .A(n12091), .B(n12092), .Z(n11814) );
  XOR U12333 ( .A(n11813), .B(n11814), .Z(n11816) );
  XOR U12334 ( .A(n11815), .B(n11816), .Z(n11808) );
  NANDN U12335 ( .A(n11797), .B(n11796), .Z(n11801) );
  NANDN U12336 ( .A(n11799), .B(n11798), .Z(n11800) );
  NAND U12337 ( .A(n11801), .B(n11800), .Z(n11807) );
  XNOR U12338 ( .A(n11808), .B(n11807), .Z(n11809) );
  XNOR U12339 ( .A(n11810), .B(n11809), .Z(n12095) );
  XNOR U12340 ( .A(sreg[135]), .B(n12095), .Z(n12097) );
  NANDN U12341 ( .A(sreg[134]), .B(n11802), .Z(n11806) );
  NAND U12342 ( .A(n11804), .B(n11803), .Z(n11805) );
  NAND U12343 ( .A(n11806), .B(n11805), .Z(n12096) );
  XNOR U12344 ( .A(n12097), .B(n12096), .Z(c[135]) );
  NANDN U12345 ( .A(n11808), .B(n11807), .Z(n11812) );
  NANDN U12346 ( .A(n11810), .B(n11809), .Z(n11811) );
  AND U12347 ( .A(n11812), .B(n11811), .Z(n12103) );
  NANDN U12348 ( .A(n11814), .B(n11813), .Z(n11818) );
  OR U12349 ( .A(n11816), .B(n11815), .Z(n11817) );
  AND U12350 ( .A(n11818), .B(n11817), .Z(n12100) );
  NANDN U12351 ( .A(n11820), .B(n11819), .Z(n11824) );
  NANDN U12352 ( .A(n11822), .B(n11821), .Z(n11823) );
  AND U12353 ( .A(n11824), .B(n11823), .Z(n12383) );
  NANDN U12354 ( .A(n11826), .B(n11825), .Z(n11830) );
  NANDN U12355 ( .A(n11828), .B(n11827), .Z(n11829) );
  NAND U12356 ( .A(n11830), .B(n11829), .Z(n12382) );
  XNOR U12357 ( .A(n12383), .B(n12382), .Z(n12385) );
  NANDN U12358 ( .A(n11832), .B(n11831), .Z(n11836) );
  OR U12359 ( .A(n11834), .B(n11833), .Z(n11835) );
  AND U12360 ( .A(n11836), .B(n11835), .Z(n12120) );
  NANDN U12361 ( .A(n11838), .B(n11837), .Z(n11842) );
  NANDN U12362 ( .A(n11840), .B(n11839), .Z(n11841) );
  AND U12363 ( .A(n11842), .B(n11841), .Z(n12119) );
  NANDN U12364 ( .A(n11844), .B(n11843), .Z(n11848) );
  OR U12365 ( .A(n11846), .B(n11845), .Z(n11847) );
  AND U12366 ( .A(n11848), .B(n11847), .Z(n12118) );
  XOR U12367 ( .A(n12119), .B(n12118), .Z(n12121) );
  XOR U12368 ( .A(n12120), .B(n12121), .Z(n12377) );
  NANDN U12369 ( .A(n11850), .B(n11849), .Z(n11854) );
  OR U12370 ( .A(n11852), .B(n11851), .Z(n11853) );
  AND U12371 ( .A(n11854), .B(n11853), .Z(n12376) );
  XNOR U12372 ( .A(n12377), .B(n12376), .Z(n12378) );
  NANDN U12373 ( .A(n11856), .B(n11855), .Z(n11860) );
  NANDN U12374 ( .A(n11858), .B(n11857), .Z(n11859) );
  AND U12375 ( .A(n11860), .B(n11859), .Z(n12115) );
  NANDN U12376 ( .A(n29499), .B(n11861), .Z(n11863) );
  XOR U12377 ( .A(b[7]), .B(a[66]), .Z(n12238) );
  NANDN U12378 ( .A(n29735), .B(n12238), .Z(n11862) );
  AND U12379 ( .A(n11863), .B(n11862), .Z(n12198) );
  NANDN U12380 ( .A(n37857), .B(n11864), .Z(n11866) );
  XOR U12381 ( .A(b[55]), .B(a[18]), .Z(n12241) );
  NANDN U12382 ( .A(n37911), .B(n12241), .Z(n11865) );
  AND U12383 ( .A(n11866), .B(n11865), .Z(n12197) );
  NANDN U12384 ( .A(n35611), .B(n11867), .Z(n11869) );
  XOR U12385 ( .A(b[35]), .B(a[38]), .Z(n12244) );
  NANDN U12386 ( .A(n35801), .B(n12244), .Z(n11868) );
  NAND U12387 ( .A(n11869), .B(n11868), .Z(n12196) );
  XOR U12388 ( .A(n12197), .B(n12196), .Z(n12199) );
  XOR U12389 ( .A(n12198), .B(n12199), .Z(n12260) );
  NANDN U12390 ( .A(n11871), .B(n11870), .Z(n11875) );
  OR U12391 ( .A(n11873), .B(n11872), .Z(n11874) );
  AND U12392 ( .A(n11875), .B(n11874), .Z(n12259) );
  XNOR U12393 ( .A(n12260), .B(n12259), .Z(n12261) );
  NANDN U12394 ( .A(n11877), .B(n11876), .Z(n11881) );
  OR U12395 ( .A(n11879), .B(n11878), .Z(n11880) );
  NAND U12396 ( .A(n11881), .B(n11880), .Z(n12262) );
  XNOR U12397 ( .A(n12261), .B(n12262), .Z(n12139) );
  NANDN U12398 ( .A(n11883), .B(n11882), .Z(n11887) );
  NANDN U12399 ( .A(n11885), .B(n11884), .Z(n11886) );
  AND U12400 ( .A(n11887), .B(n11886), .Z(n12137) );
  NANDN U12401 ( .A(n211), .B(n11888), .Z(n11890) );
  XOR U12402 ( .A(b[47]), .B(a[26]), .Z(n12214) );
  NANDN U12403 ( .A(n37172), .B(n12214), .Z(n11889) );
  AND U12404 ( .A(n11890), .B(n11889), .Z(n12255) );
  NANDN U12405 ( .A(n210), .B(n11891), .Z(n11893) );
  XOR U12406 ( .A(b[9]), .B(a[64]), .Z(n12217) );
  NANDN U12407 ( .A(n30267), .B(n12217), .Z(n11892) );
  AND U12408 ( .A(n11893), .B(n11892), .Z(n12254) );
  NANDN U12409 ( .A(n212), .B(n11894), .Z(n11896) );
  XOR U12410 ( .A(b[49]), .B(a[24]), .Z(n12220) );
  NANDN U12411 ( .A(n37432), .B(n12220), .Z(n11895) );
  NAND U12412 ( .A(n11896), .B(n11895), .Z(n12253) );
  XOR U12413 ( .A(n12254), .B(n12253), .Z(n12256) );
  XOR U12414 ( .A(n12255), .B(n12256), .Z(n12320) );
  NANDN U12415 ( .A(n36742), .B(n11897), .Z(n11899) );
  XOR U12416 ( .A(b[43]), .B(a[30]), .Z(n12223) );
  NANDN U12417 ( .A(n36891), .B(n12223), .Z(n11898) );
  AND U12418 ( .A(n11899), .B(n11898), .Z(n12234) );
  NANDN U12419 ( .A(n36991), .B(n11900), .Z(n11902) );
  XOR U12420 ( .A(b[45]), .B(a[28]), .Z(n12226) );
  NANDN U12421 ( .A(n37083), .B(n12226), .Z(n11901) );
  AND U12422 ( .A(n11902), .B(n11901), .Z(n12233) );
  NANDN U12423 ( .A(n30482), .B(n11903), .Z(n11905) );
  XOR U12424 ( .A(b[11]), .B(a[62]), .Z(n12229) );
  NANDN U12425 ( .A(n30891), .B(n12229), .Z(n11904) );
  NAND U12426 ( .A(n11905), .B(n11904), .Z(n12232) );
  XOR U12427 ( .A(n12233), .B(n12232), .Z(n12235) );
  XNOR U12428 ( .A(n12234), .B(n12235), .Z(n12319) );
  XNOR U12429 ( .A(n12320), .B(n12319), .Z(n12321) );
  NANDN U12430 ( .A(n11907), .B(n11906), .Z(n11911) );
  OR U12431 ( .A(n11909), .B(n11908), .Z(n11910) );
  NAND U12432 ( .A(n11911), .B(n11910), .Z(n12322) );
  XNOR U12433 ( .A(n12321), .B(n12322), .Z(n12136) );
  XNOR U12434 ( .A(n12137), .B(n12136), .Z(n12138) );
  XOR U12435 ( .A(n12139), .B(n12138), .Z(n12125) );
  NANDN U12436 ( .A(n11913), .B(n11912), .Z(n11917) );
  NANDN U12437 ( .A(n11915), .B(n11914), .Z(n11916) );
  AND U12438 ( .A(n11917), .B(n11916), .Z(n12145) );
  NANDN U12439 ( .A(n11919), .B(n11918), .Z(n11923) );
  NANDN U12440 ( .A(n11921), .B(n11920), .Z(n11922) );
  AND U12441 ( .A(n11923), .B(n11922), .Z(n12143) );
  NANDN U12442 ( .A(n33875), .B(n11924), .Z(n11926) );
  XOR U12443 ( .A(b[25]), .B(a[48]), .Z(n12172) );
  NANDN U12444 ( .A(n33994), .B(n12172), .Z(n11925) );
  AND U12445 ( .A(n11926), .B(n11925), .Z(n12342) );
  NANDN U12446 ( .A(n32013), .B(n11927), .Z(n11929) );
  XOR U12447 ( .A(b[17]), .B(a[56]), .Z(n12175) );
  NANDN U12448 ( .A(n32292), .B(n12175), .Z(n11928) );
  AND U12449 ( .A(n11929), .B(n11928), .Z(n12341) );
  NANDN U12450 ( .A(n31536), .B(n11930), .Z(n11932) );
  XOR U12451 ( .A(b[15]), .B(a[58]), .Z(n12178) );
  NANDN U12452 ( .A(n31925), .B(n12178), .Z(n11931) );
  NAND U12453 ( .A(n11932), .B(n11931), .Z(n12340) );
  XOR U12454 ( .A(n12341), .B(n12340), .Z(n12343) );
  XOR U12455 ( .A(n12342), .B(n12343), .Z(n12314) );
  NANDN U12456 ( .A(n37526), .B(n11933), .Z(n11935) );
  XOR U12457 ( .A(b[51]), .B(a[22]), .Z(n12181) );
  NANDN U12458 ( .A(n37605), .B(n12181), .Z(n11934) );
  AND U12459 ( .A(n11935), .B(n11934), .Z(n12366) );
  NANDN U12460 ( .A(n37705), .B(n11936), .Z(n11938) );
  XOR U12461 ( .A(b[53]), .B(a[20]), .Z(n12184) );
  NANDN U12462 ( .A(n37778), .B(n12184), .Z(n11937) );
  AND U12463 ( .A(n11938), .B(n11937), .Z(n12365) );
  NANDN U12464 ( .A(n36210), .B(n11939), .Z(n11941) );
  XOR U12465 ( .A(b[39]), .B(a[34]), .Z(n12187) );
  NANDN U12466 ( .A(n36347), .B(n12187), .Z(n11940) );
  NAND U12467 ( .A(n11941), .B(n11940), .Z(n12364) );
  XOR U12468 ( .A(n12365), .B(n12364), .Z(n12367) );
  XNOR U12469 ( .A(n12366), .B(n12367), .Z(n12313) );
  XNOR U12470 ( .A(n12314), .B(n12313), .Z(n12316) );
  NANDN U12471 ( .A(n11943), .B(n11942), .Z(n11947) );
  OR U12472 ( .A(n11945), .B(n11944), .Z(n11946) );
  AND U12473 ( .A(n11947), .B(n11946), .Z(n12315) );
  XOR U12474 ( .A(n12316), .B(n12315), .Z(n12163) );
  NANDN U12475 ( .A(n11949), .B(n11948), .Z(n11953) );
  OR U12476 ( .A(n11951), .B(n11950), .Z(n11952) );
  AND U12477 ( .A(n11953), .B(n11952), .Z(n12161) );
  NANDN U12478 ( .A(n11955), .B(n11954), .Z(n11959) );
  NANDN U12479 ( .A(n11957), .B(n11956), .Z(n11958) );
  NAND U12480 ( .A(n11959), .B(n11958), .Z(n12160) );
  XNOR U12481 ( .A(n12161), .B(n12160), .Z(n12162) );
  XNOR U12482 ( .A(n12163), .B(n12162), .Z(n12142) );
  XNOR U12483 ( .A(n12143), .B(n12142), .Z(n12144) );
  XNOR U12484 ( .A(n12145), .B(n12144), .Z(n12124) );
  XNOR U12485 ( .A(n12125), .B(n12124), .Z(n12126) );
  NANDN U12486 ( .A(n11961), .B(n11960), .Z(n11965) );
  NAND U12487 ( .A(n11963), .B(n11962), .Z(n11964) );
  NAND U12488 ( .A(n11965), .B(n11964), .Z(n12127) );
  XNOR U12489 ( .A(n12126), .B(n12127), .Z(n12112) );
  NANDN U12490 ( .A(n11967), .B(n11966), .Z(n11971) );
  NANDN U12491 ( .A(n11969), .B(n11968), .Z(n11970) );
  AND U12492 ( .A(n11971), .B(n11970), .Z(n12132) );
  NANDN U12493 ( .A(n11973), .B(n11972), .Z(n11977) );
  NANDN U12494 ( .A(n11975), .B(n11974), .Z(n11976) );
  AND U12495 ( .A(n11977), .B(n11976), .Z(n12131) );
  NANDN U12496 ( .A(n11979), .B(n11978), .Z(n11983) );
  NAND U12497 ( .A(n11981), .B(n11980), .Z(n11982) );
  AND U12498 ( .A(n11983), .B(n11982), .Z(n12130) );
  XOR U12499 ( .A(n12131), .B(n12130), .Z(n12133) );
  XOR U12500 ( .A(n12132), .B(n12133), .Z(n12151) );
  NANDN U12501 ( .A(n11985), .B(n11984), .Z(n11989) );
  NANDN U12502 ( .A(n11987), .B(n11986), .Z(n11988) );
  AND U12503 ( .A(n11989), .B(n11988), .Z(n12272) );
  NANDN U12504 ( .A(n11991), .B(n11990), .Z(n11995) );
  OR U12505 ( .A(n11993), .B(n11992), .Z(n11994) );
  NAND U12506 ( .A(n11995), .B(n11994), .Z(n12271) );
  XNOR U12507 ( .A(n12272), .B(n12271), .Z(n12274) );
  NANDN U12508 ( .A(n11997), .B(n11996), .Z(n12001) );
  OR U12509 ( .A(n11999), .B(n11998), .Z(n12000) );
  AND U12510 ( .A(n12001), .B(n12000), .Z(n12169) );
  NAND U12511 ( .A(b[0]), .B(a[72]), .Z(n12002) );
  XNOR U12512 ( .A(b[1]), .B(n12002), .Z(n12004) );
  NANDN U12513 ( .A(b[0]), .B(a[71]), .Z(n12003) );
  NAND U12514 ( .A(n12004), .B(n12003), .Z(n12205) );
  NANDN U12515 ( .A(n38278), .B(n12005), .Z(n12007) );
  XOR U12516 ( .A(b[63]), .B(a[10]), .Z(n12295) );
  NANDN U12517 ( .A(n38279), .B(n12295), .Z(n12006) );
  AND U12518 ( .A(n12007), .B(n12006), .Z(n12203) );
  NANDN U12519 ( .A(n35260), .B(n12008), .Z(n12010) );
  XOR U12520 ( .A(b[33]), .B(a[40]), .Z(n12298) );
  NANDN U12521 ( .A(n35456), .B(n12298), .Z(n12009) );
  NAND U12522 ( .A(n12010), .B(n12009), .Z(n12202) );
  XNOR U12523 ( .A(n12203), .B(n12202), .Z(n12204) );
  XNOR U12524 ( .A(n12205), .B(n12204), .Z(n12166) );
  NANDN U12525 ( .A(n37974), .B(n12011), .Z(n12013) );
  XOR U12526 ( .A(b[57]), .B(a[16]), .Z(n12304) );
  NANDN U12527 ( .A(n38031), .B(n12304), .Z(n12012) );
  AND U12528 ( .A(n12013), .B(n12012), .Z(n12280) );
  NANDN U12529 ( .A(n38090), .B(n12014), .Z(n12016) );
  XOR U12530 ( .A(b[59]), .B(a[14]), .Z(n12307) );
  NANDN U12531 ( .A(n38130), .B(n12307), .Z(n12015) );
  AND U12532 ( .A(n12016), .B(n12015), .Z(n12278) );
  NANDN U12533 ( .A(n36480), .B(n12017), .Z(n12019) );
  XOR U12534 ( .A(b[41]), .B(a[32]), .Z(n12310) );
  NANDN U12535 ( .A(n36594), .B(n12310), .Z(n12018) );
  NAND U12536 ( .A(n12019), .B(n12018), .Z(n12277) );
  XNOR U12537 ( .A(n12278), .B(n12277), .Z(n12279) );
  XOR U12538 ( .A(n12280), .B(n12279), .Z(n12167) );
  XNOR U12539 ( .A(n12166), .B(n12167), .Z(n12168) );
  XNOR U12540 ( .A(n12169), .B(n12168), .Z(n12273) );
  XOR U12541 ( .A(n12274), .B(n12273), .Z(n12155) );
  NANDN U12542 ( .A(n12021), .B(n12020), .Z(n12025) );
  NAND U12543 ( .A(n12023), .B(n12022), .Z(n12024) );
  NAND U12544 ( .A(n12025), .B(n12024), .Z(n12154) );
  XNOR U12545 ( .A(n12155), .B(n12154), .Z(n12157) );
  NANDN U12546 ( .A(n12027), .B(n12026), .Z(n12031) );
  NANDN U12547 ( .A(n12029), .B(n12028), .Z(n12030) );
  AND U12548 ( .A(n12031), .B(n12030), .Z(n12373) );
  NANDN U12549 ( .A(n32996), .B(n12032), .Z(n12034) );
  XOR U12550 ( .A(b[21]), .B(a[52]), .Z(n12325) );
  NANDN U12551 ( .A(n33271), .B(n12325), .Z(n12033) );
  AND U12552 ( .A(n12034), .B(n12033), .Z(n12291) );
  NANDN U12553 ( .A(n33866), .B(n12035), .Z(n12037) );
  XOR U12554 ( .A(b[23]), .B(a[50]), .Z(n12328) );
  NANDN U12555 ( .A(n33644), .B(n12328), .Z(n12036) );
  AND U12556 ( .A(n12037), .B(n12036), .Z(n12290) );
  NANDN U12557 ( .A(n32483), .B(n12038), .Z(n12040) );
  XOR U12558 ( .A(b[19]), .B(a[54]), .Z(n12331) );
  NANDN U12559 ( .A(n32823), .B(n12331), .Z(n12039) );
  NAND U12560 ( .A(n12040), .B(n12039), .Z(n12289) );
  XOR U12561 ( .A(n12290), .B(n12289), .Z(n12292) );
  XOR U12562 ( .A(n12291), .B(n12292), .Z(n12209) );
  NANDN U12563 ( .A(n34909), .B(n12041), .Z(n12043) );
  XOR U12564 ( .A(b[31]), .B(a[42]), .Z(n12334) );
  NANDN U12565 ( .A(n35145), .B(n12334), .Z(n12042) );
  AND U12566 ( .A(n12043), .B(n12042), .Z(n12249) );
  NANDN U12567 ( .A(n38247), .B(n12044), .Z(n12046) );
  XOR U12568 ( .A(b[61]), .B(a[12]), .Z(n12337) );
  NANDN U12569 ( .A(n38248), .B(n12337), .Z(n12045) );
  AND U12570 ( .A(n12046), .B(n12045), .Z(n12248) );
  AND U12571 ( .A(b[63]), .B(a[8]), .Z(n12247) );
  XOR U12572 ( .A(n12248), .B(n12247), .Z(n12250) );
  XNOR U12573 ( .A(n12249), .B(n12250), .Z(n12208) );
  XNOR U12574 ( .A(n12209), .B(n12208), .Z(n12210) );
  NANDN U12575 ( .A(n12048), .B(n12047), .Z(n12052) );
  OR U12576 ( .A(n12050), .B(n12049), .Z(n12051) );
  NAND U12577 ( .A(n12052), .B(n12051), .Z(n12211) );
  XNOR U12578 ( .A(n12210), .B(n12211), .Z(n12370) );
  NANDN U12579 ( .A(n34223), .B(n12053), .Z(n12055) );
  XOR U12580 ( .A(b[27]), .B(a[46]), .Z(n12346) );
  NANDN U12581 ( .A(n34458), .B(n12346), .Z(n12054) );
  AND U12582 ( .A(n12055), .B(n12054), .Z(n12192) );
  NANDN U12583 ( .A(n34634), .B(n12056), .Z(n12058) );
  XOR U12584 ( .A(b[29]), .B(a[44]), .Z(n12349) );
  NANDN U12585 ( .A(n34722), .B(n12349), .Z(n12057) );
  AND U12586 ( .A(n12058), .B(n12057), .Z(n12191) );
  NANDN U12587 ( .A(n31055), .B(n12059), .Z(n12061) );
  XOR U12588 ( .A(b[13]), .B(a[60]), .Z(n12352) );
  NANDN U12589 ( .A(n31293), .B(n12352), .Z(n12060) );
  NAND U12590 ( .A(n12061), .B(n12060), .Z(n12190) );
  XOR U12591 ( .A(n12191), .B(n12190), .Z(n12193) );
  XOR U12592 ( .A(n12192), .B(n12193), .Z(n12266) );
  NANDN U12593 ( .A(n28889), .B(n12062), .Z(n12064) );
  XOR U12594 ( .A(b[5]), .B(a[68]), .Z(n12355) );
  NANDN U12595 ( .A(n29138), .B(n12355), .Z(n12063) );
  AND U12596 ( .A(n12064), .B(n12063), .Z(n12285) );
  NANDN U12597 ( .A(n209), .B(n12065), .Z(n12067) );
  XOR U12598 ( .A(a[70]), .B(b[3]), .Z(n12358) );
  NANDN U12599 ( .A(n28941), .B(n12358), .Z(n12066) );
  AND U12600 ( .A(n12067), .B(n12066), .Z(n12284) );
  NANDN U12601 ( .A(n35936), .B(n12068), .Z(n12070) );
  XOR U12602 ( .A(b[37]), .B(a[36]), .Z(n12361) );
  NANDN U12603 ( .A(n36047), .B(n12361), .Z(n12069) );
  NAND U12604 ( .A(n12070), .B(n12069), .Z(n12283) );
  XOR U12605 ( .A(n12284), .B(n12283), .Z(n12286) );
  XNOR U12606 ( .A(n12285), .B(n12286), .Z(n12265) );
  XNOR U12607 ( .A(n12266), .B(n12265), .Z(n12267) );
  NANDN U12608 ( .A(n12072), .B(n12071), .Z(n12076) );
  OR U12609 ( .A(n12074), .B(n12073), .Z(n12075) );
  NAND U12610 ( .A(n12076), .B(n12075), .Z(n12268) );
  XOR U12611 ( .A(n12267), .B(n12268), .Z(n12371) );
  XNOR U12612 ( .A(n12370), .B(n12371), .Z(n12372) );
  XNOR U12613 ( .A(n12373), .B(n12372), .Z(n12156) );
  XOR U12614 ( .A(n12157), .B(n12156), .Z(n12149) );
  NANDN U12615 ( .A(n12078), .B(n12077), .Z(n12082) );
  NANDN U12616 ( .A(n12080), .B(n12079), .Z(n12081) );
  AND U12617 ( .A(n12082), .B(n12081), .Z(n12148) );
  XNOR U12618 ( .A(n12149), .B(n12148), .Z(n12150) );
  XOR U12619 ( .A(n12151), .B(n12150), .Z(n12113) );
  XNOR U12620 ( .A(n12112), .B(n12113), .Z(n12114) );
  XOR U12621 ( .A(n12115), .B(n12114), .Z(n12379) );
  XNOR U12622 ( .A(n12378), .B(n12379), .Z(n12384) );
  XOR U12623 ( .A(n12385), .B(n12384), .Z(n12107) );
  NANDN U12624 ( .A(n12084), .B(n12083), .Z(n12088) );
  NANDN U12625 ( .A(n12086), .B(n12085), .Z(n12087) );
  AND U12626 ( .A(n12088), .B(n12087), .Z(n12106) );
  XNOR U12627 ( .A(n12107), .B(n12106), .Z(n12108) );
  NANDN U12628 ( .A(n12090), .B(n12089), .Z(n12094) );
  NANDN U12629 ( .A(n12092), .B(n12091), .Z(n12093) );
  NAND U12630 ( .A(n12094), .B(n12093), .Z(n12109) );
  XOR U12631 ( .A(n12108), .B(n12109), .Z(n12101) );
  XNOR U12632 ( .A(n12100), .B(n12101), .Z(n12102) );
  XNOR U12633 ( .A(n12103), .B(n12102), .Z(n12388) );
  XNOR U12634 ( .A(sreg[136]), .B(n12388), .Z(n12390) );
  NANDN U12635 ( .A(sreg[135]), .B(n12095), .Z(n12099) );
  NAND U12636 ( .A(n12097), .B(n12096), .Z(n12098) );
  NAND U12637 ( .A(n12099), .B(n12098), .Z(n12389) );
  XNOR U12638 ( .A(n12390), .B(n12389), .Z(c[136]) );
  NANDN U12639 ( .A(n12101), .B(n12100), .Z(n12105) );
  NANDN U12640 ( .A(n12103), .B(n12102), .Z(n12104) );
  AND U12641 ( .A(n12105), .B(n12104), .Z(n12396) );
  NANDN U12642 ( .A(n12107), .B(n12106), .Z(n12111) );
  NANDN U12643 ( .A(n12109), .B(n12108), .Z(n12110) );
  AND U12644 ( .A(n12111), .B(n12110), .Z(n12394) );
  NANDN U12645 ( .A(n12113), .B(n12112), .Z(n12117) );
  NANDN U12646 ( .A(n12115), .B(n12114), .Z(n12116) );
  AND U12647 ( .A(n12117), .B(n12116), .Z(n12676) );
  NANDN U12648 ( .A(n12119), .B(n12118), .Z(n12123) );
  OR U12649 ( .A(n12121), .B(n12120), .Z(n12122) );
  AND U12650 ( .A(n12123), .B(n12122), .Z(n12675) );
  XNOR U12651 ( .A(n12676), .B(n12675), .Z(n12678) );
  NANDN U12652 ( .A(n12125), .B(n12124), .Z(n12129) );
  NANDN U12653 ( .A(n12127), .B(n12126), .Z(n12128) );
  AND U12654 ( .A(n12129), .B(n12128), .Z(n12670) );
  NANDN U12655 ( .A(n12131), .B(n12130), .Z(n12135) );
  OR U12656 ( .A(n12133), .B(n12132), .Z(n12134) );
  AND U12657 ( .A(n12135), .B(n12134), .Z(n12413) );
  NANDN U12658 ( .A(n12137), .B(n12136), .Z(n12141) );
  NAND U12659 ( .A(n12139), .B(n12138), .Z(n12140) );
  AND U12660 ( .A(n12141), .B(n12140), .Z(n12412) );
  NANDN U12661 ( .A(n12143), .B(n12142), .Z(n12147) );
  NANDN U12662 ( .A(n12145), .B(n12144), .Z(n12146) );
  AND U12663 ( .A(n12147), .B(n12146), .Z(n12411) );
  XOR U12664 ( .A(n12412), .B(n12411), .Z(n12414) );
  XNOR U12665 ( .A(n12413), .B(n12414), .Z(n12669) );
  XNOR U12666 ( .A(n12670), .B(n12669), .Z(n12671) );
  NANDN U12667 ( .A(n12149), .B(n12148), .Z(n12153) );
  NANDN U12668 ( .A(n12151), .B(n12150), .Z(n12152) );
  AND U12669 ( .A(n12153), .B(n12152), .Z(n12408) );
  NANDN U12670 ( .A(n12155), .B(n12154), .Z(n12159) );
  NAND U12671 ( .A(n12157), .B(n12156), .Z(n12158) );
  AND U12672 ( .A(n12159), .B(n12158), .Z(n12437) );
  NANDN U12673 ( .A(n12161), .B(n12160), .Z(n12165) );
  NANDN U12674 ( .A(n12163), .B(n12162), .Z(n12164) );
  AND U12675 ( .A(n12165), .B(n12164), .Z(n12431) );
  NANDN U12676 ( .A(n12167), .B(n12166), .Z(n12171) );
  NANDN U12677 ( .A(n12169), .B(n12168), .Z(n12170) );
  AND U12678 ( .A(n12171), .B(n12170), .Z(n12430) );
  NANDN U12679 ( .A(n33875), .B(n12172), .Z(n12174) );
  XOR U12680 ( .A(b[25]), .B(a[49]), .Z(n12465) );
  NANDN U12681 ( .A(n33994), .B(n12465), .Z(n12173) );
  AND U12682 ( .A(n12174), .B(n12173), .Z(n12635) );
  NANDN U12683 ( .A(n32013), .B(n12175), .Z(n12177) );
  XOR U12684 ( .A(b[17]), .B(a[57]), .Z(n12468) );
  NANDN U12685 ( .A(n32292), .B(n12468), .Z(n12176) );
  AND U12686 ( .A(n12177), .B(n12176), .Z(n12634) );
  NANDN U12687 ( .A(n31536), .B(n12178), .Z(n12180) );
  XOR U12688 ( .A(b[15]), .B(a[59]), .Z(n12471) );
  NANDN U12689 ( .A(n31925), .B(n12471), .Z(n12179) );
  NAND U12690 ( .A(n12180), .B(n12179), .Z(n12633) );
  XOR U12691 ( .A(n12634), .B(n12633), .Z(n12636) );
  XOR U12692 ( .A(n12635), .B(n12636), .Z(n12607) );
  NANDN U12693 ( .A(n37526), .B(n12181), .Z(n12183) );
  XOR U12694 ( .A(b[51]), .B(a[23]), .Z(n12474) );
  NANDN U12695 ( .A(n37605), .B(n12474), .Z(n12182) );
  AND U12696 ( .A(n12183), .B(n12182), .Z(n12659) );
  NANDN U12697 ( .A(n37705), .B(n12184), .Z(n12186) );
  XOR U12698 ( .A(b[53]), .B(a[21]), .Z(n12477) );
  NANDN U12699 ( .A(n37778), .B(n12477), .Z(n12185) );
  AND U12700 ( .A(n12186), .B(n12185), .Z(n12658) );
  NANDN U12701 ( .A(n36210), .B(n12187), .Z(n12189) );
  XOR U12702 ( .A(b[39]), .B(a[35]), .Z(n12480) );
  NANDN U12703 ( .A(n36347), .B(n12480), .Z(n12188) );
  NAND U12704 ( .A(n12189), .B(n12188), .Z(n12657) );
  XOR U12705 ( .A(n12658), .B(n12657), .Z(n12660) );
  XNOR U12706 ( .A(n12659), .B(n12660), .Z(n12606) );
  XNOR U12707 ( .A(n12607), .B(n12606), .Z(n12609) );
  NANDN U12708 ( .A(n12191), .B(n12190), .Z(n12195) );
  OR U12709 ( .A(n12193), .B(n12192), .Z(n12194) );
  AND U12710 ( .A(n12195), .B(n12194), .Z(n12608) );
  XOR U12711 ( .A(n12609), .B(n12608), .Z(n12456) );
  NANDN U12712 ( .A(n12197), .B(n12196), .Z(n12201) );
  OR U12713 ( .A(n12199), .B(n12198), .Z(n12200) );
  AND U12714 ( .A(n12201), .B(n12200), .Z(n12454) );
  NANDN U12715 ( .A(n12203), .B(n12202), .Z(n12207) );
  NANDN U12716 ( .A(n12205), .B(n12204), .Z(n12206) );
  NAND U12717 ( .A(n12207), .B(n12206), .Z(n12453) );
  XNOR U12718 ( .A(n12454), .B(n12453), .Z(n12455) );
  XNOR U12719 ( .A(n12456), .B(n12455), .Z(n12429) );
  XOR U12720 ( .A(n12430), .B(n12429), .Z(n12432) );
  XOR U12721 ( .A(n12431), .B(n12432), .Z(n12436) );
  NANDN U12722 ( .A(n12209), .B(n12208), .Z(n12213) );
  NANDN U12723 ( .A(n12211), .B(n12210), .Z(n12212) );
  AND U12724 ( .A(n12213), .B(n12212), .Z(n12424) );
  NANDN U12725 ( .A(n211), .B(n12214), .Z(n12216) );
  XOR U12726 ( .A(b[47]), .B(a[27]), .Z(n12507) );
  NANDN U12727 ( .A(n37172), .B(n12507), .Z(n12215) );
  AND U12728 ( .A(n12216), .B(n12215), .Z(n12548) );
  NANDN U12729 ( .A(n210), .B(n12217), .Z(n12219) );
  XOR U12730 ( .A(b[9]), .B(a[65]), .Z(n12510) );
  NANDN U12731 ( .A(n30267), .B(n12510), .Z(n12218) );
  AND U12732 ( .A(n12219), .B(n12218), .Z(n12547) );
  NANDN U12733 ( .A(n212), .B(n12220), .Z(n12222) );
  XOR U12734 ( .A(b[49]), .B(a[25]), .Z(n12513) );
  NANDN U12735 ( .A(n37432), .B(n12513), .Z(n12221) );
  NAND U12736 ( .A(n12222), .B(n12221), .Z(n12546) );
  XOR U12737 ( .A(n12547), .B(n12546), .Z(n12549) );
  XOR U12738 ( .A(n12548), .B(n12549), .Z(n12613) );
  NANDN U12739 ( .A(n36742), .B(n12223), .Z(n12225) );
  XOR U12740 ( .A(b[43]), .B(a[31]), .Z(n12516) );
  NANDN U12741 ( .A(n36891), .B(n12516), .Z(n12224) );
  AND U12742 ( .A(n12225), .B(n12224), .Z(n12527) );
  NANDN U12743 ( .A(n36991), .B(n12226), .Z(n12228) );
  XOR U12744 ( .A(b[45]), .B(a[29]), .Z(n12519) );
  NANDN U12745 ( .A(n37083), .B(n12519), .Z(n12227) );
  AND U12746 ( .A(n12228), .B(n12227), .Z(n12526) );
  NANDN U12747 ( .A(n30482), .B(n12229), .Z(n12231) );
  XOR U12748 ( .A(b[11]), .B(a[63]), .Z(n12522) );
  NANDN U12749 ( .A(n30891), .B(n12522), .Z(n12230) );
  NAND U12750 ( .A(n12231), .B(n12230), .Z(n12525) );
  XOR U12751 ( .A(n12526), .B(n12525), .Z(n12528) );
  XNOR U12752 ( .A(n12527), .B(n12528), .Z(n12612) );
  XNOR U12753 ( .A(n12613), .B(n12612), .Z(n12614) );
  NANDN U12754 ( .A(n12233), .B(n12232), .Z(n12237) );
  OR U12755 ( .A(n12235), .B(n12234), .Z(n12236) );
  NAND U12756 ( .A(n12237), .B(n12236), .Z(n12615) );
  XNOR U12757 ( .A(n12614), .B(n12615), .Z(n12423) );
  XNOR U12758 ( .A(n12424), .B(n12423), .Z(n12425) );
  NANDN U12759 ( .A(n29499), .B(n12238), .Z(n12240) );
  XOR U12760 ( .A(b[7]), .B(a[67]), .Z(n12531) );
  NANDN U12761 ( .A(n29735), .B(n12531), .Z(n12239) );
  AND U12762 ( .A(n12240), .B(n12239), .Z(n12491) );
  NANDN U12763 ( .A(n37857), .B(n12241), .Z(n12243) );
  XOR U12764 ( .A(b[55]), .B(a[19]), .Z(n12534) );
  NANDN U12765 ( .A(n37911), .B(n12534), .Z(n12242) );
  AND U12766 ( .A(n12243), .B(n12242), .Z(n12490) );
  NANDN U12767 ( .A(n35611), .B(n12244), .Z(n12246) );
  XOR U12768 ( .A(b[35]), .B(a[39]), .Z(n12537) );
  NANDN U12769 ( .A(n35801), .B(n12537), .Z(n12245) );
  NAND U12770 ( .A(n12246), .B(n12245), .Z(n12489) );
  XOR U12771 ( .A(n12490), .B(n12489), .Z(n12492) );
  XOR U12772 ( .A(n12491), .B(n12492), .Z(n12553) );
  NANDN U12773 ( .A(n12248), .B(n12247), .Z(n12252) );
  OR U12774 ( .A(n12250), .B(n12249), .Z(n12251) );
  AND U12775 ( .A(n12252), .B(n12251), .Z(n12552) );
  XNOR U12776 ( .A(n12553), .B(n12552), .Z(n12554) );
  NANDN U12777 ( .A(n12254), .B(n12253), .Z(n12258) );
  OR U12778 ( .A(n12256), .B(n12255), .Z(n12257) );
  NAND U12779 ( .A(n12258), .B(n12257), .Z(n12555) );
  XOR U12780 ( .A(n12554), .B(n12555), .Z(n12426) );
  XNOR U12781 ( .A(n12425), .B(n12426), .Z(n12435) );
  XOR U12782 ( .A(n12436), .B(n12435), .Z(n12438) );
  XOR U12783 ( .A(n12437), .B(n12438), .Z(n12406) );
  NANDN U12784 ( .A(n12260), .B(n12259), .Z(n12264) );
  NANDN U12785 ( .A(n12262), .B(n12261), .Z(n12263) );
  AND U12786 ( .A(n12264), .B(n12263), .Z(n12419) );
  NANDN U12787 ( .A(n12266), .B(n12265), .Z(n12270) );
  NANDN U12788 ( .A(n12268), .B(n12267), .Z(n12269) );
  AND U12789 ( .A(n12270), .B(n12269), .Z(n12418) );
  NANDN U12790 ( .A(n12272), .B(n12271), .Z(n12276) );
  NAND U12791 ( .A(n12274), .B(n12273), .Z(n12275) );
  AND U12792 ( .A(n12276), .B(n12275), .Z(n12417) );
  XOR U12793 ( .A(n12418), .B(n12417), .Z(n12420) );
  XOR U12794 ( .A(n12419), .B(n12420), .Z(n12444) );
  NANDN U12795 ( .A(n12278), .B(n12277), .Z(n12282) );
  NANDN U12796 ( .A(n12280), .B(n12279), .Z(n12281) );
  AND U12797 ( .A(n12282), .B(n12281), .Z(n12565) );
  NANDN U12798 ( .A(n12284), .B(n12283), .Z(n12288) );
  OR U12799 ( .A(n12286), .B(n12285), .Z(n12287) );
  NAND U12800 ( .A(n12288), .B(n12287), .Z(n12564) );
  XNOR U12801 ( .A(n12565), .B(n12564), .Z(n12567) );
  NANDN U12802 ( .A(n12290), .B(n12289), .Z(n12294) );
  OR U12803 ( .A(n12292), .B(n12291), .Z(n12293) );
  AND U12804 ( .A(n12294), .B(n12293), .Z(n12462) );
  NANDN U12805 ( .A(n38278), .B(n12295), .Z(n12297) );
  XOR U12806 ( .A(b[63]), .B(a[11]), .Z(n12591) );
  NANDN U12807 ( .A(n38279), .B(n12591), .Z(n12296) );
  AND U12808 ( .A(n12297), .B(n12296), .Z(n12496) );
  NANDN U12809 ( .A(n35260), .B(n12298), .Z(n12300) );
  XOR U12810 ( .A(b[33]), .B(a[41]), .Z(n12594) );
  NANDN U12811 ( .A(n35456), .B(n12594), .Z(n12299) );
  NAND U12812 ( .A(n12300), .B(n12299), .Z(n12495) );
  XNOR U12813 ( .A(n12496), .B(n12495), .Z(n12497) );
  NAND U12814 ( .A(b[0]), .B(a[73]), .Z(n12301) );
  XNOR U12815 ( .A(b[1]), .B(n12301), .Z(n12303) );
  NANDN U12816 ( .A(b[0]), .B(a[72]), .Z(n12302) );
  NAND U12817 ( .A(n12303), .B(n12302), .Z(n12498) );
  XNOR U12818 ( .A(n12497), .B(n12498), .Z(n12459) );
  NANDN U12819 ( .A(n37974), .B(n12304), .Z(n12306) );
  XOR U12820 ( .A(b[57]), .B(a[17]), .Z(n12597) );
  NANDN U12821 ( .A(n38031), .B(n12597), .Z(n12305) );
  AND U12822 ( .A(n12306), .B(n12305), .Z(n12573) );
  NANDN U12823 ( .A(n38090), .B(n12307), .Z(n12309) );
  XOR U12824 ( .A(b[59]), .B(a[15]), .Z(n12600) );
  NANDN U12825 ( .A(n38130), .B(n12600), .Z(n12308) );
  AND U12826 ( .A(n12309), .B(n12308), .Z(n12571) );
  NANDN U12827 ( .A(n36480), .B(n12310), .Z(n12312) );
  XOR U12828 ( .A(b[41]), .B(a[33]), .Z(n12603) );
  NANDN U12829 ( .A(n36594), .B(n12603), .Z(n12311) );
  NAND U12830 ( .A(n12312), .B(n12311), .Z(n12570) );
  XNOR U12831 ( .A(n12571), .B(n12570), .Z(n12572) );
  XOR U12832 ( .A(n12573), .B(n12572), .Z(n12460) );
  XNOR U12833 ( .A(n12459), .B(n12460), .Z(n12461) );
  XNOR U12834 ( .A(n12462), .B(n12461), .Z(n12566) );
  XOR U12835 ( .A(n12567), .B(n12566), .Z(n12448) );
  NANDN U12836 ( .A(n12314), .B(n12313), .Z(n12318) );
  NAND U12837 ( .A(n12316), .B(n12315), .Z(n12317) );
  NAND U12838 ( .A(n12318), .B(n12317), .Z(n12447) );
  XNOR U12839 ( .A(n12448), .B(n12447), .Z(n12450) );
  NANDN U12840 ( .A(n12320), .B(n12319), .Z(n12324) );
  NANDN U12841 ( .A(n12322), .B(n12321), .Z(n12323) );
  AND U12842 ( .A(n12324), .B(n12323), .Z(n12666) );
  NANDN U12843 ( .A(n32996), .B(n12325), .Z(n12327) );
  XOR U12844 ( .A(b[21]), .B(a[53]), .Z(n12618) );
  NANDN U12845 ( .A(n33271), .B(n12618), .Z(n12326) );
  AND U12846 ( .A(n12327), .B(n12326), .Z(n12584) );
  NANDN U12847 ( .A(n33866), .B(n12328), .Z(n12330) );
  XOR U12848 ( .A(b[23]), .B(a[51]), .Z(n12621) );
  NANDN U12849 ( .A(n33644), .B(n12621), .Z(n12329) );
  AND U12850 ( .A(n12330), .B(n12329), .Z(n12583) );
  NANDN U12851 ( .A(n32483), .B(n12331), .Z(n12333) );
  XOR U12852 ( .A(b[19]), .B(a[55]), .Z(n12624) );
  NANDN U12853 ( .A(n32823), .B(n12624), .Z(n12332) );
  NAND U12854 ( .A(n12333), .B(n12332), .Z(n12582) );
  XOR U12855 ( .A(n12583), .B(n12582), .Z(n12585) );
  XOR U12856 ( .A(n12584), .B(n12585), .Z(n12502) );
  NANDN U12857 ( .A(n34909), .B(n12334), .Z(n12336) );
  XOR U12858 ( .A(b[31]), .B(a[43]), .Z(n12627) );
  NANDN U12859 ( .A(n35145), .B(n12627), .Z(n12335) );
  AND U12860 ( .A(n12336), .B(n12335), .Z(n12542) );
  NANDN U12861 ( .A(n38247), .B(n12337), .Z(n12339) );
  XOR U12862 ( .A(b[61]), .B(a[13]), .Z(n12630) );
  NANDN U12863 ( .A(n38248), .B(n12630), .Z(n12338) );
  AND U12864 ( .A(n12339), .B(n12338), .Z(n12541) );
  AND U12865 ( .A(b[63]), .B(a[9]), .Z(n12540) );
  XOR U12866 ( .A(n12541), .B(n12540), .Z(n12543) );
  XNOR U12867 ( .A(n12542), .B(n12543), .Z(n12501) );
  XNOR U12868 ( .A(n12502), .B(n12501), .Z(n12503) );
  NANDN U12869 ( .A(n12341), .B(n12340), .Z(n12345) );
  OR U12870 ( .A(n12343), .B(n12342), .Z(n12344) );
  NAND U12871 ( .A(n12345), .B(n12344), .Z(n12504) );
  XNOR U12872 ( .A(n12503), .B(n12504), .Z(n12663) );
  NANDN U12873 ( .A(n34223), .B(n12346), .Z(n12348) );
  XOR U12874 ( .A(b[27]), .B(a[47]), .Z(n12639) );
  NANDN U12875 ( .A(n34458), .B(n12639), .Z(n12347) );
  AND U12876 ( .A(n12348), .B(n12347), .Z(n12485) );
  NANDN U12877 ( .A(n34634), .B(n12349), .Z(n12351) );
  XOR U12878 ( .A(b[29]), .B(a[45]), .Z(n12642) );
  NANDN U12879 ( .A(n34722), .B(n12642), .Z(n12350) );
  AND U12880 ( .A(n12351), .B(n12350), .Z(n12484) );
  NANDN U12881 ( .A(n31055), .B(n12352), .Z(n12354) );
  XOR U12882 ( .A(b[13]), .B(a[61]), .Z(n12645) );
  NANDN U12883 ( .A(n31293), .B(n12645), .Z(n12353) );
  NAND U12884 ( .A(n12354), .B(n12353), .Z(n12483) );
  XOR U12885 ( .A(n12484), .B(n12483), .Z(n12486) );
  XOR U12886 ( .A(n12485), .B(n12486), .Z(n12559) );
  NANDN U12887 ( .A(n28889), .B(n12355), .Z(n12357) );
  XOR U12888 ( .A(b[5]), .B(a[69]), .Z(n12648) );
  NANDN U12889 ( .A(n29138), .B(n12648), .Z(n12356) );
  AND U12890 ( .A(n12357), .B(n12356), .Z(n12578) );
  NANDN U12891 ( .A(n209), .B(n12358), .Z(n12360) );
  XOR U12892 ( .A(a[71]), .B(b[3]), .Z(n12651) );
  NANDN U12893 ( .A(n28941), .B(n12651), .Z(n12359) );
  AND U12894 ( .A(n12360), .B(n12359), .Z(n12577) );
  NANDN U12895 ( .A(n35936), .B(n12361), .Z(n12363) );
  XOR U12896 ( .A(b[37]), .B(a[37]), .Z(n12654) );
  NANDN U12897 ( .A(n36047), .B(n12654), .Z(n12362) );
  NAND U12898 ( .A(n12363), .B(n12362), .Z(n12576) );
  XOR U12899 ( .A(n12577), .B(n12576), .Z(n12579) );
  XNOR U12900 ( .A(n12578), .B(n12579), .Z(n12558) );
  XNOR U12901 ( .A(n12559), .B(n12558), .Z(n12560) );
  NANDN U12902 ( .A(n12365), .B(n12364), .Z(n12369) );
  OR U12903 ( .A(n12367), .B(n12366), .Z(n12368) );
  NAND U12904 ( .A(n12369), .B(n12368), .Z(n12561) );
  XOR U12905 ( .A(n12560), .B(n12561), .Z(n12664) );
  XNOR U12906 ( .A(n12663), .B(n12664), .Z(n12665) );
  XNOR U12907 ( .A(n12666), .B(n12665), .Z(n12449) );
  XOR U12908 ( .A(n12450), .B(n12449), .Z(n12442) );
  NANDN U12909 ( .A(n12371), .B(n12370), .Z(n12375) );
  NANDN U12910 ( .A(n12373), .B(n12372), .Z(n12374) );
  AND U12911 ( .A(n12375), .B(n12374), .Z(n12441) );
  XNOR U12912 ( .A(n12442), .B(n12441), .Z(n12443) );
  XNOR U12913 ( .A(n12444), .B(n12443), .Z(n12405) );
  XNOR U12914 ( .A(n12406), .B(n12405), .Z(n12407) );
  XOR U12915 ( .A(n12408), .B(n12407), .Z(n12672) );
  XNOR U12916 ( .A(n12671), .B(n12672), .Z(n12677) );
  XOR U12917 ( .A(n12678), .B(n12677), .Z(n12400) );
  NANDN U12918 ( .A(n12377), .B(n12376), .Z(n12381) );
  NANDN U12919 ( .A(n12379), .B(n12378), .Z(n12380) );
  AND U12920 ( .A(n12381), .B(n12380), .Z(n12399) );
  XNOR U12921 ( .A(n12400), .B(n12399), .Z(n12401) );
  NANDN U12922 ( .A(n12383), .B(n12382), .Z(n12387) );
  NAND U12923 ( .A(n12385), .B(n12384), .Z(n12386) );
  NAND U12924 ( .A(n12387), .B(n12386), .Z(n12402) );
  XNOR U12925 ( .A(n12401), .B(n12402), .Z(n12393) );
  XNOR U12926 ( .A(n12394), .B(n12393), .Z(n12395) );
  XNOR U12927 ( .A(n12396), .B(n12395), .Z(n12681) );
  XNOR U12928 ( .A(sreg[137]), .B(n12681), .Z(n12683) );
  NANDN U12929 ( .A(sreg[136]), .B(n12388), .Z(n12392) );
  NAND U12930 ( .A(n12390), .B(n12389), .Z(n12391) );
  NAND U12931 ( .A(n12392), .B(n12391), .Z(n12682) );
  XNOR U12932 ( .A(n12683), .B(n12682), .Z(c[137]) );
  NANDN U12933 ( .A(n12394), .B(n12393), .Z(n12398) );
  NANDN U12934 ( .A(n12396), .B(n12395), .Z(n12397) );
  AND U12935 ( .A(n12398), .B(n12397), .Z(n12689) );
  NANDN U12936 ( .A(n12400), .B(n12399), .Z(n12404) );
  NANDN U12937 ( .A(n12402), .B(n12401), .Z(n12403) );
  AND U12938 ( .A(n12404), .B(n12403), .Z(n12687) );
  NANDN U12939 ( .A(n12406), .B(n12405), .Z(n12410) );
  NANDN U12940 ( .A(n12408), .B(n12407), .Z(n12409) );
  AND U12941 ( .A(n12410), .B(n12409), .Z(n12969) );
  NANDN U12942 ( .A(n12412), .B(n12411), .Z(n12416) );
  OR U12943 ( .A(n12414), .B(n12413), .Z(n12415) );
  AND U12944 ( .A(n12416), .B(n12415), .Z(n12968) );
  XNOR U12945 ( .A(n12969), .B(n12968), .Z(n12971) );
  NANDN U12946 ( .A(n12418), .B(n12417), .Z(n12422) );
  OR U12947 ( .A(n12420), .B(n12419), .Z(n12421) );
  AND U12948 ( .A(n12422), .B(n12421), .Z(n12958) );
  NANDN U12949 ( .A(n12424), .B(n12423), .Z(n12428) );
  NANDN U12950 ( .A(n12426), .B(n12425), .Z(n12427) );
  AND U12951 ( .A(n12428), .B(n12427), .Z(n12957) );
  NANDN U12952 ( .A(n12430), .B(n12429), .Z(n12434) );
  OR U12953 ( .A(n12432), .B(n12431), .Z(n12433) );
  AND U12954 ( .A(n12434), .B(n12433), .Z(n12956) );
  XOR U12955 ( .A(n12957), .B(n12956), .Z(n12959) );
  XOR U12956 ( .A(n12958), .B(n12959), .Z(n12963) );
  NANDN U12957 ( .A(n12436), .B(n12435), .Z(n12440) );
  OR U12958 ( .A(n12438), .B(n12437), .Z(n12439) );
  AND U12959 ( .A(n12440), .B(n12439), .Z(n12962) );
  XNOR U12960 ( .A(n12963), .B(n12962), .Z(n12964) );
  NANDN U12961 ( .A(n12442), .B(n12441), .Z(n12446) );
  NANDN U12962 ( .A(n12444), .B(n12443), .Z(n12445) );
  AND U12963 ( .A(n12446), .B(n12445), .Z(n12953) );
  NANDN U12964 ( .A(n12448), .B(n12447), .Z(n12452) );
  NAND U12965 ( .A(n12450), .B(n12449), .Z(n12451) );
  AND U12966 ( .A(n12452), .B(n12451), .Z(n12718) );
  NANDN U12967 ( .A(n12454), .B(n12453), .Z(n12458) );
  NANDN U12968 ( .A(n12456), .B(n12455), .Z(n12457) );
  AND U12969 ( .A(n12458), .B(n12457), .Z(n12712) );
  NANDN U12970 ( .A(n12460), .B(n12459), .Z(n12464) );
  NANDN U12971 ( .A(n12462), .B(n12461), .Z(n12463) );
  AND U12972 ( .A(n12464), .B(n12463), .Z(n12711) );
  NANDN U12973 ( .A(n33875), .B(n12465), .Z(n12467) );
  XOR U12974 ( .A(b[25]), .B(a[50]), .Z(n12797) );
  NANDN U12975 ( .A(n33994), .B(n12797), .Z(n12466) );
  AND U12976 ( .A(n12467), .B(n12466), .Z(n12901) );
  NANDN U12977 ( .A(n32013), .B(n12468), .Z(n12470) );
  XOR U12978 ( .A(b[17]), .B(a[58]), .Z(n12800) );
  NANDN U12979 ( .A(n32292), .B(n12800), .Z(n12469) );
  AND U12980 ( .A(n12470), .B(n12469), .Z(n12900) );
  NANDN U12981 ( .A(n31536), .B(n12471), .Z(n12473) );
  XOR U12982 ( .A(b[15]), .B(a[60]), .Z(n12803) );
  NANDN U12983 ( .A(n31925), .B(n12803), .Z(n12472) );
  NAND U12984 ( .A(n12473), .B(n12472), .Z(n12899) );
  XOR U12985 ( .A(n12900), .B(n12899), .Z(n12902) );
  XOR U12986 ( .A(n12901), .B(n12902), .Z(n12888) );
  NANDN U12987 ( .A(n37526), .B(n12474), .Z(n12476) );
  XOR U12988 ( .A(b[51]), .B(a[24]), .Z(n12806) );
  NANDN U12989 ( .A(n37605), .B(n12806), .Z(n12475) );
  AND U12990 ( .A(n12476), .B(n12475), .Z(n12922) );
  NANDN U12991 ( .A(n37705), .B(n12477), .Z(n12479) );
  XOR U12992 ( .A(b[53]), .B(a[22]), .Z(n12809) );
  NANDN U12993 ( .A(n37778), .B(n12809), .Z(n12478) );
  AND U12994 ( .A(n12479), .B(n12478), .Z(n12921) );
  NANDN U12995 ( .A(n36210), .B(n12480), .Z(n12482) );
  XOR U12996 ( .A(b[39]), .B(a[36]), .Z(n12812) );
  NANDN U12997 ( .A(n36347), .B(n12812), .Z(n12481) );
  NAND U12998 ( .A(n12482), .B(n12481), .Z(n12920) );
  XOR U12999 ( .A(n12921), .B(n12920), .Z(n12923) );
  XNOR U13000 ( .A(n12922), .B(n12923), .Z(n12887) );
  XNOR U13001 ( .A(n12888), .B(n12887), .Z(n12890) );
  NANDN U13002 ( .A(n12484), .B(n12483), .Z(n12488) );
  OR U13003 ( .A(n12486), .B(n12485), .Z(n12487) );
  AND U13004 ( .A(n12488), .B(n12487), .Z(n12889) );
  XOR U13005 ( .A(n12890), .B(n12889), .Z(n12788) );
  NANDN U13006 ( .A(n12490), .B(n12489), .Z(n12494) );
  OR U13007 ( .A(n12492), .B(n12491), .Z(n12493) );
  AND U13008 ( .A(n12494), .B(n12493), .Z(n12786) );
  NANDN U13009 ( .A(n12496), .B(n12495), .Z(n12500) );
  NANDN U13010 ( .A(n12498), .B(n12497), .Z(n12499) );
  NAND U13011 ( .A(n12500), .B(n12499), .Z(n12785) );
  XNOR U13012 ( .A(n12786), .B(n12785), .Z(n12787) );
  XNOR U13013 ( .A(n12788), .B(n12787), .Z(n12710) );
  XOR U13014 ( .A(n12711), .B(n12710), .Z(n12713) );
  XOR U13015 ( .A(n12712), .B(n12713), .Z(n12717) );
  NANDN U13016 ( .A(n12502), .B(n12501), .Z(n12506) );
  NANDN U13017 ( .A(n12504), .B(n12503), .Z(n12505) );
  AND U13018 ( .A(n12506), .B(n12505), .Z(n12705) );
  NAND U13019 ( .A(n37294), .B(n12507), .Z(n12509) );
  XNOR U13020 ( .A(b[47]), .B(a[28]), .Z(n12740) );
  NANDN U13021 ( .A(n12740), .B(n37341), .Z(n12508) );
  NAND U13022 ( .A(n12509), .B(n12508), .Z(n12781) );
  NAND U13023 ( .A(n30627), .B(n12510), .Z(n12512) );
  XNOR U13024 ( .A(b[9]), .B(a[66]), .Z(n12743) );
  NANDN U13025 ( .A(n12743), .B(n30628), .Z(n12511) );
  NAND U13026 ( .A(n12512), .B(n12511), .Z(n12780) );
  NAND U13027 ( .A(n37536), .B(n12513), .Z(n12515) );
  XNOR U13028 ( .A(b[49]), .B(a[26]), .Z(n12746) );
  NANDN U13029 ( .A(n12746), .B(n37537), .Z(n12514) );
  NAND U13030 ( .A(n12515), .B(n12514), .Z(n12779) );
  XNOR U13031 ( .A(n12780), .B(n12779), .Z(n12782) );
  NANDN U13032 ( .A(n36742), .B(n12516), .Z(n12518) );
  XOR U13033 ( .A(b[43]), .B(a[32]), .Z(n12749) );
  NANDN U13034 ( .A(n36891), .B(n12749), .Z(n12517) );
  AND U13035 ( .A(n12518), .B(n12517), .Z(n12760) );
  NANDN U13036 ( .A(n36991), .B(n12519), .Z(n12521) );
  XOR U13037 ( .A(b[45]), .B(a[30]), .Z(n12752) );
  NANDN U13038 ( .A(n37083), .B(n12752), .Z(n12520) );
  AND U13039 ( .A(n12521), .B(n12520), .Z(n12759) );
  NANDN U13040 ( .A(n30482), .B(n12522), .Z(n12524) );
  XOR U13041 ( .A(b[11]), .B(a[64]), .Z(n12755) );
  NANDN U13042 ( .A(n30891), .B(n12755), .Z(n12523) );
  NAND U13043 ( .A(n12524), .B(n12523), .Z(n12758) );
  XOR U13044 ( .A(n12759), .B(n12758), .Z(n12761) );
  XNOR U13045 ( .A(n12760), .B(n12761), .Z(n12893) );
  XOR U13046 ( .A(n12894), .B(n12893), .Z(n12895) );
  NANDN U13047 ( .A(n12526), .B(n12525), .Z(n12530) );
  OR U13048 ( .A(n12528), .B(n12527), .Z(n12529) );
  NAND U13049 ( .A(n12530), .B(n12529), .Z(n12896) );
  XNOR U13050 ( .A(n12895), .B(n12896), .Z(n12704) );
  XNOR U13051 ( .A(n12705), .B(n12704), .Z(n12706) );
  NANDN U13052 ( .A(n29499), .B(n12531), .Z(n12533) );
  XOR U13053 ( .A(b[7]), .B(a[68]), .Z(n12764) );
  NANDN U13054 ( .A(n29735), .B(n12764), .Z(n12532) );
  AND U13055 ( .A(n12533), .B(n12532), .Z(n12823) );
  NANDN U13056 ( .A(n37857), .B(n12534), .Z(n12536) );
  XOR U13057 ( .A(b[55]), .B(a[20]), .Z(n12767) );
  NANDN U13058 ( .A(n37911), .B(n12767), .Z(n12535) );
  AND U13059 ( .A(n12536), .B(n12535), .Z(n12822) );
  NANDN U13060 ( .A(n35611), .B(n12537), .Z(n12539) );
  XOR U13061 ( .A(b[35]), .B(a[40]), .Z(n12770) );
  NANDN U13062 ( .A(n35801), .B(n12770), .Z(n12538) );
  NAND U13063 ( .A(n12539), .B(n12538), .Z(n12821) );
  XOR U13064 ( .A(n12822), .B(n12821), .Z(n12824) );
  XOR U13065 ( .A(n12823), .B(n12824), .Z(n12834) );
  NANDN U13066 ( .A(n12541), .B(n12540), .Z(n12545) );
  OR U13067 ( .A(n12543), .B(n12542), .Z(n12544) );
  AND U13068 ( .A(n12545), .B(n12544), .Z(n12833) );
  XNOR U13069 ( .A(n12834), .B(n12833), .Z(n12835) );
  NANDN U13070 ( .A(n12547), .B(n12546), .Z(n12551) );
  OR U13071 ( .A(n12549), .B(n12548), .Z(n12550) );
  NAND U13072 ( .A(n12551), .B(n12550), .Z(n12836) );
  XOR U13073 ( .A(n12835), .B(n12836), .Z(n12707) );
  XNOR U13074 ( .A(n12706), .B(n12707), .Z(n12716) );
  XOR U13075 ( .A(n12717), .B(n12716), .Z(n12719) );
  XOR U13076 ( .A(n12718), .B(n12719), .Z(n12951) );
  NANDN U13077 ( .A(n12553), .B(n12552), .Z(n12557) );
  NANDN U13078 ( .A(n12555), .B(n12554), .Z(n12556) );
  AND U13079 ( .A(n12557), .B(n12556), .Z(n12700) );
  NANDN U13080 ( .A(n12559), .B(n12558), .Z(n12563) );
  NANDN U13081 ( .A(n12561), .B(n12560), .Z(n12562) );
  AND U13082 ( .A(n12563), .B(n12562), .Z(n12699) );
  NANDN U13083 ( .A(n12565), .B(n12564), .Z(n12569) );
  NAND U13084 ( .A(n12567), .B(n12566), .Z(n12568) );
  AND U13085 ( .A(n12569), .B(n12568), .Z(n12698) );
  XOR U13086 ( .A(n12699), .B(n12698), .Z(n12701) );
  XOR U13087 ( .A(n12700), .B(n12701), .Z(n12725) );
  NANDN U13088 ( .A(n12571), .B(n12570), .Z(n12575) );
  NANDN U13089 ( .A(n12573), .B(n12572), .Z(n12574) );
  AND U13090 ( .A(n12575), .B(n12574), .Z(n12846) );
  NANDN U13091 ( .A(n12577), .B(n12576), .Z(n12581) );
  OR U13092 ( .A(n12579), .B(n12578), .Z(n12580) );
  NAND U13093 ( .A(n12581), .B(n12580), .Z(n12845) );
  XNOR U13094 ( .A(n12846), .B(n12845), .Z(n12848) );
  NANDN U13095 ( .A(n12583), .B(n12582), .Z(n12587) );
  OR U13096 ( .A(n12585), .B(n12584), .Z(n12586) );
  AND U13097 ( .A(n12587), .B(n12586), .Z(n12794) );
  NAND U13098 ( .A(b[0]), .B(a[74]), .Z(n12588) );
  XNOR U13099 ( .A(b[1]), .B(n12588), .Z(n12590) );
  NANDN U13100 ( .A(b[0]), .B(a[73]), .Z(n12589) );
  NAND U13101 ( .A(n12590), .B(n12589), .Z(n12830) );
  NANDN U13102 ( .A(n38278), .B(n12591), .Z(n12593) );
  XOR U13103 ( .A(b[63]), .B(a[12]), .Z(n12872) );
  NANDN U13104 ( .A(n38279), .B(n12872), .Z(n12592) );
  AND U13105 ( .A(n12593), .B(n12592), .Z(n12828) );
  NANDN U13106 ( .A(n35260), .B(n12594), .Z(n12596) );
  XOR U13107 ( .A(b[33]), .B(a[42]), .Z(n12875) );
  NANDN U13108 ( .A(n35456), .B(n12875), .Z(n12595) );
  NAND U13109 ( .A(n12596), .B(n12595), .Z(n12827) );
  XNOR U13110 ( .A(n12828), .B(n12827), .Z(n12829) );
  XNOR U13111 ( .A(n12830), .B(n12829), .Z(n12791) );
  NANDN U13112 ( .A(n37974), .B(n12597), .Z(n12599) );
  XOR U13113 ( .A(b[57]), .B(a[18]), .Z(n12878) );
  NANDN U13114 ( .A(n38031), .B(n12878), .Z(n12598) );
  AND U13115 ( .A(n12599), .B(n12598), .Z(n12854) );
  NANDN U13116 ( .A(n38090), .B(n12600), .Z(n12602) );
  XOR U13117 ( .A(b[59]), .B(a[16]), .Z(n12881) );
  NANDN U13118 ( .A(n38130), .B(n12881), .Z(n12601) );
  AND U13119 ( .A(n12602), .B(n12601), .Z(n12852) );
  NANDN U13120 ( .A(n36480), .B(n12603), .Z(n12605) );
  XOR U13121 ( .A(b[41]), .B(a[34]), .Z(n12884) );
  NANDN U13122 ( .A(n36594), .B(n12884), .Z(n12604) );
  NAND U13123 ( .A(n12605), .B(n12604), .Z(n12851) );
  XNOR U13124 ( .A(n12852), .B(n12851), .Z(n12853) );
  XOR U13125 ( .A(n12854), .B(n12853), .Z(n12792) );
  XNOR U13126 ( .A(n12791), .B(n12792), .Z(n12793) );
  XNOR U13127 ( .A(n12794), .B(n12793), .Z(n12847) );
  XOR U13128 ( .A(n12848), .B(n12847), .Z(n12729) );
  NANDN U13129 ( .A(n12607), .B(n12606), .Z(n12611) );
  NAND U13130 ( .A(n12609), .B(n12608), .Z(n12610) );
  NAND U13131 ( .A(n12611), .B(n12610), .Z(n12728) );
  XNOR U13132 ( .A(n12729), .B(n12728), .Z(n12731) );
  NANDN U13133 ( .A(n12613), .B(n12612), .Z(n12617) );
  NANDN U13134 ( .A(n12615), .B(n12614), .Z(n12616) );
  AND U13135 ( .A(n12617), .B(n12616), .Z(n12947) );
  NANDN U13136 ( .A(n32996), .B(n12618), .Z(n12620) );
  XOR U13137 ( .A(b[21]), .B(a[54]), .Z(n12905) );
  NANDN U13138 ( .A(n33271), .B(n12905), .Z(n12619) );
  AND U13139 ( .A(n12620), .B(n12619), .Z(n12865) );
  NANDN U13140 ( .A(n33866), .B(n12621), .Z(n12623) );
  XOR U13141 ( .A(b[23]), .B(a[52]), .Z(n12908) );
  NANDN U13142 ( .A(n33644), .B(n12908), .Z(n12622) );
  AND U13143 ( .A(n12623), .B(n12622), .Z(n12864) );
  NANDN U13144 ( .A(n32483), .B(n12624), .Z(n12626) );
  XOR U13145 ( .A(b[19]), .B(a[56]), .Z(n12911) );
  NANDN U13146 ( .A(n32823), .B(n12911), .Z(n12625) );
  NAND U13147 ( .A(n12626), .B(n12625), .Z(n12863) );
  XOR U13148 ( .A(n12864), .B(n12863), .Z(n12866) );
  XOR U13149 ( .A(n12865), .B(n12866), .Z(n12735) );
  NANDN U13150 ( .A(n34909), .B(n12627), .Z(n12629) );
  XOR U13151 ( .A(b[31]), .B(a[44]), .Z(n12914) );
  NANDN U13152 ( .A(n35145), .B(n12914), .Z(n12628) );
  AND U13153 ( .A(n12629), .B(n12628), .Z(n12775) );
  NANDN U13154 ( .A(n38247), .B(n12630), .Z(n12632) );
  XOR U13155 ( .A(b[61]), .B(a[14]), .Z(n12917) );
  NANDN U13156 ( .A(n38248), .B(n12917), .Z(n12631) );
  AND U13157 ( .A(n12632), .B(n12631), .Z(n12774) );
  AND U13158 ( .A(b[63]), .B(a[10]), .Z(n12773) );
  XOR U13159 ( .A(n12774), .B(n12773), .Z(n12776) );
  XNOR U13160 ( .A(n12775), .B(n12776), .Z(n12734) );
  XNOR U13161 ( .A(n12735), .B(n12734), .Z(n12736) );
  NANDN U13162 ( .A(n12634), .B(n12633), .Z(n12638) );
  OR U13163 ( .A(n12636), .B(n12635), .Z(n12637) );
  NAND U13164 ( .A(n12638), .B(n12637), .Z(n12737) );
  XNOR U13165 ( .A(n12736), .B(n12737), .Z(n12944) );
  NANDN U13166 ( .A(n34223), .B(n12639), .Z(n12641) );
  XOR U13167 ( .A(b[27]), .B(a[48]), .Z(n12926) );
  NANDN U13168 ( .A(n34458), .B(n12926), .Z(n12640) );
  AND U13169 ( .A(n12641), .B(n12640), .Z(n12817) );
  NANDN U13170 ( .A(n34634), .B(n12642), .Z(n12644) );
  XOR U13171 ( .A(b[29]), .B(a[46]), .Z(n12929) );
  NANDN U13172 ( .A(n34722), .B(n12929), .Z(n12643) );
  AND U13173 ( .A(n12644), .B(n12643), .Z(n12816) );
  NANDN U13174 ( .A(n31055), .B(n12645), .Z(n12647) );
  XOR U13175 ( .A(b[13]), .B(a[62]), .Z(n12932) );
  NANDN U13176 ( .A(n31293), .B(n12932), .Z(n12646) );
  NAND U13177 ( .A(n12647), .B(n12646), .Z(n12815) );
  XOR U13178 ( .A(n12816), .B(n12815), .Z(n12818) );
  XOR U13179 ( .A(n12817), .B(n12818), .Z(n12840) );
  NANDN U13180 ( .A(n28889), .B(n12648), .Z(n12650) );
  XOR U13181 ( .A(a[70]), .B(b[5]), .Z(n12935) );
  NANDN U13182 ( .A(n29138), .B(n12935), .Z(n12649) );
  AND U13183 ( .A(n12650), .B(n12649), .Z(n12859) );
  NANDN U13184 ( .A(n209), .B(n12651), .Z(n12653) );
  XOR U13185 ( .A(a[72]), .B(b[3]), .Z(n12938) );
  NANDN U13186 ( .A(n28941), .B(n12938), .Z(n12652) );
  AND U13187 ( .A(n12653), .B(n12652), .Z(n12858) );
  NANDN U13188 ( .A(n35936), .B(n12654), .Z(n12656) );
  XOR U13189 ( .A(b[37]), .B(a[38]), .Z(n12941) );
  NANDN U13190 ( .A(n36047), .B(n12941), .Z(n12655) );
  NAND U13191 ( .A(n12656), .B(n12655), .Z(n12857) );
  XOR U13192 ( .A(n12858), .B(n12857), .Z(n12860) );
  XNOR U13193 ( .A(n12859), .B(n12860), .Z(n12839) );
  XNOR U13194 ( .A(n12840), .B(n12839), .Z(n12841) );
  NANDN U13195 ( .A(n12658), .B(n12657), .Z(n12662) );
  OR U13196 ( .A(n12660), .B(n12659), .Z(n12661) );
  NAND U13197 ( .A(n12662), .B(n12661), .Z(n12842) );
  XOR U13198 ( .A(n12841), .B(n12842), .Z(n12945) );
  XNOR U13199 ( .A(n12944), .B(n12945), .Z(n12946) );
  XNOR U13200 ( .A(n12947), .B(n12946), .Z(n12730) );
  XOR U13201 ( .A(n12731), .B(n12730), .Z(n12723) );
  NANDN U13202 ( .A(n12664), .B(n12663), .Z(n12668) );
  NANDN U13203 ( .A(n12666), .B(n12665), .Z(n12667) );
  AND U13204 ( .A(n12668), .B(n12667), .Z(n12722) );
  XNOR U13205 ( .A(n12723), .B(n12722), .Z(n12724) );
  XNOR U13206 ( .A(n12725), .B(n12724), .Z(n12950) );
  XNOR U13207 ( .A(n12951), .B(n12950), .Z(n12952) );
  XOR U13208 ( .A(n12953), .B(n12952), .Z(n12965) );
  XNOR U13209 ( .A(n12964), .B(n12965), .Z(n12970) );
  XOR U13210 ( .A(n12971), .B(n12970), .Z(n12693) );
  NANDN U13211 ( .A(n12670), .B(n12669), .Z(n12674) );
  NANDN U13212 ( .A(n12672), .B(n12671), .Z(n12673) );
  AND U13213 ( .A(n12674), .B(n12673), .Z(n12692) );
  XNOR U13214 ( .A(n12693), .B(n12692), .Z(n12694) );
  NANDN U13215 ( .A(n12676), .B(n12675), .Z(n12680) );
  NAND U13216 ( .A(n12678), .B(n12677), .Z(n12679) );
  NAND U13217 ( .A(n12680), .B(n12679), .Z(n12695) );
  XNOR U13218 ( .A(n12694), .B(n12695), .Z(n12686) );
  XNOR U13219 ( .A(n12687), .B(n12686), .Z(n12688) );
  XNOR U13220 ( .A(n12689), .B(n12688), .Z(n12974) );
  XNOR U13221 ( .A(sreg[138]), .B(n12974), .Z(n12976) );
  NANDN U13222 ( .A(sreg[137]), .B(n12681), .Z(n12685) );
  NAND U13223 ( .A(n12683), .B(n12682), .Z(n12684) );
  NAND U13224 ( .A(n12685), .B(n12684), .Z(n12975) );
  XNOR U13225 ( .A(n12976), .B(n12975), .Z(c[138]) );
  NANDN U13226 ( .A(n12687), .B(n12686), .Z(n12691) );
  NANDN U13227 ( .A(n12689), .B(n12688), .Z(n12690) );
  AND U13228 ( .A(n12691), .B(n12690), .Z(n12982) );
  NANDN U13229 ( .A(n12693), .B(n12692), .Z(n12697) );
  NANDN U13230 ( .A(n12695), .B(n12694), .Z(n12696) );
  AND U13231 ( .A(n12697), .B(n12696), .Z(n12980) );
  NANDN U13232 ( .A(n12699), .B(n12698), .Z(n12703) );
  OR U13233 ( .A(n12701), .B(n12700), .Z(n12702) );
  AND U13234 ( .A(n12703), .B(n12702), .Z(n12999) );
  NANDN U13235 ( .A(n12705), .B(n12704), .Z(n12709) );
  NANDN U13236 ( .A(n12707), .B(n12706), .Z(n12708) );
  AND U13237 ( .A(n12709), .B(n12708), .Z(n12998) );
  NANDN U13238 ( .A(n12711), .B(n12710), .Z(n12715) );
  OR U13239 ( .A(n12713), .B(n12712), .Z(n12714) );
  AND U13240 ( .A(n12715), .B(n12714), .Z(n12997) );
  XOR U13241 ( .A(n12998), .B(n12997), .Z(n13000) );
  XOR U13242 ( .A(n12999), .B(n13000), .Z(n13254) );
  NANDN U13243 ( .A(n12717), .B(n12716), .Z(n12721) );
  OR U13244 ( .A(n12719), .B(n12718), .Z(n12720) );
  AND U13245 ( .A(n12721), .B(n12720), .Z(n13253) );
  XNOR U13246 ( .A(n13254), .B(n13253), .Z(n13255) );
  NANDN U13247 ( .A(n12723), .B(n12722), .Z(n12727) );
  NANDN U13248 ( .A(n12725), .B(n12724), .Z(n12726) );
  AND U13249 ( .A(n12727), .B(n12726), .Z(n12994) );
  NANDN U13250 ( .A(n12729), .B(n12728), .Z(n12733) );
  NAND U13251 ( .A(n12731), .B(n12730), .Z(n12732) );
  AND U13252 ( .A(n12733), .B(n12732), .Z(n13023) );
  NANDN U13253 ( .A(n12735), .B(n12734), .Z(n12739) );
  NANDN U13254 ( .A(n12737), .B(n12736), .Z(n12738) );
  AND U13255 ( .A(n12739), .B(n12738), .Z(n13010) );
  NANDN U13256 ( .A(n12740), .B(n37294), .Z(n12742) );
  XOR U13257 ( .A(b[47]), .B(a[29]), .Z(n13045) );
  NANDN U13258 ( .A(n37172), .B(n13045), .Z(n12741) );
  AND U13259 ( .A(n12742), .B(n12741), .Z(n13086) );
  NANDN U13260 ( .A(n12743), .B(n30627), .Z(n12745) );
  XOR U13261 ( .A(b[9]), .B(a[67]), .Z(n13048) );
  NANDN U13262 ( .A(n30267), .B(n13048), .Z(n12744) );
  AND U13263 ( .A(n12745), .B(n12744), .Z(n13085) );
  NANDN U13264 ( .A(n12746), .B(n37536), .Z(n12748) );
  XOR U13265 ( .A(b[49]), .B(a[27]), .Z(n13051) );
  NANDN U13266 ( .A(n37432), .B(n13051), .Z(n12747) );
  NAND U13267 ( .A(n12748), .B(n12747), .Z(n13084) );
  XOR U13268 ( .A(n13085), .B(n13084), .Z(n13087) );
  XOR U13269 ( .A(n13086), .B(n13087), .Z(n13199) );
  NANDN U13270 ( .A(n36742), .B(n12749), .Z(n12751) );
  XOR U13271 ( .A(b[43]), .B(a[33]), .Z(n13054) );
  NANDN U13272 ( .A(n36891), .B(n13054), .Z(n12750) );
  AND U13273 ( .A(n12751), .B(n12750), .Z(n13065) );
  NANDN U13274 ( .A(n36991), .B(n12752), .Z(n12754) );
  XOR U13275 ( .A(b[45]), .B(a[31]), .Z(n13057) );
  NANDN U13276 ( .A(n37083), .B(n13057), .Z(n12753) );
  AND U13277 ( .A(n12754), .B(n12753), .Z(n13064) );
  NANDN U13278 ( .A(n30482), .B(n12755), .Z(n12757) );
  XOR U13279 ( .A(b[11]), .B(a[65]), .Z(n13060) );
  NANDN U13280 ( .A(n30891), .B(n13060), .Z(n12756) );
  NAND U13281 ( .A(n12757), .B(n12756), .Z(n13063) );
  XOR U13282 ( .A(n13064), .B(n13063), .Z(n13066) );
  XNOR U13283 ( .A(n13065), .B(n13066), .Z(n13198) );
  XNOR U13284 ( .A(n13199), .B(n13198), .Z(n13200) );
  NANDN U13285 ( .A(n12759), .B(n12758), .Z(n12763) );
  OR U13286 ( .A(n12761), .B(n12760), .Z(n12762) );
  NAND U13287 ( .A(n12763), .B(n12762), .Z(n13201) );
  XNOR U13288 ( .A(n13200), .B(n13201), .Z(n13009) );
  XNOR U13289 ( .A(n13010), .B(n13009), .Z(n13012) );
  NANDN U13290 ( .A(n29499), .B(n12764), .Z(n12766) );
  XOR U13291 ( .A(b[7]), .B(a[69]), .Z(n13069) );
  NANDN U13292 ( .A(n29735), .B(n13069), .Z(n12765) );
  AND U13293 ( .A(n12766), .B(n12765), .Z(n13128) );
  NANDN U13294 ( .A(n37857), .B(n12767), .Z(n12769) );
  XOR U13295 ( .A(b[55]), .B(a[21]), .Z(n13072) );
  NANDN U13296 ( .A(n37911), .B(n13072), .Z(n12768) );
  AND U13297 ( .A(n12769), .B(n12768), .Z(n13127) );
  NANDN U13298 ( .A(n35611), .B(n12770), .Z(n12772) );
  XOR U13299 ( .A(b[35]), .B(a[41]), .Z(n13075) );
  NANDN U13300 ( .A(n35801), .B(n13075), .Z(n12771) );
  NAND U13301 ( .A(n12772), .B(n12771), .Z(n13126) );
  XOR U13302 ( .A(n13127), .B(n13126), .Z(n13129) );
  XOR U13303 ( .A(n13128), .B(n13129), .Z(n13151) );
  NANDN U13304 ( .A(n12774), .B(n12773), .Z(n12778) );
  OR U13305 ( .A(n12776), .B(n12775), .Z(n12777) );
  AND U13306 ( .A(n12778), .B(n12777), .Z(n13150) );
  XNOR U13307 ( .A(n13151), .B(n13150), .Z(n13152) );
  NAND U13308 ( .A(n12780), .B(n12779), .Z(n12784) );
  NANDN U13309 ( .A(n12782), .B(n12781), .Z(n12783) );
  NAND U13310 ( .A(n12784), .B(n12783), .Z(n13153) );
  XNOR U13311 ( .A(n13152), .B(n13153), .Z(n13011) );
  XOR U13312 ( .A(n13012), .B(n13011), .Z(n13022) );
  NANDN U13313 ( .A(n12786), .B(n12785), .Z(n12790) );
  NANDN U13314 ( .A(n12788), .B(n12787), .Z(n12789) );
  AND U13315 ( .A(n12790), .B(n12789), .Z(n13018) );
  NANDN U13316 ( .A(n12792), .B(n12791), .Z(n12796) );
  NANDN U13317 ( .A(n12794), .B(n12793), .Z(n12795) );
  AND U13318 ( .A(n12796), .B(n12795), .Z(n13016) );
  NANDN U13319 ( .A(n33875), .B(n12797), .Z(n12799) );
  XOR U13320 ( .A(b[25]), .B(a[51]), .Z(n13102) );
  NANDN U13321 ( .A(n33994), .B(n13102), .Z(n12798) );
  AND U13322 ( .A(n12799), .B(n12798), .Z(n13221) );
  NANDN U13323 ( .A(n32013), .B(n12800), .Z(n12802) );
  XOR U13324 ( .A(b[17]), .B(a[59]), .Z(n13105) );
  NANDN U13325 ( .A(n32292), .B(n13105), .Z(n12801) );
  AND U13326 ( .A(n12802), .B(n12801), .Z(n13220) );
  NANDN U13327 ( .A(n31536), .B(n12803), .Z(n12805) );
  XOR U13328 ( .A(b[15]), .B(a[61]), .Z(n13108) );
  NANDN U13329 ( .A(n31925), .B(n13108), .Z(n12804) );
  NAND U13330 ( .A(n12805), .B(n12804), .Z(n13219) );
  XOR U13331 ( .A(n13220), .B(n13219), .Z(n13222) );
  XOR U13332 ( .A(n13221), .B(n13222), .Z(n13193) );
  NANDN U13333 ( .A(n37526), .B(n12806), .Z(n12808) );
  XOR U13334 ( .A(b[51]), .B(a[25]), .Z(n13111) );
  NANDN U13335 ( .A(n37605), .B(n13111), .Z(n12807) );
  AND U13336 ( .A(n12808), .B(n12807), .Z(n13245) );
  NANDN U13337 ( .A(n37705), .B(n12809), .Z(n12811) );
  XOR U13338 ( .A(b[53]), .B(a[23]), .Z(n13114) );
  NANDN U13339 ( .A(n37778), .B(n13114), .Z(n12810) );
  AND U13340 ( .A(n12811), .B(n12810), .Z(n13244) );
  NANDN U13341 ( .A(n36210), .B(n12812), .Z(n12814) );
  XOR U13342 ( .A(b[39]), .B(a[37]), .Z(n13117) );
  NANDN U13343 ( .A(n36347), .B(n13117), .Z(n12813) );
  NAND U13344 ( .A(n12814), .B(n12813), .Z(n13243) );
  XOR U13345 ( .A(n13244), .B(n13243), .Z(n13246) );
  XNOR U13346 ( .A(n13245), .B(n13246), .Z(n13192) );
  XNOR U13347 ( .A(n13193), .B(n13192), .Z(n13195) );
  NANDN U13348 ( .A(n12816), .B(n12815), .Z(n12820) );
  OR U13349 ( .A(n12818), .B(n12817), .Z(n12819) );
  AND U13350 ( .A(n12820), .B(n12819), .Z(n13194) );
  XOR U13351 ( .A(n13195), .B(n13194), .Z(n13093) );
  NANDN U13352 ( .A(n12822), .B(n12821), .Z(n12826) );
  OR U13353 ( .A(n12824), .B(n12823), .Z(n12825) );
  AND U13354 ( .A(n12826), .B(n12825), .Z(n13091) );
  NANDN U13355 ( .A(n12828), .B(n12827), .Z(n12832) );
  NANDN U13356 ( .A(n12830), .B(n12829), .Z(n12831) );
  NAND U13357 ( .A(n12832), .B(n12831), .Z(n13090) );
  XNOR U13358 ( .A(n13091), .B(n13090), .Z(n13092) );
  XNOR U13359 ( .A(n13093), .B(n13092), .Z(n13015) );
  XNOR U13360 ( .A(n13016), .B(n13015), .Z(n13017) );
  XNOR U13361 ( .A(n13018), .B(n13017), .Z(n13021) );
  XOR U13362 ( .A(n13022), .B(n13021), .Z(n13024) );
  XNOR U13363 ( .A(n13023), .B(n13024), .Z(n12991) );
  NANDN U13364 ( .A(n12834), .B(n12833), .Z(n12838) );
  NANDN U13365 ( .A(n12836), .B(n12835), .Z(n12837) );
  AND U13366 ( .A(n12838), .B(n12837), .Z(n13005) );
  NANDN U13367 ( .A(n12840), .B(n12839), .Z(n12844) );
  NANDN U13368 ( .A(n12842), .B(n12841), .Z(n12843) );
  AND U13369 ( .A(n12844), .B(n12843), .Z(n13004) );
  NANDN U13370 ( .A(n12846), .B(n12845), .Z(n12850) );
  NAND U13371 ( .A(n12848), .B(n12847), .Z(n12849) );
  AND U13372 ( .A(n12850), .B(n12849), .Z(n13003) );
  XOR U13373 ( .A(n13004), .B(n13003), .Z(n13006) );
  XOR U13374 ( .A(n13005), .B(n13006), .Z(n13030) );
  NANDN U13375 ( .A(n12852), .B(n12851), .Z(n12856) );
  NANDN U13376 ( .A(n12854), .B(n12853), .Z(n12855) );
  AND U13377 ( .A(n12856), .B(n12855), .Z(n13145) );
  NANDN U13378 ( .A(n12858), .B(n12857), .Z(n12862) );
  OR U13379 ( .A(n12860), .B(n12859), .Z(n12861) );
  NAND U13380 ( .A(n12862), .B(n12861), .Z(n13144) );
  XNOR U13381 ( .A(n13145), .B(n13144), .Z(n13147) );
  NANDN U13382 ( .A(n12864), .B(n12863), .Z(n12868) );
  OR U13383 ( .A(n12866), .B(n12865), .Z(n12867) );
  NAND U13384 ( .A(n12868), .B(n12867), .Z(n13098) );
  AND U13385 ( .A(a[75]), .B(b[0]), .Z(n12869) );
  XOR U13386 ( .A(b[1]), .B(n12869), .Z(n12871) );
  NANDN U13387 ( .A(b[0]), .B(a[74]), .Z(n12870) );
  AND U13388 ( .A(n12871), .B(n12870), .Z(n13134) );
  NANDN U13389 ( .A(n38278), .B(n12872), .Z(n12874) );
  XOR U13390 ( .A(b[63]), .B(a[13]), .Z(n13177) );
  NANDN U13391 ( .A(n38279), .B(n13177), .Z(n12873) );
  AND U13392 ( .A(n12874), .B(n12873), .Z(n13133) );
  NANDN U13393 ( .A(n35260), .B(n12875), .Z(n12877) );
  XOR U13394 ( .A(b[33]), .B(a[43]), .Z(n13180) );
  NANDN U13395 ( .A(n35456), .B(n13180), .Z(n12876) );
  NAND U13396 ( .A(n12877), .B(n12876), .Z(n13132) );
  XOR U13397 ( .A(n13133), .B(n13132), .Z(n13135) );
  XNOR U13398 ( .A(n13134), .B(n13135), .Z(n13097) );
  NANDN U13399 ( .A(n37974), .B(n12878), .Z(n12880) );
  XOR U13400 ( .A(b[57]), .B(a[19]), .Z(n13183) );
  NANDN U13401 ( .A(n38031), .B(n13183), .Z(n12879) );
  AND U13402 ( .A(n12880), .B(n12879), .Z(n13158) );
  NANDN U13403 ( .A(n38090), .B(n12881), .Z(n12883) );
  XOR U13404 ( .A(b[59]), .B(a[17]), .Z(n13186) );
  NANDN U13405 ( .A(n38130), .B(n13186), .Z(n12882) );
  AND U13406 ( .A(n12883), .B(n12882), .Z(n13157) );
  NANDN U13407 ( .A(n36480), .B(n12884), .Z(n12886) );
  XOR U13408 ( .A(b[41]), .B(a[35]), .Z(n13189) );
  NANDN U13409 ( .A(n36594), .B(n13189), .Z(n12885) );
  NAND U13410 ( .A(n12886), .B(n12885), .Z(n13156) );
  XOR U13411 ( .A(n13157), .B(n13156), .Z(n13159) );
  XOR U13412 ( .A(n13158), .B(n13159), .Z(n13096) );
  XOR U13413 ( .A(n13097), .B(n13096), .Z(n13099) );
  XOR U13414 ( .A(n13098), .B(n13099), .Z(n13146) );
  XOR U13415 ( .A(n13147), .B(n13146), .Z(n13034) );
  NANDN U13416 ( .A(n12888), .B(n12887), .Z(n12892) );
  NAND U13417 ( .A(n12890), .B(n12889), .Z(n12891) );
  NAND U13418 ( .A(n12892), .B(n12891), .Z(n13033) );
  XNOR U13419 ( .A(n13034), .B(n13033), .Z(n13036) );
  NAND U13420 ( .A(n12894), .B(n12893), .Z(n12898) );
  NANDN U13421 ( .A(n12896), .B(n12895), .Z(n12897) );
  AND U13422 ( .A(n12898), .B(n12897), .Z(n13252) );
  NANDN U13423 ( .A(n12900), .B(n12899), .Z(n12904) );
  OR U13424 ( .A(n12902), .B(n12901), .Z(n12903) );
  AND U13425 ( .A(n12904), .B(n12903), .Z(n13041) );
  NANDN U13426 ( .A(n32996), .B(n12905), .Z(n12907) );
  XOR U13427 ( .A(b[21]), .B(a[55]), .Z(n13204) );
  NANDN U13428 ( .A(n33271), .B(n13204), .Z(n12906) );
  AND U13429 ( .A(n12907), .B(n12906), .Z(n13171) );
  NANDN U13430 ( .A(n33866), .B(n12908), .Z(n12910) );
  XOR U13431 ( .A(b[23]), .B(a[53]), .Z(n13207) );
  NANDN U13432 ( .A(n33644), .B(n13207), .Z(n12909) );
  AND U13433 ( .A(n12910), .B(n12909), .Z(n13169) );
  NANDN U13434 ( .A(n32483), .B(n12911), .Z(n12913) );
  XOR U13435 ( .A(b[19]), .B(a[57]), .Z(n13210) );
  NANDN U13436 ( .A(n32823), .B(n13210), .Z(n12912) );
  NAND U13437 ( .A(n12913), .B(n12912), .Z(n13168) );
  XNOR U13438 ( .A(n13169), .B(n13168), .Z(n13170) );
  XOR U13439 ( .A(n13171), .B(n13170), .Z(n13040) );
  NANDN U13440 ( .A(n34909), .B(n12914), .Z(n12916) );
  XOR U13441 ( .A(b[31]), .B(a[45]), .Z(n13213) );
  NANDN U13442 ( .A(n35145), .B(n13213), .Z(n12915) );
  AND U13443 ( .A(n12916), .B(n12915), .Z(n13081) );
  NANDN U13444 ( .A(n38247), .B(n12917), .Z(n12919) );
  XOR U13445 ( .A(b[61]), .B(a[15]), .Z(n13216) );
  NANDN U13446 ( .A(n38248), .B(n13216), .Z(n12918) );
  AND U13447 ( .A(n12919), .B(n12918), .Z(n13079) );
  AND U13448 ( .A(b[63]), .B(a[11]), .Z(n13078) );
  XNOR U13449 ( .A(n13079), .B(n13078), .Z(n13080) );
  XOR U13450 ( .A(n13081), .B(n13080), .Z(n13039) );
  XNOR U13451 ( .A(n13040), .B(n13039), .Z(n13042) );
  NANDN U13452 ( .A(n12921), .B(n12920), .Z(n12925) );
  OR U13453 ( .A(n12923), .B(n12922), .Z(n12924) );
  AND U13454 ( .A(n12925), .B(n12924), .Z(n13140) );
  NANDN U13455 ( .A(n34223), .B(n12926), .Z(n12928) );
  XOR U13456 ( .A(b[27]), .B(a[49]), .Z(n13225) );
  NANDN U13457 ( .A(n34458), .B(n13225), .Z(n12927) );
  AND U13458 ( .A(n12928), .B(n12927), .Z(n13123) );
  NANDN U13459 ( .A(n34634), .B(n12929), .Z(n12931) );
  XOR U13460 ( .A(b[29]), .B(a[47]), .Z(n13228) );
  NANDN U13461 ( .A(n34722), .B(n13228), .Z(n12930) );
  AND U13462 ( .A(n12931), .B(n12930), .Z(n13121) );
  NANDN U13463 ( .A(n31055), .B(n12932), .Z(n12934) );
  XOR U13464 ( .A(b[13]), .B(a[63]), .Z(n13231) );
  NANDN U13465 ( .A(n31293), .B(n13231), .Z(n12933) );
  NAND U13466 ( .A(n12934), .B(n12933), .Z(n13120) );
  XNOR U13467 ( .A(n13121), .B(n13120), .Z(n13122) );
  XOR U13468 ( .A(n13123), .B(n13122), .Z(n13139) );
  NANDN U13469 ( .A(n28889), .B(n12935), .Z(n12937) );
  XOR U13470 ( .A(a[71]), .B(b[5]), .Z(n13234) );
  NANDN U13471 ( .A(n29138), .B(n13234), .Z(n12936) );
  AND U13472 ( .A(n12937), .B(n12936), .Z(n13165) );
  NANDN U13473 ( .A(n209), .B(n12938), .Z(n12940) );
  XOR U13474 ( .A(a[73]), .B(b[3]), .Z(n13237) );
  NANDN U13475 ( .A(n28941), .B(n13237), .Z(n12939) );
  AND U13476 ( .A(n12940), .B(n12939), .Z(n13163) );
  NANDN U13477 ( .A(n35936), .B(n12941), .Z(n12943) );
  XOR U13478 ( .A(b[37]), .B(a[39]), .Z(n13240) );
  NANDN U13479 ( .A(n36047), .B(n13240), .Z(n12942) );
  NAND U13480 ( .A(n12943), .B(n12942), .Z(n13162) );
  XNOR U13481 ( .A(n13163), .B(n13162), .Z(n13164) );
  XOR U13482 ( .A(n13165), .B(n13164), .Z(n13138) );
  XNOR U13483 ( .A(n13139), .B(n13138), .Z(n13141) );
  XOR U13484 ( .A(n13250), .B(n13249), .Z(n13251) );
  XNOR U13485 ( .A(n13252), .B(n13251), .Z(n13035) );
  XOR U13486 ( .A(n13036), .B(n13035), .Z(n13028) );
  NANDN U13487 ( .A(n12945), .B(n12944), .Z(n12949) );
  NANDN U13488 ( .A(n12947), .B(n12946), .Z(n12948) );
  AND U13489 ( .A(n12949), .B(n12948), .Z(n13027) );
  XNOR U13490 ( .A(n13028), .B(n13027), .Z(n13029) );
  XOR U13491 ( .A(n13030), .B(n13029), .Z(n12992) );
  XNOR U13492 ( .A(n12991), .B(n12992), .Z(n12993) );
  XOR U13493 ( .A(n12994), .B(n12993), .Z(n13256) );
  XNOR U13494 ( .A(n13255), .B(n13256), .Z(n13262) );
  NANDN U13495 ( .A(n12951), .B(n12950), .Z(n12955) );
  NANDN U13496 ( .A(n12953), .B(n12952), .Z(n12954) );
  AND U13497 ( .A(n12955), .B(n12954), .Z(n13260) );
  NANDN U13498 ( .A(n12957), .B(n12956), .Z(n12961) );
  OR U13499 ( .A(n12959), .B(n12958), .Z(n12960) );
  AND U13500 ( .A(n12961), .B(n12960), .Z(n13259) );
  XNOR U13501 ( .A(n13260), .B(n13259), .Z(n13261) );
  XOR U13502 ( .A(n13262), .B(n13261), .Z(n12986) );
  NANDN U13503 ( .A(n12963), .B(n12962), .Z(n12967) );
  NANDN U13504 ( .A(n12965), .B(n12964), .Z(n12966) );
  AND U13505 ( .A(n12967), .B(n12966), .Z(n12985) );
  XNOR U13506 ( .A(n12986), .B(n12985), .Z(n12987) );
  NANDN U13507 ( .A(n12969), .B(n12968), .Z(n12973) );
  NAND U13508 ( .A(n12971), .B(n12970), .Z(n12972) );
  NAND U13509 ( .A(n12973), .B(n12972), .Z(n12988) );
  XNOR U13510 ( .A(n12987), .B(n12988), .Z(n12979) );
  XNOR U13511 ( .A(n12980), .B(n12979), .Z(n12981) );
  XNOR U13512 ( .A(n12982), .B(n12981), .Z(n13265) );
  XNOR U13513 ( .A(sreg[139]), .B(n13265), .Z(n13267) );
  NANDN U13514 ( .A(sreg[138]), .B(n12974), .Z(n12978) );
  NAND U13515 ( .A(n12976), .B(n12975), .Z(n12977) );
  NAND U13516 ( .A(n12978), .B(n12977), .Z(n13266) );
  XNOR U13517 ( .A(n13267), .B(n13266), .Z(c[139]) );
  NANDN U13518 ( .A(n12980), .B(n12979), .Z(n12984) );
  NANDN U13519 ( .A(n12982), .B(n12981), .Z(n12983) );
  AND U13520 ( .A(n12984), .B(n12983), .Z(n13273) );
  NANDN U13521 ( .A(n12986), .B(n12985), .Z(n12990) );
  NANDN U13522 ( .A(n12988), .B(n12987), .Z(n12989) );
  AND U13523 ( .A(n12990), .B(n12989), .Z(n13271) );
  NANDN U13524 ( .A(n12992), .B(n12991), .Z(n12996) );
  NANDN U13525 ( .A(n12994), .B(n12993), .Z(n12995) );
  AND U13526 ( .A(n12996), .B(n12995), .Z(n13553) );
  NANDN U13527 ( .A(n12998), .B(n12997), .Z(n13002) );
  OR U13528 ( .A(n13000), .B(n12999), .Z(n13001) );
  AND U13529 ( .A(n13002), .B(n13001), .Z(n13552) );
  XNOR U13530 ( .A(n13553), .B(n13552), .Z(n13555) );
  NANDN U13531 ( .A(n13004), .B(n13003), .Z(n13008) );
  OR U13532 ( .A(n13006), .B(n13005), .Z(n13007) );
  AND U13533 ( .A(n13008), .B(n13007), .Z(n13290) );
  NANDN U13534 ( .A(n13010), .B(n13009), .Z(n13014) );
  NAND U13535 ( .A(n13012), .B(n13011), .Z(n13013) );
  AND U13536 ( .A(n13014), .B(n13013), .Z(n13289) );
  NANDN U13537 ( .A(n13016), .B(n13015), .Z(n13020) );
  NANDN U13538 ( .A(n13018), .B(n13017), .Z(n13019) );
  AND U13539 ( .A(n13020), .B(n13019), .Z(n13288) );
  XOR U13540 ( .A(n13289), .B(n13288), .Z(n13291) );
  XOR U13541 ( .A(n13290), .B(n13291), .Z(n13547) );
  NANDN U13542 ( .A(n13022), .B(n13021), .Z(n13026) );
  NANDN U13543 ( .A(n13024), .B(n13023), .Z(n13025) );
  NAND U13544 ( .A(n13026), .B(n13025), .Z(n13546) );
  XNOR U13545 ( .A(n13547), .B(n13546), .Z(n13548) );
  NANDN U13546 ( .A(n13028), .B(n13027), .Z(n13032) );
  NANDN U13547 ( .A(n13030), .B(n13029), .Z(n13031) );
  AND U13548 ( .A(n13032), .B(n13031), .Z(n13285) );
  NANDN U13549 ( .A(n13034), .B(n13033), .Z(n13038) );
  NAND U13550 ( .A(n13036), .B(n13035), .Z(n13037) );
  AND U13551 ( .A(n13038), .B(n13037), .Z(n13296) );
  NAND U13552 ( .A(n13040), .B(n13039), .Z(n13044) );
  NANDN U13553 ( .A(n13042), .B(n13041), .Z(n13043) );
  AND U13554 ( .A(n13044), .B(n13043), .Z(n13307) );
  NANDN U13555 ( .A(n211), .B(n13045), .Z(n13047) );
  XOR U13556 ( .A(b[47]), .B(a[30]), .Z(n13405) );
  NANDN U13557 ( .A(n37172), .B(n13405), .Z(n13046) );
  AND U13558 ( .A(n13047), .B(n13046), .Z(n13395) );
  NANDN U13559 ( .A(n210), .B(n13048), .Z(n13050) );
  XOR U13560 ( .A(b[9]), .B(a[68]), .Z(n13408) );
  NANDN U13561 ( .A(n30267), .B(n13408), .Z(n13049) );
  AND U13562 ( .A(n13050), .B(n13049), .Z(n13394) );
  NANDN U13563 ( .A(n212), .B(n13051), .Z(n13053) );
  XOR U13564 ( .A(b[49]), .B(a[28]), .Z(n13411) );
  NANDN U13565 ( .A(n37432), .B(n13411), .Z(n13052) );
  NAND U13566 ( .A(n13053), .B(n13052), .Z(n13393) );
  XOR U13567 ( .A(n13394), .B(n13393), .Z(n13396) );
  XOR U13568 ( .A(n13395), .B(n13396), .Z(n13448) );
  NANDN U13569 ( .A(n36742), .B(n13054), .Z(n13056) );
  XOR U13570 ( .A(b[43]), .B(a[34]), .Z(n13414) );
  NANDN U13571 ( .A(n36891), .B(n13414), .Z(n13055) );
  AND U13572 ( .A(n13056), .B(n13055), .Z(n13425) );
  NANDN U13573 ( .A(n36991), .B(n13057), .Z(n13059) );
  XOR U13574 ( .A(b[45]), .B(a[32]), .Z(n13417) );
  NANDN U13575 ( .A(n37083), .B(n13417), .Z(n13058) );
  AND U13576 ( .A(n13059), .B(n13058), .Z(n13424) );
  NANDN U13577 ( .A(n30482), .B(n13060), .Z(n13062) );
  XOR U13578 ( .A(b[11]), .B(a[66]), .Z(n13420) );
  NANDN U13579 ( .A(n30891), .B(n13420), .Z(n13061) );
  NAND U13580 ( .A(n13062), .B(n13061), .Z(n13423) );
  XOR U13581 ( .A(n13424), .B(n13423), .Z(n13426) );
  XNOR U13582 ( .A(n13425), .B(n13426), .Z(n13447) );
  XNOR U13583 ( .A(n13448), .B(n13447), .Z(n13449) );
  NANDN U13584 ( .A(n13064), .B(n13063), .Z(n13068) );
  OR U13585 ( .A(n13066), .B(n13065), .Z(n13067) );
  NAND U13586 ( .A(n13068), .B(n13067), .Z(n13450) );
  XNOR U13587 ( .A(n13449), .B(n13450), .Z(n13306) );
  XNOR U13588 ( .A(n13307), .B(n13306), .Z(n13309) );
  NANDN U13589 ( .A(n29499), .B(n13069), .Z(n13071) );
  XOR U13590 ( .A(b[7]), .B(a[70]), .Z(n13378) );
  NANDN U13591 ( .A(n29735), .B(n13378), .Z(n13070) );
  AND U13592 ( .A(n13071), .B(n13070), .Z(n13368) );
  NANDN U13593 ( .A(n37857), .B(n13072), .Z(n13074) );
  XOR U13594 ( .A(b[55]), .B(a[22]), .Z(n13381) );
  NANDN U13595 ( .A(n37911), .B(n13381), .Z(n13073) );
  AND U13596 ( .A(n13074), .B(n13073), .Z(n13367) );
  NANDN U13597 ( .A(n35611), .B(n13075), .Z(n13077) );
  XOR U13598 ( .A(b[35]), .B(a[42]), .Z(n13384) );
  NANDN U13599 ( .A(n35801), .B(n13384), .Z(n13076) );
  NAND U13600 ( .A(n13077), .B(n13076), .Z(n13366) );
  XOR U13601 ( .A(n13367), .B(n13366), .Z(n13369) );
  XOR U13602 ( .A(n13368), .B(n13369), .Z(n13430) );
  NANDN U13603 ( .A(n13079), .B(n13078), .Z(n13083) );
  NANDN U13604 ( .A(n13081), .B(n13080), .Z(n13082) );
  AND U13605 ( .A(n13083), .B(n13082), .Z(n13429) );
  XNOR U13606 ( .A(n13430), .B(n13429), .Z(n13431) );
  NANDN U13607 ( .A(n13085), .B(n13084), .Z(n13089) );
  OR U13608 ( .A(n13087), .B(n13086), .Z(n13088) );
  NAND U13609 ( .A(n13089), .B(n13088), .Z(n13432) );
  XNOR U13610 ( .A(n13431), .B(n13432), .Z(n13308) );
  XOR U13611 ( .A(n13309), .B(n13308), .Z(n13295) );
  NANDN U13612 ( .A(n13091), .B(n13090), .Z(n13095) );
  NANDN U13613 ( .A(n13093), .B(n13092), .Z(n13094) );
  AND U13614 ( .A(n13095), .B(n13094), .Z(n13303) );
  NAND U13615 ( .A(n13097), .B(n13096), .Z(n13101) );
  NAND U13616 ( .A(n13099), .B(n13098), .Z(n13100) );
  AND U13617 ( .A(n13101), .B(n13100), .Z(n13301) );
  NANDN U13618 ( .A(n33875), .B(n13102), .Z(n13104) );
  XOR U13619 ( .A(b[25]), .B(a[52]), .Z(n13342) );
  NANDN U13620 ( .A(n33994), .B(n13342), .Z(n13103) );
  AND U13621 ( .A(n13104), .B(n13103), .Z(n13470) );
  NANDN U13622 ( .A(n32013), .B(n13105), .Z(n13107) );
  XOR U13623 ( .A(b[17]), .B(a[60]), .Z(n13345) );
  NANDN U13624 ( .A(n32292), .B(n13345), .Z(n13106) );
  AND U13625 ( .A(n13107), .B(n13106), .Z(n13469) );
  NANDN U13626 ( .A(n31536), .B(n13108), .Z(n13110) );
  XOR U13627 ( .A(b[15]), .B(a[62]), .Z(n13348) );
  NANDN U13628 ( .A(n31925), .B(n13348), .Z(n13109) );
  NAND U13629 ( .A(n13110), .B(n13109), .Z(n13468) );
  XOR U13630 ( .A(n13469), .B(n13468), .Z(n13471) );
  XOR U13631 ( .A(n13470), .B(n13471), .Z(n13535) );
  NANDN U13632 ( .A(n37526), .B(n13111), .Z(n13113) );
  XOR U13633 ( .A(b[51]), .B(a[26]), .Z(n13351) );
  NANDN U13634 ( .A(n37605), .B(n13351), .Z(n13112) );
  AND U13635 ( .A(n13113), .B(n13112), .Z(n13494) );
  NANDN U13636 ( .A(n37705), .B(n13114), .Z(n13116) );
  XOR U13637 ( .A(b[53]), .B(a[24]), .Z(n13354) );
  NANDN U13638 ( .A(n37778), .B(n13354), .Z(n13115) );
  AND U13639 ( .A(n13116), .B(n13115), .Z(n13493) );
  NANDN U13640 ( .A(n36210), .B(n13117), .Z(n13119) );
  XOR U13641 ( .A(b[39]), .B(a[38]), .Z(n13357) );
  NANDN U13642 ( .A(n36347), .B(n13357), .Z(n13118) );
  NAND U13643 ( .A(n13119), .B(n13118), .Z(n13492) );
  XOR U13644 ( .A(n13493), .B(n13492), .Z(n13495) );
  XNOR U13645 ( .A(n13494), .B(n13495), .Z(n13534) );
  XNOR U13646 ( .A(n13535), .B(n13534), .Z(n13537) );
  NANDN U13647 ( .A(n13121), .B(n13120), .Z(n13125) );
  NANDN U13648 ( .A(n13123), .B(n13122), .Z(n13124) );
  AND U13649 ( .A(n13125), .B(n13124), .Z(n13536) );
  XOR U13650 ( .A(n13537), .B(n13536), .Z(n13333) );
  NANDN U13651 ( .A(n13127), .B(n13126), .Z(n13131) );
  OR U13652 ( .A(n13129), .B(n13128), .Z(n13130) );
  AND U13653 ( .A(n13131), .B(n13130), .Z(n13331) );
  NANDN U13654 ( .A(n13133), .B(n13132), .Z(n13137) );
  NANDN U13655 ( .A(n13135), .B(n13134), .Z(n13136) );
  NAND U13656 ( .A(n13137), .B(n13136), .Z(n13330) );
  XNOR U13657 ( .A(n13331), .B(n13330), .Z(n13332) );
  XNOR U13658 ( .A(n13333), .B(n13332), .Z(n13300) );
  XNOR U13659 ( .A(n13301), .B(n13300), .Z(n13302) );
  XNOR U13660 ( .A(n13303), .B(n13302), .Z(n13294) );
  XOR U13661 ( .A(n13295), .B(n13294), .Z(n13297) );
  XNOR U13662 ( .A(n13296), .B(n13297), .Z(n13282) );
  NAND U13663 ( .A(n13139), .B(n13138), .Z(n13143) );
  NANDN U13664 ( .A(n13141), .B(n13140), .Z(n13142) );
  NAND U13665 ( .A(n13143), .B(n13142), .Z(n13312) );
  NANDN U13666 ( .A(n13145), .B(n13144), .Z(n13149) );
  NAND U13667 ( .A(n13147), .B(n13146), .Z(n13148) );
  AND U13668 ( .A(n13149), .B(n13148), .Z(n13313) );
  XOR U13669 ( .A(n13312), .B(n13313), .Z(n13315) );
  NANDN U13670 ( .A(n13151), .B(n13150), .Z(n13155) );
  NANDN U13671 ( .A(n13153), .B(n13152), .Z(n13154) );
  NAND U13672 ( .A(n13155), .B(n13154), .Z(n13314) );
  XOR U13673 ( .A(n13315), .B(n13314), .Z(n13321) );
  NANDN U13674 ( .A(n13157), .B(n13156), .Z(n13161) );
  OR U13675 ( .A(n13159), .B(n13158), .Z(n13160) );
  AND U13676 ( .A(n13161), .B(n13160), .Z(n13442) );
  NANDN U13677 ( .A(n13163), .B(n13162), .Z(n13167) );
  NANDN U13678 ( .A(n13165), .B(n13164), .Z(n13166) );
  NAND U13679 ( .A(n13167), .B(n13166), .Z(n13441) );
  XNOR U13680 ( .A(n13442), .B(n13441), .Z(n13444) );
  NANDN U13681 ( .A(n13169), .B(n13168), .Z(n13173) );
  NANDN U13682 ( .A(n13171), .B(n13170), .Z(n13172) );
  AND U13683 ( .A(n13173), .B(n13172), .Z(n13339) );
  NAND U13684 ( .A(b[0]), .B(a[76]), .Z(n13174) );
  XNOR U13685 ( .A(b[1]), .B(n13174), .Z(n13176) );
  NANDN U13686 ( .A(b[0]), .B(a[75]), .Z(n13175) );
  NAND U13687 ( .A(n13176), .B(n13175), .Z(n13375) );
  NANDN U13688 ( .A(n38278), .B(n13177), .Z(n13179) );
  XOR U13689 ( .A(b[63]), .B(a[14]), .Z(n13516) );
  NANDN U13690 ( .A(n38279), .B(n13516), .Z(n13178) );
  AND U13691 ( .A(n13179), .B(n13178), .Z(n13373) );
  NANDN U13692 ( .A(n35260), .B(n13180), .Z(n13182) );
  XOR U13693 ( .A(b[33]), .B(a[44]), .Z(n13519) );
  NANDN U13694 ( .A(n35456), .B(n13519), .Z(n13181) );
  NAND U13695 ( .A(n13182), .B(n13181), .Z(n13372) );
  XNOR U13696 ( .A(n13373), .B(n13372), .Z(n13374) );
  XNOR U13697 ( .A(n13375), .B(n13374), .Z(n13336) );
  NANDN U13698 ( .A(n37974), .B(n13183), .Z(n13185) );
  XOR U13699 ( .A(b[57]), .B(a[20]), .Z(n13525) );
  NANDN U13700 ( .A(n38031), .B(n13525), .Z(n13184) );
  AND U13701 ( .A(n13185), .B(n13184), .Z(n13501) );
  NANDN U13702 ( .A(n38090), .B(n13186), .Z(n13188) );
  XOR U13703 ( .A(b[59]), .B(a[18]), .Z(n13528) );
  NANDN U13704 ( .A(n38130), .B(n13528), .Z(n13187) );
  AND U13705 ( .A(n13188), .B(n13187), .Z(n13499) );
  NANDN U13706 ( .A(n36480), .B(n13189), .Z(n13191) );
  XOR U13707 ( .A(b[41]), .B(a[36]), .Z(n13531) );
  NANDN U13708 ( .A(n36594), .B(n13531), .Z(n13190) );
  NAND U13709 ( .A(n13191), .B(n13190), .Z(n13498) );
  XNOR U13710 ( .A(n13499), .B(n13498), .Z(n13500) );
  XOR U13711 ( .A(n13501), .B(n13500), .Z(n13337) );
  XNOR U13712 ( .A(n13336), .B(n13337), .Z(n13338) );
  XNOR U13713 ( .A(n13339), .B(n13338), .Z(n13443) );
  XOR U13714 ( .A(n13444), .B(n13443), .Z(n13325) );
  NANDN U13715 ( .A(n13193), .B(n13192), .Z(n13197) );
  NAND U13716 ( .A(n13195), .B(n13194), .Z(n13196) );
  NAND U13717 ( .A(n13197), .B(n13196), .Z(n13324) );
  XNOR U13718 ( .A(n13325), .B(n13324), .Z(n13327) );
  NANDN U13719 ( .A(n13199), .B(n13198), .Z(n13203) );
  NANDN U13720 ( .A(n13201), .B(n13200), .Z(n13202) );
  AND U13721 ( .A(n13203), .B(n13202), .Z(n13543) );
  NANDN U13722 ( .A(n32996), .B(n13204), .Z(n13206) );
  XOR U13723 ( .A(b[21]), .B(a[56]), .Z(n13453) );
  NANDN U13724 ( .A(n33271), .B(n13453), .Z(n13205) );
  AND U13725 ( .A(n13206), .B(n13205), .Z(n13512) );
  NANDN U13726 ( .A(n33866), .B(n13207), .Z(n13209) );
  XOR U13727 ( .A(b[23]), .B(a[54]), .Z(n13456) );
  NANDN U13728 ( .A(n33644), .B(n13456), .Z(n13208) );
  AND U13729 ( .A(n13209), .B(n13208), .Z(n13511) );
  NANDN U13730 ( .A(n32483), .B(n13210), .Z(n13212) );
  XOR U13731 ( .A(b[19]), .B(a[58]), .Z(n13459) );
  NANDN U13732 ( .A(n32823), .B(n13459), .Z(n13211) );
  NAND U13733 ( .A(n13212), .B(n13211), .Z(n13510) );
  XOR U13734 ( .A(n13511), .B(n13510), .Z(n13513) );
  XOR U13735 ( .A(n13512), .B(n13513), .Z(n13400) );
  NANDN U13736 ( .A(n34909), .B(n13213), .Z(n13215) );
  XOR U13737 ( .A(b[31]), .B(a[46]), .Z(n13462) );
  NANDN U13738 ( .A(n35145), .B(n13462), .Z(n13214) );
  AND U13739 ( .A(n13215), .B(n13214), .Z(n13389) );
  NANDN U13740 ( .A(n38247), .B(n13216), .Z(n13218) );
  XOR U13741 ( .A(b[61]), .B(a[16]), .Z(n13465) );
  NANDN U13742 ( .A(n38248), .B(n13465), .Z(n13217) );
  AND U13743 ( .A(n13218), .B(n13217), .Z(n13388) );
  AND U13744 ( .A(b[63]), .B(a[12]), .Z(n13387) );
  XOR U13745 ( .A(n13388), .B(n13387), .Z(n13390) );
  XNOR U13746 ( .A(n13389), .B(n13390), .Z(n13399) );
  XNOR U13747 ( .A(n13400), .B(n13399), .Z(n13401) );
  NANDN U13748 ( .A(n13220), .B(n13219), .Z(n13224) );
  OR U13749 ( .A(n13222), .B(n13221), .Z(n13223) );
  NAND U13750 ( .A(n13224), .B(n13223), .Z(n13402) );
  XNOR U13751 ( .A(n13401), .B(n13402), .Z(n13540) );
  NANDN U13752 ( .A(n34223), .B(n13225), .Z(n13227) );
  XOR U13753 ( .A(b[27]), .B(a[50]), .Z(n13474) );
  NANDN U13754 ( .A(n34458), .B(n13474), .Z(n13226) );
  AND U13755 ( .A(n13227), .B(n13226), .Z(n13362) );
  NANDN U13756 ( .A(n34634), .B(n13228), .Z(n13230) );
  XOR U13757 ( .A(b[29]), .B(a[48]), .Z(n13477) );
  NANDN U13758 ( .A(n34722), .B(n13477), .Z(n13229) );
  AND U13759 ( .A(n13230), .B(n13229), .Z(n13361) );
  NANDN U13760 ( .A(n31055), .B(n13231), .Z(n13233) );
  XOR U13761 ( .A(b[13]), .B(a[64]), .Z(n13480) );
  NANDN U13762 ( .A(n31293), .B(n13480), .Z(n13232) );
  NAND U13763 ( .A(n13233), .B(n13232), .Z(n13360) );
  XOR U13764 ( .A(n13361), .B(n13360), .Z(n13363) );
  XOR U13765 ( .A(n13362), .B(n13363), .Z(n13436) );
  NANDN U13766 ( .A(n28889), .B(n13234), .Z(n13236) );
  XOR U13767 ( .A(a[72]), .B(b[5]), .Z(n13483) );
  NANDN U13768 ( .A(n29138), .B(n13483), .Z(n13235) );
  AND U13769 ( .A(n13236), .B(n13235), .Z(n13506) );
  NANDN U13770 ( .A(n209), .B(n13237), .Z(n13239) );
  XOR U13771 ( .A(a[74]), .B(b[3]), .Z(n13486) );
  NANDN U13772 ( .A(n28941), .B(n13486), .Z(n13238) );
  AND U13773 ( .A(n13239), .B(n13238), .Z(n13505) );
  NANDN U13774 ( .A(n35936), .B(n13240), .Z(n13242) );
  XOR U13775 ( .A(b[37]), .B(a[40]), .Z(n13489) );
  NANDN U13776 ( .A(n36047), .B(n13489), .Z(n13241) );
  NAND U13777 ( .A(n13242), .B(n13241), .Z(n13504) );
  XOR U13778 ( .A(n13505), .B(n13504), .Z(n13507) );
  XNOR U13779 ( .A(n13506), .B(n13507), .Z(n13435) );
  XNOR U13780 ( .A(n13436), .B(n13435), .Z(n13437) );
  NANDN U13781 ( .A(n13244), .B(n13243), .Z(n13248) );
  OR U13782 ( .A(n13246), .B(n13245), .Z(n13247) );
  NAND U13783 ( .A(n13248), .B(n13247), .Z(n13438) );
  XOR U13784 ( .A(n13437), .B(n13438), .Z(n13541) );
  XNOR U13785 ( .A(n13540), .B(n13541), .Z(n13542) );
  XNOR U13786 ( .A(n13543), .B(n13542), .Z(n13326) );
  XOR U13787 ( .A(n13327), .B(n13326), .Z(n13319) );
  XNOR U13788 ( .A(n13319), .B(n13318), .Z(n13320) );
  XOR U13789 ( .A(n13321), .B(n13320), .Z(n13283) );
  XNOR U13790 ( .A(n13282), .B(n13283), .Z(n13284) );
  XOR U13791 ( .A(n13285), .B(n13284), .Z(n13549) );
  XNOR U13792 ( .A(n13548), .B(n13549), .Z(n13554) );
  XOR U13793 ( .A(n13555), .B(n13554), .Z(n13277) );
  NANDN U13794 ( .A(n13254), .B(n13253), .Z(n13258) );
  NANDN U13795 ( .A(n13256), .B(n13255), .Z(n13257) );
  AND U13796 ( .A(n13258), .B(n13257), .Z(n13276) );
  XNOR U13797 ( .A(n13277), .B(n13276), .Z(n13278) );
  NANDN U13798 ( .A(n13260), .B(n13259), .Z(n13264) );
  NAND U13799 ( .A(n13262), .B(n13261), .Z(n13263) );
  NAND U13800 ( .A(n13264), .B(n13263), .Z(n13279) );
  XNOR U13801 ( .A(n13278), .B(n13279), .Z(n13270) );
  XNOR U13802 ( .A(n13271), .B(n13270), .Z(n13272) );
  XNOR U13803 ( .A(n13273), .B(n13272), .Z(n13558) );
  XNOR U13804 ( .A(sreg[140]), .B(n13558), .Z(n13560) );
  NANDN U13805 ( .A(sreg[139]), .B(n13265), .Z(n13269) );
  NAND U13806 ( .A(n13267), .B(n13266), .Z(n13268) );
  NAND U13807 ( .A(n13269), .B(n13268), .Z(n13559) );
  XNOR U13808 ( .A(n13560), .B(n13559), .Z(c[140]) );
  NANDN U13809 ( .A(n13271), .B(n13270), .Z(n13275) );
  NANDN U13810 ( .A(n13273), .B(n13272), .Z(n13274) );
  AND U13811 ( .A(n13275), .B(n13274), .Z(n13566) );
  NANDN U13812 ( .A(n13277), .B(n13276), .Z(n13281) );
  NANDN U13813 ( .A(n13279), .B(n13278), .Z(n13280) );
  AND U13814 ( .A(n13281), .B(n13280), .Z(n13564) );
  NANDN U13815 ( .A(n13283), .B(n13282), .Z(n13287) );
  NANDN U13816 ( .A(n13285), .B(n13284), .Z(n13286) );
  AND U13817 ( .A(n13287), .B(n13286), .Z(n13846) );
  NANDN U13818 ( .A(n13289), .B(n13288), .Z(n13293) );
  OR U13819 ( .A(n13291), .B(n13290), .Z(n13292) );
  AND U13820 ( .A(n13293), .B(n13292), .Z(n13845) );
  XNOR U13821 ( .A(n13846), .B(n13845), .Z(n13848) );
  NANDN U13822 ( .A(n13295), .B(n13294), .Z(n13299) );
  NANDN U13823 ( .A(n13297), .B(n13296), .Z(n13298) );
  AND U13824 ( .A(n13299), .B(n13298), .Z(n13840) );
  NANDN U13825 ( .A(n13301), .B(n13300), .Z(n13305) );
  NANDN U13826 ( .A(n13303), .B(n13302), .Z(n13304) );
  AND U13827 ( .A(n13305), .B(n13304), .Z(n13582) );
  NANDN U13828 ( .A(n13307), .B(n13306), .Z(n13311) );
  NAND U13829 ( .A(n13309), .B(n13308), .Z(n13310) );
  AND U13830 ( .A(n13311), .B(n13310), .Z(n13581) );
  XNOR U13831 ( .A(n13582), .B(n13581), .Z(n13583) );
  NAND U13832 ( .A(n13313), .B(n13312), .Z(n13317) );
  NAND U13833 ( .A(n13315), .B(n13314), .Z(n13316) );
  NAND U13834 ( .A(n13317), .B(n13316), .Z(n13584) );
  XNOR U13835 ( .A(n13583), .B(n13584), .Z(n13839) );
  XNOR U13836 ( .A(n13840), .B(n13839), .Z(n13841) );
  NANDN U13837 ( .A(n13319), .B(n13318), .Z(n13323) );
  NANDN U13838 ( .A(n13321), .B(n13320), .Z(n13322) );
  AND U13839 ( .A(n13323), .B(n13322), .Z(n13578) );
  NANDN U13840 ( .A(n13325), .B(n13324), .Z(n13329) );
  NAND U13841 ( .A(n13327), .B(n13326), .Z(n13328) );
  AND U13842 ( .A(n13329), .B(n13328), .Z(n13607) );
  NANDN U13843 ( .A(n13331), .B(n13330), .Z(n13335) );
  NANDN U13844 ( .A(n13333), .B(n13332), .Z(n13334) );
  AND U13845 ( .A(n13335), .B(n13334), .Z(n13601) );
  NANDN U13846 ( .A(n13337), .B(n13336), .Z(n13341) );
  NANDN U13847 ( .A(n13339), .B(n13338), .Z(n13340) );
  AND U13848 ( .A(n13341), .B(n13340), .Z(n13600) );
  NANDN U13849 ( .A(n33875), .B(n13342), .Z(n13344) );
  XOR U13850 ( .A(b[25]), .B(a[53]), .Z(n13680) );
  NANDN U13851 ( .A(n33994), .B(n13680), .Z(n13343) );
  AND U13852 ( .A(n13344), .B(n13343), .Z(n13805) );
  NANDN U13853 ( .A(n32013), .B(n13345), .Z(n13347) );
  XOR U13854 ( .A(b[17]), .B(a[61]), .Z(n13683) );
  NANDN U13855 ( .A(n32292), .B(n13683), .Z(n13346) );
  AND U13856 ( .A(n13347), .B(n13346), .Z(n13804) );
  NANDN U13857 ( .A(n31536), .B(n13348), .Z(n13350) );
  XOR U13858 ( .A(b[15]), .B(a[63]), .Z(n13686) );
  NANDN U13859 ( .A(n31925), .B(n13686), .Z(n13349) );
  NAND U13860 ( .A(n13350), .B(n13349), .Z(n13803) );
  XOR U13861 ( .A(n13804), .B(n13803), .Z(n13806) );
  XOR U13862 ( .A(n13805), .B(n13806), .Z(n13777) );
  NANDN U13863 ( .A(n37526), .B(n13351), .Z(n13353) );
  XOR U13864 ( .A(b[51]), .B(a[27]), .Z(n13689) );
  NANDN U13865 ( .A(n37605), .B(n13689), .Z(n13352) );
  AND U13866 ( .A(n13353), .B(n13352), .Z(n13829) );
  NANDN U13867 ( .A(n37705), .B(n13354), .Z(n13356) );
  XOR U13868 ( .A(b[53]), .B(a[25]), .Z(n13692) );
  NANDN U13869 ( .A(n37778), .B(n13692), .Z(n13355) );
  AND U13870 ( .A(n13356), .B(n13355), .Z(n13828) );
  NANDN U13871 ( .A(n36210), .B(n13357), .Z(n13359) );
  XOR U13872 ( .A(b[39]), .B(a[39]), .Z(n13695) );
  NANDN U13873 ( .A(n36347), .B(n13695), .Z(n13358) );
  NAND U13874 ( .A(n13359), .B(n13358), .Z(n13827) );
  XOR U13875 ( .A(n13828), .B(n13827), .Z(n13830) );
  XNOR U13876 ( .A(n13829), .B(n13830), .Z(n13776) );
  XNOR U13877 ( .A(n13777), .B(n13776), .Z(n13779) );
  NANDN U13878 ( .A(n13361), .B(n13360), .Z(n13365) );
  OR U13879 ( .A(n13363), .B(n13362), .Z(n13364) );
  AND U13880 ( .A(n13365), .B(n13364), .Z(n13778) );
  XOR U13881 ( .A(n13779), .B(n13778), .Z(n13671) );
  NANDN U13882 ( .A(n13367), .B(n13366), .Z(n13371) );
  OR U13883 ( .A(n13369), .B(n13368), .Z(n13370) );
  AND U13884 ( .A(n13371), .B(n13370), .Z(n13669) );
  NANDN U13885 ( .A(n13373), .B(n13372), .Z(n13377) );
  NANDN U13886 ( .A(n13375), .B(n13374), .Z(n13376) );
  NAND U13887 ( .A(n13377), .B(n13376), .Z(n13668) );
  XNOR U13888 ( .A(n13669), .B(n13668), .Z(n13670) );
  XNOR U13889 ( .A(n13671), .B(n13670), .Z(n13599) );
  XOR U13890 ( .A(n13600), .B(n13599), .Z(n13602) );
  XOR U13891 ( .A(n13601), .B(n13602), .Z(n13606) );
  NANDN U13892 ( .A(n29499), .B(n13378), .Z(n13380) );
  XOR U13893 ( .A(b[7]), .B(a[71]), .Z(n13617) );
  NANDN U13894 ( .A(n29735), .B(n13617), .Z(n13379) );
  AND U13895 ( .A(n13380), .B(n13379), .Z(n13706) );
  NANDN U13896 ( .A(n37857), .B(n13381), .Z(n13383) );
  XOR U13897 ( .A(b[55]), .B(a[23]), .Z(n13620) );
  NANDN U13898 ( .A(n37911), .B(n13620), .Z(n13382) );
  AND U13899 ( .A(n13383), .B(n13382), .Z(n13705) );
  NANDN U13900 ( .A(n35611), .B(n13384), .Z(n13386) );
  XOR U13901 ( .A(b[35]), .B(a[43]), .Z(n13623) );
  NANDN U13902 ( .A(n35801), .B(n13623), .Z(n13385) );
  NAND U13903 ( .A(n13386), .B(n13385), .Z(n13704) );
  XOR U13904 ( .A(n13705), .B(n13704), .Z(n13707) );
  XOR U13905 ( .A(n13706), .B(n13707), .Z(n13723) );
  NANDN U13906 ( .A(n13388), .B(n13387), .Z(n13392) );
  OR U13907 ( .A(n13390), .B(n13389), .Z(n13391) );
  AND U13908 ( .A(n13392), .B(n13391), .Z(n13722) );
  XNOR U13909 ( .A(n13723), .B(n13722), .Z(n13724) );
  NANDN U13910 ( .A(n13394), .B(n13393), .Z(n13398) );
  OR U13911 ( .A(n13396), .B(n13395), .Z(n13397) );
  NAND U13912 ( .A(n13398), .B(n13397), .Z(n13725) );
  XNOR U13913 ( .A(n13724), .B(n13725), .Z(n13595) );
  NANDN U13914 ( .A(n13400), .B(n13399), .Z(n13404) );
  NANDN U13915 ( .A(n13402), .B(n13401), .Z(n13403) );
  AND U13916 ( .A(n13404), .B(n13403), .Z(n13594) );
  NANDN U13917 ( .A(n211), .B(n13405), .Z(n13407) );
  XOR U13918 ( .A(b[47]), .B(a[31]), .Z(n13644) );
  NANDN U13919 ( .A(n37172), .B(n13644), .Z(n13406) );
  AND U13920 ( .A(n13407), .B(n13406), .Z(n13634) );
  NANDN U13921 ( .A(n210), .B(n13408), .Z(n13410) );
  XOR U13922 ( .A(b[9]), .B(a[69]), .Z(n13647) );
  NANDN U13923 ( .A(n30267), .B(n13647), .Z(n13409) );
  AND U13924 ( .A(n13410), .B(n13409), .Z(n13633) );
  NANDN U13925 ( .A(n212), .B(n13411), .Z(n13413) );
  XOR U13926 ( .A(b[49]), .B(a[29]), .Z(n13650) );
  NANDN U13927 ( .A(n37432), .B(n13650), .Z(n13412) );
  NAND U13928 ( .A(n13413), .B(n13412), .Z(n13632) );
  XOR U13929 ( .A(n13633), .B(n13632), .Z(n13635) );
  XOR U13930 ( .A(n13634), .B(n13635), .Z(n13783) );
  NANDN U13931 ( .A(n36742), .B(n13414), .Z(n13416) );
  XOR U13932 ( .A(b[43]), .B(a[35]), .Z(n13653) );
  NANDN U13933 ( .A(n36891), .B(n13653), .Z(n13415) );
  AND U13934 ( .A(n13416), .B(n13415), .Z(n13664) );
  NANDN U13935 ( .A(n36991), .B(n13417), .Z(n13419) );
  XOR U13936 ( .A(b[45]), .B(a[33]), .Z(n13656) );
  NANDN U13937 ( .A(n37083), .B(n13656), .Z(n13418) );
  AND U13938 ( .A(n13419), .B(n13418), .Z(n13663) );
  NANDN U13939 ( .A(n30482), .B(n13420), .Z(n13422) );
  XOR U13940 ( .A(b[11]), .B(a[67]), .Z(n13659) );
  NANDN U13941 ( .A(n30891), .B(n13659), .Z(n13421) );
  NAND U13942 ( .A(n13422), .B(n13421), .Z(n13662) );
  XOR U13943 ( .A(n13663), .B(n13662), .Z(n13665) );
  XNOR U13944 ( .A(n13664), .B(n13665), .Z(n13782) );
  XNOR U13945 ( .A(n13783), .B(n13782), .Z(n13784) );
  NANDN U13946 ( .A(n13424), .B(n13423), .Z(n13428) );
  OR U13947 ( .A(n13426), .B(n13425), .Z(n13427) );
  NAND U13948 ( .A(n13428), .B(n13427), .Z(n13785) );
  XNOR U13949 ( .A(n13784), .B(n13785), .Z(n13593) );
  XOR U13950 ( .A(n13594), .B(n13593), .Z(n13596) );
  XNOR U13951 ( .A(n13595), .B(n13596), .Z(n13605) );
  XOR U13952 ( .A(n13606), .B(n13605), .Z(n13608) );
  XOR U13953 ( .A(n13607), .B(n13608), .Z(n13576) );
  NANDN U13954 ( .A(n13430), .B(n13429), .Z(n13434) );
  NANDN U13955 ( .A(n13432), .B(n13431), .Z(n13433) );
  AND U13956 ( .A(n13434), .B(n13433), .Z(n13589) );
  NANDN U13957 ( .A(n13436), .B(n13435), .Z(n13440) );
  NANDN U13958 ( .A(n13438), .B(n13437), .Z(n13439) );
  AND U13959 ( .A(n13440), .B(n13439), .Z(n13588) );
  NANDN U13960 ( .A(n13442), .B(n13441), .Z(n13446) );
  NAND U13961 ( .A(n13444), .B(n13443), .Z(n13445) );
  AND U13962 ( .A(n13446), .B(n13445), .Z(n13587) );
  XOR U13963 ( .A(n13588), .B(n13587), .Z(n13590) );
  XOR U13964 ( .A(n13589), .B(n13590), .Z(n13614) );
  NANDN U13965 ( .A(n13448), .B(n13447), .Z(n13452) );
  NANDN U13966 ( .A(n13450), .B(n13449), .Z(n13451) );
  AND U13967 ( .A(n13452), .B(n13451), .Z(n13836) );
  NANDN U13968 ( .A(n32996), .B(n13453), .Z(n13455) );
  XOR U13969 ( .A(b[21]), .B(a[57]), .Z(n13788) );
  NANDN U13970 ( .A(n33271), .B(n13788), .Z(n13454) );
  AND U13971 ( .A(n13455), .B(n13454), .Z(n13754) );
  NANDN U13972 ( .A(n33866), .B(n13456), .Z(n13458) );
  XOR U13973 ( .A(b[23]), .B(a[55]), .Z(n13791) );
  NANDN U13974 ( .A(n33644), .B(n13791), .Z(n13457) );
  AND U13975 ( .A(n13458), .B(n13457), .Z(n13753) );
  NANDN U13976 ( .A(n32483), .B(n13459), .Z(n13461) );
  XOR U13977 ( .A(b[19]), .B(a[59]), .Z(n13794) );
  NANDN U13978 ( .A(n32823), .B(n13794), .Z(n13460) );
  NAND U13979 ( .A(n13461), .B(n13460), .Z(n13752) );
  XOR U13980 ( .A(n13753), .B(n13752), .Z(n13755) );
  XOR U13981 ( .A(n13754), .B(n13755), .Z(n13639) );
  NANDN U13982 ( .A(n34909), .B(n13462), .Z(n13464) );
  XOR U13983 ( .A(b[31]), .B(a[47]), .Z(n13797) );
  NANDN U13984 ( .A(n35145), .B(n13797), .Z(n13463) );
  AND U13985 ( .A(n13464), .B(n13463), .Z(n13628) );
  NANDN U13986 ( .A(n38247), .B(n13465), .Z(n13467) );
  XOR U13987 ( .A(b[61]), .B(a[17]), .Z(n13800) );
  NANDN U13988 ( .A(n38248), .B(n13800), .Z(n13466) );
  AND U13989 ( .A(n13467), .B(n13466), .Z(n13627) );
  AND U13990 ( .A(b[63]), .B(a[13]), .Z(n13626) );
  XOR U13991 ( .A(n13627), .B(n13626), .Z(n13629) );
  XNOR U13992 ( .A(n13628), .B(n13629), .Z(n13638) );
  XNOR U13993 ( .A(n13639), .B(n13638), .Z(n13640) );
  NANDN U13994 ( .A(n13469), .B(n13468), .Z(n13473) );
  OR U13995 ( .A(n13471), .B(n13470), .Z(n13472) );
  NAND U13996 ( .A(n13473), .B(n13472), .Z(n13641) );
  XNOR U13997 ( .A(n13640), .B(n13641), .Z(n13833) );
  NANDN U13998 ( .A(n34223), .B(n13474), .Z(n13476) );
  XOR U13999 ( .A(b[27]), .B(a[51]), .Z(n13809) );
  NANDN U14000 ( .A(n34458), .B(n13809), .Z(n13475) );
  AND U14001 ( .A(n13476), .B(n13475), .Z(n13700) );
  NANDN U14002 ( .A(n34634), .B(n13477), .Z(n13479) );
  XOR U14003 ( .A(b[29]), .B(a[49]), .Z(n13812) );
  NANDN U14004 ( .A(n34722), .B(n13812), .Z(n13478) );
  AND U14005 ( .A(n13479), .B(n13478), .Z(n13699) );
  NANDN U14006 ( .A(n31055), .B(n13480), .Z(n13482) );
  XOR U14007 ( .A(b[13]), .B(a[65]), .Z(n13815) );
  NANDN U14008 ( .A(n31293), .B(n13815), .Z(n13481) );
  NAND U14009 ( .A(n13482), .B(n13481), .Z(n13698) );
  XOR U14010 ( .A(n13699), .B(n13698), .Z(n13701) );
  XOR U14011 ( .A(n13700), .B(n13701), .Z(n13729) );
  NANDN U14012 ( .A(n28889), .B(n13483), .Z(n13485) );
  XOR U14013 ( .A(a[73]), .B(b[5]), .Z(n13818) );
  NANDN U14014 ( .A(n29138), .B(n13818), .Z(n13484) );
  AND U14015 ( .A(n13485), .B(n13484), .Z(n13748) );
  NANDN U14016 ( .A(n209), .B(n13486), .Z(n13488) );
  XOR U14017 ( .A(a[75]), .B(b[3]), .Z(n13821) );
  NANDN U14018 ( .A(n28941), .B(n13821), .Z(n13487) );
  AND U14019 ( .A(n13488), .B(n13487), .Z(n13747) );
  NANDN U14020 ( .A(n35936), .B(n13489), .Z(n13491) );
  XOR U14021 ( .A(b[37]), .B(a[41]), .Z(n13824) );
  NANDN U14022 ( .A(n36047), .B(n13824), .Z(n13490) );
  NAND U14023 ( .A(n13491), .B(n13490), .Z(n13746) );
  XOR U14024 ( .A(n13747), .B(n13746), .Z(n13749) );
  XNOR U14025 ( .A(n13748), .B(n13749), .Z(n13728) );
  XNOR U14026 ( .A(n13729), .B(n13728), .Z(n13730) );
  NANDN U14027 ( .A(n13493), .B(n13492), .Z(n13497) );
  OR U14028 ( .A(n13495), .B(n13494), .Z(n13496) );
  NAND U14029 ( .A(n13497), .B(n13496), .Z(n13731) );
  XOR U14030 ( .A(n13730), .B(n13731), .Z(n13834) );
  XNOR U14031 ( .A(n13833), .B(n13834), .Z(n13835) );
  XNOR U14032 ( .A(n13836), .B(n13835), .Z(n13719) );
  NANDN U14033 ( .A(n13499), .B(n13498), .Z(n13503) );
  NANDN U14034 ( .A(n13501), .B(n13500), .Z(n13502) );
  AND U14035 ( .A(n13503), .B(n13502), .Z(n13735) );
  NANDN U14036 ( .A(n13505), .B(n13504), .Z(n13509) );
  OR U14037 ( .A(n13507), .B(n13506), .Z(n13508) );
  NAND U14038 ( .A(n13509), .B(n13508), .Z(n13734) );
  XNOR U14039 ( .A(n13735), .B(n13734), .Z(n13737) );
  NANDN U14040 ( .A(n13511), .B(n13510), .Z(n13515) );
  OR U14041 ( .A(n13513), .B(n13512), .Z(n13514) );
  AND U14042 ( .A(n13515), .B(n13514), .Z(n13677) );
  NANDN U14043 ( .A(n38278), .B(n13516), .Z(n13518) );
  XOR U14044 ( .A(b[63]), .B(a[15]), .Z(n13761) );
  NANDN U14045 ( .A(n38279), .B(n13761), .Z(n13517) );
  AND U14046 ( .A(n13518), .B(n13517), .Z(n13711) );
  NANDN U14047 ( .A(n35260), .B(n13519), .Z(n13521) );
  XOR U14048 ( .A(b[33]), .B(a[45]), .Z(n13764) );
  NANDN U14049 ( .A(n35456), .B(n13764), .Z(n13520) );
  NAND U14050 ( .A(n13521), .B(n13520), .Z(n13710) );
  XNOR U14051 ( .A(n13711), .B(n13710), .Z(n13712) );
  NAND U14052 ( .A(b[0]), .B(a[77]), .Z(n13522) );
  XNOR U14053 ( .A(b[1]), .B(n13522), .Z(n13524) );
  NANDN U14054 ( .A(b[0]), .B(a[76]), .Z(n13523) );
  NAND U14055 ( .A(n13524), .B(n13523), .Z(n13713) );
  XNOR U14056 ( .A(n13712), .B(n13713), .Z(n13674) );
  NANDN U14057 ( .A(n37974), .B(n13525), .Z(n13527) );
  XOR U14058 ( .A(b[57]), .B(a[21]), .Z(n13767) );
  NANDN U14059 ( .A(n38031), .B(n13767), .Z(n13526) );
  AND U14060 ( .A(n13527), .B(n13526), .Z(n13743) );
  NANDN U14061 ( .A(n38090), .B(n13528), .Z(n13530) );
  XOR U14062 ( .A(b[59]), .B(a[19]), .Z(n13770) );
  NANDN U14063 ( .A(n38130), .B(n13770), .Z(n13529) );
  AND U14064 ( .A(n13530), .B(n13529), .Z(n13741) );
  NANDN U14065 ( .A(n36480), .B(n13531), .Z(n13533) );
  XOR U14066 ( .A(b[41]), .B(a[37]), .Z(n13773) );
  NANDN U14067 ( .A(n36594), .B(n13773), .Z(n13532) );
  NAND U14068 ( .A(n13533), .B(n13532), .Z(n13740) );
  XNOR U14069 ( .A(n13741), .B(n13740), .Z(n13742) );
  XOR U14070 ( .A(n13743), .B(n13742), .Z(n13675) );
  XNOR U14071 ( .A(n13674), .B(n13675), .Z(n13676) );
  XNOR U14072 ( .A(n13677), .B(n13676), .Z(n13736) );
  XOR U14073 ( .A(n13737), .B(n13736), .Z(n13717) );
  NANDN U14074 ( .A(n13535), .B(n13534), .Z(n13539) );
  NAND U14075 ( .A(n13537), .B(n13536), .Z(n13538) );
  NAND U14076 ( .A(n13539), .B(n13538), .Z(n13716) );
  XNOR U14077 ( .A(n13717), .B(n13716), .Z(n13718) );
  XOR U14078 ( .A(n13719), .B(n13718), .Z(n13612) );
  NANDN U14079 ( .A(n13541), .B(n13540), .Z(n13545) );
  NANDN U14080 ( .A(n13543), .B(n13542), .Z(n13544) );
  AND U14081 ( .A(n13545), .B(n13544), .Z(n13611) );
  XNOR U14082 ( .A(n13612), .B(n13611), .Z(n13613) );
  XNOR U14083 ( .A(n13614), .B(n13613), .Z(n13575) );
  XNOR U14084 ( .A(n13576), .B(n13575), .Z(n13577) );
  XOR U14085 ( .A(n13578), .B(n13577), .Z(n13842) );
  XNOR U14086 ( .A(n13841), .B(n13842), .Z(n13847) );
  XOR U14087 ( .A(n13848), .B(n13847), .Z(n13570) );
  NANDN U14088 ( .A(n13547), .B(n13546), .Z(n13551) );
  NANDN U14089 ( .A(n13549), .B(n13548), .Z(n13550) );
  AND U14090 ( .A(n13551), .B(n13550), .Z(n13569) );
  XNOR U14091 ( .A(n13570), .B(n13569), .Z(n13571) );
  NANDN U14092 ( .A(n13553), .B(n13552), .Z(n13557) );
  NAND U14093 ( .A(n13555), .B(n13554), .Z(n13556) );
  NAND U14094 ( .A(n13557), .B(n13556), .Z(n13572) );
  XNOR U14095 ( .A(n13571), .B(n13572), .Z(n13563) );
  XNOR U14096 ( .A(n13564), .B(n13563), .Z(n13565) );
  XNOR U14097 ( .A(n13566), .B(n13565), .Z(n13851) );
  XNOR U14098 ( .A(sreg[141]), .B(n13851), .Z(n13853) );
  NANDN U14099 ( .A(sreg[140]), .B(n13558), .Z(n13562) );
  NAND U14100 ( .A(n13560), .B(n13559), .Z(n13561) );
  NAND U14101 ( .A(n13562), .B(n13561), .Z(n13852) );
  XNOR U14102 ( .A(n13853), .B(n13852), .Z(c[141]) );
  NANDN U14103 ( .A(n13564), .B(n13563), .Z(n13568) );
  NANDN U14104 ( .A(n13566), .B(n13565), .Z(n13567) );
  AND U14105 ( .A(n13568), .B(n13567), .Z(n13859) );
  NANDN U14106 ( .A(n13570), .B(n13569), .Z(n13574) );
  NANDN U14107 ( .A(n13572), .B(n13571), .Z(n13573) );
  AND U14108 ( .A(n13574), .B(n13573), .Z(n13857) );
  NANDN U14109 ( .A(n13576), .B(n13575), .Z(n13580) );
  NANDN U14110 ( .A(n13578), .B(n13577), .Z(n13579) );
  AND U14111 ( .A(n13580), .B(n13579), .Z(n14139) );
  NANDN U14112 ( .A(n13582), .B(n13581), .Z(n13586) );
  NANDN U14113 ( .A(n13584), .B(n13583), .Z(n13585) );
  NAND U14114 ( .A(n13586), .B(n13585), .Z(n14138) );
  XNOR U14115 ( .A(n14139), .B(n14138), .Z(n14141) );
  NANDN U14116 ( .A(n13588), .B(n13587), .Z(n13592) );
  OR U14117 ( .A(n13590), .B(n13589), .Z(n13591) );
  AND U14118 ( .A(n13592), .B(n13591), .Z(n14128) );
  NANDN U14119 ( .A(n13594), .B(n13593), .Z(n13598) );
  NANDN U14120 ( .A(n13596), .B(n13595), .Z(n13597) );
  AND U14121 ( .A(n13598), .B(n13597), .Z(n14127) );
  NANDN U14122 ( .A(n13600), .B(n13599), .Z(n13604) );
  OR U14123 ( .A(n13602), .B(n13601), .Z(n13603) );
  AND U14124 ( .A(n13604), .B(n13603), .Z(n14126) );
  XOR U14125 ( .A(n14127), .B(n14126), .Z(n14129) );
  XOR U14126 ( .A(n14128), .B(n14129), .Z(n14133) );
  NANDN U14127 ( .A(n13606), .B(n13605), .Z(n13610) );
  OR U14128 ( .A(n13608), .B(n13607), .Z(n13609) );
  AND U14129 ( .A(n13610), .B(n13609), .Z(n14132) );
  XNOR U14130 ( .A(n14133), .B(n14132), .Z(n14134) );
  NANDN U14131 ( .A(n13612), .B(n13611), .Z(n13616) );
  NANDN U14132 ( .A(n13614), .B(n13613), .Z(n13615) );
  AND U14133 ( .A(n13616), .B(n13615), .Z(n14123) );
  NANDN U14134 ( .A(n29499), .B(n13617), .Z(n13619) );
  XOR U14135 ( .A(b[7]), .B(a[72]), .Z(n13904) );
  NANDN U14136 ( .A(n29735), .B(n13904), .Z(n13618) );
  AND U14137 ( .A(n13619), .B(n13618), .Z(n13993) );
  NANDN U14138 ( .A(n37857), .B(n13620), .Z(n13622) );
  XOR U14139 ( .A(b[55]), .B(a[24]), .Z(n13907) );
  NANDN U14140 ( .A(n37911), .B(n13907), .Z(n13621) );
  AND U14141 ( .A(n13622), .B(n13621), .Z(n13992) );
  NANDN U14142 ( .A(n35611), .B(n13623), .Z(n13625) );
  XOR U14143 ( .A(b[35]), .B(a[44]), .Z(n13910) );
  NANDN U14144 ( .A(n35801), .B(n13910), .Z(n13624) );
  NAND U14145 ( .A(n13625), .B(n13624), .Z(n13991) );
  XOR U14146 ( .A(n13992), .B(n13991), .Z(n13994) );
  XOR U14147 ( .A(n13993), .B(n13994), .Z(n14004) );
  NANDN U14148 ( .A(n13627), .B(n13626), .Z(n13631) );
  OR U14149 ( .A(n13629), .B(n13628), .Z(n13630) );
  AND U14150 ( .A(n13631), .B(n13630), .Z(n14003) );
  XNOR U14151 ( .A(n14004), .B(n14003), .Z(n14005) );
  NANDN U14152 ( .A(n13633), .B(n13632), .Z(n13637) );
  OR U14153 ( .A(n13635), .B(n13634), .Z(n13636) );
  NAND U14154 ( .A(n13637), .B(n13636), .Z(n14006) );
  XNOR U14155 ( .A(n14005), .B(n14006), .Z(n13877) );
  NANDN U14156 ( .A(n13639), .B(n13638), .Z(n13643) );
  NANDN U14157 ( .A(n13641), .B(n13640), .Z(n13642) );
  AND U14158 ( .A(n13643), .B(n13642), .Z(n13875) );
  NANDN U14159 ( .A(n211), .B(n13644), .Z(n13646) );
  XOR U14160 ( .A(b[47]), .B(a[32]), .Z(n13931) );
  NANDN U14161 ( .A(n37172), .B(n13931), .Z(n13645) );
  AND U14162 ( .A(n13646), .B(n13645), .Z(n13921) );
  NANDN U14163 ( .A(n210), .B(n13647), .Z(n13649) );
  XOR U14164 ( .A(b[9]), .B(a[70]), .Z(n13934) );
  NANDN U14165 ( .A(n30267), .B(n13934), .Z(n13648) );
  AND U14166 ( .A(n13649), .B(n13648), .Z(n13920) );
  NANDN U14167 ( .A(n212), .B(n13650), .Z(n13652) );
  XOR U14168 ( .A(b[49]), .B(a[30]), .Z(n13937) );
  NANDN U14169 ( .A(n37432), .B(n13937), .Z(n13651) );
  NAND U14170 ( .A(n13652), .B(n13651), .Z(n13919) );
  XOR U14171 ( .A(n13920), .B(n13919), .Z(n13922) );
  XOR U14172 ( .A(n13921), .B(n13922), .Z(n14064) );
  NANDN U14173 ( .A(n36742), .B(n13653), .Z(n13655) );
  XOR U14174 ( .A(b[43]), .B(a[36]), .Z(n13940) );
  NANDN U14175 ( .A(n36891), .B(n13940), .Z(n13654) );
  AND U14176 ( .A(n13655), .B(n13654), .Z(n13951) );
  NANDN U14177 ( .A(n36991), .B(n13656), .Z(n13658) );
  XOR U14178 ( .A(b[45]), .B(a[34]), .Z(n13943) );
  NANDN U14179 ( .A(n37083), .B(n13943), .Z(n13657) );
  AND U14180 ( .A(n13658), .B(n13657), .Z(n13950) );
  NANDN U14181 ( .A(n30482), .B(n13659), .Z(n13661) );
  XOR U14182 ( .A(b[11]), .B(a[68]), .Z(n13946) );
  NANDN U14183 ( .A(n30891), .B(n13946), .Z(n13660) );
  NAND U14184 ( .A(n13661), .B(n13660), .Z(n13949) );
  XOR U14185 ( .A(n13950), .B(n13949), .Z(n13952) );
  XNOR U14186 ( .A(n13951), .B(n13952), .Z(n14063) );
  XNOR U14187 ( .A(n14064), .B(n14063), .Z(n14065) );
  NANDN U14188 ( .A(n13663), .B(n13662), .Z(n13667) );
  OR U14189 ( .A(n13665), .B(n13664), .Z(n13666) );
  NAND U14190 ( .A(n13667), .B(n13666), .Z(n14066) );
  XNOR U14191 ( .A(n14065), .B(n14066), .Z(n13874) );
  XNOR U14192 ( .A(n13875), .B(n13874), .Z(n13876) );
  XOR U14193 ( .A(n13877), .B(n13876), .Z(n13887) );
  NANDN U14194 ( .A(n13669), .B(n13668), .Z(n13673) );
  NANDN U14195 ( .A(n13671), .B(n13670), .Z(n13672) );
  AND U14196 ( .A(n13673), .B(n13672), .Z(n13883) );
  NANDN U14197 ( .A(n13675), .B(n13674), .Z(n13679) );
  NANDN U14198 ( .A(n13677), .B(n13676), .Z(n13678) );
  AND U14199 ( .A(n13679), .B(n13678), .Z(n13881) );
  NANDN U14200 ( .A(n33875), .B(n13680), .Z(n13682) );
  XOR U14201 ( .A(b[25]), .B(a[54]), .Z(n13967) );
  NANDN U14202 ( .A(n33994), .B(n13967), .Z(n13681) );
  AND U14203 ( .A(n13682), .B(n13681), .Z(n14086) );
  NANDN U14204 ( .A(n32013), .B(n13683), .Z(n13685) );
  XOR U14205 ( .A(b[17]), .B(a[62]), .Z(n13970) );
  NANDN U14206 ( .A(n32292), .B(n13970), .Z(n13684) );
  AND U14207 ( .A(n13685), .B(n13684), .Z(n14085) );
  NANDN U14208 ( .A(n31536), .B(n13686), .Z(n13688) );
  XOR U14209 ( .A(b[15]), .B(a[64]), .Z(n13973) );
  NANDN U14210 ( .A(n31925), .B(n13973), .Z(n13687) );
  NAND U14211 ( .A(n13688), .B(n13687), .Z(n14084) );
  XOR U14212 ( .A(n14085), .B(n14084), .Z(n14087) );
  XOR U14213 ( .A(n14086), .B(n14087), .Z(n14058) );
  NANDN U14214 ( .A(n37526), .B(n13689), .Z(n13691) );
  XOR U14215 ( .A(b[51]), .B(a[28]), .Z(n13976) );
  NANDN U14216 ( .A(n37605), .B(n13976), .Z(n13690) );
  AND U14217 ( .A(n13691), .B(n13690), .Z(n14110) );
  NANDN U14218 ( .A(n37705), .B(n13692), .Z(n13694) );
  XOR U14219 ( .A(b[53]), .B(a[26]), .Z(n13979) );
  NANDN U14220 ( .A(n37778), .B(n13979), .Z(n13693) );
  AND U14221 ( .A(n13694), .B(n13693), .Z(n14109) );
  NANDN U14222 ( .A(n36210), .B(n13695), .Z(n13697) );
  XOR U14223 ( .A(b[39]), .B(a[40]), .Z(n13982) );
  NANDN U14224 ( .A(n36347), .B(n13982), .Z(n13696) );
  NAND U14225 ( .A(n13697), .B(n13696), .Z(n14108) );
  XOR U14226 ( .A(n14109), .B(n14108), .Z(n14111) );
  XNOR U14227 ( .A(n14110), .B(n14111), .Z(n14057) );
  XNOR U14228 ( .A(n14058), .B(n14057), .Z(n14060) );
  NANDN U14229 ( .A(n13699), .B(n13698), .Z(n13703) );
  OR U14230 ( .A(n13701), .B(n13700), .Z(n13702) );
  AND U14231 ( .A(n13703), .B(n13702), .Z(n14059) );
  XOR U14232 ( .A(n14060), .B(n14059), .Z(n13958) );
  NANDN U14233 ( .A(n13705), .B(n13704), .Z(n13709) );
  OR U14234 ( .A(n13707), .B(n13706), .Z(n13708) );
  AND U14235 ( .A(n13709), .B(n13708), .Z(n13956) );
  NANDN U14236 ( .A(n13711), .B(n13710), .Z(n13715) );
  NANDN U14237 ( .A(n13713), .B(n13712), .Z(n13714) );
  NAND U14238 ( .A(n13715), .B(n13714), .Z(n13955) );
  XNOR U14239 ( .A(n13956), .B(n13955), .Z(n13957) );
  XNOR U14240 ( .A(n13958), .B(n13957), .Z(n13880) );
  XNOR U14241 ( .A(n13881), .B(n13880), .Z(n13882) );
  XNOR U14242 ( .A(n13883), .B(n13882), .Z(n13886) );
  XNOR U14243 ( .A(n13887), .B(n13886), .Z(n13888) );
  NANDN U14244 ( .A(n13717), .B(n13716), .Z(n13721) );
  NAND U14245 ( .A(n13719), .B(n13718), .Z(n13720) );
  NAND U14246 ( .A(n13721), .B(n13720), .Z(n13889) );
  XNOR U14247 ( .A(n13888), .B(n13889), .Z(n14120) );
  NANDN U14248 ( .A(n13723), .B(n13722), .Z(n13727) );
  NANDN U14249 ( .A(n13725), .B(n13724), .Z(n13726) );
  AND U14250 ( .A(n13727), .B(n13726), .Z(n13870) );
  NANDN U14251 ( .A(n13729), .B(n13728), .Z(n13733) );
  NANDN U14252 ( .A(n13731), .B(n13730), .Z(n13732) );
  AND U14253 ( .A(n13733), .B(n13732), .Z(n13869) );
  NANDN U14254 ( .A(n13735), .B(n13734), .Z(n13739) );
  NAND U14255 ( .A(n13737), .B(n13736), .Z(n13738) );
  AND U14256 ( .A(n13739), .B(n13738), .Z(n13868) );
  XOR U14257 ( .A(n13869), .B(n13868), .Z(n13871) );
  XOR U14258 ( .A(n13870), .B(n13871), .Z(n13895) );
  NANDN U14259 ( .A(n13741), .B(n13740), .Z(n13745) );
  NANDN U14260 ( .A(n13743), .B(n13742), .Z(n13744) );
  AND U14261 ( .A(n13745), .B(n13744), .Z(n14016) );
  NANDN U14262 ( .A(n13747), .B(n13746), .Z(n13751) );
  OR U14263 ( .A(n13749), .B(n13748), .Z(n13750) );
  NAND U14264 ( .A(n13751), .B(n13750), .Z(n14015) );
  XNOR U14265 ( .A(n14016), .B(n14015), .Z(n14018) );
  NANDN U14266 ( .A(n13753), .B(n13752), .Z(n13757) );
  OR U14267 ( .A(n13755), .B(n13754), .Z(n13756) );
  AND U14268 ( .A(n13757), .B(n13756), .Z(n13964) );
  NAND U14269 ( .A(b[0]), .B(a[78]), .Z(n13758) );
  XNOR U14270 ( .A(b[1]), .B(n13758), .Z(n13760) );
  NANDN U14271 ( .A(b[0]), .B(a[77]), .Z(n13759) );
  NAND U14272 ( .A(n13760), .B(n13759), .Z(n14000) );
  NANDN U14273 ( .A(n38278), .B(n13761), .Z(n13763) );
  XOR U14274 ( .A(b[63]), .B(a[16]), .Z(n14039) );
  NANDN U14275 ( .A(n38279), .B(n14039), .Z(n13762) );
  AND U14276 ( .A(n13763), .B(n13762), .Z(n13998) );
  NANDN U14277 ( .A(n35260), .B(n13764), .Z(n13766) );
  XOR U14278 ( .A(b[33]), .B(a[46]), .Z(n14042) );
  NANDN U14279 ( .A(n35456), .B(n14042), .Z(n13765) );
  NAND U14280 ( .A(n13766), .B(n13765), .Z(n13997) );
  XNOR U14281 ( .A(n13998), .B(n13997), .Z(n13999) );
  XNOR U14282 ( .A(n14000), .B(n13999), .Z(n13961) );
  NANDN U14283 ( .A(n37974), .B(n13767), .Z(n13769) );
  XOR U14284 ( .A(b[57]), .B(a[22]), .Z(n14048) );
  NANDN U14285 ( .A(n38031), .B(n14048), .Z(n13768) );
  AND U14286 ( .A(n13769), .B(n13768), .Z(n14024) );
  NANDN U14287 ( .A(n38090), .B(n13770), .Z(n13772) );
  XOR U14288 ( .A(b[59]), .B(a[20]), .Z(n14051) );
  NANDN U14289 ( .A(n38130), .B(n14051), .Z(n13771) );
  AND U14290 ( .A(n13772), .B(n13771), .Z(n14022) );
  NANDN U14291 ( .A(n36480), .B(n13773), .Z(n13775) );
  XOR U14292 ( .A(b[41]), .B(a[38]), .Z(n14054) );
  NANDN U14293 ( .A(n36594), .B(n14054), .Z(n13774) );
  NAND U14294 ( .A(n13775), .B(n13774), .Z(n14021) );
  XNOR U14295 ( .A(n14022), .B(n14021), .Z(n14023) );
  XOR U14296 ( .A(n14024), .B(n14023), .Z(n13962) );
  XNOR U14297 ( .A(n13961), .B(n13962), .Z(n13963) );
  XNOR U14298 ( .A(n13964), .B(n13963), .Z(n14017) );
  XOR U14299 ( .A(n14018), .B(n14017), .Z(n13899) );
  NANDN U14300 ( .A(n13777), .B(n13776), .Z(n13781) );
  NAND U14301 ( .A(n13779), .B(n13778), .Z(n13780) );
  NAND U14302 ( .A(n13781), .B(n13780), .Z(n13898) );
  XNOR U14303 ( .A(n13899), .B(n13898), .Z(n13901) );
  NANDN U14304 ( .A(n13783), .B(n13782), .Z(n13787) );
  NANDN U14305 ( .A(n13785), .B(n13784), .Z(n13786) );
  AND U14306 ( .A(n13787), .B(n13786), .Z(n14117) );
  NANDN U14307 ( .A(n32996), .B(n13788), .Z(n13790) );
  XOR U14308 ( .A(b[21]), .B(a[58]), .Z(n14069) );
  NANDN U14309 ( .A(n33271), .B(n14069), .Z(n13789) );
  AND U14310 ( .A(n13790), .B(n13789), .Z(n14035) );
  NANDN U14311 ( .A(n33866), .B(n13791), .Z(n13793) );
  XOR U14312 ( .A(b[23]), .B(a[56]), .Z(n14072) );
  NANDN U14313 ( .A(n33644), .B(n14072), .Z(n13792) );
  AND U14314 ( .A(n13793), .B(n13792), .Z(n14034) );
  NANDN U14315 ( .A(n32483), .B(n13794), .Z(n13796) );
  XOR U14316 ( .A(b[19]), .B(a[60]), .Z(n14075) );
  NANDN U14317 ( .A(n32823), .B(n14075), .Z(n13795) );
  NAND U14318 ( .A(n13796), .B(n13795), .Z(n14033) );
  XOR U14319 ( .A(n14034), .B(n14033), .Z(n14036) );
  XOR U14320 ( .A(n14035), .B(n14036), .Z(n13926) );
  NANDN U14321 ( .A(n34909), .B(n13797), .Z(n13799) );
  XOR U14322 ( .A(b[31]), .B(a[48]), .Z(n14078) );
  NANDN U14323 ( .A(n35145), .B(n14078), .Z(n13798) );
  AND U14324 ( .A(n13799), .B(n13798), .Z(n13915) );
  NANDN U14325 ( .A(n38247), .B(n13800), .Z(n13802) );
  XOR U14326 ( .A(b[61]), .B(a[18]), .Z(n14081) );
  NANDN U14327 ( .A(n38248), .B(n14081), .Z(n13801) );
  AND U14328 ( .A(n13802), .B(n13801), .Z(n13914) );
  AND U14329 ( .A(b[63]), .B(a[14]), .Z(n13913) );
  XOR U14330 ( .A(n13914), .B(n13913), .Z(n13916) );
  XNOR U14331 ( .A(n13915), .B(n13916), .Z(n13925) );
  XNOR U14332 ( .A(n13926), .B(n13925), .Z(n13927) );
  NANDN U14333 ( .A(n13804), .B(n13803), .Z(n13808) );
  OR U14334 ( .A(n13806), .B(n13805), .Z(n13807) );
  NAND U14335 ( .A(n13808), .B(n13807), .Z(n13928) );
  XNOR U14336 ( .A(n13927), .B(n13928), .Z(n14114) );
  NANDN U14337 ( .A(n34223), .B(n13809), .Z(n13811) );
  XOR U14338 ( .A(b[27]), .B(a[52]), .Z(n14090) );
  NANDN U14339 ( .A(n34458), .B(n14090), .Z(n13810) );
  AND U14340 ( .A(n13811), .B(n13810), .Z(n13987) );
  NANDN U14341 ( .A(n34634), .B(n13812), .Z(n13814) );
  XOR U14342 ( .A(b[29]), .B(a[50]), .Z(n14093) );
  NANDN U14343 ( .A(n34722), .B(n14093), .Z(n13813) );
  AND U14344 ( .A(n13814), .B(n13813), .Z(n13986) );
  NANDN U14345 ( .A(n31055), .B(n13815), .Z(n13817) );
  XOR U14346 ( .A(b[13]), .B(a[66]), .Z(n14096) );
  NANDN U14347 ( .A(n31293), .B(n14096), .Z(n13816) );
  NAND U14348 ( .A(n13817), .B(n13816), .Z(n13985) );
  XOR U14349 ( .A(n13986), .B(n13985), .Z(n13988) );
  XOR U14350 ( .A(n13987), .B(n13988), .Z(n14010) );
  NANDN U14351 ( .A(n28889), .B(n13818), .Z(n13820) );
  XOR U14352 ( .A(a[74]), .B(b[5]), .Z(n14099) );
  NANDN U14353 ( .A(n29138), .B(n14099), .Z(n13819) );
  AND U14354 ( .A(n13820), .B(n13819), .Z(n14029) );
  NANDN U14355 ( .A(n209), .B(n13821), .Z(n13823) );
  XOR U14356 ( .A(a[76]), .B(b[3]), .Z(n14102) );
  NANDN U14357 ( .A(n28941), .B(n14102), .Z(n13822) );
  AND U14358 ( .A(n13823), .B(n13822), .Z(n14028) );
  NANDN U14359 ( .A(n35936), .B(n13824), .Z(n13826) );
  XOR U14360 ( .A(b[37]), .B(a[42]), .Z(n14105) );
  NANDN U14361 ( .A(n36047), .B(n14105), .Z(n13825) );
  NAND U14362 ( .A(n13826), .B(n13825), .Z(n14027) );
  XOR U14363 ( .A(n14028), .B(n14027), .Z(n14030) );
  XNOR U14364 ( .A(n14029), .B(n14030), .Z(n14009) );
  XNOR U14365 ( .A(n14010), .B(n14009), .Z(n14011) );
  NANDN U14366 ( .A(n13828), .B(n13827), .Z(n13832) );
  OR U14367 ( .A(n13830), .B(n13829), .Z(n13831) );
  NAND U14368 ( .A(n13832), .B(n13831), .Z(n14012) );
  XOR U14369 ( .A(n14011), .B(n14012), .Z(n14115) );
  XNOR U14370 ( .A(n14114), .B(n14115), .Z(n14116) );
  XNOR U14371 ( .A(n14117), .B(n14116), .Z(n13900) );
  XOR U14372 ( .A(n13901), .B(n13900), .Z(n13893) );
  NANDN U14373 ( .A(n13834), .B(n13833), .Z(n13838) );
  NANDN U14374 ( .A(n13836), .B(n13835), .Z(n13837) );
  AND U14375 ( .A(n13838), .B(n13837), .Z(n13892) );
  XNOR U14376 ( .A(n13893), .B(n13892), .Z(n13894) );
  XOR U14377 ( .A(n13895), .B(n13894), .Z(n14121) );
  XNOR U14378 ( .A(n14120), .B(n14121), .Z(n14122) );
  XOR U14379 ( .A(n14123), .B(n14122), .Z(n14135) );
  XNOR U14380 ( .A(n14134), .B(n14135), .Z(n14140) );
  XOR U14381 ( .A(n14141), .B(n14140), .Z(n13863) );
  NANDN U14382 ( .A(n13840), .B(n13839), .Z(n13844) );
  NANDN U14383 ( .A(n13842), .B(n13841), .Z(n13843) );
  AND U14384 ( .A(n13844), .B(n13843), .Z(n13862) );
  XNOR U14385 ( .A(n13863), .B(n13862), .Z(n13864) );
  NANDN U14386 ( .A(n13846), .B(n13845), .Z(n13850) );
  NAND U14387 ( .A(n13848), .B(n13847), .Z(n13849) );
  NAND U14388 ( .A(n13850), .B(n13849), .Z(n13865) );
  XNOR U14389 ( .A(n13864), .B(n13865), .Z(n13856) );
  XNOR U14390 ( .A(n13857), .B(n13856), .Z(n13858) );
  XNOR U14391 ( .A(n13859), .B(n13858), .Z(n14144) );
  XNOR U14392 ( .A(sreg[142]), .B(n14144), .Z(n14146) );
  NANDN U14393 ( .A(sreg[141]), .B(n13851), .Z(n13855) );
  NAND U14394 ( .A(n13853), .B(n13852), .Z(n13854) );
  NAND U14395 ( .A(n13855), .B(n13854), .Z(n14145) );
  XNOR U14396 ( .A(n14146), .B(n14145), .Z(c[142]) );
  NANDN U14397 ( .A(n13857), .B(n13856), .Z(n13861) );
  NANDN U14398 ( .A(n13859), .B(n13858), .Z(n13860) );
  AND U14399 ( .A(n13861), .B(n13860), .Z(n14152) );
  NANDN U14400 ( .A(n13863), .B(n13862), .Z(n13867) );
  NANDN U14401 ( .A(n13865), .B(n13864), .Z(n13866) );
  AND U14402 ( .A(n13867), .B(n13866), .Z(n14150) );
  NANDN U14403 ( .A(n13869), .B(n13868), .Z(n13873) );
  OR U14404 ( .A(n13871), .B(n13870), .Z(n13872) );
  AND U14405 ( .A(n13873), .B(n13872), .Z(n14421) );
  NANDN U14406 ( .A(n13875), .B(n13874), .Z(n13879) );
  NAND U14407 ( .A(n13877), .B(n13876), .Z(n13878) );
  AND U14408 ( .A(n13879), .B(n13878), .Z(n14420) );
  NANDN U14409 ( .A(n13881), .B(n13880), .Z(n13885) );
  NANDN U14410 ( .A(n13883), .B(n13882), .Z(n13884) );
  AND U14411 ( .A(n13885), .B(n13884), .Z(n14419) );
  XOR U14412 ( .A(n14420), .B(n14419), .Z(n14422) );
  XOR U14413 ( .A(n14421), .B(n14422), .Z(n14426) );
  NANDN U14414 ( .A(n13887), .B(n13886), .Z(n13891) );
  NANDN U14415 ( .A(n13889), .B(n13888), .Z(n13890) );
  NAND U14416 ( .A(n13891), .B(n13890), .Z(n14425) );
  XNOR U14417 ( .A(n14426), .B(n14425), .Z(n14427) );
  NANDN U14418 ( .A(n13893), .B(n13892), .Z(n13897) );
  NANDN U14419 ( .A(n13895), .B(n13894), .Z(n13896) );
  AND U14420 ( .A(n13897), .B(n13896), .Z(n14416) );
  NANDN U14421 ( .A(n13899), .B(n13898), .Z(n13903) );
  NAND U14422 ( .A(n13901), .B(n13900), .Z(n13902) );
  AND U14423 ( .A(n13903), .B(n13902), .Z(n14163) );
  NANDN U14424 ( .A(n29499), .B(n13904), .Z(n13906) );
  XOR U14425 ( .A(b[7]), .B(a[73]), .Z(n14275) );
  NANDN U14426 ( .A(n29735), .B(n14275), .Z(n13905) );
  AND U14427 ( .A(n13906), .B(n13905), .Z(n14235) );
  NANDN U14428 ( .A(n37857), .B(n13907), .Z(n13909) );
  XOR U14429 ( .A(b[55]), .B(a[25]), .Z(n14278) );
  NANDN U14430 ( .A(n37911), .B(n14278), .Z(n13908) );
  AND U14431 ( .A(n13909), .B(n13908), .Z(n14234) );
  NANDN U14432 ( .A(n35611), .B(n13910), .Z(n13912) );
  XOR U14433 ( .A(b[35]), .B(a[45]), .Z(n14281) );
  NANDN U14434 ( .A(n35801), .B(n14281), .Z(n13911) );
  NAND U14435 ( .A(n13912), .B(n13911), .Z(n14233) );
  XOR U14436 ( .A(n14234), .B(n14233), .Z(n14236) );
  XOR U14437 ( .A(n14235), .B(n14236), .Z(n14297) );
  NANDN U14438 ( .A(n13914), .B(n13913), .Z(n13918) );
  OR U14439 ( .A(n13916), .B(n13915), .Z(n13917) );
  AND U14440 ( .A(n13918), .B(n13917), .Z(n14296) );
  XNOR U14441 ( .A(n14297), .B(n14296), .Z(n14298) );
  NANDN U14442 ( .A(n13920), .B(n13919), .Z(n13924) );
  OR U14443 ( .A(n13922), .B(n13921), .Z(n13923) );
  NAND U14444 ( .A(n13924), .B(n13923), .Z(n14299) );
  XNOR U14445 ( .A(n14298), .B(n14299), .Z(n14176) );
  NANDN U14446 ( .A(n13926), .B(n13925), .Z(n13930) );
  NANDN U14447 ( .A(n13928), .B(n13927), .Z(n13929) );
  AND U14448 ( .A(n13930), .B(n13929), .Z(n14174) );
  NAND U14449 ( .A(n37294), .B(n13931), .Z(n13933) );
  XNOR U14450 ( .A(b[47]), .B(a[33]), .Z(n14251) );
  NANDN U14451 ( .A(n14251), .B(n37341), .Z(n13932) );
  NAND U14452 ( .A(n13933), .B(n13932), .Z(n14292) );
  NAND U14453 ( .A(n30627), .B(n13934), .Z(n13936) );
  XNOR U14454 ( .A(b[9]), .B(a[71]), .Z(n14254) );
  NANDN U14455 ( .A(n14254), .B(n30628), .Z(n13935) );
  NAND U14456 ( .A(n13936), .B(n13935), .Z(n14291) );
  NAND U14457 ( .A(n37536), .B(n13937), .Z(n13939) );
  XNOR U14458 ( .A(b[49]), .B(a[31]), .Z(n14257) );
  NANDN U14459 ( .A(n14257), .B(n37537), .Z(n13938) );
  NAND U14460 ( .A(n13939), .B(n13938), .Z(n14290) );
  XNOR U14461 ( .A(n14291), .B(n14290), .Z(n14293) );
  NANDN U14462 ( .A(n36742), .B(n13940), .Z(n13942) );
  XOR U14463 ( .A(b[43]), .B(a[37]), .Z(n14260) );
  NANDN U14464 ( .A(n36891), .B(n14260), .Z(n13941) );
  AND U14465 ( .A(n13942), .B(n13941), .Z(n14271) );
  NANDN U14466 ( .A(n36991), .B(n13943), .Z(n13945) );
  XOR U14467 ( .A(b[45]), .B(a[35]), .Z(n14263) );
  NANDN U14468 ( .A(n37083), .B(n14263), .Z(n13944) );
  AND U14469 ( .A(n13945), .B(n13944), .Z(n14270) );
  NANDN U14470 ( .A(n30482), .B(n13946), .Z(n13948) );
  XOR U14471 ( .A(b[11]), .B(a[69]), .Z(n14266) );
  NANDN U14472 ( .A(n30891), .B(n14266), .Z(n13947) );
  NAND U14473 ( .A(n13948), .B(n13947), .Z(n14269) );
  XOR U14474 ( .A(n14270), .B(n14269), .Z(n14272) );
  XNOR U14475 ( .A(n14271), .B(n14272), .Z(n14356) );
  XOR U14476 ( .A(n14357), .B(n14356), .Z(n14358) );
  NANDN U14477 ( .A(n13950), .B(n13949), .Z(n13954) );
  OR U14478 ( .A(n13952), .B(n13951), .Z(n13953) );
  NAND U14479 ( .A(n13954), .B(n13953), .Z(n14359) );
  XNOR U14480 ( .A(n14358), .B(n14359), .Z(n14173) );
  XNOR U14481 ( .A(n14174), .B(n14173), .Z(n14175) );
  XOR U14482 ( .A(n14176), .B(n14175), .Z(n14162) );
  NANDN U14483 ( .A(n13956), .B(n13955), .Z(n13960) );
  NANDN U14484 ( .A(n13958), .B(n13957), .Z(n13959) );
  AND U14485 ( .A(n13960), .B(n13959), .Z(n14182) );
  NANDN U14486 ( .A(n13962), .B(n13961), .Z(n13966) );
  NANDN U14487 ( .A(n13964), .B(n13963), .Z(n13965) );
  AND U14488 ( .A(n13966), .B(n13965), .Z(n14180) );
  NANDN U14489 ( .A(n33875), .B(n13967), .Z(n13969) );
  XOR U14490 ( .A(b[25]), .B(a[55]), .Z(n14209) );
  NANDN U14491 ( .A(n33994), .B(n14209), .Z(n13968) );
  AND U14492 ( .A(n13969), .B(n13968), .Z(n14364) );
  NANDN U14493 ( .A(n32013), .B(n13970), .Z(n13972) );
  XOR U14494 ( .A(b[17]), .B(a[63]), .Z(n14212) );
  NANDN U14495 ( .A(n32292), .B(n14212), .Z(n13971) );
  AND U14496 ( .A(n13972), .B(n13971), .Z(n14363) );
  NANDN U14497 ( .A(n31536), .B(n13973), .Z(n13975) );
  XOR U14498 ( .A(b[15]), .B(a[65]), .Z(n14215) );
  NANDN U14499 ( .A(n31925), .B(n14215), .Z(n13974) );
  NAND U14500 ( .A(n13975), .B(n13974), .Z(n14362) );
  XOR U14501 ( .A(n14363), .B(n14362), .Z(n14365) );
  XOR U14502 ( .A(n14364), .B(n14365), .Z(n14351) );
  NANDN U14503 ( .A(n37526), .B(n13976), .Z(n13978) );
  XOR U14504 ( .A(b[51]), .B(a[29]), .Z(n14218) );
  NANDN U14505 ( .A(n37605), .B(n14218), .Z(n13977) );
  AND U14506 ( .A(n13978), .B(n13977), .Z(n14385) );
  NANDN U14507 ( .A(n37705), .B(n13979), .Z(n13981) );
  XOR U14508 ( .A(b[53]), .B(a[27]), .Z(n14221) );
  NANDN U14509 ( .A(n37778), .B(n14221), .Z(n13980) );
  AND U14510 ( .A(n13981), .B(n13980), .Z(n14384) );
  NANDN U14511 ( .A(n36210), .B(n13982), .Z(n13984) );
  XOR U14512 ( .A(b[39]), .B(a[41]), .Z(n14224) );
  NANDN U14513 ( .A(n36347), .B(n14224), .Z(n13983) );
  NAND U14514 ( .A(n13984), .B(n13983), .Z(n14383) );
  XOR U14515 ( .A(n14384), .B(n14383), .Z(n14386) );
  XNOR U14516 ( .A(n14385), .B(n14386), .Z(n14350) );
  XNOR U14517 ( .A(n14351), .B(n14350), .Z(n14353) );
  NANDN U14518 ( .A(n13986), .B(n13985), .Z(n13990) );
  OR U14519 ( .A(n13988), .B(n13987), .Z(n13989) );
  AND U14520 ( .A(n13990), .B(n13989), .Z(n14352) );
  XOR U14521 ( .A(n14353), .B(n14352), .Z(n14200) );
  NANDN U14522 ( .A(n13992), .B(n13991), .Z(n13996) );
  OR U14523 ( .A(n13994), .B(n13993), .Z(n13995) );
  AND U14524 ( .A(n13996), .B(n13995), .Z(n14198) );
  NANDN U14525 ( .A(n13998), .B(n13997), .Z(n14002) );
  NANDN U14526 ( .A(n14000), .B(n13999), .Z(n14001) );
  NAND U14527 ( .A(n14002), .B(n14001), .Z(n14197) );
  XNOR U14528 ( .A(n14198), .B(n14197), .Z(n14199) );
  XNOR U14529 ( .A(n14200), .B(n14199), .Z(n14179) );
  XNOR U14530 ( .A(n14180), .B(n14179), .Z(n14181) );
  XNOR U14531 ( .A(n14182), .B(n14181), .Z(n14161) );
  XOR U14532 ( .A(n14162), .B(n14161), .Z(n14164) );
  XNOR U14533 ( .A(n14163), .B(n14164), .Z(n14413) );
  NANDN U14534 ( .A(n14004), .B(n14003), .Z(n14008) );
  NANDN U14535 ( .A(n14006), .B(n14005), .Z(n14007) );
  AND U14536 ( .A(n14008), .B(n14007), .Z(n14169) );
  NANDN U14537 ( .A(n14010), .B(n14009), .Z(n14014) );
  NANDN U14538 ( .A(n14012), .B(n14011), .Z(n14013) );
  AND U14539 ( .A(n14014), .B(n14013), .Z(n14168) );
  NANDN U14540 ( .A(n14016), .B(n14015), .Z(n14020) );
  NAND U14541 ( .A(n14018), .B(n14017), .Z(n14019) );
  AND U14542 ( .A(n14020), .B(n14019), .Z(n14167) );
  XOR U14543 ( .A(n14168), .B(n14167), .Z(n14170) );
  XOR U14544 ( .A(n14169), .B(n14170), .Z(n14188) );
  NANDN U14545 ( .A(n14022), .B(n14021), .Z(n14026) );
  NANDN U14546 ( .A(n14024), .B(n14023), .Z(n14025) );
  AND U14547 ( .A(n14026), .B(n14025), .Z(n14309) );
  NANDN U14548 ( .A(n14028), .B(n14027), .Z(n14032) );
  OR U14549 ( .A(n14030), .B(n14029), .Z(n14031) );
  NAND U14550 ( .A(n14032), .B(n14031), .Z(n14308) );
  XNOR U14551 ( .A(n14309), .B(n14308), .Z(n14311) );
  NANDN U14552 ( .A(n14034), .B(n14033), .Z(n14038) );
  OR U14553 ( .A(n14036), .B(n14035), .Z(n14037) );
  AND U14554 ( .A(n14038), .B(n14037), .Z(n14206) );
  NANDN U14555 ( .A(n38278), .B(n14039), .Z(n14041) );
  XOR U14556 ( .A(b[63]), .B(a[17]), .Z(n14335) );
  NANDN U14557 ( .A(n38279), .B(n14335), .Z(n14040) );
  AND U14558 ( .A(n14041), .B(n14040), .Z(n14240) );
  NANDN U14559 ( .A(n35260), .B(n14042), .Z(n14044) );
  XOR U14560 ( .A(b[33]), .B(a[47]), .Z(n14338) );
  NANDN U14561 ( .A(n35456), .B(n14338), .Z(n14043) );
  NAND U14562 ( .A(n14044), .B(n14043), .Z(n14239) );
  XNOR U14563 ( .A(n14240), .B(n14239), .Z(n14241) );
  NAND U14564 ( .A(b[0]), .B(a[79]), .Z(n14045) );
  XNOR U14565 ( .A(b[1]), .B(n14045), .Z(n14047) );
  NANDN U14566 ( .A(b[0]), .B(a[78]), .Z(n14046) );
  NAND U14567 ( .A(n14047), .B(n14046), .Z(n14242) );
  XNOR U14568 ( .A(n14241), .B(n14242), .Z(n14203) );
  NANDN U14569 ( .A(n37974), .B(n14048), .Z(n14050) );
  XOR U14570 ( .A(b[57]), .B(a[23]), .Z(n14341) );
  NANDN U14571 ( .A(n38031), .B(n14341), .Z(n14049) );
  AND U14572 ( .A(n14050), .B(n14049), .Z(n14317) );
  NANDN U14573 ( .A(n38090), .B(n14051), .Z(n14053) );
  XOR U14574 ( .A(b[59]), .B(a[21]), .Z(n14344) );
  NANDN U14575 ( .A(n38130), .B(n14344), .Z(n14052) );
  AND U14576 ( .A(n14053), .B(n14052), .Z(n14315) );
  NANDN U14577 ( .A(n36480), .B(n14054), .Z(n14056) );
  XOR U14578 ( .A(b[41]), .B(a[39]), .Z(n14347) );
  NANDN U14579 ( .A(n36594), .B(n14347), .Z(n14055) );
  NAND U14580 ( .A(n14056), .B(n14055), .Z(n14314) );
  XNOR U14581 ( .A(n14315), .B(n14314), .Z(n14316) );
  XOR U14582 ( .A(n14317), .B(n14316), .Z(n14204) );
  XNOR U14583 ( .A(n14203), .B(n14204), .Z(n14205) );
  XNOR U14584 ( .A(n14206), .B(n14205), .Z(n14310) );
  XOR U14585 ( .A(n14311), .B(n14310), .Z(n14192) );
  NANDN U14586 ( .A(n14058), .B(n14057), .Z(n14062) );
  NAND U14587 ( .A(n14060), .B(n14059), .Z(n14061) );
  NAND U14588 ( .A(n14062), .B(n14061), .Z(n14191) );
  XNOR U14589 ( .A(n14192), .B(n14191), .Z(n14194) );
  NANDN U14590 ( .A(n14064), .B(n14063), .Z(n14068) );
  NANDN U14591 ( .A(n14066), .B(n14065), .Z(n14067) );
  AND U14592 ( .A(n14068), .B(n14067), .Z(n14410) );
  NANDN U14593 ( .A(n32996), .B(n14069), .Z(n14071) );
  XOR U14594 ( .A(b[21]), .B(a[59]), .Z(n14368) );
  NANDN U14595 ( .A(n33271), .B(n14368), .Z(n14070) );
  AND U14596 ( .A(n14071), .B(n14070), .Z(n14328) );
  NANDN U14597 ( .A(n33866), .B(n14072), .Z(n14074) );
  XOR U14598 ( .A(b[23]), .B(a[57]), .Z(n14371) );
  NANDN U14599 ( .A(n33644), .B(n14371), .Z(n14073) );
  AND U14600 ( .A(n14074), .B(n14073), .Z(n14327) );
  NANDN U14601 ( .A(n32483), .B(n14075), .Z(n14077) );
  XOR U14602 ( .A(b[19]), .B(a[61]), .Z(n14374) );
  NANDN U14603 ( .A(n32823), .B(n14374), .Z(n14076) );
  NAND U14604 ( .A(n14077), .B(n14076), .Z(n14326) );
  XOR U14605 ( .A(n14327), .B(n14326), .Z(n14329) );
  XOR U14606 ( .A(n14328), .B(n14329), .Z(n14246) );
  NANDN U14607 ( .A(n34909), .B(n14078), .Z(n14080) );
  XOR U14608 ( .A(b[31]), .B(a[49]), .Z(n14377) );
  NANDN U14609 ( .A(n35145), .B(n14377), .Z(n14079) );
  AND U14610 ( .A(n14080), .B(n14079), .Z(n14286) );
  NANDN U14611 ( .A(n38247), .B(n14081), .Z(n14083) );
  XOR U14612 ( .A(b[61]), .B(a[19]), .Z(n14380) );
  NANDN U14613 ( .A(n38248), .B(n14380), .Z(n14082) );
  AND U14614 ( .A(n14083), .B(n14082), .Z(n14285) );
  AND U14615 ( .A(b[63]), .B(a[15]), .Z(n14284) );
  XOR U14616 ( .A(n14285), .B(n14284), .Z(n14287) );
  XNOR U14617 ( .A(n14286), .B(n14287), .Z(n14245) );
  XNOR U14618 ( .A(n14246), .B(n14245), .Z(n14247) );
  NANDN U14619 ( .A(n14085), .B(n14084), .Z(n14089) );
  OR U14620 ( .A(n14087), .B(n14086), .Z(n14088) );
  NAND U14621 ( .A(n14089), .B(n14088), .Z(n14248) );
  XNOR U14622 ( .A(n14247), .B(n14248), .Z(n14407) );
  NANDN U14623 ( .A(n34223), .B(n14090), .Z(n14092) );
  XOR U14624 ( .A(b[27]), .B(a[53]), .Z(n14389) );
  NANDN U14625 ( .A(n34458), .B(n14389), .Z(n14091) );
  AND U14626 ( .A(n14092), .B(n14091), .Z(n14229) );
  NANDN U14627 ( .A(n34634), .B(n14093), .Z(n14095) );
  XOR U14628 ( .A(b[29]), .B(a[51]), .Z(n14392) );
  NANDN U14629 ( .A(n34722), .B(n14392), .Z(n14094) );
  AND U14630 ( .A(n14095), .B(n14094), .Z(n14228) );
  NANDN U14631 ( .A(n31055), .B(n14096), .Z(n14098) );
  XOR U14632 ( .A(b[13]), .B(a[67]), .Z(n14395) );
  NANDN U14633 ( .A(n31293), .B(n14395), .Z(n14097) );
  NAND U14634 ( .A(n14098), .B(n14097), .Z(n14227) );
  XOR U14635 ( .A(n14228), .B(n14227), .Z(n14230) );
  XOR U14636 ( .A(n14229), .B(n14230), .Z(n14303) );
  NANDN U14637 ( .A(n28889), .B(n14099), .Z(n14101) );
  XOR U14638 ( .A(a[75]), .B(b[5]), .Z(n14398) );
  NANDN U14639 ( .A(n29138), .B(n14398), .Z(n14100) );
  AND U14640 ( .A(n14101), .B(n14100), .Z(n14322) );
  NANDN U14641 ( .A(n209), .B(n14102), .Z(n14104) );
  XOR U14642 ( .A(a[77]), .B(b[3]), .Z(n14401) );
  NANDN U14643 ( .A(n28941), .B(n14401), .Z(n14103) );
  AND U14644 ( .A(n14104), .B(n14103), .Z(n14321) );
  NANDN U14645 ( .A(n35936), .B(n14105), .Z(n14107) );
  XOR U14646 ( .A(b[37]), .B(a[43]), .Z(n14404) );
  NANDN U14647 ( .A(n36047), .B(n14404), .Z(n14106) );
  NAND U14648 ( .A(n14107), .B(n14106), .Z(n14320) );
  XOR U14649 ( .A(n14321), .B(n14320), .Z(n14323) );
  XNOR U14650 ( .A(n14322), .B(n14323), .Z(n14302) );
  XNOR U14651 ( .A(n14303), .B(n14302), .Z(n14304) );
  NANDN U14652 ( .A(n14109), .B(n14108), .Z(n14113) );
  OR U14653 ( .A(n14111), .B(n14110), .Z(n14112) );
  NAND U14654 ( .A(n14113), .B(n14112), .Z(n14305) );
  XOR U14655 ( .A(n14304), .B(n14305), .Z(n14408) );
  XNOR U14656 ( .A(n14407), .B(n14408), .Z(n14409) );
  XNOR U14657 ( .A(n14410), .B(n14409), .Z(n14193) );
  XOR U14658 ( .A(n14194), .B(n14193), .Z(n14186) );
  NANDN U14659 ( .A(n14115), .B(n14114), .Z(n14119) );
  NANDN U14660 ( .A(n14117), .B(n14116), .Z(n14118) );
  AND U14661 ( .A(n14119), .B(n14118), .Z(n14185) );
  XNOR U14662 ( .A(n14186), .B(n14185), .Z(n14187) );
  XOR U14663 ( .A(n14188), .B(n14187), .Z(n14414) );
  XNOR U14664 ( .A(n14413), .B(n14414), .Z(n14415) );
  XOR U14665 ( .A(n14416), .B(n14415), .Z(n14428) );
  XNOR U14666 ( .A(n14427), .B(n14428), .Z(n14434) );
  NANDN U14667 ( .A(n14121), .B(n14120), .Z(n14125) );
  NANDN U14668 ( .A(n14123), .B(n14122), .Z(n14124) );
  AND U14669 ( .A(n14125), .B(n14124), .Z(n14432) );
  NANDN U14670 ( .A(n14127), .B(n14126), .Z(n14131) );
  OR U14671 ( .A(n14129), .B(n14128), .Z(n14130) );
  AND U14672 ( .A(n14131), .B(n14130), .Z(n14431) );
  XNOR U14673 ( .A(n14432), .B(n14431), .Z(n14433) );
  XOR U14674 ( .A(n14434), .B(n14433), .Z(n14156) );
  NANDN U14675 ( .A(n14133), .B(n14132), .Z(n14137) );
  NANDN U14676 ( .A(n14135), .B(n14134), .Z(n14136) );
  AND U14677 ( .A(n14137), .B(n14136), .Z(n14155) );
  XNOR U14678 ( .A(n14156), .B(n14155), .Z(n14157) );
  NANDN U14679 ( .A(n14139), .B(n14138), .Z(n14143) );
  NAND U14680 ( .A(n14141), .B(n14140), .Z(n14142) );
  NAND U14681 ( .A(n14143), .B(n14142), .Z(n14158) );
  XNOR U14682 ( .A(n14157), .B(n14158), .Z(n14149) );
  XNOR U14683 ( .A(n14150), .B(n14149), .Z(n14151) );
  XNOR U14684 ( .A(n14152), .B(n14151), .Z(n14437) );
  XNOR U14685 ( .A(sreg[143]), .B(n14437), .Z(n14439) );
  NANDN U14686 ( .A(sreg[142]), .B(n14144), .Z(n14148) );
  NAND U14687 ( .A(n14146), .B(n14145), .Z(n14147) );
  NAND U14688 ( .A(n14148), .B(n14147), .Z(n14438) );
  XNOR U14689 ( .A(n14439), .B(n14438), .Z(c[143]) );
  NANDN U14690 ( .A(n14150), .B(n14149), .Z(n14154) );
  NANDN U14691 ( .A(n14152), .B(n14151), .Z(n14153) );
  AND U14692 ( .A(n14154), .B(n14153), .Z(n14445) );
  NANDN U14693 ( .A(n14156), .B(n14155), .Z(n14160) );
  NANDN U14694 ( .A(n14158), .B(n14157), .Z(n14159) );
  AND U14695 ( .A(n14160), .B(n14159), .Z(n14443) );
  NANDN U14696 ( .A(n14162), .B(n14161), .Z(n14166) );
  NANDN U14697 ( .A(n14164), .B(n14163), .Z(n14165) );
  AND U14698 ( .A(n14166), .B(n14165), .Z(n14717) );
  NANDN U14699 ( .A(n14168), .B(n14167), .Z(n14172) );
  OR U14700 ( .A(n14170), .B(n14169), .Z(n14171) );
  AND U14701 ( .A(n14172), .B(n14171), .Z(n14712) );
  NANDN U14702 ( .A(n14174), .B(n14173), .Z(n14178) );
  NAND U14703 ( .A(n14176), .B(n14175), .Z(n14177) );
  AND U14704 ( .A(n14178), .B(n14177), .Z(n14711) );
  NANDN U14705 ( .A(n14180), .B(n14179), .Z(n14184) );
  NANDN U14706 ( .A(n14182), .B(n14181), .Z(n14183) );
  AND U14707 ( .A(n14184), .B(n14183), .Z(n14710) );
  XOR U14708 ( .A(n14711), .B(n14710), .Z(n14713) );
  XNOR U14709 ( .A(n14712), .B(n14713), .Z(n14716) );
  XNOR U14710 ( .A(n14717), .B(n14716), .Z(n14718) );
  NANDN U14711 ( .A(n14186), .B(n14185), .Z(n14190) );
  NANDN U14712 ( .A(n14188), .B(n14187), .Z(n14189) );
  AND U14713 ( .A(n14190), .B(n14189), .Z(n14707) );
  NANDN U14714 ( .A(n14192), .B(n14191), .Z(n14196) );
  NAND U14715 ( .A(n14194), .B(n14193), .Z(n14195) );
  AND U14716 ( .A(n14196), .B(n14195), .Z(n14682) );
  NANDN U14717 ( .A(n14198), .B(n14197), .Z(n14202) );
  NANDN U14718 ( .A(n14200), .B(n14199), .Z(n14201) );
  AND U14719 ( .A(n14202), .B(n14201), .Z(n14700) );
  NANDN U14720 ( .A(n14204), .B(n14203), .Z(n14208) );
  NANDN U14721 ( .A(n14206), .B(n14205), .Z(n14207) );
  AND U14722 ( .A(n14208), .B(n14207), .Z(n14699) );
  NANDN U14723 ( .A(n33875), .B(n14209), .Z(n14211) );
  XOR U14724 ( .A(b[25]), .B(a[56]), .Z(n14523) );
  NANDN U14725 ( .A(n33994), .B(n14523), .Z(n14210) );
  AND U14726 ( .A(n14211), .B(n14210), .Z(n14672) );
  NANDN U14727 ( .A(n32013), .B(n14212), .Z(n14214) );
  XOR U14728 ( .A(b[17]), .B(a[64]), .Z(n14526) );
  NANDN U14729 ( .A(n32292), .B(n14526), .Z(n14213) );
  AND U14730 ( .A(n14214), .B(n14213), .Z(n14671) );
  NANDN U14731 ( .A(n31536), .B(n14215), .Z(n14217) );
  XOR U14732 ( .A(b[15]), .B(a[66]), .Z(n14529) );
  NANDN U14733 ( .A(n31925), .B(n14529), .Z(n14216) );
  NAND U14734 ( .A(n14217), .B(n14216), .Z(n14670) );
  XOR U14735 ( .A(n14671), .B(n14670), .Z(n14673) );
  XOR U14736 ( .A(n14672), .B(n14673), .Z(n14620) );
  NANDN U14737 ( .A(n37526), .B(n14218), .Z(n14220) );
  XOR U14738 ( .A(b[51]), .B(a[30]), .Z(n14532) );
  NANDN U14739 ( .A(n37605), .B(n14532), .Z(n14219) );
  AND U14740 ( .A(n14220), .B(n14219), .Z(n14651) );
  NANDN U14741 ( .A(n37705), .B(n14221), .Z(n14223) );
  XOR U14742 ( .A(b[53]), .B(a[28]), .Z(n14535) );
  NANDN U14743 ( .A(n37778), .B(n14535), .Z(n14222) );
  AND U14744 ( .A(n14223), .B(n14222), .Z(n14650) );
  NANDN U14745 ( .A(n36210), .B(n14224), .Z(n14226) );
  XOR U14746 ( .A(b[39]), .B(a[42]), .Z(n14538) );
  NANDN U14747 ( .A(n36347), .B(n14538), .Z(n14225) );
  NAND U14748 ( .A(n14226), .B(n14225), .Z(n14649) );
  XOR U14749 ( .A(n14650), .B(n14649), .Z(n14652) );
  XNOR U14750 ( .A(n14651), .B(n14652), .Z(n14619) );
  XNOR U14751 ( .A(n14620), .B(n14619), .Z(n14622) );
  NANDN U14752 ( .A(n14228), .B(n14227), .Z(n14232) );
  OR U14753 ( .A(n14230), .B(n14229), .Z(n14231) );
  AND U14754 ( .A(n14232), .B(n14231), .Z(n14621) );
  XOR U14755 ( .A(n14622), .B(n14621), .Z(n14514) );
  NANDN U14756 ( .A(n14234), .B(n14233), .Z(n14238) );
  OR U14757 ( .A(n14236), .B(n14235), .Z(n14237) );
  AND U14758 ( .A(n14238), .B(n14237), .Z(n14512) );
  NANDN U14759 ( .A(n14240), .B(n14239), .Z(n14244) );
  NANDN U14760 ( .A(n14242), .B(n14241), .Z(n14243) );
  NAND U14761 ( .A(n14244), .B(n14243), .Z(n14511) );
  XNOR U14762 ( .A(n14512), .B(n14511), .Z(n14513) );
  XNOR U14763 ( .A(n14514), .B(n14513), .Z(n14698) );
  XOR U14764 ( .A(n14699), .B(n14698), .Z(n14701) );
  XOR U14765 ( .A(n14700), .B(n14701), .Z(n14681) );
  NANDN U14766 ( .A(n14246), .B(n14245), .Z(n14250) );
  NANDN U14767 ( .A(n14248), .B(n14247), .Z(n14249) );
  AND U14768 ( .A(n14250), .B(n14249), .Z(n14693) );
  NANDN U14769 ( .A(n14251), .B(n37294), .Z(n14253) );
  XOR U14770 ( .A(b[47]), .B(a[34]), .Z(n14466) );
  NANDN U14771 ( .A(n37172), .B(n14466), .Z(n14252) );
  AND U14772 ( .A(n14253), .B(n14252), .Z(n14507) );
  NANDN U14773 ( .A(n14254), .B(n30627), .Z(n14256) );
  XOR U14774 ( .A(b[9]), .B(a[72]), .Z(n14469) );
  NANDN U14775 ( .A(n30267), .B(n14469), .Z(n14255) );
  AND U14776 ( .A(n14256), .B(n14255), .Z(n14506) );
  NANDN U14777 ( .A(n14257), .B(n37536), .Z(n14259) );
  XOR U14778 ( .A(b[49]), .B(a[32]), .Z(n14472) );
  NANDN U14779 ( .A(n37432), .B(n14472), .Z(n14258) );
  NAND U14780 ( .A(n14259), .B(n14258), .Z(n14505) );
  XOR U14781 ( .A(n14506), .B(n14505), .Z(n14508) );
  XOR U14782 ( .A(n14507), .B(n14508), .Z(n14626) );
  NANDN U14783 ( .A(n36742), .B(n14260), .Z(n14262) );
  XOR U14784 ( .A(b[43]), .B(a[38]), .Z(n14475) );
  NANDN U14785 ( .A(n36891), .B(n14475), .Z(n14261) );
  AND U14786 ( .A(n14262), .B(n14261), .Z(n14486) );
  NANDN U14787 ( .A(n36991), .B(n14263), .Z(n14265) );
  XOR U14788 ( .A(b[45]), .B(a[36]), .Z(n14478) );
  NANDN U14789 ( .A(n37083), .B(n14478), .Z(n14264) );
  AND U14790 ( .A(n14265), .B(n14264), .Z(n14485) );
  NANDN U14791 ( .A(n30482), .B(n14266), .Z(n14268) );
  XOR U14792 ( .A(b[11]), .B(a[70]), .Z(n14481) );
  NANDN U14793 ( .A(n30891), .B(n14481), .Z(n14267) );
  NAND U14794 ( .A(n14268), .B(n14267), .Z(n14484) );
  XOR U14795 ( .A(n14485), .B(n14484), .Z(n14487) );
  XNOR U14796 ( .A(n14486), .B(n14487), .Z(n14625) );
  XNOR U14797 ( .A(n14626), .B(n14625), .Z(n14627) );
  NANDN U14798 ( .A(n14270), .B(n14269), .Z(n14274) );
  OR U14799 ( .A(n14272), .B(n14271), .Z(n14273) );
  NAND U14800 ( .A(n14274), .B(n14273), .Z(n14628) );
  XNOR U14801 ( .A(n14627), .B(n14628), .Z(n14692) );
  XNOR U14802 ( .A(n14693), .B(n14692), .Z(n14694) );
  NANDN U14803 ( .A(n29499), .B(n14275), .Z(n14277) );
  XOR U14804 ( .A(a[74]), .B(b[7]), .Z(n14490) );
  NANDN U14805 ( .A(n29735), .B(n14490), .Z(n14276) );
  AND U14806 ( .A(n14277), .B(n14276), .Z(n14549) );
  NANDN U14807 ( .A(n37857), .B(n14278), .Z(n14280) );
  XOR U14808 ( .A(b[55]), .B(a[26]), .Z(n14493) );
  NANDN U14809 ( .A(n37911), .B(n14493), .Z(n14279) );
  AND U14810 ( .A(n14280), .B(n14279), .Z(n14548) );
  NANDN U14811 ( .A(n35611), .B(n14281), .Z(n14283) );
  XOR U14812 ( .A(b[35]), .B(a[46]), .Z(n14496) );
  NANDN U14813 ( .A(n35801), .B(n14496), .Z(n14282) );
  NAND U14814 ( .A(n14283), .B(n14282), .Z(n14547) );
  XOR U14815 ( .A(n14548), .B(n14547), .Z(n14550) );
  XOR U14816 ( .A(n14549), .B(n14550), .Z(n14578) );
  NANDN U14817 ( .A(n14285), .B(n14284), .Z(n14289) );
  OR U14818 ( .A(n14287), .B(n14286), .Z(n14288) );
  AND U14819 ( .A(n14289), .B(n14288), .Z(n14577) );
  XNOR U14820 ( .A(n14578), .B(n14577), .Z(n14579) );
  NAND U14821 ( .A(n14291), .B(n14290), .Z(n14295) );
  NANDN U14822 ( .A(n14293), .B(n14292), .Z(n14294) );
  NAND U14823 ( .A(n14295), .B(n14294), .Z(n14580) );
  XOR U14824 ( .A(n14579), .B(n14580), .Z(n14695) );
  XNOR U14825 ( .A(n14694), .B(n14695), .Z(n14680) );
  XOR U14826 ( .A(n14681), .B(n14680), .Z(n14683) );
  XOR U14827 ( .A(n14682), .B(n14683), .Z(n14705) );
  NANDN U14828 ( .A(n14297), .B(n14296), .Z(n14301) );
  NANDN U14829 ( .A(n14299), .B(n14298), .Z(n14300) );
  AND U14830 ( .A(n14301), .B(n14300), .Z(n14688) );
  NANDN U14831 ( .A(n14303), .B(n14302), .Z(n14307) );
  NANDN U14832 ( .A(n14305), .B(n14304), .Z(n14306) );
  AND U14833 ( .A(n14307), .B(n14306), .Z(n14687) );
  NANDN U14834 ( .A(n14309), .B(n14308), .Z(n14313) );
  NAND U14835 ( .A(n14311), .B(n14310), .Z(n14312) );
  AND U14836 ( .A(n14313), .B(n14312), .Z(n14686) );
  XOR U14837 ( .A(n14687), .B(n14686), .Z(n14689) );
  XOR U14838 ( .A(n14688), .B(n14689), .Z(n14457) );
  NANDN U14839 ( .A(n14315), .B(n14314), .Z(n14319) );
  NANDN U14840 ( .A(n14317), .B(n14316), .Z(n14318) );
  AND U14841 ( .A(n14319), .B(n14318), .Z(n14572) );
  NANDN U14842 ( .A(n14321), .B(n14320), .Z(n14325) );
  OR U14843 ( .A(n14323), .B(n14322), .Z(n14324) );
  NAND U14844 ( .A(n14325), .B(n14324), .Z(n14571) );
  XNOR U14845 ( .A(n14572), .B(n14571), .Z(n14574) );
  NANDN U14846 ( .A(n14327), .B(n14326), .Z(n14331) );
  OR U14847 ( .A(n14329), .B(n14328), .Z(n14330) );
  NAND U14848 ( .A(n14331), .B(n14330), .Z(n14519) );
  NAND U14849 ( .A(b[0]), .B(a[80]), .Z(n14332) );
  XNOR U14850 ( .A(b[1]), .B(n14332), .Z(n14334) );
  NANDN U14851 ( .A(b[0]), .B(a[79]), .Z(n14333) );
  NAND U14852 ( .A(n14334), .B(n14333), .Z(n14556) );
  NANDN U14853 ( .A(n38278), .B(n14335), .Z(n14337) );
  XOR U14854 ( .A(b[63]), .B(a[18]), .Z(n14604) );
  NANDN U14855 ( .A(n38279), .B(n14604), .Z(n14336) );
  AND U14856 ( .A(n14337), .B(n14336), .Z(n14554) );
  NANDN U14857 ( .A(n35260), .B(n14338), .Z(n14340) );
  XOR U14858 ( .A(b[33]), .B(a[48]), .Z(n14607) );
  NANDN U14859 ( .A(n35456), .B(n14607), .Z(n14339) );
  NAND U14860 ( .A(n14340), .B(n14339), .Z(n14553) );
  XNOR U14861 ( .A(n14554), .B(n14553), .Z(n14555) );
  XNOR U14862 ( .A(n14556), .B(n14555), .Z(n14518) );
  NANDN U14863 ( .A(n37974), .B(n14341), .Z(n14343) );
  XOR U14864 ( .A(b[57]), .B(a[24]), .Z(n14610) );
  NANDN U14865 ( .A(n38031), .B(n14610), .Z(n14342) );
  AND U14866 ( .A(n14343), .B(n14342), .Z(n14585) );
  NANDN U14867 ( .A(n38090), .B(n14344), .Z(n14346) );
  XOR U14868 ( .A(b[59]), .B(a[22]), .Z(n14613) );
  NANDN U14869 ( .A(n38130), .B(n14613), .Z(n14345) );
  AND U14870 ( .A(n14346), .B(n14345), .Z(n14584) );
  NANDN U14871 ( .A(n36480), .B(n14347), .Z(n14349) );
  XOR U14872 ( .A(b[41]), .B(a[40]), .Z(n14616) );
  NANDN U14873 ( .A(n36594), .B(n14616), .Z(n14348) );
  NAND U14874 ( .A(n14349), .B(n14348), .Z(n14583) );
  XOR U14875 ( .A(n14584), .B(n14583), .Z(n14586) );
  XOR U14876 ( .A(n14585), .B(n14586), .Z(n14517) );
  XOR U14877 ( .A(n14518), .B(n14517), .Z(n14520) );
  XOR U14878 ( .A(n14519), .B(n14520), .Z(n14573) );
  XOR U14879 ( .A(n14574), .B(n14573), .Z(n14560) );
  NANDN U14880 ( .A(n14351), .B(n14350), .Z(n14355) );
  NAND U14881 ( .A(n14353), .B(n14352), .Z(n14354) );
  NAND U14882 ( .A(n14355), .B(n14354), .Z(n14559) );
  XNOR U14883 ( .A(n14560), .B(n14559), .Z(n14562) );
  NAND U14884 ( .A(n14357), .B(n14356), .Z(n14361) );
  NANDN U14885 ( .A(n14359), .B(n14358), .Z(n14360) );
  AND U14886 ( .A(n14361), .B(n14360), .Z(n14679) );
  NANDN U14887 ( .A(n14363), .B(n14362), .Z(n14367) );
  OR U14888 ( .A(n14365), .B(n14364), .Z(n14366) );
  AND U14889 ( .A(n14367), .B(n14366), .Z(n14462) );
  NANDN U14890 ( .A(n32996), .B(n14368), .Z(n14370) );
  XOR U14891 ( .A(b[21]), .B(a[60]), .Z(n14655) );
  NANDN U14892 ( .A(n33271), .B(n14655), .Z(n14369) );
  AND U14893 ( .A(n14370), .B(n14369), .Z(n14598) );
  NANDN U14894 ( .A(n33866), .B(n14371), .Z(n14373) );
  XOR U14895 ( .A(b[23]), .B(a[58]), .Z(n14658) );
  NANDN U14896 ( .A(n33644), .B(n14658), .Z(n14372) );
  AND U14897 ( .A(n14373), .B(n14372), .Z(n14596) );
  NANDN U14898 ( .A(n32483), .B(n14374), .Z(n14376) );
  XOR U14899 ( .A(b[19]), .B(a[62]), .Z(n14661) );
  NANDN U14900 ( .A(n32823), .B(n14661), .Z(n14375) );
  NAND U14901 ( .A(n14376), .B(n14375), .Z(n14595) );
  XNOR U14902 ( .A(n14596), .B(n14595), .Z(n14597) );
  XOR U14903 ( .A(n14598), .B(n14597), .Z(n14461) );
  NANDN U14904 ( .A(n34909), .B(n14377), .Z(n14379) );
  XOR U14905 ( .A(b[31]), .B(a[50]), .Z(n14664) );
  NANDN U14906 ( .A(n35145), .B(n14664), .Z(n14378) );
  AND U14907 ( .A(n14379), .B(n14378), .Z(n14502) );
  NANDN U14908 ( .A(n38247), .B(n14380), .Z(n14382) );
  XOR U14909 ( .A(b[61]), .B(a[20]), .Z(n14667) );
  NANDN U14910 ( .A(n38248), .B(n14667), .Z(n14381) );
  AND U14911 ( .A(n14382), .B(n14381), .Z(n14500) );
  AND U14912 ( .A(b[63]), .B(a[16]), .Z(n14499) );
  XNOR U14913 ( .A(n14500), .B(n14499), .Z(n14501) );
  XOR U14914 ( .A(n14502), .B(n14501), .Z(n14460) );
  XNOR U14915 ( .A(n14461), .B(n14460), .Z(n14463) );
  NANDN U14916 ( .A(n14384), .B(n14383), .Z(n14388) );
  OR U14917 ( .A(n14386), .B(n14385), .Z(n14387) );
  AND U14918 ( .A(n14388), .B(n14387), .Z(n14567) );
  NANDN U14919 ( .A(n34223), .B(n14389), .Z(n14391) );
  XOR U14920 ( .A(b[27]), .B(a[54]), .Z(n14631) );
  NANDN U14921 ( .A(n34458), .B(n14631), .Z(n14390) );
  AND U14922 ( .A(n14391), .B(n14390), .Z(n14544) );
  NANDN U14923 ( .A(n34634), .B(n14392), .Z(n14394) );
  XOR U14924 ( .A(b[29]), .B(a[52]), .Z(n14634) );
  NANDN U14925 ( .A(n34722), .B(n14634), .Z(n14393) );
  AND U14926 ( .A(n14394), .B(n14393), .Z(n14542) );
  NANDN U14927 ( .A(n31055), .B(n14395), .Z(n14397) );
  XOR U14928 ( .A(b[13]), .B(a[68]), .Z(n14637) );
  NANDN U14929 ( .A(n31293), .B(n14637), .Z(n14396) );
  NAND U14930 ( .A(n14397), .B(n14396), .Z(n14541) );
  XNOR U14931 ( .A(n14542), .B(n14541), .Z(n14543) );
  XOR U14932 ( .A(n14544), .B(n14543), .Z(n14566) );
  NANDN U14933 ( .A(n28889), .B(n14398), .Z(n14400) );
  XOR U14934 ( .A(a[76]), .B(b[5]), .Z(n14640) );
  NANDN U14935 ( .A(n29138), .B(n14640), .Z(n14399) );
  AND U14936 ( .A(n14400), .B(n14399), .Z(n14592) );
  NANDN U14937 ( .A(n209), .B(n14401), .Z(n14403) );
  XOR U14938 ( .A(a[78]), .B(b[3]), .Z(n14643) );
  NANDN U14939 ( .A(n28941), .B(n14643), .Z(n14402) );
  AND U14940 ( .A(n14403), .B(n14402), .Z(n14590) );
  NANDN U14941 ( .A(n35936), .B(n14404), .Z(n14406) );
  XOR U14942 ( .A(b[37]), .B(a[44]), .Z(n14646) );
  NANDN U14943 ( .A(n36047), .B(n14646), .Z(n14405) );
  NAND U14944 ( .A(n14406), .B(n14405), .Z(n14589) );
  XNOR U14945 ( .A(n14590), .B(n14589), .Z(n14591) );
  XOR U14946 ( .A(n14592), .B(n14591), .Z(n14565) );
  XNOR U14947 ( .A(n14566), .B(n14565), .Z(n14568) );
  XOR U14948 ( .A(n14677), .B(n14676), .Z(n14678) );
  XNOR U14949 ( .A(n14679), .B(n14678), .Z(n14561) );
  XOR U14950 ( .A(n14562), .B(n14561), .Z(n14455) );
  NANDN U14951 ( .A(n14408), .B(n14407), .Z(n14412) );
  NANDN U14952 ( .A(n14410), .B(n14409), .Z(n14411) );
  AND U14953 ( .A(n14412), .B(n14411), .Z(n14454) );
  XNOR U14954 ( .A(n14455), .B(n14454), .Z(n14456) );
  XNOR U14955 ( .A(n14457), .B(n14456), .Z(n14704) );
  XNOR U14956 ( .A(n14705), .B(n14704), .Z(n14706) );
  XOR U14957 ( .A(n14707), .B(n14706), .Z(n14719) );
  XNOR U14958 ( .A(n14718), .B(n14719), .Z(n14725) );
  NANDN U14959 ( .A(n14414), .B(n14413), .Z(n14418) );
  NANDN U14960 ( .A(n14416), .B(n14415), .Z(n14417) );
  AND U14961 ( .A(n14418), .B(n14417), .Z(n14723) );
  NANDN U14962 ( .A(n14420), .B(n14419), .Z(n14424) );
  OR U14963 ( .A(n14422), .B(n14421), .Z(n14423) );
  AND U14964 ( .A(n14424), .B(n14423), .Z(n14722) );
  XNOR U14965 ( .A(n14723), .B(n14722), .Z(n14724) );
  XOR U14966 ( .A(n14725), .B(n14724), .Z(n14449) );
  NANDN U14967 ( .A(n14426), .B(n14425), .Z(n14430) );
  NANDN U14968 ( .A(n14428), .B(n14427), .Z(n14429) );
  AND U14969 ( .A(n14430), .B(n14429), .Z(n14448) );
  XNOR U14970 ( .A(n14449), .B(n14448), .Z(n14450) );
  NANDN U14971 ( .A(n14432), .B(n14431), .Z(n14436) );
  NAND U14972 ( .A(n14434), .B(n14433), .Z(n14435) );
  NAND U14973 ( .A(n14436), .B(n14435), .Z(n14451) );
  XNOR U14974 ( .A(n14450), .B(n14451), .Z(n14442) );
  XNOR U14975 ( .A(n14443), .B(n14442), .Z(n14444) );
  XNOR U14976 ( .A(n14445), .B(n14444), .Z(n14728) );
  XNOR U14977 ( .A(sreg[144]), .B(n14728), .Z(n14730) );
  NANDN U14978 ( .A(sreg[143]), .B(n14437), .Z(n14441) );
  NAND U14979 ( .A(n14439), .B(n14438), .Z(n14440) );
  NAND U14980 ( .A(n14441), .B(n14440), .Z(n14729) );
  XNOR U14981 ( .A(n14730), .B(n14729), .Z(c[144]) );
  NANDN U14982 ( .A(n14443), .B(n14442), .Z(n14447) );
  NANDN U14983 ( .A(n14445), .B(n14444), .Z(n14446) );
  AND U14984 ( .A(n14447), .B(n14446), .Z(n14736) );
  NANDN U14985 ( .A(n14449), .B(n14448), .Z(n14453) );
  NANDN U14986 ( .A(n14451), .B(n14450), .Z(n14452) );
  AND U14987 ( .A(n14453), .B(n14452), .Z(n14734) );
  NANDN U14988 ( .A(n14455), .B(n14454), .Z(n14459) );
  NANDN U14989 ( .A(n14457), .B(n14456), .Z(n14458) );
  AND U14990 ( .A(n14459), .B(n14458), .Z(n14747) );
  NAND U14991 ( .A(n14461), .B(n14460), .Z(n14465) );
  NANDN U14992 ( .A(n14463), .B(n14462), .Z(n14464) );
  AND U14993 ( .A(n14465), .B(n14464), .Z(n14776) );
  NAND U14994 ( .A(n37294), .B(n14466), .Z(n14468) );
  XNOR U14995 ( .A(b[47]), .B(a[35]), .Z(n14847) );
  NANDN U14996 ( .A(n14847), .B(n37341), .Z(n14467) );
  NAND U14997 ( .A(n14468), .B(n14467), .Z(n14888) );
  NAND U14998 ( .A(n30627), .B(n14469), .Z(n14471) );
  XNOR U14999 ( .A(b[9]), .B(a[73]), .Z(n14850) );
  NANDN U15000 ( .A(n14850), .B(n30628), .Z(n14470) );
  NAND U15001 ( .A(n14471), .B(n14470), .Z(n14887) );
  NAND U15002 ( .A(n37536), .B(n14472), .Z(n14474) );
  XNOR U15003 ( .A(b[49]), .B(a[33]), .Z(n14853) );
  NANDN U15004 ( .A(n14853), .B(n37537), .Z(n14473) );
  NAND U15005 ( .A(n14474), .B(n14473), .Z(n14886) );
  XNOR U15006 ( .A(n14887), .B(n14886), .Z(n14889) );
  NANDN U15007 ( .A(n36742), .B(n14475), .Z(n14477) );
  XOR U15008 ( .A(b[43]), .B(a[39]), .Z(n14856) );
  NANDN U15009 ( .A(n36891), .B(n14856), .Z(n14476) );
  AND U15010 ( .A(n14477), .B(n14476), .Z(n14867) );
  NANDN U15011 ( .A(n36991), .B(n14478), .Z(n14480) );
  XOR U15012 ( .A(b[45]), .B(a[37]), .Z(n14859) );
  NANDN U15013 ( .A(n37083), .B(n14859), .Z(n14479) );
  AND U15014 ( .A(n14480), .B(n14479), .Z(n14866) );
  NANDN U15015 ( .A(n30482), .B(n14481), .Z(n14483) );
  XOR U15016 ( .A(b[11]), .B(a[71]), .Z(n14862) );
  NANDN U15017 ( .A(n30891), .B(n14862), .Z(n14482) );
  NAND U15018 ( .A(n14483), .B(n14482), .Z(n14865) );
  XOR U15019 ( .A(n14866), .B(n14865), .Z(n14868) );
  XNOR U15020 ( .A(n14867), .B(n14868), .Z(n14952) );
  XOR U15021 ( .A(n14953), .B(n14952), .Z(n14954) );
  NANDN U15022 ( .A(n14485), .B(n14484), .Z(n14489) );
  OR U15023 ( .A(n14487), .B(n14486), .Z(n14488) );
  NAND U15024 ( .A(n14489), .B(n14488), .Z(n14955) );
  XNOR U15025 ( .A(n14954), .B(n14955), .Z(n14775) );
  XNOR U15026 ( .A(n14776), .B(n14775), .Z(n14778) );
  NANDN U15027 ( .A(n29499), .B(n14490), .Z(n14492) );
  XOR U15028 ( .A(a[75]), .B(b[7]), .Z(n14871) );
  NANDN U15029 ( .A(n29735), .B(n14871), .Z(n14491) );
  AND U15030 ( .A(n14492), .B(n14491), .Z(n14831) );
  NANDN U15031 ( .A(n37857), .B(n14493), .Z(n14495) );
  XOR U15032 ( .A(b[55]), .B(a[27]), .Z(n14874) );
  NANDN U15033 ( .A(n37911), .B(n14874), .Z(n14494) );
  AND U15034 ( .A(n14495), .B(n14494), .Z(n14830) );
  NANDN U15035 ( .A(n35611), .B(n14496), .Z(n14498) );
  XOR U15036 ( .A(b[35]), .B(a[47]), .Z(n14877) );
  NANDN U15037 ( .A(n35801), .B(n14877), .Z(n14497) );
  NAND U15038 ( .A(n14498), .B(n14497), .Z(n14829) );
  XOR U15039 ( .A(n14830), .B(n14829), .Z(n14832) );
  XOR U15040 ( .A(n14831), .B(n14832), .Z(n14893) );
  NANDN U15041 ( .A(n14500), .B(n14499), .Z(n14504) );
  NANDN U15042 ( .A(n14502), .B(n14501), .Z(n14503) );
  AND U15043 ( .A(n14504), .B(n14503), .Z(n14892) );
  XNOR U15044 ( .A(n14893), .B(n14892), .Z(n14894) );
  NANDN U15045 ( .A(n14506), .B(n14505), .Z(n14510) );
  OR U15046 ( .A(n14508), .B(n14507), .Z(n14509) );
  NAND U15047 ( .A(n14510), .B(n14509), .Z(n14895) );
  XNOR U15048 ( .A(n14894), .B(n14895), .Z(n14777) );
  XOR U15049 ( .A(n14778), .B(n14777), .Z(n14758) );
  NANDN U15050 ( .A(n14512), .B(n14511), .Z(n14516) );
  NANDN U15051 ( .A(n14514), .B(n14513), .Z(n14515) );
  AND U15052 ( .A(n14516), .B(n14515), .Z(n14772) );
  NAND U15053 ( .A(n14518), .B(n14517), .Z(n14522) );
  NAND U15054 ( .A(n14520), .B(n14519), .Z(n14521) );
  AND U15055 ( .A(n14522), .B(n14521), .Z(n14770) );
  NANDN U15056 ( .A(n33875), .B(n14523), .Z(n14525) );
  XOR U15057 ( .A(b[25]), .B(a[57]), .Z(n14805) );
  NANDN U15058 ( .A(n33994), .B(n14805), .Z(n14524) );
  AND U15059 ( .A(n14525), .B(n14524), .Z(n14960) );
  NANDN U15060 ( .A(n32013), .B(n14526), .Z(n14528) );
  XOR U15061 ( .A(b[17]), .B(a[65]), .Z(n14808) );
  NANDN U15062 ( .A(n32292), .B(n14808), .Z(n14527) );
  AND U15063 ( .A(n14528), .B(n14527), .Z(n14959) );
  NANDN U15064 ( .A(n31536), .B(n14529), .Z(n14531) );
  XOR U15065 ( .A(b[15]), .B(a[67]), .Z(n14811) );
  NANDN U15066 ( .A(n31925), .B(n14811), .Z(n14530) );
  NAND U15067 ( .A(n14531), .B(n14530), .Z(n14958) );
  XOR U15068 ( .A(n14959), .B(n14958), .Z(n14961) );
  XOR U15069 ( .A(n14960), .B(n14961), .Z(n14947) );
  NANDN U15070 ( .A(n37526), .B(n14532), .Z(n14534) );
  XOR U15071 ( .A(b[51]), .B(a[31]), .Z(n14814) );
  NANDN U15072 ( .A(n37605), .B(n14814), .Z(n14533) );
  AND U15073 ( .A(n14534), .B(n14533), .Z(n14981) );
  NANDN U15074 ( .A(n37705), .B(n14535), .Z(n14537) );
  XOR U15075 ( .A(b[53]), .B(a[29]), .Z(n14817) );
  NANDN U15076 ( .A(n37778), .B(n14817), .Z(n14536) );
  AND U15077 ( .A(n14537), .B(n14536), .Z(n14980) );
  NANDN U15078 ( .A(n36210), .B(n14538), .Z(n14540) );
  XOR U15079 ( .A(b[39]), .B(a[43]), .Z(n14820) );
  NANDN U15080 ( .A(n36347), .B(n14820), .Z(n14539) );
  NAND U15081 ( .A(n14540), .B(n14539), .Z(n14979) );
  XOR U15082 ( .A(n14980), .B(n14979), .Z(n14982) );
  XNOR U15083 ( .A(n14981), .B(n14982), .Z(n14946) );
  XNOR U15084 ( .A(n14947), .B(n14946), .Z(n14949) );
  NANDN U15085 ( .A(n14542), .B(n14541), .Z(n14546) );
  NANDN U15086 ( .A(n14544), .B(n14543), .Z(n14545) );
  AND U15087 ( .A(n14546), .B(n14545), .Z(n14948) );
  XOR U15088 ( .A(n14949), .B(n14948), .Z(n14796) );
  NANDN U15089 ( .A(n14548), .B(n14547), .Z(n14552) );
  OR U15090 ( .A(n14550), .B(n14549), .Z(n14551) );
  AND U15091 ( .A(n14552), .B(n14551), .Z(n14794) );
  NANDN U15092 ( .A(n14554), .B(n14553), .Z(n14558) );
  NANDN U15093 ( .A(n14556), .B(n14555), .Z(n14557) );
  NAND U15094 ( .A(n14558), .B(n14557), .Z(n14793) );
  XNOR U15095 ( .A(n14794), .B(n14793), .Z(n14795) );
  XNOR U15096 ( .A(n14796), .B(n14795), .Z(n14769) );
  XNOR U15097 ( .A(n14770), .B(n14769), .Z(n14771) );
  XNOR U15098 ( .A(n14772), .B(n14771), .Z(n14757) );
  XNOR U15099 ( .A(n14758), .B(n14757), .Z(n14759) );
  NANDN U15100 ( .A(n14560), .B(n14559), .Z(n14564) );
  NAND U15101 ( .A(n14562), .B(n14561), .Z(n14563) );
  NAND U15102 ( .A(n14564), .B(n14563), .Z(n14760) );
  XNOR U15103 ( .A(n14759), .B(n14760), .Z(n14745) );
  NAND U15104 ( .A(n14566), .B(n14565), .Z(n14570) );
  NANDN U15105 ( .A(n14568), .B(n14567), .Z(n14569) );
  NAND U15106 ( .A(n14570), .B(n14569), .Z(n14763) );
  NANDN U15107 ( .A(n14572), .B(n14571), .Z(n14576) );
  NAND U15108 ( .A(n14574), .B(n14573), .Z(n14575) );
  AND U15109 ( .A(n14576), .B(n14575), .Z(n14764) );
  XOR U15110 ( .A(n14763), .B(n14764), .Z(n14766) );
  NANDN U15111 ( .A(n14578), .B(n14577), .Z(n14582) );
  NANDN U15112 ( .A(n14580), .B(n14579), .Z(n14581) );
  NAND U15113 ( .A(n14582), .B(n14581), .Z(n14765) );
  XOR U15114 ( .A(n14766), .B(n14765), .Z(n14784) );
  NANDN U15115 ( .A(n14584), .B(n14583), .Z(n14588) );
  OR U15116 ( .A(n14586), .B(n14585), .Z(n14587) );
  AND U15117 ( .A(n14588), .B(n14587), .Z(n14905) );
  NANDN U15118 ( .A(n14590), .B(n14589), .Z(n14594) );
  NANDN U15119 ( .A(n14592), .B(n14591), .Z(n14593) );
  NAND U15120 ( .A(n14594), .B(n14593), .Z(n14904) );
  XNOR U15121 ( .A(n14905), .B(n14904), .Z(n14907) );
  NANDN U15122 ( .A(n14596), .B(n14595), .Z(n14600) );
  NANDN U15123 ( .A(n14598), .B(n14597), .Z(n14599) );
  AND U15124 ( .A(n14600), .B(n14599), .Z(n14802) );
  NAND U15125 ( .A(b[0]), .B(a[81]), .Z(n14601) );
  XNOR U15126 ( .A(b[1]), .B(n14601), .Z(n14603) );
  NANDN U15127 ( .A(b[0]), .B(a[80]), .Z(n14602) );
  NAND U15128 ( .A(n14603), .B(n14602), .Z(n14838) );
  NANDN U15129 ( .A(n38278), .B(n14604), .Z(n14606) );
  XOR U15130 ( .A(b[63]), .B(a[19]), .Z(n14931) );
  NANDN U15131 ( .A(n38279), .B(n14931), .Z(n14605) );
  AND U15132 ( .A(n14606), .B(n14605), .Z(n14836) );
  NANDN U15133 ( .A(n35260), .B(n14607), .Z(n14609) );
  XOR U15134 ( .A(b[33]), .B(a[49]), .Z(n14934) );
  NANDN U15135 ( .A(n35456), .B(n14934), .Z(n14608) );
  NAND U15136 ( .A(n14609), .B(n14608), .Z(n14835) );
  XNOR U15137 ( .A(n14836), .B(n14835), .Z(n14837) );
  XNOR U15138 ( .A(n14838), .B(n14837), .Z(n14799) );
  NANDN U15139 ( .A(n37974), .B(n14610), .Z(n14612) );
  XOR U15140 ( .A(b[57]), .B(a[25]), .Z(n14937) );
  NANDN U15141 ( .A(n38031), .B(n14937), .Z(n14611) );
  AND U15142 ( .A(n14612), .B(n14611), .Z(n14913) );
  NANDN U15143 ( .A(n38090), .B(n14613), .Z(n14615) );
  XOR U15144 ( .A(b[59]), .B(a[23]), .Z(n14940) );
  NANDN U15145 ( .A(n38130), .B(n14940), .Z(n14614) );
  AND U15146 ( .A(n14615), .B(n14614), .Z(n14911) );
  NANDN U15147 ( .A(n36480), .B(n14616), .Z(n14618) );
  XOR U15148 ( .A(b[41]), .B(a[41]), .Z(n14943) );
  NANDN U15149 ( .A(n36594), .B(n14943), .Z(n14617) );
  NAND U15150 ( .A(n14618), .B(n14617), .Z(n14910) );
  XNOR U15151 ( .A(n14911), .B(n14910), .Z(n14912) );
  XOR U15152 ( .A(n14913), .B(n14912), .Z(n14800) );
  XNOR U15153 ( .A(n14799), .B(n14800), .Z(n14801) );
  XNOR U15154 ( .A(n14802), .B(n14801), .Z(n14906) );
  XOR U15155 ( .A(n14907), .B(n14906), .Z(n14788) );
  NANDN U15156 ( .A(n14620), .B(n14619), .Z(n14624) );
  NAND U15157 ( .A(n14622), .B(n14621), .Z(n14623) );
  NAND U15158 ( .A(n14624), .B(n14623), .Z(n14787) );
  XNOR U15159 ( .A(n14788), .B(n14787), .Z(n14790) );
  NANDN U15160 ( .A(n14626), .B(n14625), .Z(n14630) );
  NANDN U15161 ( .A(n14628), .B(n14627), .Z(n14629) );
  AND U15162 ( .A(n14630), .B(n14629), .Z(n15006) );
  NANDN U15163 ( .A(n34223), .B(n14631), .Z(n14633) );
  XOR U15164 ( .A(b[27]), .B(a[55]), .Z(n14985) );
  NANDN U15165 ( .A(n34458), .B(n14985), .Z(n14632) );
  AND U15166 ( .A(n14633), .B(n14632), .Z(n14825) );
  NANDN U15167 ( .A(n34634), .B(n14634), .Z(n14636) );
  XOR U15168 ( .A(b[29]), .B(a[53]), .Z(n14988) );
  NANDN U15169 ( .A(n34722), .B(n14988), .Z(n14635) );
  AND U15170 ( .A(n14636), .B(n14635), .Z(n14824) );
  NANDN U15171 ( .A(n31055), .B(n14637), .Z(n14639) );
  XOR U15172 ( .A(b[13]), .B(a[69]), .Z(n14991) );
  NANDN U15173 ( .A(n31293), .B(n14991), .Z(n14638) );
  NAND U15174 ( .A(n14639), .B(n14638), .Z(n14823) );
  XOR U15175 ( .A(n14824), .B(n14823), .Z(n14826) );
  XOR U15176 ( .A(n14825), .B(n14826), .Z(n14899) );
  NANDN U15177 ( .A(n28889), .B(n14640), .Z(n14642) );
  XOR U15178 ( .A(a[77]), .B(b[5]), .Z(n14994) );
  NANDN U15179 ( .A(n29138), .B(n14994), .Z(n14641) );
  AND U15180 ( .A(n14642), .B(n14641), .Z(n14918) );
  NANDN U15181 ( .A(n209), .B(n14643), .Z(n14645) );
  XOR U15182 ( .A(a[79]), .B(b[3]), .Z(n14997) );
  NANDN U15183 ( .A(n28941), .B(n14997), .Z(n14644) );
  AND U15184 ( .A(n14645), .B(n14644), .Z(n14917) );
  NANDN U15185 ( .A(n35936), .B(n14646), .Z(n14648) );
  XOR U15186 ( .A(b[37]), .B(a[45]), .Z(n15000) );
  NANDN U15187 ( .A(n36047), .B(n15000), .Z(n14647) );
  NAND U15188 ( .A(n14648), .B(n14647), .Z(n14916) );
  XOR U15189 ( .A(n14917), .B(n14916), .Z(n14919) );
  XNOR U15190 ( .A(n14918), .B(n14919), .Z(n14898) );
  XNOR U15191 ( .A(n14899), .B(n14898), .Z(n14900) );
  NANDN U15192 ( .A(n14650), .B(n14649), .Z(n14654) );
  OR U15193 ( .A(n14652), .B(n14651), .Z(n14653) );
  NAND U15194 ( .A(n14654), .B(n14653), .Z(n14901) );
  XNOR U15195 ( .A(n14900), .B(n14901), .Z(n15003) );
  NANDN U15196 ( .A(n32996), .B(n14655), .Z(n14657) );
  XOR U15197 ( .A(b[21]), .B(a[61]), .Z(n14964) );
  NANDN U15198 ( .A(n33271), .B(n14964), .Z(n14656) );
  AND U15199 ( .A(n14657), .B(n14656), .Z(n14924) );
  NANDN U15200 ( .A(n33866), .B(n14658), .Z(n14660) );
  XOR U15201 ( .A(b[23]), .B(a[59]), .Z(n14967) );
  NANDN U15202 ( .A(n33644), .B(n14967), .Z(n14659) );
  AND U15203 ( .A(n14660), .B(n14659), .Z(n14923) );
  NANDN U15204 ( .A(n32483), .B(n14661), .Z(n14663) );
  XOR U15205 ( .A(b[19]), .B(a[63]), .Z(n14970) );
  NANDN U15206 ( .A(n32823), .B(n14970), .Z(n14662) );
  NAND U15207 ( .A(n14663), .B(n14662), .Z(n14922) );
  XOR U15208 ( .A(n14923), .B(n14922), .Z(n14925) );
  XOR U15209 ( .A(n14924), .B(n14925), .Z(n14842) );
  NANDN U15210 ( .A(n34909), .B(n14664), .Z(n14666) );
  XOR U15211 ( .A(b[31]), .B(a[51]), .Z(n14973) );
  NANDN U15212 ( .A(n35145), .B(n14973), .Z(n14665) );
  AND U15213 ( .A(n14666), .B(n14665), .Z(n14882) );
  NANDN U15214 ( .A(n38247), .B(n14667), .Z(n14669) );
  XOR U15215 ( .A(b[61]), .B(a[21]), .Z(n14976) );
  NANDN U15216 ( .A(n38248), .B(n14976), .Z(n14668) );
  AND U15217 ( .A(n14669), .B(n14668), .Z(n14881) );
  AND U15218 ( .A(b[63]), .B(a[17]), .Z(n14880) );
  XOR U15219 ( .A(n14881), .B(n14880), .Z(n14883) );
  XNOR U15220 ( .A(n14882), .B(n14883), .Z(n14841) );
  XNOR U15221 ( .A(n14842), .B(n14841), .Z(n14843) );
  NANDN U15222 ( .A(n14671), .B(n14670), .Z(n14675) );
  OR U15223 ( .A(n14673), .B(n14672), .Z(n14674) );
  NAND U15224 ( .A(n14675), .B(n14674), .Z(n14844) );
  XOR U15225 ( .A(n14843), .B(n14844), .Z(n15004) );
  XNOR U15226 ( .A(n15003), .B(n15004), .Z(n15005) );
  XNOR U15227 ( .A(n15006), .B(n15005), .Z(n14789) );
  XOR U15228 ( .A(n14790), .B(n14789), .Z(n14782) );
  XNOR U15229 ( .A(n14782), .B(n14781), .Z(n14783) );
  XOR U15230 ( .A(n14784), .B(n14783), .Z(n14746) );
  XOR U15231 ( .A(n14745), .B(n14746), .Z(n14748) );
  XOR U15232 ( .A(n14747), .B(n14748), .Z(n15011) );
  NANDN U15233 ( .A(n14681), .B(n14680), .Z(n14685) );
  OR U15234 ( .A(n14683), .B(n14682), .Z(n14684) );
  AND U15235 ( .A(n14685), .B(n14684), .Z(n15010) );
  NANDN U15236 ( .A(n14687), .B(n14686), .Z(n14691) );
  OR U15237 ( .A(n14689), .B(n14688), .Z(n14690) );
  AND U15238 ( .A(n14691), .B(n14690), .Z(n14754) );
  NANDN U15239 ( .A(n14693), .B(n14692), .Z(n14697) );
  NANDN U15240 ( .A(n14695), .B(n14694), .Z(n14696) );
  AND U15241 ( .A(n14697), .B(n14696), .Z(n14752) );
  NANDN U15242 ( .A(n14699), .B(n14698), .Z(n14703) );
  OR U15243 ( .A(n14701), .B(n14700), .Z(n14702) );
  AND U15244 ( .A(n14703), .B(n14702), .Z(n14751) );
  XNOR U15245 ( .A(n14752), .B(n14751), .Z(n14753) );
  XNOR U15246 ( .A(n14754), .B(n14753), .Z(n15009) );
  XOR U15247 ( .A(n15010), .B(n15009), .Z(n15012) );
  XOR U15248 ( .A(n15011), .B(n15012), .Z(n15017) );
  NANDN U15249 ( .A(n14705), .B(n14704), .Z(n14709) );
  NANDN U15250 ( .A(n14707), .B(n14706), .Z(n14708) );
  AND U15251 ( .A(n14709), .B(n14708), .Z(n15016) );
  NANDN U15252 ( .A(n14711), .B(n14710), .Z(n14715) );
  OR U15253 ( .A(n14713), .B(n14712), .Z(n14714) );
  AND U15254 ( .A(n14715), .B(n14714), .Z(n15015) );
  XOR U15255 ( .A(n15016), .B(n15015), .Z(n15018) );
  XOR U15256 ( .A(n15017), .B(n15018), .Z(n14740) );
  NANDN U15257 ( .A(n14717), .B(n14716), .Z(n14721) );
  NANDN U15258 ( .A(n14719), .B(n14718), .Z(n14720) );
  AND U15259 ( .A(n14721), .B(n14720), .Z(n14739) );
  XNOR U15260 ( .A(n14740), .B(n14739), .Z(n14741) );
  NANDN U15261 ( .A(n14723), .B(n14722), .Z(n14727) );
  NAND U15262 ( .A(n14725), .B(n14724), .Z(n14726) );
  NAND U15263 ( .A(n14727), .B(n14726), .Z(n14742) );
  XNOR U15264 ( .A(n14741), .B(n14742), .Z(n14733) );
  XNOR U15265 ( .A(n14734), .B(n14733), .Z(n14735) );
  XNOR U15266 ( .A(n14736), .B(n14735), .Z(n15021) );
  XNOR U15267 ( .A(sreg[145]), .B(n15021), .Z(n15023) );
  NANDN U15268 ( .A(sreg[144]), .B(n14728), .Z(n14732) );
  NAND U15269 ( .A(n14730), .B(n14729), .Z(n14731) );
  NAND U15270 ( .A(n14732), .B(n14731), .Z(n15022) );
  XNOR U15271 ( .A(n15023), .B(n15022), .Z(c[145]) );
  NANDN U15272 ( .A(n14734), .B(n14733), .Z(n14738) );
  NANDN U15273 ( .A(n14736), .B(n14735), .Z(n14737) );
  AND U15274 ( .A(n14738), .B(n14737), .Z(n15033) );
  NANDN U15275 ( .A(n14740), .B(n14739), .Z(n14744) );
  NANDN U15276 ( .A(n14742), .B(n14741), .Z(n14743) );
  AND U15277 ( .A(n14744), .B(n14743), .Z(n15032) );
  NANDN U15278 ( .A(n14746), .B(n14745), .Z(n14750) );
  OR U15279 ( .A(n14748), .B(n14747), .Z(n14749) );
  AND U15280 ( .A(n14750), .B(n14749), .Z(n15038) );
  NANDN U15281 ( .A(n14752), .B(n14751), .Z(n14756) );
  NANDN U15282 ( .A(n14754), .B(n14753), .Z(n14755) );
  AND U15283 ( .A(n14756), .B(n14755), .Z(n15037) );
  XNOR U15284 ( .A(n15038), .B(n15037), .Z(n15040) );
  NANDN U15285 ( .A(n14758), .B(n14757), .Z(n14762) );
  NANDN U15286 ( .A(n14760), .B(n14759), .Z(n14761) );
  AND U15287 ( .A(n14762), .B(n14761), .Z(n15044) );
  NAND U15288 ( .A(n14764), .B(n14763), .Z(n14768) );
  NAND U15289 ( .A(n14766), .B(n14765), .Z(n14767) );
  AND U15290 ( .A(n14768), .B(n14767), .Z(n15307) );
  NANDN U15291 ( .A(n14770), .B(n14769), .Z(n14774) );
  NANDN U15292 ( .A(n14772), .B(n14771), .Z(n14773) );
  AND U15293 ( .A(n14774), .B(n14773), .Z(n15306) );
  NANDN U15294 ( .A(n14776), .B(n14775), .Z(n14780) );
  NAND U15295 ( .A(n14778), .B(n14777), .Z(n14779) );
  AND U15296 ( .A(n14780), .B(n14779), .Z(n15305) );
  XOR U15297 ( .A(n15306), .B(n15305), .Z(n15308) );
  XNOR U15298 ( .A(n15307), .B(n15308), .Z(n15043) );
  XNOR U15299 ( .A(n15044), .B(n15043), .Z(n15045) );
  NANDN U15300 ( .A(n14782), .B(n14781), .Z(n14786) );
  NANDN U15301 ( .A(n14784), .B(n14783), .Z(n14785) );
  AND U15302 ( .A(n14786), .B(n14785), .Z(n15302) );
  NANDN U15303 ( .A(n14788), .B(n14787), .Z(n14792) );
  NAND U15304 ( .A(n14790), .B(n14789), .Z(n14791) );
  AND U15305 ( .A(n14792), .B(n14791), .Z(n15277) );
  NANDN U15306 ( .A(n14794), .B(n14793), .Z(n14798) );
  NANDN U15307 ( .A(n14796), .B(n14795), .Z(n14797) );
  AND U15308 ( .A(n14798), .B(n14797), .Z(n15295) );
  NANDN U15309 ( .A(n14800), .B(n14799), .Z(n14804) );
  NANDN U15310 ( .A(n14802), .B(n14801), .Z(n14803) );
  AND U15311 ( .A(n14804), .B(n14803), .Z(n15294) );
  NANDN U15312 ( .A(n33875), .B(n14805), .Z(n14807) );
  XOR U15313 ( .A(b[25]), .B(a[58]), .Z(n15073) );
  NANDN U15314 ( .A(n33994), .B(n15073), .Z(n14806) );
  AND U15315 ( .A(n14807), .B(n14806), .Z(n15243) );
  NANDN U15316 ( .A(n32013), .B(n14808), .Z(n14810) );
  XOR U15317 ( .A(b[17]), .B(a[66]), .Z(n15076) );
  NANDN U15318 ( .A(n32292), .B(n15076), .Z(n14809) );
  AND U15319 ( .A(n14810), .B(n14809), .Z(n15242) );
  NANDN U15320 ( .A(n31536), .B(n14811), .Z(n14813) );
  XOR U15321 ( .A(b[15]), .B(a[68]), .Z(n15079) );
  NANDN U15322 ( .A(n31925), .B(n15079), .Z(n14812) );
  NAND U15323 ( .A(n14813), .B(n14812), .Z(n15241) );
  XOR U15324 ( .A(n15242), .B(n15241), .Z(n15244) );
  XOR U15325 ( .A(n15243), .B(n15244), .Z(n15215) );
  NANDN U15326 ( .A(n37526), .B(n14814), .Z(n14816) );
  XOR U15327 ( .A(b[51]), .B(a[32]), .Z(n15082) );
  NANDN U15328 ( .A(n37605), .B(n15082), .Z(n14815) );
  AND U15329 ( .A(n14816), .B(n14815), .Z(n15267) );
  NANDN U15330 ( .A(n37705), .B(n14817), .Z(n14819) );
  XOR U15331 ( .A(b[53]), .B(a[30]), .Z(n15085) );
  NANDN U15332 ( .A(n37778), .B(n15085), .Z(n14818) );
  AND U15333 ( .A(n14819), .B(n14818), .Z(n15266) );
  NANDN U15334 ( .A(n36210), .B(n14820), .Z(n14822) );
  XOR U15335 ( .A(b[39]), .B(a[44]), .Z(n15088) );
  NANDN U15336 ( .A(n36347), .B(n15088), .Z(n14821) );
  NAND U15337 ( .A(n14822), .B(n14821), .Z(n15265) );
  XOR U15338 ( .A(n15266), .B(n15265), .Z(n15268) );
  XNOR U15339 ( .A(n15267), .B(n15268), .Z(n15214) );
  XNOR U15340 ( .A(n15215), .B(n15214), .Z(n15217) );
  NANDN U15341 ( .A(n14824), .B(n14823), .Z(n14828) );
  OR U15342 ( .A(n14826), .B(n14825), .Z(n14827) );
  AND U15343 ( .A(n14828), .B(n14827), .Z(n15216) );
  XOR U15344 ( .A(n15217), .B(n15216), .Z(n15064) );
  NANDN U15345 ( .A(n14830), .B(n14829), .Z(n14834) );
  OR U15346 ( .A(n14832), .B(n14831), .Z(n14833) );
  AND U15347 ( .A(n14834), .B(n14833), .Z(n15062) );
  NANDN U15348 ( .A(n14836), .B(n14835), .Z(n14840) );
  NANDN U15349 ( .A(n14838), .B(n14837), .Z(n14839) );
  NAND U15350 ( .A(n14840), .B(n14839), .Z(n15061) );
  XNOR U15351 ( .A(n15062), .B(n15061), .Z(n15063) );
  XNOR U15352 ( .A(n15064), .B(n15063), .Z(n15293) );
  XOR U15353 ( .A(n15294), .B(n15293), .Z(n15296) );
  XOR U15354 ( .A(n15295), .B(n15296), .Z(n15276) );
  NANDN U15355 ( .A(n14842), .B(n14841), .Z(n14846) );
  NANDN U15356 ( .A(n14844), .B(n14843), .Z(n14845) );
  AND U15357 ( .A(n14846), .B(n14845), .Z(n15288) );
  NANDN U15358 ( .A(n14847), .B(n37294), .Z(n14849) );
  XOR U15359 ( .A(b[47]), .B(a[36]), .Z(n15115) );
  NANDN U15360 ( .A(n37172), .B(n15115), .Z(n14848) );
  AND U15361 ( .A(n14849), .B(n14848), .Z(n15156) );
  NANDN U15362 ( .A(n14850), .B(n30627), .Z(n14852) );
  XOR U15363 ( .A(b[9]), .B(a[74]), .Z(n15118) );
  NANDN U15364 ( .A(n30267), .B(n15118), .Z(n14851) );
  AND U15365 ( .A(n14852), .B(n14851), .Z(n15155) );
  NANDN U15366 ( .A(n14853), .B(n37536), .Z(n14855) );
  XOR U15367 ( .A(b[49]), .B(a[34]), .Z(n15121) );
  NANDN U15368 ( .A(n37432), .B(n15121), .Z(n14854) );
  NAND U15369 ( .A(n14855), .B(n14854), .Z(n15154) );
  XOR U15370 ( .A(n15155), .B(n15154), .Z(n15157) );
  XOR U15371 ( .A(n15156), .B(n15157), .Z(n15221) );
  NANDN U15372 ( .A(n36742), .B(n14856), .Z(n14858) );
  XOR U15373 ( .A(b[43]), .B(a[40]), .Z(n15124) );
  NANDN U15374 ( .A(n36891), .B(n15124), .Z(n14857) );
  AND U15375 ( .A(n14858), .B(n14857), .Z(n15135) );
  NANDN U15376 ( .A(n36991), .B(n14859), .Z(n14861) );
  XOR U15377 ( .A(b[45]), .B(a[38]), .Z(n15127) );
  NANDN U15378 ( .A(n37083), .B(n15127), .Z(n14860) );
  AND U15379 ( .A(n14861), .B(n14860), .Z(n15134) );
  NANDN U15380 ( .A(n30482), .B(n14862), .Z(n14864) );
  XOR U15381 ( .A(b[11]), .B(a[72]), .Z(n15130) );
  NANDN U15382 ( .A(n30891), .B(n15130), .Z(n14863) );
  NAND U15383 ( .A(n14864), .B(n14863), .Z(n15133) );
  XOR U15384 ( .A(n15134), .B(n15133), .Z(n15136) );
  XNOR U15385 ( .A(n15135), .B(n15136), .Z(n15220) );
  XNOR U15386 ( .A(n15221), .B(n15220), .Z(n15222) );
  NANDN U15387 ( .A(n14866), .B(n14865), .Z(n14870) );
  OR U15388 ( .A(n14868), .B(n14867), .Z(n14869) );
  NAND U15389 ( .A(n14870), .B(n14869), .Z(n15223) );
  XNOR U15390 ( .A(n15222), .B(n15223), .Z(n15287) );
  XNOR U15391 ( .A(n15288), .B(n15287), .Z(n15289) );
  NANDN U15392 ( .A(n29499), .B(n14871), .Z(n14873) );
  XOR U15393 ( .A(a[76]), .B(b[7]), .Z(n15139) );
  NANDN U15394 ( .A(n29735), .B(n15139), .Z(n14872) );
  AND U15395 ( .A(n14873), .B(n14872), .Z(n15099) );
  NANDN U15396 ( .A(n37857), .B(n14874), .Z(n14876) );
  XOR U15397 ( .A(b[55]), .B(a[28]), .Z(n15142) );
  NANDN U15398 ( .A(n37911), .B(n15142), .Z(n14875) );
  AND U15399 ( .A(n14876), .B(n14875), .Z(n15098) );
  NANDN U15400 ( .A(n35611), .B(n14877), .Z(n14879) );
  XOR U15401 ( .A(b[35]), .B(a[48]), .Z(n15145) );
  NANDN U15402 ( .A(n35801), .B(n15145), .Z(n14878) );
  NAND U15403 ( .A(n14879), .B(n14878), .Z(n15097) );
  XOR U15404 ( .A(n15098), .B(n15097), .Z(n15100) );
  XOR U15405 ( .A(n15099), .B(n15100), .Z(n15173) );
  NANDN U15406 ( .A(n14881), .B(n14880), .Z(n14885) );
  OR U15407 ( .A(n14883), .B(n14882), .Z(n14884) );
  AND U15408 ( .A(n14885), .B(n14884), .Z(n15172) );
  XNOR U15409 ( .A(n15173), .B(n15172), .Z(n15174) );
  NAND U15410 ( .A(n14887), .B(n14886), .Z(n14891) );
  NANDN U15411 ( .A(n14889), .B(n14888), .Z(n14890) );
  NAND U15412 ( .A(n14891), .B(n14890), .Z(n15175) );
  XOR U15413 ( .A(n15174), .B(n15175), .Z(n15290) );
  XNOR U15414 ( .A(n15289), .B(n15290), .Z(n15275) );
  XOR U15415 ( .A(n15276), .B(n15275), .Z(n15278) );
  XOR U15416 ( .A(n15277), .B(n15278), .Z(n15300) );
  NANDN U15417 ( .A(n14893), .B(n14892), .Z(n14897) );
  NANDN U15418 ( .A(n14895), .B(n14894), .Z(n14896) );
  AND U15419 ( .A(n14897), .B(n14896), .Z(n15283) );
  NANDN U15420 ( .A(n14899), .B(n14898), .Z(n14903) );
  NANDN U15421 ( .A(n14901), .B(n14900), .Z(n14902) );
  AND U15422 ( .A(n14903), .B(n14902), .Z(n15282) );
  NANDN U15423 ( .A(n14905), .B(n14904), .Z(n14909) );
  NAND U15424 ( .A(n14907), .B(n14906), .Z(n14908) );
  AND U15425 ( .A(n14909), .B(n14908), .Z(n15281) );
  XOR U15426 ( .A(n15282), .B(n15281), .Z(n15284) );
  XOR U15427 ( .A(n15283), .B(n15284), .Z(n15052) );
  NANDN U15428 ( .A(n14911), .B(n14910), .Z(n14915) );
  NANDN U15429 ( .A(n14913), .B(n14912), .Z(n14914) );
  AND U15430 ( .A(n14915), .B(n14914), .Z(n15167) );
  NANDN U15431 ( .A(n14917), .B(n14916), .Z(n14921) );
  OR U15432 ( .A(n14919), .B(n14918), .Z(n14920) );
  NAND U15433 ( .A(n14921), .B(n14920), .Z(n15166) );
  XNOR U15434 ( .A(n15167), .B(n15166), .Z(n15169) );
  NANDN U15435 ( .A(n14923), .B(n14922), .Z(n14927) );
  OR U15436 ( .A(n14925), .B(n14924), .Z(n14926) );
  NAND U15437 ( .A(n14927), .B(n14926), .Z(n15069) );
  NAND U15438 ( .A(b[0]), .B(a[82]), .Z(n14928) );
  XNOR U15439 ( .A(b[1]), .B(n14928), .Z(n14930) );
  NANDN U15440 ( .A(b[0]), .B(a[81]), .Z(n14929) );
  NAND U15441 ( .A(n14930), .B(n14929), .Z(n15106) );
  NANDN U15442 ( .A(n38278), .B(n14931), .Z(n14933) );
  XOR U15443 ( .A(b[63]), .B(a[20]), .Z(n15199) );
  NANDN U15444 ( .A(n38279), .B(n15199), .Z(n14932) );
  AND U15445 ( .A(n14933), .B(n14932), .Z(n15104) );
  NANDN U15446 ( .A(n35260), .B(n14934), .Z(n14936) );
  XOR U15447 ( .A(b[33]), .B(a[50]), .Z(n15202) );
  NANDN U15448 ( .A(n35456), .B(n15202), .Z(n14935) );
  NAND U15449 ( .A(n14936), .B(n14935), .Z(n15103) );
  XNOR U15450 ( .A(n15104), .B(n15103), .Z(n15105) );
  XNOR U15451 ( .A(n15106), .B(n15105), .Z(n15068) );
  NANDN U15452 ( .A(n37974), .B(n14937), .Z(n14939) );
  XOR U15453 ( .A(b[57]), .B(a[26]), .Z(n15205) );
  NANDN U15454 ( .A(n38031), .B(n15205), .Z(n14938) );
  AND U15455 ( .A(n14939), .B(n14938), .Z(n15180) );
  NANDN U15456 ( .A(n38090), .B(n14940), .Z(n14942) );
  XOR U15457 ( .A(b[59]), .B(a[24]), .Z(n15208) );
  NANDN U15458 ( .A(n38130), .B(n15208), .Z(n14941) );
  AND U15459 ( .A(n14942), .B(n14941), .Z(n15179) );
  NANDN U15460 ( .A(n36480), .B(n14943), .Z(n14945) );
  XOR U15461 ( .A(b[41]), .B(a[42]), .Z(n15211) );
  NANDN U15462 ( .A(n36594), .B(n15211), .Z(n14944) );
  NAND U15463 ( .A(n14945), .B(n14944), .Z(n15178) );
  XOR U15464 ( .A(n15179), .B(n15178), .Z(n15181) );
  XOR U15465 ( .A(n15180), .B(n15181), .Z(n15067) );
  XOR U15466 ( .A(n15068), .B(n15067), .Z(n15070) );
  XOR U15467 ( .A(n15069), .B(n15070), .Z(n15168) );
  XOR U15468 ( .A(n15169), .B(n15168), .Z(n15056) );
  NANDN U15469 ( .A(n14947), .B(n14946), .Z(n14951) );
  NAND U15470 ( .A(n14949), .B(n14948), .Z(n14950) );
  NAND U15471 ( .A(n14951), .B(n14950), .Z(n15055) );
  XNOR U15472 ( .A(n15056), .B(n15055), .Z(n15058) );
  NAND U15473 ( .A(n14953), .B(n14952), .Z(n14957) );
  NANDN U15474 ( .A(n14955), .B(n14954), .Z(n14956) );
  AND U15475 ( .A(n14957), .B(n14956), .Z(n15274) );
  NANDN U15476 ( .A(n14959), .B(n14958), .Z(n14963) );
  OR U15477 ( .A(n14961), .B(n14960), .Z(n14962) );
  AND U15478 ( .A(n14963), .B(n14962), .Z(n15111) );
  NANDN U15479 ( .A(n32996), .B(n14964), .Z(n14966) );
  XOR U15480 ( .A(b[21]), .B(a[62]), .Z(n15226) );
  NANDN U15481 ( .A(n33271), .B(n15226), .Z(n14965) );
  AND U15482 ( .A(n14966), .B(n14965), .Z(n15193) );
  NANDN U15483 ( .A(n33866), .B(n14967), .Z(n14969) );
  XOR U15484 ( .A(b[23]), .B(a[60]), .Z(n15229) );
  NANDN U15485 ( .A(n33644), .B(n15229), .Z(n14968) );
  AND U15486 ( .A(n14969), .B(n14968), .Z(n15191) );
  NANDN U15487 ( .A(n32483), .B(n14970), .Z(n14972) );
  XOR U15488 ( .A(b[19]), .B(a[64]), .Z(n15232) );
  NANDN U15489 ( .A(n32823), .B(n15232), .Z(n14971) );
  NAND U15490 ( .A(n14972), .B(n14971), .Z(n15190) );
  XNOR U15491 ( .A(n15191), .B(n15190), .Z(n15192) );
  XOR U15492 ( .A(n15193), .B(n15192), .Z(n15110) );
  NANDN U15493 ( .A(n34909), .B(n14973), .Z(n14975) );
  XOR U15494 ( .A(b[31]), .B(a[52]), .Z(n15235) );
  NANDN U15495 ( .A(n35145), .B(n15235), .Z(n14974) );
  AND U15496 ( .A(n14975), .B(n14974), .Z(n15151) );
  NANDN U15497 ( .A(n38247), .B(n14976), .Z(n14978) );
  XOR U15498 ( .A(b[61]), .B(a[22]), .Z(n15238) );
  NANDN U15499 ( .A(n38248), .B(n15238), .Z(n14977) );
  AND U15500 ( .A(n14978), .B(n14977), .Z(n15149) );
  AND U15501 ( .A(b[63]), .B(a[18]), .Z(n15148) );
  XNOR U15502 ( .A(n15149), .B(n15148), .Z(n15150) );
  XOR U15503 ( .A(n15151), .B(n15150), .Z(n15109) );
  XNOR U15504 ( .A(n15110), .B(n15109), .Z(n15112) );
  NANDN U15505 ( .A(n14980), .B(n14979), .Z(n14984) );
  OR U15506 ( .A(n14982), .B(n14981), .Z(n14983) );
  AND U15507 ( .A(n14984), .B(n14983), .Z(n15162) );
  NANDN U15508 ( .A(n34223), .B(n14985), .Z(n14987) );
  XOR U15509 ( .A(b[27]), .B(a[56]), .Z(n15247) );
  NANDN U15510 ( .A(n34458), .B(n15247), .Z(n14986) );
  AND U15511 ( .A(n14987), .B(n14986), .Z(n15094) );
  NANDN U15512 ( .A(n34634), .B(n14988), .Z(n14990) );
  XOR U15513 ( .A(b[29]), .B(a[54]), .Z(n15250) );
  NANDN U15514 ( .A(n34722), .B(n15250), .Z(n14989) );
  AND U15515 ( .A(n14990), .B(n14989), .Z(n15092) );
  NANDN U15516 ( .A(n31055), .B(n14991), .Z(n14993) );
  XOR U15517 ( .A(b[13]), .B(a[70]), .Z(n15253) );
  NANDN U15518 ( .A(n31293), .B(n15253), .Z(n14992) );
  NAND U15519 ( .A(n14993), .B(n14992), .Z(n15091) );
  XNOR U15520 ( .A(n15092), .B(n15091), .Z(n15093) );
  XOR U15521 ( .A(n15094), .B(n15093), .Z(n15161) );
  NANDN U15522 ( .A(n28889), .B(n14994), .Z(n14996) );
  XOR U15523 ( .A(a[78]), .B(b[5]), .Z(n15256) );
  NANDN U15524 ( .A(n29138), .B(n15256), .Z(n14995) );
  AND U15525 ( .A(n14996), .B(n14995), .Z(n15187) );
  NANDN U15526 ( .A(n209), .B(n14997), .Z(n14999) );
  XOR U15527 ( .A(a[80]), .B(b[3]), .Z(n15259) );
  NANDN U15528 ( .A(n28941), .B(n15259), .Z(n14998) );
  AND U15529 ( .A(n14999), .B(n14998), .Z(n15185) );
  NANDN U15530 ( .A(n35936), .B(n15000), .Z(n15002) );
  XOR U15531 ( .A(b[37]), .B(a[46]), .Z(n15262) );
  NANDN U15532 ( .A(n36047), .B(n15262), .Z(n15001) );
  NAND U15533 ( .A(n15002), .B(n15001), .Z(n15184) );
  XNOR U15534 ( .A(n15185), .B(n15184), .Z(n15186) );
  XOR U15535 ( .A(n15187), .B(n15186), .Z(n15160) );
  XNOR U15536 ( .A(n15161), .B(n15160), .Z(n15163) );
  XOR U15537 ( .A(n15272), .B(n15271), .Z(n15273) );
  XNOR U15538 ( .A(n15274), .B(n15273), .Z(n15057) );
  XOR U15539 ( .A(n15058), .B(n15057), .Z(n15050) );
  NANDN U15540 ( .A(n15004), .B(n15003), .Z(n15008) );
  NANDN U15541 ( .A(n15006), .B(n15005), .Z(n15007) );
  AND U15542 ( .A(n15008), .B(n15007), .Z(n15049) );
  XNOR U15543 ( .A(n15050), .B(n15049), .Z(n15051) );
  XNOR U15544 ( .A(n15052), .B(n15051), .Z(n15299) );
  XNOR U15545 ( .A(n15300), .B(n15299), .Z(n15301) );
  XOR U15546 ( .A(n15302), .B(n15301), .Z(n15046) );
  XNOR U15547 ( .A(n15045), .B(n15046), .Z(n15039) );
  XOR U15548 ( .A(n15040), .B(n15039), .Z(n15312) );
  NANDN U15549 ( .A(n15010), .B(n15009), .Z(n15014) );
  OR U15550 ( .A(n15012), .B(n15011), .Z(n15013) );
  NAND U15551 ( .A(n15014), .B(n15013), .Z(n15311) );
  XNOR U15552 ( .A(n15312), .B(n15311), .Z(n15313) );
  NANDN U15553 ( .A(n15016), .B(n15015), .Z(n15020) );
  OR U15554 ( .A(n15018), .B(n15017), .Z(n15019) );
  NAND U15555 ( .A(n15020), .B(n15019), .Z(n15314) );
  XNOR U15556 ( .A(n15313), .B(n15314), .Z(n15031) );
  XOR U15557 ( .A(n15032), .B(n15031), .Z(n15034) );
  XOR U15558 ( .A(n15033), .B(n15034), .Z(n15026) );
  XNOR U15559 ( .A(n15026), .B(sreg[146]), .Z(n15028) );
  NANDN U15560 ( .A(sreg[145]), .B(n15021), .Z(n15025) );
  NAND U15561 ( .A(n15023), .B(n15022), .Z(n15024) );
  AND U15562 ( .A(n15025), .B(n15024), .Z(n15027) );
  XOR U15563 ( .A(n15028), .B(n15027), .Z(c[146]) );
  NANDN U15564 ( .A(n15026), .B(sreg[146]), .Z(n15030) );
  NAND U15565 ( .A(n15028), .B(n15027), .Z(n15029) );
  AND U15566 ( .A(n15030), .B(n15029), .Z(n15607) );
  NANDN U15567 ( .A(n15032), .B(n15031), .Z(n15036) );
  OR U15568 ( .A(n15034), .B(n15033), .Z(n15035) );
  AND U15569 ( .A(n15036), .B(n15035), .Z(n15320) );
  NANDN U15570 ( .A(n15038), .B(n15037), .Z(n15042) );
  NAND U15571 ( .A(n15040), .B(n15039), .Z(n15041) );
  AND U15572 ( .A(n15042), .B(n15041), .Z(n15325) );
  NANDN U15573 ( .A(n15044), .B(n15043), .Z(n15048) );
  NANDN U15574 ( .A(n15046), .B(n15045), .Z(n15047) );
  AND U15575 ( .A(n15048), .B(n15047), .Z(n15324) );
  NANDN U15576 ( .A(n15050), .B(n15049), .Z(n15054) );
  NANDN U15577 ( .A(n15052), .B(n15051), .Z(n15053) );
  AND U15578 ( .A(n15054), .B(n15053), .Z(n15331) );
  NANDN U15579 ( .A(n15056), .B(n15055), .Z(n15060) );
  NAND U15580 ( .A(n15058), .B(n15057), .Z(n15059) );
  AND U15581 ( .A(n15060), .B(n15059), .Z(n15343) );
  NANDN U15582 ( .A(n15062), .B(n15061), .Z(n15066) );
  NANDN U15583 ( .A(n15064), .B(n15063), .Z(n15065) );
  AND U15584 ( .A(n15066), .B(n15065), .Z(n15349) );
  NAND U15585 ( .A(n15068), .B(n15067), .Z(n15072) );
  NAND U15586 ( .A(n15070), .B(n15069), .Z(n15071) );
  AND U15587 ( .A(n15072), .B(n15071), .Z(n15348) );
  NANDN U15588 ( .A(n33875), .B(n15073), .Z(n15075) );
  XOR U15589 ( .A(b[25]), .B(a[59]), .Z(n15440) );
  NANDN U15590 ( .A(n33994), .B(n15440), .Z(n15074) );
  AND U15591 ( .A(n15075), .B(n15074), .Z(n15544) );
  NANDN U15592 ( .A(n32013), .B(n15076), .Z(n15078) );
  XOR U15593 ( .A(b[17]), .B(a[67]), .Z(n15443) );
  NANDN U15594 ( .A(n32292), .B(n15443), .Z(n15077) );
  AND U15595 ( .A(n15078), .B(n15077), .Z(n15543) );
  NANDN U15596 ( .A(n31536), .B(n15079), .Z(n15081) );
  XOR U15597 ( .A(b[15]), .B(a[69]), .Z(n15446) );
  NANDN U15598 ( .A(n31925), .B(n15446), .Z(n15080) );
  NAND U15599 ( .A(n15081), .B(n15080), .Z(n15542) );
  XOR U15600 ( .A(n15543), .B(n15542), .Z(n15545) );
  XOR U15601 ( .A(n15544), .B(n15545), .Z(n15531) );
  NANDN U15602 ( .A(n37526), .B(n15082), .Z(n15084) );
  XOR U15603 ( .A(b[51]), .B(a[33]), .Z(n15449) );
  NANDN U15604 ( .A(n37605), .B(n15449), .Z(n15083) );
  AND U15605 ( .A(n15084), .B(n15083), .Z(n15565) );
  NANDN U15606 ( .A(n37705), .B(n15085), .Z(n15087) );
  XOR U15607 ( .A(b[53]), .B(a[31]), .Z(n15452) );
  NANDN U15608 ( .A(n37778), .B(n15452), .Z(n15086) );
  AND U15609 ( .A(n15087), .B(n15086), .Z(n15564) );
  NANDN U15610 ( .A(n36210), .B(n15088), .Z(n15090) );
  XOR U15611 ( .A(b[39]), .B(a[45]), .Z(n15455) );
  NANDN U15612 ( .A(n36347), .B(n15455), .Z(n15089) );
  NAND U15613 ( .A(n15090), .B(n15089), .Z(n15563) );
  XOR U15614 ( .A(n15564), .B(n15563), .Z(n15566) );
  XNOR U15615 ( .A(n15565), .B(n15566), .Z(n15530) );
  XNOR U15616 ( .A(n15531), .B(n15530), .Z(n15533) );
  NANDN U15617 ( .A(n15092), .B(n15091), .Z(n15096) );
  NANDN U15618 ( .A(n15094), .B(n15093), .Z(n15095) );
  AND U15619 ( .A(n15096), .B(n15095), .Z(n15532) );
  XOR U15620 ( .A(n15533), .B(n15532), .Z(n15431) );
  NANDN U15621 ( .A(n15098), .B(n15097), .Z(n15102) );
  OR U15622 ( .A(n15100), .B(n15099), .Z(n15101) );
  AND U15623 ( .A(n15102), .B(n15101), .Z(n15429) );
  NANDN U15624 ( .A(n15104), .B(n15103), .Z(n15108) );
  NANDN U15625 ( .A(n15106), .B(n15105), .Z(n15107) );
  NAND U15626 ( .A(n15108), .B(n15107), .Z(n15428) );
  XNOR U15627 ( .A(n15429), .B(n15428), .Z(n15430) );
  XNOR U15628 ( .A(n15431), .B(n15430), .Z(n15347) );
  XOR U15629 ( .A(n15348), .B(n15347), .Z(n15350) );
  XOR U15630 ( .A(n15349), .B(n15350), .Z(n15342) );
  NAND U15631 ( .A(n15110), .B(n15109), .Z(n15114) );
  NANDN U15632 ( .A(n15112), .B(n15111), .Z(n15113) );
  AND U15633 ( .A(n15114), .B(n15113), .Z(n15354) );
  NAND U15634 ( .A(n37294), .B(n15115), .Z(n15117) );
  XNOR U15635 ( .A(b[47]), .B(a[37]), .Z(n15383) );
  NANDN U15636 ( .A(n15383), .B(n37341), .Z(n15116) );
  NAND U15637 ( .A(n15117), .B(n15116), .Z(n15424) );
  NAND U15638 ( .A(n30627), .B(n15118), .Z(n15120) );
  XNOR U15639 ( .A(b[9]), .B(a[75]), .Z(n15386) );
  NANDN U15640 ( .A(n15386), .B(n30628), .Z(n15119) );
  NAND U15641 ( .A(n15120), .B(n15119), .Z(n15423) );
  NAND U15642 ( .A(n37536), .B(n15121), .Z(n15123) );
  XNOR U15643 ( .A(b[49]), .B(a[35]), .Z(n15389) );
  NANDN U15644 ( .A(n15389), .B(n37537), .Z(n15122) );
  NAND U15645 ( .A(n15123), .B(n15122), .Z(n15422) );
  XNOR U15646 ( .A(n15423), .B(n15422), .Z(n15425) );
  NANDN U15647 ( .A(n36742), .B(n15124), .Z(n15126) );
  XOR U15648 ( .A(b[43]), .B(a[41]), .Z(n15392) );
  NANDN U15649 ( .A(n36891), .B(n15392), .Z(n15125) );
  AND U15650 ( .A(n15126), .B(n15125), .Z(n15403) );
  NANDN U15651 ( .A(n36991), .B(n15127), .Z(n15129) );
  XOR U15652 ( .A(b[45]), .B(a[39]), .Z(n15395) );
  NANDN U15653 ( .A(n37083), .B(n15395), .Z(n15128) );
  AND U15654 ( .A(n15129), .B(n15128), .Z(n15402) );
  NANDN U15655 ( .A(n30482), .B(n15130), .Z(n15132) );
  XOR U15656 ( .A(b[11]), .B(a[73]), .Z(n15398) );
  NANDN U15657 ( .A(n30891), .B(n15398), .Z(n15131) );
  NAND U15658 ( .A(n15132), .B(n15131), .Z(n15401) );
  XOR U15659 ( .A(n15402), .B(n15401), .Z(n15404) );
  XNOR U15660 ( .A(n15403), .B(n15404), .Z(n15536) );
  XOR U15661 ( .A(n15537), .B(n15536), .Z(n15538) );
  NANDN U15662 ( .A(n15134), .B(n15133), .Z(n15138) );
  OR U15663 ( .A(n15136), .B(n15135), .Z(n15137) );
  NAND U15664 ( .A(n15138), .B(n15137), .Z(n15539) );
  XNOR U15665 ( .A(n15538), .B(n15539), .Z(n15353) );
  XNOR U15666 ( .A(n15354), .B(n15353), .Z(n15355) );
  NANDN U15667 ( .A(n29499), .B(n15139), .Z(n15141) );
  XOR U15668 ( .A(a[77]), .B(b[7]), .Z(n15407) );
  NANDN U15669 ( .A(n29735), .B(n15407), .Z(n15140) );
  AND U15670 ( .A(n15141), .B(n15140), .Z(n15466) );
  NANDN U15671 ( .A(n37857), .B(n15142), .Z(n15144) );
  XOR U15672 ( .A(b[55]), .B(a[29]), .Z(n15410) );
  NANDN U15673 ( .A(n37911), .B(n15410), .Z(n15143) );
  AND U15674 ( .A(n15144), .B(n15143), .Z(n15465) );
  NANDN U15675 ( .A(n35611), .B(n15145), .Z(n15147) );
  XOR U15676 ( .A(b[35]), .B(a[49]), .Z(n15413) );
  NANDN U15677 ( .A(n35801), .B(n15413), .Z(n15146) );
  NAND U15678 ( .A(n15147), .B(n15146), .Z(n15464) );
  XOR U15679 ( .A(n15465), .B(n15464), .Z(n15467) );
  XOR U15680 ( .A(n15466), .B(n15467), .Z(n15477) );
  NANDN U15681 ( .A(n15149), .B(n15148), .Z(n15153) );
  NANDN U15682 ( .A(n15151), .B(n15150), .Z(n15152) );
  AND U15683 ( .A(n15153), .B(n15152), .Z(n15476) );
  XNOR U15684 ( .A(n15477), .B(n15476), .Z(n15478) );
  NANDN U15685 ( .A(n15155), .B(n15154), .Z(n15159) );
  OR U15686 ( .A(n15157), .B(n15156), .Z(n15158) );
  NAND U15687 ( .A(n15159), .B(n15158), .Z(n15479) );
  XOR U15688 ( .A(n15478), .B(n15479), .Z(n15356) );
  XNOR U15689 ( .A(n15355), .B(n15356), .Z(n15341) );
  XOR U15690 ( .A(n15342), .B(n15341), .Z(n15344) );
  XOR U15691 ( .A(n15343), .B(n15344), .Z(n15330) );
  NAND U15692 ( .A(n15161), .B(n15160), .Z(n15165) );
  NANDN U15693 ( .A(n15163), .B(n15162), .Z(n15164) );
  NAND U15694 ( .A(n15165), .B(n15164), .Z(n15359) );
  NANDN U15695 ( .A(n15167), .B(n15166), .Z(n15171) );
  NAND U15696 ( .A(n15169), .B(n15168), .Z(n15170) );
  AND U15697 ( .A(n15171), .B(n15170), .Z(n15360) );
  XOR U15698 ( .A(n15359), .B(n15360), .Z(n15362) );
  NANDN U15699 ( .A(n15173), .B(n15172), .Z(n15177) );
  NANDN U15700 ( .A(n15175), .B(n15174), .Z(n15176) );
  NAND U15701 ( .A(n15177), .B(n15176), .Z(n15361) );
  XOR U15702 ( .A(n15362), .B(n15361), .Z(n15368) );
  NANDN U15703 ( .A(n15179), .B(n15178), .Z(n15183) );
  OR U15704 ( .A(n15181), .B(n15180), .Z(n15182) );
  AND U15705 ( .A(n15183), .B(n15182), .Z(n15489) );
  NANDN U15706 ( .A(n15185), .B(n15184), .Z(n15189) );
  NANDN U15707 ( .A(n15187), .B(n15186), .Z(n15188) );
  NAND U15708 ( .A(n15189), .B(n15188), .Z(n15488) );
  XNOR U15709 ( .A(n15489), .B(n15488), .Z(n15491) );
  NANDN U15710 ( .A(n15191), .B(n15190), .Z(n15195) );
  NANDN U15711 ( .A(n15193), .B(n15192), .Z(n15194) );
  AND U15712 ( .A(n15195), .B(n15194), .Z(n15437) );
  NAND U15713 ( .A(b[0]), .B(a[83]), .Z(n15196) );
  XNOR U15714 ( .A(b[1]), .B(n15196), .Z(n15198) );
  NANDN U15715 ( .A(b[0]), .B(a[82]), .Z(n15197) );
  NAND U15716 ( .A(n15198), .B(n15197), .Z(n15473) );
  NANDN U15717 ( .A(n38278), .B(n15199), .Z(n15201) );
  XOR U15718 ( .A(b[63]), .B(a[21]), .Z(n15515) );
  NANDN U15719 ( .A(n38279), .B(n15515), .Z(n15200) );
  AND U15720 ( .A(n15201), .B(n15200), .Z(n15471) );
  NANDN U15721 ( .A(n35260), .B(n15202), .Z(n15204) );
  XOR U15722 ( .A(b[33]), .B(a[51]), .Z(n15518) );
  NANDN U15723 ( .A(n35456), .B(n15518), .Z(n15203) );
  NAND U15724 ( .A(n15204), .B(n15203), .Z(n15470) );
  XNOR U15725 ( .A(n15471), .B(n15470), .Z(n15472) );
  XNOR U15726 ( .A(n15473), .B(n15472), .Z(n15434) );
  NANDN U15727 ( .A(n37974), .B(n15205), .Z(n15207) );
  XOR U15728 ( .A(b[57]), .B(a[27]), .Z(n15521) );
  NANDN U15729 ( .A(n38031), .B(n15521), .Z(n15206) );
  AND U15730 ( .A(n15207), .B(n15206), .Z(n15497) );
  NANDN U15731 ( .A(n38090), .B(n15208), .Z(n15210) );
  XOR U15732 ( .A(b[59]), .B(a[25]), .Z(n15524) );
  NANDN U15733 ( .A(n38130), .B(n15524), .Z(n15209) );
  AND U15734 ( .A(n15210), .B(n15209), .Z(n15495) );
  NANDN U15735 ( .A(n36480), .B(n15211), .Z(n15213) );
  XOR U15736 ( .A(b[41]), .B(a[43]), .Z(n15527) );
  NANDN U15737 ( .A(n36594), .B(n15527), .Z(n15212) );
  NAND U15738 ( .A(n15213), .B(n15212), .Z(n15494) );
  XNOR U15739 ( .A(n15495), .B(n15494), .Z(n15496) );
  XOR U15740 ( .A(n15497), .B(n15496), .Z(n15435) );
  XNOR U15741 ( .A(n15434), .B(n15435), .Z(n15436) );
  XNOR U15742 ( .A(n15437), .B(n15436), .Z(n15490) );
  XOR U15743 ( .A(n15491), .B(n15490), .Z(n15372) );
  NANDN U15744 ( .A(n15215), .B(n15214), .Z(n15219) );
  NAND U15745 ( .A(n15217), .B(n15216), .Z(n15218) );
  NAND U15746 ( .A(n15219), .B(n15218), .Z(n15371) );
  XNOR U15747 ( .A(n15372), .B(n15371), .Z(n15374) );
  NANDN U15748 ( .A(n15221), .B(n15220), .Z(n15225) );
  NANDN U15749 ( .A(n15223), .B(n15222), .Z(n15224) );
  AND U15750 ( .A(n15225), .B(n15224), .Z(n15590) );
  NANDN U15751 ( .A(n32996), .B(n15226), .Z(n15228) );
  XOR U15752 ( .A(b[21]), .B(a[63]), .Z(n15548) );
  NANDN U15753 ( .A(n33271), .B(n15548), .Z(n15227) );
  AND U15754 ( .A(n15228), .B(n15227), .Z(n15508) );
  NANDN U15755 ( .A(n33866), .B(n15229), .Z(n15231) );
  XOR U15756 ( .A(b[23]), .B(a[61]), .Z(n15551) );
  NANDN U15757 ( .A(n33644), .B(n15551), .Z(n15230) );
  AND U15758 ( .A(n15231), .B(n15230), .Z(n15507) );
  NANDN U15759 ( .A(n32483), .B(n15232), .Z(n15234) );
  XOR U15760 ( .A(b[19]), .B(a[65]), .Z(n15554) );
  NANDN U15761 ( .A(n32823), .B(n15554), .Z(n15233) );
  NAND U15762 ( .A(n15234), .B(n15233), .Z(n15506) );
  XOR U15763 ( .A(n15507), .B(n15506), .Z(n15509) );
  XOR U15764 ( .A(n15508), .B(n15509), .Z(n15378) );
  NANDN U15765 ( .A(n34909), .B(n15235), .Z(n15237) );
  XOR U15766 ( .A(b[31]), .B(a[53]), .Z(n15557) );
  NANDN U15767 ( .A(n35145), .B(n15557), .Z(n15236) );
  AND U15768 ( .A(n15237), .B(n15236), .Z(n15418) );
  NANDN U15769 ( .A(n38247), .B(n15238), .Z(n15240) );
  XOR U15770 ( .A(b[61]), .B(a[23]), .Z(n15560) );
  NANDN U15771 ( .A(n38248), .B(n15560), .Z(n15239) );
  AND U15772 ( .A(n15240), .B(n15239), .Z(n15417) );
  AND U15773 ( .A(b[63]), .B(a[19]), .Z(n15416) );
  XOR U15774 ( .A(n15417), .B(n15416), .Z(n15419) );
  XNOR U15775 ( .A(n15418), .B(n15419), .Z(n15377) );
  XNOR U15776 ( .A(n15378), .B(n15377), .Z(n15379) );
  NANDN U15777 ( .A(n15242), .B(n15241), .Z(n15246) );
  OR U15778 ( .A(n15244), .B(n15243), .Z(n15245) );
  NAND U15779 ( .A(n15246), .B(n15245), .Z(n15380) );
  XNOR U15780 ( .A(n15379), .B(n15380), .Z(n15587) );
  NANDN U15781 ( .A(n34223), .B(n15247), .Z(n15249) );
  XOR U15782 ( .A(b[27]), .B(a[57]), .Z(n15569) );
  NANDN U15783 ( .A(n34458), .B(n15569), .Z(n15248) );
  AND U15784 ( .A(n15249), .B(n15248), .Z(n15460) );
  NANDN U15785 ( .A(n34634), .B(n15250), .Z(n15252) );
  XOR U15786 ( .A(b[29]), .B(a[55]), .Z(n15572) );
  NANDN U15787 ( .A(n34722), .B(n15572), .Z(n15251) );
  AND U15788 ( .A(n15252), .B(n15251), .Z(n15459) );
  NANDN U15789 ( .A(n31055), .B(n15253), .Z(n15255) );
  XOR U15790 ( .A(b[13]), .B(a[71]), .Z(n15575) );
  NANDN U15791 ( .A(n31293), .B(n15575), .Z(n15254) );
  NAND U15792 ( .A(n15255), .B(n15254), .Z(n15458) );
  XOR U15793 ( .A(n15459), .B(n15458), .Z(n15461) );
  XOR U15794 ( .A(n15460), .B(n15461), .Z(n15483) );
  NANDN U15795 ( .A(n28889), .B(n15256), .Z(n15258) );
  XOR U15796 ( .A(a[79]), .B(b[5]), .Z(n15578) );
  NANDN U15797 ( .A(n29138), .B(n15578), .Z(n15257) );
  AND U15798 ( .A(n15258), .B(n15257), .Z(n15502) );
  NANDN U15799 ( .A(n209), .B(n15259), .Z(n15261) );
  XOR U15800 ( .A(a[81]), .B(b[3]), .Z(n15581) );
  NANDN U15801 ( .A(n28941), .B(n15581), .Z(n15260) );
  AND U15802 ( .A(n15261), .B(n15260), .Z(n15501) );
  NANDN U15803 ( .A(n35936), .B(n15262), .Z(n15264) );
  XOR U15804 ( .A(b[37]), .B(a[47]), .Z(n15584) );
  NANDN U15805 ( .A(n36047), .B(n15584), .Z(n15263) );
  NAND U15806 ( .A(n15264), .B(n15263), .Z(n15500) );
  XOR U15807 ( .A(n15501), .B(n15500), .Z(n15503) );
  XNOR U15808 ( .A(n15502), .B(n15503), .Z(n15482) );
  XNOR U15809 ( .A(n15483), .B(n15482), .Z(n15484) );
  NANDN U15810 ( .A(n15266), .B(n15265), .Z(n15270) );
  OR U15811 ( .A(n15268), .B(n15267), .Z(n15269) );
  NAND U15812 ( .A(n15270), .B(n15269), .Z(n15485) );
  XOR U15813 ( .A(n15484), .B(n15485), .Z(n15588) );
  XNOR U15814 ( .A(n15587), .B(n15588), .Z(n15589) );
  XNOR U15815 ( .A(n15590), .B(n15589), .Z(n15373) );
  XOR U15816 ( .A(n15374), .B(n15373), .Z(n15366) );
  XNOR U15817 ( .A(n15366), .B(n15365), .Z(n15367) );
  XNOR U15818 ( .A(n15368), .B(n15367), .Z(n15329) );
  XOR U15819 ( .A(n15330), .B(n15329), .Z(n15332) );
  XOR U15820 ( .A(n15331), .B(n15332), .Z(n15595) );
  NANDN U15821 ( .A(n15276), .B(n15275), .Z(n15280) );
  OR U15822 ( .A(n15278), .B(n15277), .Z(n15279) );
  AND U15823 ( .A(n15280), .B(n15279), .Z(n15594) );
  NANDN U15824 ( .A(n15282), .B(n15281), .Z(n15286) );
  OR U15825 ( .A(n15284), .B(n15283), .Z(n15285) );
  AND U15826 ( .A(n15286), .B(n15285), .Z(n15338) );
  NANDN U15827 ( .A(n15288), .B(n15287), .Z(n15292) );
  NANDN U15828 ( .A(n15290), .B(n15289), .Z(n15291) );
  AND U15829 ( .A(n15292), .B(n15291), .Z(n15336) );
  NANDN U15830 ( .A(n15294), .B(n15293), .Z(n15298) );
  OR U15831 ( .A(n15296), .B(n15295), .Z(n15297) );
  AND U15832 ( .A(n15298), .B(n15297), .Z(n15335) );
  XNOR U15833 ( .A(n15336), .B(n15335), .Z(n15337) );
  XNOR U15834 ( .A(n15338), .B(n15337), .Z(n15593) );
  XOR U15835 ( .A(n15594), .B(n15593), .Z(n15596) );
  XOR U15836 ( .A(n15595), .B(n15596), .Z(n15602) );
  NANDN U15837 ( .A(n15300), .B(n15299), .Z(n15304) );
  NANDN U15838 ( .A(n15302), .B(n15301), .Z(n15303) );
  AND U15839 ( .A(n15304), .B(n15303), .Z(n15600) );
  NANDN U15840 ( .A(n15306), .B(n15305), .Z(n15310) );
  NANDN U15841 ( .A(n15308), .B(n15307), .Z(n15309) );
  NAND U15842 ( .A(n15310), .B(n15309), .Z(n15599) );
  XNOR U15843 ( .A(n15600), .B(n15599), .Z(n15601) );
  XNOR U15844 ( .A(n15602), .B(n15601), .Z(n15323) );
  XOR U15845 ( .A(n15324), .B(n15323), .Z(n15326) );
  XOR U15846 ( .A(n15325), .B(n15326), .Z(n15318) );
  NANDN U15847 ( .A(n15312), .B(n15311), .Z(n15316) );
  NANDN U15848 ( .A(n15314), .B(n15313), .Z(n15315) );
  NAND U15849 ( .A(n15316), .B(n15315), .Z(n15317) );
  XNOR U15850 ( .A(n15318), .B(n15317), .Z(n15319) );
  XNOR U15851 ( .A(n15320), .B(n15319), .Z(n15605) );
  XNOR U15852 ( .A(sreg[147]), .B(n15605), .Z(n15606) );
  XNOR U15853 ( .A(n15607), .B(n15606), .Z(c[147]) );
  NANDN U15854 ( .A(n15318), .B(n15317), .Z(n15322) );
  NANDN U15855 ( .A(n15320), .B(n15319), .Z(n15321) );
  AND U15856 ( .A(n15322), .B(n15321), .Z(n15613) );
  NANDN U15857 ( .A(n15324), .B(n15323), .Z(n15328) );
  OR U15858 ( .A(n15326), .B(n15325), .Z(n15327) );
  AND U15859 ( .A(n15328), .B(n15327), .Z(n15610) );
  NANDN U15860 ( .A(n15330), .B(n15329), .Z(n15334) );
  OR U15861 ( .A(n15332), .B(n15331), .Z(n15333) );
  AND U15862 ( .A(n15334), .B(n15333), .Z(n15891) );
  NANDN U15863 ( .A(n15336), .B(n15335), .Z(n15340) );
  NANDN U15864 ( .A(n15338), .B(n15337), .Z(n15339) );
  AND U15865 ( .A(n15340), .B(n15339), .Z(n15890) );
  XNOR U15866 ( .A(n15891), .B(n15890), .Z(n15893) );
  NANDN U15867 ( .A(n15342), .B(n15341), .Z(n15346) );
  OR U15868 ( .A(n15344), .B(n15343), .Z(n15345) );
  AND U15869 ( .A(n15346), .B(n15345), .Z(n15884) );
  NANDN U15870 ( .A(n15348), .B(n15347), .Z(n15352) );
  OR U15871 ( .A(n15350), .B(n15349), .Z(n15351) );
  AND U15872 ( .A(n15352), .B(n15351), .Z(n15629) );
  NANDN U15873 ( .A(n15354), .B(n15353), .Z(n15358) );
  NANDN U15874 ( .A(n15356), .B(n15355), .Z(n15357) );
  AND U15875 ( .A(n15358), .B(n15357), .Z(n15628) );
  XNOR U15876 ( .A(n15629), .B(n15628), .Z(n15630) );
  NAND U15877 ( .A(n15360), .B(n15359), .Z(n15364) );
  NAND U15878 ( .A(n15362), .B(n15361), .Z(n15363) );
  NAND U15879 ( .A(n15364), .B(n15363), .Z(n15631) );
  XOR U15880 ( .A(n15630), .B(n15631), .Z(n15885) );
  XNOR U15881 ( .A(n15884), .B(n15885), .Z(n15886) );
  NANDN U15882 ( .A(n15366), .B(n15365), .Z(n15370) );
  NANDN U15883 ( .A(n15368), .B(n15367), .Z(n15369) );
  AND U15884 ( .A(n15370), .B(n15369), .Z(n15625) );
  NANDN U15885 ( .A(n15372), .B(n15371), .Z(n15376) );
  NAND U15886 ( .A(n15374), .B(n15373), .Z(n15375) );
  AND U15887 ( .A(n15376), .B(n15375), .Z(n15636) );
  NANDN U15888 ( .A(n15378), .B(n15377), .Z(n15382) );
  NANDN U15889 ( .A(n15380), .B(n15379), .Z(n15381) );
  AND U15890 ( .A(n15382), .B(n15381), .Z(n15647) );
  NANDN U15891 ( .A(n15383), .B(n37294), .Z(n15385) );
  XNOR U15892 ( .A(b[47]), .B(a[38]), .Z(n15724) );
  NANDN U15893 ( .A(n15724), .B(n37341), .Z(n15384) );
  NAND U15894 ( .A(n15385), .B(n15384), .Z(n15765) );
  NANDN U15895 ( .A(n15386), .B(n30627), .Z(n15388) );
  XNOR U15896 ( .A(a[76]), .B(b[9]), .Z(n15727) );
  NANDN U15897 ( .A(n15727), .B(n30628), .Z(n15387) );
  NAND U15898 ( .A(n15388), .B(n15387), .Z(n15764) );
  NANDN U15899 ( .A(n15389), .B(n37536), .Z(n15391) );
  XNOR U15900 ( .A(b[49]), .B(a[36]), .Z(n15730) );
  NANDN U15901 ( .A(n15730), .B(n37537), .Z(n15390) );
  NAND U15902 ( .A(n15391), .B(n15390), .Z(n15763) );
  XNOR U15903 ( .A(n15764), .B(n15763), .Z(n15766) );
  NANDN U15904 ( .A(n36742), .B(n15392), .Z(n15394) );
  XOR U15905 ( .A(b[43]), .B(a[42]), .Z(n15733) );
  NANDN U15906 ( .A(n36891), .B(n15733), .Z(n15393) );
  AND U15907 ( .A(n15394), .B(n15393), .Z(n15744) );
  NANDN U15908 ( .A(n36991), .B(n15395), .Z(n15397) );
  XOR U15909 ( .A(b[45]), .B(a[40]), .Z(n15736) );
  NANDN U15910 ( .A(n37083), .B(n15736), .Z(n15396) );
  AND U15911 ( .A(n15397), .B(n15396), .Z(n15743) );
  NANDN U15912 ( .A(n30482), .B(n15398), .Z(n15400) );
  XOR U15913 ( .A(b[11]), .B(a[74]), .Z(n15739) );
  NANDN U15914 ( .A(n30891), .B(n15739), .Z(n15399) );
  NAND U15915 ( .A(n15400), .B(n15399), .Z(n15742) );
  XOR U15916 ( .A(n15743), .B(n15742), .Z(n15745) );
  XNOR U15917 ( .A(n15744), .B(n15745), .Z(n15787) );
  XOR U15918 ( .A(n15788), .B(n15787), .Z(n15789) );
  NANDN U15919 ( .A(n15402), .B(n15401), .Z(n15406) );
  OR U15920 ( .A(n15404), .B(n15403), .Z(n15405) );
  NAND U15921 ( .A(n15406), .B(n15405), .Z(n15790) );
  XNOR U15922 ( .A(n15789), .B(n15790), .Z(n15646) );
  XNOR U15923 ( .A(n15647), .B(n15646), .Z(n15649) );
  NANDN U15924 ( .A(n29499), .B(n15407), .Z(n15409) );
  XOR U15925 ( .A(a[78]), .B(b[7]), .Z(n15748) );
  NANDN U15926 ( .A(n29735), .B(n15748), .Z(n15408) );
  AND U15927 ( .A(n15409), .B(n15408), .Z(n15708) );
  NANDN U15928 ( .A(n37857), .B(n15410), .Z(n15412) );
  XOR U15929 ( .A(b[55]), .B(a[30]), .Z(n15751) );
  NANDN U15930 ( .A(n37911), .B(n15751), .Z(n15411) );
  AND U15931 ( .A(n15412), .B(n15411), .Z(n15707) );
  NANDN U15932 ( .A(n35611), .B(n15413), .Z(n15415) );
  XOR U15933 ( .A(b[35]), .B(a[50]), .Z(n15754) );
  NANDN U15934 ( .A(n35801), .B(n15754), .Z(n15414) );
  NAND U15935 ( .A(n15415), .B(n15414), .Z(n15706) );
  XOR U15936 ( .A(n15707), .B(n15706), .Z(n15709) );
  XOR U15937 ( .A(n15708), .B(n15709), .Z(n15782) );
  NANDN U15938 ( .A(n15417), .B(n15416), .Z(n15421) );
  OR U15939 ( .A(n15419), .B(n15418), .Z(n15420) );
  AND U15940 ( .A(n15421), .B(n15420), .Z(n15781) );
  XNOR U15941 ( .A(n15782), .B(n15781), .Z(n15783) );
  NAND U15942 ( .A(n15423), .B(n15422), .Z(n15427) );
  NANDN U15943 ( .A(n15425), .B(n15424), .Z(n15426) );
  NAND U15944 ( .A(n15427), .B(n15426), .Z(n15784) );
  XNOR U15945 ( .A(n15783), .B(n15784), .Z(n15648) );
  XOR U15946 ( .A(n15649), .B(n15648), .Z(n15635) );
  NANDN U15947 ( .A(n15429), .B(n15428), .Z(n15433) );
  NANDN U15948 ( .A(n15431), .B(n15430), .Z(n15432) );
  AND U15949 ( .A(n15433), .B(n15432), .Z(n15655) );
  NANDN U15950 ( .A(n15435), .B(n15434), .Z(n15439) );
  NANDN U15951 ( .A(n15437), .B(n15436), .Z(n15438) );
  AND U15952 ( .A(n15439), .B(n15438), .Z(n15653) );
  NANDN U15953 ( .A(n33875), .B(n15440), .Z(n15442) );
  XOR U15954 ( .A(b[25]), .B(a[60]), .Z(n15682) );
  NANDN U15955 ( .A(n33994), .B(n15682), .Z(n15441) );
  AND U15956 ( .A(n15442), .B(n15441), .Z(n15795) );
  NANDN U15957 ( .A(n32013), .B(n15443), .Z(n15445) );
  XOR U15958 ( .A(b[17]), .B(a[68]), .Z(n15685) );
  NANDN U15959 ( .A(n32292), .B(n15685), .Z(n15444) );
  AND U15960 ( .A(n15445), .B(n15444), .Z(n15794) );
  NANDN U15961 ( .A(n31536), .B(n15446), .Z(n15448) );
  XOR U15962 ( .A(b[15]), .B(a[70]), .Z(n15688) );
  NANDN U15963 ( .A(n31925), .B(n15688), .Z(n15447) );
  NAND U15964 ( .A(n15448), .B(n15447), .Z(n15793) );
  XOR U15965 ( .A(n15794), .B(n15793), .Z(n15796) );
  XOR U15966 ( .A(n15795), .B(n15796), .Z(n15875) );
  NANDN U15967 ( .A(n37526), .B(n15449), .Z(n15451) );
  XOR U15968 ( .A(b[51]), .B(a[34]), .Z(n15691) );
  NANDN U15969 ( .A(n37605), .B(n15691), .Z(n15450) );
  AND U15970 ( .A(n15451), .B(n15450), .Z(n15816) );
  NANDN U15971 ( .A(n37705), .B(n15452), .Z(n15454) );
  XOR U15972 ( .A(b[53]), .B(a[32]), .Z(n15694) );
  NANDN U15973 ( .A(n37778), .B(n15694), .Z(n15453) );
  AND U15974 ( .A(n15454), .B(n15453), .Z(n15815) );
  NANDN U15975 ( .A(n36210), .B(n15455), .Z(n15457) );
  XOR U15976 ( .A(b[39]), .B(a[46]), .Z(n15697) );
  NANDN U15977 ( .A(n36347), .B(n15697), .Z(n15456) );
  NAND U15978 ( .A(n15457), .B(n15456), .Z(n15814) );
  XOR U15979 ( .A(n15815), .B(n15814), .Z(n15817) );
  XNOR U15980 ( .A(n15816), .B(n15817), .Z(n15874) );
  XNOR U15981 ( .A(n15875), .B(n15874), .Z(n15877) );
  NANDN U15982 ( .A(n15459), .B(n15458), .Z(n15463) );
  OR U15983 ( .A(n15461), .B(n15460), .Z(n15462) );
  AND U15984 ( .A(n15463), .B(n15462), .Z(n15876) );
  XOR U15985 ( .A(n15877), .B(n15876), .Z(n15673) );
  NANDN U15986 ( .A(n15465), .B(n15464), .Z(n15469) );
  OR U15987 ( .A(n15467), .B(n15466), .Z(n15468) );
  AND U15988 ( .A(n15469), .B(n15468), .Z(n15671) );
  NANDN U15989 ( .A(n15471), .B(n15470), .Z(n15475) );
  NANDN U15990 ( .A(n15473), .B(n15472), .Z(n15474) );
  NAND U15991 ( .A(n15475), .B(n15474), .Z(n15670) );
  XNOR U15992 ( .A(n15671), .B(n15670), .Z(n15672) );
  XNOR U15993 ( .A(n15673), .B(n15672), .Z(n15652) );
  XNOR U15994 ( .A(n15653), .B(n15652), .Z(n15654) );
  XNOR U15995 ( .A(n15655), .B(n15654), .Z(n15634) );
  XOR U15996 ( .A(n15635), .B(n15634), .Z(n15637) );
  XNOR U15997 ( .A(n15636), .B(n15637), .Z(n15622) );
  NANDN U15998 ( .A(n15477), .B(n15476), .Z(n15481) );
  NANDN U15999 ( .A(n15479), .B(n15478), .Z(n15480) );
  AND U16000 ( .A(n15481), .B(n15480), .Z(n15642) );
  NANDN U16001 ( .A(n15483), .B(n15482), .Z(n15487) );
  NANDN U16002 ( .A(n15485), .B(n15484), .Z(n15486) );
  AND U16003 ( .A(n15487), .B(n15486), .Z(n15641) );
  NANDN U16004 ( .A(n15489), .B(n15488), .Z(n15493) );
  NAND U16005 ( .A(n15491), .B(n15490), .Z(n15492) );
  AND U16006 ( .A(n15493), .B(n15492), .Z(n15640) );
  XOR U16007 ( .A(n15641), .B(n15640), .Z(n15643) );
  XOR U16008 ( .A(n15642), .B(n15643), .Z(n15661) );
  NANDN U16009 ( .A(n15495), .B(n15494), .Z(n15499) );
  NANDN U16010 ( .A(n15497), .B(n15496), .Z(n15498) );
  AND U16011 ( .A(n15499), .B(n15498), .Z(n15776) );
  NANDN U16012 ( .A(n15501), .B(n15500), .Z(n15505) );
  OR U16013 ( .A(n15503), .B(n15502), .Z(n15504) );
  NAND U16014 ( .A(n15505), .B(n15504), .Z(n15775) );
  XNOR U16015 ( .A(n15776), .B(n15775), .Z(n15778) );
  NANDN U16016 ( .A(n15507), .B(n15506), .Z(n15511) );
  OR U16017 ( .A(n15509), .B(n15508), .Z(n15510) );
  NAND U16018 ( .A(n15511), .B(n15510), .Z(n15678) );
  NAND U16019 ( .A(b[0]), .B(a[84]), .Z(n15512) );
  XNOR U16020 ( .A(b[1]), .B(n15512), .Z(n15514) );
  NANDN U16021 ( .A(b[0]), .B(a[83]), .Z(n15513) );
  NAND U16022 ( .A(n15514), .B(n15513), .Z(n15715) );
  NANDN U16023 ( .A(n38278), .B(n15515), .Z(n15517) );
  XOR U16024 ( .A(b[63]), .B(a[22]), .Z(n15859) );
  NANDN U16025 ( .A(n38279), .B(n15859), .Z(n15516) );
  AND U16026 ( .A(n15517), .B(n15516), .Z(n15713) );
  NANDN U16027 ( .A(n35260), .B(n15518), .Z(n15520) );
  XOR U16028 ( .A(b[33]), .B(a[52]), .Z(n15862) );
  NANDN U16029 ( .A(n35456), .B(n15862), .Z(n15519) );
  NAND U16030 ( .A(n15520), .B(n15519), .Z(n15712) );
  XNOR U16031 ( .A(n15713), .B(n15712), .Z(n15714) );
  XNOR U16032 ( .A(n15715), .B(n15714), .Z(n15677) );
  NANDN U16033 ( .A(n37974), .B(n15521), .Z(n15523) );
  XOR U16034 ( .A(b[57]), .B(a[28]), .Z(n15865) );
  NANDN U16035 ( .A(n38031), .B(n15865), .Z(n15522) );
  AND U16036 ( .A(n15523), .B(n15522), .Z(n15840) );
  NANDN U16037 ( .A(n38090), .B(n15524), .Z(n15526) );
  XOR U16038 ( .A(b[59]), .B(a[26]), .Z(n15868) );
  NANDN U16039 ( .A(n38130), .B(n15868), .Z(n15525) );
  AND U16040 ( .A(n15526), .B(n15525), .Z(n15839) );
  NANDN U16041 ( .A(n36480), .B(n15527), .Z(n15529) );
  XOR U16042 ( .A(b[41]), .B(a[44]), .Z(n15871) );
  NANDN U16043 ( .A(n36594), .B(n15871), .Z(n15528) );
  NAND U16044 ( .A(n15529), .B(n15528), .Z(n15838) );
  XOR U16045 ( .A(n15839), .B(n15838), .Z(n15841) );
  XOR U16046 ( .A(n15840), .B(n15841), .Z(n15676) );
  XOR U16047 ( .A(n15677), .B(n15676), .Z(n15679) );
  XOR U16048 ( .A(n15678), .B(n15679), .Z(n15777) );
  XOR U16049 ( .A(n15778), .B(n15777), .Z(n15665) );
  NANDN U16050 ( .A(n15531), .B(n15530), .Z(n15535) );
  NAND U16051 ( .A(n15533), .B(n15532), .Z(n15534) );
  NAND U16052 ( .A(n15535), .B(n15534), .Z(n15664) );
  XNOR U16053 ( .A(n15665), .B(n15664), .Z(n15667) );
  NAND U16054 ( .A(n15537), .B(n15536), .Z(n15541) );
  NANDN U16055 ( .A(n15539), .B(n15538), .Z(n15540) );
  AND U16056 ( .A(n15541), .B(n15540), .Z(n15883) );
  NANDN U16057 ( .A(n15543), .B(n15542), .Z(n15547) );
  OR U16058 ( .A(n15545), .B(n15544), .Z(n15546) );
  AND U16059 ( .A(n15547), .B(n15546), .Z(n15720) );
  NANDN U16060 ( .A(n32996), .B(n15548), .Z(n15550) );
  XOR U16061 ( .A(b[21]), .B(a[64]), .Z(n15799) );
  NANDN U16062 ( .A(n33271), .B(n15799), .Z(n15549) );
  AND U16063 ( .A(n15550), .B(n15549), .Z(n15853) );
  NANDN U16064 ( .A(n33866), .B(n15551), .Z(n15553) );
  XOR U16065 ( .A(b[23]), .B(a[62]), .Z(n15802) );
  NANDN U16066 ( .A(n33644), .B(n15802), .Z(n15552) );
  AND U16067 ( .A(n15553), .B(n15552), .Z(n15851) );
  NANDN U16068 ( .A(n32483), .B(n15554), .Z(n15556) );
  XOR U16069 ( .A(b[19]), .B(a[66]), .Z(n15805) );
  NANDN U16070 ( .A(n32823), .B(n15805), .Z(n15555) );
  NAND U16071 ( .A(n15556), .B(n15555), .Z(n15850) );
  XNOR U16072 ( .A(n15851), .B(n15850), .Z(n15852) );
  XOR U16073 ( .A(n15853), .B(n15852), .Z(n15719) );
  NANDN U16074 ( .A(n34909), .B(n15557), .Z(n15559) );
  XOR U16075 ( .A(b[31]), .B(a[54]), .Z(n15808) );
  NANDN U16076 ( .A(n35145), .B(n15808), .Z(n15558) );
  AND U16077 ( .A(n15559), .B(n15558), .Z(n15760) );
  NANDN U16078 ( .A(n38247), .B(n15560), .Z(n15562) );
  XOR U16079 ( .A(b[61]), .B(a[24]), .Z(n15811) );
  NANDN U16080 ( .A(n38248), .B(n15811), .Z(n15561) );
  AND U16081 ( .A(n15562), .B(n15561), .Z(n15758) );
  AND U16082 ( .A(b[63]), .B(a[20]), .Z(n15757) );
  XNOR U16083 ( .A(n15758), .B(n15757), .Z(n15759) );
  XOR U16084 ( .A(n15760), .B(n15759), .Z(n15718) );
  XNOR U16085 ( .A(n15719), .B(n15718), .Z(n15721) );
  NANDN U16086 ( .A(n15564), .B(n15563), .Z(n15568) );
  OR U16087 ( .A(n15566), .B(n15565), .Z(n15567) );
  AND U16088 ( .A(n15568), .B(n15567), .Z(n15771) );
  NANDN U16089 ( .A(n34223), .B(n15569), .Z(n15571) );
  XOR U16090 ( .A(b[27]), .B(a[58]), .Z(n15820) );
  NANDN U16091 ( .A(n34458), .B(n15820), .Z(n15570) );
  AND U16092 ( .A(n15571), .B(n15570), .Z(n15703) );
  NANDN U16093 ( .A(n34634), .B(n15572), .Z(n15574) );
  XOR U16094 ( .A(b[29]), .B(a[56]), .Z(n15823) );
  NANDN U16095 ( .A(n34722), .B(n15823), .Z(n15573) );
  AND U16096 ( .A(n15574), .B(n15573), .Z(n15701) );
  NANDN U16097 ( .A(n31055), .B(n15575), .Z(n15577) );
  XOR U16098 ( .A(b[13]), .B(a[72]), .Z(n15826) );
  NANDN U16099 ( .A(n31293), .B(n15826), .Z(n15576) );
  NAND U16100 ( .A(n15577), .B(n15576), .Z(n15700) );
  XNOR U16101 ( .A(n15701), .B(n15700), .Z(n15702) );
  XOR U16102 ( .A(n15703), .B(n15702), .Z(n15770) );
  NANDN U16103 ( .A(n28889), .B(n15578), .Z(n15580) );
  XOR U16104 ( .A(a[80]), .B(b[5]), .Z(n15829) );
  NANDN U16105 ( .A(n29138), .B(n15829), .Z(n15579) );
  AND U16106 ( .A(n15580), .B(n15579), .Z(n15847) );
  NANDN U16107 ( .A(n209), .B(n15581), .Z(n15583) );
  XOR U16108 ( .A(a[82]), .B(b[3]), .Z(n15832) );
  NANDN U16109 ( .A(n28941), .B(n15832), .Z(n15582) );
  AND U16110 ( .A(n15583), .B(n15582), .Z(n15845) );
  NANDN U16111 ( .A(n35936), .B(n15584), .Z(n15586) );
  XOR U16112 ( .A(b[37]), .B(a[48]), .Z(n15835) );
  NANDN U16113 ( .A(n36047), .B(n15835), .Z(n15585) );
  NAND U16114 ( .A(n15586), .B(n15585), .Z(n15844) );
  XNOR U16115 ( .A(n15845), .B(n15844), .Z(n15846) );
  XOR U16116 ( .A(n15847), .B(n15846), .Z(n15769) );
  XNOR U16117 ( .A(n15770), .B(n15769), .Z(n15772) );
  XOR U16118 ( .A(n15881), .B(n15880), .Z(n15882) );
  XNOR U16119 ( .A(n15883), .B(n15882), .Z(n15666) );
  XOR U16120 ( .A(n15667), .B(n15666), .Z(n15659) );
  NANDN U16121 ( .A(n15588), .B(n15587), .Z(n15592) );
  NANDN U16122 ( .A(n15590), .B(n15589), .Z(n15591) );
  AND U16123 ( .A(n15592), .B(n15591), .Z(n15658) );
  XNOR U16124 ( .A(n15659), .B(n15658), .Z(n15660) );
  XOR U16125 ( .A(n15661), .B(n15660), .Z(n15623) );
  XNOR U16126 ( .A(n15622), .B(n15623), .Z(n15624) );
  XOR U16127 ( .A(n15625), .B(n15624), .Z(n15887) );
  XNOR U16128 ( .A(n15886), .B(n15887), .Z(n15892) );
  XOR U16129 ( .A(n15893), .B(n15892), .Z(n15617) );
  NANDN U16130 ( .A(n15594), .B(n15593), .Z(n15598) );
  OR U16131 ( .A(n15596), .B(n15595), .Z(n15597) );
  NAND U16132 ( .A(n15598), .B(n15597), .Z(n15616) );
  XNOR U16133 ( .A(n15617), .B(n15616), .Z(n15618) );
  NANDN U16134 ( .A(n15600), .B(n15599), .Z(n15604) );
  NANDN U16135 ( .A(n15602), .B(n15601), .Z(n15603) );
  NAND U16136 ( .A(n15604), .B(n15603), .Z(n15619) );
  XOR U16137 ( .A(n15618), .B(n15619), .Z(n15611) );
  XNOR U16138 ( .A(n15610), .B(n15611), .Z(n15612) );
  XNOR U16139 ( .A(n15613), .B(n15612), .Z(n15896) );
  XNOR U16140 ( .A(sreg[148]), .B(n15896), .Z(n15898) );
  NANDN U16141 ( .A(sreg[147]), .B(n15605), .Z(n15609) );
  NAND U16142 ( .A(n15607), .B(n15606), .Z(n15608) );
  NAND U16143 ( .A(n15609), .B(n15608), .Z(n15897) );
  XNOR U16144 ( .A(n15898), .B(n15897), .Z(c[148]) );
  NANDN U16145 ( .A(n15611), .B(n15610), .Z(n15615) );
  NANDN U16146 ( .A(n15613), .B(n15612), .Z(n15614) );
  AND U16147 ( .A(n15615), .B(n15614), .Z(n15908) );
  NANDN U16148 ( .A(n15617), .B(n15616), .Z(n15621) );
  NANDN U16149 ( .A(n15619), .B(n15618), .Z(n15620) );
  AND U16150 ( .A(n15621), .B(n15620), .Z(n15907) );
  NANDN U16151 ( .A(n15623), .B(n15622), .Z(n15627) );
  NANDN U16152 ( .A(n15625), .B(n15624), .Z(n15626) );
  AND U16153 ( .A(n15627), .B(n15626), .Z(n16187) );
  NANDN U16154 ( .A(n15629), .B(n15628), .Z(n15633) );
  NANDN U16155 ( .A(n15631), .B(n15630), .Z(n15632) );
  NAND U16156 ( .A(n15633), .B(n15632), .Z(n16186) );
  XNOR U16157 ( .A(n16187), .B(n16186), .Z(n16189) );
  NANDN U16158 ( .A(n15635), .B(n15634), .Z(n15639) );
  NANDN U16159 ( .A(n15637), .B(n15636), .Z(n15638) );
  AND U16160 ( .A(n15639), .B(n15638), .Z(n16181) );
  NANDN U16161 ( .A(n15641), .B(n15640), .Z(n15645) );
  OR U16162 ( .A(n15643), .B(n15642), .Z(n15644) );
  AND U16163 ( .A(n15645), .B(n15644), .Z(n16176) );
  NANDN U16164 ( .A(n15647), .B(n15646), .Z(n15651) );
  NAND U16165 ( .A(n15649), .B(n15648), .Z(n15650) );
  AND U16166 ( .A(n15651), .B(n15650), .Z(n16175) );
  NANDN U16167 ( .A(n15653), .B(n15652), .Z(n15657) );
  NANDN U16168 ( .A(n15655), .B(n15654), .Z(n15656) );
  AND U16169 ( .A(n15657), .B(n15656), .Z(n16174) );
  XOR U16170 ( .A(n16175), .B(n16174), .Z(n16177) );
  XNOR U16171 ( .A(n16176), .B(n16177), .Z(n16180) );
  XNOR U16172 ( .A(n16181), .B(n16180), .Z(n16182) );
  NANDN U16173 ( .A(n15659), .B(n15658), .Z(n15663) );
  NANDN U16174 ( .A(n15661), .B(n15660), .Z(n15662) );
  AND U16175 ( .A(n15663), .B(n15662), .Z(n16171) );
  NANDN U16176 ( .A(n15665), .B(n15664), .Z(n15669) );
  NAND U16177 ( .A(n15667), .B(n15666), .Z(n15668) );
  AND U16178 ( .A(n15669), .B(n15668), .Z(n16164) );
  NANDN U16179 ( .A(n15671), .B(n15670), .Z(n15675) );
  NANDN U16180 ( .A(n15673), .B(n15672), .Z(n15674) );
  AND U16181 ( .A(n15675), .B(n15674), .Z(n16152) );
  NAND U16182 ( .A(n15677), .B(n15676), .Z(n15681) );
  NAND U16183 ( .A(n15679), .B(n15678), .Z(n15680) );
  AND U16184 ( .A(n15681), .B(n15680), .Z(n16151) );
  NANDN U16185 ( .A(n33875), .B(n15682), .Z(n15684) );
  XOR U16186 ( .A(b[25]), .B(a[61]), .Z(n15987) );
  NANDN U16187 ( .A(n33994), .B(n15987), .Z(n15683) );
  AND U16188 ( .A(n15684), .B(n15683), .Z(n16112) );
  NANDN U16189 ( .A(n32013), .B(n15685), .Z(n15687) );
  XOR U16190 ( .A(b[17]), .B(a[69]), .Z(n15990) );
  NANDN U16191 ( .A(n32292), .B(n15990), .Z(n15686) );
  AND U16192 ( .A(n15687), .B(n15686), .Z(n16111) );
  NANDN U16193 ( .A(n31536), .B(n15688), .Z(n15690) );
  XOR U16194 ( .A(b[15]), .B(a[71]), .Z(n15993) );
  NANDN U16195 ( .A(n31925), .B(n15993), .Z(n15689) );
  NAND U16196 ( .A(n15690), .B(n15689), .Z(n16110) );
  XOR U16197 ( .A(n16111), .B(n16110), .Z(n16113) );
  XOR U16198 ( .A(n16112), .B(n16113), .Z(n16084) );
  NANDN U16199 ( .A(n37526), .B(n15691), .Z(n15693) );
  XOR U16200 ( .A(b[51]), .B(a[35]), .Z(n15996) );
  NANDN U16201 ( .A(n37605), .B(n15996), .Z(n15692) );
  AND U16202 ( .A(n15693), .B(n15692), .Z(n16136) );
  NANDN U16203 ( .A(n37705), .B(n15694), .Z(n15696) );
  XOR U16204 ( .A(b[53]), .B(a[33]), .Z(n15999) );
  NANDN U16205 ( .A(n37778), .B(n15999), .Z(n15695) );
  AND U16206 ( .A(n15696), .B(n15695), .Z(n16135) );
  NANDN U16207 ( .A(n36210), .B(n15697), .Z(n15699) );
  XOR U16208 ( .A(b[39]), .B(a[47]), .Z(n16002) );
  NANDN U16209 ( .A(n36347), .B(n16002), .Z(n15698) );
  NAND U16210 ( .A(n15699), .B(n15698), .Z(n16134) );
  XOR U16211 ( .A(n16135), .B(n16134), .Z(n16137) );
  XNOR U16212 ( .A(n16136), .B(n16137), .Z(n16083) );
  XNOR U16213 ( .A(n16084), .B(n16083), .Z(n16086) );
  NANDN U16214 ( .A(n15701), .B(n15700), .Z(n15705) );
  NANDN U16215 ( .A(n15703), .B(n15702), .Z(n15704) );
  AND U16216 ( .A(n15705), .B(n15704), .Z(n16085) );
  XOR U16217 ( .A(n16086), .B(n16085), .Z(n15978) );
  NANDN U16218 ( .A(n15707), .B(n15706), .Z(n15711) );
  OR U16219 ( .A(n15709), .B(n15708), .Z(n15710) );
  AND U16220 ( .A(n15711), .B(n15710), .Z(n15976) );
  NANDN U16221 ( .A(n15713), .B(n15712), .Z(n15717) );
  NANDN U16222 ( .A(n15715), .B(n15714), .Z(n15716) );
  NAND U16223 ( .A(n15717), .B(n15716), .Z(n15975) );
  XNOR U16224 ( .A(n15976), .B(n15975), .Z(n15977) );
  XNOR U16225 ( .A(n15978), .B(n15977), .Z(n16150) );
  XOR U16226 ( .A(n16151), .B(n16150), .Z(n16153) );
  XOR U16227 ( .A(n16152), .B(n16153), .Z(n16163) );
  NAND U16228 ( .A(n15719), .B(n15718), .Z(n15723) );
  NANDN U16229 ( .A(n15721), .B(n15720), .Z(n15722) );
  AND U16230 ( .A(n15723), .B(n15722), .Z(n16157) );
  NANDN U16231 ( .A(n15724), .B(n37294), .Z(n15726) );
  XOR U16232 ( .A(b[47]), .B(a[39]), .Z(n15930) );
  NANDN U16233 ( .A(n37172), .B(n15930), .Z(n15725) );
  AND U16234 ( .A(n15726), .B(n15725), .Z(n15971) );
  NANDN U16235 ( .A(n15727), .B(n30627), .Z(n15729) );
  XOR U16236 ( .A(a[77]), .B(b[9]), .Z(n15933) );
  NANDN U16237 ( .A(n30267), .B(n15933), .Z(n15728) );
  AND U16238 ( .A(n15729), .B(n15728), .Z(n15970) );
  NANDN U16239 ( .A(n15730), .B(n37536), .Z(n15732) );
  XOR U16240 ( .A(b[49]), .B(a[37]), .Z(n15936) );
  NANDN U16241 ( .A(n37432), .B(n15936), .Z(n15731) );
  NAND U16242 ( .A(n15732), .B(n15731), .Z(n15969) );
  XOR U16243 ( .A(n15970), .B(n15969), .Z(n15972) );
  XOR U16244 ( .A(n15971), .B(n15972), .Z(n16090) );
  NANDN U16245 ( .A(n36742), .B(n15733), .Z(n15735) );
  XOR U16246 ( .A(b[43]), .B(a[43]), .Z(n15939) );
  NANDN U16247 ( .A(n36891), .B(n15939), .Z(n15734) );
  AND U16248 ( .A(n15735), .B(n15734), .Z(n15950) );
  NANDN U16249 ( .A(n36991), .B(n15736), .Z(n15738) );
  XOR U16250 ( .A(b[45]), .B(a[41]), .Z(n15942) );
  NANDN U16251 ( .A(n37083), .B(n15942), .Z(n15737) );
  AND U16252 ( .A(n15738), .B(n15737), .Z(n15949) );
  NANDN U16253 ( .A(n30482), .B(n15739), .Z(n15741) );
  XOR U16254 ( .A(b[11]), .B(a[75]), .Z(n15945) );
  NANDN U16255 ( .A(n30891), .B(n15945), .Z(n15740) );
  NAND U16256 ( .A(n15741), .B(n15740), .Z(n15948) );
  XOR U16257 ( .A(n15949), .B(n15948), .Z(n15951) );
  XNOR U16258 ( .A(n15950), .B(n15951), .Z(n16089) );
  XNOR U16259 ( .A(n16090), .B(n16089), .Z(n16091) );
  NANDN U16260 ( .A(n15743), .B(n15742), .Z(n15747) );
  OR U16261 ( .A(n15745), .B(n15744), .Z(n15746) );
  NAND U16262 ( .A(n15747), .B(n15746), .Z(n16092) );
  XNOR U16263 ( .A(n16091), .B(n16092), .Z(n16156) );
  XNOR U16264 ( .A(n16157), .B(n16156), .Z(n16158) );
  NANDN U16265 ( .A(n29499), .B(n15748), .Z(n15750) );
  XOR U16266 ( .A(a[79]), .B(b[7]), .Z(n15954) );
  NANDN U16267 ( .A(n29735), .B(n15954), .Z(n15749) );
  AND U16268 ( .A(n15750), .B(n15749), .Z(n16013) );
  NANDN U16269 ( .A(n37857), .B(n15751), .Z(n15753) );
  XOR U16270 ( .A(b[55]), .B(a[31]), .Z(n15957) );
  NANDN U16271 ( .A(n37911), .B(n15957), .Z(n15752) );
  AND U16272 ( .A(n15753), .B(n15752), .Z(n16012) );
  NANDN U16273 ( .A(n35611), .B(n15754), .Z(n15756) );
  XOR U16274 ( .A(b[35]), .B(a[51]), .Z(n15960) );
  NANDN U16275 ( .A(n35801), .B(n15960), .Z(n15755) );
  NAND U16276 ( .A(n15756), .B(n15755), .Z(n16011) );
  XOR U16277 ( .A(n16012), .B(n16011), .Z(n16014) );
  XOR U16278 ( .A(n16013), .B(n16014), .Z(n16042) );
  NANDN U16279 ( .A(n15758), .B(n15757), .Z(n15762) );
  NANDN U16280 ( .A(n15760), .B(n15759), .Z(n15761) );
  AND U16281 ( .A(n15762), .B(n15761), .Z(n16041) );
  XNOR U16282 ( .A(n16042), .B(n16041), .Z(n16043) );
  NAND U16283 ( .A(n15764), .B(n15763), .Z(n15768) );
  NANDN U16284 ( .A(n15766), .B(n15765), .Z(n15767) );
  NAND U16285 ( .A(n15768), .B(n15767), .Z(n16044) );
  XOR U16286 ( .A(n16043), .B(n16044), .Z(n16159) );
  XNOR U16287 ( .A(n16158), .B(n16159), .Z(n16162) );
  XOR U16288 ( .A(n16163), .B(n16162), .Z(n16165) );
  XOR U16289 ( .A(n16164), .B(n16165), .Z(n16169) );
  NAND U16290 ( .A(n15770), .B(n15769), .Z(n15774) );
  NANDN U16291 ( .A(n15772), .B(n15771), .Z(n15773) );
  NAND U16292 ( .A(n15774), .B(n15773), .Z(n16144) );
  NANDN U16293 ( .A(n15776), .B(n15775), .Z(n15780) );
  NAND U16294 ( .A(n15778), .B(n15777), .Z(n15779) );
  AND U16295 ( .A(n15780), .B(n15779), .Z(n16145) );
  XOR U16296 ( .A(n16144), .B(n16145), .Z(n16147) );
  NANDN U16297 ( .A(n15782), .B(n15781), .Z(n15786) );
  NANDN U16298 ( .A(n15784), .B(n15783), .Z(n15785) );
  NAND U16299 ( .A(n15786), .B(n15785), .Z(n16146) );
  XOR U16300 ( .A(n16147), .B(n16146), .Z(n15921) );
  NAND U16301 ( .A(n15788), .B(n15787), .Z(n15792) );
  NANDN U16302 ( .A(n15790), .B(n15789), .Z(n15791) );
  AND U16303 ( .A(n15792), .B(n15791), .Z(n16143) );
  NANDN U16304 ( .A(n15794), .B(n15793), .Z(n15798) );
  OR U16305 ( .A(n15796), .B(n15795), .Z(n15797) );
  AND U16306 ( .A(n15798), .B(n15797), .Z(n15926) );
  NANDN U16307 ( .A(n32996), .B(n15799), .Z(n15801) );
  XOR U16308 ( .A(b[21]), .B(a[65]), .Z(n16095) );
  NANDN U16309 ( .A(n33271), .B(n16095), .Z(n15800) );
  AND U16310 ( .A(n15801), .B(n15800), .Z(n16062) );
  NANDN U16311 ( .A(n33866), .B(n15802), .Z(n15804) );
  XOR U16312 ( .A(b[23]), .B(a[63]), .Z(n16098) );
  NANDN U16313 ( .A(n33644), .B(n16098), .Z(n15803) );
  AND U16314 ( .A(n15804), .B(n15803), .Z(n16060) );
  NANDN U16315 ( .A(n32483), .B(n15805), .Z(n15807) );
  XOR U16316 ( .A(b[19]), .B(a[67]), .Z(n16101) );
  NANDN U16317 ( .A(n32823), .B(n16101), .Z(n15806) );
  NAND U16318 ( .A(n15807), .B(n15806), .Z(n16059) );
  XNOR U16319 ( .A(n16060), .B(n16059), .Z(n16061) );
  XOR U16320 ( .A(n16062), .B(n16061), .Z(n15925) );
  NANDN U16321 ( .A(n34909), .B(n15808), .Z(n15810) );
  XOR U16322 ( .A(b[31]), .B(a[55]), .Z(n16104) );
  NANDN U16323 ( .A(n35145), .B(n16104), .Z(n15809) );
  AND U16324 ( .A(n15810), .B(n15809), .Z(n15966) );
  NANDN U16325 ( .A(n38247), .B(n15811), .Z(n15813) );
  XOR U16326 ( .A(b[61]), .B(a[25]), .Z(n16107) );
  NANDN U16327 ( .A(n38248), .B(n16107), .Z(n15812) );
  AND U16328 ( .A(n15813), .B(n15812), .Z(n15964) );
  AND U16329 ( .A(b[63]), .B(a[21]), .Z(n15963) );
  XNOR U16330 ( .A(n15964), .B(n15963), .Z(n15965) );
  XOR U16331 ( .A(n15966), .B(n15965), .Z(n15924) );
  XNOR U16332 ( .A(n15925), .B(n15924), .Z(n15927) );
  NANDN U16333 ( .A(n15815), .B(n15814), .Z(n15819) );
  OR U16334 ( .A(n15817), .B(n15816), .Z(n15818) );
  AND U16335 ( .A(n15819), .B(n15818), .Z(n16031) );
  NANDN U16336 ( .A(n34223), .B(n15820), .Z(n15822) );
  XOR U16337 ( .A(b[27]), .B(a[59]), .Z(n16116) );
  NANDN U16338 ( .A(n34458), .B(n16116), .Z(n15821) );
  AND U16339 ( .A(n15822), .B(n15821), .Z(n16008) );
  NANDN U16340 ( .A(n34634), .B(n15823), .Z(n15825) );
  XOR U16341 ( .A(b[29]), .B(a[57]), .Z(n16119) );
  NANDN U16342 ( .A(n34722), .B(n16119), .Z(n15824) );
  AND U16343 ( .A(n15825), .B(n15824), .Z(n16006) );
  NANDN U16344 ( .A(n31055), .B(n15826), .Z(n15828) );
  XOR U16345 ( .A(b[13]), .B(a[73]), .Z(n16122) );
  NANDN U16346 ( .A(n31293), .B(n16122), .Z(n15827) );
  NAND U16347 ( .A(n15828), .B(n15827), .Z(n16005) );
  XNOR U16348 ( .A(n16006), .B(n16005), .Z(n16007) );
  XOR U16349 ( .A(n16008), .B(n16007), .Z(n16030) );
  NANDN U16350 ( .A(n28889), .B(n15829), .Z(n15831) );
  XOR U16351 ( .A(a[81]), .B(b[5]), .Z(n16125) );
  NANDN U16352 ( .A(n29138), .B(n16125), .Z(n15830) );
  AND U16353 ( .A(n15831), .B(n15830), .Z(n16056) );
  NANDN U16354 ( .A(n209), .B(n15832), .Z(n15834) );
  XOR U16355 ( .A(a[83]), .B(b[3]), .Z(n16128) );
  NANDN U16356 ( .A(n28941), .B(n16128), .Z(n15833) );
  AND U16357 ( .A(n15834), .B(n15833), .Z(n16054) );
  NANDN U16358 ( .A(n35936), .B(n15835), .Z(n15837) );
  XOR U16359 ( .A(b[37]), .B(a[49]), .Z(n16131) );
  NANDN U16360 ( .A(n36047), .B(n16131), .Z(n15836) );
  NAND U16361 ( .A(n15837), .B(n15836), .Z(n16053) );
  XNOR U16362 ( .A(n16054), .B(n16053), .Z(n16055) );
  XOR U16363 ( .A(n16056), .B(n16055), .Z(n16029) );
  XNOR U16364 ( .A(n16030), .B(n16029), .Z(n16032) );
  XOR U16365 ( .A(n16141), .B(n16140), .Z(n16142) );
  XNOR U16366 ( .A(n16143), .B(n16142), .Z(n16026) );
  NANDN U16367 ( .A(n15839), .B(n15838), .Z(n15843) );
  OR U16368 ( .A(n15841), .B(n15840), .Z(n15842) );
  AND U16369 ( .A(n15843), .B(n15842), .Z(n16036) );
  NANDN U16370 ( .A(n15845), .B(n15844), .Z(n15849) );
  NANDN U16371 ( .A(n15847), .B(n15846), .Z(n15848) );
  NAND U16372 ( .A(n15849), .B(n15848), .Z(n16035) );
  XNOR U16373 ( .A(n16036), .B(n16035), .Z(n16038) );
  NANDN U16374 ( .A(n15851), .B(n15850), .Z(n15855) );
  NANDN U16375 ( .A(n15853), .B(n15852), .Z(n15854) );
  NAND U16376 ( .A(n15855), .B(n15854), .Z(n15983) );
  NAND U16377 ( .A(b[0]), .B(a[85]), .Z(n15856) );
  XNOR U16378 ( .A(b[1]), .B(n15856), .Z(n15858) );
  NANDN U16379 ( .A(b[0]), .B(a[84]), .Z(n15857) );
  NAND U16380 ( .A(n15858), .B(n15857), .Z(n16020) );
  NANDN U16381 ( .A(n38278), .B(n15859), .Z(n15861) );
  XOR U16382 ( .A(b[63]), .B(a[23]), .Z(n16068) );
  NANDN U16383 ( .A(n38279), .B(n16068), .Z(n15860) );
  AND U16384 ( .A(n15861), .B(n15860), .Z(n16018) );
  NANDN U16385 ( .A(n35260), .B(n15862), .Z(n15864) );
  XOR U16386 ( .A(b[33]), .B(a[53]), .Z(n16071) );
  NANDN U16387 ( .A(n35456), .B(n16071), .Z(n15863) );
  NAND U16388 ( .A(n15864), .B(n15863), .Z(n16017) );
  XNOR U16389 ( .A(n16018), .B(n16017), .Z(n16019) );
  XNOR U16390 ( .A(n16020), .B(n16019), .Z(n15982) );
  NANDN U16391 ( .A(n37974), .B(n15865), .Z(n15867) );
  XOR U16392 ( .A(b[57]), .B(a[29]), .Z(n16074) );
  NANDN U16393 ( .A(n38031), .B(n16074), .Z(n15866) );
  AND U16394 ( .A(n15867), .B(n15866), .Z(n16049) );
  NANDN U16395 ( .A(n38090), .B(n15868), .Z(n15870) );
  XOR U16396 ( .A(b[59]), .B(a[27]), .Z(n16077) );
  NANDN U16397 ( .A(n38130), .B(n16077), .Z(n15869) );
  AND U16398 ( .A(n15870), .B(n15869), .Z(n16048) );
  NANDN U16399 ( .A(n36480), .B(n15871), .Z(n15873) );
  XOR U16400 ( .A(b[41]), .B(a[45]), .Z(n16080) );
  NANDN U16401 ( .A(n36594), .B(n16080), .Z(n15872) );
  NAND U16402 ( .A(n15873), .B(n15872), .Z(n16047) );
  XOR U16403 ( .A(n16048), .B(n16047), .Z(n16050) );
  XOR U16404 ( .A(n16049), .B(n16050), .Z(n15981) );
  XOR U16405 ( .A(n15982), .B(n15981), .Z(n15984) );
  XOR U16406 ( .A(n15983), .B(n15984), .Z(n16037) );
  XOR U16407 ( .A(n16038), .B(n16037), .Z(n16024) );
  NANDN U16408 ( .A(n15875), .B(n15874), .Z(n15879) );
  NAND U16409 ( .A(n15877), .B(n15876), .Z(n15878) );
  NAND U16410 ( .A(n15879), .B(n15878), .Z(n16023) );
  XNOR U16411 ( .A(n16024), .B(n16023), .Z(n16025) );
  XOR U16412 ( .A(n16026), .B(n16025), .Z(n15919) );
  XNOR U16413 ( .A(n15919), .B(n15918), .Z(n15920) );
  XNOR U16414 ( .A(n15921), .B(n15920), .Z(n16168) );
  XNOR U16415 ( .A(n16169), .B(n16168), .Z(n16170) );
  XOR U16416 ( .A(n16171), .B(n16170), .Z(n16183) );
  XNOR U16417 ( .A(n16182), .B(n16183), .Z(n16188) );
  XOR U16418 ( .A(n16189), .B(n16188), .Z(n15913) );
  NANDN U16419 ( .A(n15885), .B(n15884), .Z(n15889) );
  NANDN U16420 ( .A(n15887), .B(n15886), .Z(n15888) );
  AND U16421 ( .A(n15889), .B(n15888), .Z(n15912) );
  XNOR U16422 ( .A(n15913), .B(n15912), .Z(n15914) );
  NANDN U16423 ( .A(n15891), .B(n15890), .Z(n15895) );
  NAND U16424 ( .A(n15893), .B(n15892), .Z(n15894) );
  NAND U16425 ( .A(n15895), .B(n15894), .Z(n15915) );
  XNOR U16426 ( .A(n15914), .B(n15915), .Z(n15906) );
  XOR U16427 ( .A(n15907), .B(n15906), .Z(n15909) );
  XOR U16428 ( .A(n15908), .B(n15909), .Z(n15901) );
  XNOR U16429 ( .A(n15901), .B(sreg[149]), .Z(n15903) );
  NANDN U16430 ( .A(sreg[148]), .B(n15896), .Z(n15900) );
  NAND U16431 ( .A(n15898), .B(n15897), .Z(n15899) );
  AND U16432 ( .A(n15900), .B(n15899), .Z(n15902) );
  XOR U16433 ( .A(n15903), .B(n15902), .Z(c[149]) );
  NANDN U16434 ( .A(n15901), .B(sreg[149]), .Z(n15905) );
  NAND U16435 ( .A(n15903), .B(n15902), .Z(n15904) );
  AND U16436 ( .A(n15905), .B(n15904), .Z(n16482) );
  NANDN U16437 ( .A(n15907), .B(n15906), .Z(n15911) );
  OR U16438 ( .A(n15909), .B(n15908), .Z(n15910) );
  AND U16439 ( .A(n15911), .B(n15910), .Z(n16195) );
  NANDN U16440 ( .A(n15913), .B(n15912), .Z(n15917) );
  NANDN U16441 ( .A(n15915), .B(n15914), .Z(n15916) );
  AND U16442 ( .A(n15917), .B(n15916), .Z(n16193) );
  NANDN U16443 ( .A(n15919), .B(n15918), .Z(n15923) );
  NANDN U16444 ( .A(n15921), .B(n15920), .Z(n15922) );
  AND U16445 ( .A(n15923), .B(n15922), .Z(n16470) );
  NAND U16446 ( .A(n15925), .B(n15924), .Z(n15929) );
  NANDN U16447 ( .A(n15927), .B(n15926), .Z(n15928) );
  AND U16448 ( .A(n15929), .B(n15928), .Z(n16235) );
  NANDN U16449 ( .A(n211), .B(n15930), .Z(n15932) );
  XOR U16450 ( .A(b[47]), .B(a[40]), .Z(n16327) );
  NANDN U16451 ( .A(n37172), .B(n16327), .Z(n15931) );
  AND U16452 ( .A(n15932), .B(n15931), .Z(n16317) );
  NANDN U16453 ( .A(n210), .B(n15933), .Z(n15935) );
  XOR U16454 ( .A(a[78]), .B(b[9]), .Z(n16330) );
  NANDN U16455 ( .A(n30267), .B(n16330), .Z(n15934) );
  AND U16456 ( .A(n15935), .B(n15934), .Z(n16316) );
  NANDN U16457 ( .A(n212), .B(n15936), .Z(n15938) );
  XOR U16458 ( .A(b[49]), .B(a[38]), .Z(n16333) );
  NANDN U16459 ( .A(n37432), .B(n16333), .Z(n15937) );
  NAND U16460 ( .A(n15938), .B(n15937), .Z(n16315) );
  XOR U16461 ( .A(n16316), .B(n16315), .Z(n16318) );
  XOR U16462 ( .A(n16317), .B(n16318), .Z(n16412) );
  NANDN U16463 ( .A(n36742), .B(n15939), .Z(n15941) );
  XOR U16464 ( .A(b[43]), .B(a[44]), .Z(n16336) );
  NANDN U16465 ( .A(n36891), .B(n16336), .Z(n15940) );
  AND U16466 ( .A(n15941), .B(n15940), .Z(n16347) );
  NANDN U16467 ( .A(n36991), .B(n15942), .Z(n15944) );
  XOR U16468 ( .A(b[45]), .B(a[42]), .Z(n16339) );
  NANDN U16469 ( .A(n37083), .B(n16339), .Z(n15943) );
  AND U16470 ( .A(n15944), .B(n15943), .Z(n16346) );
  NANDN U16471 ( .A(n30482), .B(n15945), .Z(n15947) );
  XOR U16472 ( .A(a[76]), .B(b[11]), .Z(n16342) );
  NANDN U16473 ( .A(n30891), .B(n16342), .Z(n15946) );
  NAND U16474 ( .A(n15947), .B(n15946), .Z(n16345) );
  XOR U16475 ( .A(n16346), .B(n16345), .Z(n16348) );
  XNOR U16476 ( .A(n16347), .B(n16348), .Z(n16411) );
  XNOR U16477 ( .A(n16412), .B(n16411), .Z(n16413) );
  NANDN U16478 ( .A(n15949), .B(n15948), .Z(n15953) );
  OR U16479 ( .A(n15951), .B(n15950), .Z(n15952) );
  NAND U16480 ( .A(n15953), .B(n15952), .Z(n16414) );
  XNOR U16481 ( .A(n16413), .B(n16414), .Z(n16234) );
  XNOR U16482 ( .A(n16235), .B(n16234), .Z(n16237) );
  NANDN U16483 ( .A(n29499), .B(n15954), .Z(n15956) );
  XOR U16484 ( .A(a[80]), .B(b[7]), .Z(n16300) );
  NANDN U16485 ( .A(n29735), .B(n16300), .Z(n15955) );
  AND U16486 ( .A(n15956), .B(n15955), .Z(n16290) );
  NANDN U16487 ( .A(n37857), .B(n15957), .Z(n15959) );
  XOR U16488 ( .A(b[55]), .B(a[32]), .Z(n16303) );
  NANDN U16489 ( .A(n37911), .B(n16303), .Z(n15958) );
  AND U16490 ( .A(n15959), .B(n15958), .Z(n16289) );
  NANDN U16491 ( .A(n35611), .B(n15960), .Z(n15962) );
  XOR U16492 ( .A(b[35]), .B(a[52]), .Z(n16306) );
  NANDN U16493 ( .A(n35801), .B(n16306), .Z(n15961) );
  NAND U16494 ( .A(n15962), .B(n15961), .Z(n16288) );
  XOR U16495 ( .A(n16289), .B(n16288), .Z(n16291) );
  XOR U16496 ( .A(n16290), .B(n16291), .Z(n16352) );
  NANDN U16497 ( .A(n15964), .B(n15963), .Z(n15968) );
  NANDN U16498 ( .A(n15966), .B(n15965), .Z(n15967) );
  AND U16499 ( .A(n15968), .B(n15967), .Z(n16351) );
  XNOR U16500 ( .A(n16352), .B(n16351), .Z(n16353) );
  NANDN U16501 ( .A(n15970), .B(n15969), .Z(n15974) );
  OR U16502 ( .A(n15972), .B(n15971), .Z(n15973) );
  NAND U16503 ( .A(n15974), .B(n15973), .Z(n16354) );
  XNOR U16504 ( .A(n16353), .B(n16354), .Z(n16236) );
  XOR U16505 ( .A(n16237), .B(n16236), .Z(n16217) );
  NANDN U16506 ( .A(n15976), .B(n15975), .Z(n15980) );
  NANDN U16507 ( .A(n15978), .B(n15977), .Z(n15979) );
  AND U16508 ( .A(n15980), .B(n15979), .Z(n16231) );
  NAND U16509 ( .A(n15982), .B(n15981), .Z(n15986) );
  NAND U16510 ( .A(n15984), .B(n15983), .Z(n15985) );
  AND U16511 ( .A(n15986), .B(n15985), .Z(n16229) );
  NANDN U16512 ( .A(n33875), .B(n15987), .Z(n15989) );
  XOR U16513 ( .A(b[25]), .B(a[62]), .Z(n16264) );
  NANDN U16514 ( .A(n33994), .B(n16264), .Z(n15988) );
  AND U16515 ( .A(n15989), .B(n15988), .Z(n16434) );
  NANDN U16516 ( .A(n32013), .B(n15990), .Z(n15992) );
  XOR U16517 ( .A(b[17]), .B(a[70]), .Z(n16267) );
  NANDN U16518 ( .A(n32292), .B(n16267), .Z(n15991) );
  AND U16519 ( .A(n15992), .B(n15991), .Z(n16433) );
  NANDN U16520 ( .A(n31536), .B(n15993), .Z(n15995) );
  XOR U16521 ( .A(b[15]), .B(a[72]), .Z(n16270) );
  NANDN U16522 ( .A(n31925), .B(n16270), .Z(n15994) );
  NAND U16523 ( .A(n15995), .B(n15994), .Z(n16432) );
  XOR U16524 ( .A(n16433), .B(n16432), .Z(n16435) );
  XOR U16525 ( .A(n16434), .B(n16435), .Z(n16406) );
  NANDN U16526 ( .A(n37526), .B(n15996), .Z(n15998) );
  XOR U16527 ( .A(b[51]), .B(a[36]), .Z(n16273) );
  NANDN U16528 ( .A(n37605), .B(n16273), .Z(n15997) );
  AND U16529 ( .A(n15998), .B(n15997), .Z(n16458) );
  NANDN U16530 ( .A(n37705), .B(n15999), .Z(n16001) );
  XOR U16531 ( .A(b[53]), .B(a[34]), .Z(n16276) );
  NANDN U16532 ( .A(n37778), .B(n16276), .Z(n16000) );
  AND U16533 ( .A(n16001), .B(n16000), .Z(n16457) );
  NANDN U16534 ( .A(n36210), .B(n16002), .Z(n16004) );
  XOR U16535 ( .A(b[39]), .B(a[48]), .Z(n16279) );
  NANDN U16536 ( .A(n36347), .B(n16279), .Z(n16003) );
  NAND U16537 ( .A(n16004), .B(n16003), .Z(n16456) );
  XOR U16538 ( .A(n16457), .B(n16456), .Z(n16459) );
  XNOR U16539 ( .A(n16458), .B(n16459), .Z(n16405) );
  XNOR U16540 ( .A(n16406), .B(n16405), .Z(n16408) );
  NANDN U16541 ( .A(n16006), .B(n16005), .Z(n16010) );
  NANDN U16542 ( .A(n16008), .B(n16007), .Z(n16009) );
  AND U16543 ( .A(n16010), .B(n16009), .Z(n16407) );
  XOR U16544 ( .A(n16408), .B(n16407), .Z(n16255) );
  NANDN U16545 ( .A(n16012), .B(n16011), .Z(n16016) );
  OR U16546 ( .A(n16014), .B(n16013), .Z(n16015) );
  AND U16547 ( .A(n16016), .B(n16015), .Z(n16253) );
  NANDN U16548 ( .A(n16018), .B(n16017), .Z(n16022) );
  NANDN U16549 ( .A(n16020), .B(n16019), .Z(n16021) );
  NAND U16550 ( .A(n16022), .B(n16021), .Z(n16252) );
  XNOR U16551 ( .A(n16253), .B(n16252), .Z(n16254) );
  XNOR U16552 ( .A(n16255), .B(n16254), .Z(n16228) );
  XNOR U16553 ( .A(n16229), .B(n16228), .Z(n16230) );
  XNOR U16554 ( .A(n16231), .B(n16230), .Z(n16216) );
  XNOR U16555 ( .A(n16217), .B(n16216), .Z(n16218) );
  NANDN U16556 ( .A(n16024), .B(n16023), .Z(n16028) );
  NAND U16557 ( .A(n16026), .B(n16025), .Z(n16027) );
  NAND U16558 ( .A(n16028), .B(n16027), .Z(n16219) );
  XNOR U16559 ( .A(n16218), .B(n16219), .Z(n16468) );
  NAND U16560 ( .A(n16030), .B(n16029), .Z(n16034) );
  NANDN U16561 ( .A(n16032), .B(n16031), .Z(n16033) );
  NAND U16562 ( .A(n16034), .B(n16033), .Z(n16222) );
  NANDN U16563 ( .A(n16036), .B(n16035), .Z(n16040) );
  NAND U16564 ( .A(n16038), .B(n16037), .Z(n16039) );
  AND U16565 ( .A(n16040), .B(n16039), .Z(n16223) );
  XOR U16566 ( .A(n16222), .B(n16223), .Z(n16225) );
  NANDN U16567 ( .A(n16042), .B(n16041), .Z(n16046) );
  NANDN U16568 ( .A(n16044), .B(n16043), .Z(n16045) );
  NAND U16569 ( .A(n16046), .B(n16045), .Z(n16224) );
  XOR U16570 ( .A(n16225), .B(n16224), .Z(n16243) );
  NANDN U16571 ( .A(n16048), .B(n16047), .Z(n16052) );
  OR U16572 ( .A(n16050), .B(n16049), .Z(n16051) );
  AND U16573 ( .A(n16052), .B(n16051), .Z(n16364) );
  NANDN U16574 ( .A(n16054), .B(n16053), .Z(n16058) );
  NANDN U16575 ( .A(n16056), .B(n16055), .Z(n16057) );
  NAND U16576 ( .A(n16058), .B(n16057), .Z(n16363) );
  XNOR U16577 ( .A(n16364), .B(n16363), .Z(n16366) );
  NANDN U16578 ( .A(n16060), .B(n16059), .Z(n16064) );
  NANDN U16579 ( .A(n16062), .B(n16061), .Z(n16063) );
  AND U16580 ( .A(n16064), .B(n16063), .Z(n16261) );
  NAND U16581 ( .A(b[0]), .B(a[86]), .Z(n16065) );
  XNOR U16582 ( .A(b[1]), .B(n16065), .Z(n16067) );
  NANDN U16583 ( .A(b[0]), .B(a[85]), .Z(n16066) );
  NAND U16584 ( .A(n16067), .B(n16066), .Z(n16297) );
  NANDN U16585 ( .A(n38278), .B(n16068), .Z(n16070) );
  XOR U16586 ( .A(b[63]), .B(a[24]), .Z(n16387) );
  NANDN U16587 ( .A(n38279), .B(n16387), .Z(n16069) );
  AND U16588 ( .A(n16070), .B(n16069), .Z(n16295) );
  NANDN U16589 ( .A(n35260), .B(n16071), .Z(n16073) );
  XOR U16590 ( .A(b[33]), .B(a[54]), .Z(n16390) );
  NANDN U16591 ( .A(n35456), .B(n16390), .Z(n16072) );
  NAND U16592 ( .A(n16073), .B(n16072), .Z(n16294) );
  XNOR U16593 ( .A(n16295), .B(n16294), .Z(n16296) );
  XNOR U16594 ( .A(n16297), .B(n16296), .Z(n16258) );
  NANDN U16595 ( .A(n37974), .B(n16074), .Z(n16076) );
  XOR U16596 ( .A(b[57]), .B(a[30]), .Z(n16396) );
  NANDN U16597 ( .A(n38031), .B(n16396), .Z(n16075) );
  AND U16598 ( .A(n16076), .B(n16075), .Z(n16372) );
  NANDN U16599 ( .A(n38090), .B(n16077), .Z(n16079) );
  XOR U16600 ( .A(b[59]), .B(a[28]), .Z(n16399) );
  NANDN U16601 ( .A(n38130), .B(n16399), .Z(n16078) );
  AND U16602 ( .A(n16079), .B(n16078), .Z(n16370) );
  NANDN U16603 ( .A(n36480), .B(n16080), .Z(n16082) );
  XOR U16604 ( .A(b[41]), .B(a[46]), .Z(n16402) );
  NANDN U16605 ( .A(n36594), .B(n16402), .Z(n16081) );
  NAND U16606 ( .A(n16082), .B(n16081), .Z(n16369) );
  XNOR U16607 ( .A(n16370), .B(n16369), .Z(n16371) );
  XOR U16608 ( .A(n16372), .B(n16371), .Z(n16259) );
  XNOR U16609 ( .A(n16258), .B(n16259), .Z(n16260) );
  XNOR U16610 ( .A(n16261), .B(n16260), .Z(n16365) );
  XOR U16611 ( .A(n16366), .B(n16365), .Z(n16247) );
  NANDN U16612 ( .A(n16084), .B(n16083), .Z(n16088) );
  NAND U16613 ( .A(n16086), .B(n16085), .Z(n16087) );
  NAND U16614 ( .A(n16088), .B(n16087), .Z(n16246) );
  XNOR U16615 ( .A(n16247), .B(n16246), .Z(n16249) );
  NANDN U16616 ( .A(n16090), .B(n16089), .Z(n16094) );
  NANDN U16617 ( .A(n16092), .B(n16091), .Z(n16093) );
  AND U16618 ( .A(n16094), .B(n16093), .Z(n16465) );
  NANDN U16619 ( .A(n32996), .B(n16095), .Z(n16097) );
  XOR U16620 ( .A(b[21]), .B(a[66]), .Z(n16417) );
  NANDN U16621 ( .A(n33271), .B(n16417), .Z(n16096) );
  AND U16622 ( .A(n16097), .B(n16096), .Z(n16383) );
  NANDN U16623 ( .A(n33866), .B(n16098), .Z(n16100) );
  XOR U16624 ( .A(b[23]), .B(a[64]), .Z(n16420) );
  NANDN U16625 ( .A(n33644), .B(n16420), .Z(n16099) );
  AND U16626 ( .A(n16100), .B(n16099), .Z(n16382) );
  NANDN U16627 ( .A(n32483), .B(n16101), .Z(n16103) );
  XOR U16628 ( .A(b[19]), .B(a[68]), .Z(n16423) );
  NANDN U16629 ( .A(n32823), .B(n16423), .Z(n16102) );
  NAND U16630 ( .A(n16103), .B(n16102), .Z(n16381) );
  XOR U16631 ( .A(n16382), .B(n16381), .Z(n16384) );
  XOR U16632 ( .A(n16383), .B(n16384), .Z(n16322) );
  NANDN U16633 ( .A(n34909), .B(n16104), .Z(n16106) );
  XOR U16634 ( .A(b[31]), .B(a[56]), .Z(n16426) );
  NANDN U16635 ( .A(n35145), .B(n16426), .Z(n16105) );
  AND U16636 ( .A(n16106), .B(n16105), .Z(n16311) );
  NANDN U16637 ( .A(n38247), .B(n16107), .Z(n16109) );
  XOR U16638 ( .A(b[61]), .B(a[26]), .Z(n16429) );
  NANDN U16639 ( .A(n38248), .B(n16429), .Z(n16108) );
  AND U16640 ( .A(n16109), .B(n16108), .Z(n16310) );
  AND U16641 ( .A(b[63]), .B(a[22]), .Z(n16309) );
  XOR U16642 ( .A(n16310), .B(n16309), .Z(n16312) );
  XNOR U16643 ( .A(n16311), .B(n16312), .Z(n16321) );
  XNOR U16644 ( .A(n16322), .B(n16321), .Z(n16323) );
  NANDN U16645 ( .A(n16111), .B(n16110), .Z(n16115) );
  OR U16646 ( .A(n16113), .B(n16112), .Z(n16114) );
  NAND U16647 ( .A(n16115), .B(n16114), .Z(n16324) );
  XNOR U16648 ( .A(n16323), .B(n16324), .Z(n16462) );
  NANDN U16649 ( .A(n34223), .B(n16116), .Z(n16118) );
  XOR U16650 ( .A(b[27]), .B(a[60]), .Z(n16438) );
  NANDN U16651 ( .A(n34458), .B(n16438), .Z(n16117) );
  AND U16652 ( .A(n16118), .B(n16117), .Z(n16284) );
  NANDN U16653 ( .A(n34634), .B(n16119), .Z(n16121) );
  XOR U16654 ( .A(b[29]), .B(a[58]), .Z(n16441) );
  NANDN U16655 ( .A(n34722), .B(n16441), .Z(n16120) );
  AND U16656 ( .A(n16121), .B(n16120), .Z(n16283) );
  NANDN U16657 ( .A(n31055), .B(n16122), .Z(n16124) );
  XOR U16658 ( .A(b[13]), .B(a[74]), .Z(n16444) );
  NANDN U16659 ( .A(n31293), .B(n16444), .Z(n16123) );
  NAND U16660 ( .A(n16124), .B(n16123), .Z(n16282) );
  XOR U16661 ( .A(n16283), .B(n16282), .Z(n16285) );
  XOR U16662 ( .A(n16284), .B(n16285), .Z(n16358) );
  NANDN U16663 ( .A(n28889), .B(n16125), .Z(n16127) );
  XOR U16664 ( .A(a[82]), .B(b[5]), .Z(n16447) );
  NANDN U16665 ( .A(n29138), .B(n16447), .Z(n16126) );
  AND U16666 ( .A(n16127), .B(n16126), .Z(n16377) );
  NANDN U16667 ( .A(n209), .B(n16128), .Z(n16130) );
  XOR U16668 ( .A(a[84]), .B(b[3]), .Z(n16450) );
  NANDN U16669 ( .A(n28941), .B(n16450), .Z(n16129) );
  AND U16670 ( .A(n16130), .B(n16129), .Z(n16376) );
  NANDN U16671 ( .A(n35936), .B(n16131), .Z(n16133) );
  XOR U16672 ( .A(b[37]), .B(a[50]), .Z(n16453) );
  NANDN U16673 ( .A(n36047), .B(n16453), .Z(n16132) );
  NAND U16674 ( .A(n16133), .B(n16132), .Z(n16375) );
  XOR U16675 ( .A(n16376), .B(n16375), .Z(n16378) );
  XNOR U16676 ( .A(n16377), .B(n16378), .Z(n16357) );
  XNOR U16677 ( .A(n16358), .B(n16357), .Z(n16359) );
  NANDN U16678 ( .A(n16135), .B(n16134), .Z(n16139) );
  OR U16679 ( .A(n16137), .B(n16136), .Z(n16138) );
  NAND U16680 ( .A(n16139), .B(n16138), .Z(n16360) );
  XOR U16681 ( .A(n16359), .B(n16360), .Z(n16463) );
  XNOR U16682 ( .A(n16462), .B(n16463), .Z(n16464) );
  XNOR U16683 ( .A(n16465), .B(n16464), .Z(n16248) );
  XOR U16684 ( .A(n16249), .B(n16248), .Z(n16241) );
  XNOR U16685 ( .A(n16241), .B(n16240), .Z(n16242) );
  XOR U16686 ( .A(n16243), .B(n16242), .Z(n16469) );
  XOR U16687 ( .A(n16468), .B(n16469), .Z(n16471) );
  XOR U16688 ( .A(n16470), .B(n16471), .Z(n16212) );
  NAND U16689 ( .A(n16145), .B(n16144), .Z(n16149) );
  NAND U16690 ( .A(n16147), .B(n16146), .Z(n16148) );
  AND U16691 ( .A(n16149), .B(n16148), .Z(n16477) );
  NANDN U16692 ( .A(n16151), .B(n16150), .Z(n16155) );
  OR U16693 ( .A(n16153), .B(n16152), .Z(n16154) );
  AND U16694 ( .A(n16155), .B(n16154), .Z(n16475) );
  NANDN U16695 ( .A(n16157), .B(n16156), .Z(n16161) );
  NANDN U16696 ( .A(n16159), .B(n16158), .Z(n16160) );
  AND U16697 ( .A(n16161), .B(n16160), .Z(n16474) );
  XNOR U16698 ( .A(n16475), .B(n16474), .Z(n16476) );
  XOR U16699 ( .A(n16477), .B(n16476), .Z(n16211) );
  NANDN U16700 ( .A(n16163), .B(n16162), .Z(n16167) );
  OR U16701 ( .A(n16165), .B(n16164), .Z(n16166) );
  NAND U16702 ( .A(n16167), .B(n16166), .Z(n16210) );
  XOR U16703 ( .A(n16211), .B(n16210), .Z(n16213) );
  XOR U16704 ( .A(n16212), .B(n16213), .Z(n16206) );
  NANDN U16705 ( .A(n16169), .B(n16168), .Z(n16173) );
  NANDN U16706 ( .A(n16171), .B(n16170), .Z(n16172) );
  AND U16707 ( .A(n16173), .B(n16172), .Z(n16205) );
  NANDN U16708 ( .A(n16175), .B(n16174), .Z(n16179) );
  OR U16709 ( .A(n16177), .B(n16176), .Z(n16178) );
  AND U16710 ( .A(n16179), .B(n16178), .Z(n16204) );
  XOR U16711 ( .A(n16205), .B(n16204), .Z(n16207) );
  XOR U16712 ( .A(n16206), .B(n16207), .Z(n16199) );
  NANDN U16713 ( .A(n16181), .B(n16180), .Z(n16185) );
  NANDN U16714 ( .A(n16183), .B(n16182), .Z(n16184) );
  AND U16715 ( .A(n16185), .B(n16184), .Z(n16198) );
  XNOR U16716 ( .A(n16199), .B(n16198), .Z(n16200) );
  NANDN U16717 ( .A(n16187), .B(n16186), .Z(n16191) );
  NAND U16718 ( .A(n16189), .B(n16188), .Z(n16190) );
  NAND U16719 ( .A(n16191), .B(n16190), .Z(n16201) );
  XNOR U16720 ( .A(n16200), .B(n16201), .Z(n16192) );
  XNOR U16721 ( .A(n16193), .B(n16192), .Z(n16194) );
  XNOR U16722 ( .A(n16195), .B(n16194), .Z(n16480) );
  XNOR U16723 ( .A(sreg[150]), .B(n16480), .Z(n16481) );
  XNOR U16724 ( .A(n16482), .B(n16481), .Z(c[150]) );
  NANDN U16725 ( .A(n16193), .B(n16192), .Z(n16197) );
  NANDN U16726 ( .A(n16195), .B(n16194), .Z(n16196) );
  AND U16727 ( .A(n16197), .B(n16196), .Z(n16488) );
  NANDN U16728 ( .A(n16199), .B(n16198), .Z(n16203) );
  NANDN U16729 ( .A(n16201), .B(n16200), .Z(n16202) );
  AND U16730 ( .A(n16203), .B(n16202), .Z(n16486) );
  NANDN U16731 ( .A(n16205), .B(n16204), .Z(n16209) );
  OR U16732 ( .A(n16207), .B(n16206), .Z(n16208) );
  AND U16733 ( .A(n16209), .B(n16208), .Z(n16769) );
  NANDN U16734 ( .A(n16211), .B(n16210), .Z(n16215) );
  OR U16735 ( .A(n16213), .B(n16212), .Z(n16214) );
  AND U16736 ( .A(n16215), .B(n16214), .Z(n16767) );
  NANDN U16737 ( .A(n16217), .B(n16216), .Z(n16221) );
  NANDN U16738 ( .A(n16219), .B(n16218), .Z(n16220) );
  AND U16739 ( .A(n16221), .B(n16220), .Z(n16756) );
  NAND U16740 ( .A(n16223), .B(n16222), .Z(n16227) );
  NAND U16741 ( .A(n16225), .B(n16224), .Z(n16226) );
  AND U16742 ( .A(n16227), .B(n16226), .Z(n16751) );
  NANDN U16743 ( .A(n16229), .B(n16228), .Z(n16233) );
  NANDN U16744 ( .A(n16231), .B(n16230), .Z(n16232) );
  AND U16745 ( .A(n16233), .B(n16232), .Z(n16750) );
  NANDN U16746 ( .A(n16235), .B(n16234), .Z(n16239) );
  NAND U16747 ( .A(n16237), .B(n16236), .Z(n16238) );
  AND U16748 ( .A(n16239), .B(n16238), .Z(n16749) );
  XOR U16749 ( .A(n16750), .B(n16749), .Z(n16752) );
  XNOR U16750 ( .A(n16751), .B(n16752), .Z(n16755) );
  XNOR U16751 ( .A(n16756), .B(n16755), .Z(n16757) );
  NANDN U16752 ( .A(n16241), .B(n16240), .Z(n16245) );
  NANDN U16753 ( .A(n16243), .B(n16242), .Z(n16244) );
  AND U16754 ( .A(n16245), .B(n16244), .Z(n16746) );
  NANDN U16755 ( .A(n16247), .B(n16246), .Z(n16251) );
  NAND U16756 ( .A(n16249), .B(n16248), .Z(n16250) );
  AND U16757 ( .A(n16251), .B(n16250), .Z(n16511) );
  NANDN U16758 ( .A(n16253), .B(n16252), .Z(n16257) );
  NANDN U16759 ( .A(n16255), .B(n16254), .Z(n16256) );
  AND U16760 ( .A(n16257), .B(n16256), .Z(n16505) );
  NANDN U16761 ( .A(n16259), .B(n16258), .Z(n16263) );
  NANDN U16762 ( .A(n16261), .B(n16260), .Z(n16262) );
  AND U16763 ( .A(n16263), .B(n16262), .Z(n16504) );
  NANDN U16764 ( .A(n33875), .B(n16264), .Z(n16266) );
  XOR U16765 ( .A(b[25]), .B(a[63]), .Z(n16584) );
  NANDN U16766 ( .A(n33994), .B(n16584), .Z(n16265) );
  AND U16767 ( .A(n16266), .B(n16265), .Z(n16673) );
  NANDN U16768 ( .A(n32013), .B(n16267), .Z(n16269) );
  XOR U16769 ( .A(b[17]), .B(a[71]), .Z(n16587) );
  NANDN U16770 ( .A(n32292), .B(n16587), .Z(n16268) );
  AND U16771 ( .A(n16269), .B(n16268), .Z(n16672) );
  NANDN U16772 ( .A(n31536), .B(n16270), .Z(n16272) );
  XOR U16773 ( .A(b[15]), .B(a[73]), .Z(n16590) );
  NANDN U16774 ( .A(n31925), .B(n16590), .Z(n16271) );
  NAND U16775 ( .A(n16272), .B(n16271), .Z(n16671) );
  XOR U16776 ( .A(n16672), .B(n16671), .Z(n16674) );
  XOR U16777 ( .A(n16673), .B(n16674), .Z(n16702) );
  NANDN U16778 ( .A(n37526), .B(n16273), .Z(n16275) );
  XOR U16779 ( .A(b[51]), .B(a[37]), .Z(n16593) );
  NANDN U16780 ( .A(n37605), .B(n16593), .Z(n16274) );
  AND U16781 ( .A(n16275), .B(n16274), .Z(n16697) );
  NANDN U16782 ( .A(n37705), .B(n16276), .Z(n16278) );
  XOR U16783 ( .A(b[53]), .B(a[35]), .Z(n16596) );
  NANDN U16784 ( .A(n37778), .B(n16596), .Z(n16277) );
  AND U16785 ( .A(n16278), .B(n16277), .Z(n16696) );
  NANDN U16786 ( .A(n36210), .B(n16279), .Z(n16281) );
  XOR U16787 ( .A(b[39]), .B(a[49]), .Z(n16599) );
  NANDN U16788 ( .A(n36347), .B(n16599), .Z(n16280) );
  NAND U16789 ( .A(n16281), .B(n16280), .Z(n16695) );
  XOR U16790 ( .A(n16696), .B(n16695), .Z(n16698) );
  XNOR U16791 ( .A(n16697), .B(n16698), .Z(n16701) );
  XNOR U16792 ( .A(n16702), .B(n16701), .Z(n16704) );
  NANDN U16793 ( .A(n16283), .B(n16282), .Z(n16287) );
  OR U16794 ( .A(n16285), .B(n16284), .Z(n16286) );
  AND U16795 ( .A(n16287), .B(n16286), .Z(n16703) );
  XOR U16796 ( .A(n16704), .B(n16703), .Z(n16575) );
  NANDN U16797 ( .A(n16289), .B(n16288), .Z(n16293) );
  OR U16798 ( .A(n16291), .B(n16290), .Z(n16292) );
  AND U16799 ( .A(n16293), .B(n16292), .Z(n16573) );
  NANDN U16800 ( .A(n16295), .B(n16294), .Z(n16299) );
  NANDN U16801 ( .A(n16297), .B(n16296), .Z(n16298) );
  NAND U16802 ( .A(n16299), .B(n16298), .Z(n16572) );
  XNOR U16803 ( .A(n16573), .B(n16572), .Z(n16574) );
  XNOR U16804 ( .A(n16575), .B(n16574), .Z(n16503) );
  XOR U16805 ( .A(n16504), .B(n16503), .Z(n16506) );
  XOR U16806 ( .A(n16505), .B(n16506), .Z(n16510) );
  NANDN U16807 ( .A(n29499), .B(n16300), .Z(n16302) );
  XOR U16808 ( .A(a[81]), .B(b[7]), .Z(n16551) );
  NANDN U16809 ( .A(n29735), .B(n16551), .Z(n16301) );
  AND U16810 ( .A(n16302), .B(n16301), .Z(n16610) );
  NANDN U16811 ( .A(n37857), .B(n16303), .Z(n16305) );
  XOR U16812 ( .A(b[55]), .B(a[33]), .Z(n16554) );
  NANDN U16813 ( .A(n37911), .B(n16554), .Z(n16304) );
  AND U16814 ( .A(n16305), .B(n16304), .Z(n16609) );
  NANDN U16815 ( .A(n35611), .B(n16306), .Z(n16308) );
  XOR U16816 ( .A(b[35]), .B(a[53]), .Z(n16557) );
  NANDN U16817 ( .A(n35801), .B(n16557), .Z(n16307) );
  NAND U16818 ( .A(n16308), .B(n16307), .Z(n16608) );
  XOR U16819 ( .A(n16609), .B(n16608), .Z(n16611) );
  XOR U16820 ( .A(n16610), .B(n16611), .Z(n16627) );
  NANDN U16821 ( .A(n16310), .B(n16309), .Z(n16314) );
  OR U16822 ( .A(n16312), .B(n16311), .Z(n16313) );
  AND U16823 ( .A(n16314), .B(n16313), .Z(n16626) );
  XNOR U16824 ( .A(n16627), .B(n16626), .Z(n16628) );
  NANDN U16825 ( .A(n16316), .B(n16315), .Z(n16320) );
  OR U16826 ( .A(n16318), .B(n16317), .Z(n16319) );
  NAND U16827 ( .A(n16320), .B(n16319), .Z(n16629) );
  XNOR U16828 ( .A(n16628), .B(n16629), .Z(n16499) );
  NANDN U16829 ( .A(n16322), .B(n16321), .Z(n16326) );
  NANDN U16830 ( .A(n16324), .B(n16323), .Z(n16325) );
  AND U16831 ( .A(n16326), .B(n16325), .Z(n16498) );
  NANDN U16832 ( .A(n211), .B(n16327), .Z(n16329) );
  XOR U16833 ( .A(b[47]), .B(a[41]), .Z(n16527) );
  NANDN U16834 ( .A(n37172), .B(n16527), .Z(n16328) );
  AND U16835 ( .A(n16329), .B(n16328), .Z(n16568) );
  NANDN U16836 ( .A(n210), .B(n16330), .Z(n16332) );
  XOR U16837 ( .A(a[79]), .B(b[9]), .Z(n16530) );
  NANDN U16838 ( .A(n30267), .B(n16530), .Z(n16331) );
  AND U16839 ( .A(n16332), .B(n16331), .Z(n16567) );
  NANDN U16840 ( .A(n212), .B(n16333), .Z(n16335) );
  XOR U16841 ( .A(b[49]), .B(a[39]), .Z(n16533) );
  NANDN U16842 ( .A(n37432), .B(n16533), .Z(n16334) );
  NAND U16843 ( .A(n16335), .B(n16334), .Z(n16566) );
  XOR U16844 ( .A(n16567), .B(n16566), .Z(n16569) );
  XOR U16845 ( .A(n16568), .B(n16569), .Z(n16651) );
  NANDN U16846 ( .A(n36742), .B(n16336), .Z(n16338) );
  XOR U16847 ( .A(b[43]), .B(a[45]), .Z(n16536) );
  NANDN U16848 ( .A(n36891), .B(n16536), .Z(n16337) );
  AND U16849 ( .A(n16338), .B(n16337), .Z(n16547) );
  NANDN U16850 ( .A(n36991), .B(n16339), .Z(n16341) );
  XOR U16851 ( .A(b[45]), .B(a[43]), .Z(n16539) );
  NANDN U16852 ( .A(n37083), .B(n16539), .Z(n16340) );
  AND U16853 ( .A(n16341), .B(n16340), .Z(n16546) );
  NANDN U16854 ( .A(n30482), .B(n16342), .Z(n16344) );
  XOR U16855 ( .A(a[77]), .B(b[11]), .Z(n16542) );
  NANDN U16856 ( .A(n30891), .B(n16542), .Z(n16343) );
  NAND U16857 ( .A(n16344), .B(n16343), .Z(n16545) );
  XOR U16858 ( .A(n16546), .B(n16545), .Z(n16548) );
  XNOR U16859 ( .A(n16547), .B(n16548), .Z(n16650) );
  XNOR U16860 ( .A(n16651), .B(n16650), .Z(n16652) );
  NANDN U16861 ( .A(n16346), .B(n16345), .Z(n16350) );
  OR U16862 ( .A(n16348), .B(n16347), .Z(n16349) );
  NAND U16863 ( .A(n16350), .B(n16349), .Z(n16653) );
  XNOR U16864 ( .A(n16652), .B(n16653), .Z(n16497) );
  XOR U16865 ( .A(n16498), .B(n16497), .Z(n16500) );
  XNOR U16866 ( .A(n16499), .B(n16500), .Z(n16509) );
  XOR U16867 ( .A(n16510), .B(n16509), .Z(n16512) );
  XOR U16868 ( .A(n16511), .B(n16512), .Z(n16744) );
  NANDN U16869 ( .A(n16352), .B(n16351), .Z(n16356) );
  NANDN U16870 ( .A(n16354), .B(n16353), .Z(n16355) );
  AND U16871 ( .A(n16356), .B(n16355), .Z(n16493) );
  NANDN U16872 ( .A(n16358), .B(n16357), .Z(n16362) );
  NANDN U16873 ( .A(n16360), .B(n16359), .Z(n16361) );
  AND U16874 ( .A(n16362), .B(n16361), .Z(n16492) );
  NANDN U16875 ( .A(n16364), .B(n16363), .Z(n16368) );
  NAND U16876 ( .A(n16366), .B(n16365), .Z(n16367) );
  AND U16877 ( .A(n16368), .B(n16367), .Z(n16491) );
  XOR U16878 ( .A(n16492), .B(n16491), .Z(n16494) );
  XOR U16879 ( .A(n16493), .B(n16494), .Z(n16518) );
  NANDN U16880 ( .A(n16370), .B(n16369), .Z(n16374) );
  NANDN U16881 ( .A(n16372), .B(n16371), .Z(n16373) );
  AND U16882 ( .A(n16374), .B(n16373), .Z(n16639) );
  NANDN U16883 ( .A(n16376), .B(n16375), .Z(n16380) );
  OR U16884 ( .A(n16378), .B(n16377), .Z(n16379) );
  NAND U16885 ( .A(n16380), .B(n16379), .Z(n16638) );
  XNOR U16886 ( .A(n16639), .B(n16638), .Z(n16641) );
  NANDN U16887 ( .A(n16382), .B(n16381), .Z(n16386) );
  OR U16888 ( .A(n16384), .B(n16383), .Z(n16385) );
  AND U16889 ( .A(n16386), .B(n16385), .Z(n16581) );
  NANDN U16890 ( .A(n38278), .B(n16387), .Z(n16389) );
  XOR U16891 ( .A(b[63]), .B(a[25]), .Z(n16725) );
  NANDN U16892 ( .A(n38279), .B(n16725), .Z(n16388) );
  AND U16893 ( .A(n16389), .B(n16388), .Z(n16615) );
  NANDN U16894 ( .A(n35260), .B(n16390), .Z(n16392) );
  XOR U16895 ( .A(b[33]), .B(a[55]), .Z(n16728) );
  NANDN U16896 ( .A(n35456), .B(n16728), .Z(n16391) );
  NAND U16897 ( .A(n16392), .B(n16391), .Z(n16614) );
  XNOR U16898 ( .A(n16615), .B(n16614), .Z(n16616) );
  NAND U16899 ( .A(b[0]), .B(a[87]), .Z(n16393) );
  XNOR U16900 ( .A(b[1]), .B(n16393), .Z(n16395) );
  NANDN U16901 ( .A(b[0]), .B(a[86]), .Z(n16394) );
  NAND U16902 ( .A(n16395), .B(n16394), .Z(n16617) );
  XNOR U16903 ( .A(n16616), .B(n16617), .Z(n16578) );
  NANDN U16904 ( .A(n37974), .B(n16396), .Z(n16398) );
  XOR U16905 ( .A(b[57]), .B(a[31]), .Z(n16734) );
  NANDN U16906 ( .A(n38031), .B(n16734), .Z(n16397) );
  AND U16907 ( .A(n16398), .B(n16397), .Z(n16710) );
  NANDN U16908 ( .A(n38090), .B(n16399), .Z(n16401) );
  XOR U16909 ( .A(b[59]), .B(a[29]), .Z(n16737) );
  NANDN U16910 ( .A(n38130), .B(n16737), .Z(n16400) );
  AND U16911 ( .A(n16401), .B(n16400), .Z(n16708) );
  NANDN U16912 ( .A(n36480), .B(n16402), .Z(n16404) );
  XOR U16913 ( .A(b[41]), .B(a[47]), .Z(n16740) );
  NANDN U16914 ( .A(n36594), .B(n16740), .Z(n16403) );
  NAND U16915 ( .A(n16404), .B(n16403), .Z(n16707) );
  XNOR U16916 ( .A(n16708), .B(n16707), .Z(n16709) );
  XOR U16917 ( .A(n16710), .B(n16709), .Z(n16579) );
  XNOR U16918 ( .A(n16578), .B(n16579), .Z(n16580) );
  XNOR U16919 ( .A(n16581), .B(n16580), .Z(n16640) );
  XOR U16920 ( .A(n16641), .B(n16640), .Z(n16621) );
  NANDN U16921 ( .A(n16406), .B(n16405), .Z(n16410) );
  NAND U16922 ( .A(n16408), .B(n16407), .Z(n16409) );
  NAND U16923 ( .A(n16410), .B(n16409), .Z(n16620) );
  XNOR U16924 ( .A(n16621), .B(n16620), .Z(n16623) );
  NANDN U16925 ( .A(n16412), .B(n16411), .Z(n16416) );
  NANDN U16926 ( .A(n16414), .B(n16413), .Z(n16415) );
  AND U16927 ( .A(n16416), .B(n16415), .Z(n16647) );
  NANDN U16928 ( .A(n32996), .B(n16417), .Z(n16419) );
  XOR U16929 ( .A(b[21]), .B(a[67]), .Z(n16656) );
  NANDN U16930 ( .A(n33271), .B(n16656), .Z(n16418) );
  AND U16931 ( .A(n16419), .B(n16418), .Z(n16721) );
  NANDN U16932 ( .A(n33866), .B(n16420), .Z(n16422) );
  XOR U16933 ( .A(b[23]), .B(a[65]), .Z(n16659) );
  NANDN U16934 ( .A(n33644), .B(n16659), .Z(n16421) );
  AND U16935 ( .A(n16422), .B(n16421), .Z(n16720) );
  NANDN U16936 ( .A(n32483), .B(n16423), .Z(n16425) );
  XOR U16937 ( .A(b[19]), .B(a[69]), .Z(n16662) );
  NANDN U16938 ( .A(n32823), .B(n16662), .Z(n16424) );
  NAND U16939 ( .A(n16425), .B(n16424), .Z(n16719) );
  XOR U16940 ( .A(n16720), .B(n16719), .Z(n16722) );
  XOR U16941 ( .A(n16721), .B(n16722), .Z(n16522) );
  NANDN U16942 ( .A(n34909), .B(n16426), .Z(n16428) );
  XOR U16943 ( .A(b[31]), .B(a[57]), .Z(n16665) );
  NANDN U16944 ( .A(n35145), .B(n16665), .Z(n16427) );
  AND U16945 ( .A(n16428), .B(n16427), .Z(n16562) );
  NANDN U16946 ( .A(n38247), .B(n16429), .Z(n16431) );
  XOR U16947 ( .A(b[61]), .B(a[27]), .Z(n16668) );
  NANDN U16948 ( .A(n38248), .B(n16668), .Z(n16430) );
  AND U16949 ( .A(n16431), .B(n16430), .Z(n16561) );
  AND U16950 ( .A(b[63]), .B(a[23]), .Z(n16560) );
  XOR U16951 ( .A(n16561), .B(n16560), .Z(n16563) );
  XNOR U16952 ( .A(n16562), .B(n16563), .Z(n16521) );
  XNOR U16953 ( .A(n16522), .B(n16521), .Z(n16523) );
  NANDN U16954 ( .A(n16433), .B(n16432), .Z(n16437) );
  OR U16955 ( .A(n16435), .B(n16434), .Z(n16436) );
  NAND U16956 ( .A(n16437), .B(n16436), .Z(n16524) );
  XNOR U16957 ( .A(n16523), .B(n16524), .Z(n16644) );
  NANDN U16958 ( .A(n34223), .B(n16438), .Z(n16440) );
  XOR U16959 ( .A(b[27]), .B(a[61]), .Z(n16677) );
  NANDN U16960 ( .A(n34458), .B(n16677), .Z(n16439) );
  AND U16961 ( .A(n16440), .B(n16439), .Z(n16604) );
  NANDN U16962 ( .A(n34634), .B(n16441), .Z(n16443) );
  XOR U16963 ( .A(b[29]), .B(a[59]), .Z(n16680) );
  NANDN U16964 ( .A(n34722), .B(n16680), .Z(n16442) );
  AND U16965 ( .A(n16443), .B(n16442), .Z(n16603) );
  NANDN U16966 ( .A(n31055), .B(n16444), .Z(n16446) );
  XOR U16967 ( .A(b[13]), .B(a[75]), .Z(n16683) );
  NANDN U16968 ( .A(n31293), .B(n16683), .Z(n16445) );
  NAND U16969 ( .A(n16446), .B(n16445), .Z(n16602) );
  XOR U16970 ( .A(n16603), .B(n16602), .Z(n16605) );
  XOR U16971 ( .A(n16604), .B(n16605), .Z(n16633) );
  NANDN U16972 ( .A(n28889), .B(n16447), .Z(n16449) );
  XOR U16973 ( .A(a[83]), .B(b[5]), .Z(n16686) );
  NANDN U16974 ( .A(n29138), .B(n16686), .Z(n16448) );
  AND U16975 ( .A(n16449), .B(n16448), .Z(n16715) );
  NANDN U16976 ( .A(n209), .B(n16450), .Z(n16452) );
  XOR U16977 ( .A(a[85]), .B(b[3]), .Z(n16689) );
  NANDN U16978 ( .A(n28941), .B(n16689), .Z(n16451) );
  AND U16979 ( .A(n16452), .B(n16451), .Z(n16714) );
  NANDN U16980 ( .A(n35936), .B(n16453), .Z(n16455) );
  XOR U16981 ( .A(b[37]), .B(a[51]), .Z(n16692) );
  NANDN U16982 ( .A(n36047), .B(n16692), .Z(n16454) );
  NAND U16983 ( .A(n16455), .B(n16454), .Z(n16713) );
  XOR U16984 ( .A(n16714), .B(n16713), .Z(n16716) );
  XNOR U16985 ( .A(n16715), .B(n16716), .Z(n16632) );
  XNOR U16986 ( .A(n16633), .B(n16632), .Z(n16634) );
  NANDN U16987 ( .A(n16457), .B(n16456), .Z(n16461) );
  OR U16988 ( .A(n16459), .B(n16458), .Z(n16460) );
  NAND U16989 ( .A(n16461), .B(n16460), .Z(n16635) );
  XOR U16990 ( .A(n16634), .B(n16635), .Z(n16645) );
  XNOR U16991 ( .A(n16644), .B(n16645), .Z(n16646) );
  XNOR U16992 ( .A(n16647), .B(n16646), .Z(n16622) );
  XOR U16993 ( .A(n16623), .B(n16622), .Z(n16516) );
  NANDN U16994 ( .A(n16463), .B(n16462), .Z(n16467) );
  NANDN U16995 ( .A(n16465), .B(n16464), .Z(n16466) );
  AND U16996 ( .A(n16467), .B(n16466), .Z(n16515) );
  XNOR U16997 ( .A(n16516), .B(n16515), .Z(n16517) );
  XNOR U16998 ( .A(n16518), .B(n16517), .Z(n16743) );
  XNOR U16999 ( .A(n16744), .B(n16743), .Z(n16745) );
  XOR U17000 ( .A(n16746), .B(n16745), .Z(n16758) );
  XNOR U17001 ( .A(n16757), .B(n16758), .Z(n16763) );
  NANDN U17002 ( .A(n16469), .B(n16468), .Z(n16473) );
  OR U17003 ( .A(n16471), .B(n16470), .Z(n16472) );
  AND U17004 ( .A(n16473), .B(n16472), .Z(n16762) );
  NANDN U17005 ( .A(n16475), .B(n16474), .Z(n16479) );
  NAND U17006 ( .A(n16477), .B(n16476), .Z(n16478) );
  NAND U17007 ( .A(n16479), .B(n16478), .Z(n16761) );
  XOR U17008 ( .A(n16762), .B(n16761), .Z(n16764) );
  XOR U17009 ( .A(n16763), .B(n16764), .Z(n16768) );
  XOR U17010 ( .A(n16767), .B(n16768), .Z(n16770) );
  XNOR U17011 ( .A(n16769), .B(n16770), .Z(n16485) );
  XNOR U17012 ( .A(n16486), .B(n16485), .Z(n16487) );
  XNOR U17013 ( .A(n16488), .B(n16487), .Z(n16773) );
  XNOR U17014 ( .A(sreg[151]), .B(n16773), .Z(n16775) );
  NANDN U17015 ( .A(sreg[150]), .B(n16480), .Z(n16484) );
  NAND U17016 ( .A(n16482), .B(n16481), .Z(n16483) );
  NAND U17017 ( .A(n16484), .B(n16483), .Z(n16774) );
  XNOR U17018 ( .A(n16775), .B(n16774), .Z(c[151]) );
  NANDN U17019 ( .A(n16486), .B(n16485), .Z(n16490) );
  NANDN U17020 ( .A(n16488), .B(n16487), .Z(n16489) );
  AND U17021 ( .A(n16490), .B(n16489), .Z(n16781) );
  NANDN U17022 ( .A(n16492), .B(n16491), .Z(n16496) );
  OR U17023 ( .A(n16494), .B(n16493), .Z(n16495) );
  AND U17024 ( .A(n16496), .B(n16495), .Z(n17050) );
  NANDN U17025 ( .A(n16498), .B(n16497), .Z(n16502) );
  NANDN U17026 ( .A(n16500), .B(n16499), .Z(n16501) );
  AND U17027 ( .A(n16502), .B(n16501), .Z(n17049) );
  NANDN U17028 ( .A(n16504), .B(n16503), .Z(n16508) );
  OR U17029 ( .A(n16506), .B(n16505), .Z(n16507) );
  AND U17030 ( .A(n16508), .B(n16507), .Z(n17048) );
  XOR U17031 ( .A(n17049), .B(n17048), .Z(n17051) );
  XOR U17032 ( .A(n17050), .B(n17051), .Z(n17055) );
  NANDN U17033 ( .A(n16510), .B(n16509), .Z(n16514) );
  OR U17034 ( .A(n16512), .B(n16511), .Z(n16513) );
  AND U17035 ( .A(n16514), .B(n16513), .Z(n17054) );
  XNOR U17036 ( .A(n17055), .B(n17054), .Z(n17056) );
  NANDN U17037 ( .A(n16516), .B(n16515), .Z(n16520) );
  NANDN U17038 ( .A(n16518), .B(n16517), .Z(n16519) );
  AND U17039 ( .A(n16520), .B(n16519), .Z(n17045) );
  NANDN U17040 ( .A(n16522), .B(n16521), .Z(n16526) );
  NANDN U17041 ( .A(n16524), .B(n16523), .Z(n16525) );
  AND U17042 ( .A(n16526), .B(n16525), .Z(n17031) );
  NANDN U17043 ( .A(n211), .B(n16527), .Z(n16529) );
  XOR U17044 ( .A(b[47]), .B(a[42]), .Z(n16850) );
  NANDN U17045 ( .A(n37172), .B(n16850), .Z(n16528) );
  AND U17046 ( .A(n16529), .B(n16528), .Z(n16891) );
  NANDN U17047 ( .A(n210), .B(n16530), .Z(n16532) );
  XOR U17048 ( .A(a[80]), .B(b[9]), .Z(n16853) );
  NANDN U17049 ( .A(n30267), .B(n16853), .Z(n16531) );
  AND U17050 ( .A(n16532), .B(n16531), .Z(n16890) );
  NANDN U17051 ( .A(n212), .B(n16533), .Z(n16535) );
  XOR U17052 ( .A(b[49]), .B(a[40]), .Z(n16856) );
  NANDN U17053 ( .A(n37432), .B(n16856), .Z(n16534) );
  NAND U17054 ( .A(n16535), .B(n16534), .Z(n16889) );
  XOR U17055 ( .A(n16890), .B(n16889), .Z(n16892) );
  XOR U17056 ( .A(n16891), .B(n16892), .Z(n16962) );
  NANDN U17057 ( .A(n36742), .B(n16536), .Z(n16538) );
  XOR U17058 ( .A(b[43]), .B(a[46]), .Z(n16859) );
  NANDN U17059 ( .A(n36891), .B(n16859), .Z(n16537) );
  AND U17060 ( .A(n16538), .B(n16537), .Z(n16870) );
  NANDN U17061 ( .A(n36991), .B(n16539), .Z(n16541) );
  XOR U17062 ( .A(b[45]), .B(a[44]), .Z(n16862) );
  NANDN U17063 ( .A(n37083), .B(n16862), .Z(n16540) );
  AND U17064 ( .A(n16541), .B(n16540), .Z(n16869) );
  NANDN U17065 ( .A(n30482), .B(n16542), .Z(n16544) );
  XOR U17066 ( .A(a[78]), .B(b[11]), .Z(n16865) );
  NANDN U17067 ( .A(n30891), .B(n16865), .Z(n16543) );
  NAND U17068 ( .A(n16544), .B(n16543), .Z(n16868) );
  XOR U17069 ( .A(n16869), .B(n16868), .Z(n16871) );
  XNOR U17070 ( .A(n16870), .B(n16871), .Z(n16961) );
  XNOR U17071 ( .A(n16962), .B(n16961), .Z(n16963) );
  NANDN U17072 ( .A(n16546), .B(n16545), .Z(n16550) );
  OR U17073 ( .A(n16548), .B(n16547), .Z(n16549) );
  NAND U17074 ( .A(n16550), .B(n16549), .Z(n16964) );
  XNOR U17075 ( .A(n16963), .B(n16964), .Z(n17030) );
  XNOR U17076 ( .A(n17031), .B(n17030), .Z(n17033) );
  NANDN U17077 ( .A(n29499), .B(n16551), .Z(n16553) );
  XOR U17078 ( .A(a[82]), .B(b[7]), .Z(n16874) );
  NANDN U17079 ( .A(n29735), .B(n16874), .Z(n16552) );
  AND U17080 ( .A(n16553), .B(n16552), .Z(n16834) );
  NANDN U17081 ( .A(n37857), .B(n16554), .Z(n16556) );
  XOR U17082 ( .A(b[55]), .B(a[34]), .Z(n16877) );
  NANDN U17083 ( .A(n37911), .B(n16877), .Z(n16555) );
  AND U17084 ( .A(n16556), .B(n16555), .Z(n16833) );
  NANDN U17085 ( .A(n35611), .B(n16557), .Z(n16559) );
  XOR U17086 ( .A(b[35]), .B(a[54]), .Z(n16880) );
  NANDN U17087 ( .A(n35801), .B(n16880), .Z(n16558) );
  NAND U17088 ( .A(n16559), .B(n16558), .Z(n16832) );
  XOR U17089 ( .A(n16833), .B(n16832), .Z(n16835) );
  XOR U17090 ( .A(n16834), .B(n16835), .Z(n16902) );
  NANDN U17091 ( .A(n16561), .B(n16560), .Z(n16565) );
  OR U17092 ( .A(n16563), .B(n16562), .Z(n16564) );
  AND U17093 ( .A(n16565), .B(n16564), .Z(n16901) );
  XNOR U17094 ( .A(n16902), .B(n16901), .Z(n16903) );
  NANDN U17095 ( .A(n16567), .B(n16566), .Z(n16571) );
  OR U17096 ( .A(n16569), .B(n16568), .Z(n16570) );
  NAND U17097 ( .A(n16571), .B(n16570), .Z(n16904) );
  XNOR U17098 ( .A(n16903), .B(n16904), .Z(n17032) );
  XOR U17099 ( .A(n17033), .B(n17032), .Z(n17019) );
  NANDN U17100 ( .A(n16573), .B(n16572), .Z(n16577) );
  NANDN U17101 ( .A(n16575), .B(n16574), .Z(n16576) );
  AND U17102 ( .A(n16577), .B(n16576), .Z(n17039) );
  NANDN U17103 ( .A(n16579), .B(n16578), .Z(n16583) );
  NANDN U17104 ( .A(n16581), .B(n16580), .Z(n16582) );
  AND U17105 ( .A(n16583), .B(n16582), .Z(n17037) );
  NANDN U17106 ( .A(n33875), .B(n16584), .Z(n16586) );
  XOR U17107 ( .A(b[25]), .B(a[64]), .Z(n16808) );
  NANDN U17108 ( .A(n33994), .B(n16808), .Z(n16585) );
  AND U17109 ( .A(n16586), .B(n16585), .Z(n16984) );
  NANDN U17110 ( .A(n32013), .B(n16587), .Z(n16589) );
  XOR U17111 ( .A(b[17]), .B(a[72]), .Z(n16811) );
  NANDN U17112 ( .A(n32292), .B(n16811), .Z(n16588) );
  AND U17113 ( .A(n16589), .B(n16588), .Z(n16983) );
  NANDN U17114 ( .A(n31536), .B(n16590), .Z(n16592) );
  XOR U17115 ( .A(b[15]), .B(a[74]), .Z(n16814) );
  NANDN U17116 ( .A(n31925), .B(n16814), .Z(n16591) );
  NAND U17117 ( .A(n16592), .B(n16591), .Z(n16982) );
  XOR U17118 ( .A(n16983), .B(n16982), .Z(n16985) );
  XOR U17119 ( .A(n16984), .B(n16985), .Z(n16956) );
  NANDN U17120 ( .A(n37526), .B(n16593), .Z(n16595) );
  XOR U17121 ( .A(b[51]), .B(a[38]), .Z(n16817) );
  NANDN U17122 ( .A(n37605), .B(n16817), .Z(n16594) );
  AND U17123 ( .A(n16595), .B(n16594), .Z(n17008) );
  NANDN U17124 ( .A(n37705), .B(n16596), .Z(n16598) );
  XOR U17125 ( .A(b[53]), .B(a[36]), .Z(n16820) );
  NANDN U17126 ( .A(n37778), .B(n16820), .Z(n16597) );
  AND U17127 ( .A(n16598), .B(n16597), .Z(n17007) );
  NANDN U17128 ( .A(n36210), .B(n16599), .Z(n16601) );
  XOR U17129 ( .A(b[39]), .B(a[50]), .Z(n16823) );
  NANDN U17130 ( .A(n36347), .B(n16823), .Z(n16600) );
  NAND U17131 ( .A(n16601), .B(n16600), .Z(n17006) );
  XOR U17132 ( .A(n17007), .B(n17006), .Z(n17009) );
  XNOR U17133 ( .A(n17008), .B(n17009), .Z(n16955) );
  XNOR U17134 ( .A(n16956), .B(n16955), .Z(n16958) );
  NANDN U17135 ( .A(n16603), .B(n16602), .Z(n16607) );
  OR U17136 ( .A(n16605), .B(n16604), .Z(n16606) );
  AND U17137 ( .A(n16607), .B(n16606), .Z(n16957) );
  XOR U17138 ( .A(n16958), .B(n16957), .Z(n16799) );
  NANDN U17139 ( .A(n16609), .B(n16608), .Z(n16613) );
  OR U17140 ( .A(n16611), .B(n16610), .Z(n16612) );
  AND U17141 ( .A(n16613), .B(n16612), .Z(n16797) );
  NANDN U17142 ( .A(n16615), .B(n16614), .Z(n16619) );
  NANDN U17143 ( .A(n16617), .B(n16616), .Z(n16618) );
  NAND U17144 ( .A(n16619), .B(n16618), .Z(n16796) );
  XNOR U17145 ( .A(n16797), .B(n16796), .Z(n16798) );
  XNOR U17146 ( .A(n16799), .B(n16798), .Z(n17036) );
  XNOR U17147 ( .A(n17037), .B(n17036), .Z(n17038) );
  XNOR U17148 ( .A(n17039), .B(n17038), .Z(n17018) );
  XNOR U17149 ( .A(n17019), .B(n17018), .Z(n17020) );
  NANDN U17150 ( .A(n16621), .B(n16620), .Z(n16625) );
  NAND U17151 ( .A(n16623), .B(n16622), .Z(n16624) );
  NAND U17152 ( .A(n16625), .B(n16624), .Z(n17021) );
  XNOR U17153 ( .A(n17020), .B(n17021), .Z(n17042) );
  NANDN U17154 ( .A(n16627), .B(n16626), .Z(n16631) );
  NANDN U17155 ( .A(n16629), .B(n16628), .Z(n16630) );
  AND U17156 ( .A(n16631), .B(n16630), .Z(n17026) );
  NANDN U17157 ( .A(n16633), .B(n16632), .Z(n16637) );
  NANDN U17158 ( .A(n16635), .B(n16634), .Z(n16636) );
  AND U17159 ( .A(n16637), .B(n16636), .Z(n17025) );
  NANDN U17160 ( .A(n16639), .B(n16638), .Z(n16643) );
  NAND U17161 ( .A(n16641), .B(n16640), .Z(n16642) );
  AND U17162 ( .A(n16643), .B(n16642), .Z(n17024) );
  XOR U17163 ( .A(n17025), .B(n17024), .Z(n17027) );
  XOR U17164 ( .A(n17026), .B(n17027), .Z(n16793) );
  NANDN U17165 ( .A(n16645), .B(n16644), .Z(n16649) );
  NANDN U17166 ( .A(n16647), .B(n16646), .Z(n16648) );
  AND U17167 ( .A(n16649), .B(n16648), .Z(n16790) );
  NANDN U17168 ( .A(n16651), .B(n16650), .Z(n16655) );
  NANDN U17169 ( .A(n16653), .B(n16652), .Z(n16654) );
  AND U17170 ( .A(n16655), .B(n16654), .Z(n17014) );
  NANDN U17171 ( .A(n32996), .B(n16656), .Z(n16658) );
  XOR U17172 ( .A(b[21]), .B(a[68]), .Z(n16967) );
  NANDN U17173 ( .A(n33271), .B(n16967), .Z(n16657) );
  AND U17174 ( .A(n16658), .B(n16657), .Z(n16933) );
  NANDN U17175 ( .A(n33866), .B(n16659), .Z(n16661) );
  XOR U17176 ( .A(b[23]), .B(a[66]), .Z(n16970) );
  NANDN U17177 ( .A(n33644), .B(n16970), .Z(n16660) );
  AND U17178 ( .A(n16661), .B(n16660), .Z(n16932) );
  NANDN U17179 ( .A(n32483), .B(n16662), .Z(n16664) );
  XOR U17180 ( .A(b[19]), .B(a[70]), .Z(n16973) );
  NANDN U17181 ( .A(n32823), .B(n16973), .Z(n16663) );
  NAND U17182 ( .A(n16664), .B(n16663), .Z(n16931) );
  XOR U17183 ( .A(n16932), .B(n16931), .Z(n16934) );
  XOR U17184 ( .A(n16933), .B(n16934), .Z(n16845) );
  NANDN U17185 ( .A(n34909), .B(n16665), .Z(n16667) );
  XOR U17186 ( .A(b[31]), .B(a[58]), .Z(n16976) );
  NANDN U17187 ( .A(n35145), .B(n16976), .Z(n16666) );
  AND U17188 ( .A(n16667), .B(n16666), .Z(n16885) );
  NANDN U17189 ( .A(n38247), .B(n16668), .Z(n16670) );
  XOR U17190 ( .A(b[61]), .B(a[28]), .Z(n16979) );
  NANDN U17191 ( .A(n38248), .B(n16979), .Z(n16669) );
  AND U17192 ( .A(n16670), .B(n16669), .Z(n16884) );
  AND U17193 ( .A(b[63]), .B(a[24]), .Z(n16883) );
  XOR U17194 ( .A(n16884), .B(n16883), .Z(n16886) );
  XNOR U17195 ( .A(n16885), .B(n16886), .Z(n16844) );
  XNOR U17196 ( .A(n16845), .B(n16844), .Z(n16846) );
  NANDN U17197 ( .A(n16672), .B(n16671), .Z(n16676) );
  OR U17198 ( .A(n16674), .B(n16673), .Z(n16675) );
  NAND U17199 ( .A(n16676), .B(n16675), .Z(n16847) );
  XNOR U17200 ( .A(n16846), .B(n16847), .Z(n17012) );
  NANDN U17201 ( .A(n34223), .B(n16677), .Z(n16679) );
  XOR U17202 ( .A(b[27]), .B(a[62]), .Z(n16988) );
  NANDN U17203 ( .A(n34458), .B(n16988), .Z(n16678) );
  AND U17204 ( .A(n16679), .B(n16678), .Z(n16828) );
  NANDN U17205 ( .A(n34634), .B(n16680), .Z(n16682) );
  XOR U17206 ( .A(b[29]), .B(a[60]), .Z(n16991) );
  NANDN U17207 ( .A(n34722), .B(n16991), .Z(n16681) );
  AND U17208 ( .A(n16682), .B(n16681), .Z(n16827) );
  NANDN U17209 ( .A(n31055), .B(n16683), .Z(n16685) );
  XOR U17210 ( .A(b[13]), .B(a[76]), .Z(n16994) );
  NANDN U17211 ( .A(n31293), .B(n16994), .Z(n16684) );
  NAND U17212 ( .A(n16685), .B(n16684), .Z(n16826) );
  XOR U17213 ( .A(n16827), .B(n16826), .Z(n16829) );
  XOR U17214 ( .A(n16828), .B(n16829), .Z(n16908) );
  NANDN U17215 ( .A(n28889), .B(n16686), .Z(n16688) );
  XOR U17216 ( .A(a[84]), .B(b[5]), .Z(n16997) );
  NANDN U17217 ( .A(n29138), .B(n16997), .Z(n16687) );
  AND U17218 ( .A(n16688), .B(n16687), .Z(n16927) );
  NANDN U17219 ( .A(n209), .B(n16689), .Z(n16691) );
  XOR U17220 ( .A(a[86]), .B(b[3]), .Z(n17000) );
  NANDN U17221 ( .A(n28941), .B(n17000), .Z(n16690) );
  AND U17222 ( .A(n16691), .B(n16690), .Z(n16926) );
  NANDN U17223 ( .A(n35936), .B(n16692), .Z(n16694) );
  XOR U17224 ( .A(b[37]), .B(a[52]), .Z(n17003) );
  NANDN U17225 ( .A(n36047), .B(n17003), .Z(n16693) );
  NAND U17226 ( .A(n16694), .B(n16693), .Z(n16925) );
  XOR U17227 ( .A(n16926), .B(n16925), .Z(n16928) );
  XNOR U17228 ( .A(n16927), .B(n16928), .Z(n16907) );
  XNOR U17229 ( .A(n16908), .B(n16907), .Z(n16909) );
  NANDN U17230 ( .A(n16696), .B(n16695), .Z(n16700) );
  OR U17231 ( .A(n16698), .B(n16697), .Z(n16699) );
  NAND U17232 ( .A(n16700), .B(n16699), .Z(n16910) );
  XOR U17233 ( .A(n16909), .B(n16910), .Z(n17013) );
  XOR U17234 ( .A(n17012), .B(n17013), .Z(n17015) );
  XOR U17235 ( .A(n17014), .B(n17015), .Z(n16898) );
  NANDN U17236 ( .A(n16702), .B(n16701), .Z(n16706) );
  NAND U17237 ( .A(n16704), .B(n16703), .Z(n16705) );
  AND U17238 ( .A(n16706), .B(n16705), .Z(n16895) );
  NANDN U17239 ( .A(n16708), .B(n16707), .Z(n16712) );
  NANDN U17240 ( .A(n16710), .B(n16709), .Z(n16711) );
  AND U17241 ( .A(n16712), .B(n16711), .Z(n16914) );
  NANDN U17242 ( .A(n16714), .B(n16713), .Z(n16718) );
  OR U17243 ( .A(n16716), .B(n16715), .Z(n16717) );
  NAND U17244 ( .A(n16718), .B(n16717), .Z(n16913) );
  XNOR U17245 ( .A(n16914), .B(n16913), .Z(n16915) );
  NANDN U17246 ( .A(n16720), .B(n16719), .Z(n16724) );
  OR U17247 ( .A(n16722), .B(n16721), .Z(n16723) );
  AND U17248 ( .A(n16724), .B(n16723), .Z(n16805) );
  NANDN U17249 ( .A(n38278), .B(n16725), .Z(n16727) );
  XOR U17250 ( .A(b[63]), .B(a[26]), .Z(n16940) );
  NANDN U17251 ( .A(n38279), .B(n16940), .Z(n16726) );
  AND U17252 ( .A(n16727), .B(n16726), .Z(n16839) );
  NANDN U17253 ( .A(n35260), .B(n16728), .Z(n16730) );
  XOR U17254 ( .A(b[33]), .B(a[56]), .Z(n16943) );
  NANDN U17255 ( .A(n35456), .B(n16943), .Z(n16729) );
  NAND U17256 ( .A(n16730), .B(n16729), .Z(n16838) );
  XNOR U17257 ( .A(n16839), .B(n16838), .Z(n16840) );
  NAND U17258 ( .A(b[0]), .B(a[88]), .Z(n16731) );
  XNOR U17259 ( .A(b[1]), .B(n16731), .Z(n16733) );
  NANDN U17260 ( .A(b[0]), .B(a[87]), .Z(n16732) );
  NAND U17261 ( .A(n16733), .B(n16732), .Z(n16841) );
  XNOR U17262 ( .A(n16840), .B(n16841), .Z(n16802) );
  NANDN U17263 ( .A(n37974), .B(n16734), .Z(n16736) );
  XOR U17264 ( .A(b[57]), .B(a[32]), .Z(n16946) );
  NANDN U17265 ( .A(n38031), .B(n16946), .Z(n16735) );
  AND U17266 ( .A(n16736), .B(n16735), .Z(n16922) );
  NANDN U17267 ( .A(n38090), .B(n16737), .Z(n16739) );
  XOR U17268 ( .A(b[59]), .B(a[30]), .Z(n16949) );
  NANDN U17269 ( .A(n38130), .B(n16949), .Z(n16738) );
  AND U17270 ( .A(n16739), .B(n16738), .Z(n16920) );
  NANDN U17271 ( .A(n36480), .B(n16740), .Z(n16742) );
  XOR U17272 ( .A(b[41]), .B(a[48]), .Z(n16952) );
  NANDN U17273 ( .A(n36594), .B(n16952), .Z(n16741) );
  NAND U17274 ( .A(n16742), .B(n16741), .Z(n16919) );
  XNOR U17275 ( .A(n16920), .B(n16919), .Z(n16921) );
  XOR U17276 ( .A(n16922), .B(n16921), .Z(n16803) );
  XNOR U17277 ( .A(n16802), .B(n16803), .Z(n16804) );
  XOR U17278 ( .A(n16805), .B(n16804), .Z(n16916) );
  XOR U17279 ( .A(n16915), .B(n16916), .Z(n16896) );
  XNOR U17280 ( .A(n16895), .B(n16896), .Z(n16897) );
  XOR U17281 ( .A(n16898), .B(n16897), .Z(n16791) );
  XNOR U17282 ( .A(n16790), .B(n16791), .Z(n16792) );
  XOR U17283 ( .A(n16793), .B(n16792), .Z(n17043) );
  XNOR U17284 ( .A(n17042), .B(n17043), .Z(n17044) );
  XOR U17285 ( .A(n17045), .B(n17044), .Z(n17057) );
  XNOR U17286 ( .A(n17056), .B(n17057), .Z(n17063) );
  NANDN U17287 ( .A(n16744), .B(n16743), .Z(n16748) );
  NANDN U17288 ( .A(n16746), .B(n16745), .Z(n16747) );
  AND U17289 ( .A(n16748), .B(n16747), .Z(n17061) );
  NANDN U17290 ( .A(n16750), .B(n16749), .Z(n16754) );
  NANDN U17291 ( .A(n16752), .B(n16751), .Z(n16753) );
  NAND U17292 ( .A(n16754), .B(n16753), .Z(n17060) );
  XNOR U17293 ( .A(n17061), .B(n17060), .Z(n17062) );
  XOR U17294 ( .A(n17063), .B(n17062), .Z(n16785) );
  NANDN U17295 ( .A(n16756), .B(n16755), .Z(n16760) );
  NANDN U17296 ( .A(n16758), .B(n16757), .Z(n16759) );
  AND U17297 ( .A(n16760), .B(n16759), .Z(n16784) );
  XNOR U17298 ( .A(n16785), .B(n16784), .Z(n16786) );
  NANDN U17299 ( .A(n16762), .B(n16761), .Z(n16766) );
  NANDN U17300 ( .A(n16764), .B(n16763), .Z(n16765) );
  NAND U17301 ( .A(n16766), .B(n16765), .Z(n16787) );
  XNOR U17302 ( .A(n16786), .B(n16787), .Z(n16778) );
  NANDN U17303 ( .A(n16768), .B(n16767), .Z(n16772) );
  OR U17304 ( .A(n16770), .B(n16769), .Z(n16771) );
  NAND U17305 ( .A(n16772), .B(n16771), .Z(n16779) );
  XNOR U17306 ( .A(n16778), .B(n16779), .Z(n16780) );
  XNOR U17307 ( .A(n16781), .B(n16780), .Z(n17066) );
  XNOR U17308 ( .A(sreg[152]), .B(n17066), .Z(n17068) );
  NANDN U17309 ( .A(sreg[151]), .B(n16773), .Z(n16777) );
  NAND U17310 ( .A(n16775), .B(n16774), .Z(n16776) );
  NAND U17311 ( .A(n16777), .B(n16776), .Z(n17067) );
  XNOR U17312 ( .A(n17068), .B(n17067), .Z(c[152]) );
  NANDN U17313 ( .A(n16779), .B(n16778), .Z(n16783) );
  NANDN U17314 ( .A(n16781), .B(n16780), .Z(n16782) );
  AND U17315 ( .A(n16783), .B(n16782), .Z(n17074) );
  NANDN U17316 ( .A(n16785), .B(n16784), .Z(n16789) );
  NANDN U17317 ( .A(n16787), .B(n16786), .Z(n16788) );
  AND U17318 ( .A(n16789), .B(n16788), .Z(n17072) );
  NANDN U17319 ( .A(n16791), .B(n16790), .Z(n16795) );
  NANDN U17320 ( .A(n16793), .B(n16792), .Z(n16794) );
  AND U17321 ( .A(n16795), .B(n16794), .Z(n17337) );
  NANDN U17322 ( .A(n16797), .B(n16796), .Z(n16801) );
  NANDN U17323 ( .A(n16799), .B(n16798), .Z(n16800) );
  AND U17324 ( .A(n16801), .B(n16800), .Z(n17097) );
  NANDN U17325 ( .A(n16803), .B(n16802), .Z(n16807) );
  NANDN U17326 ( .A(n16805), .B(n16804), .Z(n16806) );
  AND U17327 ( .A(n16807), .B(n16806), .Z(n17096) );
  NANDN U17328 ( .A(n33875), .B(n16808), .Z(n16810) );
  XOR U17329 ( .A(b[25]), .B(a[65]), .Z(n17182) );
  NANDN U17330 ( .A(n33994), .B(n17182), .Z(n16809) );
  AND U17331 ( .A(n16810), .B(n16809), .Z(n17259) );
  NANDN U17332 ( .A(n32013), .B(n16811), .Z(n16813) );
  XOR U17333 ( .A(b[17]), .B(a[73]), .Z(n17185) );
  NANDN U17334 ( .A(n32292), .B(n17185), .Z(n16812) );
  AND U17335 ( .A(n16813), .B(n16812), .Z(n17258) );
  NANDN U17336 ( .A(n31536), .B(n16814), .Z(n16816) );
  XOR U17337 ( .A(b[15]), .B(a[75]), .Z(n17188) );
  NANDN U17338 ( .A(n31925), .B(n17188), .Z(n16815) );
  NAND U17339 ( .A(n16816), .B(n16815), .Z(n17257) );
  XOR U17340 ( .A(n17258), .B(n17257), .Z(n17260) );
  XOR U17341 ( .A(n17259), .B(n17260), .Z(n17324) );
  NANDN U17342 ( .A(n37526), .B(n16817), .Z(n16819) );
  XOR U17343 ( .A(b[51]), .B(a[39]), .Z(n17191) );
  NANDN U17344 ( .A(n37605), .B(n17191), .Z(n16818) );
  AND U17345 ( .A(n16819), .B(n16818), .Z(n17283) );
  NANDN U17346 ( .A(n37705), .B(n16820), .Z(n16822) );
  XOR U17347 ( .A(b[53]), .B(a[37]), .Z(n17194) );
  NANDN U17348 ( .A(n37778), .B(n17194), .Z(n16821) );
  AND U17349 ( .A(n16822), .B(n16821), .Z(n17282) );
  NANDN U17350 ( .A(n36210), .B(n16823), .Z(n16825) );
  XOR U17351 ( .A(b[39]), .B(a[51]), .Z(n17197) );
  NANDN U17352 ( .A(n36347), .B(n17197), .Z(n16824) );
  NAND U17353 ( .A(n16825), .B(n16824), .Z(n17281) );
  XOR U17354 ( .A(n17282), .B(n17281), .Z(n17284) );
  XNOR U17355 ( .A(n17283), .B(n17284), .Z(n17323) );
  XNOR U17356 ( .A(n17324), .B(n17323), .Z(n17326) );
  NANDN U17357 ( .A(n16827), .B(n16826), .Z(n16831) );
  OR U17358 ( .A(n16829), .B(n16828), .Z(n16830) );
  AND U17359 ( .A(n16831), .B(n16830), .Z(n17325) );
  XOR U17360 ( .A(n17326), .B(n17325), .Z(n17173) );
  NANDN U17361 ( .A(n16833), .B(n16832), .Z(n16837) );
  OR U17362 ( .A(n16835), .B(n16834), .Z(n16836) );
  AND U17363 ( .A(n16837), .B(n16836), .Z(n17171) );
  NANDN U17364 ( .A(n16839), .B(n16838), .Z(n16843) );
  NANDN U17365 ( .A(n16841), .B(n16840), .Z(n16842) );
  NAND U17366 ( .A(n16843), .B(n16842), .Z(n17170) );
  XNOR U17367 ( .A(n17171), .B(n17170), .Z(n17172) );
  XNOR U17368 ( .A(n17173), .B(n17172), .Z(n17095) );
  XOR U17369 ( .A(n17096), .B(n17095), .Z(n17098) );
  XOR U17370 ( .A(n17097), .B(n17098), .Z(n17102) );
  NANDN U17371 ( .A(n16845), .B(n16844), .Z(n16849) );
  NANDN U17372 ( .A(n16847), .B(n16846), .Z(n16848) );
  AND U17373 ( .A(n16849), .B(n16848), .Z(n17090) );
  NANDN U17374 ( .A(n211), .B(n16850), .Z(n16852) );
  XOR U17375 ( .A(b[47]), .B(a[43]), .Z(n17125) );
  NANDN U17376 ( .A(n37172), .B(n17125), .Z(n16851) );
  AND U17377 ( .A(n16852), .B(n16851), .Z(n17166) );
  NANDN U17378 ( .A(n210), .B(n16853), .Z(n16855) );
  XOR U17379 ( .A(a[81]), .B(b[9]), .Z(n17128) );
  NANDN U17380 ( .A(n30267), .B(n17128), .Z(n16854) );
  AND U17381 ( .A(n16855), .B(n16854), .Z(n17165) );
  NANDN U17382 ( .A(n212), .B(n16856), .Z(n16858) );
  XOR U17383 ( .A(b[49]), .B(a[41]), .Z(n17131) );
  NANDN U17384 ( .A(n37432), .B(n17131), .Z(n16857) );
  NAND U17385 ( .A(n16858), .B(n16857), .Z(n17164) );
  XOR U17386 ( .A(n17165), .B(n17164), .Z(n17167) );
  XOR U17387 ( .A(n17166), .B(n17167), .Z(n17237) );
  NANDN U17388 ( .A(n36742), .B(n16859), .Z(n16861) );
  XOR U17389 ( .A(b[43]), .B(a[47]), .Z(n17134) );
  NANDN U17390 ( .A(n36891), .B(n17134), .Z(n16860) );
  AND U17391 ( .A(n16861), .B(n16860), .Z(n17145) );
  NANDN U17392 ( .A(n36991), .B(n16862), .Z(n16864) );
  XOR U17393 ( .A(b[45]), .B(a[45]), .Z(n17137) );
  NANDN U17394 ( .A(n37083), .B(n17137), .Z(n16863) );
  AND U17395 ( .A(n16864), .B(n16863), .Z(n17144) );
  NANDN U17396 ( .A(n30482), .B(n16865), .Z(n16867) );
  XOR U17397 ( .A(a[79]), .B(b[11]), .Z(n17140) );
  NANDN U17398 ( .A(n30891), .B(n17140), .Z(n16866) );
  NAND U17399 ( .A(n16867), .B(n16866), .Z(n17143) );
  XOR U17400 ( .A(n17144), .B(n17143), .Z(n17146) );
  XNOR U17401 ( .A(n17145), .B(n17146), .Z(n17236) );
  XNOR U17402 ( .A(n17237), .B(n17236), .Z(n17238) );
  NANDN U17403 ( .A(n16869), .B(n16868), .Z(n16873) );
  OR U17404 ( .A(n16871), .B(n16870), .Z(n16872) );
  NAND U17405 ( .A(n16873), .B(n16872), .Z(n17239) );
  XNOR U17406 ( .A(n17238), .B(n17239), .Z(n17089) );
  XNOR U17407 ( .A(n17090), .B(n17089), .Z(n17091) );
  NANDN U17408 ( .A(n29499), .B(n16874), .Z(n16876) );
  XOR U17409 ( .A(a[83]), .B(b[7]), .Z(n17149) );
  NANDN U17410 ( .A(n29735), .B(n17149), .Z(n16875) );
  AND U17411 ( .A(n16876), .B(n16875), .Z(n17208) );
  NANDN U17412 ( .A(n37857), .B(n16877), .Z(n16879) );
  XOR U17413 ( .A(b[55]), .B(a[35]), .Z(n17152) );
  NANDN U17414 ( .A(n37911), .B(n17152), .Z(n16878) );
  AND U17415 ( .A(n16879), .B(n16878), .Z(n17207) );
  NANDN U17416 ( .A(n35611), .B(n16880), .Z(n16882) );
  XOR U17417 ( .A(b[35]), .B(a[55]), .Z(n17155) );
  NANDN U17418 ( .A(n35801), .B(n17155), .Z(n16881) );
  NAND U17419 ( .A(n16882), .B(n16881), .Z(n17206) );
  XOR U17420 ( .A(n17207), .B(n17206), .Z(n17209) );
  XOR U17421 ( .A(n17208), .B(n17209), .Z(n17219) );
  NANDN U17422 ( .A(n16884), .B(n16883), .Z(n16888) );
  OR U17423 ( .A(n16886), .B(n16885), .Z(n16887) );
  AND U17424 ( .A(n16888), .B(n16887), .Z(n17218) );
  XNOR U17425 ( .A(n17219), .B(n17218), .Z(n17220) );
  NANDN U17426 ( .A(n16890), .B(n16889), .Z(n16894) );
  OR U17427 ( .A(n16892), .B(n16891), .Z(n16893) );
  NAND U17428 ( .A(n16894), .B(n16893), .Z(n17221) );
  XOR U17429 ( .A(n17220), .B(n17221), .Z(n17092) );
  XNOR U17430 ( .A(n17091), .B(n17092), .Z(n17101) );
  XNOR U17431 ( .A(n17102), .B(n17101), .Z(n17104) );
  NANDN U17432 ( .A(n16896), .B(n16895), .Z(n16900) );
  NANDN U17433 ( .A(n16898), .B(n16897), .Z(n16899) );
  AND U17434 ( .A(n16900), .B(n16899), .Z(n17103) );
  XOR U17435 ( .A(n17104), .B(n17103), .Z(n17336) );
  NANDN U17436 ( .A(n16902), .B(n16901), .Z(n16906) );
  NANDN U17437 ( .A(n16904), .B(n16903), .Z(n16905) );
  AND U17438 ( .A(n16906), .B(n16905), .Z(n17085) );
  NANDN U17439 ( .A(n16908), .B(n16907), .Z(n16912) );
  NANDN U17440 ( .A(n16910), .B(n16909), .Z(n16911) );
  AND U17441 ( .A(n16912), .B(n16911), .Z(n17084) );
  NANDN U17442 ( .A(n16914), .B(n16913), .Z(n16918) );
  NANDN U17443 ( .A(n16916), .B(n16915), .Z(n16917) );
  AND U17444 ( .A(n16918), .B(n16917), .Z(n17083) );
  XOR U17445 ( .A(n17084), .B(n17083), .Z(n17086) );
  XOR U17446 ( .A(n17085), .B(n17086), .Z(n17110) );
  NANDN U17447 ( .A(n16920), .B(n16919), .Z(n16924) );
  NANDN U17448 ( .A(n16922), .B(n16921), .Z(n16923) );
  AND U17449 ( .A(n16924), .B(n16923), .Z(n17231) );
  NANDN U17450 ( .A(n16926), .B(n16925), .Z(n16930) );
  OR U17451 ( .A(n16928), .B(n16927), .Z(n16929) );
  NAND U17452 ( .A(n16930), .B(n16929), .Z(n17230) );
  XNOR U17453 ( .A(n17231), .B(n17230), .Z(n17233) );
  NANDN U17454 ( .A(n16932), .B(n16931), .Z(n16936) );
  OR U17455 ( .A(n16934), .B(n16933), .Z(n16935) );
  AND U17456 ( .A(n16936), .B(n16935), .Z(n17179) );
  NAND U17457 ( .A(b[0]), .B(a[89]), .Z(n16937) );
  XNOR U17458 ( .A(b[1]), .B(n16937), .Z(n16939) );
  NANDN U17459 ( .A(b[0]), .B(a[88]), .Z(n16938) );
  NAND U17460 ( .A(n16939), .B(n16938), .Z(n17215) );
  NANDN U17461 ( .A(n38278), .B(n16940), .Z(n16942) );
  XOR U17462 ( .A(b[63]), .B(a[27]), .Z(n17305) );
  NANDN U17463 ( .A(n38279), .B(n17305), .Z(n16941) );
  AND U17464 ( .A(n16942), .B(n16941), .Z(n17213) );
  NANDN U17465 ( .A(n35260), .B(n16943), .Z(n16945) );
  XOR U17466 ( .A(b[33]), .B(a[57]), .Z(n17308) );
  NANDN U17467 ( .A(n35456), .B(n17308), .Z(n16944) );
  NAND U17468 ( .A(n16945), .B(n16944), .Z(n17212) );
  XNOR U17469 ( .A(n17213), .B(n17212), .Z(n17214) );
  XNOR U17470 ( .A(n17215), .B(n17214), .Z(n17176) );
  NANDN U17471 ( .A(n37974), .B(n16946), .Z(n16948) );
  XOR U17472 ( .A(b[57]), .B(a[33]), .Z(n17314) );
  NANDN U17473 ( .A(n38031), .B(n17314), .Z(n16947) );
  AND U17474 ( .A(n16948), .B(n16947), .Z(n17290) );
  NANDN U17475 ( .A(n38090), .B(n16949), .Z(n16951) );
  XOR U17476 ( .A(b[59]), .B(a[31]), .Z(n17317) );
  NANDN U17477 ( .A(n38130), .B(n17317), .Z(n16950) );
  AND U17478 ( .A(n16951), .B(n16950), .Z(n17288) );
  NANDN U17479 ( .A(n36480), .B(n16952), .Z(n16954) );
  XOR U17480 ( .A(b[41]), .B(a[49]), .Z(n17320) );
  NANDN U17481 ( .A(n36594), .B(n17320), .Z(n16953) );
  NAND U17482 ( .A(n16954), .B(n16953), .Z(n17287) );
  XNOR U17483 ( .A(n17288), .B(n17287), .Z(n17289) );
  XOR U17484 ( .A(n17290), .B(n17289), .Z(n17177) );
  XNOR U17485 ( .A(n17176), .B(n17177), .Z(n17178) );
  XNOR U17486 ( .A(n17179), .B(n17178), .Z(n17232) );
  XOR U17487 ( .A(n17233), .B(n17232), .Z(n17114) );
  NANDN U17488 ( .A(n16956), .B(n16955), .Z(n16960) );
  NAND U17489 ( .A(n16958), .B(n16957), .Z(n16959) );
  NAND U17490 ( .A(n16960), .B(n16959), .Z(n17113) );
  XNOR U17491 ( .A(n17114), .B(n17113), .Z(n17116) );
  NANDN U17492 ( .A(n16962), .B(n16961), .Z(n16966) );
  NANDN U17493 ( .A(n16964), .B(n16963), .Z(n16965) );
  AND U17494 ( .A(n16966), .B(n16965), .Z(n17332) );
  NANDN U17495 ( .A(n32996), .B(n16967), .Z(n16969) );
  XOR U17496 ( .A(b[21]), .B(a[69]), .Z(n17242) );
  NANDN U17497 ( .A(n33271), .B(n17242), .Z(n16968) );
  AND U17498 ( .A(n16969), .B(n16968), .Z(n17301) );
  NANDN U17499 ( .A(n33866), .B(n16970), .Z(n16972) );
  XOR U17500 ( .A(b[23]), .B(a[67]), .Z(n17245) );
  NANDN U17501 ( .A(n33644), .B(n17245), .Z(n16971) );
  AND U17502 ( .A(n16972), .B(n16971), .Z(n17300) );
  NANDN U17503 ( .A(n32483), .B(n16973), .Z(n16975) );
  XOR U17504 ( .A(b[19]), .B(a[71]), .Z(n17248) );
  NANDN U17505 ( .A(n32823), .B(n17248), .Z(n16974) );
  NAND U17506 ( .A(n16975), .B(n16974), .Z(n17299) );
  XOR U17507 ( .A(n17300), .B(n17299), .Z(n17302) );
  XOR U17508 ( .A(n17301), .B(n17302), .Z(n17120) );
  NANDN U17509 ( .A(n34909), .B(n16976), .Z(n16978) );
  XOR U17510 ( .A(b[31]), .B(a[59]), .Z(n17251) );
  NANDN U17511 ( .A(n35145), .B(n17251), .Z(n16977) );
  AND U17512 ( .A(n16978), .B(n16977), .Z(n17160) );
  NANDN U17513 ( .A(n38247), .B(n16979), .Z(n16981) );
  XOR U17514 ( .A(b[61]), .B(a[29]), .Z(n17254) );
  NANDN U17515 ( .A(n38248), .B(n17254), .Z(n16980) );
  AND U17516 ( .A(n16981), .B(n16980), .Z(n17159) );
  AND U17517 ( .A(b[63]), .B(a[25]), .Z(n17158) );
  XOR U17518 ( .A(n17159), .B(n17158), .Z(n17161) );
  XNOR U17519 ( .A(n17160), .B(n17161), .Z(n17119) );
  XNOR U17520 ( .A(n17120), .B(n17119), .Z(n17121) );
  NANDN U17521 ( .A(n16983), .B(n16982), .Z(n16987) );
  OR U17522 ( .A(n16985), .B(n16984), .Z(n16986) );
  NAND U17523 ( .A(n16987), .B(n16986), .Z(n17122) );
  XNOR U17524 ( .A(n17121), .B(n17122), .Z(n17329) );
  NANDN U17525 ( .A(n34223), .B(n16988), .Z(n16990) );
  XOR U17526 ( .A(b[27]), .B(a[63]), .Z(n17263) );
  NANDN U17527 ( .A(n34458), .B(n17263), .Z(n16989) );
  AND U17528 ( .A(n16990), .B(n16989), .Z(n17202) );
  NANDN U17529 ( .A(n34634), .B(n16991), .Z(n16993) );
  XOR U17530 ( .A(b[29]), .B(a[61]), .Z(n17266) );
  NANDN U17531 ( .A(n34722), .B(n17266), .Z(n16992) );
  AND U17532 ( .A(n16993), .B(n16992), .Z(n17201) );
  NANDN U17533 ( .A(n31055), .B(n16994), .Z(n16996) );
  XOR U17534 ( .A(b[13]), .B(a[77]), .Z(n17269) );
  NANDN U17535 ( .A(n31293), .B(n17269), .Z(n16995) );
  NAND U17536 ( .A(n16996), .B(n16995), .Z(n17200) );
  XOR U17537 ( .A(n17201), .B(n17200), .Z(n17203) );
  XOR U17538 ( .A(n17202), .B(n17203), .Z(n17225) );
  NANDN U17539 ( .A(n28889), .B(n16997), .Z(n16999) );
  XOR U17540 ( .A(a[85]), .B(b[5]), .Z(n17272) );
  NANDN U17541 ( .A(n29138), .B(n17272), .Z(n16998) );
  AND U17542 ( .A(n16999), .B(n16998), .Z(n17295) );
  NANDN U17543 ( .A(n209), .B(n17000), .Z(n17002) );
  XOR U17544 ( .A(a[87]), .B(b[3]), .Z(n17275) );
  NANDN U17545 ( .A(n28941), .B(n17275), .Z(n17001) );
  AND U17546 ( .A(n17002), .B(n17001), .Z(n17294) );
  NANDN U17547 ( .A(n35936), .B(n17003), .Z(n17005) );
  XOR U17548 ( .A(b[37]), .B(a[53]), .Z(n17278) );
  NANDN U17549 ( .A(n36047), .B(n17278), .Z(n17004) );
  NAND U17550 ( .A(n17005), .B(n17004), .Z(n17293) );
  XOR U17551 ( .A(n17294), .B(n17293), .Z(n17296) );
  XNOR U17552 ( .A(n17295), .B(n17296), .Z(n17224) );
  XNOR U17553 ( .A(n17225), .B(n17224), .Z(n17226) );
  NANDN U17554 ( .A(n17007), .B(n17006), .Z(n17011) );
  OR U17555 ( .A(n17009), .B(n17008), .Z(n17010) );
  NAND U17556 ( .A(n17011), .B(n17010), .Z(n17227) );
  XOR U17557 ( .A(n17226), .B(n17227), .Z(n17330) );
  XNOR U17558 ( .A(n17329), .B(n17330), .Z(n17331) );
  XNOR U17559 ( .A(n17332), .B(n17331), .Z(n17115) );
  XOR U17560 ( .A(n17116), .B(n17115), .Z(n17108) );
  NANDN U17561 ( .A(n17013), .B(n17012), .Z(n17017) );
  OR U17562 ( .A(n17015), .B(n17014), .Z(n17016) );
  AND U17563 ( .A(n17017), .B(n17016), .Z(n17107) );
  XNOR U17564 ( .A(n17108), .B(n17107), .Z(n17109) );
  XNOR U17565 ( .A(n17110), .B(n17109), .Z(n17335) );
  XOR U17566 ( .A(n17336), .B(n17335), .Z(n17338) );
  XOR U17567 ( .A(n17337), .B(n17338), .Z(n17349) );
  NANDN U17568 ( .A(n17019), .B(n17018), .Z(n17023) );
  NANDN U17569 ( .A(n17021), .B(n17020), .Z(n17022) );
  AND U17570 ( .A(n17023), .B(n17022), .Z(n17347) );
  NANDN U17571 ( .A(n17025), .B(n17024), .Z(n17029) );
  OR U17572 ( .A(n17027), .B(n17026), .Z(n17028) );
  AND U17573 ( .A(n17029), .B(n17028), .Z(n17344) );
  NANDN U17574 ( .A(n17031), .B(n17030), .Z(n17035) );
  NAND U17575 ( .A(n17033), .B(n17032), .Z(n17034) );
  AND U17576 ( .A(n17035), .B(n17034), .Z(n17342) );
  NANDN U17577 ( .A(n17037), .B(n17036), .Z(n17041) );
  NANDN U17578 ( .A(n17039), .B(n17038), .Z(n17040) );
  AND U17579 ( .A(n17041), .B(n17040), .Z(n17341) );
  XNOR U17580 ( .A(n17342), .B(n17341), .Z(n17343) );
  XOR U17581 ( .A(n17344), .B(n17343), .Z(n17348) );
  XOR U17582 ( .A(n17347), .B(n17348), .Z(n17350) );
  XOR U17583 ( .A(n17349), .B(n17350), .Z(n17079) );
  NANDN U17584 ( .A(n17043), .B(n17042), .Z(n17047) );
  NANDN U17585 ( .A(n17045), .B(n17044), .Z(n17046) );
  AND U17586 ( .A(n17047), .B(n17046), .Z(n17078) );
  NANDN U17587 ( .A(n17049), .B(n17048), .Z(n17053) );
  OR U17588 ( .A(n17051), .B(n17050), .Z(n17052) );
  AND U17589 ( .A(n17053), .B(n17052), .Z(n17077) );
  XOR U17590 ( .A(n17078), .B(n17077), .Z(n17080) );
  XOR U17591 ( .A(n17079), .B(n17080), .Z(n17355) );
  NANDN U17592 ( .A(n17055), .B(n17054), .Z(n17059) );
  NANDN U17593 ( .A(n17057), .B(n17056), .Z(n17058) );
  AND U17594 ( .A(n17059), .B(n17058), .Z(n17354) );
  XNOR U17595 ( .A(n17355), .B(n17354), .Z(n17356) );
  NANDN U17596 ( .A(n17061), .B(n17060), .Z(n17065) );
  NAND U17597 ( .A(n17063), .B(n17062), .Z(n17064) );
  NAND U17598 ( .A(n17065), .B(n17064), .Z(n17357) );
  XNOR U17599 ( .A(n17356), .B(n17357), .Z(n17071) );
  XNOR U17600 ( .A(n17072), .B(n17071), .Z(n17073) );
  XNOR U17601 ( .A(n17074), .B(n17073), .Z(n17360) );
  XNOR U17602 ( .A(sreg[153]), .B(n17360), .Z(n17362) );
  NANDN U17603 ( .A(sreg[152]), .B(n17066), .Z(n17070) );
  NAND U17604 ( .A(n17068), .B(n17067), .Z(n17069) );
  NAND U17605 ( .A(n17070), .B(n17069), .Z(n17361) );
  XNOR U17606 ( .A(n17362), .B(n17361), .Z(c[153]) );
  NANDN U17607 ( .A(n17072), .B(n17071), .Z(n17076) );
  NANDN U17608 ( .A(n17074), .B(n17073), .Z(n17075) );
  AND U17609 ( .A(n17076), .B(n17075), .Z(n17368) );
  NANDN U17610 ( .A(n17078), .B(n17077), .Z(n17082) );
  OR U17611 ( .A(n17080), .B(n17079), .Z(n17081) );
  AND U17612 ( .A(n17082), .B(n17081), .Z(n17373) );
  NANDN U17613 ( .A(n17084), .B(n17083), .Z(n17088) );
  OR U17614 ( .A(n17086), .B(n17085), .Z(n17087) );
  AND U17615 ( .A(n17088), .B(n17087), .Z(n17634) );
  NANDN U17616 ( .A(n17090), .B(n17089), .Z(n17094) );
  NANDN U17617 ( .A(n17092), .B(n17091), .Z(n17093) );
  AND U17618 ( .A(n17094), .B(n17093), .Z(n17633) );
  NANDN U17619 ( .A(n17096), .B(n17095), .Z(n17100) );
  OR U17620 ( .A(n17098), .B(n17097), .Z(n17099) );
  AND U17621 ( .A(n17100), .B(n17099), .Z(n17632) );
  XOR U17622 ( .A(n17633), .B(n17632), .Z(n17635) );
  XOR U17623 ( .A(n17634), .B(n17635), .Z(n17639) );
  NANDN U17624 ( .A(n17102), .B(n17101), .Z(n17106) );
  NAND U17625 ( .A(n17104), .B(n17103), .Z(n17105) );
  AND U17626 ( .A(n17106), .B(n17105), .Z(n17638) );
  XNOR U17627 ( .A(n17639), .B(n17638), .Z(n17640) );
  NANDN U17628 ( .A(n17108), .B(n17107), .Z(n17112) );
  NANDN U17629 ( .A(n17110), .B(n17109), .Z(n17111) );
  AND U17630 ( .A(n17112), .B(n17111), .Z(n17629) );
  NANDN U17631 ( .A(n17114), .B(n17113), .Z(n17118) );
  NAND U17632 ( .A(n17116), .B(n17115), .Z(n17117) );
  AND U17633 ( .A(n17118), .B(n17117), .Z(n17394) );
  NANDN U17634 ( .A(n17120), .B(n17119), .Z(n17124) );
  NANDN U17635 ( .A(n17122), .B(n17121), .Z(n17123) );
  AND U17636 ( .A(n17124), .B(n17123), .Z(n17381) );
  NANDN U17637 ( .A(n211), .B(n17125), .Z(n17127) );
  XOR U17638 ( .A(b[47]), .B(a[44]), .Z(n17464) );
  NANDN U17639 ( .A(n37172), .B(n17464), .Z(n17126) );
  AND U17640 ( .A(n17127), .B(n17126), .Z(n17505) );
  NANDN U17641 ( .A(n210), .B(n17128), .Z(n17130) );
  XOR U17642 ( .A(a[82]), .B(b[9]), .Z(n17467) );
  NANDN U17643 ( .A(n30267), .B(n17467), .Z(n17129) );
  AND U17644 ( .A(n17130), .B(n17129), .Z(n17504) );
  NANDN U17645 ( .A(n212), .B(n17131), .Z(n17133) );
  XOR U17646 ( .A(b[49]), .B(a[42]), .Z(n17470) );
  NANDN U17647 ( .A(n37432), .B(n17470), .Z(n17132) );
  NAND U17648 ( .A(n17133), .B(n17132), .Z(n17503) );
  XOR U17649 ( .A(n17504), .B(n17503), .Z(n17506) );
  XOR U17650 ( .A(n17505), .B(n17506), .Z(n17528) );
  NANDN U17651 ( .A(n36742), .B(n17134), .Z(n17136) );
  XOR U17652 ( .A(b[43]), .B(a[48]), .Z(n17473) );
  NANDN U17653 ( .A(n36891), .B(n17473), .Z(n17135) );
  AND U17654 ( .A(n17136), .B(n17135), .Z(n17484) );
  NANDN U17655 ( .A(n36991), .B(n17137), .Z(n17139) );
  XOR U17656 ( .A(b[45]), .B(a[46]), .Z(n17476) );
  NANDN U17657 ( .A(n37083), .B(n17476), .Z(n17138) );
  AND U17658 ( .A(n17139), .B(n17138), .Z(n17483) );
  NANDN U17659 ( .A(n30482), .B(n17140), .Z(n17142) );
  XOR U17660 ( .A(a[80]), .B(b[11]), .Z(n17479) );
  NANDN U17661 ( .A(n30891), .B(n17479), .Z(n17141) );
  NAND U17662 ( .A(n17142), .B(n17141), .Z(n17482) );
  XOR U17663 ( .A(n17483), .B(n17482), .Z(n17485) );
  XNOR U17664 ( .A(n17484), .B(n17485), .Z(n17527) );
  XNOR U17665 ( .A(n17528), .B(n17527), .Z(n17529) );
  NANDN U17666 ( .A(n17144), .B(n17143), .Z(n17148) );
  OR U17667 ( .A(n17146), .B(n17145), .Z(n17147) );
  NAND U17668 ( .A(n17148), .B(n17147), .Z(n17530) );
  XNOR U17669 ( .A(n17529), .B(n17530), .Z(n17380) );
  XNOR U17670 ( .A(n17381), .B(n17380), .Z(n17383) );
  NANDN U17671 ( .A(n29499), .B(n17149), .Z(n17151) );
  XOR U17672 ( .A(a[84]), .B(b[7]), .Z(n17488) );
  NANDN U17673 ( .A(n29735), .B(n17488), .Z(n17150) );
  AND U17674 ( .A(n17151), .B(n17150), .Z(n17448) );
  NANDN U17675 ( .A(n37857), .B(n17152), .Z(n17154) );
  XOR U17676 ( .A(b[55]), .B(a[36]), .Z(n17491) );
  NANDN U17677 ( .A(n37911), .B(n17491), .Z(n17153) );
  AND U17678 ( .A(n17154), .B(n17153), .Z(n17447) );
  NANDN U17679 ( .A(n35611), .B(n17155), .Z(n17157) );
  XOR U17680 ( .A(b[35]), .B(a[56]), .Z(n17494) );
  NANDN U17681 ( .A(n35801), .B(n17494), .Z(n17156) );
  NAND U17682 ( .A(n17157), .B(n17156), .Z(n17446) );
  XOR U17683 ( .A(n17447), .B(n17446), .Z(n17449) );
  XOR U17684 ( .A(n17448), .B(n17449), .Z(n17510) );
  NANDN U17685 ( .A(n17159), .B(n17158), .Z(n17163) );
  OR U17686 ( .A(n17161), .B(n17160), .Z(n17162) );
  AND U17687 ( .A(n17163), .B(n17162), .Z(n17509) );
  XNOR U17688 ( .A(n17510), .B(n17509), .Z(n17511) );
  NANDN U17689 ( .A(n17165), .B(n17164), .Z(n17169) );
  OR U17690 ( .A(n17167), .B(n17166), .Z(n17168) );
  NAND U17691 ( .A(n17169), .B(n17168), .Z(n17512) );
  XNOR U17692 ( .A(n17511), .B(n17512), .Z(n17382) );
  XOR U17693 ( .A(n17383), .B(n17382), .Z(n17393) );
  NANDN U17694 ( .A(n17171), .B(n17170), .Z(n17175) );
  NANDN U17695 ( .A(n17173), .B(n17172), .Z(n17174) );
  AND U17696 ( .A(n17175), .B(n17174), .Z(n17389) );
  NANDN U17697 ( .A(n17177), .B(n17176), .Z(n17181) );
  NANDN U17698 ( .A(n17179), .B(n17178), .Z(n17180) );
  AND U17699 ( .A(n17181), .B(n17180), .Z(n17387) );
  NANDN U17700 ( .A(n33875), .B(n17182), .Z(n17184) );
  XOR U17701 ( .A(b[25]), .B(a[66]), .Z(n17422) );
  NANDN U17702 ( .A(n33994), .B(n17422), .Z(n17183) );
  AND U17703 ( .A(n17184), .B(n17183), .Z(n17550) );
  NANDN U17704 ( .A(n32013), .B(n17185), .Z(n17187) );
  XOR U17705 ( .A(b[17]), .B(a[74]), .Z(n17425) );
  NANDN U17706 ( .A(n32292), .B(n17425), .Z(n17186) );
  AND U17707 ( .A(n17187), .B(n17186), .Z(n17549) );
  NANDN U17708 ( .A(n31536), .B(n17188), .Z(n17190) );
  XOR U17709 ( .A(b[15]), .B(a[76]), .Z(n17428) );
  NANDN U17710 ( .A(n31925), .B(n17428), .Z(n17189) );
  NAND U17711 ( .A(n17190), .B(n17189), .Z(n17548) );
  XOR U17712 ( .A(n17549), .B(n17548), .Z(n17551) );
  XOR U17713 ( .A(n17550), .B(n17551), .Z(n17615) );
  NANDN U17714 ( .A(n37526), .B(n17191), .Z(n17193) );
  XOR U17715 ( .A(b[51]), .B(a[40]), .Z(n17431) );
  NANDN U17716 ( .A(n37605), .B(n17431), .Z(n17192) );
  AND U17717 ( .A(n17193), .B(n17192), .Z(n17574) );
  NANDN U17718 ( .A(n37705), .B(n17194), .Z(n17196) );
  XOR U17719 ( .A(b[53]), .B(a[38]), .Z(n17434) );
  NANDN U17720 ( .A(n37778), .B(n17434), .Z(n17195) );
  AND U17721 ( .A(n17196), .B(n17195), .Z(n17573) );
  NANDN U17722 ( .A(n36210), .B(n17197), .Z(n17199) );
  XOR U17723 ( .A(b[39]), .B(a[52]), .Z(n17437) );
  NANDN U17724 ( .A(n36347), .B(n17437), .Z(n17198) );
  NAND U17725 ( .A(n17199), .B(n17198), .Z(n17572) );
  XOR U17726 ( .A(n17573), .B(n17572), .Z(n17575) );
  XNOR U17727 ( .A(n17574), .B(n17575), .Z(n17614) );
  XNOR U17728 ( .A(n17615), .B(n17614), .Z(n17617) );
  NANDN U17729 ( .A(n17201), .B(n17200), .Z(n17205) );
  OR U17730 ( .A(n17203), .B(n17202), .Z(n17204) );
  AND U17731 ( .A(n17205), .B(n17204), .Z(n17616) );
  XOR U17732 ( .A(n17617), .B(n17616), .Z(n17413) );
  NANDN U17733 ( .A(n17207), .B(n17206), .Z(n17211) );
  OR U17734 ( .A(n17209), .B(n17208), .Z(n17210) );
  AND U17735 ( .A(n17211), .B(n17210), .Z(n17411) );
  NANDN U17736 ( .A(n17213), .B(n17212), .Z(n17217) );
  NANDN U17737 ( .A(n17215), .B(n17214), .Z(n17216) );
  NAND U17738 ( .A(n17217), .B(n17216), .Z(n17410) );
  XNOR U17739 ( .A(n17411), .B(n17410), .Z(n17412) );
  XNOR U17740 ( .A(n17413), .B(n17412), .Z(n17386) );
  XNOR U17741 ( .A(n17387), .B(n17386), .Z(n17388) );
  XNOR U17742 ( .A(n17389), .B(n17388), .Z(n17392) );
  XOR U17743 ( .A(n17393), .B(n17392), .Z(n17395) );
  XNOR U17744 ( .A(n17394), .B(n17395), .Z(n17626) );
  NANDN U17745 ( .A(n17219), .B(n17218), .Z(n17223) );
  NANDN U17746 ( .A(n17221), .B(n17220), .Z(n17222) );
  AND U17747 ( .A(n17223), .B(n17222), .Z(n17376) );
  NANDN U17748 ( .A(n17225), .B(n17224), .Z(n17229) );
  NANDN U17749 ( .A(n17227), .B(n17226), .Z(n17228) );
  AND U17750 ( .A(n17229), .B(n17228), .Z(n17375) );
  NANDN U17751 ( .A(n17231), .B(n17230), .Z(n17235) );
  NAND U17752 ( .A(n17233), .B(n17232), .Z(n17234) );
  AND U17753 ( .A(n17235), .B(n17234), .Z(n17374) );
  XOR U17754 ( .A(n17375), .B(n17374), .Z(n17377) );
  XOR U17755 ( .A(n17376), .B(n17377), .Z(n17401) );
  NANDN U17756 ( .A(n17237), .B(n17236), .Z(n17241) );
  NANDN U17757 ( .A(n17239), .B(n17238), .Z(n17240) );
  AND U17758 ( .A(n17241), .B(n17240), .Z(n17623) );
  NANDN U17759 ( .A(n32996), .B(n17242), .Z(n17244) );
  XOR U17760 ( .A(b[21]), .B(a[70]), .Z(n17533) );
  NANDN U17761 ( .A(n33271), .B(n17533), .Z(n17243) );
  AND U17762 ( .A(n17244), .B(n17243), .Z(n17592) );
  NANDN U17763 ( .A(n33866), .B(n17245), .Z(n17247) );
  XOR U17764 ( .A(b[23]), .B(a[68]), .Z(n17536) );
  NANDN U17765 ( .A(n33644), .B(n17536), .Z(n17246) );
  AND U17766 ( .A(n17247), .B(n17246), .Z(n17591) );
  NANDN U17767 ( .A(n32483), .B(n17248), .Z(n17250) );
  XOR U17768 ( .A(b[19]), .B(a[72]), .Z(n17539) );
  NANDN U17769 ( .A(n32823), .B(n17539), .Z(n17249) );
  NAND U17770 ( .A(n17250), .B(n17249), .Z(n17590) );
  XOR U17771 ( .A(n17591), .B(n17590), .Z(n17593) );
  XOR U17772 ( .A(n17592), .B(n17593), .Z(n17459) );
  NANDN U17773 ( .A(n34909), .B(n17251), .Z(n17253) );
  XOR U17774 ( .A(b[31]), .B(a[60]), .Z(n17542) );
  NANDN U17775 ( .A(n35145), .B(n17542), .Z(n17252) );
  AND U17776 ( .A(n17253), .B(n17252), .Z(n17499) );
  NANDN U17777 ( .A(n38247), .B(n17254), .Z(n17256) );
  XOR U17778 ( .A(b[61]), .B(a[30]), .Z(n17545) );
  NANDN U17779 ( .A(n38248), .B(n17545), .Z(n17255) );
  AND U17780 ( .A(n17256), .B(n17255), .Z(n17498) );
  AND U17781 ( .A(b[63]), .B(a[26]), .Z(n17497) );
  XOR U17782 ( .A(n17498), .B(n17497), .Z(n17500) );
  XNOR U17783 ( .A(n17499), .B(n17500), .Z(n17458) );
  XNOR U17784 ( .A(n17459), .B(n17458), .Z(n17460) );
  NANDN U17785 ( .A(n17258), .B(n17257), .Z(n17262) );
  OR U17786 ( .A(n17260), .B(n17259), .Z(n17261) );
  NAND U17787 ( .A(n17262), .B(n17261), .Z(n17461) );
  XNOR U17788 ( .A(n17460), .B(n17461), .Z(n17620) );
  NANDN U17789 ( .A(n34223), .B(n17263), .Z(n17265) );
  XOR U17790 ( .A(b[27]), .B(a[64]), .Z(n17554) );
  NANDN U17791 ( .A(n34458), .B(n17554), .Z(n17264) );
  AND U17792 ( .A(n17265), .B(n17264), .Z(n17442) );
  NANDN U17793 ( .A(n34634), .B(n17266), .Z(n17268) );
  XOR U17794 ( .A(b[29]), .B(a[62]), .Z(n17557) );
  NANDN U17795 ( .A(n34722), .B(n17557), .Z(n17267) );
  AND U17796 ( .A(n17268), .B(n17267), .Z(n17441) );
  NANDN U17797 ( .A(n31055), .B(n17269), .Z(n17271) );
  XOR U17798 ( .A(b[13]), .B(a[78]), .Z(n17560) );
  NANDN U17799 ( .A(n31293), .B(n17560), .Z(n17270) );
  NAND U17800 ( .A(n17271), .B(n17270), .Z(n17440) );
  XOR U17801 ( .A(n17441), .B(n17440), .Z(n17443) );
  XOR U17802 ( .A(n17442), .B(n17443), .Z(n17516) );
  NANDN U17803 ( .A(n28889), .B(n17272), .Z(n17274) );
  XOR U17804 ( .A(a[86]), .B(b[5]), .Z(n17563) );
  NANDN U17805 ( .A(n29138), .B(n17563), .Z(n17273) );
  AND U17806 ( .A(n17274), .B(n17273), .Z(n17586) );
  NANDN U17807 ( .A(n209), .B(n17275), .Z(n17277) );
  XOR U17808 ( .A(a[88]), .B(b[3]), .Z(n17566) );
  NANDN U17809 ( .A(n28941), .B(n17566), .Z(n17276) );
  AND U17810 ( .A(n17277), .B(n17276), .Z(n17585) );
  NANDN U17811 ( .A(n35936), .B(n17278), .Z(n17280) );
  XOR U17812 ( .A(b[37]), .B(a[54]), .Z(n17569) );
  NANDN U17813 ( .A(n36047), .B(n17569), .Z(n17279) );
  NAND U17814 ( .A(n17280), .B(n17279), .Z(n17584) );
  XOR U17815 ( .A(n17585), .B(n17584), .Z(n17587) );
  XNOR U17816 ( .A(n17586), .B(n17587), .Z(n17515) );
  XNOR U17817 ( .A(n17516), .B(n17515), .Z(n17517) );
  NANDN U17818 ( .A(n17282), .B(n17281), .Z(n17286) );
  OR U17819 ( .A(n17284), .B(n17283), .Z(n17285) );
  NAND U17820 ( .A(n17286), .B(n17285), .Z(n17518) );
  XOR U17821 ( .A(n17517), .B(n17518), .Z(n17621) );
  XNOR U17822 ( .A(n17620), .B(n17621), .Z(n17622) );
  XNOR U17823 ( .A(n17623), .B(n17622), .Z(n17407) );
  NANDN U17824 ( .A(n17288), .B(n17287), .Z(n17292) );
  NANDN U17825 ( .A(n17290), .B(n17289), .Z(n17291) );
  AND U17826 ( .A(n17292), .B(n17291), .Z(n17522) );
  NANDN U17827 ( .A(n17294), .B(n17293), .Z(n17298) );
  OR U17828 ( .A(n17296), .B(n17295), .Z(n17297) );
  NAND U17829 ( .A(n17298), .B(n17297), .Z(n17521) );
  XNOR U17830 ( .A(n17522), .B(n17521), .Z(n17524) );
  NANDN U17831 ( .A(n17300), .B(n17299), .Z(n17304) );
  OR U17832 ( .A(n17302), .B(n17301), .Z(n17303) );
  AND U17833 ( .A(n17304), .B(n17303), .Z(n17419) );
  NANDN U17834 ( .A(n38278), .B(n17305), .Z(n17307) );
  XOR U17835 ( .A(b[63]), .B(a[28]), .Z(n17599) );
  NANDN U17836 ( .A(n38279), .B(n17599), .Z(n17306) );
  AND U17837 ( .A(n17307), .B(n17306), .Z(n17453) );
  NANDN U17838 ( .A(n35260), .B(n17308), .Z(n17310) );
  XOR U17839 ( .A(b[33]), .B(a[58]), .Z(n17602) );
  NANDN U17840 ( .A(n35456), .B(n17602), .Z(n17309) );
  NAND U17841 ( .A(n17310), .B(n17309), .Z(n17452) );
  XNOR U17842 ( .A(n17453), .B(n17452), .Z(n17454) );
  NAND U17843 ( .A(b[0]), .B(a[90]), .Z(n17311) );
  XNOR U17844 ( .A(b[1]), .B(n17311), .Z(n17313) );
  NANDN U17845 ( .A(b[0]), .B(a[89]), .Z(n17312) );
  NAND U17846 ( .A(n17313), .B(n17312), .Z(n17455) );
  XNOR U17847 ( .A(n17454), .B(n17455), .Z(n17416) );
  NANDN U17848 ( .A(n37974), .B(n17314), .Z(n17316) );
  XOR U17849 ( .A(b[57]), .B(a[34]), .Z(n17605) );
  NANDN U17850 ( .A(n38031), .B(n17605), .Z(n17315) );
  AND U17851 ( .A(n17316), .B(n17315), .Z(n17581) );
  NANDN U17852 ( .A(n38090), .B(n17317), .Z(n17319) );
  XOR U17853 ( .A(b[59]), .B(a[32]), .Z(n17608) );
  NANDN U17854 ( .A(n38130), .B(n17608), .Z(n17318) );
  AND U17855 ( .A(n17319), .B(n17318), .Z(n17579) );
  NANDN U17856 ( .A(n36480), .B(n17320), .Z(n17322) );
  XOR U17857 ( .A(b[41]), .B(a[50]), .Z(n17611) );
  NANDN U17858 ( .A(n36594), .B(n17611), .Z(n17321) );
  NAND U17859 ( .A(n17322), .B(n17321), .Z(n17578) );
  XNOR U17860 ( .A(n17579), .B(n17578), .Z(n17580) );
  XOR U17861 ( .A(n17581), .B(n17580), .Z(n17417) );
  XNOR U17862 ( .A(n17416), .B(n17417), .Z(n17418) );
  XNOR U17863 ( .A(n17419), .B(n17418), .Z(n17523) );
  XOR U17864 ( .A(n17524), .B(n17523), .Z(n17405) );
  NANDN U17865 ( .A(n17324), .B(n17323), .Z(n17328) );
  NAND U17866 ( .A(n17326), .B(n17325), .Z(n17327) );
  NAND U17867 ( .A(n17328), .B(n17327), .Z(n17404) );
  XNOR U17868 ( .A(n17405), .B(n17404), .Z(n17406) );
  XOR U17869 ( .A(n17407), .B(n17406), .Z(n17399) );
  NANDN U17870 ( .A(n17330), .B(n17329), .Z(n17334) );
  NANDN U17871 ( .A(n17332), .B(n17331), .Z(n17333) );
  AND U17872 ( .A(n17334), .B(n17333), .Z(n17398) );
  XNOR U17873 ( .A(n17399), .B(n17398), .Z(n17400) );
  XOR U17874 ( .A(n17401), .B(n17400), .Z(n17627) );
  XNOR U17875 ( .A(n17626), .B(n17627), .Z(n17628) );
  XOR U17876 ( .A(n17629), .B(n17628), .Z(n17641) );
  XNOR U17877 ( .A(n17640), .B(n17641), .Z(n17646) );
  NANDN U17878 ( .A(n17336), .B(n17335), .Z(n17340) );
  OR U17879 ( .A(n17338), .B(n17337), .Z(n17339) );
  AND U17880 ( .A(n17340), .B(n17339), .Z(n17645) );
  NANDN U17881 ( .A(n17342), .B(n17341), .Z(n17346) );
  NANDN U17882 ( .A(n17344), .B(n17343), .Z(n17345) );
  AND U17883 ( .A(n17346), .B(n17345), .Z(n17644) );
  XOR U17884 ( .A(n17645), .B(n17644), .Z(n17647) );
  XNOR U17885 ( .A(n17646), .B(n17647), .Z(n17372) );
  NANDN U17886 ( .A(n17348), .B(n17347), .Z(n17352) );
  OR U17887 ( .A(n17350), .B(n17349), .Z(n17351) );
  NAND U17888 ( .A(n17352), .B(n17351), .Z(n17371) );
  XOR U17889 ( .A(n17372), .B(n17371), .Z(n17353) );
  XNOR U17890 ( .A(n17373), .B(n17353), .Z(n17365) );
  NANDN U17891 ( .A(n17355), .B(n17354), .Z(n17359) );
  NANDN U17892 ( .A(n17357), .B(n17356), .Z(n17358) );
  AND U17893 ( .A(n17359), .B(n17358), .Z(n17366) );
  XNOR U17894 ( .A(n17365), .B(n17366), .Z(n17367) );
  XNOR U17895 ( .A(n17368), .B(n17367), .Z(n17650) );
  XNOR U17896 ( .A(sreg[154]), .B(n17650), .Z(n17652) );
  NANDN U17897 ( .A(sreg[153]), .B(n17360), .Z(n17364) );
  NAND U17898 ( .A(n17362), .B(n17361), .Z(n17363) );
  NAND U17899 ( .A(n17364), .B(n17363), .Z(n17651) );
  XNOR U17900 ( .A(n17652), .B(n17651), .Z(c[154]) );
  NANDN U17901 ( .A(n17366), .B(n17365), .Z(n17370) );
  NANDN U17902 ( .A(n17368), .B(n17367), .Z(n17369) );
  AND U17903 ( .A(n17370), .B(n17369), .Z(n17658) );
  NANDN U17904 ( .A(n17375), .B(n17374), .Z(n17379) );
  OR U17905 ( .A(n17377), .B(n17376), .Z(n17378) );
  AND U17906 ( .A(n17379), .B(n17378), .Z(n17675) );
  NANDN U17907 ( .A(n17381), .B(n17380), .Z(n17385) );
  NAND U17908 ( .A(n17383), .B(n17382), .Z(n17384) );
  AND U17909 ( .A(n17385), .B(n17384), .Z(n17674) );
  NANDN U17910 ( .A(n17387), .B(n17386), .Z(n17391) );
  NANDN U17911 ( .A(n17389), .B(n17388), .Z(n17390) );
  AND U17912 ( .A(n17391), .B(n17390), .Z(n17673) );
  XOR U17913 ( .A(n17674), .B(n17673), .Z(n17676) );
  XOR U17914 ( .A(n17675), .B(n17676), .Z(n17932) );
  NANDN U17915 ( .A(n17393), .B(n17392), .Z(n17397) );
  NANDN U17916 ( .A(n17395), .B(n17394), .Z(n17396) );
  NAND U17917 ( .A(n17397), .B(n17396), .Z(n17931) );
  XNOR U17918 ( .A(n17932), .B(n17931), .Z(n17933) );
  NANDN U17919 ( .A(n17399), .B(n17398), .Z(n17403) );
  NANDN U17920 ( .A(n17401), .B(n17400), .Z(n17402) );
  AND U17921 ( .A(n17403), .B(n17402), .Z(n17670) );
  NANDN U17922 ( .A(n17405), .B(n17404), .Z(n17409) );
  NAND U17923 ( .A(n17407), .B(n17406), .Z(n17408) );
  AND U17924 ( .A(n17409), .B(n17408), .Z(n17699) );
  NANDN U17925 ( .A(n17411), .B(n17410), .Z(n17415) );
  NANDN U17926 ( .A(n17413), .B(n17412), .Z(n17414) );
  AND U17927 ( .A(n17415), .B(n17414), .Z(n17693) );
  NANDN U17928 ( .A(n17417), .B(n17416), .Z(n17421) );
  NANDN U17929 ( .A(n17419), .B(n17418), .Z(n17420) );
  AND U17930 ( .A(n17421), .B(n17420), .Z(n17692) );
  NANDN U17931 ( .A(n33875), .B(n17422), .Z(n17424) );
  XOR U17932 ( .A(b[25]), .B(a[67]), .Z(n17727) );
  NANDN U17933 ( .A(n33994), .B(n17727), .Z(n17423) );
  AND U17934 ( .A(n17424), .B(n17423), .Z(n17897) );
  NANDN U17935 ( .A(n32013), .B(n17425), .Z(n17427) );
  XOR U17936 ( .A(b[17]), .B(a[75]), .Z(n17730) );
  NANDN U17937 ( .A(n32292), .B(n17730), .Z(n17426) );
  AND U17938 ( .A(n17427), .B(n17426), .Z(n17896) );
  NANDN U17939 ( .A(n31536), .B(n17428), .Z(n17430) );
  XOR U17940 ( .A(b[15]), .B(a[77]), .Z(n17733) );
  NANDN U17941 ( .A(n31925), .B(n17733), .Z(n17429) );
  NAND U17942 ( .A(n17430), .B(n17429), .Z(n17895) );
  XOR U17943 ( .A(n17896), .B(n17895), .Z(n17898) );
  XOR U17944 ( .A(n17897), .B(n17898), .Z(n17869) );
  NANDN U17945 ( .A(n37526), .B(n17431), .Z(n17433) );
  XOR U17946 ( .A(b[51]), .B(a[41]), .Z(n17736) );
  NANDN U17947 ( .A(n37605), .B(n17736), .Z(n17432) );
  AND U17948 ( .A(n17433), .B(n17432), .Z(n17921) );
  NANDN U17949 ( .A(n37705), .B(n17434), .Z(n17436) );
  XOR U17950 ( .A(b[53]), .B(a[39]), .Z(n17739) );
  NANDN U17951 ( .A(n37778), .B(n17739), .Z(n17435) );
  AND U17952 ( .A(n17436), .B(n17435), .Z(n17920) );
  NANDN U17953 ( .A(n36210), .B(n17437), .Z(n17439) );
  XOR U17954 ( .A(b[39]), .B(a[53]), .Z(n17742) );
  NANDN U17955 ( .A(n36347), .B(n17742), .Z(n17438) );
  NAND U17956 ( .A(n17439), .B(n17438), .Z(n17919) );
  XOR U17957 ( .A(n17920), .B(n17919), .Z(n17922) );
  XNOR U17958 ( .A(n17921), .B(n17922), .Z(n17868) );
  XNOR U17959 ( .A(n17869), .B(n17868), .Z(n17871) );
  NANDN U17960 ( .A(n17441), .B(n17440), .Z(n17445) );
  OR U17961 ( .A(n17443), .B(n17442), .Z(n17444) );
  AND U17962 ( .A(n17445), .B(n17444), .Z(n17870) );
  XOR U17963 ( .A(n17871), .B(n17870), .Z(n17718) );
  NANDN U17964 ( .A(n17447), .B(n17446), .Z(n17451) );
  OR U17965 ( .A(n17449), .B(n17448), .Z(n17450) );
  AND U17966 ( .A(n17451), .B(n17450), .Z(n17716) );
  NANDN U17967 ( .A(n17453), .B(n17452), .Z(n17457) );
  NANDN U17968 ( .A(n17455), .B(n17454), .Z(n17456) );
  NAND U17969 ( .A(n17457), .B(n17456), .Z(n17715) );
  XNOR U17970 ( .A(n17716), .B(n17715), .Z(n17717) );
  XNOR U17971 ( .A(n17718), .B(n17717), .Z(n17691) );
  XOR U17972 ( .A(n17692), .B(n17691), .Z(n17694) );
  XOR U17973 ( .A(n17693), .B(n17694), .Z(n17698) );
  NANDN U17974 ( .A(n17459), .B(n17458), .Z(n17463) );
  NANDN U17975 ( .A(n17461), .B(n17460), .Z(n17462) );
  AND U17976 ( .A(n17463), .B(n17462), .Z(n17686) );
  NANDN U17977 ( .A(n211), .B(n17464), .Z(n17466) );
  XOR U17978 ( .A(b[47]), .B(a[45]), .Z(n17790) );
  NANDN U17979 ( .A(n37172), .B(n17790), .Z(n17465) );
  AND U17980 ( .A(n17466), .B(n17465), .Z(n17780) );
  NANDN U17981 ( .A(n210), .B(n17467), .Z(n17469) );
  XOR U17982 ( .A(a[83]), .B(b[9]), .Z(n17793) );
  NANDN U17983 ( .A(n30267), .B(n17793), .Z(n17468) );
  AND U17984 ( .A(n17469), .B(n17468), .Z(n17779) );
  NANDN U17985 ( .A(n212), .B(n17470), .Z(n17472) );
  XOR U17986 ( .A(b[49]), .B(a[43]), .Z(n17796) );
  NANDN U17987 ( .A(n37432), .B(n17796), .Z(n17471) );
  NAND U17988 ( .A(n17472), .B(n17471), .Z(n17778) );
  XOR U17989 ( .A(n17779), .B(n17778), .Z(n17781) );
  XOR U17990 ( .A(n17780), .B(n17781), .Z(n17875) );
  NANDN U17991 ( .A(n36742), .B(n17473), .Z(n17475) );
  XOR U17992 ( .A(b[43]), .B(a[49]), .Z(n17799) );
  NANDN U17993 ( .A(n36891), .B(n17799), .Z(n17474) );
  AND U17994 ( .A(n17475), .B(n17474), .Z(n17810) );
  NANDN U17995 ( .A(n36991), .B(n17476), .Z(n17478) );
  XOR U17996 ( .A(b[45]), .B(a[47]), .Z(n17802) );
  NANDN U17997 ( .A(n37083), .B(n17802), .Z(n17477) );
  AND U17998 ( .A(n17478), .B(n17477), .Z(n17809) );
  NANDN U17999 ( .A(n30482), .B(n17479), .Z(n17481) );
  XOR U18000 ( .A(a[81]), .B(b[11]), .Z(n17805) );
  NANDN U18001 ( .A(n30891), .B(n17805), .Z(n17480) );
  NAND U18002 ( .A(n17481), .B(n17480), .Z(n17808) );
  XOR U18003 ( .A(n17809), .B(n17808), .Z(n17811) );
  XNOR U18004 ( .A(n17810), .B(n17811), .Z(n17874) );
  XNOR U18005 ( .A(n17875), .B(n17874), .Z(n17876) );
  NANDN U18006 ( .A(n17483), .B(n17482), .Z(n17487) );
  OR U18007 ( .A(n17485), .B(n17484), .Z(n17486) );
  NAND U18008 ( .A(n17487), .B(n17486), .Z(n17877) );
  XNOR U18009 ( .A(n17876), .B(n17877), .Z(n17685) );
  XNOR U18010 ( .A(n17686), .B(n17685), .Z(n17687) );
  NANDN U18011 ( .A(n29499), .B(n17488), .Z(n17490) );
  XOR U18012 ( .A(a[85]), .B(b[7]), .Z(n17763) );
  NANDN U18013 ( .A(n29735), .B(n17763), .Z(n17489) );
  AND U18014 ( .A(n17490), .B(n17489), .Z(n17753) );
  NANDN U18015 ( .A(n37857), .B(n17491), .Z(n17493) );
  XOR U18016 ( .A(b[55]), .B(a[37]), .Z(n17766) );
  NANDN U18017 ( .A(n37911), .B(n17766), .Z(n17492) );
  AND U18018 ( .A(n17493), .B(n17492), .Z(n17752) );
  NANDN U18019 ( .A(n35611), .B(n17494), .Z(n17496) );
  XOR U18020 ( .A(b[35]), .B(a[57]), .Z(n17769) );
  NANDN U18021 ( .A(n35801), .B(n17769), .Z(n17495) );
  NAND U18022 ( .A(n17496), .B(n17495), .Z(n17751) );
  XOR U18023 ( .A(n17752), .B(n17751), .Z(n17754) );
  XOR U18024 ( .A(n17753), .B(n17754), .Z(n17815) );
  NANDN U18025 ( .A(n17498), .B(n17497), .Z(n17502) );
  OR U18026 ( .A(n17500), .B(n17499), .Z(n17501) );
  AND U18027 ( .A(n17502), .B(n17501), .Z(n17814) );
  XNOR U18028 ( .A(n17815), .B(n17814), .Z(n17816) );
  NANDN U18029 ( .A(n17504), .B(n17503), .Z(n17508) );
  OR U18030 ( .A(n17506), .B(n17505), .Z(n17507) );
  NAND U18031 ( .A(n17508), .B(n17507), .Z(n17817) );
  XOR U18032 ( .A(n17816), .B(n17817), .Z(n17688) );
  XNOR U18033 ( .A(n17687), .B(n17688), .Z(n17697) );
  XOR U18034 ( .A(n17698), .B(n17697), .Z(n17700) );
  XOR U18035 ( .A(n17699), .B(n17700), .Z(n17668) );
  NANDN U18036 ( .A(n17510), .B(n17509), .Z(n17514) );
  NANDN U18037 ( .A(n17512), .B(n17511), .Z(n17513) );
  AND U18038 ( .A(n17514), .B(n17513), .Z(n17681) );
  NANDN U18039 ( .A(n17516), .B(n17515), .Z(n17520) );
  NANDN U18040 ( .A(n17518), .B(n17517), .Z(n17519) );
  AND U18041 ( .A(n17520), .B(n17519), .Z(n17680) );
  NANDN U18042 ( .A(n17522), .B(n17521), .Z(n17526) );
  NAND U18043 ( .A(n17524), .B(n17523), .Z(n17525) );
  AND U18044 ( .A(n17526), .B(n17525), .Z(n17679) );
  XOR U18045 ( .A(n17680), .B(n17679), .Z(n17682) );
  XOR U18046 ( .A(n17681), .B(n17682), .Z(n17706) );
  NANDN U18047 ( .A(n17528), .B(n17527), .Z(n17532) );
  NANDN U18048 ( .A(n17530), .B(n17529), .Z(n17531) );
  AND U18049 ( .A(n17532), .B(n17531), .Z(n17928) );
  NANDN U18050 ( .A(n32996), .B(n17533), .Z(n17535) );
  XOR U18051 ( .A(b[21]), .B(a[71]), .Z(n17880) );
  NANDN U18052 ( .A(n33271), .B(n17880), .Z(n17534) );
  AND U18053 ( .A(n17535), .B(n17534), .Z(n17846) );
  NANDN U18054 ( .A(n33866), .B(n17536), .Z(n17538) );
  XOR U18055 ( .A(b[23]), .B(a[69]), .Z(n17883) );
  NANDN U18056 ( .A(n33644), .B(n17883), .Z(n17537) );
  AND U18057 ( .A(n17538), .B(n17537), .Z(n17845) );
  NANDN U18058 ( .A(n32483), .B(n17539), .Z(n17541) );
  XOR U18059 ( .A(b[19]), .B(a[73]), .Z(n17886) );
  NANDN U18060 ( .A(n32823), .B(n17886), .Z(n17540) );
  NAND U18061 ( .A(n17541), .B(n17540), .Z(n17844) );
  XOR U18062 ( .A(n17845), .B(n17844), .Z(n17847) );
  XOR U18063 ( .A(n17846), .B(n17847), .Z(n17785) );
  NANDN U18064 ( .A(n34909), .B(n17542), .Z(n17544) );
  XOR U18065 ( .A(b[31]), .B(a[61]), .Z(n17889) );
  NANDN U18066 ( .A(n35145), .B(n17889), .Z(n17543) );
  AND U18067 ( .A(n17544), .B(n17543), .Z(n17774) );
  NANDN U18068 ( .A(n38247), .B(n17545), .Z(n17547) );
  XOR U18069 ( .A(b[61]), .B(a[31]), .Z(n17892) );
  NANDN U18070 ( .A(n38248), .B(n17892), .Z(n17546) );
  AND U18071 ( .A(n17547), .B(n17546), .Z(n17773) );
  AND U18072 ( .A(b[63]), .B(a[27]), .Z(n17772) );
  XOR U18073 ( .A(n17773), .B(n17772), .Z(n17775) );
  XNOR U18074 ( .A(n17774), .B(n17775), .Z(n17784) );
  XNOR U18075 ( .A(n17785), .B(n17784), .Z(n17786) );
  NANDN U18076 ( .A(n17549), .B(n17548), .Z(n17553) );
  OR U18077 ( .A(n17551), .B(n17550), .Z(n17552) );
  NAND U18078 ( .A(n17553), .B(n17552), .Z(n17787) );
  XNOR U18079 ( .A(n17786), .B(n17787), .Z(n17925) );
  NANDN U18080 ( .A(n34223), .B(n17554), .Z(n17556) );
  XOR U18081 ( .A(b[27]), .B(a[65]), .Z(n17901) );
  NANDN U18082 ( .A(n34458), .B(n17901), .Z(n17555) );
  AND U18083 ( .A(n17556), .B(n17555), .Z(n17747) );
  NANDN U18084 ( .A(n34634), .B(n17557), .Z(n17559) );
  XOR U18085 ( .A(b[29]), .B(a[63]), .Z(n17904) );
  NANDN U18086 ( .A(n34722), .B(n17904), .Z(n17558) );
  AND U18087 ( .A(n17559), .B(n17558), .Z(n17746) );
  NANDN U18088 ( .A(n31055), .B(n17560), .Z(n17562) );
  XOR U18089 ( .A(b[13]), .B(a[79]), .Z(n17907) );
  NANDN U18090 ( .A(n31293), .B(n17907), .Z(n17561) );
  NAND U18091 ( .A(n17562), .B(n17561), .Z(n17745) );
  XOR U18092 ( .A(n17746), .B(n17745), .Z(n17748) );
  XOR U18093 ( .A(n17747), .B(n17748), .Z(n17821) );
  NANDN U18094 ( .A(n28889), .B(n17563), .Z(n17565) );
  XOR U18095 ( .A(a[87]), .B(b[5]), .Z(n17910) );
  NANDN U18096 ( .A(n29138), .B(n17910), .Z(n17564) );
  AND U18097 ( .A(n17565), .B(n17564), .Z(n17840) );
  NANDN U18098 ( .A(n209), .B(n17566), .Z(n17568) );
  XOR U18099 ( .A(a[89]), .B(b[3]), .Z(n17913) );
  NANDN U18100 ( .A(n28941), .B(n17913), .Z(n17567) );
  AND U18101 ( .A(n17568), .B(n17567), .Z(n17839) );
  NANDN U18102 ( .A(n35936), .B(n17569), .Z(n17571) );
  XOR U18103 ( .A(b[37]), .B(a[55]), .Z(n17916) );
  NANDN U18104 ( .A(n36047), .B(n17916), .Z(n17570) );
  NAND U18105 ( .A(n17571), .B(n17570), .Z(n17838) );
  XOR U18106 ( .A(n17839), .B(n17838), .Z(n17841) );
  XNOR U18107 ( .A(n17840), .B(n17841), .Z(n17820) );
  XNOR U18108 ( .A(n17821), .B(n17820), .Z(n17822) );
  NANDN U18109 ( .A(n17573), .B(n17572), .Z(n17577) );
  OR U18110 ( .A(n17575), .B(n17574), .Z(n17576) );
  NAND U18111 ( .A(n17577), .B(n17576), .Z(n17823) );
  XOR U18112 ( .A(n17822), .B(n17823), .Z(n17926) );
  XNOR U18113 ( .A(n17925), .B(n17926), .Z(n17927) );
  XNOR U18114 ( .A(n17928), .B(n17927), .Z(n17712) );
  NANDN U18115 ( .A(n17579), .B(n17578), .Z(n17583) );
  NANDN U18116 ( .A(n17581), .B(n17580), .Z(n17582) );
  AND U18117 ( .A(n17583), .B(n17582), .Z(n17827) );
  NANDN U18118 ( .A(n17585), .B(n17584), .Z(n17589) );
  OR U18119 ( .A(n17587), .B(n17586), .Z(n17588) );
  NAND U18120 ( .A(n17589), .B(n17588), .Z(n17826) );
  XNOR U18121 ( .A(n17827), .B(n17826), .Z(n17829) );
  NANDN U18122 ( .A(n17591), .B(n17590), .Z(n17595) );
  OR U18123 ( .A(n17593), .B(n17592), .Z(n17594) );
  AND U18124 ( .A(n17595), .B(n17594), .Z(n17724) );
  NAND U18125 ( .A(b[0]), .B(a[91]), .Z(n17596) );
  XNOR U18126 ( .A(b[1]), .B(n17596), .Z(n17598) );
  NANDN U18127 ( .A(b[0]), .B(a[90]), .Z(n17597) );
  NAND U18128 ( .A(n17598), .B(n17597), .Z(n17760) );
  NANDN U18129 ( .A(n38278), .B(n17599), .Z(n17601) );
  XOR U18130 ( .A(b[63]), .B(a[29]), .Z(n17853) );
  NANDN U18131 ( .A(n38279), .B(n17853), .Z(n17600) );
  AND U18132 ( .A(n17601), .B(n17600), .Z(n17758) );
  NANDN U18133 ( .A(n35260), .B(n17602), .Z(n17604) );
  XOR U18134 ( .A(b[33]), .B(a[59]), .Z(n17856) );
  NANDN U18135 ( .A(n35456), .B(n17856), .Z(n17603) );
  NAND U18136 ( .A(n17604), .B(n17603), .Z(n17757) );
  XNOR U18137 ( .A(n17758), .B(n17757), .Z(n17759) );
  XNOR U18138 ( .A(n17760), .B(n17759), .Z(n17721) );
  NANDN U18139 ( .A(n37974), .B(n17605), .Z(n17607) );
  XOR U18140 ( .A(b[57]), .B(a[35]), .Z(n17859) );
  NANDN U18141 ( .A(n38031), .B(n17859), .Z(n17606) );
  AND U18142 ( .A(n17607), .B(n17606), .Z(n17835) );
  NANDN U18143 ( .A(n38090), .B(n17608), .Z(n17610) );
  XOR U18144 ( .A(b[59]), .B(a[33]), .Z(n17862) );
  NANDN U18145 ( .A(n38130), .B(n17862), .Z(n17609) );
  AND U18146 ( .A(n17610), .B(n17609), .Z(n17833) );
  NANDN U18147 ( .A(n36480), .B(n17611), .Z(n17613) );
  XOR U18148 ( .A(b[41]), .B(a[51]), .Z(n17865) );
  NANDN U18149 ( .A(n36594), .B(n17865), .Z(n17612) );
  NAND U18150 ( .A(n17613), .B(n17612), .Z(n17832) );
  XNOR U18151 ( .A(n17833), .B(n17832), .Z(n17834) );
  XOR U18152 ( .A(n17835), .B(n17834), .Z(n17722) );
  XNOR U18153 ( .A(n17721), .B(n17722), .Z(n17723) );
  XNOR U18154 ( .A(n17724), .B(n17723), .Z(n17828) );
  XOR U18155 ( .A(n17829), .B(n17828), .Z(n17710) );
  NANDN U18156 ( .A(n17615), .B(n17614), .Z(n17619) );
  NAND U18157 ( .A(n17617), .B(n17616), .Z(n17618) );
  NAND U18158 ( .A(n17619), .B(n17618), .Z(n17709) );
  XNOR U18159 ( .A(n17710), .B(n17709), .Z(n17711) );
  XOR U18160 ( .A(n17712), .B(n17711), .Z(n17704) );
  NANDN U18161 ( .A(n17621), .B(n17620), .Z(n17625) );
  NANDN U18162 ( .A(n17623), .B(n17622), .Z(n17624) );
  AND U18163 ( .A(n17625), .B(n17624), .Z(n17703) );
  XNOR U18164 ( .A(n17704), .B(n17703), .Z(n17705) );
  XNOR U18165 ( .A(n17706), .B(n17705), .Z(n17667) );
  XNOR U18166 ( .A(n17668), .B(n17667), .Z(n17669) );
  XOR U18167 ( .A(n17670), .B(n17669), .Z(n17934) );
  XNOR U18168 ( .A(n17933), .B(n17934), .Z(n17940) );
  NANDN U18169 ( .A(n17627), .B(n17626), .Z(n17631) );
  NANDN U18170 ( .A(n17629), .B(n17628), .Z(n17630) );
  AND U18171 ( .A(n17631), .B(n17630), .Z(n17938) );
  NANDN U18172 ( .A(n17633), .B(n17632), .Z(n17637) );
  OR U18173 ( .A(n17635), .B(n17634), .Z(n17636) );
  AND U18174 ( .A(n17637), .B(n17636), .Z(n17937) );
  XNOR U18175 ( .A(n17938), .B(n17937), .Z(n17939) );
  XOR U18176 ( .A(n17940), .B(n17939), .Z(n17662) );
  NANDN U18177 ( .A(n17639), .B(n17638), .Z(n17643) );
  NANDN U18178 ( .A(n17641), .B(n17640), .Z(n17642) );
  AND U18179 ( .A(n17643), .B(n17642), .Z(n17661) );
  XNOR U18180 ( .A(n17662), .B(n17661), .Z(n17663) );
  NANDN U18181 ( .A(n17645), .B(n17644), .Z(n17649) );
  NANDN U18182 ( .A(n17647), .B(n17646), .Z(n17648) );
  NAND U18183 ( .A(n17649), .B(n17648), .Z(n17664) );
  XNOR U18184 ( .A(n17663), .B(n17664), .Z(n17655) );
  XNOR U18185 ( .A(n17656), .B(n17655), .Z(n17657) );
  XNOR U18186 ( .A(n17658), .B(n17657), .Z(n17943) );
  XNOR U18187 ( .A(sreg[155]), .B(n17943), .Z(n17945) );
  NANDN U18188 ( .A(sreg[154]), .B(n17650), .Z(n17654) );
  NAND U18189 ( .A(n17652), .B(n17651), .Z(n17653) );
  NAND U18190 ( .A(n17654), .B(n17653), .Z(n17944) );
  XNOR U18191 ( .A(n17945), .B(n17944), .Z(c[155]) );
  NANDN U18192 ( .A(n17656), .B(n17655), .Z(n17660) );
  NANDN U18193 ( .A(n17658), .B(n17657), .Z(n17659) );
  AND U18194 ( .A(n17660), .B(n17659), .Z(n17951) );
  NANDN U18195 ( .A(n17662), .B(n17661), .Z(n17666) );
  NANDN U18196 ( .A(n17664), .B(n17663), .Z(n17665) );
  AND U18197 ( .A(n17666), .B(n17665), .Z(n17949) );
  NANDN U18198 ( .A(n17668), .B(n17667), .Z(n17672) );
  NANDN U18199 ( .A(n17670), .B(n17669), .Z(n17671) );
  AND U18200 ( .A(n17672), .B(n17671), .Z(n18231) );
  NANDN U18201 ( .A(n17674), .B(n17673), .Z(n17678) );
  OR U18202 ( .A(n17676), .B(n17675), .Z(n17677) );
  AND U18203 ( .A(n17678), .B(n17677), .Z(n18230) );
  XNOR U18204 ( .A(n18231), .B(n18230), .Z(n18233) );
  NANDN U18205 ( .A(n17680), .B(n17679), .Z(n17684) );
  OR U18206 ( .A(n17682), .B(n17681), .Z(n17683) );
  AND U18207 ( .A(n17684), .B(n17683), .Z(n17968) );
  NANDN U18208 ( .A(n17686), .B(n17685), .Z(n17690) );
  NANDN U18209 ( .A(n17688), .B(n17687), .Z(n17689) );
  AND U18210 ( .A(n17690), .B(n17689), .Z(n17967) );
  NANDN U18211 ( .A(n17692), .B(n17691), .Z(n17696) );
  OR U18212 ( .A(n17694), .B(n17693), .Z(n17695) );
  AND U18213 ( .A(n17696), .B(n17695), .Z(n17966) );
  XOR U18214 ( .A(n17967), .B(n17966), .Z(n17969) );
  XOR U18215 ( .A(n17968), .B(n17969), .Z(n18225) );
  NANDN U18216 ( .A(n17698), .B(n17697), .Z(n17702) );
  OR U18217 ( .A(n17700), .B(n17699), .Z(n17701) );
  AND U18218 ( .A(n17702), .B(n17701), .Z(n18224) );
  XNOR U18219 ( .A(n18225), .B(n18224), .Z(n18226) );
  NANDN U18220 ( .A(n17704), .B(n17703), .Z(n17708) );
  NANDN U18221 ( .A(n17706), .B(n17705), .Z(n17707) );
  AND U18222 ( .A(n17708), .B(n17707), .Z(n17963) );
  NANDN U18223 ( .A(n17710), .B(n17709), .Z(n17714) );
  NAND U18224 ( .A(n17712), .B(n17711), .Z(n17713) );
  AND U18225 ( .A(n17714), .B(n17713), .Z(n17992) );
  NANDN U18226 ( .A(n17716), .B(n17715), .Z(n17720) );
  NANDN U18227 ( .A(n17718), .B(n17717), .Z(n17719) );
  AND U18228 ( .A(n17720), .B(n17719), .Z(n17986) );
  NANDN U18229 ( .A(n17722), .B(n17721), .Z(n17726) );
  NANDN U18230 ( .A(n17724), .B(n17723), .Z(n17725) );
  AND U18231 ( .A(n17726), .B(n17725), .Z(n17985) );
  NANDN U18232 ( .A(n33875), .B(n17727), .Z(n17729) );
  XOR U18233 ( .A(b[25]), .B(a[68]), .Z(n18020) );
  NANDN U18234 ( .A(n33994), .B(n18020), .Z(n17728) );
  AND U18235 ( .A(n17729), .B(n17728), .Z(n18190) );
  NANDN U18236 ( .A(n32013), .B(n17730), .Z(n17732) );
  XOR U18237 ( .A(b[17]), .B(a[76]), .Z(n18023) );
  NANDN U18238 ( .A(n32292), .B(n18023), .Z(n17731) );
  AND U18239 ( .A(n17732), .B(n17731), .Z(n18189) );
  NANDN U18240 ( .A(n31536), .B(n17733), .Z(n17735) );
  XOR U18241 ( .A(b[15]), .B(a[78]), .Z(n18026) );
  NANDN U18242 ( .A(n31925), .B(n18026), .Z(n17734) );
  NAND U18243 ( .A(n17735), .B(n17734), .Z(n18188) );
  XOR U18244 ( .A(n18189), .B(n18188), .Z(n18191) );
  XOR U18245 ( .A(n18190), .B(n18191), .Z(n18162) );
  NANDN U18246 ( .A(n37526), .B(n17736), .Z(n17738) );
  XOR U18247 ( .A(b[51]), .B(a[42]), .Z(n18029) );
  NANDN U18248 ( .A(n37605), .B(n18029), .Z(n17737) );
  AND U18249 ( .A(n17738), .B(n17737), .Z(n18214) );
  NANDN U18250 ( .A(n37705), .B(n17739), .Z(n17741) );
  XOR U18251 ( .A(b[53]), .B(a[40]), .Z(n18032) );
  NANDN U18252 ( .A(n37778), .B(n18032), .Z(n17740) );
  AND U18253 ( .A(n17741), .B(n17740), .Z(n18213) );
  NANDN U18254 ( .A(n36210), .B(n17742), .Z(n17744) );
  XOR U18255 ( .A(b[39]), .B(a[54]), .Z(n18035) );
  NANDN U18256 ( .A(n36347), .B(n18035), .Z(n17743) );
  NAND U18257 ( .A(n17744), .B(n17743), .Z(n18212) );
  XOR U18258 ( .A(n18213), .B(n18212), .Z(n18215) );
  XNOR U18259 ( .A(n18214), .B(n18215), .Z(n18161) );
  XNOR U18260 ( .A(n18162), .B(n18161), .Z(n18164) );
  NANDN U18261 ( .A(n17746), .B(n17745), .Z(n17750) );
  OR U18262 ( .A(n17748), .B(n17747), .Z(n17749) );
  AND U18263 ( .A(n17750), .B(n17749), .Z(n18163) );
  XOR U18264 ( .A(n18164), .B(n18163), .Z(n18011) );
  NANDN U18265 ( .A(n17752), .B(n17751), .Z(n17756) );
  OR U18266 ( .A(n17754), .B(n17753), .Z(n17755) );
  AND U18267 ( .A(n17756), .B(n17755), .Z(n18009) );
  NANDN U18268 ( .A(n17758), .B(n17757), .Z(n17762) );
  NANDN U18269 ( .A(n17760), .B(n17759), .Z(n17761) );
  NAND U18270 ( .A(n17762), .B(n17761), .Z(n18008) );
  XNOR U18271 ( .A(n18009), .B(n18008), .Z(n18010) );
  XNOR U18272 ( .A(n18011), .B(n18010), .Z(n17984) );
  XOR U18273 ( .A(n17985), .B(n17984), .Z(n17987) );
  XOR U18274 ( .A(n17986), .B(n17987), .Z(n17991) );
  NANDN U18275 ( .A(n29499), .B(n17763), .Z(n17765) );
  XOR U18276 ( .A(a[86]), .B(b[7]), .Z(n18086) );
  NANDN U18277 ( .A(n29735), .B(n18086), .Z(n17764) );
  AND U18278 ( .A(n17765), .B(n17764), .Z(n18046) );
  NANDN U18279 ( .A(n37857), .B(n17766), .Z(n17768) );
  XOR U18280 ( .A(b[55]), .B(a[38]), .Z(n18089) );
  NANDN U18281 ( .A(n37911), .B(n18089), .Z(n17767) );
  AND U18282 ( .A(n17768), .B(n17767), .Z(n18045) );
  NANDN U18283 ( .A(n35611), .B(n17769), .Z(n17771) );
  XOR U18284 ( .A(b[35]), .B(a[58]), .Z(n18092) );
  NANDN U18285 ( .A(n35801), .B(n18092), .Z(n17770) );
  NAND U18286 ( .A(n17771), .B(n17770), .Z(n18044) );
  XOR U18287 ( .A(n18045), .B(n18044), .Z(n18047) );
  XOR U18288 ( .A(n18046), .B(n18047), .Z(n18108) );
  NANDN U18289 ( .A(n17773), .B(n17772), .Z(n17777) );
  OR U18290 ( .A(n17775), .B(n17774), .Z(n17776) );
  AND U18291 ( .A(n17777), .B(n17776), .Z(n18107) );
  XNOR U18292 ( .A(n18108), .B(n18107), .Z(n18109) );
  NANDN U18293 ( .A(n17779), .B(n17778), .Z(n17783) );
  OR U18294 ( .A(n17781), .B(n17780), .Z(n17782) );
  NAND U18295 ( .A(n17783), .B(n17782), .Z(n18110) );
  XNOR U18296 ( .A(n18109), .B(n18110), .Z(n17980) );
  NANDN U18297 ( .A(n17785), .B(n17784), .Z(n17789) );
  NANDN U18298 ( .A(n17787), .B(n17786), .Z(n17788) );
  AND U18299 ( .A(n17789), .B(n17788), .Z(n17979) );
  NANDN U18300 ( .A(n211), .B(n17790), .Z(n17792) );
  XOR U18301 ( .A(b[47]), .B(a[46]), .Z(n18062) );
  NANDN U18302 ( .A(n37172), .B(n18062), .Z(n17791) );
  AND U18303 ( .A(n17792), .B(n17791), .Z(n18103) );
  NANDN U18304 ( .A(n210), .B(n17793), .Z(n17795) );
  XOR U18305 ( .A(a[84]), .B(b[9]), .Z(n18065) );
  NANDN U18306 ( .A(n30267), .B(n18065), .Z(n17794) );
  AND U18307 ( .A(n17795), .B(n17794), .Z(n18102) );
  NANDN U18308 ( .A(n212), .B(n17796), .Z(n17798) );
  XOR U18309 ( .A(b[49]), .B(a[44]), .Z(n18068) );
  NANDN U18310 ( .A(n37432), .B(n18068), .Z(n17797) );
  NAND U18311 ( .A(n17798), .B(n17797), .Z(n18101) );
  XOR U18312 ( .A(n18102), .B(n18101), .Z(n18104) );
  XOR U18313 ( .A(n18103), .B(n18104), .Z(n18168) );
  NANDN U18314 ( .A(n36742), .B(n17799), .Z(n17801) );
  XOR U18315 ( .A(b[43]), .B(a[50]), .Z(n18071) );
  NANDN U18316 ( .A(n36891), .B(n18071), .Z(n17800) );
  AND U18317 ( .A(n17801), .B(n17800), .Z(n18082) );
  NANDN U18318 ( .A(n36991), .B(n17802), .Z(n17804) );
  XOR U18319 ( .A(b[45]), .B(a[48]), .Z(n18074) );
  NANDN U18320 ( .A(n37083), .B(n18074), .Z(n17803) );
  AND U18321 ( .A(n17804), .B(n17803), .Z(n18081) );
  NANDN U18322 ( .A(n30482), .B(n17805), .Z(n17807) );
  XOR U18323 ( .A(a[82]), .B(b[11]), .Z(n18077) );
  NANDN U18324 ( .A(n30891), .B(n18077), .Z(n17806) );
  NAND U18325 ( .A(n17807), .B(n17806), .Z(n18080) );
  XOR U18326 ( .A(n18081), .B(n18080), .Z(n18083) );
  XNOR U18327 ( .A(n18082), .B(n18083), .Z(n18167) );
  XNOR U18328 ( .A(n18168), .B(n18167), .Z(n18169) );
  NANDN U18329 ( .A(n17809), .B(n17808), .Z(n17813) );
  OR U18330 ( .A(n17811), .B(n17810), .Z(n17812) );
  NAND U18331 ( .A(n17813), .B(n17812), .Z(n18170) );
  XNOR U18332 ( .A(n18169), .B(n18170), .Z(n17978) );
  XOR U18333 ( .A(n17979), .B(n17978), .Z(n17981) );
  XNOR U18334 ( .A(n17980), .B(n17981), .Z(n17990) );
  XOR U18335 ( .A(n17991), .B(n17990), .Z(n17993) );
  XOR U18336 ( .A(n17992), .B(n17993), .Z(n17961) );
  NANDN U18337 ( .A(n17815), .B(n17814), .Z(n17819) );
  NANDN U18338 ( .A(n17817), .B(n17816), .Z(n17818) );
  AND U18339 ( .A(n17819), .B(n17818), .Z(n17974) );
  NANDN U18340 ( .A(n17821), .B(n17820), .Z(n17825) );
  NANDN U18341 ( .A(n17823), .B(n17822), .Z(n17824) );
  AND U18342 ( .A(n17825), .B(n17824), .Z(n17973) );
  NANDN U18343 ( .A(n17827), .B(n17826), .Z(n17831) );
  NAND U18344 ( .A(n17829), .B(n17828), .Z(n17830) );
  AND U18345 ( .A(n17831), .B(n17830), .Z(n17972) );
  XOR U18346 ( .A(n17973), .B(n17972), .Z(n17975) );
  XOR U18347 ( .A(n17974), .B(n17975), .Z(n17999) );
  NANDN U18348 ( .A(n17833), .B(n17832), .Z(n17837) );
  NANDN U18349 ( .A(n17835), .B(n17834), .Z(n17836) );
  AND U18350 ( .A(n17837), .B(n17836), .Z(n18120) );
  NANDN U18351 ( .A(n17839), .B(n17838), .Z(n17843) );
  OR U18352 ( .A(n17841), .B(n17840), .Z(n17842) );
  NAND U18353 ( .A(n17843), .B(n17842), .Z(n18119) );
  XNOR U18354 ( .A(n18120), .B(n18119), .Z(n18122) );
  NANDN U18355 ( .A(n17845), .B(n17844), .Z(n17849) );
  OR U18356 ( .A(n17847), .B(n17846), .Z(n17848) );
  AND U18357 ( .A(n17849), .B(n17848), .Z(n18017) );
  NAND U18358 ( .A(b[0]), .B(a[92]), .Z(n17850) );
  XNOR U18359 ( .A(b[1]), .B(n17850), .Z(n17852) );
  NANDN U18360 ( .A(b[0]), .B(a[91]), .Z(n17851) );
  NAND U18361 ( .A(n17852), .B(n17851), .Z(n18053) );
  NANDN U18362 ( .A(n38278), .B(n17853), .Z(n17855) );
  XOR U18363 ( .A(b[63]), .B(a[30]), .Z(n18146) );
  NANDN U18364 ( .A(n38279), .B(n18146), .Z(n17854) );
  AND U18365 ( .A(n17855), .B(n17854), .Z(n18051) );
  NANDN U18366 ( .A(n35260), .B(n17856), .Z(n17858) );
  XOR U18367 ( .A(b[33]), .B(a[60]), .Z(n18149) );
  NANDN U18368 ( .A(n35456), .B(n18149), .Z(n17857) );
  NAND U18369 ( .A(n17858), .B(n17857), .Z(n18050) );
  XNOR U18370 ( .A(n18051), .B(n18050), .Z(n18052) );
  XNOR U18371 ( .A(n18053), .B(n18052), .Z(n18014) );
  NANDN U18372 ( .A(n37974), .B(n17859), .Z(n17861) );
  XOR U18373 ( .A(b[57]), .B(a[36]), .Z(n18152) );
  NANDN U18374 ( .A(n38031), .B(n18152), .Z(n17860) );
  AND U18375 ( .A(n17861), .B(n17860), .Z(n18128) );
  NANDN U18376 ( .A(n38090), .B(n17862), .Z(n17864) );
  XOR U18377 ( .A(b[59]), .B(a[34]), .Z(n18155) );
  NANDN U18378 ( .A(n38130), .B(n18155), .Z(n17863) );
  AND U18379 ( .A(n17864), .B(n17863), .Z(n18126) );
  NANDN U18380 ( .A(n36480), .B(n17865), .Z(n17867) );
  XOR U18381 ( .A(b[41]), .B(a[52]), .Z(n18158) );
  NANDN U18382 ( .A(n36594), .B(n18158), .Z(n17866) );
  NAND U18383 ( .A(n17867), .B(n17866), .Z(n18125) );
  XNOR U18384 ( .A(n18126), .B(n18125), .Z(n18127) );
  XOR U18385 ( .A(n18128), .B(n18127), .Z(n18015) );
  XNOR U18386 ( .A(n18014), .B(n18015), .Z(n18016) );
  XNOR U18387 ( .A(n18017), .B(n18016), .Z(n18121) );
  XOR U18388 ( .A(n18122), .B(n18121), .Z(n18003) );
  NANDN U18389 ( .A(n17869), .B(n17868), .Z(n17873) );
  NAND U18390 ( .A(n17871), .B(n17870), .Z(n17872) );
  NAND U18391 ( .A(n17873), .B(n17872), .Z(n18002) );
  XNOR U18392 ( .A(n18003), .B(n18002), .Z(n18005) );
  NANDN U18393 ( .A(n17875), .B(n17874), .Z(n17879) );
  NANDN U18394 ( .A(n17877), .B(n17876), .Z(n17878) );
  AND U18395 ( .A(n17879), .B(n17878), .Z(n18221) );
  NANDN U18396 ( .A(n32996), .B(n17880), .Z(n17882) );
  XOR U18397 ( .A(b[21]), .B(a[72]), .Z(n18173) );
  NANDN U18398 ( .A(n33271), .B(n18173), .Z(n17881) );
  AND U18399 ( .A(n17882), .B(n17881), .Z(n18139) );
  NANDN U18400 ( .A(n33866), .B(n17883), .Z(n17885) );
  XOR U18401 ( .A(b[23]), .B(a[70]), .Z(n18176) );
  NANDN U18402 ( .A(n33644), .B(n18176), .Z(n17884) );
  AND U18403 ( .A(n17885), .B(n17884), .Z(n18138) );
  NANDN U18404 ( .A(n32483), .B(n17886), .Z(n17888) );
  XOR U18405 ( .A(b[19]), .B(a[74]), .Z(n18179) );
  NANDN U18406 ( .A(n32823), .B(n18179), .Z(n17887) );
  NAND U18407 ( .A(n17888), .B(n17887), .Z(n18137) );
  XOR U18408 ( .A(n18138), .B(n18137), .Z(n18140) );
  XOR U18409 ( .A(n18139), .B(n18140), .Z(n18057) );
  NANDN U18410 ( .A(n34909), .B(n17889), .Z(n17891) );
  XOR U18411 ( .A(b[31]), .B(a[62]), .Z(n18182) );
  NANDN U18412 ( .A(n35145), .B(n18182), .Z(n17890) );
  AND U18413 ( .A(n17891), .B(n17890), .Z(n18097) );
  NANDN U18414 ( .A(n38247), .B(n17892), .Z(n17894) );
  XOR U18415 ( .A(b[61]), .B(a[32]), .Z(n18185) );
  NANDN U18416 ( .A(n38248), .B(n18185), .Z(n17893) );
  AND U18417 ( .A(n17894), .B(n17893), .Z(n18096) );
  AND U18418 ( .A(b[63]), .B(a[28]), .Z(n18095) );
  XOR U18419 ( .A(n18096), .B(n18095), .Z(n18098) );
  XNOR U18420 ( .A(n18097), .B(n18098), .Z(n18056) );
  XNOR U18421 ( .A(n18057), .B(n18056), .Z(n18058) );
  NANDN U18422 ( .A(n17896), .B(n17895), .Z(n17900) );
  OR U18423 ( .A(n17898), .B(n17897), .Z(n17899) );
  NAND U18424 ( .A(n17900), .B(n17899), .Z(n18059) );
  XNOR U18425 ( .A(n18058), .B(n18059), .Z(n18218) );
  NANDN U18426 ( .A(n34223), .B(n17901), .Z(n17903) );
  XOR U18427 ( .A(b[27]), .B(a[66]), .Z(n18194) );
  NANDN U18428 ( .A(n34458), .B(n18194), .Z(n17902) );
  AND U18429 ( .A(n17903), .B(n17902), .Z(n18040) );
  NANDN U18430 ( .A(n34634), .B(n17904), .Z(n17906) );
  XOR U18431 ( .A(b[29]), .B(a[64]), .Z(n18197) );
  NANDN U18432 ( .A(n34722), .B(n18197), .Z(n17905) );
  AND U18433 ( .A(n17906), .B(n17905), .Z(n18039) );
  NANDN U18434 ( .A(n31055), .B(n17907), .Z(n17909) );
  XOR U18435 ( .A(a[80]), .B(b[13]), .Z(n18200) );
  NANDN U18436 ( .A(n31293), .B(n18200), .Z(n17908) );
  NAND U18437 ( .A(n17909), .B(n17908), .Z(n18038) );
  XOR U18438 ( .A(n18039), .B(n18038), .Z(n18041) );
  XOR U18439 ( .A(n18040), .B(n18041), .Z(n18114) );
  NANDN U18440 ( .A(n28889), .B(n17910), .Z(n17912) );
  XOR U18441 ( .A(a[88]), .B(b[5]), .Z(n18203) );
  NANDN U18442 ( .A(n29138), .B(n18203), .Z(n17911) );
  AND U18443 ( .A(n17912), .B(n17911), .Z(n18133) );
  NANDN U18444 ( .A(n209), .B(n17913), .Z(n17915) );
  XOR U18445 ( .A(a[90]), .B(b[3]), .Z(n18206) );
  NANDN U18446 ( .A(n28941), .B(n18206), .Z(n17914) );
  AND U18447 ( .A(n17915), .B(n17914), .Z(n18132) );
  NANDN U18448 ( .A(n35936), .B(n17916), .Z(n17918) );
  XOR U18449 ( .A(b[37]), .B(a[56]), .Z(n18209) );
  NANDN U18450 ( .A(n36047), .B(n18209), .Z(n17917) );
  NAND U18451 ( .A(n17918), .B(n17917), .Z(n18131) );
  XOR U18452 ( .A(n18132), .B(n18131), .Z(n18134) );
  XNOR U18453 ( .A(n18133), .B(n18134), .Z(n18113) );
  XNOR U18454 ( .A(n18114), .B(n18113), .Z(n18115) );
  NANDN U18455 ( .A(n17920), .B(n17919), .Z(n17924) );
  OR U18456 ( .A(n17922), .B(n17921), .Z(n17923) );
  NAND U18457 ( .A(n17924), .B(n17923), .Z(n18116) );
  XOR U18458 ( .A(n18115), .B(n18116), .Z(n18219) );
  XNOR U18459 ( .A(n18218), .B(n18219), .Z(n18220) );
  XNOR U18460 ( .A(n18221), .B(n18220), .Z(n18004) );
  XOR U18461 ( .A(n18005), .B(n18004), .Z(n17997) );
  NANDN U18462 ( .A(n17926), .B(n17925), .Z(n17930) );
  NANDN U18463 ( .A(n17928), .B(n17927), .Z(n17929) );
  AND U18464 ( .A(n17930), .B(n17929), .Z(n17996) );
  XNOR U18465 ( .A(n17997), .B(n17996), .Z(n17998) );
  XNOR U18466 ( .A(n17999), .B(n17998), .Z(n17960) );
  XNOR U18467 ( .A(n17961), .B(n17960), .Z(n17962) );
  XOR U18468 ( .A(n17963), .B(n17962), .Z(n18227) );
  XNOR U18469 ( .A(n18226), .B(n18227), .Z(n18232) );
  XOR U18470 ( .A(n18233), .B(n18232), .Z(n17955) );
  NANDN U18471 ( .A(n17932), .B(n17931), .Z(n17936) );
  NANDN U18472 ( .A(n17934), .B(n17933), .Z(n17935) );
  AND U18473 ( .A(n17936), .B(n17935), .Z(n17954) );
  XNOR U18474 ( .A(n17955), .B(n17954), .Z(n17956) );
  NANDN U18475 ( .A(n17938), .B(n17937), .Z(n17942) );
  NAND U18476 ( .A(n17940), .B(n17939), .Z(n17941) );
  NAND U18477 ( .A(n17942), .B(n17941), .Z(n17957) );
  XNOR U18478 ( .A(n17956), .B(n17957), .Z(n17948) );
  XNOR U18479 ( .A(n17949), .B(n17948), .Z(n17950) );
  XNOR U18480 ( .A(n17951), .B(n17950), .Z(n18236) );
  XNOR U18481 ( .A(sreg[156]), .B(n18236), .Z(n18238) );
  NANDN U18482 ( .A(sreg[155]), .B(n17943), .Z(n17947) );
  NAND U18483 ( .A(n17945), .B(n17944), .Z(n17946) );
  NAND U18484 ( .A(n17947), .B(n17946), .Z(n18237) );
  XNOR U18485 ( .A(n18238), .B(n18237), .Z(c[156]) );
  NANDN U18486 ( .A(n17949), .B(n17948), .Z(n17953) );
  NANDN U18487 ( .A(n17951), .B(n17950), .Z(n17952) );
  AND U18488 ( .A(n17953), .B(n17952), .Z(n18244) );
  NANDN U18489 ( .A(n17955), .B(n17954), .Z(n17959) );
  NANDN U18490 ( .A(n17957), .B(n17956), .Z(n17958) );
  AND U18491 ( .A(n17959), .B(n17958), .Z(n18242) );
  NANDN U18492 ( .A(n17961), .B(n17960), .Z(n17965) );
  NANDN U18493 ( .A(n17963), .B(n17962), .Z(n17964) );
  AND U18494 ( .A(n17965), .B(n17964), .Z(n18524) );
  NANDN U18495 ( .A(n17967), .B(n17966), .Z(n17971) );
  OR U18496 ( .A(n17969), .B(n17968), .Z(n17970) );
  AND U18497 ( .A(n17971), .B(n17970), .Z(n18523) );
  XNOR U18498 ( .A(n18524), .B(n18523), .Z(n18526) );
  NANDN U18499 ( .A(n17973), .B(n17972), .Z(n17977) );
  OR U18500 ( .A(n17975), .B(n17974), .Z(n17976) );
  AND U18501 ( .A(n17977), .B(n17976), .Z(n18261) );
  NANDN U18502 ( .A(n17979), .B(n17978), .Z(n17983) );
  NANDN U18503 ( .A(n17981), .B(n17980), .Z(n17982) );
  AND U18504 ( .A(n17983), .B(n17982), .Z(n18260) );
  NANDN U18505 ( .A(n17985), .B(n17984), .Z(n17989) );
  OR U18506 ( .A(n17987), .B(n17986), .Z(n17988) );
  AND U18507 ( .A(n17989), .B(n17988), .Z(n18259) );
  XOR U18508 ( .A(n18260), .B(n18259), .Z(n18262) );
  XOR U18509 ( .A(n18261), .B(n18262), .Z(n18518) );
  NANDN U18510 ( .A(n17991), .B(n17990), .Z(n17995) );
  OR U18511 ( .A(n17993), .B(n17992), .Z(n17994) );
  AND U18512 ( .A(n17995), .B(n17994), .Z(n18517) );
  XNOR U18513 ( .A(n18518), .B(n18517), .Z(n18519) );
  NANDN U18514 ( .A(n17997), .B(n17996), .Z(n18001) );
  NANDN U18515 ( .A(n17999), .B(n17998), .Z(n18000) );
  AND U18516 ( .A(n18001), .B(n18000), .Z(n18256) );
  NANDN U18517 ( .A(n18003), .B(n18002), .Z(n18007) );
  NAND U18518 ( .A(n18005), .B(n18004), .Z(n18006) );
  AND U18519 ( .A(n18007), .B(n18006), .Z(n18285) );
  NANDN U18520 ( .A(n18009), .B(n18008), .Z(n18013) );
  NANDN U18521 ( .A(n18011), .B(n18010), .Z(n18012) );
  AND U18522 ( .A(n18013), .B(n18012), .Z(n18279) );
  NANDN U18523 ( .A(n18015), .B(n18014), .Z(n18019) );
  NANDN U18524 ( .A(n18017), .B(n18016), .Z(n18018) );
  AND U18525 ( .A(n18019), .B(n18018), .Z(n18278) );
  NANDN U18526 ( .A(n33875), .B(n18020), .Z(n18022) );
  XOR U18527 ( .A(b[25]), .B(a[69]), .Z(n18313) );
  NANDN U18528 ( .A(n33994), .B(n18313), .Z(n18021) );
  AND U18529 ( .A(n18022), .B(n18021), .Z(n18483) );
  NANDN U18530 ( .A(n32013), .B(n18023), .Z(n18025) );
  XOR U18531 ( .A(b[17]), .B(a[77]), .Z(n18316) );
  NANDN U18532 ( .A(n32292), .B(n18316), .Z(n18024) );
  AND U18533 ( .A(n18025), .B(n18024), .Z(n18482) );
  NANDN U18534 ( .A(n31536), .B(n18026), .Z(n18028) );
  XOR U18535 ( .A(b[15]), .B(a[79]), .Z(n18319) );
  NANDN U18536 ( .A(n31925), .B(n18319), .Z(n18027) );
  NAND U18537 ( .A(n18028), .B(n18027), .Z(n18481) );
  XOR U18538 ( .A(n18482), .B(n18481), .Z(n18484) );
  XOR U18539 ( .A(n18483), .B(n18484), .Z(n18455) );
  NANDN U18540 ( .A(n37526), .B(n18029), .Z(n18031) );
  XOR U18541 ( .A(b[51]), .B(a[43]), .Z(n18322) );
  NANDN U18542 ( .A(n37605), .B(n18322), .Z(n18030) );
  AND U18543 ( .A(n18031), .B(n18030), .Z(n18507) );
  NANDN U18544 ( .A(n37705), .B(n18032), .Z(n18034) );
  XOR U18545 ( .A(b[53]), .B(a[41]), .Z(n18325) );
  NANDN U18546 ( .A(n37778), .B(n18325), .Z(n18033) );
  AND U18547 ( .A(n18034), .B(n18033), .Z(n18506) );
  NANDN U18548 ( .A(n36210), .B(n18035), .Z(n18037) );
  XOR U18549 ( .A(b[39]), .B(a[55]), .Z(n18328) );
  NANDN U18550 ( .A(n36347), .B(n18328), .Z(n18036) );
  NAND U18551 ( .A(n18037), .B(n18036), .Z(n18505) );
  XOR U18552 ( .A(n18506), .B(n18505), .Z(n18508) );
  XNOR U18553 ( .A(n18507), .B(n18508), .Z(n18454) );
  XNOR U18554 ( .A(n18455), .B(n18454), .Z(n18457) );
  NANDN U18555 ( .A(n18039), .B(n18038), .Z(n18043) );
  OR U18556 ( .A(n18041), .B(n18040), .Z(n18042) );
  AND U18557 ( .A(n18043), .B(n18042), .Z(n18456) );
  XOR U18558 ( .A(n18457), .B(n18456), .Z(n18304) );
  NANDN U18559 ( .A(n18045), .B(n18044), .Z(n18049) );
  OR U18560 ( .A(n18047), .B(n18046), .Z(n18048) );
  AND U18561 ( .A(n18049), .B(n18048), .Z(n18302) );
  NANDN U18562 ( .A(n18051), .B(n18050), .Z(n18055) );
  NANDN U18563 ( .A(n18053), .B(n18052), .Z(n18054) );
  NAND U18564 ( .A(n18055), .B(n18054), .Z(n18301) );
  XNOR U18565 ( .A(n18302), .B(n18301), .Z(n18303) );
  XNOR U18566 ( .A(n18304), .B(n18303), .Z(n18277) );
  XOR U18567 ( .A(n18278), .B(n18277), .Z(n18280) );
  XOR U18568 ( .A(n18279), .B(n18280), .Z(n18284) );
  NANDN U18569 ( .A(n18057), .B(n18056), .Z(n18061) );
  NANDN U18570 ( .A(n18059), .B(n18058), .Z(n18060) );
  AND U18571 ( .A(n18061), .B(n18060), .Z(n18272) );
  NANDN U18572 ( .A(n211), .B(n18062), .Z(n18064) );
  XOR U18573 ( .A(b[47]), .B(a[47]), .Z(n18355) );
  NANDN U18574 ( .A(n37172), .B(n18355), .Z(n18063) );
  AND U18575 ( .A(n18064), .B(n18063), .Z(n18396) );
  NANDN U18576 ( .A(n210), .B(n18065), .Z(n18067) );
  XOR U18577 ( .A(a[85]), .B(b[9]), .Z(n18358) );
  NANDN U18578 ( .A(n30267), .B(n18358), .Z(n18066) );
  AND U18579 ( .A(n18067), .B(n18066), .Z(n18395) );
  NANDN U18580 ( .A(n212), .B(n18068), .Z(n18070) );
  XOR U18581 ( .A(b[49]), .B(a[45]), .Z(n18361) );
  NANDN U18582 ( .A(n37432), .B(n18361), .Z(n18069) );
  NAND U18583 ( .A(n18070), .B(n18069), .Z(n18394) );
  XOR U18584 ( .A(n18395), .B(n18394), .Z(n18397) );
  XOR U18585 ( .A(n18396), .B(n18397), .Z(n18461) );
  NANDN U18586 ( .A(n36742), .B(n18071), .Z(n18073) );
  XOR U18587 ( .A(b[43]), .B(a[51]), .Z(n18364) );
  NANDN U18588 ( .A(n36891), .B(n18364), .Z(n18072) );
  AND U18589 ( .A(n18073), .B(n18072), .Z(n18375) );
  NANDN U18590 ( .A(n36991), .B(n18074), .Z(n18076) );
  XOR U18591 ( .A(b[45]), .B(a[49]), .Z(n18367) );
  NANDN U18592 ( .A(n37083), .B(n18367), .Z(n18075) );
  AND U18593 ( .A(n18076), .B(n18075), .Z(n18374) );
  NANDN U18594 ( .A(n30482), .B(n18077), .Z(n18079) );
  XOR U18595 ( .A(a[83]), .B(b[11]), .Z(n18370) );
  NANDN U18596 ( .A(n30891), .B(n18370), .Z(n18078) );
  NAND U18597 ( .A(n18079), .B(n18078), .Z(n18373) );
  XOR U18598 ( .A(n18374), .B(n18373), .Z(n18376) );
  XNOR U18599 ( .A(n18375), .B(n18376), .Z(n18460) );
  XNOR U18600 ( .A(n18461), .B(n18460), .Z(n18462) );
  NANDN U18601 ( .A(n18081), .B(n18080), .Z(n18085) );
  OR U18602 ( .A(n18083), .B(n18082), .Z(n18084) );
  NAND U18603 ( .A(n18085), .B(n18084), .Z(n18463) );
  XNOR U18604 ( .A(n18462), .B(n18463), .Z(n18271) );
  XNOR U18605 ( .A(n18272), .B(n18271), .Z(n18273) );
  NANDN U18606 ( .A(n29499), .B(n18086), .Z(n18088) );
  XOR U18607 ( .A(a[87]), .B(b[7]), .Z(n18379) );
  NANDN U18608 ( .A(n29735), .B(n18379), .Z(n18087) );
  AND U18609 ( .A(n18088), .B(n18087), .Z(n18339) );
  NANDN U18610 ( .A(n37857), .B(n18089), .Z(n18091) );
  XOR U18611 ( .A(b[55]), .B(a[39]), .Z(n18382) );
  NANDN U18612 ( .A(n37911), .B(n18382), .Z(n18090) );
  AND U18613 ( .A(n18091), .B(n18090), .Z(n18338) );
  NANDN U18614 ( .A(n35611), .B(n18092), .Z(n18094) );
  XOR U18615 ( .A(b[35]), .B(a[59]), .Z(n18385) );
  NANDN U18616 ( .A(n35801), .B(n18385), .Z(n18093) );
  NAND U18617 ( .A(n18094), .B(n18093), .Z(n18337) );
  XOR U18618 ( .A(n18338), .B(n18337), .Z(n18340) );
  XOR U18619 ( .A(n18339), .B(n18340), .Z(n18401) );
  NANDN U18620 ( .A(n18096), .B(n18095), .Z(n18100) );
  OR U18621 ( .A(n18098), .B(n18097), .Z(n18099) );
  AND U18622 ( .A(n18100), .B(n18099), .Z(n18400) );
  XNOR U18623 ( .A(n18401), .B(n18400), .Z(n18402) );
  NANDN U18624 ( .A(n18102), .B(n18101), .Z(n18106) );
  OR U18625 ( .A(n18104), .B(n18103), .Z(n18105) );
  NAND U18626 ( .A(n18106), .B(n18105), .Z(n18403) );
  XOR U18627 ( .A(n18402), .B(n18403), .Z(n18274) );
  XNOR U18628 ( .A(n18273), .B(n18274), .Z(n18283) );
  XOR U18629 ( .A(n18284), .B(n18283), .Z(n18286) );
  XOR U18630 ( .A(n18285), .B(n18286), .Z(n18254) );
  NANDN U18631 ( .A(n18108), .B(n18107), .Z(n18112) );
  NANDN U18632 ( .A(n18110), .B(n18109), .Z(n18111) );
  AND U18633 ( .A(n18112), .B(n18111), .Z(n18267) );
  NANDN U18634 ( .A(n18114), .B(n18113), .Z(n18118) );
  NANDN U18635 ( .A(n18116), .B(n18115), .Z(n18117) );
  AND U18636 ( .A(n18118), .B(n18117), .Z(n18266) );
  NANDN U18637 ( .A(n18120), .B(n18119), .Z(n18124) );
  NAND U18638 ( .A(n18122), .B(n18121), .Z(n18123) );
  AND U18639 ( .A(n18124), .B(n18123), .Z(n18265) );
  XOR U18640 ( .A(n18266), .B(n18265), .Z(n18268) );
  XOR U18641 ( .A(n18267), .B(n18268), .Z(n18292) );
  NANDN U18642 ( .A(n18126), .B(n18125), .Z(n18130) );
  NANDN U18643 ( .A(n18128), .B(n18127), .Z(n18129) );
  AND U18644 ( .A(n18130), .B(n18129), .Z(n18413) );
  NANDN U18645 ( .A(n18132), .B(n18131), .Z(n18136) );
  OR U18646 ( .A(n18134), .B(n18133), .Z(n18135) );
  NAND U18647 ( .A(n18136), .B(n18135), .Z(n18412) );
  XNOR U18648 ( .A(n18413), .B(n18412), .Z(n18415) );
  NANDN U18649 ( .A(n18138), .B(n18137), .Z(n18142) );
  OR U18650 ( .A(n18140), .B(n18139), .Z(n18141) );
  AND U18651 ( .A(n18142), .B(n18141), .Z(n18310) );
  NAND U18652 ( .A(b[0]), .B(a[93]), .Z(n18143) );
  XNOR U18653 ( .A(b[1]), .B(n18143), .Z(n18145) );
  NANDN U18654 ( .A(b[0]), .B(a[92]), .Z(n18144) );
  NAND U18655 ( .A(n18145), .B(n18144), .Z(n18346) );
  NANDN U18656 ( .A(n38278), .B(n18146), .Z(n18148) );
  XOR U18657 ( .A(b[63]), .B(a[31]), .Z(n18439) );
  NANDN U18658 ( .A(n38279), .B(n18439), .Z(n18147) );
  AND U18659 ( .A(n18148), .B(n18147), .Z(n18344) );
  NANDN U18660 ( .A(n35260), .B(n18149), .Z(n18151) );
  XOR U18661 ( .A(b[33]), .B(a[61]), .Z(n18442) );
  NANDN U18662 ( .A(n35456), .B(n18442), .Z(n18150) );
  NAND U18663 ( .A(n18151), .B(n18150), .Z(n18343) );
  XNOR U18664 ( .A(n18344), .B(n18343), .Z(n18345) );
  XNOR U18665 ( .A(n18346), .B(n18345), .Z(n18307) );
  NANDN U18666 ( .A(n37974), .B(n18152), .Z(n18154) );
  XOR U18667 ( .A(b[57]), .B(a[37]), .Z(n18445) );
  NANDN U18668 ( .A(n38031), .B(n18445), .Z(n18153) );
  AND U18669 ( .A(n18154), .B(n18153), .Z(n18421) );
  NANDN U18670 ( .A(n38090), .B(n18155), .Z(n18157) );
  XOR U18671 ( .A(b[59]), .B(a[35]), .Z(n18448) );
  NANDN U18672 ( .A(n38130), .B(n18448), .Z(n18156) );
  AND U18673 ( .A(n18157), .B(n18156), .Z(n18419) );
  NANDN U18674 ( .A(n36480), .B(n18158), .Z(n18160) );
  XOR U18675 ( .A(b[41]), .B(a[53]), .Z(n18451) );
  NANDN U18676 ( .A(n36594), .B(n18451), .Z(n18159) );
  NAND U18677 ( .A(n18160), .B(n18159), .Z(n18418) );
  XNOR U18678 ( .A(n18419), .B(n18418), .Z(n18420) );
  XOR U18679 ( .A(n18421), .B(n18420), .Z(n18308) );
  XNOR U18680 ( .A(n18307), .B(n18308), .Z(n18309) );
  XNOR U18681 ( .A(n18310), .B(n18309), .Z(n18414) );
  XOR U18682 ( .A(n18415), .B(n18414), .Z(n18296) );
  NANDN U18683 ( .A(n18162), .B(n18161), .Z(n18166) );
  NAND U18684 ( .A(n18164), .B(n18163), .Z(n18165) );
  NAND U18685 ( .A(n18166), .B(n18165), .Z(n18295) );
  XNOR U18686 ( .A(n18296), .B(n18295), .Z(n18298) );
  NANDN U18687 ( .A(n18168), .B(n18167), .Z(n18172) );
  NANDN U18688 ( .A(n18170), .B(n18169), .Z(n18171) );
  AND U18689 ( .A(n18172), .B(n18171), .Z(n18514) );
  NANDN U18690 ( .A(n32996), .B(n18173), .Z(n18175) );
  XOR U18691 ( .A(b[21]), .B(a[73]), .Z(n18466) );
  NANDN U18692 ( .A(n33271), .B(n18466), .Z(n18174) );
  AND U18693 ( .A(n18175), .B(n18174), .Z(n18432) );
  NANDN U18694 ( .A(n33866), .B(n18176), .Z(n18178) );
  XOR U18695 ( .A(b[23]), .B(a[71]), .Z(n18469) );
  NANDN U18696 ( .A(n33644), .B(n18469), .Z(n18177) );
  AND U18697 ( .A(n18178), .B(n18177), .Z(n18431) );
  NANDN U18698 ( .A(n32483), .B(n18179), .Z(n18181) );
  XOR U18699 ( .A(b[19]), .B(a[75]), .Z(n18472) );
  NANDN U18700 ( .A(n32823), .B(n18472), .Z(n18180) );
  NAND U18701 ( .A(n18181), .B(n18180), .Z(n18430) );
  XOR U18702 ( .A(n18431), .B(n18430), .Z(n18433) );
  XOR U18703 ( .A(n18432), .B(n18433), .Z(n18350) );
  NANDN U18704 ( .A(n34909), .B(n18182), .Z(n18184) );
  XOR U18705 ( .A(b[31]), .B(a[63]), .Z(n18475) );
  NANDN U18706 ( .A(n35145), .B(n18475), .Z(n18183) );
  AND U18707 ( .A(n18184), .B(n18183), .Z(n18390) );
  NANDN U18708 ( .A(n38247), .B(n18185), .Z(n18187) );
  XOR U18709 ( .A(b[61]), .B(a[33]), .Z(n18478) );
  NANDN U18710 ( .A(n38248), .B(n18478), .Z(n18186) );
  AND U18711 ( .A(n18187), .B(n18186), .Z(n18389) );
  AND U18712 ( .A(b[63]), .B(a[29]), .Z(n18388) );
  XOR U18713 ( .A(n18389), .B(n18388), .Z(n18391) );
  XNOR U18714 ( .A(n18390), .B(n18391), .Z(n18349) );
  XNOR U18715 ( .A(n18350), .B(n18349), .Z(n18351) );
  NANDN U18716 ( .A(n18189), .B(n18188), .Z(n18193) );
  OR U18717 ( .A(n18191), .B(n18190), .Z(n18192) );
  NAND U18718 ( .A(n18193), .B(n18192), .Z(n18352) );
  XNOR U18719 ( .A(n18351), .B(n18352), .Z(n18511) );
  NANDN U18720 ( .A(n34223), .B(n18194), .Z(n18196) );
  XOR U18721 ( .A(b[27]), .B(a[67]), .Z(n18487) );
  NANDN U18722 ( .A(n34458), .B(n18487), .Z(n18195) );
  AND U18723 ( .A(n18196), .B(n18195), .Z(n18333) );
  NANDN U18724 ( .A(n34634), .B(n18197), .Z(n18199) );
  XOR U18725 ( .A(b[29]), .B(a[65]), .Z(n18490) );
  NANDN U18726 ( .A(n34722), .B(n18490), .Z(n18198) );
  AND U18727 ( .A(n18199), .B(n18198), .Z(n18332) );
  NANDN U18728 ( .A(n31055), .B(n18200), .Z(n18202) );
  XOR U18729 ( .A(a[81]), .B(b[13]), .Z(n18493) );
  NANDN U18730 ( .A(n31293), .B(n18493), .Z(n18201) );
  NAND U18731 ( .A(n18202), .B(n18201), .Z(n18331) );
  XOR U18732 ( .A(n18332), .B(n18331), .Z(n18334) );
  XOR U18733 ( .A(n18333), .B(n18334), .Z(n18407) );
  NANDN U18734 ( .A(n28889), .B(n18203), .Z(n18205) );
  XOR U18735 ( .A(a[89]), .B(b[5]), .Z(n18496) );
  NANDN U18736 ( .A(n29138), .B(n18496), .Z(n18204) );
  AND U18737 ( .A(n18205), .B(n18204), .Z(n18426) );
  NANDN U18738 ( .A(n209), .B(n18206), .Z(n18208) );
  XOR U18739 ( .A(a[91]), .B(b[3]), .Z(n18499) );
  NANDN U18740 ( .A(n28941), .B(n18499), .Z(n18207) );
  AND U18741 ( .A(n18208), .B(n18207), .Z(n18425) );
  NANDN U18742 ( .A(n35936), .B(n18209), .Z(n18211) );
  XOR U18743 ( .A(b[37]), .B(a[57]), .Z(n18502) );
  NANDN U18744 ( .A(n36047), .B(n18502), .Z(n18210) );
  NAND U18745 ( .A(n18211), .B(n18210), .Z(n18424) );
  XOR U18746 ( .A(n18425), .B(n18424), .Z(n18427) );
  XNOR U18747 ( .A(n18426), .B(n18427), .Z(n18406) );
  XNOR U18748 ( .A(n18407), .B(n18406), .Z(n18408) );
  NANDN U18749 ( .A(n18213), .B(n18212), .Z(n18217) );
  OR U18750 ( .A(n18215), .B(n18214), .Z(n18216) );
  NAND U18751 ( .A(n18217), .B(n18216), .Z(n18409) );
  XOR U18752 ( .A(n18408), .B(n18409), .Z(n18512) );
  XNOR U18753 ( .A(n18511), .B(n18512), .Z(n18513) );
  XNOR U18754 ( .A(n18514), .B(n18513), .Z(n18297) );
  XOR U18755 ( .A(n18298), .B(n18297), .Z(n18290) );
  NANDN U18756 ( .A(n18219), .B(n18218), .Z(n18223) );
  NANDN U18757 ( .A(n18221), .B(n18220), .Z(n18222) );
  AND U18758 ( .A(n18223), .B(n18222), .Z(n18289) );
  XNOR U18759 ( .A(n18290), .B(n18289), .Z(n18291) );
  XNOR U18760 ( .A(n18292), .B(n18291), .Z(n18253) );
  XNOR U18761 ( .A(n18254), .B(n18253), .Z(n18255) );
  XOR U18762 ( .A(n18256), .B(n18255), .Z(n18520) );
  XNOR U18763 ( .A(n18519), .B(n18520), .Z(n18525) );
  XOR U18764 ( .A(n18526), .B(n18525), .Z(n18248) );
  NANDN U18765 ( .A(n18225), .B(n18224), .Z(n18229) );
  NANDN U18766 ( .A(n18227), .B(n18226), .Z(n18228) );
  AND U18767 ( .A(n18229), .B(n18228), .Z(n18247) );
  XNOR U18768 ( .A(n18248), .B(n18247), .Z(n18249) );
  NANDN U18769 ( .A(n18231), .B(n18230), .Z(n18235) );
  NAND U18770 ( .A(n18233), .B(n18232), .Z(n18234) );
  NAND U18771 ( .A(n18235), .B(n18234), .Z(n18250) );
  XNOR U18772 ( .A(n18249), .B(n18250), .Z(n18241) );
  XNOR U18773 ( .A(n18242), .B(n18241), .Z(n18243) );
  XNOR U18774 ( .A(n18244), .B(n18243), .Z(n18529) );
  XNOR U18775 ( .A(sreg[157]), .B(n18529), .Z(n18531) );
  NANDN U18776 ( .A(sreg[156]), .B(n18236), .Z(n18240) );
  NAND U18777 ( .A(n18238), .B(n18237), .Z(n18239) );
  NAND U18778 ( .A(n18240), .B(n18239), .Z(n18530) );
  XNOR U18779 ( .A(n18531), .B(n18530), .Z(c[157]) );
  NANDN U18780 ( .A(n18242), .B(n18241), .Z(n18246) );
  NANDN U18781 ( .A(n18244), .B(n18243), .Z(n18245) );
  AND U18782 ( .A(n18246), .B(n18245), .Z(n18537) );
  NANDN U18783 ( .A(n18248), .B(n18247), .Z(n18252) );
  NANDN U18784 ( .A(n18250), .B(n18249), .Z(n18251) );
  AND U18785 ( .A(n18252), .B(n18251), .Z(n18535) );
  NANDN U18786 ( .A(n18254), .B(n18253), .Z(n18258) );
  NANDN U18787 ( .A(n18256), .B(n18255), .Z(n18257) );
  AND U18788 ( .A(n18258), .B(n18257), .Z(n18547) );
  NANDN U18789 ( .A(n18260), .B(n18259), .Z(n18264) );
  OR U18790 ( .A(n18262), .B(n18261), .Z(n18263) );
  AND U18791 ( .A(n18264), .B(n18263), .Z(n18546) );
  XNOR U18792 ( .A(n18547), .B(n18546), .Z(n18549) );
  NANDN U18793 ( .A(n18266), .B(n18265), .Z(n18270) );
  OR U18794 ( .A(n18268), .B(n18267), .Z(n18269) );
  AND U18795 ( .A(n18270), .B(n18269), .Z(n18818) );
  NANDN U18796 ( .A(n18272), .B(n18271), .Z(n18276) );
  NANDN U18797 ( .A(n18274), .B(n18273), .Z(n18275) );
  AND U18798 ( .A(n18276), .B(n18275), .Z(n18817) );
  NANDN U18799 ( .A(n18278), .B(n18277), .Z(n18282) );
  OR U18800 ( .A(n18280), .B(n18279), .Z(n18281) );
  AND U18801 ( .A(n18282), .B(n18281), .Z(n18816) );
  XOR U18802 ( .A(n18817), .B(n18816), .Z(n18819) );
  XOR U18803 ( .A(n18818), .B(n18819), .Z(n18553) );
  NANDN U18804 ( .A(n18284), .B(n18283), .Z(n18288) );
  OR U18805 ( .A(n18286), .B(n18285), .Z(n18287) );
  AND U18806 ( .A(n18288), .B(n18287), .Z(n18552) );
  XNOR U18807 ( .A(n18553), .B(n18552), .Z(n18554) );
  NANDN U18808 ( .A(n18290), .B(n18289), .Z(n18294) );
  NANDN U18809 ( .A(n18292), .B(n18291), .Z(n18293) );
  AND U18810 ( .A(n18294), .B(n18293), .Z(n18813) );
  NANDN U18811 ( .A(n18296), .B(n18295), .Z(n18300) );
  NAND U18812 ( .A(n18298), .B(n18297), .Z(n18299) );
  AND U18813 ( .A(n18300), .B(n18299), .Z(n18788) );
  NANDN U18814 ( .A(n18302), .B(n18301), .Z(n18306) );
  NANDN U18815 ( .A(n18304), .B(n18303), .Z(n18305) );
  AND U18816 ( .A(n18306), .B(n18305), .Z(n18806) );
  NANDN U18817 ( .A(n18308), .B(n18307), .Z(n18312) );
  NANDN U18818 ( .A(n18310), .B(n18309), .Z(n18311) );
  AND U18819 ( .A(n18312), .B(n18311), .Z(n18805) );
  NANDN U18820 ( .A(n33875), .B(n18313), .Z(n18315) );
  XOR U18821 ( .A(b[25]), .B(a[70]), .Z(n18582) );
  NANDN U18822 ( .A(n33994), .B(n18582), .Z(n18314) );
  AND U18823 ( .A(n18315), .B(n18314), .Z(n18776) );
  NANDN U18824 ( .A(n32013), .B(n18316), .Z(n18318) );
  XOR U18825 ( .A(b[17]), .B(a[78]), .Z(n18585) );
  NANDN U18826 ( .A(n32292), .B(n18585), .Z(n18317) );
  AND U18827 ( .A(n18318), .B(n18317), .Z(n18775) );
  NANDN U18828 ( .A(n31536), .B(n18319), .Z(n18321) );
  XOR U18829 ( .A(a[80]), .B(b[15]), .Z(n18588) );
  NANDN U18830 ( .A(n31925), .B(n18588), .Z(n18320) );
  NAND U18831 ( .A(n18321), .B(n18320), .Z(n18774) );
  XOR U18832 ( .A(n18775), .B(n18774), .Z(n18777) );
  XOR U18833 ( .A(n18776), .B(n18777), .Z(n18724) );
  NANDN U18834 ( .A(n37526), .B(n18322), .Z(n18324) );
  XOR U18835 ( .A(b[51]), .B(a[44]), .Z(n18591) );
  NANDN U18836 ( .A(n37605), .B(n18591), .Z(n18323) );
  AND U18837 ( .A(n18324), .B(n18323), .Z(n18755) );
  NANDN U18838 ( .A(n37705), .B(n18325), .Z(n18327) );
  XOR U18839 ( .A(b[53]), .B(a[42]), .Z(n18594) );
  NANDN U18840 ( .A(n37778), .B(n18594), .Z(n18326) );
  AND U18841 ( .A(n18327), .B(n18326), .Z(n18754) );
  NANDN U18842 ( .A(n36210), .B(n18328), .Z(n18330) );
  XOR U18843 ( .A(b[39]), .B(a[56]), .Z(n18597) );
  NANDN U18844 ( .A(n36347), .B(n18597), .Z(n18329) );
  NAND U18845 ( .A(n18330), .B(n18329), .Z(n18753) );
  XOR U18846 ( .A(n18754), .B(n18753), .Z(n18756) );
  XNOR U18847 ( .A(n18755), .B(n18756), .Z(n18723) );
  XNOR U18848 ( .A(n18724), .B(n18723), .Z(n18726) );
  NANDN U18849 ( .A(n18332), .B(n18331), .Z(n18336) );
  OR U18850 ( .A(n18334), .B(n18333), .Z(n18335) );
  AND U18851 ( .A(n18336), .B(n18335), .Z(n18725) );
  XOR U18852 ( .A(n18726), .B(n18725), .Z(n18573) );
  NANDN U18853 ( .A(n18338), .B(n18337), .Z(n18342) );
  OR U18854 ( .A(n18340), .B(n18339), .Z(n18341) );
  AND U18855 ( .A(n18342), .B(n18341), .Z(n18571) );
  NANDN U18856 ( .A(n18344), .B(n18343), .Z(n18348) );
  NANDN U18857 ( .A(n18346), .B(n18345), .Z(n18347) );
  NAND U18858 ( .A(n18348), .B(n18347), .Z(n18570) );
  XNOR U18859 ( .A(n18571), .B(n18570), .Z(n18572) );
  XNOR U18860 ( .A(n18573), .B(n18572), .Z(n18804) );
  XOR U18861 ( .A(n18805), .B(n18804), .Z(n18807) );
  XOR U18862 ( .A(n18806), .B(n18807), .Z(n18787) );
  NANDN U18863 ( .A(n18350), .B(n18349), .Z(n18354) );
  NANDN U18864 ( .A(n18352), .B(n18351), .Z(n18353) );
  AND U18865 ( .A(n18354), .B(n18353), .Z(n18799) );
  NANDN U18866 ( .A(n211), .B(n18355), .Z(n18357) );
  XOR U18867 ( .A(b[47]), .B(a[48]), .Z(n18645) );
  NANDN U18868 ( .A(n37172), .B(n18645), .Z(n18356) );
  AND U18869 ( .A(n18357), .B(n18356), .Z(n18635) );
  NANDN U18870 ( .A(n210), .B(n18358), .Z(n18360) );
  XOR U18871 ( .A(a[86]), .B(b[9]), .Z(n18648) );
  NANDN U18872 ( .A(n30267), .B(n18648), .Z(n18359) );
  AND U18873 ( .A(n18360), .B(n18359), .Z(n18634) );
  NANDN U18874 ( .A(n212), .B(n18361), .Z(n18363) );
  XOR U18875 ( .A(b[49]), .B(a[46]), .Z(n18651) );
  NANDN U18876 ( .A(n37432), .B(n18651), .Z(n18362) );
  NAND U18877 ( .A(n18363), .B(n18362), .Z(n18633) );
  XOR U18878 ( .A(n18634), .B(n18633), .Z(n18636) );
  XOR U18879 ( .A(n18635), .B(n18636), .Z(n18730) );
  NANDN U18880 ( .A(n36742), .B(n18364), .Z(n18366) );
  XOR U18881 ( .A(b[43]), .B(a[52]), .Z(n18654) );
  NANDN U18882 ( .A(n36891), .B(n18654), .Z(n18365) );
  AND U18883 ( .A(n18366), .B(n18365), .Z(n18665) );
  NANDN U18884 ( .A(n36991), .B(n18367), .Z(n18369) );
  XOR U18885 ( .A(b[45]), .B(a[50]), .Z(n18657) );
  NANDN U18886 ( .A(n37083), .B(n18657), .Z(n18368) );
  AND U18887 ( .A(n18369), .B(n18368), .Z(n18664) );
  NANDN U18888 ( .A(n30482), .B(n18370), .Z(n18372) );
  XOR U18889 ( .A(a[84]), .B(b[11]), .Z(n18660) );
  NANDN U18890 ( .A(n30891), .B(n18660), .Z(n18371) );
  NAND U18891 ( .A(n18372), .B(n18371), .Z(n18663) );
  XOR U18892 ( .A(n18664), .B(n18663), .Z(n18666) );
  XNOR U18893 ( .A(n18665), .B(n18666), .Z(n18729) );
  XNOR U18894 ( .A(n18730), .B(n18729), .Z(n18731) );
  NANDN U18895 ( .A(n18374), .B(n18373), .Z(n18378) );
  OR U18896 ( .A(n18376), .B(n18375), .Z(n18377) );
  NAND U18897 ( .A(n18378), .B(n18377), .Z(n18732) );
  XNOR U18898 ( .A(n18731), .B(n18732), .Z(n18798) );
  XNOR U18899 ( .A(n18799), .B(n18798), .Z(n18800) );
  NANDN U18900 ( .A(n29499), .B(n18379), .Z(n18381) );
  XOR U18901 ( .A(a[88]), .B(b[7]), .Z(n18618) );
  NANDN U18902 ( .A(n29735), .B(n18618), .Z(n18380) );
  AND U18903 ( .A(n18381), .B(n18380), .Z(n18608) );
  NANDN U18904 ( .A(n37857), .B(n18382), .Z(n18384) );
  XOR U18905 ( .A(b[55]), .B(a[40]), .Z(n18621) );
  NANDN U18906 ( .A(n37911), .B(n18621), .Z(n18383) );
  AND U18907 ( .A(n18384), .B(n18383), .Z(n18607) );
  NANDN U18908 ( .A(n35611), .B(n18385), .Z(n18387) );
  XOR U18909 ( .A(b[35]), .B(a[60]), .Z(n18624) );
  NANDN U18910 ( .A(n35801), .B(n18624), .Z(n18386) );
  NAND U18911 ( .A(n18387), .B(n18386), .Z(n18606) );
  XOR U18912 ( .A(n18607), .B(n18606), .Z(n18609) );
  XOR U18913 ( .A(n18608), .B(n18609), .Z(n18670) );
  NANDN U18914 ( .A(n18389), .B(n18388), .Z(n18393) );
  OR U18915 ( .A(n18391), .B(n18390), .Z(n18392) );
  AND U18916 ( .A(n18393), .B(n18392), .Z(n18669) );
  XNOR U18917 ( .A(n18670), .B(n18669), .Z(n18671) );
  NANDN U18918 ( .A(n18395), .B(n18394), .Z(n18399) );
  OR U18919 ( .A(n18397), .B(n18396), .Z(n18398) );
  NAND U18920 ( .A(n18399), .B(n18398), .Z(n18672) );
  XOR U18921 ( .A(n18671), .B(n18672), .Z(n18801) );
  XNOR U18922 ( .A(n18800), .B(n18801), .Z(n18786) );
  XOR U18923 ( .A(n18787), .B(n18786), .Z(n18789) );
  XOR U18924 ( .A(n18788), .B(n18789), .Z(n18811) );
  NANDN U18925 ( .A(n18401), .B(n18400), .Z(n18405) );
  NANDN U18926 ( .A(n18403), .B(n18402), .Z(n18404) );
  AND U18927 ( .A(n18405), .B(n18404), .Z(n18794) );
  NANDN U18928 ( .A(n18407), .B(n18406), .Z(n18411) );
  NANDN U18929 ( .A(n18409), .B(n18408), .Z(n18410) );
  AND U18930 ( .A(n18411), .B(n18410), .Z(n18793) );
  NANDN U18931 ( .A(n18413), .B(n18412), .Z(n18417) );
  NAND U18932 ( .A(n18415), .B(n18414), .Z(n18416) );
  AND U18933 ( .A(n18417), .B(n18416), .Z(n18792) );
  XOR U18934 ( .A(n18793), .B(n18792), .Z(n18795) );
  XOR U18935 ( .A(n18794), .B(n18795), .Z(n18561) );
  NANDN U18936 ( .A(n18419), .B(n18418), .Z(n18423) );
  NANDN U18937 ( .A(n18421), .B(n18420), .Z(n18422) );
  AND U18938 ( .A(n18423), .B(n18422), .Z(n18682) );
  NANDN U18939 ( .A(n18425), .B(n18424), .Z(n18429) );
  OR U18940 ( .A(n18427), .B(n18426), .Z(n18428) );
  NAND U18941 ( .A(n18429), .B(n18428), .Z(n18681) );
  XNOR U18942 ( .A(n18682), .B(n18681), .Z(n18684) );
  NANDN U18943 ( .A(n18431), .B(n18430), .Z(n18435) );
  OR U18944 ( .A(n18433), .B(n18432), .Z(n18434) );
  AND U18945 ( .A(n18435), .B(n18434), .Z(n18579) );
  NAND U18946 ( .A(b[0]), .B(a[94]), .Z(n18436) );
  XNOR U18947 ( .A(b[1]), .B(n18436), .Z(n18438) );
  NANDN U18948 ( .A(b[0]), .B(a[93]), .Z(n18437) );
  NAND U18949 ( .A(n18438), .B(n18437), .Z(n18615) );
  NANDN U18950 ( .A(n38278), .B(n18439), .Z(n18441) );
  XOR U18951 ( .A(b[63]), .B(a[32]), .Z(n18708) );
  NANDN U18952 ( .A(n38279), .B(n18708), .Z(n18440) );
  AND U18953 ( .A(n18441), .B(n18440), .Z(n18613) );
  NANDN U18954 ( .A(n35260), .B(n18442), .Z(n18444) );
  XOR U18955 ( .A(b[33]), .B(a[62]), .Z(n18711) );
  NANDN U18956 ( .A(n35456), .B(n18711), .Z(n18443) );
  NAND U18957 ( .A(n18444), .B(n18443), .Z(n18612) );
  XNOR U18958 ( .A(n18613), .B(n18612), .Z(n18614) );
  XNOR U18959 ( .A(n18615), .B(n18614), .Z(n18576) );
  NANDN U18960 ( .A(n37974), .B(n18445), .Z(n18447) );
  XOR U18961 ( .A(b[57]), .B(a[38]), .Z(n18714) );
  NANDN U18962 ( .A(n38031), .B(n18714), .Z(n18446) );
  AND U18963 ( .A(n18447), .B(n18446), .Z(n18690) );
  NANDN U18964 ( .A(n38090), .B(n18448), .Z(n18450) );
  XOR U18965 ( .A(b[59]), .B(a[36]), .Z(n18717) );
  NANDN U18966 ( .A(n38130), .B(n18717), .Z(n18449) );
  AND U18967 ( .A(n18450), .B(n18449), .Z(n18688) );
  NANDN U18968 ( .A(n36480), .B(n18451), .Z(n18453) );
  XOR U18969 ( .A(b[41]), .B(a[54]), .Z(n18720) );
  NANDN U18970 ( .A(n36594), .B(n18720), .Z(n18452) );
  NAND U18971 ( .A(n18453), .B(n18452), .Z(n18687) );
  XNOR U18972 ( .A(n18688), .B(n18687), .Z(n18689) );
  XOR U18973 ( .A(n18690), .B(n18689), .Z(n18577) );
  XNOR U18974 ( .A(n18576), .B(n18577), .Z(n18578) );
  XNOR U18975 ( .A(n18579), .B(n18578), .Z(n18683) );
  XOR U18976 ( .A(n18684), .B(n18683), .Z(n18565) );
  NANDN U18977 ( .A(n18455), .B(n18454), .Z(n18459) );
  NAND U18978 ( .A(n18457), .B(n18456), .Z(n18458) );
  NAND U18979 ( .A(n18459), .B(n18458), .Z(n18564) );
  XNOR U18980 ( .A(n18565), .B(n18564), .Z(n18567) );
  NANDN U18981 ( .A(n18461), .B(n18460), .Z(n18465) );
  NANDN U18982 ( .A(n18463), .B(n18462), .Z(n18464) );
  AND U18983 ( .A(n18465), .B(n18464), .Z(n18783) );
  NANDN U18984 ( .A(n32996), .B(n18466), .Z(n18468) );
  XOR U18985 ( .A(b[21]), .B(a[74]), .Z(n18759) );
  NANDN U18986 ( .A(n33271), .B(n18759), .Z(n18467) );
  AND U18987 ( .A(n18468), .B(n18467), .Z(n18701) );
  NANDN U18988 ( .A(n33866), .B(n18469), .Z(n18471) );
  XOR U18989 ( .A(b[23]), .B(a[72]), .Z(n18762) );
  NANDN U18990 ( .A(n33644), .B(n18762), .Z(n18470) );
  AND U18991 ( .A(n18471), .B(n18470), .Z(n18700) );
  NANDN U18992 ( .A(n32483), .B(n18472), .Z(n18474) );
  XOR U18993 ( .A(b[19]), .B(a[76]), .Z(n18765) );
  NANDN U18994 ( .A(n32823), .B(n18765), .Z(n18473) );
  NAND U18995 ( .A(n18474), .B(n18473), .Z(n18699) );
  XOR U18996 ( .A(n18700), .B(n18699), .Z(n18702) );
  XOR U18997 ( .A(n18701), .B(n18702), .Z(n18640) );
  NANDN U18998 ( .A(n34909), .B(n18475), .Z(n18477) );
  XOR U18999 ( .A(b[31]), .B(a[64]), .Z(n18768) );
  NANDN U19000 ( .A(n35145), .B(n18768), .Z(n18476) );
  AND U19001 ( .A(n18477), .B(n18476), .Z(n18629) );
  NANDN U19002 ( .A(n38247), .B(n18478), .Z(n18480) );
  XOR U19003 ( .A(b[61]), .B(a[34]), .Z(n18771) );
  NANDN U19004 ( .A(n38248), .B(n18771), .Z(n18479) );
  AND U19005 ( .A(n18480), .B(n18479), .Z(n18628) );
  AND U19006 ( .A(b[63]), .B(a[30]), .Z(n18627) );
  XOR U19007 ( .A(n18628), .B(n18627), .Z(n18630) );
  XNOR U19008 ( .A(n18629), .B(n18630), .Z(n18639) );
  XNOR U19009 ( .A(n18640), .B(n18639), .Z(n18641) );
  NANDN U19010 ( .A(n18482), .B(n18481), .Z(n18486) );
  OR U19011 ( .A(n18484), .B(n18483), .Z(n18485) );
  NAND U19012 ( .A(n18486), .B(n18485), .Z(n18642) );
  XNOR U19013 ( .A(n18641), .B(n18642), .Z(n18780) );
  NANDN U19014 ( .A(n34223), .B(n18487), .Z(n18489) );
  XOR U19015 ( .A(b[27]), .B(a[68]), .Z(n18735) );
  NANDN U19016 ( .A(n34458), .B(n18735), .Z(n18488) );
  AND U19017 ( .A(n18489), .B(n18488), .Z(n18602) );
  NANDN U19018 ( .A(n34634), .B(n18490), .Z(n18492) );
  XOR U19019 ( .A(b[29]), .B(a[66]), .Z(n18738) );
  NANDN U19020 ( .A(n34722), .B(n18738), .Z(n18491) );
  AND U19021 ( .A(n18492), .B(n18491), .Z(n18601) );
  NANDN U19022 ( .A(n31055), .B(n18493), .Z(n18495) );
  XOR U19023 ( .A(a[82]), .B(b[13]), .Z(n18741) );
  NANDN U19024 ( .A(n31293), .B(n18741), .Z(n18494) );
  NAND U19025 ( .A(n18495), .B(n18494), .Z(n18600) );
  XOR U19026 ( .A(n18601), .B(n18600), .Z(n18603) );
  XOR U19027 ( .A(n18602), .B(n18603), .Z(n18676) );
  NANDN U19028 ( .A(n28889), .B(n18496), .Z(n18498) );
  XOR U19029 ( .A(a[90]), .B(b[5]), .Z(n18744) );
  NANDN U19030 ( .A(n29138), .B(n18744), .Z(n18497) );
  AND U19031 ( .A(n18498), .B(n18497), .Z(n18695) );
  NANDN U19032 ( .A(n209), .B(n18499), .Z(n18501) );
  XOR U19033 ( .A(a[92]), .B(b[3]), .Z(n18747) );
  NANDN U19034 ( .A(n28941), .B(n18747), .Z(n18500) );
  AND U19035 ( .A(n18501), .B(n18500), .Z(n18694) );
  NANDN U19036 ( .A(n35936), .B(n18502), .Z(n18504) );
  XOR U19037 ( .A(b[37]), .B(a[58]), .Z(n18750) );
  NANDN U19038 ( .A(n36047), .B(n18750), .Z(n18503) );
  NAND U19039 ( .A(n18504), .B(n18503), .Z(n18693) );
  XOR U19040 ( .A(n18694), .B(n18693), .Z(n18696) );
  XNOR U19041 ( .A(n18695), .B(n18696), .Z(n18675) );
  XNOR U19042 ( .A(n18676), .B(n18675), .Z(n18677) );
  NANDN U19043 ( .A(n18506), .B(n18505), .Z(n18510) );
  OR U19044 ( .A(n18508), .B(n18507), .Z(n18509) );
  NAND U19045 ( .A(n18510), .B(n18509), .Z(n18678) );
  XOR U19046 ( .A(n18677), .B(n18678), .Z(n18781) );
  XNOR U19047 ( .A(n18780), .B(n18781), .Z(n18782) );
  XNOR U19048 ( .A(n18783), .B(n18782), .Z(n18566) );
  XOR U19049 ( .A(n18567), .B(n18566), .Z(n18559) );
  NANDN U19050 ( .A(n18512), .B(n18511), .Z(n18516) );
  NANDN U19051 ( .A(n18514), .B(n18513), .Z(n18515) );
  AND U19052 ( .A(n18516), .B(n18515), .Z(n18558) );
  XNOR U19053 ( .A(n18559), .B(n18558), .Z(n18560) );
  XNOR U19054 ( .A(n18561), .B(n18560), .Z(n18810) );
  XNOR U19055 ( .A(n18811), .B(n18810), .Z(n18812) );
  XOR U19056 ( .A(n18813), .B(n18812), .Z(n18555) );
  XNOR U19057 ( .A(n18554), .B(n18555), .Z(n18548) );
  XOR U19058 ( .A(n18549), .B(n18548), .Z(n18541) );
  NANDN U19059 ( .A(n18518), .B(n18517), .Z(n18522) );
  NANDN U19060 ( .A(n18520), .B(n18519), .Z(n18521) );
  AND U19061 ( .A(n18522), .B(n18521), .Z(n18540) );
  XNOR U19062 ( .A(n18541), .B(n18540), .Z(n18542) );
  NANDN U19063 ( .A(n18524), .B(n18523), .Z(n18528) );
  NAND U19064 ( .A(n18526), .B(n18525), .Z(n18527) );
  NAND U19065 ( .A(n18528), .B(n18527), .Z(n18543) );
  XNOR U19066 ( .A(n18542), .B(n18543), .Z(n18534) );
  XNOR U19067 ( .A(n18535), .B(n18534), .Z(n18536) );
  XNOR U19068 ( .A(n18537), .B(n18536), .Z(n18822) );
  XNOR U19069 ( .A(sreg[158]), .B(n18822), .Z(n18824) );
  NANDN U19070 ( .A(sreg[157]), .B(n18529), .Z(n18533) );
  NAND U19071 ( .A(n18531), .B(n18530), .Z(n18532) );
  NAND U19072 ( .A(n18533), .B(n18532), .Z(n18823) );
  XNOR U19073 ( .A(n18824), .B(n18823), .Z(c[158]) );
  NANDN U19074 ( .A(n18535), .B(n18534), .Z(n18539) );
  NANDN U19075 ( .A(n18537), .B(n18536), .Z(n18538) );
  AND U19076 ( .A(n18539), .B(n18538), .Z(n18830) );
  NANDN U19077 ( .A(n18541), .B(n18540), .Z(n18545) );
  NANDN U19078 ( .A(n18543), .B(n18542), .Z(n18544) );
  AND U19079 ( .A(n18545), .B(n18544), .Z(n18828) );
  NANDN U19080 ( .A(n18547), .B(n18546), .Z(n18551) );
  NAND U19081 ( .A(n18549), .B(n18548), .Z(n18550) );
  AND U19082 ( .A(n18551), .B(n18550), .Z(n18835) );
  NANDN U19083 ( .A(n18553), .B(n18552), .Z(n18557) );
  NANDN U19084 ( .A(n18555), .B(n18554), .Z(n18556) );
  AND U19085 ( .A(n18557), .B(n18556), .Z(n18834) );
  NANDN U19086 ( .A(n18559), .B(n18558), .Z(n18563) );
  NANDN U19087 ( .A(n18561), .B(n18560), .Z(n18562) );
  AND U19088 ( .A(n18563), .B(n18562), .Z(n19093) );
  NANDN U19089 ( .A(n18565), .B(n18564), .Z(n18569) );
  NAND U19090 ( .A(n18567), .B(n18566), .Z(n18568) );
  AND U19091 ( .A(n18569), .B(n18568), .Z(n19069) );
  NANDN U19092 ( .A(n18571), .B(n18570), .Z(n18575) );
  NANDN U19093 ( .A(n18573), .B(n18572), .Z(n18574) );
  AND U19094 ( .A(n18575), .B(n18574), .Z(n19087) );
  NANDN U19095 ( .A(n18577), .B(n18576), .Z(n18581) );
  NANDN U19096 ( .A(n18579), .B(n18578), .Z(n18580) );
  AND U19097 ( .A(n18581), .B(n18580), .Z(n19086) );
  NANDN U19098 ( .A(n33875), .B(n18582), .Z(n18584) );
  XOR U19099 ( .A(b[25]), .B(a[71]), .Z(n18863) );
  NANDN U19100 ( .A(n33994), .B(n18863), .Z(n18583) );
  AND U19101 ( .A(n18584), .B(n18583), .Z(n19033) );
  NANDN U19102 ( .A(n32013), .B(n18585), .Z(n18587) );
  XOR U19103 ( .A(b[17]), .B(a[79]), .Z(n18866) );
  NANDN U19104 ( .A(n32292), .B(n18866), .Z(n18586) );
  AND U19105 ( .A(n18587), .B(n18586), .Z(n19032) );
  NANDN U19106 ( .A(n31536), .B(n18588), .Z(n18590) );
  XOR U19107 ( .A(a[81]), .B(b[15]), .Z(n18869) );
  NANDN U19108 ( .A(n31925), .B(n18869), .Z(n18589) );
  NAND U19109 ( .A(n18590), .B(n18589), .Z(n19031) );
  XOR U19110 ( .A(n19032), .B(n19031), .Z(n19034) );
  XOR U19111 ( .A(n19033), .B(n19034), .Z(n19005) );
  NANDN U19112 ( .A(n37526), .B(n18591), .Z(n18593) );
  XOR U19113 ( .A(b[51]), .B(a[45]), .Z(n18872) );
  NANDN U19114 ( .A(n37605), .B(n18872), .Z(n18592) );
  AND U19115 ( .A(n18593), .B(n18592), .Z(n19057) );
  NANDN U19116 ( .A(n37705), .B(n18594), .Z(n18596) );
  XOR U19117 ( .A(b[53]), .B(a[43]), .Z(n18875) );
  NANDN U19118 ( .A(n37778), .B(n18875), .Z(n18595) );
  AND U19119 ( .A(n18596), .B(n18595), .Z(n19056) );
  NANDN U19120 ( .A(n36210), .B(n18597), .Z(n18599) );
  XOR U19121 ( .A(b[39]), .B(a[57]), .Z(n18878) );
  NANDN U19122 ( .A(n36347), .B(n18878), .Z(n18598) );
  NAND U19123 ( .A(n18599), .B(n18598), .Z(n19055) );
  XOR U19124 ( .A(n19056), .B(n19055), .Z(n19058) );
  XNOR U19125 ( .A(n19057), .B(n19058), .Z(n19004) );
  XNOR U19126 ( .A(n19005), .B(n19004), .Z(n19007) );
  NANDN U19127 ( .A(n18601), .B(n18600), .Z(n18605) );
  OR U19128 ( .A(n18603), .B(n18602), .Z(n18604) );
  AND U19129 ( .A(n18605), .B(n18604), .Z(n19006) );
  XOR U19130 ( .A(n19007), .B(n19006), .Z(n18854) );
  NANDN U19131 ( .A(n18607), .B(n18606), .Z(n18611) );
  OR U19132 ( .A(n18609), .B(n18608), .Z(n18610) );
  AND U19133 ( .A(n18611), .B(n18610), .Z(n18852) );
  NANDN U19134 ( .A(n18613), .B(n18612), .Z(n18617) );
  NANDN U19135 ( .A(n18615), .B(n18614), .Z(n18616) );
  NAND U19136 ( .A(n18617), .B(n18616), .Z(n18851) );
  XNOR U19137 ( .A(n18852), .B(n18851), .Z(n18853) );
  XNOR U19138 ( .A(n18854), .B(n18853), .Z(n19085) );
  XOR U19139 ( .A(n19086), .B(n19085), .Z(n19088) );
  XOR U19140 ( .A(n19087), .B(n19088), .Z(n19068) );
  NANDN U19141 ( .A(n29499), .B(n18618), .Z(n18620) );
  XOR U19142 ( .A(a[89]), .B(b[7]), .Z(n18929) );
  NANDN U19143 ( .A(n29735), .B(n18929), .Z(n18619) );
  AND U19144 ( .A(n18620), .B(n18619), .Z(n18889) );
  NANDN U19145 ( .A(n37857), .B(n18621), .Z(n18623) );
  XOR U19146 ( .A(b[55]), .B(a[41]), .Z(n18932) );
  NANDN U19147 ( .A(n37911), .B(n18932), .Z(n18622) );
  AND U19148 ( .A(n18623), .B(n18622), .Z(n18888) );
  NANDN U19149 ( .A(n35611), .B(n18624), .Z(n18626) );
  XOR U19150 ( .A(b[35]), .B(a[61]), .Z(n18935) );
  NANDN U19151 ( .A(n35801), .B(n18935), .Z(n18625) );
  NAND U19152 ( .A(n18626), .B(n18625), .Z(n18887) );
  XOR U19153 ( .A(n18888), .B(n18887), .Z(n18890) );
  XOR U19154 ( .A(n18889), .B(n18890), .Z(n18951) );
  NANDN U19155 ( .A(n18628), .B(n18627), .Z(n18632) );
  OR U19156 ( .A(n18630), .B(n18629), .Z(n18631) );
  AND U19157 ( .A(n18632), .B(n18631), .Z(n18950) );
  XNOR U19158 ( .A(n18951), .B(n18950), .Z(n18952) );
  NANDN U19159 ( .A(n18634), .B(n18633), .Z(n18638) );
  OR U19160 ( .A(n18636), .B(n18635), .Z(n18637) );
  NAND U19161 ( .A(n18638), .B(n18637), .Z(n18953) );
  XNOR U19162 ( .A(n18952), .B(n18953), .Z(n19081) );
  NANDN U19163 ( .A(n18640), .B(n18639), .Z(n18644) );
  NANDN U19164 ( .A(n18642), .B(n18641), .Z(n18643) );
  AND U19165 ( .A(n18644), .B(n18643), .Z(n19080) );
  NANDN U19166 ( .A(n211), .B(n18645), .Z(n18647) );
  XOR U19167 ( .A(b[47]), .B(a[49]), .Z(n18905) );
  NANDN U19168 ( .A(n37172), .B(n18905), .Z(n18646) );
  AND U19169 ( .A(n18647), .B(n18646), .Z(n18946) );
  NANDN U19170 ( .A(n210), .B(n18648), .Z(n18650) );
  XOR U19171 ( .A(a[87]), .B(b[9]), .Z(n18908) );
  NANDN U19172 ( .A(n30267), .B(n18908), .Z(n18649) );
  AND U19173 ( .A(n18650), .B(n18649), .Z(n18945) );
  NANDN U19174 ( .A(n212), .B(n18651), .Z(n18653) );
  XOR U19175 ( .A(b[49]), .B(a[47]), .Z(n18911) );
  NANDN U19176 ( .A(n37432), .B(n18911), .Z(n18652) );
  NAND U19177 ( .A(n18653), .B(n18652), .Z(n18944) );
  XOR U19178 ( .A(n18945), .B(n18944), .Z(n18947) );
  XOR U19179 ( .A(n18946), .B(n18947), .Z(n19011) );
  NANDN U19180 ( .A(n36742), .B(n18654), .Z(n18656) );
  XOR U19181 ( .A(b[43]), .B(a[53]), .Z(n18914) );
  NANDN U19182 ( .A(n36891), .B(n18914), .Z(n18655) );
  AND U19183 ( .A(n18656), .B(n18655), .Z(n18925) );
  NANDN U19184 ( .A(n36991), .B(n18657), .Z(n18659) );
  XOR U19185 ( .A(b[45]), .B(a[51]), .Z(n18917) );
  NANDN U19186 ( .A(n37083), .B(n18917), .Z(n18658) );
  AND U19187 ( .A(n18659), .B(n18658), .Z(n18924) );
  NANDN U19188 ( .A(n30482), .B(n18660), .Z(n18662) );
  XOR U19189 ( .A(a[85]), .B(b[11]), .Z(n18920) );
  NANDN U19190 ( .A(n30891), .B(n18920), .Z(n18661) );
  NAND U19191 ( .A(n18662), .B(n18661), .Z(n18923) );
  XOR U19192 ( .A(n18924), .B(n18923), .Z(n18926) );
  XNOR U19193 ( .A(n18925), .B(n18926), .Z(n19010) );
  XNOR U19194 ( .A(n19011), .B(n19010), .Z(n19012) );
  NANDN U19195 ( .A(n18664), .B(n18663), .Z(n18668) );
  OR U19196 ( .A(n18666), .B(n18665), .Z(n18667) );
  NAND U19197 ( .A(n18668), .B(n18667), .Z(n19013) );
  XNOR U19198 ( .A(n19012), .B(n19013), .Z(n19079) );
  XOR U19199 ( .A(n19080), .B(n19079), .Z(n19082) );
  XNOR U19200 ( .A(n19081), .B(n19082), .Z(n19067) );
  XOR U19201 ( .A(n19068), .B(n19067), .Z(n19070) );
  XOR U19202 ( .A(n19069), .B(n19070), .Z(n19092) );
  NANDN U19203 ( .A(n18670), .B(n18669), .Z(n18674) );
  NANDN U19204 ( .A(n18672), .B(n18671), .Z(n18673) );
  AND U19205 ( .A(n18674), .B(n18673), .Z(n19075) );
  NANDN U19206 ( .A(n18676), .B(n18675), .Z(n18680) );
  NANDN U19207 ( .A(n18678), .B(n18677), .Z(n18679) );
  AND U19208 ( .A(n18680), .B(n18679), .Z(n19074) );
  NANDN U19209 ( .A(n18682), .B(n18681), .Z(n18686) );
  NAND U19210 ( .A(n18684), .B(n18683), .Z(n18685) );
  AND U19211 ( .A(n18686), .B(n18685), .Z(n19073) );
  XOR U19212 ( .A(n19074), .B(n19073), .Z(n19076) );
  XOR U19213 ( .A(n19075), .B(n19076), .Z(n18842) );
  NANDN U19214 ( .A(n18688), .B(n18687), .Z(n18692) );
  NANDN U19215 ( .A(n18690), .B(n18689), .Z(n18691) );
  AND U19216 ( .A(n18692), .B(n18691), .Z(n18963) );
  NANDN U19217 ( .A(n18694), .B(n18693), .Z(n18698) );
  OR U19218 ( .A(n18696), .B(n18695), .Z(n18697) );
  NAND U19219 ( .A(n18698), .B(n18697), .Z(n18962) );
  XNOR U19220 ( .A(n18963), .B(n18962), .Z(n18965) );
  NANDN U19221 ( .A(n18700), .B(n18699), .Z(n18704) );
  OR U19222 ( .A(n18702), .B(n18701), .Z(n18703) );
  AND U19223 ( .A(n18704), .B(n18703), .Z(n18860) );
  NAND U19224 ( .A(b[0]), .B(a[95]), .Z(n18705) );
  XNOR U19225 ( .A(b[1]), .B(n18705), .Z(n18707) );
  NANDN U19226 ( .A(b[0]), .B(a[94]), .Z(n18706) );
  NAND U19227 ( .A(n18707), .B(n18706), .Z(n18896) );
  NANDN U19228 ( .A(n38278), .B(n18708), .Z(n18710) );
  XOR U19229 ( .A(b[63]), .B(a[33]), .Z(n18989) );
  NANDN U19230 ( .A(n38279), .B(n18989), .Z(n18709) );
  AND U19231 ( .A(n18710), .B(n18709), .Z(n18894) );
  NANDN U19232 ( .A(n35260), .B(n18711), .Z(n18713) );
  XOR U19233 ( .A(b[33]), .B(a[63]), .Z(n18992) );
  NANDN U19234 ( .A(n35456), .B(n18992), .Z(n18712) );
  NAND U19235 ( .A(n18713), .B(n18712), .Z(n18893) );
  XNOR U19236 ( .A(n18894), .B(n18893), .Z(n18895) );
  XNOR U19237 ( .A(n18896), .B(n18895), .Z(n18857) );
  NANDN U19238 ( .A(n37974), .B(n18714), .Z(n18716) );
  XOR U19239 ( .A(b[57]), .B(a[39]), .Z(n18995) );
  NANDN U19240 ( .A(n38031), .B(n18995), .Z(n18715) );
  AND U19241 ( .A(n18716), .B(n18715), .Z(n18971) );
  NANDN U19242 ( .A(n38090), .B(n18717), .Z(n18719) );
  XOR U19243 ( .A(b[59]), .B(a[37]), .Z(n18998) );
  NANDN U19244 ( .A(n38130), .B(n18998), .Z(n18718) );
  AND U19245 ( .A(n18719), .B(n18718), .Z(n18969) );
  NANDN U19246 ( .A(n36480), .B(n18720), .Z(n18722) );
  XOR U19247 ( .A(b[41]), .B(a[55]), .Z(n19001) );
  NANDN U19248 ( .A(n36594), .B(n19001), .Z(n18721) );
  NAND U19249 ( .A(n18722), .B(n18721), .Z(n18968) );
  XNOR U19250 ( .A(n18969), .B(n18968), .Z(n18970) );
  XOR U19251 ( .A(n18971), .B(n18970), .Z(n18858) );
  XNOR U19252 ( .A(n18857), .B(n18858), .Z(n18859) );
  XNOR U19253 ( .A(n18860), .B(n18859), .Z(n18964) );
  XOR U19254 ( .A(n18965), .B(n18964), .Z(n18846) );
  NANDN U19255 ( .A(n18724), .B(n18723), .Z(n18728) );
  NAND U19256 ( .A(n18726), .B(n18725), .Z(n18727) );
  NAND U19257 ( .A(n18728), .B(n18727), .Z(n18845) );
  XNOR U19258 ( .A(n18846), .B(n18845), .Z(n18848) );
  NANDN U19259 ( .A(n18730), .B(n18729), .Z(n18734) );
  NANDN U19260 ( .A(n18732), .B(n18731), .Z(n18733) );
  AND U19261 ( .A(n18734), .B(n18733), .Z(n19064) );
  NANDN U19262 ( .A(n34223), .B(n18735), .Z(n18737) );
  XOR U19263 ( .A(b[27]), .B(a[69]), .Z(n19037) );
  NANDN U19264 ( .A(n34458), .B(n19037), .Z(n18736) );
  AND U19265 ( .A(n18737), .B(n18736), .Z(n18883) );
  NANDN U19266 ( .A(n34634), .B(n18738), .Z(n18740) );
  XOR U19267 ( .A(b[29]), .B(a[67]), .Z(n19040) );
  NANDN U19268 ( .A(n34722), .B(n19040), .Z(n18739) );
  AND U19269 ( .A(n18740), .B(n18739), .Z(n18882) );
  NANDN U19270 ( .A(n31055), .B(n18741), .Z(n18743) );
  XOR U19271 ( .A(a[83]), .B(b[13]), .Z(n19043) );
  NANDN U19272 ( .A(n31293), .B(n19043), .Z(n18742) );
  NAND U19273 ( .A(n18743), .B(n18742), .Z(n18881) );
  XOR U19274 ( .A(n18882), .B(n18881), .Z(n18884) );
  XOR U19275 ( .A(n18883), .B(n18884), .Z(n18957) );
  NANDN U19276 ( .A(n28889), .B(n18744), .Z(n18746) );
  XOR U19277 ( .A(a[91]), .B(b[5]), .Z(n19046) );
  NANDN U19278 ( .A(n29138), .B(n19046), .Z(n18745) );
  AND U19279 ( .A(n18746), .B(n18745), .Z(n18976) );
  NANDN U19280 ( .A(n209), .B(n18747), .Z(n18749) );
  XOR U19281 ( .A(a[93]), .B(b[3]), .Z(n19049) );
  NANDN U19282 ( .A(n28941), .B(n19049), .Z(n18748) );
  AND U19283 ( .A(n18749), .B(n18748), .Z(n18975) );
  NANDN U19284 ( .A(n35936), .B(n18750), .Z(n18752) );
  XOR U19285 ( .A(b[37]), .B(a[59]), .Z(n19052) );
  NANDN U19286 ( .A(n36047), .B(n19052), .Z(n18751) );
  NAND U19287 ( .A(n18752), .B(n18751), .Z(n18974) );
  XOR U19288 ( .A(n18975), .B(n18974), .Z(n18977) );
  XNOR U19289 ( .A(n18976), .B(n18977), .Z(n18956) );
  XNOR U19290 ( .A(n18957), .B(n18956), .Z(n18958) );
  NANDN U19291 ( .A(n18754), .B(n18753), .Z(n18758) );
  OR U19292 ( .A(n18756), .B(n18755), .Z(n18757) );
  NAND U19293 ( .A(n18758), .B(n18757), .Z(n18959) );
  XNOR U19294 ( .A(n18958), .B(n18959), .Z(n19061) );
  NANDN U19295 ( .A(n32996), .B(n18759), .Z(n18761) );
  XOR U19296 ( .A(b[21]), .B(a[75]), .Z(n19016) );
  NANDN U19297 ( .A(n33271), .B(n19016), .Z(n18760) );
  AND U19298 ( .A(n18761), .B(n18760), .Z(n18982) );
  NANDN U19299 ( .A(n33866), .B(n18762), .Z(n18764) );
  XOR U19300 ( .A(b[23]), .B(a[73]), .Z(n19019) );
  NANDN U19301 ( .A(n33644), .B(n19019), .Z(n18763) );
  AND U19302 ( .A(n18764), .B(n18763), .Z(n18981) );
  NANDN U19303 ( .A(n32483), .B(n18765), .Z(n18767) );
  XOR U19304 ( .A(b[19]), .B(a[77]), .Z(n19022) );
  NANDN U19305 ( .A(n32823), .B(n19022), .Z(n18766) );
  NAND U19306 ( .A(n18767), .B(n18766), .Z(n18980) );
  XOR U19307 ( .A(n18981), .B(n18980), .Z(n18983) );
  XOR U19308 ( .A(n18982), .B(n18983), .Z(n18900) );
  NANDN U19309 ( .A(n34909), .B(n18768), .Z(n18770) );
  XOR U19310 ( .A(b[31]), .B(a[65]), .Z(n19025) );
  NANDN U19311 ( .A(n35145), .B(n19025), .Z(n18769) );
  AND U19312 ( .A(n18770), .B(n18769), .Z(n18940) );
  NANDN U19313 ( .A(n38247), .B(n18771), .Z(n18773) );
  XOR U19314 ( .A(b[61]), .B(a[35]), .Z(n19028) );
  NANDN U19315 ( .A(n38248), .B(n19028), .Z(n18772) );
  AND U19316 ( .A(n18773), .B(n18772), .Z(n18939) );
  AND U19317 ( .A(b[63]), .B(a[31]), .Z(n18938) );
  XOR U19318 ( .A(n18939), .B(n18938), .Z(n18941) );
  XNOR U19319 ( .A(n18940), .B(n18941), .Z(n18899) );
  XNOR U19320 ( .A(n18900), .B(n18899), .Z(n18901) );
  NANDN U19321 ( .A(n18775), .B(n18774), .Z(n18779) );
  OR U19322 ( .A(n18777), .B(n18776), .Z(n18778) );
  NAND U19323 ( .A(n18779), .B(n18778), .Z(n18902) );
  XOR U19324 ( .A(n18901), .B(n18902), .Z(n19062) );
  XNOR U19325 ( .A(n19061), .B(n19062), .Z(n19063) );
  XNOR U19326 ( .A(n19064), .B(n19063), .Z(n18847) );
  XOR U19327 ( .A(n18848), .B(n18847), .Z(n18840) );
  NANDN U19328 ( .A(n18781), .B(n18780), .Z(n18785) );
  NANDN U19329 ( .A(n18783), .B(n18782), .Z(n18784) );
  AND U19330 ( .A(n18785), .B(n18784), .Z(n18839) );
  XNOR U19331 ( .A(n18840), .B(n18839), .Z(n18841) );
  XNOR U19332 ( .A(n18842), .B(n18841), .Z(n19091) );
  XOR U19333 ( .A(n19092), .B(n19091), .Z(n19094) );
  XOR U19334 ( .A(n19093), .B(n19094), .Z(n19105) );
  NANDN U19335 ( .A(n18787), .B(n18786), .Z(n18791) );
  OR U19336 ( .A(n18789), .B(n18788), .Z(n18790) );
  AND U19337 ( .A(n18791), .B(n18790), .Z(n19104) );
  NANDN U19338 ( .A(n18793), .B(n18792), .Z(n18797) );
  OR U19339 ( .A(n18795), .B(n18794), .Z(n18796) );
  AND U19340 ( .A(n18797), .B(n18796), .Z(n19100) );
  NANDN U19341 ( .A(n18799), .B(n18798), .Z(n18803) );
  NANDN U19342 ( .A(n18801), .B(n18800), .Z(n18802) );
  AND U19343 ( .A(n18803), .B(n18802), .Z(n19098) );
  NANDN U19344 ( .A(n18805), .B(n18804), .Z(n18809) );
  OR U19345 ( .A(n18807), .B(n18806), .Z(n18808) );
  AND U19346 ( .A(n18809), .B(n18808), .Z(n19097) );
  XNOR U19347 ( .A(n19098), .B(n19097), .Z(n19099) );
  XNOR U19348 ( .A(n19100), .B(n19099), .Z(n19103) );
  XOR U19349 ( .A(n19104), .B(n19103), .Z(n19106) );
  XOR U19350 ( .A(n19105), .B(n19106), .Z(n19112) );
  NANDN U19351 ( .A(n18811), .B(n18810), .Z(n18815) );
  NANDN U19352 ( .A(n18813), .B(n18812), .Z(n18814) );
  AND U19353 ( .A(n18815), .B(n18814), .Z(n19110) );
  NANDN U19354 ( .A(n18817), .B(n18816), .Z(n18821) );
  OR U19355 ( .A(n18819), .B(n18818), .Z(n18820) );
  AND U19356 ( .A(n18821), .B(n18820), .Z(n19109) );
  XNOR U19357 ( .A(n19110), .B(n19109), .Z(n19111) );
  XNOR U19358 ( .A(n19112), .B(n19111), .Z(n18833) );
  XOR U19359 ( .A(n18834), .B(n18833), .Z(n18836) );
  XNOR U19360 ( .A(n18835), .B(n18836), .Z(n18827) );
  XNOR U19361 ( .A(n18828), .B(n18827), .Z(n18829) );
  XNOR U19362 ( .A(n18830), .B(n18829), .Z(n19115) );
  XNOR U19363 ( .A(sreg[159]), .B(n19115), .Z(n19117) );
  NANDN U19364 ( .A(sreg[158]), .B(n18822), .Z(n18826) );
  NAND U19365 ( .A(n18824), .B(n18823), .Z(n18825) );
  NAND U19366 ( .A(n18826), .B(n18825), .Z(n19116) );
  XNOR U19367 ( .A(n19117), .B(n19116), .Z(c[159]) );
  NANDN U19368 ( .A(n18828), .B(n18827), .Z(n18832) );
  NANDN U19369 ( .A(n18830), .B(n18829), .Z(n18831) );
  AND U19370 ( .A(n18832), .B(n18831), .Z(n19123) );
  NANDN U19371 ( .A(n18834), .B(n18833), .Z(n18838) );
  OR U19372 ( .A(n18836), .B(n18835), .Z(n18837) );
  AND U19373 ( .A(n18838), .B(n18837), .Z(n19120) );
  NANDN U19374 ( .A(n18840), .B(n18839), .Z(n18844) );
  NANDN U19375 ( .A(n18842), .B(n18841), .Z(n18843) );
  AND U19376 ( .A(n18844), .B(n18843), .Z(n19140) );
  NANDN U19377 ( .A(n18846), .B(n18845), .Z(n18850) );
  NAND U19378 ( .A(n18848), .B(n18847), .Z(n18849) );
  AND U19379 ( .A(n18850), .B(n18849), .Z(n19170) );
  NANDN U19380 ( .A(n18852), .B(n18851), .Z(n18856) );
  NANDN U19381 ( .A(n18854), .B(n18853), .Z(n18855) );
  AND U19382 ( .A(n18856), .B(n18855), .Z(n19164) );
  NANDN U19383 ( .A(n18858), .B(n18857), .Z(n18862) );
  NANDN U19384 ( .A(n18860), .B(n18859), .Z(n18861) );
  AND U19385 ( .A(n18862), .B(n18861), .Z(n19163) );
  NANDN U19386 ( .A(n33875), .B(n18863), .Z(n18865) );
  XOR U19387 ( .A(b[25]), .B(a[72]), .Z(n19249) );
  NANDN U19388 ( .A(n33994), .B(n19249), .Z(n18864) );
  AND U19389 ( .A(n18865), .B(n18864), .Z(n19368) );
  NANDN U19390 ( .A(n32013), .B(n18866), .Z(n18868) );
  XOR U19391 ( .A(b[17]), .B(a[80]), .Z(n19252) );
  NANDN U19392 ( .A(n32292), .B(n19252), .Z(n18867) );
  AND U19393 ( .A(n18868), .B(n18867), .Z(n19367) );
  NANDN U19394 ( .A(n31536), .B(n18869), .Z(n18871) );
  XOR U19395 ( .A(a[82]), .B(b[15]), .Z(n19255) );
  NANDN U19396 ( .A(n31925), .B(n19255), .Z(n18870) );
  NAND U19397 ( .A(n18871), .B(n18870), .Z(n19366) );
  XOR U19398 ( .A(n19367), .B(n19366), .Z(n19369) );
  XOR U19399 ( .A(n19368), .B(n19369), .Z(n19340) );
  NANDN U19400 ( .A(n37526), .B(n18872), .Z(n18874) );
  XOR U19401 ( .A(b[51]), .B(a[46]), .Z(n19258) );
  NANDN U19402 ( .A(n37605), .B(n19258), .Z(n18873) );
  AND U19403 ( .A(n18874), .B(n18873), .Z(n19392) );
  NANDN U19404 ( .A(n37705), .B(n18875), .Z(n18877) );
  XOR U19405 ( .A(b[53]), .B(a[44]), .Z(n19261) );
  NANDN U19406 ( .A(n37778), .B(n19261), .Z(n18876) );
  AND U19407 ( .A(n18877), .B(n18876), .Z(n19391) );
  NANDN U19408 ( .A(n36210), .B(n18878), .Z(n18880) );
  XOR U19409 ( .A(b[39]), .B(a[58]), .Z(n19264) );
  NANDN U19410 ( .A(n36347), .B(n19264), .Z(n18879) );
  NAND U19411 ( .A(n18880), .B(n18879), .Z(n19390) );
  XOR U19412 ( .A(n19391), .B(n19390), .Z(n19393) );
  XNOR U19413 ( .A(n19392), .B(n19393), .Z(n19339) );
  XNOR U19414 ( .A(n19340), .B(n19339), .Z(n19342) );
  NANDN U19415 ( .A(n18882), .B(n18881), .Z(n18886) );
  OR U19416 ( .A(n18884), .B(n18883), .Z(n18885) );
  AND U19417 ( .A(n18886), .B(n18885), .Z(n19341) );
  XOR U19418 ( .A(n19342), .B(n19341), .Z(n19240) );
  NANDN U19419 ( .A(n18888), .B(n18887), .Z(n18892) );
  OR U19420 ( .A(n18890), .B(n18889), .Z(n18891) );
  AND U19421 ( .A(n18892), .B(n18891), .Z(n19238) );
  NANDN U19422 ( .A(n18894), .B(n18893), .Z(n18898) );
  NANDN U19423 ( .A(n18896), .B(n18895), .Z(n18897) );
  NAND U19424 ( .A(n18898), .B(n18897), .Z(n19237) );
  XNOR U19425 ( .A(n19238), .B(n19237), .Z(n19239) );
  XNOR U19426 ( .A(n19240), .B(n19239), .Z(n19162) );
  XOR U19427 ( .A(n19163), .B(n19162), .Z(n19165) );
  XOR U19428 ( .A(n19164), .B(n19165), .Z(n19169) );
  NANDN U19429 ( .A(n18900), .B(n18899), .Z(n18904) );
  NANDN U19430 ( .A(n18902), .B(n18901), .Z(n18903) );
  AND U19431 ( .A(n18904), .B(n18903), .Z(n19157) );
  NANDN U19432 ( .A(n211), .B(n18905), .Z(n18907) );
  XOR U19433 ( .A(b[47]), .B(a[50]), .Z(n19192) );
  NANDN U19434 ( .A(n37172), .B(n19192), .Z(n18906) );
  AND U19435 ( .A(n18907), .B(n18906), .Z(n19233) );
  NANDN U19436 ( .A(n210), .B(n18908), .Z(n18910) );
  XOR U19437 ( .A(a[88]), .B(b[9]), .Z(n19195) );
  NANDN U19438 ( .A(n30267), .B(n19195), .Z(n18909) );
  AND U19439 ( .A(n18910), .B(n18909), .Z(n19232) );
  NANDN U19440 ( .A(n212), .B(n18911), .Z(n18913) );
  XOR U19441 ( .A(b[49]), .B(a[48]), .Z(n19198) );
  NANDN U19442 ( .A(n37432), .B(n19198), .Z(n18912) );
  NAND U19443 ( .A(n18913), .B(n18912), .Z(n19231) );
  XOR U19444 ( .A(n19232), .B(n19231), .Z(n19234) );
  XOR U19445 ( .A(n19233), .B(n19234), .Z(n19346) );
  NANDN U19446 ( .A(n36742), .B(n18914), .Z(n18916) );
  XOR U19447 ( .A(b[43]), .B(a[54]), .Z(n19201) );
  NANDN U19448 ( .A(n36891), .B(n19201), .Z(n18915) );
  AND U19449 ( .A(n18916), .B(n18915), .Z(n19212) );
  NANDN U19450 ( .A(n36991), .B(n18917), .Z(n18919) );
  XOR U19451 ( .A(b[45]), .B(a[52]), .Z(n19204) );
  NANDN U19452 ( .A(n37083), .B(n19204), .Z(n18918) );
  AND U19453 ( .A(n18919), .B(n18918), .Z(n19211) );
  NANDN U19454 ( .A(n30482), .B(n18920), .Z(n18922) );
  XOR U19455 ( .A(a[86]), .B(b[11]), .Z(n19207) );
  NANDN U19456 ( .A(n30891), .B(n19207), .Z(n18921) );
  NAND U19457 ( .A(n18922), .B(n18921), .Z(n19210) );
  XOR U19458 ( .A(n19211), .B(n19210), .Z(n19213) );
  XNOR U19459 ( .A(n19212), .B(n19213), .Z(n19345) );
  XNOR U19460 ( .A(n19346), .B(n19345), .Z(n19347) );
  NANDN U19461 ( .A(n18924), .B(n18923), .Z(n18928) );
  OR U19462 ( .A(n18926), .B(n18925), .Z(n18927) );
  NAND U19463 ( .A(n18928), .B(n18927), .Z(n19348) );
  XNOR U19464 ( .A(n19347), .B(n19348), .Z(n19156) );
  XNOR U19465 ( .A(n19157), .B(n19156), .Z(n19158) );
  NANDN U19466 ( .A(n29499), .B(n18929), .Z(n18931) );
  XOR U19467 ( .A(a[90]), .B(b[7]), .Z(n19216) );
  NANDN U19468 ( .A(n29735), .B(n19216), .Z(n18930) );
  AND U19469 ( .A(n18931), .B(n18930), .Z(n19275) );
  NANDN U19470 ( .A(n37857), .B(n18932), .Z(n18934) );
  XOR U19471 ( .A(b[55]), .B(a[42]), .Z(n19219) );
  NANDN U19472 ( .A(n37911), .B(n19219), .Z(n18933) );
  AND U19473 ( .A(n18934), .B(n18933), .Z(n19274) );
  NANDN U19474 ( .A(n35611), .B(n18935), .Z(n18937) );
  XOR U19475 ( .A(b[35]), .B(a[62]), .Z(n19222) );
  NANDN U19476 ( .A(n35801), .B(n19222), .Z(n18936) );
  NAND U19477 ( .A(n18937), .B(n18936), .Z(n19273) );
  XOR U19478 ( .A(n19274), .B(n19273), .Z(n19276) );
  XOR U19479 ( .A(n19275), .B(n19276), .Z(n19286) );
  NANDN U19480 ( .A(n18939), .B(n18938), .Z(n18943) );
  OR U19481 ( .A(n18941), .B(n18940), .Z(n18942) );
  AND U19482 ( .A(n18943), .B(n18942), .Z(n19285) );
  XNOR U19483 ( .A(n19286), .B(n19285), .Z(n19287) );
  NANDN U19484 ( .A(n18945), .B(n18944), .Z(n18949) );
  OR U19485 ( .A(n18947), .B(n18946), .Z(n18948) );
  NAND U19486 ( .A(n18949), .B(n18948), .Z(n19288) );
  XOR U19487 ( .A(n19287), .B(n19288), .Z(n19159) );
  XNOR U19488 ( .A(n19158), .B(n19159), .Z(n19168) );
  XOR U19489 ( .A(n19169), .B(n19168), .Z(n19171) );
  XOR U19490 ( .A(n19170), .B(n19171), .Z(n19139) );
  NANDN U19491 ( .A(n18951), .B(n18950), .Z(n18955) );
  NANDN U19492 ( .A(n18953), .B(n18952), .Z(n18954) );
  AND U19493 ( .A(n18955), .B(n18954), .Z(n19152) );
  NANDN U19494 ( .A(n18957), .B(n18956), .Z(n18961) );
  NANDN U19495 ( .A(n18959), .B(n18958), .Z(n18960) );
  AND U19496 ( .A(n18961), .B(n18960), .Z(n19151) );
  NANDN U19497 ( .A(n18963), .B(n18962), .Z(n18967) );
  NAND U19498 ( .A(n18965), .B(n18964), .Z(n18966) );
  AND U19499 ( .A(n18967), .B(n18966), .Z(n19150) );
  XOR U19500 ( .A(n19151), .B(n19150), .Z(n19153) );
  XOR U19501 ( .A(n19152), .B(n19153), .Z(n19177) );
  NANDN U19502 ( .A(n18969), .B(n18968), .Z(n18973) );
  NANDN U19503 ( .A(n18971), .B(n18970), .Z(n18972) );
  AND U19504 ( .A(n18973), .B(n18972), .Z(n19298) );
  NANDN U19505 ( .A(n18975), .B(n18974), .Z(n18979) );
  OR U19506 ( .A(n18977), .B(n18976), .Z(n18978) );
  NAND U19507 ( .A(n18979), .B(n18978), .Z(n19297) );
  XNOR U19508 ( .A(n19298), .B(n19297), .Z(n19300) );
  NANDN U19509 ( .A(n18981), .B(n18980), .Z(n18985) );
  OR U19510 ( .A(n18983), .B(n18982), .Z(n18984) );
  AND U19511 ( .A(n18985), .B(n18984), .Z(n19246) );
  NAND U19512 ( .A(b[0]), .B(a[96]), .Z(n18986) );
  XNOR U19513 ( .A(b[1]), .B(n18986), .Z(n18988) );
  NANDN U19514 ( .A(b[0]), .B(a[95]), .Z(n18987) );
  NAND U19515 ( .A(n18988), .B(n18987), .Z(n19282) );
  NANDN U19516 ( .A(n38278), .B(n18989), .Z(n18991) );
  XOR U19517 ( .A(b[63]), .B(a[34]), .Z(n19324) );
  NANDN U19518 ( .A(n38279), .B(n19324), .Z(n18990) );
  AND U19519 ( .A(n18991), .B(n18990), .Z(n19280) );
  NANDN U19520 ( .A(n35260), .B(n18992), .Z(n18994) );
  XOR U19521 ( .A(b[33]), .B(a[64]), .Z(n19327) );
  NANDN U19522 ( .A(n35456), .B(n19327), .Z(n18993) );
  NAND U19523 ( .A(n18994), .B(n18993), .Z(n19279) );
  XNOR U19524 ( .A(n19280), .B(n19279), .Z(n19281) );
  XNOR U19525 ( .A(n19282), .B(n19281), .Z(n19243) );
  NANDN U19526 ( .A(n37974), .B(n18995), .Z(n18997) );
  XOR U19527 ( .A(b[57]), .B(a[40]), .Z(n19330) );
  NANDN U19528 ( .A(n38031), .B(n19330), .Z(n18996) );
  AND U19529 ( .A(n18997), .B(n18996), .Z(n19306) );
  NANDN U19530 ( .A(n38090), .B(n18998), .Z(n19000) );
  XOR U19531 ( .A(b[59]), .B(a[38]), .Z(n19333) );
  NANDN U19532 ( .A(n38130), .B(n19333), .Z(n18999) );
  AND U19533 ( .A(n19000), .B(n18999), .Z(n19304) );
  NANDN U19534 ( .A(n36480), .B(n19001), .Z(n19003) );
  XOR U19535 ( .A(b[41]), .B(a[56]), .Z(n19336) );
  NANDN U19536 ( .A(n36594), .B(n19336), .Z(n19002) );
  NAND U19537 ( .A(n19003), .B(n19002), .Z(n19303) );
  XNOR U19538 ( .A(n19304), .B(n19303), .Z(n19305) );
  XOR U19539 ( .A(n19306), .B(n19305), .Z(n19244) );
  XNOR U19540 ( .A(n19243), .B(n19244), .Z(n19245) );
  XNOR U19541 ( .A(n19246), .B(n19245), .Z(n19299) );
  XOR U19542 ( .A(n19300), .B(n19299), .Z(n19181) );
  NANDN U19543 ( .A(n19005), .B(n19004), .Z(n19009) );
  NAND U19544 ( .A(n19007), .B(n19006), .Z(n19008) );
  NAND U19545 ( .A(n19009), .B(n19008), .Z(n19180) );
  XNOR U19546 ( .A(n19181), .B(n19180), .Z(n19183) );
  NANDN U19547 ( .A(n19011), .B(n19010), .Z(n19015) );
  NANDN U19548 ( .A(n19013), .B(n19012), .Z(n19014) );
  AND U19549 ( .A(n19015), .B(n19014), .Z(n19399) );
  NANDN U19550 ( .A(n32996), .B(n19016), .Z(n19018) );
  XOR U19551 ( .A(b[21]), .B(a[76]), .Z(n19351) );
  NANDN U19552 ( .A(n33271), .B(n19351), .Z(n19017) );
  AND U19553 ( .A(n19018), .B(n19017), .Z(n19317) );
  NANDN U19554 ( .A(n33866), .B(n19019), .Z(n19021) );
  XOR U19555 ( .A(b[23]), .B(a[74]), .Z(n19354) );
  NANDN U19556 ( .A(n33644), .B(n19354), .Z(n19020) );
  AND U19557 ( .A(n19021), .B(n19020), .Z(n19316) );
  NANDN U19558 ( .A(n32483), .B(n19022), .Z(n19024) );
  XOR U19559 ( .A(b[19]), .B(a[78]), .Z(n19357) );
  NANDN U19560 ( .A(n32823), .B(n19357), .Z(n19023) );
  NAND U19561 ( .A(n19024), .B(n19023), .Z(n19315) );
  XOR U19562 ( .A(n19316), .B(n19315), .Z(n19318) );
  XOR U19563 ( .A(n19317), .B(n19318), .Z(n19187) );
  NANDN U19564 ( .A(n34909), .B(n19025), .Z(n19027) );
  XOR U19565 ( .A(b[31]), .B(a[66]), .Z(n19360) );
  NANDN U19566 ( .A(n35145), .B(n19360), .Z(n19026) );
  AND U19567 ( .A(n19027), .B(n19026), .Z(n19227) );
  NANDN U19568 ( .A(n38247), .B(n19028), .Z(n19030) );
  XOR U19569 ( .A(b[61]), .B(a[36]), .Z(n19363) );
  NANDN U19570 ( .A(n38248), .B(n19363), .Z(n19029) );
  AND U19571 ( .A(n19030), .B(n19029), .Z(n19226) );
  AND U19572 ( .A(b[63]), .B(a[32]), .Z(n19225) );
  XOR U19573 ( .A(n19226), .B(n19225), .Z(n19228) );
  XNOR U19574 ( .A(n19227), .B(n19228), .Z(n19186) );
  XNOR U19575 ( .A(n19187), .B(n19186), .Z(n19188) );
  NANDN U19576 ( .A(n19032), .B(n19031), .Z(n19036) );
  OR U19577 ( .A(n19034), .B(n19033), .Z(n19035) );
  NAND U19578 ( .A(n19036), .B(n19035), .Z(n19189) );
  XNOR U19579 ( .A(n19188), .B(n19189), .Z(n19396) );
  NANDN U19580 ( .A(n34223), .B(n19037), .Z(n19039) );
  XOR U19581 ( .A(b[27]), .B(a[70]), .Z(n19372) );
  NANDN U19582 ( .A(n34458), .B(n19372), .Z(n19038) );
  AND U19583 ( .A(n19039), .B(n19038), .Z(n19269) );
  NANDN U19584 ( .A(n34634), .B(n19040), .Z(n19042) );
  XOR U19585 ( .A(b[29]), .B(a[68]), .Z(n19375) );
  NANDN U19586 ( .A(n34722), .B(n19375), .Z(n19041) );
  AND U19587 ( .A(n19042), .B(n19041), .Z(n19268) );
  NANDN U19588 ( .A(n31055), .B(n19043), .Z(n19045) );
  XOR U19589 ( .A(a[84]), .B(b[13]), .Z(n19378) );
  NANDN U19590 ( .A(n31293), .B(n19378), .Z(n19044) );
  NAND U19591 ( .A(n19045), .B(n19044), .Z(n19267) );
  XOR U19592 ( .A(n19268), .B(n19267), .Z(n19270) );
  XOR U19593 ( .A(n19269), .B(n19270), .Z(n19292) );
  NANDN U19594 ( .A(n28889), .B(n19046), .Z(n19048) );
  XOR U19595 ( .A(a[92]), .B(b[5]), .Z(n19381) );
  NANDN U19596 ( .A(n29138), .B(n19381), .Z(n19047) );
  AND U19597 ( .A(n19048), .B(n19047), .Z(n19311) );
  NANDN U19598 ( .A(n209), .B(n19049), .Z(n19051) );
  XOR U19599 ( .A(a[94]), .B(b[3]), .Z(n19384) );
  NANDN U19600 ( .A(n28941), .B(n19384), .Z(n19050) );
  AND U19601 ( .A(n19051), .B(n19050), .Z(n19310) );
  NANDN U19602 ( .A(n35936), .B(n19052), .Z(n19054) );
  XOR U19603 ( .A(b[37]), .B(a[60]), .Z(n19387) );
  NANDN U19604 ( .A(n36047), .B(n19387), .Z(n19053) );
  NAND U19605 ( .A(n19054), .B(n19053), .Z(n19309) );
  XOR U19606 ( .A(n19310), .B(n19309), .Z(n19312) );
  XNOR U19607 ( .A(n19311), .B(n19312), .Z(n19291) );
  XNOR U19608 ( .A(n19292), .B(n19291), .Z(n19293) );
  NANDN U19609 ( .A(n19056), .B(n19055), .Z(n19060) );
  OR U19610 ( .A(n19058), .B(n19057), .Z(n19059) );
  NAND U19611 ( .A(n19060), .B(n19059), .Z(n19294) );
  XOR U19612 ( .A(n19293), .B(n19294), .Z(n19397) );
  XNOR U19613 ( .A(n19396), .B(n19397), .Z(n19398) );
  XNOR U19614 ( .A(n19399), .B(n19398), .Z(n19182) );
  XOR U19615 ( .A(n19183), .B(n19182), .Z(n19175) );
  NANDN U19616 ( .A(n19062), .B(n19061), .Z(n19066) );
  NANDN U19617 ( .A(n19064), .B(n19063), .Z(n19065) );
  AND U19618 ( .A(n19066), .B(n19065), .Z(n19174) );
  XNOR U19619 ( .A(n19175), .B(n19174), .Z(n19176) );
  XNOR U19620 ( .A(n19177), .B(n19176), .Z(n19138) );
  XOR U19621 ( .A(n19139), .B(n19138), .Z(n19141) );
  XOR U19622 ( .A(n19140), .B(n19141), .Z(n19134) );
  NANDN U19623 ( .A(n19068), .B(n19067), .Z(n19072) );
  OR U19624 ( .A(n19070), .B(n19069), .Z(n19071) );
  AND U19625 ( .A(n19072), .B(n19071), .Z(n19133) );
  NANDN U19626 ( .A(n19074), .B(n19073), .Z(n19078) );
  OR U19627 ( .A(n19076), .B(n19075), .Z(n19077) );
  AND U19628 ( .A(n19078), .B(n19077), .Z(n19147) );
  NANDN U19629 ( .A(n19080), .B(n19079), .Z(n19084) );
  NANDN U19630 ( .A(n19082), .B(n19081), .Z(n19083) );
  AND U19631 ( .A(n19084), .B(n19083), .Z(n19145) );
  NANDN U19632 ( .A(n19086), .B(n19085), .Z(n19090) );
  OR U19633 ( .A(n19088), .B(n19087), .Z(n19089) );
  AND U19634 ( .A(n19090), .B(n19089), .Z(n19144) );
  XNOR U19635 ( .A(n19145), .B(n19144), .Z(n19146) );
  XNOR U19636 ( .A(n19147), .B(n19146), .Z(n19132) );
  XOR U19637 ( .A(n19133), .B(n19132), .Z(n19135) );
  XOR U19638 ( .A(n19134), .B(n19135), .Z(n19128) );
  NANDN U19639 ( .A(n19092), .B(n19091), .Z(n19096) );
  OR U19640 ( .A(n19094), .B(n19093), .Z(n19095) );
  AND U19641 ( .A(n19096), .B(n19095), .Z(n19127) );
  NANDN U19642 ( .A(n19098), .B(n19097), .Z(n19102) );
  NANDN U19643 ( .A(n19100), .B(n19099), .Z(n19101) );
  AND U19644 ( .A(n19102), .B(n19101), .Z(n19126) );
  XOR U19645 ( .A(n19127), .B(n19126), .Z(n19129) );
  XOR U19646 ( .A(n19128), .B(n19129), .Z(n19403) );
  NANDN U19647 ( .A(n19104), .B(n19103), .Z(n19108) );
  OR U19648 ( .A(n19106), .B(n19105), .Z(n19107) );
  NAND U19649 ( .A(n19108), .B(n19107), .Z(n19402) );
  XNOR U19650 ( .A(n19403), .B(n19402), .Z(n19404) );
  NANDN U19651 ( .A(n19110), .B(n19109), .Z(n19114) );
  NANDN U19652 ( .A(n19112), .B(n19111), .Z(n19113) );
  NAND U19653 ( .A(n19114), .B(n19113), .Z(n19405) );
  XOR U19654 ( .A(n19404), .B(n19405), .Z(n19121) );
  XNOR U19655 ( .A(n19120), .B(n19121), .Z(n19122) );
  XNOR U19656 ( .A(n19123), .B(n19122), .Z(n19408) );
  XNOR U19657 ( .A(sreg[160]), .B(n19408), .Z(n19410) );
  NANDN U19658 ( .A(sreg[159]), .B(n19115), .Z(n19119) );
  NAND U19659 ( .A(n19117), .B(n19116), .Z(n19118) );
  NAND U19660 ( .A(n19119), .B(n19118), .Z(n19409) );
  XNOR U19661 ( .A(n19410), .B(n19409), .Z(c[160]) );
  NANDN U19662 ( .A(n19121), .B(n19120), .Z(n19125) );
  NANDN U19663 ( .A(n19123), .B(n19122), .Z(n19124) );
  AND U19664 ( .A(n19125), .B(n19124), .Z(n19416) );
  NANDN U19665 ( .A(n19127), .B(n19126), .Z(n19131) );
  OR U19666 ( .A(n19129), .B(n19128), .Z(n19130) );
  AND U19667 ( .A(n19131), .B(n19130), .Z(n19697) );
  NANDN U19668 ( .A(n19133), .B(n19132), .Z(n19137) );
  OR U19669 ( .A(n19135), .B(n19134), .Z(n19136) );
  AND U19670 ( .A(n19137), .B(n19136), .Z(n19695) );
  NANDN U19671 ( .A(n19139), .B(n19138), .Z(n19143) );
  OR U19672 ( .A(n19141), .B(n19140), .Z(n19142) );
  AND U19673 ( .A(n19143), .B(n19142), .Z(n19690) );
  NANDN U19674 ( .A(n19145), .B(n19144), .Z(n19149) );
  NANDN U19675 ( .A(n19147), .B(n19146), .Z(n19148) );
  AND U19676 ( .A(n19149), .B(n19148), .Z(n19689) );
  XNOR U19677 ( .A(n19690), .B(n19689), .Z(n19691) );
  NANDN U19678 ( .A(n19151), .B(n19150), .Z(n19155) );
  OR U19679 ( .A(n19153), .B(n19152), .Z(n19154) );
  AND U19680 ( .A(n19155), .B(n19154), .Z(n19679) );
  NANDN U19681 ( .A(n19157), .B(n19156), .Z(n19161) );
  NANDN U19682 ( .A(n19159), .B(n19158), .Z(n19160) );
  AND U19683 ( .A(n19161), .B(n19160), .Z(n19678) );
  NANDN U19684 ( .A(n19163), .B(n19162), .Z(n19167) );
  OR U19685 ( .A(n19165), .B(n19164), .Z(n19166) );
  AND U19686 ( .A(n19167), .B(n19166), .Z(n19677) );
  XOR U19687 ( .A(n19678), .B(n19677), .Z(n19680) );
  XOR U19688 ( .A(n19679), .B(n19680), .Z(n19684) );
  NANDN U19689 ( .A(n19169), .B(n19168), .Z(n19173) );
  OR U19690 ( .A(n19171), .B(n19170), .Z(n19172) );
  AND U19691 ( .A(n19173), .B(n19172), .Z(n19683) );
  XNOR U19692 ( .A(n19684), .B(n19683), .Z(n19685) );
  NANDN U19693 ( .A(n19175), .B(n19174), .Z(n19179) );
  NANDN U19694 ( .A(n19177), .B(n19176), .Z(n19178) );
  AND U19695 ( .A(n19179), .B(n19178), .Z(n19674) );
  NANDN U19696 ( .A(n19181), .B(n19180), .Z(n19185) );
  NAND U19697 ( .A(n19183), .B(n19182), .Z(n19184) );
  AND U19698 ( .A(n19185), .B(n19184), .Z(n19439) );
  NANDN U19699 ( .A(n19187), .B(n19186), .Z(n19191) );
  NANDN U19700 ( .A(n19189), .B(n19188), .Z(n19190) );
  AND U19701 ( .A(n19191), .B(n19190), .Z(n19426) );
  NANDN U19702 ( .A(n211), .B(n19192), .Z(n19194) );
  XOR U19703 ( .A(b[47]), .B(a[51]), .Z(n19509) );
  NANDN U19704 ( .A(n37172), .B(n19509), .Z(n19193) );
  AND U19705 ( .A(n19194), .B(n19193), .Z(n19550) );
  NANDN U19706 ( .A(n210), .B(n19195), .Z(n19197) );
  XOR U19707 ( .A(a[89]), .B(b[9]), .Z(n19512) );
  NANDN U19708 ( .A(n30267), .B(n19512), .Z(n19196) );
  AND U19709 ( .A(n19197), .B(n19196), .Z(n19549) );
  NANDN U19710 ( .A(n212), .B(n19198), .Z(n19200) );
  XOR U19711 ( .A(b[49]), .B(a[49]), .Z(n19515) );
  NANDN U19712 ( .A(n37432), .B(n19515), .Z(n19199) );
  NAND U19713 ( .A(n19200), .B(n19199), .Z(n19548) );
  XOR U19714 ( .A(n19549), .B(n19548), .Z(n19551) );
  XOR U19715 ( .A(n19550), .B(n19551), .Z(n19615) );
  NANDN U19716 ( .A(n36742), .B(n19201), .Z(n19203) );
  XOR U19717 ( .A(b[43]), .B(a[55]), .Z(n19518) );
  NANDN U19718 ( .A(n36891), .B(n19518), .Z(n19202) );
  AND U19719 ( .A(n19203), .B(n19202), .Z(n19529) );
  NANDN U19720 ( .A(n36991), .B(n19204), .Z(n19206) );
  XOR U19721 ( .A(b[45]), .B(a[53]), .Z(n19521) );
  NANDN U19722 ( .A(n37083), .B(n19521), .Z(n19205) );
  AND U19723 ( .A(n19206), .B(n19205), .Z(n19528) );
  NANDN U19724 ( .A(n30482), .B(n19207), .Z(n19209) );
  XOR U19725 ( .A(a[87]), .B(b[11]), .Z(n19524) );
  NANDN U19726 ( .A(n30891), .B(n19524), .Z(n19208) );
  NAND U19727 ( .A(n19209), .B(n19208), .Z(n19527) );
  XOR U19728 ( .A(n19528), .B(n19527), .Z(n19530) );
  XNOR U19729 ( .A(n19529), .B(n19530), .Z(n19614) );
  XNOR U19730 ( .A(n19615), .B(n19614), .Z(n19616) );
  NANDN U19731 ( .A(n19211), .B(n19210), .Z(n19215) );
  OR U19732 ( .A(n19213), .B(n19212), .Z(n19214) );
  NAND U19733 ( .A(n19215), .B(n19214), .Z(n19617) );
  XNOR U19734 ( .A(n19616), .B(n19617), .Z(n19425) );
  XNOR U19735 ( .A(n19426), .B(n19425), .Z(n19428) );
  NANDN U19736 ( .A(n29499), .B(n19216), .Z(n19218) );
  XOR U19737 ( .A(a[91]), .B(b[7]), .Z(n19533) );
  NANDN U19738 ( .A(n29735), .B(n19533), .Z(n19217) );
  AND U19739 ( .A(n19218), .B(n19217), .Z(n19493) );
  NANDN U19740 ( .A(n37857), .B(n19219), .Z(n19221) );
  XOR U19741 ( .A(b[55]), .B(a[43]), .Z(n19536) );
  NANDN U19742 ( .A(n37911), .B(n19536), .Z(n19220) );
  AND U19743 ( .A(n19221), .B(n19220), .Z(n19492) );
  NANDN U19744 ( .A(n35611), .B(n19222), .Z(n19224) );
  XOR U19745 ( .A(b[35]), .B(a[63]), .Z(n19539) );
  NANDN U19746 ( .A(n35801), .B(n19539), .Z(n19223) );
  NAND U19747 ( .A(n19224), .B(n19223), .Z(n19491) );
  XOR U19748 ( .A(n19492), .B(n19491), .Z(n19494) );
  XOR U19749 ( .A(n19493), .B(n19494), .Z(n19555) );
  NANDN U19750 ( .A(n19226), .B(n19225), .Z(n19230) );
  OR U19751 ( .A(n19228), .B(n19227), .Z(n19229) );
  AND U19752 ( .A(n19230), .B(n19229), .Z(n19554) );
  XNOR U19753 ( .A(n19555), .B(n19554), .Z(n19556) );
  NANDN U19754 ( .A(n19232), .B(n19231), .Z(n19236) );
  OR U19755 ( .A(n19234), .B(n19233), .Z(n19235) );
  NAND U19756 ( .A(n19236), .B(n19235), .Z(n19557) );
  XNOR U19757 ( .A(n19556), .B(n19557), .Z(n19427) );
  XOR U19758 ( .A(n19428), .B(n19427), .Z(n19438) );
  NANDN U19759 ( .A(n19238), .B(n19237), .Z(n19242) );
  NANDN U19760 ( .A(n19240), .B(n19239), .Z(n19241) );
  AND U19761 ( .A(n19242), .B(n19241), .Z(n19434) );
  NANDN U19762 ( .A(n19244), .B(n19243), .Z(n19248) );
  NANDN U19763 ( .A(n19246), .B(n19245), .Z(n19247) );
  AND U19764 ( .A(n19248), .B(n19247), .Z(n19432) );
  NANDN U19765 ( .A(n33875), .B(n19249), .Z(n19251) );
  XOR U19766 ( .A(b[25]), .B(a[73]), .Z(n19467) );
  NANDN U19767 ( .A(n33994), .B(n19467), .Z(n19250) );
  AND U19768 ( .A(n19251), .B(n19250), .Z(n19637) );
  NANDN U19769 ( .A(n32013), .B(n19252), .Z(n19254) );
  XOR U19770 ( .A(b[17]), .B(a[81]), .Z(n19470) );
  NANDN U19771 ( .A(n32292), .B(n19470), .Z(n19253) );
  AND U19772 ( .A(n19254), .B(n19253), .Z(n19636) );
  NANDN U19773 ( .A(n31536), .B(n19255), .Z(n19257) );
  XOR U19774 ( .A(a[83]), .B(b[15]), .Z(n19473) );
  NANDN U19775 ( .A(n31925), .B(n19473), .Z(n19256) );
  NAND U19776 ( .A(n19257), .B(n19256), .Z(n19635) );
  XOR U19777 ( .A(n19636), .B(n19635), .Z(n19638) );
  XOR U19778 ( .A(n19637), .B(n19638), .Z(n19609) );
  NANDN U19779 ( .A(n37526), .B(n19258), .Z(n19260) );
  XOR U19780 ( .A(b[51]), .B(a[47]), .Z(n19476) );
  NANDN U19781 ( .A(n37605), .B(n19476), .Z(n19259) );
  AND U19782 ( .A(n19260), .B(n19259), .Z(n19661) );
  NANDN U19783 ( .A(n37705), .B(n19261), .Z(n19263) );
  XOR U19784 ( .A(b[53]), .B(a[45]), .Z(n19479) );
  NANDN U19785 ( .A(n37778), .B(n19479), .Z(n19262) );
  AND U19786 ( .A(n19263), .B(n19262), .Z(n19660) );
  NANDN U19787 ( .A(n36210), .B(n19264), .Z(n19266) );
  XOR U19788 ( .A(b[39]), .B(a[59]), .Z(n19482) );
  NANDN U19789 ( .A(n36347), .B(n19482), .Z(n19265) );
  NAND U19790 ( .A(n19266), .B(n19265), .Z(n19659) );
  XOR U19791 ( .A(n19660), .B(n19659), .Z(n19662) );
  XNOR U19792 ( .A(n19661), .B(n19662), .Z(n19608) );
  XNOR U19793 ( .A(n19609), .B(n19608), .Z(n19611) );
  NANDN U19794 ( .A(n19268), .B(n19267), .Z(n19272) );
  OR U19795 ( .A(n19270), .B(n19269), .Z(n19271) );
  AND U19796 ( .A(n19272), .B(n19271), .Z(n19610) );
  XOR U19797 ( .A(n19611), .B(n19610), .Z(n19458) );
  NANDN U19798 ( .A(n19274), .B(n19273), .Z(n19278) );
  OR U19799 ( .A(n19276), .B(n19275), .Z(n19277) );
  AND U19800 ( .A(n19278), .B(n19277), .Z(n19456) );
  NANDN U19801 ( .A(n19280), .B(n19279), .Z(n19284) );
  NANDN U19802 ( .A(n19282), .B(n19281), .Z(n19283) );
  NAND U19803 ( .A(n19284), .B(n19283), .Z(n19455) );
  XNOR U19804 ( .A(n19456), .B(n19455), .Z(n19457) );
  XNOR U19805 ( .A(n19458), .B(n19457), .Z(n19431) );
  XNOR U19806 ( .A(n19432), .B(n19431), .Z(n19433) );
  XNOR U19807 ( .A(n19434), .B(n19433), .Z(n19437) );
  XOR U19808 ( .A(n19438), .B(n19437), .Z(n19440) );
  XNOR U19809 ( .A(n19439), .B(n19440), .Z(n19671) );
  NANDN U19810 ( .A(n19286), .B(n19285), .Z(n19290) );
  NANDN U19811 ( .A(n19288), .B(n19287), .Z(n19289) );
  AND U19812 ( .A(n19290), .B(n19289), .Z(n19421) );
  NANDN U19813 ( .A(n19292), .B(n19291), .Z(n19296) );
  NANDN U19814 ( .A(n19294), .B(n19293), .Z(n19295) );
  AND U19815 ( .A(n19296), .B(n19295), .Z(n19420) );
  NANDN U19816 ( .A(n19298), .B(n19297), .Z(n19302) );
  NAND U19817 ( .A(n19300), .B(n19299), .Z(n19301) );
  AND U19818 ( .A(n19302), .B(n19301), .Z(n19419) );
  XOR U19819 ( .A(n19420), .B(n19419), .Z(n19422) );
  XOR U19820 ( .A(n19421), .B(n19422), .Z(n19446) );
  NANDN U19821 ( .A(n19304), .B(n19303), .Z(n19308) );
  NANDN U19822 ( .A(n19306), .B(n19305), .Z(n19307) );
  AND U19823 ( .A(n19308), .B(n19307), .Z(n19567) );
  NANDN U19824 ( .A(n19310), .B(n19309), .Z(n19314) );
  OR U19825 ( .A(n19312), .B(n19311), .Z(n19313) );
  NAND U19826 ( .A(n19314), .B(n19313), .Z(n19566) );
  XNOR U19827 ( .A(n19567), .B(n19566), .Z(n19569) );
  NANDN U19828 ( .A(n19316), .B(n19315), .Z(n19320) );
  OR U19829 ( .A(n19318), .B(n19317), .Z(n19319) );
  AND U19830 ( .A(n19320), .B(n19319), .Z(n19464) );
  NAND U19831 ( .A(b[0]), .B(a[97]), .Z(n19321) );
  XNOR U19832 ( .A(b[1]), .B(n19321), .Z(n19323) );
  NANDN U19833 ( .A(b[0]), .B(a[96]), .Z(n19322) );
  NAND U19834 ( .A(n19323), .B(n19322), .Z(n19500) );
  NANDN U19835 ( .A(n38278), .B(n19324), .Z(n19326) );
  XOR U19836 ( .A(b[63]), .B(a[35]), .Z(n19593) );
  NANDN U19837 ( .A(n38279), .B(n19593), .Z(n19325) );
  AND U19838 ( .A(n19326), .B(n19325), .Z(n19498) );
  NANDN U19839 ( .A(n35260), .B(n19327), .Z(n19329) );
  XOR U19840 ( .A(b[33]), .B(a[65]), .Z(n19596) );
  NANDN U19841 ( .A(n35456), .B(n19596), .Z(n19328) );
  NAND U19842 ( .A(n19329), .B(n19328), .Z(n19497) );
  XNOR U19843 ( .A(n19498), .B(n19497), .Z(n19499) );
  XNOR U19844 ( .A(n19500), .B(n19499), .Z(n19461) );
  NANDN U19845 ( .A(n37974), .B(n19330), .Z(n19332) );
  XOR U19846 ( .A(b[57]), .B(a[41]), .Z(n19599) );
  NANDN U19847 ( .A(n38031), .B(n19599), .Z(n19331) );
  AND U19848 ( .A(n19332), .B(n19331), .Z(n19575) );
  NANDN U19849 ( .A(n38090), .B(n19333), .Z(n19335) );
  XOR U19850 ( .A(b[59]), .B(a[39]), .Z(n19602) );
  NANDN U19851 ( .A(n38130), .B(n19602), .Z(n19334) );
  AND U19852 ( .A(n19335), .B(n19334), .Z(n19573) );
  NANDN U19853 ( .A(n36480), .B(n19336), .Z(n19338) );
  XOR U19854 ( .A(b[41]), .B(a[57]), .Z(n19605) );
  NANDN U19855 ( .A(n36594), .B(n19605), .Z(n19337) );
  NAND U19856 ( .A(n19338), .B(n19337), .Z(n19572) );
  XNOR U19857 ( .A(n19573), .B(n19572), .Z(n19574) );
  XOR U19858 ( .A(n19575), .B(n19574), .Z(n19462) );
  XNOR U19859 ( .A(n19461), .B(n19462), .Z(n19463) );
  XNOR U19860 ( .A(n19464), .B(n19463), .Z(n19568) );
  XOR U19861 ( .A(n19569), .B(n19568), .Z(n19450) );
  NANDN U19862 ( .A(n19340), .B(n19339), .Z(n19344) );
  NAND U19863 ( .A(n19342), .B(n19341), .Z(n19343) );
  NAND U19864 ( .A(n19344), .B(n19343), .Z(n19449) );
  XNOR U19865 ( .A(n19450), .B(n19449), .Z(n19452) );
  NANDN U19866 ( .A(n19346), .B(n19345), .Z(n19350) );
  NANDN U19867 ( .A(n19348), .B(n19347), .Z(n19349) );
  AND U19868 ( .A(n19350), .B(n19349), .Z(n19668) );
  NANDN U19869 ( .A(n32996), .B(n19351), .Z(n19353) );
  XOR U19870 ( .A(b[21]), .B(a[77]), .Z(n19620) );
  NANDN U19871 ( .A(n33271), .B(n19620), .Z(n19352) );
  AND U19872 ( .A(n19353), .B(n19352), .Z(n19586) );
  NANDN U19873 ( .A(n33866), .B(n19354), .Z(n19356) );
  XOR U19874 ( .A(b[23]), .B(a[75]), .Z(n19623) );
  NANDN U19875 ( .A(n33644), .B(n19623), .Z(n19355) );
  AND U19876 ( .A(n19356), .B(n19355), .Z(n19585) );
  NANDN U19877 ( .A(n32483), .B(n19357), .Z(n19359) );
  XOR U19878 ( .A(b[19]), .B(a[79]), .Z(n19626) );
  NANDN U19879 ( .A(n32823), .B(n19626), .Z(n19358) );
  NAND U19880 ( .A(n19359), .B(n19358), .Z(n19584) );
  XOR U19881 ( .A(n19585), .B(n19584), .Z(n19587) );
  XOR U19882 ( .A(n19586), .B(n19587), .Z(n19504) );
  NANDN U19883 ( .A(n34909), .B(n19360), .Z(n19362) );
  XOR U19884 ( .A(b[31]), .B(a[67]), .Z(n19629) );
  NANDN U19885 ( .A(n35145), .B(n19629), .Z(n19361) );
  AND U19886 ( .A(n19362), .B(n19361), .Z(n19544) );
  NANDN U19887 ( .A(n38247), .B(n19363), .Z(n19365) );
  XOR U19888 ( .A(b[61]), .B(a[37]), .Z(n19632) );
  NANDN U19889 ( .A(n38248), .B(n19632), .Z(n19364) );
  AND U19890 ( .A(n19365), .B(n19364), .Z(n19543) );
  AND U19891 ( .A(b[63]), .B(a[33]), .Z(n19542) );
  XOR U19892 ( .A(n19543), .B(n19542), .Z(n19545) );
  XNOR U19893 ( .A(n19544), .B(n19545), .Z(n19503) );
  XNOR U19894 ( .A(n19504), .B(n19503), .Z(n19505) );
  NANDN U19895 ( .A(n19367), .B(n19366), .Z(n19371) );
  OR U19896 ( .A(n19369), .B(n19368), .Z(n19370) );
  NAND U19897 ( .A(n19371), .B(n19370), .Z(n19506) );
  XNOR U19898 ( .A(n19505), .B(n19506), .Z(n19665) );
  NANDN U19899 ( .A(n34223), .B(n19372), .Z(n19374) );
  XOR U19900 ( .A(b[27]), .B(a[71]), .Z(n19641) );
  NANDN U19901 ( .A(n34458), .B(n19641), .Z(n19373) );
  AND U19902 ( .A(n19374), .B(n19373), .Z(n19487) );
  NANDN U19903 ( .A(n34634), .B(n19375), .Z(n19377) );
  XOR U19904 ( .A(b[29]), .B(a[69]), .Z(n19644) );
  NANDN U19905 ( .A(n34722), .B(n19644), .Z(n19376) );
  AND U19906 ( .A(n19377), .B(n19376), .Z(n19486) );
  NANDN U19907 ( .A(n31055), .B(n19378), .Z(n19380) );
  XOR U19908 ( .A(a[85]), .B(b[13]), .Z(n19647) );
  NANDN U19909 ( .A(n31293), .B(n19647), .Z(n19379) );
  NAND U19910 ( .A(n19380), .B(n19379), .Z(n19485) );
  XOR U19911 ( .A(n19486), .B(n19485), .Z(n19488) );
  XOR U19912 ( .A(n19487), .B(n19488), .Z(n19561) );
  NANDN U19913 ( .A(n28889), .B(n19381), .Z(n19383) );
  XOR U19914 ( .A(a[93]), .B(b[5]), .Z(n19650) );
  NANDN U19915 ( .A(n29138), .B(n19650), .Z(n19382) );
  AND U19916 ( .A(n19383), .B(n19382), .Z(n19580) );
  NANDN U19917 ( .A(n209), .B(n19384), .Z(n19386) );
  XOR U19918 ( .A(a[95]), .B(b[3]), .Z(n19653) );
  NANDN U19919 ( .A(n28941), .B(n19653), .Z(n19385) );
  AND U19920 ( .A(n19386), .B(n19385), .Z(n19579) );
  NANDN U19921 ( .A(n35936), .B(n19387), .Z(n19389) );
  XOR U19922 ( .A(b[37]), .B(a[61]), .Z(n19656) );
  NANDN U19923 ( .A(n36047), .B(n19656), .Z(n19388) );
  NAND U19924 ( .A(n19389), .B(n19388), .Z(n19578) );
  XOR U19925 ( .A(n19579), .B(n19578), .Z(n19581) );
  XNOR U19926 ( .A(n19580), .B(n19581), .Z(n19560) );
  XNOR U19927 ( .A(n19561), .B(n19560), .Z(n19562) );
  NANDN U19928 ( .A(n19391), .B(n19390), .Z(n19395) );
  OR U19929 ( .A(n19393), .B(n19392), .Z(n19394) );
  NAND U19930 ( .A(n19395), .B(n19394), .Z(n19563) );
  XOR U19931 ( .A(n19562), .B(n19563), .Z(n19666) );
  XNOR U19932 ( .A(n19665), .B(n19666), .Z(n19667) );
  XNOR U19933 ( .A(n19668), .B(n19667), .Z(n19451) );
  XOR U19934 ( .A(n19452), .B(n19451), .Z(n19444) );
  NANDN U19935 ( .A(n19397), .B(n19396), .Z(n19401) );
  NANDN U19936 ( .A(n19399), .B(n19398), .Z(n19400) );
  AND U19937 ( .A(n19401), .B(n19400), .Z(n19443) );
  XNOR U19938 ( .A(n19444), .B(n19443), .Z(n19445) );
  XOR U19939 ( .A(n19446), .B(n19445), .Z(n19672) );
  XNOR U19940 ( .A(n19671), .B(n19672), .Z(n19673) );
  XOR U19941 ( .A(n19674), .B(n19673), .Z(n19686) );
  XOR U19942 ( .A(n19685), .B(n19686), .Z(n19692) );
  XOR U19943 ( .A(n19691), .B(n19692), .Z(n19696) );
  XOR U19944 ( .A(n19695), .B(n19696), .Z(n19698) );
  XOR U19945 ( .A(n19697), .B(n19698), .Z(n19414) );
  NANDN U19946 ( .A(n19403), .B(n19402), .Z(n19407) );
  NANDN U19947 ( .A(n19405), .B(n19404), .Z(n19406) );
  NAND U19948 ( .A(n19407), .B(n19406), .Z(n19413) );
  XNOR U19949 ( .A(n19414), .B(n19413), .Z(n19415) );
  XNOR U19950 ( .A(n19416), .B(n19415), .Z(n19701) );
  XNOR U19951 ( .A(sreg[161]), .B(n19701), .Z(n19703) );
  NANDN U19952 ( .A(sreg[160]), .B(n19408), .Z(n19412) );
  NAND U19953 ( .A(n19410), .B(n19409), .Z(n19411) );
  NAND U19954 ( .A(n19412), .B(n19411), .Z(n19702) );
  XNOR U19955 ( .A(n19703), .B(n19702), .Z(c[161]) );
  NANDN U19956 ( .A(n19414), .B(n19413), .Z(n19418) );
  NANDN U19957 ( .A(n19416), .B(n19415), .Z(n19417) );
  AND U19958 ( .A(n19418), .B(n19417), .Z(n19709) );
  NANDN U19959 ( .A(n19420), .B(n19419), .Z(n19424) );
  OR U19960 ( .A(n19422), .B(n19421), .Z(n19423) );
  AND U19961 ( .A(n19424), .B(n19423), .Z(n19978) );
  NANDN U19962 ( .A(n19426), .B(n19425), .Z(n19430) );
  NAND U19963 ( .A(n19428), .B(n19427), .Z(n19429) );
  AND U19964 ( .A(n19430), .B(n19429), .Z(n19977) );
  NANDN U19965 ( .A(n19432), .B(n19431), .Z(n19436) );
  NANDN U19966 ( .A(n19434), .B(n19433), .Z(n19435) );
  AND U19967 ( .A(n19436), .B(n19435), .Z(n19976) );
  XOR U19968 ( .A(n19977), .B(n19976), .Z(n19979) );
  XOR U19969 ( .A(n19978), .B(n19979), .Z(n19983) );
  NANDN U19970 ( .A(n19438), .B(n19437), .Z(n19442) );
  NANDN U19971 ( .A(n19440), .B(n19439), .Z(n19441) );
  NAND U19972 ( .A(n19442), .B(n19441), .Z(n19982) );
  XNOR U19973 ( .A(n19983), .B(n19982), .Z(n19984) );
  NANDN U19974 ( .A(n19444), .B(n19443), .Z(n19448) );
  NANDN U19975 ( .A(n19446), .B(n19445), .Z(n19447) );
  AND U19976 ( .A(n19448), .B(n19447), .Z(n19973) );
  NANDN U19977 ( .A(n19450), .B(n19449), .Z(n19454) );
  NAND U19978 ( .A(n19452), .B(n19451), .Z(n19453) );
  AND U19979 ( .A(n19454), .B(n19453), .Z(n19948) );
  NANDN U19980 ( .A(n19456), .B(n19455), .Z(n19460) );
  NANDN U19981 ( .A(n19458), .B(n19457), .Z(n19459) );
  AND U19982 ( .A(n19460), .B(n19459), .Z(n19966) );
  NANDN U19983 ( .A(n19462), .B(n19461), .Z(n19466) );
  NANDN U19984 ( .A(n19464), .B(n19463), .Z(n19465) );
  AND U19985 ( .A(n19466), .B(n19465), .Z(n19965) );
  NANDN U19986 ( .A(n33875), .B(n19467), .Z(n19469) );
  XOR U19987 ( .A(b[25]), .B(a[74]), .Z(n19742) );
  NANDN U19988 ( .A(n33994), .B(n19742), .Z(n19468) );
  AND U19989 ( .A(n19469), .B(n19468), .Z(n19876) );
  NANDN U19990 ( .A(n32013), .B(n19470), .Z(n19472) );
  XOR U19991 ( .A(a[82]), .B(b[17]), .Z(n19745) );
  NANDN U19992 ( .A(n32292), .B(n19745), .Z(n19471) );
  AND U19993 ( .A(n19472), .B(n19471), .Z(n19875) );
  NANDN U19994 ( .A(n31536), .B(n19473), .Z(n19475) );
  XOR U19995 ( .A(a[84]), .B(b[15]), .Z(n19748) );
  NANDN U19996 ( .A(n31925), .B(n19748), .Z(n19474) );
  NAND U19997 ( .A(n19475), .B(n19474), .Z(n19874) );
  XOR U19998 ( .A(n19875), .B(n19874), .Z(n19877) );
  XOR U19999 ( .A(n19876), .B(n19877), .Z(n19905) );
  NANDN U20000 ( .A(n37526), .B(n19476), .Z(n19478) );
  XOR U20001 ( .A(b[51]), .B(a[48]), .Z(n19751) );
  NANDN U20002 ( .A(n37605), .B(n19751), .Z(n19477) );
  AND U20003 ( .A(n19478), .B(n19477), .Z(n19900) );
  NANDN U20004 ( .A(n37705), .B(n19479), .Z(n19481) );
  XOR U20005 ( .A(b[53]), .B(a[46]), .Z(n19754) );
  NANDN U20006 ( .A(n37778), .B(n19754), .Z(n19480) );
  AND U20007 ( .A(n19481), .B(n19480), .Z(n19899) );
  NANDN U20008 ( .A(n36210), .B(n19482), .Z(n19484) );
  XOR U20009 ( .A(b[39]), .B(a[60]), .Z(n19757) );
  NANDN U20010 ( .A(n36347), .B(n19757), .Z(n19483) );
  NAND U20011 ( .A(n19484), .B(n19483), .Z(n19898) );
  XOR U20012 ( .A(n19899), .B(n19898), .Z(n19901) );
  XNOR U20013 ( .A(n19900), .B(n19901), .Z(n19904) );
  XNOR U20014 ( .A(n19905), .B(n19904), .Z(n19907) );
  NANDN U20015 ( .A(n19486), .B(n19485), .Z(n19490) );
  OR U20016 ( .A(n19488), .B(n19487), .Z(n19489) );
  AND U20017 ( .A(n19490), .B(n19489), .Z(n19906) );
  XOR U20018 ( .A(n19907), .B(n19906), .Z(n19733) );
  NANDN U20019 ( .A(n19492), .B(n19491), .Z(n19496) );
  OR U20020 ( .A(n19494), .B(n19493), .Z(n19495) );
  AND U20021 ( .A(n19496), .B(n19495), .Z(n19731) );
  NANDN U20022 ( .A(n19498), .B(n19497), .Z(n19502) );
  NANDN U20023 ( .A(n19500), .B(n19499), .Z(n19501) );
  NAND U20024 ( .A(n19502), .B(n19501), .Z(n19730) );
  XNOR U20025 ( .A(n19731), .B(n19730), .Z(n19732) );
  XNOR U20026 ( .A(n19733), .B(n19732), .Z(n19964) );
  XOR U20027 ( .A(n19965), .B(n19964), .Z(n19967) );
  XOR U20028 ( .A(n19966), .B(n19967), .Z(n19947) );
  NANDN U20029 ( .A(n19504), .B(n19503), .Z(n19508) );
  NANDN U20030 ( .A(n19506), .B(n19505), .Z(n19507) );
  AND U20031 ( .A(n19508), .B(n19507), .Z(n19959) );
  NANDN U20032 ( .A(n211), .B(n19509), .Z(n19511) );
  XOR U20033 ( .A(b[47]), .B(a[52]), .Z(n19784) );
  NANDN U20034 ( .A(n37172), .B(n19784), .Z(n19510) );
  AND U20035 ( .A(n19511), .B(n19510), .Z(n19825) );
  NANDN U20036 ( .A(n210), .B(n19512), .Z(n19514) );
  XOR U20037 ( .A(a[90]), .B(b[9]), .Z(n19787) );
  NANDN U20038 ( .A(n30267), .B(n19787), .Z(n19513) );
  AND U20039 ( .A(n19514), .B(n19513), .Z(n19824) );
  NANDN U20040 ( .A(n212), .B(n19515), .Z(n19517) );
  XOR U20041 ( .A(b[49]), .B(a[50]), .Z(n19790) );
  NANDN U20042 ( .A(n37432), .B(n19790), .Z(n19516) );
  NAND U20043 ( .A(n19517), .B(n19516), .Z(n19823) );
  XOR U20044 ( .A(n19824), .B(n19823), .Z(n19826) );
  XOR U20045 ( .A(n19825), .B(n19826), .Z(n19854) );
  NANDN U20046 ( .A(n36742), .B(n19518), .Z(n19520) );
  XOR U20047 ( .A(b[43]), .B(a[56]), .Z(n19793) );
  NANDN U20048 ( .A(n36891), .B(n19793), .Z(n19519) );
  AND U20049 ( .A(n19520), .B(n19519), .Z(n19804) );
  NANDN U20050 ( .A(n36991), .B(n19521), .Z(n19523) );
  XOR U20051 ( .A(b[45]), .B(a[54]), .Z(n19796) );
  NANDN U20052 ( .A(n37083), .B(n19796), .Z(n19522) );
  AND U20053 ( .A(n19523), .B(n19522), .Z(n19803) );
  NANDN U20054 ( .A(n30482), .B(n19524), .Z(n19526) );
  XOR U20055 ( .A(a[88]), .B(b[11]), .Z(n19799) );
  NANDN U20056 ( .A(n30891), .B(n19799), .Z(n19525) );
  NAND U20057 ( .A(n19526), .B(n19525), .Z(n19802) );
  XOR U20058 ( .A(n19803), .B(n19802), .Z(n19805) );
  XNOR U20059 ( .A(n19804), .B(n19805), .Z(n19853) );
  XNOR U20060 ( .A(n19854), .B(n19853), .Z(n19855) );
  NANDN U20061 ( .A(n19528), .B(n19527), .Z(n19532) );
  OR U20062 ( .A(n19530), .B(n19529), .Z(n19531) );
  NAND U20063 ( .A(n19532), .B(n19531), .Z(n19856) );
  XNOR U20064 ( .A(n19855), .B(n19856), .Z(n19958) );
  XNOR U20065 ( .A(n19959), .B(n19958), .Z(n19960) );
  NANDN U20066 ( .A(n29499), .B(n19533), .Z(n19535) );
  XOR U20067 ( .A(a[92]), .B(b[7]), .Z(n19808) );
  NANDN U20068 ( .A(n29735), .B(n19808), .Z(n19534) );
  AND U20069 ( .A(n19535), .B(n19534), .Z(n19768) );
  NANDN U20070 ( .A(n37857), .B(n19536), .Z(n19538) );
  XOR U20071 ( .A(b[55]), .B(a[44]), .Z(n19811) );
  NANDN U20072 ( .A(n37911), .B(n19811), .Z(n19537) );
  AND U20073 ( .A(n19538), .B(n19537), .Z(n19767) );
  NANDN U20074 ( .A(n35611), .B(n19539), .Z(n19541) );
  XOR U20075 ( .A(b[35]), .B(a[64]), .Z(n19814) );
  NANDN U20076 ( .A(n35801), .B(n19814), .Z(n19540) );
  NAND U20077 ( .A(n19541), .B(n19540), .Z(n19766) );
  XOR U20078 ( .A(n19767), .B(n19766), .Z(n19769) );
  XOR U20079 ( .A(n19768), .B(n19769), .Z(n19830) );
  NANDN U20080 ( .A(n19543), .B(n19542), .Z(n19547) );
  OR U20081 ( .A(n19545), .B(n19544), .Z(n19546) );
  AND U20082 ( .A(n19547), .B(n19546), .Z(n19829) );
  XNOR U20083 ( .A(n19830), .B(n19829), .Z(n19831) );
  NANDN U20084 ( .A(n19549), .B(n19548), .Z(n19553) );
  OR U20085 ( .A(n19551), .B(n19550), .Z(n19552) );
  NAND U20086 ( .A(n19553), .B(n19552), .Z(n19832) );
  XOR U20087 ( .A(n19831), .B(n19832), .Z(n19961) );
  XNOR U20088 ( .A(n19960), .B(n19961), .Z(n19946) );
  XOR U20089 ( .A(n19947), .B(n19946), .Z(n19949) );
  XOR U20090 ( .A(n19948), .B(n19949), .Z(n19971) );
  NANDN U20091 ( .A(n19555), .B(n19554), .Z(n19559) );
  NANDN U20092 ( .A(n19557), .B(n19556), .Z(n19558) );
  AND U20093 ( .A(n19559), .B(n19558), .Z(n19954) );
  NANDN U20094 ( .A(n19561), .B(n19560), .Z(n19565) );
  NANDN U20095 ( .A(n19563), .B(n19562), .Z(n19564) );
  AND U20096 ( .A(n19565), .B(n19564), .Z(n19953) );
  NANDN U20097 ( .A(n19567), .B(n19566), .Z(n19571) );
  NAND U20098 ( .A(n19569), .B(n19568), .Z(n19570) );
  AND U20099 ( .A(n19571), .B(n19570), .Z(n19952) );
  XOR U20100 ( .A(n19953), .B(n19952), .Z(n19955) );
  XOR U20101 ( .A(n19954), .B(n19955), .Z(n19721) );
  NANDN U20102 ( .A(n19573), .B(n19572), .Z(n19577) );
  NANDN U20103 ( .A(n19575), .B(n19574), .Z(n19576) );
  AND U20104 ( .A(n19577), .B(n19576), .Z(n19842) );
  NANDN U20105 ( .A(n19579), .B(n19578), .Z(n19583) );
  OR U20106 ( .A(n19581), .B(n19580), .Z(n19582) );
  NAND U20107 ( .A(n19583), .B(n19582), .Z(n19841) );
  XNOR U20108 ( .A(n19842), .B(n19841), .Z(n19844) );
  NANDN U20109 ( .A(n19585), .B(n19584), .Z(n19589) );
  OR U20110 ( .A(n19587), .B(n19586), .Z(n19588) );
  AND U20111 ( .A(n19589), .B(n19588), .Z(n19739) );
  NAND U20112 ( .A(b[0]), .B(a[98]), .Z(n19590) );
  XNOR U20113 ( .A(b[1]), .B(n19590), .Z(n19592) );
  NANDN U20114 ( .A(b[0]), .B(a[97]), .Z(n19591) );
  NAND U20115 ( .A(n19592), .B(n19591), .Z(n19775) );
  NANDN U20116 ( .A(n38278), .B(n19593), .Z(n19595) );
  XOR U20117 ( .A(b[63]), .B(a[36]), .Z(n19928) );
  NANDN U20118 ( .A(n38279), .B(n19928), .Z(n19594) );
  AND U20119 ( .A(n19595), .B(n19594), .Z(n19773) );
  NANDN U20120 ( .A(n35260), .B(n19596), .Z(n19598) );
  XOR U20121 ( .A(b[33]), .B(a[66]), .Z(n19931) );
  NANDN U20122 ( .A(n35456), .B(n19931), .Z(n19597) );
  NAND U20123 ( .A(n19598), .B(n19597), .Z(n19772) );
  XNOR U20124 ( .A(n19773), .B(n19772), .Z(n19774) );
  XNOR U20125 ( .A(n19775), .B(n19774), .Z(n19736) );
  NANDN U20126 ( .A(n37974), .B(n19599), .Z(n19601) );
  XOR U20127 ( .A(b[57]), .B(a[42]), .Z(n19937) );
  NANDN U20128 ( .A(n38031), .B(n19937), .Z(n19600) );
  AND U20129 ( .A(n19601), .B(n19600), .Z(n19913) );
  NANDN U20130 ( .A(n38090), .B(n19602), .Z(n19604) );
  XOR U20131 ( .A(b[59]), .B(a[40]), .Z(n19940) );
  NANDN U20132 ( .A(n38130), .B(n19940), .Z(n19603) );
  AND U20133 ( .A(n19604), .B(n19603), .Z(n19911) );
  NANDN U20134 ( .A(n36480), .B(n19605), .Z(n19607) );
  XOR U20135 ( .A(b[41]), .B(a[58]), .Z(n19943) );
  NANDN U20136 ( .A(n36594), .B(n19943), .Z(n19606) );
  NAND U20137 ( .A(n19607), .B(n19606), .Z(n19910) );
  XNOR U20138 ( .A(n19911), .B(n19910), .Z(n19912) );
  XOR U20139 ( .A(n19913), .B(n19912), .Z(n19737) );
  XNOR U20140 ( .A(n19736), .B(n19737), .Z(n19738) );
  XNOR U20141 ( .A(n19739), .B(n19738), .Z(n19843) );
  XOR U20142 ( .A(n19844), .B(n19843), .Z(n19725) );
  NANDN U20143 ( .A(n19609), .B(n19608), .Z(n19613) );
  NAND U20144 ( .A(n19611), .B(n19610), .Z(n19612) );
  NAND U20145 ( .A(n19613), .B(n19612), .Z(n19724) );
  XNOR U20146 ( .A(n19725), .B(n19724), .Z(n19727) );
  NANDN U20147 ( .A(n19615), .B(n19614), .Z(n19619) );
  NANDN U20148 ( .A(n19617), .B(n19616), .Z(n19618) );
  AND U20149 ( .A(n19619), .B(n19618), .Z(n19850) );
  NANDN U20150 ( .A(n32996), .B(n19620), .Z(n19622) );
  XOR U20151 ( .A(b[21]), .B(a[78]), .Z(n19859) );
  NANDN U20152 ( .A(n33271), .B(n19859), .Z(n19621) );
  AND U20153 ( .A(n19622), .B(n19621), .Z(n19924) );
  NANDN U20154 ( .A(n33866), .B(n19623), .Z(n19625) );
  XOR U20155 ( .A(b[23]), .B(a[76]), .Z(n19862) );
  NANDN U20156 ( .A(n33644), .B(n19862), .Z(n19624) );
  AND U20157 ( .A(n19625), .B(n19624), .Z(n19923) );
  NANDN U20158 ( .A(n32483), .B(n19626), .Z(n19628) );
  XOR U20159 ( .A(b[19]), .B(a[80]), .Z(n19865) );
  NANDN U20160 ( .A(n32823), .B(n19865), .Z(n19627) );
  NAND U20161 ( .A(n19628), .B(n19627), .Z(n19922) );
  XOR U20162 ( .A(n19923), .B(n19922), .Z(n19925) );
  XOR U20163 ( .A(n19924), .B(n19925), .Z(n19779) );
  NANDN U20164 ( .A(n34909), .B(n19629), .Z(n19631) );
  XOR U20165 ( .A(b[31]), .B(a[68]), .Z(n19868) );
  NANDN U20166 ( .A(n35145), .B(n19868), .Z(n19630) );
  AND U20167 ( .A(n19631), .B(n19630), .Z(n19819) );
  NANDN U20168 ( .A(n38247), .B(n19632), .Z(n19634) );
  XOR U20169 ( .A(b[61]), .B(a[38]), .Z(n19871) );
  NANDN U20170 ( .A(n38248), .B(n19871), .Z(n19633) );
  AND U20171 ( .A(n19634), .B(n19633), .Z(n19818) );
  AND U20172 ( .A(b[63]), .B(a[34]), .Z(n19817) );
  XOR U20173 ( .A(n19818), .B(n19817), .Z(n19820) );
  XNOR U20174 ( .A(n19819), .B(n19820), .Z(n19778) );
  XNOR U20175 ( .A(n19779), .B(n19778), .Z(n19780) );
  NANDN U20176 ( .A(n19636), .B(n19635), .Z(n19640) );
  OR U20177 ( .A(n19638), .B(n19637), .Z(n19639) );
  NAND U20178 ( .A(n19640), .B(n19639), .Z(n19781) );
  XNOR U20179 ( .A(n19780), .B(n19781), .Z(n19847) );
  NANDN U20180 ( .A(n34223), .B(n19641), .Z(n19643) );
  XOR U20181 ( .A(b[27]), .B(a[72]), .Z(n19880) );
  NANDN U20182 ( .A(n34458), .B(n19880), .Z(n19642) );
  AND U20183 ( .A(n19643), .B(n19642), .Z(n19762) );
  NANDN U20184 ( .A(n34634), .B(n19644), .Z(n19646) );
  XOR U20185 ( .A(b[29]), .B(a[70]), .Z(n19883) );
  NANDN U20186 ( .A(n34722), .B(n19883), .Z(n19645) );
  AND U20187 ( .A(n19646), .B(n19645), .Z(n19761) );
  NANDN U20188 ( .A(n31055), .B(n19647), .Z(n19649) );
  XOR U20189 ( .A(a[86]), .B(b[13]), .Z(n19886) );
  NANDN U20190 ( .A(n31293), .B(n19886), .Z(n19648) );
  NAND U20191 ( .A(n19649), .B(n19648), .Z(n19760) );
  XOR U20192 ( .A(n19761), .B(n19760), .Z(n19763) );
  XOR U20193 ( .A(n19762), .B(n19763), .Z(n19836) );
  NANDN U20194 ( .A(n28889), .B(n19650), .Z(n19652) );
  XOR U20195 ( .A(a[94]), .B(b[5]), .Z(n19889) );
  NANDN U20196 ( .A(n29138), .B(n19889), .Z(n19651) );
  AND U20197 ( .A(n19652), .B(n19651), .Z(n19918) );
  NANDN U20198 ( .A(n209), .B(n19653), .Z(n19655) );
  XOR U20199 ( .A(a[96]), .B(b[3]), .Z(n19892) );
  NANDN U20200 ( .A(n28941), .B(n19892), .Z(n19654) );
  AND U20201 ( .A(n19655), .B(n19654), .Z(n19917) );
  NANDN U20202 ( .A(n35936), .B(n19656), .Z(n19658) );
  XOR U20203 ( .A(b[37]), .B(a[62]), .Z(n19895) );
  NANDN U20204 ( .A(n36047), .B(n19895), .Z(n19657) );
  NAND U20205 ( .A(n19658), .B(n19657), .Z(n19916) );
  XOR U20206 ( .A(n19917), .B(n19916), .Z(n19919) );
  XNOR U20207 ( .A(n19918), .B(n19919), .Z(n19835) );
  XNOR U20208 ( .A(n19836), .B(n19835), .Z(n19837) );
  NANDN U20209 ( .A(n19660), .B(n19659), .Z(n19664) );
  OR U20210 ( .A(n19662), .B(n19661), .Z(n19663) );
  NAND U20211 ( .A(n19664), .B(n19663), .Z(n19838) );
  XOR U20212 ( .A(n19837), .B(n19838), .Z(n19848) );
  XNOR U20213 ( .A(n19847), .B(n19848), .Z(n19849) );
  XNOR U20214 ( .A(n19850), .B(n19849), .Z(n19726) );
  XOR U20215 ( .A(n19727), .B(n19726), .Z(n19719) );
  NANDN U20216 ( .A(n19666), .B(n19665), .Z(n19670) );
  NANDN U20217 ( .A(n19668), .B(n19667), .Z(n19669) );
  AND U20218 ( .A(n19670), .B(n19669), .Z(n19718) );
  XNOR U20219 ( .A(n19719), .B(n19718), .Z(n19720) );
  XNOR U20220 ( .A(n19721), .B(n19720), .Z(n19970) );
  XNOR U20221 ( .A(n19971), .B(n19970), .Z(n19972) );
  XOR U20222 ( .A(n19973), .B(n19972), .Z(n19985) );
  XNOR U20223 ( .A(n19984), .B(n19985), .Z(n19991) );
  NANDN U20224 ( .A(n19672), .B(n19671), .Z(n19676) );
  NANDN U20225 ( .A(n19674), .B(n19673), .Z(n19675) );
  AND U20226 ( .A(n19676), .B(n19675), .Z(n19989) );
  NANDN U20227 ( .A(n19678), .B(n19677), .Z(n19682) );
  OR U20228 ( .A(n19680), .B(n19679), .Z(n19681) );
  AND U20229 ( .A(n19682), .B(n19681), .Z(n19988) );
  XNOR U20230 ( .A(n19989), .B(n19988), .Z(n19990) );
  XOR U20231 ( .A(n19991), .B(n19990), .Z(n19713) );
  NANDN U20232 ( .A(n19684), .B(n19683), .Z(n19688) );
  NANDN U20233 ( .A(n19686), .B(n19685), .Z(n19687) );
  AND U20234 ( .A(n19688), .B(n19687), .Z(n19712) );
  XNOR U20235 ( .A(n19713), .B(n19712), .Z(n19714) );
  NANDN U20236 ( .A(n19690), .B(n19689), .Z(n19694) );
  NANDN U20237 ( .A(n19692), .B(n19691), .Z(n19693) );
  NAND U20238 ( .A(n19694), .B(n19693), .Z(n19715) );
  XNOR U20239 ( .A(n19714), .B(n19715), .Z(n19706) );
  NANDN U20240 ( .A(n19696), .B(n19695), .Z(n19700) );
  OR U20241 ( .A(n19698), .B(n19697), .Z(n19699) );
  NAND U20242 ( .A(n19700), .B(n19699), .Z(n19707) );
  XNOR U20243 ( .A(n19706), .B(n19707), .Z(n19708) );
  XNOR U20244 ( .A(n19709), .B(n19708), .Z(n19994) );
  XNOR U20245 ( .A(sreg[162]), .B(n19994), .Z(n19996) );
  NANDN U20246 ( .A(sreg[161]), .B(n19701), .Z(n19705) );
  NAND U20247 ( .A(n19703), .B(n19702), .Z(n19704) );
  NAND U20248 ( .A(n19705), .B(n19704), .Z(n19995) );
  XNOR U20249 ( .A(n19996), .B(n19995), .Z(c[162]) );
  NANDN U20250 ( .A(n19707), .B(n19706), .Z(n19711) );
  NANDN U20251 ( .A(n19709), .B(n19708), .Z(n19710) );
  AND U20252 ( .A(n19711), .B(n19710), .Z(n20002) );
  NANDN U20253 ( .A(n19713), .B(n19712), .Z(n19717) );
  NANDN U20254 ( .A(n19715), .B(n19714), .Z(n19716) );
  AND U20255 ( .A(n19717), .B(n19716), .Z(n20000) );
  NANDN U20256 ( .A(n19719), .B(n19718), .Z(n19723) );
  NANDN U20257 ( .A(n19721), .B(n19720), .Z(n19722) );
  AND U20258 ( .A(n19723), .B(n19722), .Z(n20271) );
  NANDN U20259 ( .A(n19725), .B(n19724), .Z(n19729) );
  NAND U20260 ( .A(n19727), .B(n19726), .Z(n19728) );
  AND U20261 ( .A(n19729), .B(n19728), .Z(n20247) );
  NANDN U20262 ( .A(n19731), .B(n19730), .Z(n19735) );
  NANDN U20263 ( .A(n19733), .B(n19732), .Z(n19734) );
  AND U20264 ( .A(n19735), .B(n19734), .Z(n20265) );
  NANDN U20265 ( .A(n19737), .B(n19736), .Z(n19741) );
  NANDN U20266 ( .A(n19739), .B(n19738), .Z(n19740) );
  AND U20267 ( .A(n19741), .B(n19740), .Z(n20264) );
  NANDN U20268 ( .A(n33875), .B(n19742), .Z(n19744) );
  XOR U20269 ( .A(b[25]), .B(a[75]), .Z(n20092) );
  NANDN U20270 ( .A(n33994), .B(n20092), .Z(n19743) );
  AND U20271 ( .A(n19744), .B(n19743), .Z(n20196) );
  NANDN U20272 ( .A(n32013), .B(n19745), .Z(n19747) );
  XOR U20273 ( .A(a[83]), .B(b[17]), .Z(n20095) );
  NANDN U20274 ( .A(n32292), .B(n20095), .Z(n19746) );
  AND U20275 ( .A(n19747), .B(n19746), .Z(n20195) );
  NANDN U20276 ( .A(n31536), .B(n19748), .Z(n19750) );
  XOR U20277 ( .A(a[85]), .B(b[15]), .Z(n20098) );
  NANDN U20278 ( .A(n31925), .B(n20098), .Z(n19749) );
  NAND U20279 ( .A(n19750), .B(n19749), .Z(n20194) );
  XOR U20280 ( .A(n20195), .B(n20194), .Z(n20197) );
  XOR U20281 ( .A(n20196), .B(n20197), .Z(n20183) );
  NANDN U20282 ( .A(n37526), .B(n19751), .Z(n19753) );
  XOR U20283 ( .A(b[51]), .B(a[49]), .Z(n20101) );
  NANDN U20284 ( .A(n37605), .B(n20101), .Z(n19752) );
  AND U20285 ( .A(n19753), .B(n19752), .Z(n20217) );
  NANDN U20286 ( .A(n37705), .B(n19754), .Z(n19756) );
  XOR U20287 ( .A(b[53]), .B(a[47]), .Z(n20104) );
  NANDN U20288 ( .A(n37778), .B(n20104), .Z(n19755) );
  AND U20289 ( .A(n19756), .B(n19755), .Z(n20216) );
  NANDN U20290 ( .A(n36210), .B(n19757), .Z(n19759) );
  XOR U20291 ( .A(b[39]), .B(a[61]), .Z(n20107) );
  NANDN U20292 ( .A(n36347), .B(n20107), .Z(n19758) );
  NAND U20293 ( .A(n19759), .B(n19758), .Z(n20215) );
  XOR U20294 ( .A(n20216), .B(n20215), .Z(n20218) );
  XNOR U20295 ( .A(n20217), .B(n20218), .Z(n20182) );
  XNOR U20296 ( .A(n20183), .B(n20182), .Z(n20185) );
  NANDN U20297 ( .A(n19761), .B(n19760), .Z(n19765) );
  OR U20298 ( .A(n19763), .B(n19762), .Z(n19764) );
  AND U20299 ( .A(n19765), .B(n19764), .Z(n20184) );
  XOR U20300 ( .A(n20185), .B(n20184), .Z(n20083) );
  NANDN U20301 ( .A(n19767), .B(n19766), .Z(n19771) );
  OR U20302 ( .A(n19769), .B(n19768), .Z(n19770) );
  AND U20303 ( .A(n19771), .B(n19770), .Z(n20081) );
  NANDN U20304 ( .A(n19773), .B(n19772), .Z(n19777) );
  NANDN U20305 ( .A(n19775), .B(n19774), .Z(n19776) );
  NAND U20306 ( .A(n19777), .B(n19776), .Z(n20080) );
  XNOR U20307 ( .A(n20081), .B(n20080), .Z(n20082) );
  XNOR U20308 ( .A(n20083), .B(n20082), .Z(n20263) );
  XOR U20309 ( .A(n20264), .B(n20263), .Z(n20266) );
  XOR U20310 ( .A(n20265), .B(n20266), .Z(n20246) );
  NANDN U20311 ( .A(n19779), .B(n19778), .Z(n19783) );
  NANDN U20312 ( .A(n19781), .B(n19780), .Z(n19782) );
  AND U20313 ( .A(n19783), .B(n19782), .Z(n20258) );
  NAND U20314 ( .A(n37294), .B(n19784), .Z(n19786) );
  XNOR U20315 ( .A(b[47]), .B(a[53]), .Z(n20035) );
  NANDN U20316 ( .A(n20035), .B(n37341), .Z(n19785) );
  NAND U20317 ( .A(n19786), .B(n19785), .Z(n20076) );
  NAND U20318 ( .A(n30627), .B(n19787), .Z(n19789) );
  XNOR U20319 ( .A(a[91]), .B(b[9]), .Z(n20038) );
  NANDN U20320 ( .A(n20038), .B(n30628), .Z(n19788) );
  NAND U20321 ( .A(n19789), .B(n19788), .Z(n20075) );
  NAND U20322 ( .A(n37536), .B(n19790), .Z(n19792) );
  XNOR U20323 ( .A(b[49]), .B(a[51]), .Z(n20041) );
  NANDN U20324 ( .A(n20041), .B(n37537), .Z(n19791) );
  NAND U20325 ( .A(n19792), .B(n19791), .Z(n20074) );
  XNOR U20326 ( .A(n20075), .B(n20074), .Z(n20077) );
  NANDN U20327 ( .A(n36742), .B(n19793), .Z(n19795) );
  XOR U20328 ( .A(b[43]), .B(a[57]), .Z(n20044) );
  NANDN U20329 ( .A(n36891), .B(n20044), .Z(n19794) );
  AND U20330 ( .A(n19795), .B(n19794), .Z(n20055) );
  NANDN U20331 ( .A(n36991), .B(n19796), .Z(n19798) );
  XOR U20332 ( .A(b[45]), .B(a[55]), .Z(n20047) );
  NANDN U20333 ( .A(n37083), .B(n20047), .Z(n19797) );
  AND U20334 ( .A(n19798), .B(n19797), .Z(n20054) );
  NANDN U20335 ( .A(n30482), .B(n19799), .Z(n19801) );
  XOR U20336 ( .A(a[89]), .B(b[11]), .Z(n20050) );
  NANDN U20337 ( .A(n30891), .B(n20050), .Z(n19800) );
  NAND U20338 ( .A(n19801), .B(n19800), .Z(n20053) );
  XOR U20339 ( .A(n20054), .B(n20053), .Z(n20056) );
  XNOR U20340 ( .A(n20055), .B(n20056), .Z(n20188) );
  XOR U20341 ( .A(n20189), .B(n20188), .Z(n20190) );
  NANDN U20342 ( .A(n19803), .B(n19802), .Z(n19807) );
  OR U20343 ( .A(n19805), .B(n19804), .Z(n19806) );
  NAND U20344 ( .A(n19807), .B(n19806), .Z(n20191) );
  XNOR U20345 ( .A(n20190), .B(n20191), .Z(n20257) );
  XNOR U20346 ( .A(n20258), .B(n20257), .Z(n20259) );
  NANDN U20347 ( .A(n29499), .B(n19808), .Z(n19810) );
  XOR U20348 ( .A(a[93]), .B(b[7]), .Z(n20059) );
  NANDN U20349 ( .A(n29735), .B(n20059), .Z(n19809) );
  AND U20350 ( .A(n19810), .B(n19809), .Z(n20118) );
  NANDN U20351 ( .A(n37857), .B(n19811), .Z(n19813) );
  XOR U20352 ( .A(b[55]), .B(a[45]), .Z(n20062) );
  NANDN U20353 ( .A(n37911), .B(n20062), .Z(n19812) );
  AND U20354 ( .A(n19813), .B(n19812), .Z(n20117) );
  NANDN U20355 ( .A(n35611), .B(n19814), .Z(n19816) );
  XOR U20356 ( .A(b[35]), .B(a[65]), .Z(n20065) );
  NANDN U20357 ( .A(n35801), .B(n20065), .Z(n19815) );
  NAND U20358 ( .A(n19816), .B(n19815), .Z(n20116) );
  XOR U20359 ( .A(n20117), .B(n20116), .Z(n20119) );
  XOR U20360 ( .A(n20118), .B(n20119), .Z(n20129) );
  NANDN U20361 ( .A(n19818), .B(n19817), .Z(n19822) );
  OR U20362 ( .A(n19820), .B(n19819), .Z(n19821) );
  AND U20363 ( .A(n19822), .B(n19821), .Z(n20128) );
  XNOR U20364 ( .A(n20129), .B(n20128), .Z(n20130) );
  NANDN U20365 ( .A(n19824), .B(n19823), .Z(n19828) );
  OR U20366 ( .A(n19826), .B(n19825), .Z(n19827) );
  NAND U20367 ( .A(n19828), .B(n19827), .Z(n20131) );
  XOR U20368 ( .A(n20130), .B(n20131), .Z(n20260) );
  XNOR U20369 ( .A(n20259), .B(n20260), .Z(n20245) );
  XOR U20370 ( .A(n20246), .B(n20245), .Z(n20248) );
  XOR U20371 ( .A(n20247), .B(n20248), .Z(n20270) );
  NANDN U20372 ( .A(n19830), .B(n19829), .Z(n19834) );
  NANDN U20373 ( .A(n19832), .B(n19831), .Z(n19833) );
  AND U20374 ( .A(n19834), .B(n19833), .Z(n20253) );
  NANDN U20375 ( .A(n19836), .B(n19835), .Z(n19840) );
  NANDN U20376 ( .A(n19838), .B(n19837), .Z(n19839) );
  AND U20377 ( .A(n19840), .B(n19839), .Z(n20252) );
  NANDN U20378 ( .A(n19842), .B(n19841), .Z(n19846) );
  NAND U20379 ( .A(n19844), .B(n19843), .Z(n19845) );
  AND U20380 ( .A(n19846), .B(n19845), .Z(n20251) );
  XOR U20381 ( .A(n20252), .B(n20251), .Z(n20254) );
  XOR U20382 ( .A(n20253), .B(n20254), .Z(n20020) );
  NANDN U20383 ( .A(n19848), .B(n19847), .Z(n19852) );
  NANDN U20384 ( .A(n19850), .B(n19849), .Z(n19851) );
  AND U20385 ( .A(n19852), .B(n19851), .Z(n20017) );
  NANDN U20386 ( .A(n19854), .B(n19853), .Z(n19858) );
  NANDN U20387 ( .A(n19856), .B(n19855), .Z(n19857) );
  AND U20388 ( .A(n19858), .B(n19857), .Z(n20241) );
  NANDN U20389 ( .A(n32996), .B(n19859), .Z(n19861) );
  XOR U20390 ( .A(b[21]), .B(a[79]), .Z(n20200) );
  NANDN U20391 ( .A(n33271), .B(n20200), .Z(n19860) );
  AND U20392 ( .A(n19861), .B(n19860), .Z(n20160) );
  NANDN U20393 ( .A(n33866), .B(n19862), .Z(n19864) );
  XOR U20394 ( .A(b[23]), .B(a[77]), .Z(n20203) );
  NANDN U20395 ( .A(n33644), .B(n20203), .Z(n19863) );
  AND U20396 ( .A(n19864), .B(n19863), .Z(n20159) );
  NANDN U20397 ( .A(n32483), .B(n19865), .Z(n19867) );
  XOR U20398 ( .A(b[19]), .B(a[81]), .Z(n20206) );
  NANDN U20399 ( .A(n32823), .B(n20206), .Z(n19866) );
  NAND U20400 ( .A(n19867), .B(n19866), .Z(n20158) );
  XOR U20401 ( .A(n20159), .B(n20158), .Z(n20161) );
  XOR U20402 ( .A(n20160), .B(n20161), .Z(n20030) );
  NANDN U20403 ( .A(n34909), .B(n19868), .Z(n19870) );
  XOR U20404 ( .A(b[31]), .B(a[69]), .Z(n20209) );
  NANDN U20405 ( .A(n35145), .B(n20209), .Z(n19869) );
  AND U20406 ( .A(n19870), .B(n19869), .Z(n20070) );
  NANDN U20407 ( .A(n38247), .B(n19871), .Z(n19873) );
  XOR U20408 ( .A(b[61]), .B(a[39]), .Z(n20212) );
  NANDN U20409 ( .A(n38248), .B(n20212), .Z(n19872) );
  AND U20410 ( .A(n19873), .B(n19872), .Z(n20069) );
  AND U20411 ( .A(b[63]), .B(a[35]), .Z(n20068) );
  XOR U20412 ( .A(n20069), .B(n20068), .Z(n20071) );
  XNOR U20413 ( .A(n20070), .B(n20071), .Z(n20029) );
  XNOR U20414 ( .A(n20030), .B(n20029), .Z(n20031) );
  NANDN U20415 ( .A(n19875), .B(n19874), .Z(n19879) );
  OR U20416 ( .A(n19877), .B(n19876), .Z(n19878) );
  NAND U20417 ( .A(n19879), .B(n19878), .Z(n20032) );
  XNOR U20418 ( .A(n20031), .B(n20032), .Z(n20239) );
  NANDN U20419 ( .A(n34223), .B(n19880), .Z(n19882) );
  XOR U20420 ( .A(b[27]), .B(a[73]), .Z(n20221) );
  NANDN U20421 ( .A(n34458), .B(n20221), .Z(n19881) );
  AND U20422 ( .A(n19882), .B(n19881), .Z(n20112) );
  NANDN U20423 ( .A(n34634), .B(n19883), .Z(n19885) );
  XOR U20424 ( .A(b[29]), .B(a[71]), .Z(n20224) );
  NANDN U20425 ( .A(n34722), .B(n20224), .Z(n19884) );
  AND U20426 ( .A(n19885), .B(n19884), .Z(n20111) );
  NANDN U20427 ( .A(n31055), .B(n19886), .Z(n19888) );
  XOR U20428 ( .A(a[87]), .B(b[13]), .Z(n20227) );
  NANDN U20429 ( .A(n31293), .B(n20227), .Z(n19887) );
  NAND U20430 ( .A(n19888), .B(n19887), .Z(n20110) );
  XOR U20431 ( .A(n20111), .B(n20110), .Z(n20113) );
  XOR U20432 ( .A(n20112), .B(n20113), .Z(n20135) );
  NANDN U20433 ( .A(n28889), .B(n19889), .Z(n19891) );
  XOR U20434 ( .A(a[95]), .B(b[5]), .Z(n20230) );
  NANDN U20435 ( .A(n29138), .B(n20230), .Z(n19890) );
  AND U20436 ( .A(n19891), .B(n19890), .Z(n20154) );
  NANDN U20437 ( .A(n209), .B(n19892), .Z(n19894) );
  XOR U20438 ( .A(a[97]), .B(b[3]), .Z(n20233) );
  NANDN U20439 ( .A(n28941), .B(n20233), .Z(n19893) );
  AND U20440 ( .A(n19894), .B(n19893), .Z(n20153) );
  NANDN U20441 ( .A(n35936), .B(n19895), .Z(n19897) );
  XOR U20442 ( .A(b[37]), .B(a[63]), .Z(n20236) );
  NANDN U20443 ( .A(n36047), .B(n20236), .Z(n19896) );
  NAND U20444 ( .A(n19897), .B(n19896), .Z(n20152) );
  XOR U20445 ( .A(n20153), .B(n20152), .Z(n20155) );
  XNOR U20446 ( .A(n20154), .B(n20155), .Z(n20134) );
  XNOR U20447 ( .A(n20135), .B(n20134), .Z(n20136) );
  NANDN U20448 ( .A(n19899), .B(n19898), .Z(n19903) );
  OR U20449 ( .A(n19901), .B(n19900), .Z(n19902) );
  NAND U20450 ( .A(n19903), .B(n19902), .Z(n20137) );
  XOR U20451 ( .A(n20136), .B(n20137), .Z(n20240) );
  XOR U20452 ( .A(n20239), .B(n20240), .Z(n20242) );
  XOR U20453 ( .A(n20241), .B(n20242), .Z(n20026) );
  NANDN U20454 ( .A(n19905), .B(n19904), .Z(n19909) );
  NAND U20455 ( .A(n19907), .B(n19906), .Z(n19908) );
  AND U20456 ( .A(n19909), .B(n19908), .Z(n20023) );
  NANDN U20457 ( .A(n19911), .B(n19910), .Z(n19915) );
  NANDN U20458 ( .A(n19913), .B(n19912), .Z(n19914) );
  AND U20459 ( .A(n19915), .B(n19914), .Z(n20141) );
  NANDN U20460 ( .A(n19917), .B(n19916), .Z(n19921) );
  OR U20461 ( .A(n19919), .B(n19918), .Z(n19920) );
  NAND U20462 ( .A(n19921), .B(n19920), .Z(n20140) );
  XNOR U20463 ( .A(n20141), .B(n20140), .Z(n20142) );
  NANDN U20464 ( .A(n19923), .B(n19922), .Z(n19927) );
  OR U20465 ( .A(n19925), .B(n19924), .Z(n19926) );
  AND U20466 ( .A(n19927), .B(n19926), .Z(n20089) );
  NANDN U20467 ( .A(n38278), .B(n19928), .Z(n19930) );
  XOR U20468 ( .A(b[63]), .B(a[37]), .Z(n20167) );
  NANDN U20469 ( .A(n38279), .B(n20167), .Z(n19929) );
  AND U20470 ( .A(n19930), .B(n19929), .Z(n20123) );
  NANDN U20471 ( .A(n35260), .B(n19931), .Z(n19933) );
  XOR U20472 ( .A(b[33]), .B(a[67]), .Z(n20170) );
  NANDN U20473 ( .A(n35456), .B(n20170), .Z(n19932) );
  NAND U20474 ( .A(n19933), .B(n19932), .Z(n20122) );
  XNOR U20475 ( .A(n20123), .B(n20122), .Z(n20124) );
  NAND U20476 ( .A(b[0]), .B(a[99]), .Z(n19934) );
  XNOR U20477 ( .A(b[1]), .B(n19934), .Z(n19936) );
  NANDN U20478 ( .A(b[0]), .B(a[98]), .Z(n19935) );
  NAND U20479 ( .A(n19936), .B(n19935), .Z(n20125) );
  XNOR U20480 ( .A(n20124), .B(n20125), .Z(n20086) );
  NANDN U20481 ( .A(n37974), .B(n19937), .Z(n19939) );
  XOR U20482 ( .A(b[57]), .B(a[43]), .Z(n20173) );
  NANDN U20483 ( .A(n38031), .B(n20173), .Z(n19938) );
  AND U20484 ( .A(n19939), .B(n19938), .Z(n20149) );
  NANDN U20485 ( .A(n38090), .B(n19940), .Z(n19942) );
  XOR U20486 ( .A(b[59]), .B(a[41]), .Z(n20176) );
  NANDN U20487 ( .A(n38130), .B(n20176), .Z(n19941) );
  AND U20488 ( .A(n19942), .B(n19941), .Z(n20147) );
  NANDN U20489 ( .A(n36480), .B(n19943), .Z(n19945) );
  XOR U20490 ( .A(b[41]), .B(a[59]), .Z(n20179) );
  NANDN U20491 ( .A(n36594), .B(n20179), .Z(n19944) );
  NAND U20492 ( .A(n19945), .B(n19944), .Z(n20146) );
  XNOR U20493 ( .A(n20147), .B(n20146), .Z(n20148) );
  XOR U20494 ( .A(n20149), .B(n20148), .Z(n20087) );
  XNOR U20495 ( .A(n20086), .B(n20087), .Z(n20088) );
  XOR U20496 ( .A(n20089), .B(n20088), .Z(n20143) );
  XOR U20497 ( .A(n20142), .B(n20143), .Z(n20024) );
  XNOR U20498 ( .A(n20023), .B(n20024), .Z(n20025) );
  XOR U20499 ( .A(n20026), .B(n20025), .Z(n20018) );
  XNOR U20500 ( .A(n20017), .B(n20018), .Z(n20019) );
  XNOR U20501 ( .A(n20020), .B(n20019), .Z(n20269) );
  XOR U20502 ( .A(n20270), .B(n20269), .Z(n20272) );
  XOR U20503 ( .A(n20271), .B(n20272), .Z(n20013) );
  NANDN U20504 ( .A(n19947), .B(n19946), .Z(n19951) );
  OR U20505 ( .A(n19949), .B(n19948), .Z(n19950) );
  AND U20506 ( .A(n19951), .B(n19950), .Z(n20012) );
  NANDN U20507 ( .A(n19953), .B(n19952), .Z(n19957) );
  OR U20508 ( .A(n19955), .B(n19954), .Z(n19956) );
  AND U20509 ( .A(n19957), .B(n19956), .Z(n20278) );
  NANDN U20510 ( .A(n19959), .B(n19958), .Z(n19963) );
  NANDN U20511 ( .A(n19961), .B(n19960), .Z(n19962) );
  AND U20512 ( .A(n19963), .B(n19962), .Z(n20276) );
  NANDN U20513 ( .A(n19965), .B(n19964), .Z(n19969) );
  OR U20514 ( .A(n19967), .B(n19966), .Z(n19968) );
  AND U20515 ( .A(n19969), .B(n19968), .Z(n20275) );
  XNOR U20516 ( .A(n20276), .B(n20275), .Z(n20277) );
  XNOR U20517 ( .A(n20278), .B(n20277), .Z(n20011) );
  XOR U20518 ( .A(n20012), .B(n20011), .Z(n20014) );
  XOR U20519 ( .A(n20013), .B(n20014), .Z(n20007) );
  NANDN U20520 ( .A(n19971), .B(n19970), .Z(n19975) );
  NANDN U20521 ( .A(n19973), .B(n19972), .Z(n19974) );
  AND U20522 ( .A(n19975), .B(n19974), .Z(n20006) );
  NANDN U20523 ( .A(n19977), .B(n19976), .Z(n19981) );
  OR U20524 ( .A(n19979), .B(n19978), .Z(n19980) );
  AND U20525 ( .A(n19981), .B(n19980), .Z(n20005) );
  XOR U20526 ( .A(n20006), .B(n20005), .Z(n20008) );
  XOR U20527 ( .A(n20007), .B(n20008), .Z(n20282) );
  NANDN U20528 ( .A(n19983), .B(n19982), .Z(n19987) );
  NANDN U20529 ( .A(n19985), .B(n19984), .Z(n19986) );
  AND U20530 ( .A(n19987), .B(n19986), .Z(n20281) );
  XNOR U20531 ( .A(n20282), .B(n20281), .Z(n20283) );
  NANDN U20532 ( .A(n19989), .B(n19988), .Z(n19993) );
  NAND U20533 ( .A(n19991), .B(n19990), .Z(n19992) );
  NAND U20534 ( .A(n19993), .B(n19992), .Z(n20284) );
  XNOR U20535 ( .A(n20283), .B(n20284), .Z(n19999) );
  XNOR U20536 ( .A(n20000), .B(n19999), .Z(n20001) );
  XNOR U20537 ( .A(n20002), .B(n20001), .Z(n20287) );
  XNOR U20538 ( .A(sreg[163]), .B(n20287), .Z(n20289) );
  NANDN U20539 ( .A(sreg[162]), .B(n19994), .Z(n19998) );
  NAND U20540 ( .A(n19996), .B(n19995), .Z(n19997) );
  NAND U20541 ( .A(n19998), .B(n19997), .Z(n20288) );
  XNOR U20542 ( .A(n20289), .B(n20288), .Z(c[163]) );
  NANDN U20543 ( .A(n20000), .B(n19999), .Z(n20004) );
  NANDN U20544 ( .A(n20002), .B(n20001), .Z(n20003) );
  AND U20545 ( .A(n20004), .B(n20003), .Z(n20295) );
  NANDN U20546 ( .A(n20006), .B(n20005), .Z(n20010) );
  OR U20547 ( .A(n20008), .B(n20007), .Z(n20009) );
  AND U20548 ( .A(n20010), .B(n20009), .Z(n20574) );
  NANDN U20549 ( .A(n20012), .B(n20011), .Z(n20016) );
  OR U20550 ( .A(n20014), .B(n20013), .Z(n20015) );
  AND U20551 ( .A(n20016), .B(n20015), .Z(n20572) );
  NANDN U20552 ( .A(n20018), .B(n20017), .Z(n20022) );
  NANDN U20553 ( .A(n20020), .B(n20019), .Z(n20021) );
  AND U20554 ( .A(n20022), .B(n20021), .Z(n20550) );
  NANDN U20555 ( .A(n20024), .B(n20023), .Z(n20028) );
  NANDN U20556 ( .A(n20026), .B(n20025), .Z(n20027) );
  AND U20557 ( .A(n20028), .B(n20027), .Z(n20301) );
  NANDN U20558 ( .A(n20030), .B(n20029), .Z(n20034) );
  NANDN U20559 ( .A(n20032), .B(n20031), .Z(n20033) );
  AND U20560 ( .A(n20034), .B(n20033), .Z(n20311) );
  NANDN U20561 ( .A(n20035), .B(n37294), .Z(n20037) );
  XNOR U20562 ( .A(b[47]), .B(a[54]), .Z(n20388) );
  NANDN U20563 ( .A(n20388), .B(n37341), .Z(n20036) );
  NAND U20564 ( .A(n20037), .B(n20036), .Z(n20429) );
  NANDN U20565 ( .A(n20038), .B(n30627), .Z(n20040) );
  XNOR U20566 ( .A(a[92]), .B(b[9]), .Z(n20391) );
  NANDN U20567 ( .A(n20391), .B(n30628), .Z(n20039) );
  NAND U20568 ( .A(n20040), .B(n20039), .Z(n20428) );
  NANDN U20569 ( .A(n20041), .B(n37536), .Z(n20043) );
  XNOR U20570 ( .A(b[49]), .B(a[52]), .Z(n20394) );
  NANDN U20571 ( .A(n20394), .B(n37537), .Z(n20042) );
  NAND U20572 ( .A(n20043), .B(n20042), .Z(n20427) );
  XNOR U20573 ( .A(n20428), .B(n20427), .Z(n20430) );
  NANDN U20574 ( .A(n36742), .B(n20044), .Z(n20046) );
  XOR U20575 ( .A(b[43]), .B(a[58]), .Z(n20397) );
  NANDN U20576 ( .A(n36891), .B(n20397), .Z(n20045) );
  AND U20577 ( .A(n20046), .B(n20045), .Z(n20408) );
  NANDN U20578 ( .A(n36991), .B(n20047), .Z(n20049) );
  XOR U20579 ( .A(b[45]), .B(a[56]), .Z(n20400) );
  NANDN U20580 ( .A(n37083), .B(n20400), .Z(n20048) );
  AND U20581 ( .A(n20049), .B(n20048), .Z(n20407) );
  NANDN U20582 ( .A(n30482), .B(n20050), .Z(n20052) );
  XOR U20583 ( .A(a[90]), .B(b[11]), .Z(n20403) );
  NANDN U20584 ( .A(n30891), .B(n20403), .Z(n20051) );
  NAND U20585 ( .A(n20052), .B(n20051), .Z(n20406) );
  XOR U20586 ( .A(n20407), .B(n20406), .Z(n20409) );
  XNOR U20587 ( .A(n20408), .B(n20409), .Z(n20493) );
  XOR U20588 ( .A(n20494), .B(n20493), .Z(n20495) );
  NANDN U20589 ( .A(n20054), .B(n20053), .Z(n20058) );
  OR U20590 ( .A(n20056), .B(n20055), .Z(n20057) );
  NAND U20591 ( .A(n20058), .B(n20057), .Z(n20496) );
  XNOR U20592 ( .A(n20495), .B(n20496), .Z(n20310) );
  XNOR U20593 ( .A(n20311), .B(n20310), .Z(n20313) );
  NANDN U20594 ( .A(n29499), .B(n20059), .Z(n20061) );
  XOR U20595 ( .A(a[94]), .B(b[7]), .Z(n20412) );
  NANDN U20596 ( .A(n29735), .B(n20412), .Z(n20060) );
  AND U20597 ( .A(n20061), .B(n20060), .Z(n20372) );
  NANDN U20598 ( .A(n37857), .B(n20062), .Z(n20064) );
  XOR U20599 ( .A(b[55]), .B(a[46]), .Z(n20415) );
  NANDN U20600 ( .A(n37911), .B(n20415), .Z(n20063) );
  AND U20601 ( .A(n20064), .B(n20063), .Z(n20371) );
  NANDN U20602 ( .A(n35611), .B(n20065), .Z(n20067) );
  XOR U20603 ( .A(b[35]), .B(a[66]), .Z(n20418) );
  NANDN U20604 ( .A(n35801), .B(n20418), .Z(n20066) );
  NAND U20605 ( .A(n20067), .B(n20066), .Z(n20370) );
  XOR U20606 ( .A(n20371), .B(n20370), .Z(n20373) );
  XOR U20607 ( .A(n20372), .B(n20373), .Z(n20446) );
  NANDN U20608 ( .A(n20069), .B(n20068), .Z(n20073) );
  OR U20609 ( .A(n20071), .B(n20070), .Z(n20072) );
  AND U20610 ( .A(n20073), .B(n20072), .Z(n20445) );
  XNOR U20611 ( .A(n20446), .B(n20445), .Z(n20447) );
  NAND U20612 ( .A(n20075), .B(n20074), .Z(n20079) );
  NANDN U20613 ( .A(n20077), .B(n20076), .Z(n20078) );
  NAND U20614 ( .A(n20079), .B(n20078), .Z(n20448) );
  XNOR U20615 ( .A(n20447), .B(n20448), .Z(n20312) );
  XOR U20616 ( .A(n20313), .B(n20312), .Z(n20299) );
  NANDN U20617 ( .A(n20081), .B(n20080), .Z(n20085) );
  NANDN U20618 ( .A(n20083), .B(n20082), .Z(n20084) );
  AND U20619 ( .A(n20085), .B(n20084), .Z(n20319) );
  NANDN U20620 ( .A(n20087), .B(n20086), .Z(n20091) );
  NANDN U20621 ( .A(n20089), .B(n20088), .Z(n20090) );
  AND U20622 ( .A(n20091), .B(n20090), .Z(n20317) );
  NANDN U20623 ( .A(n33875), .B(n20092), .Z(n20094) );
  XOR U20624 ( .A(b[25]), .B(a[76]), .Z(n20346) );
  NANDN U20625 ( .A(n33994), .B(n20346), .Z(n20093) );
  AND U20626 ( .A(n20094), .B(n20093), .Z(n20501) );
  NANDN U20627 ( .A(n32013), .B(n20095), .Z(n20097) );
  XOR U20628 ( .A(a[84]), .B(b[17]), .Z(n20349) );
  NANDN U20629 ( .A(n32292), .B(n20349), .Z(n20096) );
  AND U20630 ( .A(n20097), .B(n20096), .Z(n20500) );
  NANDN U20631 ( .A(n31536), .B(n20098), .Z(n20100) );
  XOR U20632 ( .A(a[86]), .B(b[15]), .Z(n20352) );
  NANDN U20633 ( .A(n31925), .B(n20352), .Z(n20099) );
  NAND U20634 ( .A(n20100), .B(n20099), .Z(n20499) );
  XOR U20635 ( .A(n20500), .B(n20499), .Z(n20502) );
  XOR U20636 ( .A(n20501), .B(n20502), .Z(n20488) );
  NANDN U20637 ( .A(n37526), .B(n20101), .Z(n20103) );
  XOR U20638 ( .A(b[51]), .B(a[50]), .Z(n20355) );
  NANDN U20639 ( .A(n37605), .B(n20355), .Z(n20102) );
  AND U20640 ( .A(n20103), .B(n20102), .Z(n20522) );
  NANDN U20641 ( .A(n37705), .B(n20104), .Z(n20106) );
  XOR U20642 ( .A(b[53]), .B(a[48]), .Z(n20358) );
  NANDN U20643 ( .A(n37778), .B(n20358), .Z(n20105) );
  AND U20644 ( .A(n20106), .B(n20105), .Z(n20521) );
  NANDN U20645 ( .A(n36210), .B(n20107), .Z(n20109) );
  XOR U20646 ( .A(b[39]), .B(a[62]), .Z(n20361) );
  NANDN U20647 ( .A(n36347), .B(n20361), .Z(n20108) );
  NAND U20648 ( .A(n20109), .B(n20108), .Z(n20520) );
  XOR U20649 ( .A(n20521), .B(n20520), .Z(n20523) );
  XNOR U20650 ( .A(n20522), .B(n20523), .Z(n20487) );
  XNOR U20651 ( .A(n20488), .B(n20487), .Z(n20490) );
  NANDN U20652 ( .A(n20111), .B(n20110), .Z(n20115) );
  OR U20653 ( .A(n20113), .B(n20112), .Z(n20114) );
  AND U20654 ( .A(n20115), .B(n20114), .Z(n20489) );
  XOR U20655 ( .A(n20490), .B(n20489), .Z(n20337) );
  NANDN U20656 ( .A(n20117), .B(n20116), .Z(n20121) );
  OR U20657 ( .A(n20119), .B(n20118), .Z(n20120) );
  AND U20658 ( .A(n20121), .B(n20120), .Z(n20335) );
  NANDN U20659 ( .A(n20123), .B(n20122), .Z(n20127) );
  NANDN U20660 ( .A(n20125), .B(n20124), .Z(n20126) );
  NAND U20661 ( .A(n20127), .B(n20126), .Z(n20334) );
  XNOR U20662 ( .A(n20335), .B(n20334), .Z(n20336) );
  XNOR U20663 ( .A(n20337), .B(n20336), .Z(n20316) );
  XNOR U20664 ( .A(n20317), .B(n20316), .Z(n20318) );
  XNOR U20665 ( .A(n20319), .B(n20318), .Z(n20298) );
  XNOR U20666 ( .A(n20299), .B(n20298), .Z(n20300) );
  XNOR U20667 ( .A(n20301), .B(n20300), .Z(n20548) );
  NANDN U20668 ( .A(n20129), .B(n20128), .Z(n20133) );
  NANDN U20669 ( .A(n20131), .B(n20130), .Z(n20132) );
  AND U20670 ( .A(n20133), .B(n20132), .Z(n20306) );
  NANDN U20671 ( .A(n20135), .B(n20134), .Z(n20139) );
  NANDN U20672 ( .A(n20137), .B(n20136), .Z(n20138) );
  AND U20673 ( .A(n20139), .B(n20138), .Z(n20305) );
  NANDN U20674 ( .A(n20141), .B(n20140), .Z(n20145) );
  NANDN U20675 ( .A(n20143), .B(n20142), .Z(n20144) );
  AND U20676 ( .A(n20145), .B(n20144), .Z(n20304) );
  XOR U20677 ( .A(n20305), .B(n20304), .Z(n20307) );
  XOR U20678 ( .A(n20306), .B(n20307), .Z(n20325) );
  NANDN U20679 ( .A(n20147), .B(n20146), .Z(n20151) );
  NANDN U20680 ( .A(n20149), .B(n20148), .Z(n20150) );
  AND U20681 ( .A(n20151), .B(n20150), .Z(n20440) );
  NANDN U20682 ( .A(n20153), .B(n20152), .Z(n20157) );
  OR U20683 ( .A(n20155), .B(n20154), .Z(n20156) );
  NAND U20684 ( .A(n20157), .B(n20156), .Z(n20439) );
  XNOR U20685 ( .A(n20440), .B(n20439), .Z(n20442) );
  NANDN U20686 ( .A(n20159), .B(n20158), .Z(n20163) );
  OR U20687 ( .A(n20161), .B(n20160), .Z(n20162) );
  NAND U20688 ( .A(n20163), .B(n20162), .Z(n20342) );
  NAND U20689 ( .A(b[0]), .B(a[100]), .Z(n20164) );
  XNOR U20690 ( .A(b[1]), .B(n20164), .Z(n20166) );
  NANDN U20691 ( .A(b[0]), .B(a[99]), .Z(n20165) );
  NAND U20692 ( .A(n20166), .B(n20165), .Z(n20379) );
  NANDN U20693 ( .A(n38278), .B(n20167), .Z(n20169) );
  XOR U20694 ( .A(b[63]), .B(a[38]), .Z(n20472) );
  NANDN U20695 ( .A(n38279), .B(n20472), .Z(n20168) );
  AND U20696 ( .A(n20169), .B(n20168), .Z(n20377) );
  NANDN U20697 ( .A(n35260), .B(n20170), .Z(n20172) );
  XOR U20698 ( .A(b[33]), .B(a[68]), .Z(n20475) );
  NANDN U20699 ( .A(n35456), .B(n20475), .Z(n20171) );
  NAND U20700 ( .A(n20172), .B(n20171), .Z(n20376) );
  XNOR U20701 ( .A(n20377), .B(n20376), .Z(n20378) );
  XNOR U20702 ( .A(n20379), .B(n20378), .Z(n20341) );
  NANDN U20703 ( .A(n37974), .B(n20173), .Z(n20175) );
  XOR U20704 ( .A(b[57]), .B(a[44]), .Z(n20478) );
  NANDN U20705 ( .A(n38031), .B(n20478), .Z(n20174) );
  AND U20706 ( .A(n20175), .B(n20174), .Z(n20453) );
  NANDN U20707 ( .A(n38090), .B(n20176), .Z(n20178) );
  XOR U20708 ( .A(b[59]), .B(a[42]), .Z(n20481) );
  NANDN U20709 ( .A(n38130), .B(n20481), .Z(n20177) );
  AND U20710 ( .A(n20178), .B(n20177), .Z(n20452) );
  NANDN U20711 ( .A(n36480), .B(n20179), .Z(n20181) );
  XOR U20712 ( .A(b[41]), .B(a[60]), .Z(n20484) );
  NANDN U20713 ( .A(n36594), .B(n20484), .Z(n20180) );
  NAND U20714 ( .A(n20181), .B(n20180), .Z(n20451) );
  XOR U20715 ( .A(n20452), .B(n20451), .Z(n20454) );
  XOR U20716 ( .A(n20453), .B(n20454), .Z(n20340) );
  XOR U20717 ( .A(n20341), .B(n20340), .Z(n20343) );
  XOR U20718 ( .A(n20342), .B(n20343), .Z(n20441) );
  XOR U20719 ( .A(n20442), .B(n20441), .Z(n20329) );
  NANDN U20720 ( .A(n20183), .B(n20182), .Z(n20187) );
  NAND U20721 ( .A(n20185), .B(n20184), .Z(n20186) );
  NAND U20722 ( .A(n20187), .B(n20186), .Z(n20328) );
  XNOR U20723 ( .A(n20329), .B(n20328), .Z(n20331) );
  NAND U20724 ( .A(n20189), .B(n20188), .Z(n20193) );
  NANDN U20725 ( .A(n20191), .B(n20190), .Z(n20192) );
  AND U20726 ( .A(n20193), .B(n20192), .Z(n20547) );
  NANDN U20727 ( .A(n20195), .B(n20194), .Z(n20199) );
  OR U20728 ( .A(n20197), .B(n20196), .Z(n20198) );
  AND U20729 ( .A(n20199), .B(n20198), .Z(n20384) );
  NANDN U20730 ( .A(n32996), .B(n20200), .Z(n20202) );
  XOR U20731 ( .A(b[21]), .B(a[80]), .Z(n20505) );
  NANDN U20732 ( .A(n33271), .B(n20505), .Z(n20201) );
  AND U20733 ( .A(n20202), .B(n20201), .Z(n20466) );
  NANDN U20734 ( .A(n33866), .B(n20203), .Z(n20205) );
  XOR U20735 ( .A(b[23]), .B(a[78]), .Z(n20508) );
  NANDN U20736 ( .A(n33644), .B(n20508), .Z(n20204) );
  AND U20737 ( .A(n20205), .B(n20204), .Z(n20464) );
  NANDN U20738 ( .A(n32483), .B(n20206), .Z(n20208) );
  XOR U20739 ( .A(b[19]), .B(a[82]), .Z(n20511) );
  NANDN U20740 ( .A(n32823), .B(n20511), .Z(n20207) );
  NAND U20741 ( .A(n20208), .B(n20207), .Z(n20463) );
  XNOR U20742 ( .A(n20464), .B(n20463), .Z(n20465) );
  XOR U20743 ( .A(n20466), .B(n20465), .Z(n20383) );
  NANDN U20744 ( .A(n34909), .B(n20209), .Z(n20211) );
  XOR U20745 ( .A(b[31]), .B(a[70]), .Z(n20514) );
  NANDN U20746 ( .A(n35145), .B(n20514), .Z(n20210) );
  AND U20747 ( .A(n20211), .B(n20210), .Z(n20424) );
  NANDN U20748 ( .A(n38247), .B(n20212), .Z(n20214) );
  XOR U20749 ( .A(b[61]), .B(a[40]), .Z(n20517) );
  NANDN U20750 ( .A(n38248), .B(n20517), .Z(n20213) );
  AND U20751 ( .A(n20214), .B(n20213), .Z(n20422) );
  AND U20752 ( .A(b[63]), .B(a[36]), .Z(n20421) );
  XNOR U20753 ( .A(n20422), .B(n20421), .Z(n20423) );
  XOR U20754 ( .A(n20424), .B(n20423), .Z(n20382) );
  XNOR U20755 ( .A(n20383), .B(n20382), .Z(n20385) );
  NANDN U20756 ( .A(n20216), .B(n20215), .Z(n20220) );
  OR U20757 ( .A(n20218), .B(n20217), .Z(n20219) );
  AND U20758 ( .A(n20220), .B(n20219), .Z(n20435) );
  NANDN U20759 ( .A(n34223), .B(n20221), .Z(n20223) );
  XOR U20760 ( .A(b[27]), .B(a[74]), .Z(n20526) );
  NANDN U20761 ( .A(n34458), .B(n20526), .Z(n20222) );
  AND U20762 ( .A(n20223), .B(n20222), .Z(n20367) );
  NANDN U20763 ( .A(n34634), .B(n20224), .Z(n20226) );
  XOR U20764 ( .A(b[29]), .B(a[72]), .Z(n20529) );
  NANDN U20765 ( .A(n34722), .B(n20529), .Z(n20225) );
  AND U20766 ( .A(n20226), .B(n20225), .Z(n20365) );
  NANDN U20767 ( .A(n31055), .B(n20227), .Z(n20229) );
  XOR U20768 ( .A(a[88]), .B(b[13]), .Z(n20532) );
  NANDN U20769 ( .A(n31293), .B(n20532), .Z(n20228) );
  NAND U20770 ( .A(n20229), .B(n20228), .Z(n20364) );
  XNOR U20771 ( .A(n20365), .B(n20364), .Z(n20366) );
  XOR U20772 ( .A(n20367), .B(n20366), .Z(n20434) );
  NANDN U20773 ( .A(n28889), .B(n20230), .Z(n20232) );
  XOR U20774 ( .A(a[96]), .B(b[5]), .Z(n20535) );
  NANDN U20775 ( .A(n29138), .B(n20535), .Z(n20231) );
  AND U20776 ( .A(n20232), .B(n20231), .Z(n20460) );
  NANDN U20777 ( .A(n209), .B(n20233), .Z(n20235) );
  XOR U20778 ( .A(a[98]), .B(b[3]), .Z(n20538) );
  NANDN U20779 ( .A(n28941), .B(n20538), .Z(n20234) );
  AND U20780 ( .A(n20235), .B(n20234), .Z(n20458) );
  NANDN U20781 ( .A(n35936), .B(n20236), .Z(n20238) );
  XOR U20782 ( .A(b[37]), .B(a[64]), .Z(n20541) );
  NANDN U20783 ( .A(n36047), .B(n20541), .Z(n20237) );
  NAND U20784 ( .A(n20238), .B(n20237), .Z(n20457) );
  XNOR U20785 ( .A(n20458), .B(n20457), .Z(n20459) );
  XOR U20786 ( .A(n20460), .B(n20459), .Z(n20433) );
  XNOR U20787 ( .A(n20434), .B(n20433), .Z(n20436) );
  XOR U20788 ( .A(n20545), .B(n20544), .Z(n20546) );
  XNOR U20789 ( .A(n20547), .B(n20546), .Z(n20330) );
  XOR U20790 ( .A(n20331), .B(n20330), .Z(n20323) );
  NANDN U20791 ( .A(n20240), .B(n20239), .Z(n20244) );
  OR U20792 ( .A(n20242), .B(n20241), .Z(n20243) );
  AND U20793 ( .A(n20244), .B(n20243), .Z(n20322) );
  XNOR U20794 ( .A(n20323), .B(n20322), .Z(n20324) );
  XOR U20795 ( .A(n20325), .B(n20324), .Z(n20549) );
  XOR U20796 ( .A(n20548), .B(n20549), .Z(n20551) );
  XOR U20797 ( .A(n20550), .B(n20551), .Z(n20562) );
  NANDN U20798 ( .A(n20246), .B(n20245), .Z(n20250) );
  OR U20799 ( .A(n20248), .B(n20247), .Z(n20249) );
  AND U20800 ( .A(n20250), .B(n20249), .Z(n20561) );
  NANDN U20801 ( .A(n20252), .B(n20251), .Z(n20256) );
  OR U20802 ( .A(n20254), .B(n20253), .Z(n20255) );
  AND U20803 ( .A(n20256), .B(n20255), .Z(n20557) );
  NANDN U20804 ( .A(n20258), .B(n20257), .Z(n20262) );
  NANDN U20805 ( .A(n20260), .B(n20259), .Z(n20261) );
  AND U20806 ( .A(n20262), .B(n20261), .Z(n20555) );
  NANDN U20807 ( .A(n20264), .B(n20263), .Z(n20268) );
  OR U20808 ( .A(n20266), .B(n20265), .Z(n20267) );
  AND U20809 ( .A(n20268), .B(n20267), .Z(n20554) );
  XNOR U20810 ( .A(n20555), .B(n20554), .Z(n20556) );
  XNOR U20811 ( .A(n20557), .B(n20556), .Z(n20560) );
  XOR U20812 ( .A(n20561), .B(n20560), .Z(n20563) );
  XOR U20813 ( .A(n20562), .B(n20563), .Z(n20569) );
  NANDN U20814 ( .A(n20270), .B(n20269), .Z(n20274) );
  OR U20815 ( .A(n20272), .B(n20271), .Z(n20273) );
  AND U20816 ( .A(n20274), .B(n20273), .Z(n20567) );
  NANDN U20817 ( .A(n20276), .B(n20275), .Z(n20280) );
  NANDN U20818 ( .A(n20278), .B(n20277), .Z(n20279) );
  AND U20819 ( .A(n20280), .B(n20279), .Z(n20566) );
  XNOR U20820 ( .A(n20567), .B(n20566), .Z(n20568) );
  XOR U20821 ( .A(n20569), .B(n20568), .Z(n20573) );
  XOR U20822 ( .A(n20572), .B(n20573), .Z(n20575) );
  XOR U20823 ( .A(n20574), .B(n20575), .Z(n20293) );
  NANDN U20824 ( .A(n20282), .B(n20281), .Z(n20286) );
  NANDN U20825 ( .A(n20284), .B(n20283), .Z(n20285) );
  NAND U20826 ( .A(n20286), .B(n20285), .Z(n20292) );
  XNOR U20827 ( .A(n20293), .B(n20292), .Z(n20294) );
  XNOR U20828 ( .A(n20295), .B(n20294), .Z(n20578) );
  XNOR U20829 ( .A(sreg[164]), .B(n20578), .Z(n20580) );
  NANDN U20830 ( .A(sreg[163]), .B(n20287), .Z(n20291) );
  NAND U20831 ( .A(n20289), .B(n20288), .Z(n20290) );
  NAND U20832 ( .A(n20291), .B(n20290), .Z(n20579) );
  XNOR U20833 ( .A(n20580), .B(n20579), .Z(c[164]) );
  NANDN U20834 ( .A(n20293), .B(n20292), .Z(n20297) );
  NANDN U20835 ( .A(n20295), .B(n20294), .Z(n20296) );
  AND U20836 ( .A(n20297), .B(n20296), .Z(n20586) );
  NANDN U20837 ( .A(n20299), .B(n20298), .Z(n20303) );
  NANDN U20838 ( .A(n20301), .B(n20300), .Z(n20302) );
  AND U20839 ( .A(n20303), .B(n20302), .Z(n20858) );
  NANDN U20840 ( .A(n20305), .B(n20304), .Z(n20309) );
  OR U20841 ( .A(n20307), .B(n20306), .Z(n20308) );
  AND U20842 ( .A(n20309), .B(n20308), .Z(n20603) );
  NANDN U20843 ( .A(n20311), .B(n20310), .Z(n20315) );
  NAND U20844 ( .A(n20313), .B(n20312), .Z(n20314) );
  AND U20845 ( .A(n20315), .B(n20314), .Z(n20602) );
  NANDN U20846 ( .A(n20317), .B(n20316), .Z(n20321) );
  NANDN U20847 ( .A(n20319), .B(n20318), .Z(n20320) );
  AND U20848 ( .A(n20321), .B(n20320), .Z(n20601) );
  XOR U20849 ( .A(n20602), .B(n20601), .Z(n20604) );
  XNOR U20850 ( .A(n20603), .B(n20604), .Z(n20857) );
  XNOR U20851 ( .A(n20858), .B(n20857), .Z(n20859) );
  NANDN U20852 ( .A(n20323), .B(n20322), .Z(n20327) );
  NANDN U20853 ( .A(n20325), .B(n20324), .Z(n20326) );
  AND U20854 ( .A(n20327), .B(n20326), .Z(n20598) );
  NANDN U20855 ( .A(n20329), .B(n20328), .Z(n20333) );
  NAND U20856 ( .A(n20331), .B(n20330), .Z(n20332) );
  AND U20857 ( .A(n20333), .B(n20332), .Z(n20609) );
  NANDN U20858 ( .A(n20335), .B(n20334), .Z(n20339) );
  NANDN U20859 ( .A(n20337), .B(n20336), .Z(n20338) );
  AND U20860 ( .A(n20339), .B(n20338), .Z(n20621) );
  NAND U20861 ( .A(n20341), .B(n20340), .Z(n20345) );
  NAND U20862 ( .A(n20343), .B(n20342), .Z(n20344) );
  AND U20863 ( .A(n20345), .B(n20344), .Z(n20620) );
  NANDN U20864 ( .A(n33875), .B(n20346), .Z(n20348) );
  XOR U20865 ( .A(b[25]), .B(a[77]), .Z(n20655) );
  NANDN U20866 ( .A(n33994), .B(n20655), .Z(n20347) );
  AND U20867 ( .A(n20348), .B(n20347), .Z(n20825) );
  NANDN U20868 ( .A(n32013), .B(n20349), .Z(n20351) );
  XOR U20869 ( .A(a[85]), .B(b[17]), .Z(n20658) );
  NANDN U20870 ( .A(n32292), .B(n20658), .Z(n20350) );
  AND U20871 ( .A(n20351), .B(n20350), .Z(n20824) );
  NANDN U20872 ( .A(n31536), .B(n20352), .Z(n20354) );
  XOR U20873 ( .A(a[87]), .B(b[15]), .Z(n20661) );
  NANDN U20874 ( .A(n31925), .B(n20661), .Z(n20353) );
  NAND U20875 ( .A(n20354), .B(n20353), .Z(n20823) );
  XOR U20876 ( .A(n20824), .B(n20823), .Z(n20826) );
  XOR U20877 ( .A(n20825), .B(n20826), .Z(n20797) );
  NANDN U20878 ( .A(n37526), .B(n20355), .Z(n20357) );
  XOR U20879 ( .A(b[51]), .B(a[51]), .Z(n20664) );
  NANDN U20880 ( .A(n37605), .B(n20664), .Z(n20356) );
  AND U20881 ( .A(n20357), .B(n20356), .Z(n20849) );
  NANDN U20882 ( .A(n37705), .B(n20358), .Z(n20360) );
  XOR U20883 ( .A(b[53]), .B(a[49]), .Z(n20667) );
  NANDN U20884 ( .A(n37778), .B(n20667), .Z(n20359) );
  AND U20885 ( .A(n20360), .B(n20359), .Z(n20848) );
  NANDN U20886 ( .A(n36210), .B(n20361), .Z(n20363) );
  XOR U20887 ( .A(b[39]), .B(a[63]), .Z(n20670) );
  NANDN U20888 ( .A(n36347), .B(n20670), .Z(n20362) );
  NAND U20889 ( .A(n20363), .B(n20362), .Z(n20847) );
  XOR U20890 ( .A(n20848), .B(n20847), .Z(n20850) );
  XNOR U20891 ( .A(n20849), .B(n20850), .Z(n20796) );
  XNOR U20892 ( .A(n20797), .B(n20796), .Z(n20799) );
  NANDN U20893 ( .A(n20365), .B(n20364), .Z(n20369) );
  NANDN U20894 ( .A(n20367), .B(n20366), .Z(n20368) );
  AND U20895 ( .A(n20369), .B(n20368), .Z(n20798) );
  XOR U20896 ( .A(n20799), .B(n20798), .Z(n20646) );
  NANDN U20897 ( .A(n20371), .B(n20370), .Z(n20375) );
  OR U20898 ( .A(n20373), .B(n20372), .Z(n20374) );
  AND U20899 ( .A(n20375), .B(n20374), .Z(n20644) );
  NANDN U20900 ( .A(n20377), .B(n20376), .Z(n20381) );
  NANDN U20901 ( .A(n20379), .B(n20378), .Z(n20380) );
  NAND U20902 ( .A(n20381), .B(n20380), .Z(n20643) );
  XNOR U20903 ( .A(n20644), .B(n20643), .Z(n20645) );
  XNOR U20904 ( .A(n20646), .B(n20645), .Z(n20619) );
  XOR U20905 ( .A(n20620), .B(n20619), .Z(n20622) );
  XOR U20906 ( .A(n20621), .B(n20622), .Z(n20608) );
  NAND U20907 ( .A(n20383), .B(n20382), .Z(n20387) );
  NANDN U20908 ( .A(n20385), .B(n20384), .Z(n20386) );
  AND U20909 ( .A(n20387), .B(n20386), .Z(n20626) );
  NANDN U20910 ( .A(n20388), .B(n37294), .Z(n20390) );
  XOR U20911 ( .A(b[47]), .B(a[55]), .Z(n20718) );
  NANDN U20912 ( .A(n37172), .B(n20718), .Z(n20389) );
  AND U20913 ( .A(n20390), .B(n20389), .Z(n20708) );
  NANDN U20914 ( .A(n20391), .B(n30627), .Z(n20393) );
  XOR U20915 ( .A(a[93]), .B(b[9]), .Z(n20721) );
  NANDN U20916 ( .A(n30267), .B(n20721), .Z(n20392) );
  AND U20917 ( .A(n20393), .B(n20392), .Z(n20707) );
  NANDN U20918 ( .A(n20394), .B(n37536), .Z(n20396) );
  XOR U20919 ( .A(b[49]), .B(a[53]), .Z(n20724) );
  NANDN U20920 ( .A(n37432), .B(n20724), .Z(n20395) );
  NAND U20921 ( .A(n20396), .B(n20395), .Z(n20706) );
  XOR U20922 ( .A(n20707), .B(n20706), .Z(n20709) );
  XOR U20923 ( .A(n20708), .B(n20709), .Z(n20803) );
  NANDN U20924 ( .A(n36742), .B(n20397), .Z(n20399) );
  XOR U20925 ( .A(b[43]), .B(a[59]), .Z(n20727) );
  NANDN U20926 ( .A(n36891), .B(n20727), .Z(n20398) );
  AND U20927 ( .A(n20399), .B(n20398), .Z(n20738) );
  NANDN U20928 ( .A(n36991), .B(n20400), .Z(n20402) );
  XOR U20929 ( .A(b[45]), .B(a[57]), .Z(n20730) );
  NANDN U20930 ( .A(n37083), .B(n20730), .Z(n20401) );
  AND U20931 ( .A(n20402), .B(n20401), .Z(n20737) );
  NANDN U20932 ( .A(n30482), .B(n20403), .Z(n20405) );
  XOR U20933 ( .A(a[91]), .B(b[11]), .Z(n20733) );
  NANDN U20934 ( .A(n30891), .B(n20733), .Z(n20404) );
  NAND U20935 ( .A(n20405), .B(n20404), .Z(n20736) );
  XOR U20936 ( .A(n20737), .B(n20736), .Z(n20739) );
  XNOR U20937 ( .A(n20738), .B(n20739), .Z(n20802) );
  XNOR U20938 ( .A(n20803), .B(n20802), .Z(n20804) );
  NANDN U20939 ( .A(n20407), .B(n20406), .Z(n20411) );
  OR U20940 ( .A(n20409), .B(n20408), .Z(n20410) );
  NAND U20941 ( .A(n20411), .B(n20410), .Z(n20805) );
  XNOR U20942 ( .A(n20804), .B(n20805), .Z(n20625) );
  XNOR U20943 ( .A(n20626), .B(n20625), .Z(n20627) );
  NANDN U20944 ( .A(n29499), .B(n20412), .Z(n20414) );
  XOR U20945 ( .A(a[95]), .B(b[7]), .Z(n20691) );
  NANDN U20946 ( .A(n29735), .B(n20691), .Z(n20413) );
  AND U20947 ( .A(n20414), .B(n20413), .Z(n20681) );
  NANDN U20948 ( .A(n37857), .B(n20415), .Z(n20417) );
  XOR U20949 ( .A(b[55]), .B(a[47]), .Z(n20694) );
  NANDN U20950 ( .A(n37911), .B(n20694), .Z(n20416) );
  AND U20951 ( .A(n20417), .B(n20416), .Z(n20680) );
  NANDN U20952 ( .A(n35611), .B(n20418), .Z(n20420) );
  XOR U20953 ( .A(b[35]), .B(a[67]), .Z(n20697) );
  NANDN U20954 ( .A(n35801), .B(n20697), .Z(n20419) );
  NAND U20955 ( .A(n20420), .B(n20419), .Z(n20679) );
  XOR U20956 ( .A(n20680), .B(n20679), .Z(n20682) );
  XOR U20957 ( .A(n20681), .B(n20682), .Z(n20755) );
  NANDN U20958 ( .A(n20422), .B(n20421), .Z(n20426) );
  NANDN U20959 ( .A(n20424), .B(n20423), .Z(n20425) );
  AND U20960 ( .A(n20426), .B(n20425), .Z(n20754) );
  XNOR U20961 ( .A(n20755), .B(n20754), .Z(n20756) );
  NAND U20962 ( .A(n20428), .B(n20427), .Z(n20432) );
  NANDN U20963 ( .A(n20430), .B(n20429), .Z(n20431) );
  NAND U20964 ( .A(n20432), .B(n20431), .Z(n20757) );
  XOR U20965 ( .A(n20756), .B(n20757), .Z(n20628) );
  XNOR U20966 ( .A(n20627), .B(n20628), .Z(n20607) );
  XOR U20967 ( .A(n20608), .B(n20607), .Z(n20610) );
  XOR U20968 ( .A(n20609), .B(n20610), .Z(n20596) );
  NAND U20969 ( .A(n20434), .B(n20433), .Z(n20438) );
  NANDN U20970 ( .A(n20436), .B(n20435), .Z(n20437) );
  NAND U20971 ( .A(n20438), .B(n20437), .Z(n20613) );
  NANDN U20972 ( .A(n20440), .B(n20439), .Z(n20444) );
  NAND U20973 ( .A(n20442), .B(n20441), .Z(n20443) );
  AND U20974 ( .A(n20444), .B(n20443), .Z(n20614) );
  XOR U20975 ( .A(n20613), .B(n20614), .Z(n20616) );
  NANDN U20976 ( .A(n20446), .B(n20445), .Z(n20450) );
  NANDN U20977 ( .A(n20448), .B(n20447), .Z(n20449) );
  NAND U20978 ( .A(n20450), .B(n20449), .Z(n20615) );
  XOR U20979 ( .A(n20616), .B(n20615), .Z(n20634) );
  NANDN U20980 ( .A(n20452), .B(n20451), .Z(n20456) );
  OR U20981 ( .A(n20454), .B(n20453), .Z(n20455) );
  AND U20982 ( .A(n20456), .B(n20455), .Z(n20749) );
  NANDN U20983 ( .A(n20458), .B(n20457), .Z(n20462) );
  NANDN U20984 ( .A(n20460), .B(n20459), .Z(n20461) );
  NAND U20985 ( .A(n20462), .B(n20461), .Z(n20748) );
  XNOR U20986 ( .A(n20749), .B(n20748), .Z(n20751) );
  NANDN U20987 ( .A(n20464), .B(n20463), .Z(n20468) );
  NANDN U20988 ( .A(n20466), .B(n20465), .Z(n20467) );
  NAND U20989 ( .A(n20468), .B(n20467), .Z(n20651) );
  NAND U20990 ( .A(b[0]), .B(a[101]), .Z(n20469) );
  XNOR U20991 ( .A(b[1]), .B(n20469), .Z(n20471) );
  NANDN U20992 ( .A(b[0]), .B(a[100]), .Z(n20470) );
  NAND U20993 ( .A(n20471), .B(n20470), .Z(n20688) );
  NANDN U20994 ( .A(n38278), .B(n20472), .Z(n20474) );
  XOR U20995 ( .A(b[63]), .B(a[39]), .Z(n20781) );
  NANDN U20996 ( .A(n38279), .B(n20781), .Z(n20473) );
  AND U20997 ( .A(n20474), .B(n20473), .Z(n20686) );
  NANDN U20998 ( .A(n35260), .B(n20475), .Z(n20477) );
  XOR U20999 ( .A(b[33]), .B(a[69]), .Z(n20784) );
  NANDN U21000 ( .A(n35456), .B(n20784), .Z(n20476) );
  NAND U21001 ( .A(n20477), .B(n20476), .Z(n20685) );
  XNOR U21002 ( .A(n20686), .B(n20685), .Z(n20687) );
  XNOR U21003 ( .A(n20688), .B(n20687), .Z(n20650) );
  NANDN U21004 ( .A(n37974), .B(n20478), .Z(n20480) );
  XOR U21005 ( .A(b[57]), .B(a[45]), .Z(n20787) );
  NANDN U21006 ( .A(n38031), .B(n20787), .Z(n20479) );
  AND U21007 ( .A(n20480), .B(n20479), .Z(n20762) );
  NANDN U21008 ( .A(n38090), .B(n20481), .Z(n20483) );
  XOR U21009 ( .A(b[59]), .B(a[43]), .Z(n20790) );
  NANDN U21010 ( .A(n38130), .B(n20790), .Z(n20482) );
  AND U21011 ( .A(n20483), .B(n20482), .Z(n20761) );
  NANDN U21012 ( .A(n36480), .B(n20484), .Z(n20486) );
  XOR U21013 ( .A(b[41]), .B(a[61]), .Z(n20793) );
  NANDN U21014 ( .A(n36594), .B(n20793), .Z(n20485) );
  NAND U21015 ( .A(n20486), .B(n20485), .Z(n20760) );
  XOR U21016 ( .A(n20761), .B(n20760), .Z(n20763) );
  XOR U21017 ( .A(n20762), .B(n20763), .Z(n20649) );
  XOR U21018 ( .A(n20650), .B(n20649), .Z(n20652) );
  XOR U21019 ( .A(n20651), .B(n20652), .Z(n20750) );
  XOR U21020 ( .A(n20751), .B(n20750), .Z(n20638) );
  NANDN U21021 ( .A(n20488), .B(n20487), .Z(n20492) );
  NAND U21022 ( .A(n20490), .B(n20489), .Z(n20491) );
  NAND U21023 ( .A(n20492), .B(n20491), .Z(n20637) );
  XNOR U21024 ( .A(n20638), .B(n20637), .Z(n20640) );
  NAND U21025 ( .A(n20494), .B(n20493), .Z(n20498) );
  NANDN U21026 ( .A(n20496), .B(n20495), .Z(n20497) );
  AND U21027 ( .A(n20498), .B(n20497), .Z(n20856) );
  NANDN U21028 ( .A(n20500), .B(n20499), .Z(n20504) );
  OR U21029 ( .A(n20502), .B(n20501), .Z(n20503) );
  AND U21030 ( .A(n20504), .B(n20503), .Z(n20714) );
  NANDN U21031 ( .A(n32996), .B(n20505), .Z(n20507) );
  XOR U21032 ( .A(b[21]), .B(a[81]), .Z(n20808) );
  NANDN U21033 ( .A(n33271), .B(n20808), .Z(n20506) );
  AND U21034 ( .A(n20507), .B(n20506), .Z(n20775) );
  NANDN U21035 ( .A(n33866), .B(n20508), .Z(n20510) );
  XOR U21036 ( .A(b[23]), .B(a[79]), .Z(n20811) );
  NANDN U21037 ( .A(n33644), .B(n20811), .Z(n20509) );
  AND U21038 ( .A(n20510), .B(n20509), .Z(n20773) );
  NANDN U21039 ( .A(n32483), .B(n20511), .Z(n20513) );
  XOR U21040 ( .A(b[19]), .B(a[83]), .Z(n20814) );
  NANDN U21041 ( .A(n32823), .B(n20814), .Z(n20512) );
  NAND U21042 ( .A(n20513), .B(n20512), .Z(n20772) );
  XNOR U21043 ( .A(n20773), .B(n20772), .Z(n20774) );
  XOR U21044 ( .A(n20775), .B(n20774), .Z(n20713) );
  NANDN U21045 ( .A(n34909), .B(n20514), .Z(n20516) );
  XOR U21046 ( .A(b[31]), .B(a[71]), .Z(n20817) );
  NANDN U21047 ( .A(n35145), .B(n20817), .Z(n20515) );
  AND U21048 ( .A(n20516), .B(n20515), .Z(n20703) );
  NANDN U21049 ( .A(n38247), .B(n20517), .Z(n20519) );
  XOR U21050 ( .A(b[61]), .B(a[41]), .Z(n20820) );
  NANDN U21051 ( .A(n38248), .B(n20820), .Z(n20518) );
  AND U21052 ( .A(n20519), .B(n20518), .Z(n20701) );
  AND U21053 ( .A(b[63]), .B(a[37]), .Z(n20700) );
  XNOR U21054 ( .A(n20701), .B(n20700), .Z(n20702) );
  XOR U21055 ( .A(n20703), .B(n20702), .Z(n20712) );
  XNOR U21056 ( .A(n20713), .B(n20712), .Z(n20715) );
  NANDN U21057 ( .A(n20521), .B(n20520), .Z(n20525) );
  OR U21058 ( .A(n20523), .B(n20522), .Z(n20524) );
  AND U21059 ( .A(n20525), .B(n20524), .Z(n20744) );
  NANDN U21060 ( .A(n34223), .B(n20526), .Z(n20528) );
  XOR U21061 ( .A(b[27]), .B(a[75]), .Z(n20829) );
  NANDN U21062 ( .A(n34458), .B(n20829), .Z(n20527) );
  AND U21063 ( .A(n20528), .B(n20527), .Z(n20676) );
  NANDN U21064 ( .A(n34634), .B(n20529), .Z(n20531) );
  XOR U21065 ( .A(b[29]), .B(a[73]), .Z(n20832) );
  NANDN U21066 ( .A(n34722), .B(n20832), .Z(n20530) );
  AND U21067 ( .A(n20531), .B(n20530), .Z(n20674) );
  NANDN U21068 ( .A(n31055), .B(n20532), .Z(n20534) );
  XOR U21069 ( .A(a[89]), .B(b[13]), .Z(n20835) );
  NANDN U21070 ( .A(n31293), .B(n20835), .Z(n20533) );
  NAND U21071 ( .A(n20534), .B(n20533), .Z(n20673) );
  XNOR U21072 ( .A(n20674), .B(n20673), .Z(n20675) );
  XOR U21073 ( .A(n20676), .B(n20675), .Z(n20743) );
  NANDN U21074 ( .A(n28889), .B(n20535), .Z(n20537) );
  XOR U21075 ( .A(a[97]), .B(b[5]), .Z(n20838) );
  NANDN U21076 ( .A(n29138), .B(n20838), .Z(n20536) );
  AND U21077 ( .A(n20537), .B(n20536), .Z(n20769) );
  NANDN U21078 ( .A(n209), .B(n20538), .Z(n20540) );
  XOR U21079 ( .A(a[99]), .B(b[3]), .Z(n20841) );
  NANDN U21080 ( .A(n28941), .B(n20841), .Z(n20539) );
  AND U21081 ( .A(n20540), .B(n20539), .Z(n20767) );
  NANDN U21082 ( .A(n35936), .B(n20541), .Z(n20543) );
  XOR U21083 ( .A(b[37]), .B(a[65]), .Z(n20844) );
  NANDN U21084 ( .A(n36047), .B(n20844), .Z(n20542) );
  NAND U21085 ( .A(n20543), .B(n20542), .Z(n20766) );
  XNOR U21086 ( .A(n20767), .B(n20766), .Z(n20768) );
  XOR U21087 ( .A(n20769), .B(n20768), .Z(n20742) );
  XNOR U21088 ( .A(n20743), .B(n20742), .Z(n20745) );
  XOR U21089 ( .A(n20854), .B(n20853), .Z(n20855) );
  XNOR U21090 ( .A(n20856), .B(n20855), .Z(n20639) );
  XOR U21091 ( .A(n20640), .B(n20639), .Z(n20632) );
  XNOR U21092 ( .A(n20632), .B(n20631), .Z(n20633) );
  XNOR U21093 ( .A(n20634), .B(n20633), .Z(n20595) );
  XNOR U21094 ( .A(n20596), .B(n20595), .Z(n20597) );
  XOR U21095 ( .A(n20598), .B(n20597), .Z(n20860) );
  XNOR U21096 ( .A(n20859), .B(n20860), .Z(n20866) );
  NANDN U21097 ( .A(n20549), .B(n20548), .Z(n20553) );
  OR U21098 ( .A(n20551), .B(n20550), .Z(n20552) );
  AND U21099 ( .A(n20553), .B(n20552), .Z(n20864) );
  NANDN U21100 ( .A(n20555), .B(n20554), .Z(n20559) );
  NANDN U21101 ( .A(n20557), .B(n20556), .Z(n20558) );
  AND U21102 ( .A(n20559), .B(n20558), .Z(n20863) );
  XNOR U21103 ( .A(n20864), .B(n20863), .Z(n20865) );
  XOR U21104 ( .A(n20866), .B(n20865), .Z(n20590) );
  NANDN U21105 ( .A(n20561), .B(n20560), .Z(n20565) );
  OR U21106 ( .A(n20563), .B(n20562), .Z(n20564) );
  NAND U21107 ( .A(n20565), .B(n20564), .Z(n20589) );
  XNOR U21108 ( .A(n20590), .B(n20589), .Z(n20591) );
  NANDN U21109 ( .A(n20567), .B(n20566), .Z(n20571) );
  NANDN U21110 ( .A(n20569), .B(n20568), .Z(n20570) );
  NAND U21111 ( .A(n20571), .B(n20570), .Z(n20592) );
  XNOR U21112 ( .A(n20591), .B(n20592), .Z(n20583) );
  NANDN U21113 ( .A(n20573), .B(n20572), .Z(n20577) );
  OR U21114 ( .A(n20575), .B(n20574), .Z(n20576) );
  NAND U21115 ( .A(n20577), .B(n20576), .Z(n20584) );
  XNOR U21116 ( .A(n20583), .B(n20584), .Z(n20585) );
  XNOR U21117 ( .A(n20586), .B(n20585), .Z(n20869) );
  XNOR U21118 ( .A(sreg[165]), .B(n20869), .Z(n20871) );
  NANDN U21119 ( .A(sreg[164]), .B(n20578), .Z(n20582) );
  NAND U21120 ( .A(n20580), .B(n20579), .Z(n20581) );
  NAND U21121 ( .A(n20582), .B(n20581), .Z(n20870) );
  XNOR U21122 ( .A(n20871), .B(n20870), .Z(c[165]) );
  NANDN U21123 ( .A(n20584), .B(n20583), .Z(n20588) );
  NANDN U21124 ( .A(n20586), .B(n20585), .Z(n20587) );
  AND U21125 ( .A(n20588), .B(n20587), .Z(n20877) );
  NANDN U21126 ( .A(n20590), .B(n20589), .Z(n20594) );
  NANDN U21127 ( .A(n20592), .B(n20591), .Z(n20593) );
  AND U21128 ( .A(n20594), .B(n20593), .Z(n20875) );
  NANDN U21129 ( .A(n20596), .B(n20595), .Z(n20600) );
  NANDN U21130 ( .A(n20598), .B(n20597), .Z(n20599) );
  AND U21131 ( .A(n20600), .B(n20599), .Z(n21157) );
  NANDN U21132 ( .A(n20602), .B(n20601), .Z(n20606) );
  OR U21133 ( .A(n20604), .B(n20603), .Z(n20605) );
  AND U21134 ( .A(n20606), .B(n20605), .Z(n21156) );
  XNOR U21135 ( .A(n21157), .B(n21156), .Z(n21159) );
  NANDN U21136 ( .A(n20608), .B(n20607), .Z(n20612) );
  OR U21137 ( .A(n20610), .B(n20609), .Z(n20611) );
  AND U21138 ( .A(n20612), .B(n20611), .Z(n21150) );
  NAND U21139 ( .A(n20614), .B(n20613), .Z(n20618) );
  NAND U21140 ( .A(n20616), .B(n20615), .Z(n20617) );
  AND U21141 ( .A(n20618), .B(n20617), .Z(n20894) );
  NANDN U21142 ( .A(n20620), .B(n20619), .Z(n20624) );
  OR U21143 ( .A(n20622), .B(n20621), .Z(n20623) );
  AND U21144 ( .A(n20624), .B(n20623), .Z(n20893) );
  NANDN U21145 ( .A(n20626), .B(n20625), .Z(n20630) );
  NANDN U21146 ( .A(n20628), .B(n20627), .Z(n20629) );
  AND U21147 ( .A(n20630), .B(n20629), .Z(n20892) );
  XOR U21148 ( .A(n20893), .B(n20892), .Z(n20895) );
  XOR U21149 ( .A(n20894), .B(n20895), .Z(n21151) );
  XNOR U21150 ( .A(n21150), .B(n21151), .Z(n21152) );
  NANDN U21151 ( .A(n20632), .B(n20631), .Z(n20636) );
  NANDN U21152 ( .A(n20634), .B(n20633), .Z(n20635) );
  AND U21153 ( .A(n20636), .B(n20635), .Z(n20889) );
  NANDN U21154 ( .A(n20638), .B(n20637), .Z(n20642) );
  NAND U21155 ( .A(n20640), .B(n20639), .Z(n20641) );
  AND U21156 ( .A(n20642), .B(n20641), .Z(n20900) );
  NANDN U21157 ( .A(n20644), .B(n20643), .Z(n20648) );
  NANDN U21158 ( .A(n20646), .B(n20645), .Z(n20647) );
  AND U21159 ( .A(n20648), .B(n20647), .Z(n20912) );
  NAND U21160 ( .A(n20650), .B(n20649), .Z(n20654) );
  NAND U21161 ( .A(n20652), .B(n20651), .Z(n20653) );
  AND U21162 ( .A(n20654), .B(n20653), .Z(n20911) );
  NANDN U21163 ( .A(n33875), .B(n20655), .Z(n20657) );
  XOR U21164 ( .A(b[25]), .B(a[78]), .Z(n20946) );
  NANDN U21165 ( .A(n33994), .B(n20946), .Z(n20656) );
  AND U21166 ( .A(n20657), .B(n20656), .Z(n21116) );
  NANDN U21167 ( .A(n32013), .B(n20658), .Z(n20660) );
  XOR U21168 ( .A(a[86]), .B(b[17]), .Z(n20949) );
  NANDN U21169 ( .A(n32292), .B(n20949), .Z(n20659) );
  AND U21170 ( .A(n20660), .B(n20659), .Z(n21115) );
  NANDN U21171 ( .A(n31536), .B(n20661), .Z(n20663) );
  XOR U21172 ( .A(a[88]), .B(b[15]), .Z(n20952) );
  NANDN U21173 ( .A(n31925), .B(n20952), .Z(n20662) );
  NAND U21174 ( .A(n20663), .B(n20662), .Z(n21114) );
  XOR U21175 ( .A(n21115), .B(n21114), .Z(n21117) );
  XOR U21176 ( .A(n21116), .B(n21117), .Z(n21088) );
  NANDN U21177 ( .A(n37526), .B(n20664), .Z(n20666) );
  XOR U21178 ( .A(b[51]), .B(a[52]), .Z(n20955) );
  NANDN U21179 ( .A(n37605), .B(n20955), .Z(n20665) );
  AND U21180 ( .A(n20666), .B(n20665), .Z(n21140) );
  NANDN U21181 ( .A(n37705), .B(n20667), .Z(n20669) );
  XOR U21182 ( .A(b[53]), .B(a[50]), .Z(n20958) );
  NANDN U21183 ( .A(n37778), .B(n20958), .Z(n20668) );
  AND U21184 ( .A(n20669), .B(n20668), .Z(n21139) );
  NANDN U21185 ( .A(n36210), .B(n20670), .Z(n20672) );
  XOR U21186 ( .A(b[39]), .B(a[64]), .Z(n20961) );
  NANDN U21187 ( .A(n36347), .B(n20961), .Z(n20671) );
  NAND U21188 ( .A(n20672), .B(n20671), .Z(n21138) );
  XOR U21189 ( .A(n21139), .B(n21138), .Z(n21141) );
  XNOR U21190 ( .A(n21140), .B(n21141), .Z(n21087) );
  XNOR U21191 ( .A(n21088), .B(n21087), .Z(n21090) );
  NANDN U21192 ( .A(n20674), .B(n20673), .Z(n20678) );
  NANDN U21193 ( .A(n20676), .B(n20675), .Z(n20677) );
  AND U21194 ( .A(n20678), .B(n20677), .Z(n21089) );
  XOR U21195 ( .A(n21090), .B(n21089), .Z(n20937) );
  NANDN U21196 ( .A(n20680), .B(n20679), .Z(n20684) );
  OR U21197 ( .A(n20682), .B(n20681), .Z(n20683) );
  AND U21198 ( .A(n20684), .B(n20683), .Z(n20935) );
  NANDN U21199 ( .A(n20686), .B(n20685), .Z(n20690) );
  NANDN U21200 ( .A(n20688), .B(n20687), .Z(n20689) );
  NAND U21201 ( .A(n20690), .B(n20689), .Z(n20934) );
  XNOR U21202 ( .A(n20935), .B(n20934), .Z(n20936) );
  XNOR U21203 ( .A(n20937), .B(n20936), .Z(n20910) );
  XOR U21204 ( .A(n20911), .B(n20910), .Z(n20913) );
  XOR U21205 ( .A(n20912), .B(n20913), .Z(n20899) );
  NANDN U21206 ( .A(n29499), .B(n20691), .Z(n20693) );
  XOR U21207 ( .A(a[96]), .B(b[7]), .Z(n21012) );
  NANDN U21208 ( .A(n29735), .B(n21012), .Z(n20692) );
  AND U21209 ( .A(n20693), .B(n20692), .Z(n20972) );
  NANDN U21210 ( .A(n37857), .B(n20694), .Z(n20696) );
  XOR U21211 ( .A(b[55]), .B(a[48]), .Z(n21015) );
  NANDN U21212 ( .A(n37911), .B(n21015), .Z(n20695) );
  AND U21213 ( .A(n20696), .B(n20695), .Z(n20971) );
  NANDN U21214 ( .A(n35611), .B(n20697), .Z(n20699) );
  XOR U21215 ( .A(b[35]), .B(a[68]), .Z(n21018) );
  NANDN U21216 ( .A(n35801), .B(n21018), .Z(n20698) );
  NAND U21217 ( .A(n20699), .B(n20698), .Z(n20970) );
  XOR U21218 ( .A(n20971), .B(n20970), .Z(n20973) );
  XOR U21219 ( .A(n20972), .B(n20973), .Z(n21034) );
  NANDN U21220 ( .A(n20701), .B(n20700), .Z(n20705) );
  NANDN U21221 ( .A(n20703), .B(n20702), .Z(n20704) );
  AND U21222 ( .A(n20705), .B(n20704), .Z(n21033) );
  XNOR U21223 ( .A(n21034), .B(n21033), .Z(n21035) );
  NANDN U21224 ( .A(n20707), .B(n20706), .Z(n20711) );
  OR U21225 ( .A(n20709), .B(n20708), .Z(n20710) );
  NAND U21226 ( .A(n20711), .B(n20710), .Z(n21036) );
  XNOR U21227 ( .A(n21035), .B(n21036), .Z(n20918) );
  NAND U21228 ( .A(n20713), .B(n20712), .Z(n20717) );
  NANDN U21229 ( .A(n20715), .B(n20714), .Z(n20716) );
  AND U21230 ( .A(n20717), .B(n20716), .Z(n20917) );
  NANDN U21231 ( .A(n211), .B(n20718), .Z(n20720) );
  XOR U21232 ( .A(b[47]), .B(a[56]), .Z(n20988) );
  NANDN U21233 ( .A(n37172), .B(n20988), .Z(n20719) );
  AND U21234 ( .A(n20720), .B(n20719), .Z(n21029) );
  NANDN U21235 ( .A(n210), .B(n20721), .Z(n20723) );
  XOR U21236 ( .A(a[94]), .B(b[9]), .Z(n20991) );
  NANDN U21237 ( .A(n30267), .B(n20991), .Z(n20722) );
  AND U21238 ( .A(n20723), .B(n20722), .Z(n21028) );
  NANDN U21239 ( .A(n212), .B(n20724), .Z(n20726) );
  XOR U21240 ( .A(b[49]), .B(a[54]), .Z(n20994) );
  NANDN U21241 ( .A(n37432), .B(n20994), .Z(n20725) );
  NAND U21242 ( .A(n20726), .B(n20725), .Z(n21027) );
  XOR U21243 ( .A(n21028), .B(n21027), .Z(n21030) );
  XOR U21244 ( .A(n21029), .B(n21030), .Z(n21094) );
  NANDN U21245 ( .A(n36742), .B(n20727), .Z(n20729) );
  XOR U21246 ( .A(b[43]), .B(a[60]), .Z(n20997) );
  NANDN U21247 ( .A(n36891), .B(n20997), .Z(n20728) );
  AND U21248 ( .A(n20729), .B(n20728), .Z(n21008) );
  NANDN U21249 ( .A(n36991), .B(n20730), .Z(n20732) );
  XOR U21250 ( .A(b[45]), .B(a[58]), .Z(n21000) );
  NANDN U21251 ( .A(n37083), .B(n21000), .Z(n20731) );
  AND U21252 ( .A(n20732), .B(n20731), .Z(n21007) );
  NANDN U21253 ( .A(n30482), .B(n20733), .Z(n20735) );
  XOR U21254 ( .A(a[92]), .B(b[11]), .Z(n21003) );
  NANDN U21255 ( .A(n30891), .B(n21003), .Z(n20734) );
  NAND U21256 ( .A(n20735), .B(n20734), .Z(n21006) );
  XOR U21257 ( .A(n21007), .B(n21006), .Z(n21009) );
  XNOR U21258 ( .A(n21008), .B(n21009), .Z(n21093) );
  XNOR U21259 ( .A(n21094), .B(n21093), .Z(n21095) );
  NANDN U21260 ( .A(n20737), .B(n20736), .Z(n20741) );
  OR U21261 ( .A(n20739), .B(n20738), .Z(n20740) );
  NAND U21262 ( .A(n20741), .B(n20740), .Z(n21096) );
  XNOR U21263 ( .A(n21095), .B(n21096), .Z(n20916) );
  XOR U21264 ( .A(n20917), .B(n20916), .Z(n20919) );
  XNOR U21265 ( .A(n20918), .B(n20919), .Z(n20898) );
  XOR U21266 ( .A(n20899), .B(n20898), .Z(n20901) );
  XOR U21267 ( .A(n20900), .B(n20901), .Z(n20887) );
  NAND U21268 ( .A(n20743), .B(n20742), .Z(n20747) );
  NANDN U21269 ( .A(n20745), .B(n20744), .Z(n20746) );
  NAND U21270 ( .A(n20747), .B(n20746), .Z(n20904) );
  NANDN U21271 ( .A(n20749), .B(n20748), .Z(n20753) );
  NAND U21272 ( .A(n20751), .B(n20750), .Z(n20752) );
  AND U21273 ( .A(n20753), .B(n20752), .Z(n20905) );
  XOR U21274 ( .A(n20904), .B(n20905), .Z(n20907) );
  NANDN U21275 ( .A(n20755), .B(n20754), .Z(n20759) );
  NANDN U21276 ( .A(n20757), .B(n20756), .Z(n20758) );
  NAND U21277 ( .A(n20759), .B(n20758), .Z(n20906) );
  XOR U21278 ( .A(n20907), .B(n20906), .Z(n20925) );
  NANDN U21279 ( .A(n20761), .B(n20760), .Z(n20765) );
  OR U21280 ( .A(n20763), .B(n20762), .Z(n20764) );
  AND U21281 ( .A(n20765), .B(n20764), .Z(n21046) );
  NANDN U21282 ( .A(n20767), .B(n20766), .Z(n20771) );
  NANDN U21283 ( .A(n20769), .B(n20768), .Z(n20770) );
  NAND U21284 ( .A(n20771), .B(n20770), .Z(n21045) );
  XNOR U21285 ( .A(n21046), .B(n21045), .Z(n21048) );
  NANDN U21286 ( .A(n20773), .B(n20772), .Z(n20777) );
  NANDN U21287 ( .A(n20775), .B(n20774), .Z(n20776) );
  AND U21288 ( .A(n20777), .B(n20776), .Z(n20943) );
  NAND U21289 ( .A(b[0]), .B(a[102]), .Z(n20778) );
  XNOR U21290 ( .A(b[1]), .B(n20778), .Z(n20780) );
  NANDN U21291 ( .A(b[0]), .B(a[101]), .Z(n20779) );
  NAND U21292 ( .A(n20780), .B(n20779), .Z(n20979) );
  NANDN U21293 ( .A(n38278), .B(n20781), .Z(n20783) );
  XOR U21294 ( .A(b[63]), .B(a[40]), .Z(n21072) );
  NANDN U21295 ( .A(n38279), .B(n21072), .Z(n20782) );
  AND U21296 ( .A(n20783), .B(n20782), .Z(n20977) );
  NANDN U21297 ( .A(n35260), .B(n20784), .Z(n20786) );
  XOR U21298 ( .A(b[33]), .B(a[70]), .Z(n21075) );
  NANDN U21299 ( .A(n35456), .B(n21075), .Z(n20785) );
  NAND U21300 ( .A(n20786), .B(n20785), .Z(n20976) );
  XNOR U21301 ( .A(n20977), .B(n20976), .Z(n20978) );
  XNOR U21302 ( .A(n20979), .B(n20978), .Z(n20940) );
  NANDN U21303 ( .A(n37974), .B(n20787), .Z(n20789) );
  XOR U21304 ( .A(b[57]), .B(a[46]), .Z(n21078) );
  NANDN U21305 ( .A(n38031), .B(n21078), .Z(n20788) );
  AND U21306 ( .A(n20789), .B(n20788), .Z(n21054) );
  NANDN U21307 ( .A(n38090), .B(n20790), .Z(n20792) );
  XOR U21308 ( .A(b[59]), .B(a[44]), .Z(n21081) );
  NANDN U21309 ( .A(n38130), .B(n21081), .Z(n20791) );
  AND U21310 ( .A(n20792), .B(n20791), .Z(n21052) );
  NANDN U21311 ( .A(n36480), .B(n20793), .Z(n20795) );
  XOR U21312 ( .A(b[41]), .B(a[62]), .Z(n21084) );
  NANDN U21313 ( .A(n36594), .B(n21084), .Z(n20794) );
  NAND U21314 ( .A(n20795), .B(n20794), .Z(n21051) );
  XNOR U21315 ( .A(n21052), .B(n21051), .Z(n21053) );
  XOR U21316 ( .A(n21054), .B(n21053), .Z(n20941) );
  XNOR U21317 ( .A(n20940), .B(n20941), .Z(n20942) );
  XNOR U21318 ( .A(n20943), .B(n20942), .Z(n21047) );
  XOR U21319 ( .A(n21048), .B(n21047), .Z(n20929) );
  NANDN U21320 ( .A(n20797), .B(n20796), .Z(n20801) );
  NAND U21321 ( .A(n20799), .B(n20798), .Z(n20800) );
  NAND U21322 ( .A(n20801), .B(n20800), .Z(n20928) );
  XNOR U21323 ( .A(n20929), .B(n20928), .Z(n20931) );
  NANDN U21324 ( .A(n20803), .B(n20802), .Z(n20807) );
  NANDN U21325 ( .A(n20805), .B(n20804), .Z(n20806) );
  AND U21326 ( .A(n20807), .B(n20806), .Z(n21147) );
  NANDN U21327 ( .A(n32996), .B(n20808), .Z(n20810) );
  XOR U21328 ( .A(b[21]), .B(a[82]), .Z(n21099) );
  NANDN U21329 ( .A(n33271), .B(n21099), .Z(n20809) );
  AND U21330 ( .A(n20810), .B(n20809), .Z(n21065) );
  NANDN U21331 ( .A(n33866), .B(n20811), .Z(n20813) );
  XOR U21332 ( .A(b[23]), .B(a[80]), .Z(n21102) );
  NANDN U21333 ( .A(n33644), .B(n21102), .Z(n20812) );
  AND U21334 ( .A(n20813), .B(n20812), .Z(n21064) );
  NANDN U21335 ( .A(n32483), .B(n20814), .Z(n20816) );
  XOR U21336 ( .A(b[19]), .B(a[84]), .Z(n21105) );
  NANDN U21337 ( .A(n32823), .B(n21105), .Z(n20815) );
  NAND U21338 ( .A(n20816), .B(n20815), .Z(n21063) );
  XOR U21339 ( .A(n21064), .B(n21063), .Z(n21066) );
  XOR U21340 ( .A(n21065), .B(n21066), .Z(n20983) );
  NANDN U21341 ( .A(n34909), .B(n20817), .Z(n20819) );
  XOR U21342 ( .A(b[31]), .B(a[72]), .Z(n21108) );
  NANDN U21343 ( .A(n35145), .B(n21108), .Z(n20818) );
  AND U21344 ( .A(n20819), .B(n20818), .Z(n21023) );
  NANDN U21345 ( .A(n38247), .B(n20820), .Z(n20822) );
  XOR U21346 ( .A(b[61]), .B(a[42]), .Z(n21111) );
  NANDN U21347 ( .A(n38248), .B(n21111), .Z(n20821) );
  AND U21348 ( .A(n20822), .B(n20821), .Z(n21022) );
  AND U21349 ( .A(b[63]), .B(a[38]), .Z(n21021) );
  XOR U21350 ( .A(n21022), .B(n21021), .Z(n21024) );
  XNOR U21351 ( .A(n21023), .B(n21024), .Z(n20982) );
  XNOR U21352 ( .A(n20983), .B(n20982), .Z(n20984) );
  NANDN U21353 ( .A(n20824), .B(n20823), .Z(n20828) );
  OR U21354 ( .A(n20826), .B(n20825), .Z(n20827) );
  NAND U21355 ( .A(n20828), .B(n20827), .Z(n20985) );
  XNOR U21356 ( .A(n20984), .B(n20985), .Z(n21144) );
  NANDN U21357 ( .A(n34223), .B(n20829), .Z(n20831) );
  XOR U21358 ( .A(b[27]), .B(a[76]), .Z(n21120) );
  NANDN U21359 ( .A(n34458), .B(n21120), .Z(n20830) );
  AND U21360 ( .A(n20831), .B(n20830), .Z(n20966) );
  NANDN U21361 ( .A(n34634), .B(n20832), .Z(n20834) );
  XOR U21362 ( .A(b[29]), .B(a[74]), .Z(n21123) );
  NANDN U21363 ( .A(n34722), .B(n21123), .Z(n20833) );
  AND U21364 ( .A(n20834), .B(n20833), .Z(n20965) );
  NANDN U21365 ( .A(n31055), .B(n20835), .Z(n20837) );
  XOR U21366 ( .A(a[90]), .B(b[13]), .Z(n21126) );
  NANDN U21367 ( .A(n31293), .B(n21126), .Z(n20836) );
  NAND U21368 ( .A(n20837), .B(n20836), .Z(n20964) );
  XOR U21369 ( .A(n20965), .B(n20964), .Z(n20967) );
  XOR U21370 ( .A(n20966), .B(n20967), .Z(n21040) );
  NANDN U21371 ( .A(n28889), .B(n20838), .Z(n20840) );
  XOR U21372 ( .A(a[98]), .B(b[5]), .Z(n21129) );
  NANDN U21373 ( .A(n29138), .B(n21129), .Z(n20839) );
  AND U21374 ( .A(n20840), .B(n20839), .Z(n21059) );
  NANDN U21375 ( .A(n209), .B(n20841), .Z(n20843) );
  XOR U21376 ( .A(a[100]), .B(b[3]), .Z(n21132) );
  NANDN U21377 ( .A(n28941), .B(n21132), .Z(n20842) );
  AND U21378 ( .A(n20843), .B(n20842), .Z(n21058) );
  NANDN U21379 ( .A(n35936), .B(n20844), .Z(n20846) );
  XOR U21380 ( .A(b[37]), .B(a[66]), .Z(n21135) );
  NANDN U21381 ( .A(n36047), .B(n21135), .Z(n20845) );
  NAND U21382 ( .A(n20846), .B(n20845), .Z(n21057) );
  XOR U21383 ( .A(n21058), .B(n21057), .Z(n21060) );
  XNOR U21384 ( .A(n21059), .B(n21060), .Z(n21039) );
  XNOR U21385 ( .A(n21040), .B(n21039), .Z(n21041) );
  NANDN U21386 ( .A(n20848), .B(n20847), .Z(n20852) );
  OR U21387 ( .A(n20850), .B(n20849), .Z(n20851) );
  NAND U21388 ( .A(n20852), .B(n20851), .Z(n21042) );
  XOR U21389 ( .A(n21041), .B(n21042), .Z(n21145) );
  XNOR U21390 ( .A(n21144), .B(n21145), .Z(n21146) );
  XNOR U21391 ( .A(n21147), .B(n21146), .Z(n20930) );
  XOR U21392 ( .A(n20931), .B(n20930), .Z(n20923) );
  XNOR U21393 ( .A(n20923), .B(n20922), .Z(n20924) );
  XNOR U21394 ( .A(n20925), .B(n20924), .Z(n20886) );
  XNOR U21395 ( .A(n20887), .B(n20886), .Z(n20888) );
  XOR U21396 ( .A(n20889), .B(n20888), .Z(n21153) );
  XNOR U21397 ( .A(n21152), .B(n21153), .Z(n21158) );
  XOR U21398 ( .A(n21159), .B(n21158), .Z(n20881) );
  NANDN U21399 ( .A(n20858), .B(n20857), .Z(n20862) );
  NANDN U21400 ( .A(n20860), .B(n20859), .Z(n20861) );
  AND U21401 ( .A(n20862), .B(n20861), .Z(n20880) );
  XNOR U21402 ( .A(n20881), .B(n20880), .Z(n20882) );
  NANDN U21403 ( .A(n20864), .B(n20863), .Z(n20868) );
  NAND U21404 ( .A(n20866), .B(n20865), .Z(n20867) );
  NAND U21405 ( .A(n20868), .B(n20867), .Z(n20883) );
  XNOR U21406 ( .A(n20882), .B(n20883), .Z(n20874) );
  XNOR U21407 ( .A(n20875), .B(n20874), .Z(n20876) );
  XNOR U21408 ( .A(n20877), .B(n20876), .Z(n21162) );
  XNOR U21409 ( .A(sreg[166]), .B(n21162), .Z(n21164) );
  NANDN U21410 ( .A(sreg[165]), .B(n20869), .Z(n20873) );
  NAND U21411 ( .A(n20871), .B(n20870), .Z(n20872) );
  NAND U21412 ( .A(n20873), .B(n20872), .Z(n21163) );
  XNOR U21413 ( .A(n21164), .B(n21163), .Z(c[166]) );
  NANDN U21414 ( .A(n20875), .B(n20874), .Z(n20879) );
  NANDN U21415 ( .A(n20877), .B(n20876), .Z(n20878) );
  AND U21416 ( .A(n20879), .B(n20878), .Z(n21170) );
  NANDN U21417 ( .A(n20881), .B(n20880), .Z(n20885) );
  NANDN U21418 ( .A(n20883), .B(n20882), .Z(n20884) );
  AND U21419 ( .A(n20885), .B(n20884), .Z(n21168) );
  NANDN U21420 ( .A(n20887), .B(n20886), .Z(n20891) );
  NANDN U21421 ( .A(n20889), .B(n20888), .Z(n20890) );
  AND U21422 ( .A(n20891), .B(n20890), .Z(n21180) );
  NANDN U21423 ( .A(n20893), .B(n20892), .Z(n20897) );
  NANDN U21424 ( .A(n20895), .B(n20894), .Z(n20896) );
  NAND U21425 ( .A(n20897), .B(n20896), .Z(n21179) );
  XNOR U21426 ( .A(n21180), .B(n21179), .Z(n21182) );
  NANDN U21427 ( .A(n20899), .B(n20898), .Z(n20903) );
  OR U21428 ( .A(n20901), .B(n20900), .Z(n20902) );
  AND U21429 ( .A(n20903), .B(n20902), .Z(n21185) );
  NAND U21430 ( .A(n20905), .B(n20904), .Z(n20909) );
  NAND U21431 ( .A(n20907), .B(n20906), .Z(n20908) );
  AND U21432 ( .A(n20909), .B(n20908), .Z(n21451) );
  NANDN U21433 ( .A(n20911), .B(n20910), .Z(n20915) );
  OR U21434 ( .A(n20913), .B(n20912), .Z(n20914) );
  AND U21435 ( .A(n20915), .B(n20914), .Z(n21450) );
  NANDN U21436 ( .A(n20917), .B(n20916), .Z(n20921) );
  NANDN U21437 ( .A(n20919), .B(n20918), .Z(n20920) );
  AND U21438 ( .A(n20921), .B(n20920), .Z(n21449) );
  XOR U21439 ( .A(n21450), .B(n21449), .Z(n21452) );
  XOR U21440 ( .A(n21451), .B(n21452), .Z(n21186) );
  XNOR U21441 ( .A(n21185), .B(n21186), .Z(n21187) );
  NANDN U21442 ( .A(n20923), .B(n20922), .Z(n20927) );
  NANDN U21443 ( .A(n20925), .B(n20924), .Z(n20926) );
  AND U21444 ( .A(n20927), .B(n20926), .Z(n21446) );
  NANDN U21445 ( .A(n20929), .B(n20928), .Z(n20933) );
  NAND U21446 ( .A(n20931), .B(n20930), .Z(n20932) );
  AND U21447 ( .A(n20933), .B(n20932), .Z(n21421) );
  NANDN U21448 ( .A(n20935), .B(n20934), .Z(n20939) );
  NANDN U21449 ( .A(n20937), .B(n20936), .Z(n20938) );
  AND U21450 ( .A(n20939), .B(n20938), .Z(n21439) );
  NANDN U21451 ( .A(n20941), .B(n20940), .Z(n20945) );
  NANDN U21452 ( .A(n20943), .B(n20942), .Z(n20944) );
  AND U21453 ( .A(n20945), .B(n20944), .Z(n21438) );
  NANDN U21454 ( .A(n33875), .B(n20946), .Z(n20948) );
  XOR U21455 ( .A(b[25]), .B(a[79]), .Z(n21215) );
  NANDN U21456 ( .A(n33994), .B(n21215), .Z(n20947) );
  AND U21457 ( .A(n20948), .B(n20947), .Z(n21328) );
  NANDN U21458 ( .A(n32013), .B(n20949), .Z(n20951) );
  XOR U21459 ( .A(a[87]), .B(b[17]), .Z(n21218) );
  NANDN U21460 ( .A(n32292), .B(n21218), .Z(n20950) );
  AND U21461 ( .A(n20951), .B(n20950), .Z(n21327) );
  NANDN U21462 ( .A(n31536), .B(n20952), .Z(n20954) );
  XOR U21463 ( .A(a[89]), .B(b[15]), .Z(n21221) );
  NANDN U21464 ( .A(n31925), .B(n21221), .Z(n20953) );
  NAND U21465 ( .A(n20954), .B(n20953), .Z(n21326) );
  XOR U21466 ( .A(n21327), .B(n21326), .Z(n21329) );
  XOR U21467 ( .A(n21328), .B(n21329), .Z(n21408) );
  NANDN U21468 ( .A(n37526), .B(n20955), .Z(n20957) );
  XOR U21469 ( .A(b[51]), .B(a[53]), .Z(n21224) );
  NANDN U21470 ( .A(n37605), .B(n21224), .Z(n20956) );
  AND U21471 ( .A(n20957), .B(n20956), .Z(n21349) );
  NANDN U21472 ( .A(n37705), .B(n20958), .Z(n20960) );
  XOR U21473 ( .A(b[53]), .B(a[51]), .Z(n21227) );
  NANDN U21474 ( .A(n37778), .B(n21227), .Z(n20959) );
  AND U21475 ( .A(n20960), .B(n20959), .Z(n21348) );
  NANDN U21476 ( .A(n36210), .B(n20961), .Z(n20963) );
  XOR U21477 ( .A(b[39]), .B(a[65]), .Z(n21230) );
  NANDN U21478 ( .A(n36347), .B(n21230), .Z(n20962) );
  NAND U21479 ( .A(n20963), .B(n20962), .Z(n21347) );
  XOR U21480 ( .A(n21348), .B(n21347), .Z(n21350) );
  XNOR U21481 ( .A(n21349), .B(n21350), .Z(n21407) );
  XNOR U21482 ( .A(n21408), .B(n21407), .Z(n21410) );
  NANDN U21483 ( .A(n20965), .B(n20964), .Z(n20969) );
  OR U21484 ( .A(n20967), .B(n20966), .Z(n20968) );
  AND U21485 ( .A(n20969), .B(n20968), .Z(n21409) );
  XOR U21486 ( .A(n21410), .B(n21409), .Z(n21206) );
  NANDN U21487 ( .A(n20971), .B(n20970), .Z(n20975) );
  OR U21488 ( .A(n20973), .B(n20972), .Z(n20974) );
  AND U21489 ( .A(n20975), .B(n20974), .Z(n21204) );
  NANDN U21490 ( .A(n20977), .B(n20976), .Z(n20981) );
  NANDN U21491 ( .A(n20979), .B(n20978), .Z(n20980) );
  NAND U21492 ( .A(n20981), .B(n20980), .Z(n21203) );
  XNOR U21493 ( .A(n21204), .B(n21203), .Z(n21205) );
  XNOR U21494 ( .A(n21206), .B(n21205), .Z(n21437) );
  XOR U21495 ( .A(n21438), .B(n21437), .Z(n21440) );
  XOR U21496 ( .A(n21439), .B(n21440), .Z(n21420) );
  NANDN U21497 ( .A(n20983), .B(n20982), .Z(n20987) );
  NANDN U21498 ( .A(n20985), .B(n20984), .Z(n20986) );
  AND U21499 ( .A(n20987), .B(n20986), .Z(n21432) );
  NAND U21500 ( .A(n37294), .B(n20988), .Z(n20990) );
  XNOR U21501 ( .A(b[47]), .B(a[57]), .Z(n21257) );
  NANDN U21502 ( .A(n21257), .B(n37341), .Z(n20989) );
  NAND U21503 ( .A(n20990), .B(n20989), .Z(n21298) );
  NAND U21504 ( .A(n30627), .B(n20991), .Z(n20993) );
  XNOR U21505 ( .A(a[95]), .B(b[9]), .Z(n21260) );
  NANDN U21506 ( .A(n21260), .B(n30628), .Z(n20992) );
  NAND U21507 ( .A(n20993), .B(n20992), .Z(n21297) );
  NAND U21508 ( .A(n37536), .B(n20994), .Z(n20996) );
  XNOR U21509 ( .A(b[49]), .B(a[55]), .Z(n21263) );
  NANDN U21510 ( .A(n21263), .B(n37537), .Z(n20995) );
  NAND U21511 ( .A(n20996), .B(n20995), .Z(n21296) );
  XNOR U21512 ( .A(n21297), .B(n21296), .Z(n21299) );
  NANDN U21513 ( .A(n36742), .B(n20997), .Z(n20999) );
  XOR U21514 ( .A(b[43]), .B(a[61]), .Z(n21266) );
  NANDN U21515 ( .A(n36891), .B(n21266), .Z(n20998) );
  AND U21516 ( .A(n20999), .B(n20998), .Z(n21277) );
  NANDN U21517 ( .A(n36991), .B(n21000), .Z(n21002) );
  XOR U21518 ( .A(b[45]), .B(a[59]), .Z(n21269) );
  NANDN U21519 ( .A(n37083), .B(n21269), .Z(n21001) );
  AND U21520 ( .A(n21002), .B(n21001), .Z(n21276) );
  NANDN U21521 ( .A(n30482), .B(n21003), .Z(n21005) );
  XOR U21522 ( .A(a[93]), .B(b[11]), .Z(n21272) );
  NANDN U21523 ( .A(n30891), .B(n21272), .Z(n21004) );
  NAND U21524 ( .A(n21005), .B(n21004), .Z(n21275) );
  XOR U21525 ( .A(n21276), .B(n21275), .Z(n21278) );
  XNOR U21526 ( .A(n21277), .B(n21278), .Z(n21320) );
  XOR U21527 ( .A(n21321), .B(n21320), .Z(n21322) );
  NANDN U21528 ( .A(n21007), .B(n21006), .Z(n21011) );
  OR U21529 ( .A(n21009), .B(n21008), .Z(n21010) );
  NAND U21530 ( .A(n21011), .B(n21010), .Z(n21323) );
  XNOR U21531 ( .A(n21322), .B(n21323), .Z(n21431) );
  XNOR U21532 ( .A(n21432), .B(n21431), .Z(n21433) );
  NANDN U21533 ( .A(n29499), .B(n21012), .Z(n21014) );
  XOR U21534 ( .A(a[97]), .B(b[7]), .Z(n21281) );
  NANDN U21535 ( .A(n29735), .B(n21281), .Z(n21013) );
  AND U21536 ( .A(n21014), .B(n21013), .Z(n21241) );
  NANDN U21537 ( .A(n37857), .B(n21015), .Z(n21017) );
  XOR U21538 ( .A(b[55]), .B(a[49]), .Z(n21284) );
  NANDN U21539 ( .A(n37911), .B(n21284), .Z(n21016) );
  AND U21540 ( .A(n21017), .B(n21016), .Z(n21240) );
  NANDN U21541 ( .A(n35611), .B(n21018), .Z(n21020) );
  XOR U21542 ( .A(b[35]), .B(a[69]), .Z(n21287) );
  NANDN U21543 ( .A(n35801), .B(n21287), .Z(n21019) );
  NAND U21544 ( .A(n21020), .B(n21019), .Z(n21239) );
  XOR U21545 ( .A(n21240), .B(n21239), .Z(n21242) );
  XOR U21546 ( .A(n21241), .B(n21242), .Z(n21303) );
  NANDN U21547 ( .A(n21022), .B(n21021), .Z(n21026) );
  OR U21548 ( .A(n21024), .B(n21023), .Z(n21025) );
  AND U21549 ( .A(n21026), .B(n21025), .Z(n21302) );
  XNOR U21550 ( .A(n21303), .B(n21302), .Z(n21304) );
  NANDN U21551 ( .A(n21028), .B(n21027), .Z(n21032) );
  OR U21552 ( .A(n21030), .B(n21029), .Z(n21031) );
  NAND U21553 ( .A(n21032), .B(n21031), .Z(n21305) );
  XOR U21554 ( .A(n21304), .B(n21305), .Z(n21434) );
  XNOR U21555 ( .A(n21433), .B(n21434), .Z(n21419) );
  XOR U21556 ( .A(n21420), .B(n21419), .Z(n21422) );
  XOR U21557 ( .A(n21421), .B(n21422), .Z(n21444) );
  NANDN U21558 ( .A(n21034), .B(n21033), .Z(n21038) );
  NANDN U21559 ( .A(n21036), .B(n21035), .Z(n21037) );
  AND U21560 ( .A(n21038), .B(n21037), .Z(n21427) );
  NANDN U21561 ( .A(n21040), .B(n21039), .Z(n21044) );
  NANDN U21562 ( .A(n21042), .B(n21041), .Z(n21043) );
  AND U21563 ( .A(n21044), .B(n21043), .Z(n21426) );
  NANDN U21564 ( .A(n21046), .B(n21045), .Z(n21050) );
  NAND U21565 ( .A(n21048), .B(n21047), .Z(n21049) );
  AND U21566 ( .A(n21050), .B(n21049), .Z(n21425) );
  XOR U21567 ( .A(n21426), .B(n21425), .Z(n21428) );
  XOR U21568 ( .A(n21427), .B(n21428), .Z(n21194) );
  NANDN U21569 ( .A(n21052), .B(n21051), .Z(n21056) );
  NANDN U21570 ( .A(n21054), .B(n21053), .Z(n21055) );
  AND U21571 ( .A(n21056), .B(n21055), .Z(n21315) );
  NANDN U21572 ( .A(n21058), .B(n21057), .Z(n21062) );
  OR U21573 ( .A(n21060), .B(n21059), .Z(n21061) );
  NAND U21574 ( .A(n21062), .B(n21061), .Z(n21314) );
  XNOR U21575 ( .A(n21315), .B(n21314), .Z(n21317) );
  NANDN U21576 ( .A(n21064), .B(n21063), .Z(n21068) );
  OR U21577 ( .A(n21066), .B(n21065), .Z(n21067) );
  AND U21578 ( .A(n21068), .B(n21067), .Z(n21212) );
  NAND U21579 ( .A(b[0]), .B(a[103]), .Z(n21069) );
  XNOR U21580 ( .A(b[1]), .B(n21069), .Z(n21071) );
  NANDN U21581 ( .A(b[0]), .B(a[102]), .Z(n21070) );
  NAND U21582 ( .A(n21071), .B(n21070), .Z(n21248) );
  NANDN U21583 ( .A(n38278), .B(n21072), .Z(n21074) );
  XOR U21584 ( .A(b[63]), .B(a[41]), .Z(n21389) );
  NANDN U21585 ( .A(n38279), .B(n21389), .Z(n21073) );
  AND U21586 ( .A(n21074), .B(n21073), .Z(n21246) );
  NANDN U21587 ( .A(n35260), .B(n21075), .Z(n21077) );
  XOR U21588 ( .A(b[33]), .B(a[71]), .Z(n21392) );
  NANDN U21589 ( .A(n35456), .B(n21392), .Z(n21076) );
  NAND U21590 ( .A(n21077), .B(n21076), .Z(n21245) );
  XNOR U21591 ( .A(n21246), .B(n21245), .Z(n21247) );
  XNOR U21592 ( .A(n21248), .B(n21247), .Z(n21209) );
  NANDN U21593 ( .A(n37974), .B(n21078), .Z(n21080) );
  XOR U21594 ( .A(b[57]), .B(a[47]), .Z(n21398) );
  NANDN U21595 ( .A(n38031), .B(n21398), .Z(n21079) );
  AND U21596 ( .A(n21080), .B(n21079), .Z(n21374) );
  NANDN U21597 ( .A(n38090), .B(n21081), .Z(n21083) );
  XOR U21598 ( .A(b[59]), .B(a[45]), .Z(n21401) );
  NANDN U21599 ( .A(n38130), .B(n21401), .Z(n21082) );
  AND U21600 ( .A(n21083), .B(n21082), .Z(n21372) );
  NANDN U21601 ( .A(n36480), .B(n21084), .Z(n21086) );
  XOR U21602 ( .A(b[41]), .B(a[63]), .Z(n21404) );
  NANDN U21603 ( .A(n36594), .B(n21404), .Z(n21085) );
  NAND U21604 ( .A(n21086), .B(n21085), .Z(n21371) );
  XNOR U21605 ( .A(n21372), .B(n21371), .Z(n21373) );
  XOR U21606 ( .A(n21374), .B(n21373), .Z(n21210) );
  XNOR U21607 ( .A(n21209), .B(n21210), .Z(n21211) );
  XNOR U21608 ( .A(n21212), .B(n21211), .Z(n21316) );
  XOR U21609 ( .A(n21317), .B(n21316), .Z(n21198) );
  NANDN U21610 ( .A(n21088), .B(n21087), .Z(n21092) );
  NAND U21611 ( .A(n21090), .B(n21089), .Z(n21091) );
  NAND U21612 ( .A(n21092), .B(n21091), .Z(n21197) );
  XNOR U21613 ( .A(n21198), .B(n21197), .Z(n21200) );
  NANDN U21614 ( .A(n21094), .B(n21093), .Z(n21098) );
  NANDN U21615 ( .A(n21096), .B(n21095), .Z(n21097) );
  AND U21616 ( .A(n21098), .B(n21097), .Z(n21416) );
  NANDN U21617 ( .A(n32996), .B(n21099), .Z(n21101) );
  XOR U21618 ( .A(b[21]), .B(a[83]), .Z(n21332) );
  NANDN U21619 ( .A(n33271), .B(n21332), .Z(n21100) );
  AND U21620 ( .A(n21101), .B(n21100), .Z(n21385) );
  NANDN U21621 ( .A(n33866), .B(n21102), .Z(n21104) );
  XOR U21622 ( .A(b[23]), .B(a[81]), .Z(n21335) );
  NANDN U21623 ( .A(n33644), .B(n21335), .Z(n21103) );
  AND U21624 ( .A(n21104), .B(n21103), .Z(n21384) );
  NANDN U21625 ( .A(n32483), .B(n21105), .Z(n21107) );
  XOR U21626 ( .A(b[19]), .B(a[85]), .Z(n21338) );
  NANDN U21627 ( .A(n32823), .B(n21338), .Z(n21106) );
  NAND U21628 ( .A(n21107), .B(n21106), .Z(n21383) );
  XOR U21629 ( .A(n21384), .B(n21383), .Z(n21386) );
  XOR U21630 ( .A(n21385), .B(n21386), .Z(n21252) );
  NANDN U21631 ( .A(n34909), .B(n21108), .Z(n21110) );
  XOR U21632 ( .A(b[31]), .B(a[73]), .Z(n21341) );
  NANDN U21633 ( .A(n35145), .B(n21341), .Z(n21109) );
  AND U21634 ( .A(n21110), .B(n21109), .Z(n21292) );
  NANDN U21635 ( .A(n38247), .B(n21111), .Z(n21113) );
  XOR U21636 ( .A(b[61]), .B(a[43]), .Z(n21344) );
  NANDN U21637 ( .A(n38248), .B(n21344), .Z(n21112) );
  AND U21638 ( .A(n21113), .B(n21112), .Z(n21291) );
  AND U21639 ( .A(b[63]), .B(a[39]), .Z(n21290) );
  XOR U21640 ( .A(n21291), .B(n21290), .Z(n21293) );
  XNOR U21641 ( .A(n21292), .B(n21293), .Z(n21251) );
  XNOR U21642 ( .A(n21252), .B(n21251), .Z(n21253) );
  NANDN U21643 ( .A(n21115), .B(n21114), .Z(n21119) );
  OR U21644 ( .A(n21117), .B(n21116), .Z(n21118) );
  NAND U21645 ( .A(n21119), .B(n21118), .Z(n21254) );
  XNOR U21646 ( .A(n21253), .B(n21254), .Z(n21413) );
  NANDN U21647 ( .A(n34223), .B(n21120), .Z(n21122) );
  XOR U21648 ( .A(b[27]), .B(a[77]), .Z(n21353) );
  NANDN U21649 ( .A(n34458), .B(n21353), .Z(n21121) );
  AND U21650 ( .A(n21122), .B(n21121), .Z(n21235) );
  NANDN U21651 ( .A(n34634), .B(n21123), .Z(n21125) );
  XOR U21652 ( .A(b[29]), .B(a[75]), .Z(n21356) );
  NANDN U21653 ( .A(n34722), .B(n21356), .Z(n21124) );
  AND U21654 ( .A(n21125), .B(n21124), .Z(n21234) );
  NANDN U21655 ( .A(n31055), .B(n21126), .Z(n21128) );
  XOR U21656 ( .A(a[91]), .B(b[13]), .Z(n21359) );
  NANDN U21657 ( .A(n31293), .B(n21359), .Z(n21127) );
  NAND U21658 ( .A(n21128), .B(n21127), .Z(n21233) );
  XOR U21659 ( .A(n21234), .B(n21233), .Z(n21236) );
  XOR U21660 ( .A(n21235), .B(n21236), .Z(n21309) );
  NANDN U21661 ( .A(n28889), .B(n21129), .Z(n21131) );
  XOR U21662 ( .A(a[99]), .B(b[5]), .Z(n21362) );
  NANDN U21663 ( .A(n29138), .B(n21362), .Z(n21130) );
  AND U21664 ( .A(n21131), .B(n21130), .Z(n21379) );
  NANDN U21665 ( .A(n209), .B(n21132), .Z(n21134) );
  XOR U21666 ( .A(a[101]), .B(b[3]), .Z(n21365) );
  NANDN U21667 ( .A(n28941), .B(n21365), .Z(n21133) );
  AND U21668 ( .A(n21134), .B(n21133), .Z(n21378) );
  NANDN U21669 ( .A(n35936), .B(n21135), .Z(n21137) );
  XOR U21670 ( .A(b[37]), .B(a[67]), .Z(n21368) );
  NANDN U21671 ( .A(n36047), .B(n21368), .Z(n21136) );
  NAND U21672 ( .A(n21137), .B(n21136), .Z(n21377) );
  XOR U21673 ( .A(n21378), .B(n21377), .Z(n21380) );
  XNOR U21674 ( .A(n21379), .B(n21380), .Z(n21308) );
  XNOR U21675 ( .A(n21309), .B(n21308), .Z(n21310) );
  NANDN U21676 ( .A(n21139), .B(n21138), .Z(n21143) );
  OR U21677 ( .A(n21141), .B(n21140), .Z(n21142) );
  NAND U21678 ( .A(n21143), .B(n21142), .Z(n21311) );
  XOR U21679 ( .A(n21310), .B(n21311), .Z(n21414) );
  XNOR U21680 ( .A(n21413), .B(n21414), .Z(n21415) );
  XNOR U21681 ( .A(n21416), .B(n21415), .Z(n21199) );
  XOR U21682 ( .A(n21200), .B(n21199), .Z(n21192) );
  NANDN U21683 ( .A(n21145), .B(n21144), .Z(n21149) );
  NANDN U21684 ( .A(n21147), .B(n21146), .Z(n21148) );
  AND U21685 ( .A(n21149), .B(n21148), .Z(n21191) );
  XNOR U21686 ( .A(n21192), .B(n21191), .Z(n21193) );
  XNOR U21687 ( .A(n21194), .B(n21193), .Z(n21443) );
  XNOR U21688 ( .A(n21444), .B(n21443), .Z(n21445) );
  XOR U21689 ( .A(n21446), .B(n21445), .Z(n21188) );
  XNOR U21690 ( .A(n21187), .B(n21188), .Z(n21181) );
  XOR U21691 ( .A(n21182), .B(n21181), .Z(n21174) );
  NANDN U21692 ( .A(n21151), .B(n21150), .Z(n21155) );
  NANDN U21693 ( .A(n21153), .B(n21152), .Z(n21154) );
  AND U21694 ( .A(n21155), .B(n21154), .Z(n21173) );
  XNOR U21695 ( .A(n21174), .B(n21173), .Z(n21175) );
  NANDN U21696 ( .A(n21157), .B(n21156), .Z(n21161) );
  NAND U21697 ( .A(n21159), .B(n21158), .Z(n21160) );
  NAND U21698 ( .A(n21161), .B(n21160), .Z(n21176) );
  XNOR U21699 ( .A(n21175), .B(n21176), .Z(n21167) );
  XNOR U21700 ( .A(n21168), .B(n21167), .Z(n21169) );
  XNOR U21701 ( .A(n21170), .B(n21169), .Z(n21455) );
  XNOR U21702 ( .A(sreg[167]), .B(n21455), .Z(n21457) );
  NANDN U21703 ( .A(sreg[166]), .B(n21162), .Z(n21166) );
  NAND U21704 ( .A(n21164), .B(n21163), .Z(n21165) );
  NAND U21705 ( .A(n21166), .B(n21165), .Z(n21456) );
  XNOR U21706 ( .A(n21457), .B(n21456), .Z(c[167]) );
  NANDN U21707 ( .A(n21168), .B(n21167), .Z(n21172) );
  NANDN U21708 ( .A(n21170), .B(n21169), .Z(n21171) );
  AND U21709 ( .A(n21172), .B(n21171), .Z(n21463) );
  NANDN U21710 ( .A(n21174), .B(n21173), .Z(n21178) );
  NANDN U21711 ( .A(n21176), .B(n21175), .Z(n21177) );
  AND U21712 ( .A(n21178), .B(n21177), .Z(n21461) );
  NANDN U21713 ( .A(n21180), .B(n21179), .Z(n21184) );
  NAND U21714 ( .A(n21182), .B(n21181), .Z(n21183) );
  AND U21715 ( .A(n21184), .B(n21183), .Z(n21468) );
  NANDN U21716 ( .A(n21186), .B(n21185), .Z(n21190) );
  NANDN U21717 ( .A(n21188), .B(n21187), .Z(n21189) );
  AND U21718 ( .A(n21190), .B(n21189), .Z(n21467) );
  NANDN U21719 ( .A(n21192), .B(n21191), .Z(n21196) );
  NANDN U21720 ( .A(n21194), .B(n21193), .Z(n21195) );
  AND U21721 ( .A(n21196), .B(n21195), .Z(n21474) );
  NANDN U21722 ( .A(n21198), .B(n21197), .Z(n21202) );
  NAND U21723 ( .A(n21200), .B(n21199), .Z(n21201) );
  AND U21724 ( .A(n21202), .B(n21201), .Z(n21504) );
  NANDN U21725 ( .A(n21204), .B(n21203), .Z(n21208) );
  NANDN U21726 ( .A(n21206), .B(n21205), .Z(n21207) );
  AND U21727 ( .A(n21208), .B(n21207), .Z(n21498) );
  NANDN U21728 ( .A(n21210), .B(n21209), .Z(n21214) );
  NANDN U21729 ( .A(n21212), .B(n21211), .Z(n21213) );
  AND U21730 ( .A(n21214), .B(n21213), .Z(n21497) );
  NANDN U21731 ( .A(n33875), .B(n21215), .Z(n21217) );
  XOR U21732 ( .A(b[25]), .B(a[80]), .Z(n21532) );
  NANDN U21733 ( .A(n33994), .B(n21532), .Z(n21216) );
  AND U21734 ( .A(n21217), .B(n21216), .Z(n21660) );
  NANDN U21735 ( .A(n32013), .B(n21218), .Z(n21220) );
  XOR U21736 ( .A(a[88]), .B(b[17]), .Z(n21535) );
  NANDN U21737 ( .A(n32292), .B(n21535), .Z(n21219) );
  AND U21738 ( .A(n21220), .B(n21219), .Z(n21659) );
  NANDN U21739 ( .A(n31536), .B(n21221), .Z(n21223) );
  XOR U21740 ( .A(a[90]), .B(b[15]), .Z(n21538) );
  NANDN U21741 ( .A(n31925), .B(n21538), .Z(n21222) );
  NAND U21742 ( .A(n21223), .B(n21222), .Z(n21658) );
  XOR U21743 ( .A(n21659), .B(n21658), .Z(n21661) );
  XOR U21744 ( .A(n21660), .B(n21661), .Z(n21725) );
  NANDN U21745 ( .A(n37526), .B(n21224), .Z(n21226) );
  XOR U21746 ( .A(b[51]), .B(a[54]), .Z(n21541) );
  NANDN U21747 ( .A(n37605), .B(n21541), .Z(n21225) );
  AND U21748 ( .A(n21226), .B(n21225), .Z(n21684) );
  NANDN U21749 ( .A(n37705), .B(n21227), .Z(n21229) );
  XOR U21750 ( .A(b[53]), .B(a[52]), .Z(n21544) );
  NANDN U21751 ( .A(n37778), .B(n21544), .Z(n21228) );
  AND U21752 ( .A(n21229), .B(n21228), .Z(n21683) );
  NANDN U21753 ( .A(n36210), .B(n21230), .Z(n21232) );
  XOR U21754 ( .A(b[39]), .B(a[66]), .Z(n21547) );
  NANDN U21755 ( .A(n36347), .B(n21547), .Z(n21231) );
  NAND U21756 ( .A(n21232), .B(n21231), .Z(n21682) );
  XOR U21757 ( .A(n21683), .B(n21682), .Z(n21685) );
  XNOR U21758 ( .A(n21684), .B(n21685), .Z(n21724) );
  XNOR U21759 ( .A(n21725), .B(n21724), .Z(n21727) );
  NANDN U21760 ( .A(n21234), .B(n21233), .Z(n21238) );
  OR U21761 ( .A(n21236), .B(n21235), .Z(n21237) );
  AND U21762 ( .A(n21238), .B(n21237), .Z(n21726) );
  XOR U21763 ( .A(n21727), .B(n21726), .Z(n21523) );
  NANDN U21764 ( .A(n21240), .B(n21239), .Z(n21244) );
  OR U21765 ( .A(n21242), .B(n21241), .Z(n21243) );
  AND U21766 ( .A(n21244), .B(n21243), .Z(n21521) );
  NANDN U21767 ( .A(n21246), .B(n21245), .Z(n21250) );
  NANDN U21768 ( .A(n21248), .B(n21247), .Z(n21249) );
  NAND U21769 ( .A(n21250), .B(n21249), .Z(n21520) );
  XNOR U21770 ( .A(n21521), .B(n21520), .Z(n21522) );
  XNOR U21771 ( .A(n21523), .B(n21522), .Z(n21496) );
  XOR U21772 ( .A(n21497), .B(n21496), .Z(n21499) );
  XOR U21773 ( .A(n21498), .B(n21499), .Z(n21503) );
  NANDN U21774 ( .A(n21252), .B(n21251), .Z(n21256) );
  NANDN U21775 ( .A(n21254), .B(n21253), .Z(n21255) );
  AND U21776 ( .A(n21256), .B(n21255), .Z(n21491) );
  NANDN U21777 ( .A(n21257), .B(n37294), .Z(n21259) );
  XOR U21778 ( .A(b[47]), .B(a[58]), .Z(n21574) );
  NANDN U21779 ( .A(n37172), .B(n21574), .Z(n21258) );
  AND U21780 ( .A(n21259), .B(n21258), .Z(n21615) );
  NANDN U21781 ( .A(n21260), .B(n30627), .Z(n21262) );
  XOR U21782 ( .A(a[96]), .B(b[9]), .Z(n21577) );
  NANDN U21783 ( .A(n30267), .B(n21577), .Z(n21261) );
  AND U21784 ( .A(n21262), .B(n21261), .Z(n21614) );
  NANDN U21785 ( .A(n21263), .B(n37536), .Z(n21265) );
  XOR U21786 ( .A(b[49]), .B(a[56]), .Z(n21580) );
  NANDN U21787 ( .A(n37432), .B(n21580), .Z(n21264) );
  NAND U21788 ( .A(n21265), .B(n21264), .Z(n21613) );
  XOR U21789 ( .A(n21614), .B(n21613), .Z(n21616) );
  XOR U21790 ( .A(n21615), .B(n21616), .Z(n21638) );
  NANDN U21791 ( .A(n36742), .B(n21266), .Z(n21268) );
  XOR U21792 ( .A(b[43]), .B(a[62]), .Z(n21583) );
  NANDN U21793 ( .A(n36891), .B(n21583), .Z(n21267) );
  AND U21794 ( .A(n21268), .B(n21267), .Z(n21594) );
  NANDN U21795 ( .A(n36991), .B(n21269), .Z(n21271) );
  XOR U21796 ( .A(b[45]), .B(a[60]), .Z(n21586) );
  NANDN U21797 ( .A(n37083), .B(n21586), .Z(n21270) );
  AND U21798 ( .A(n21271), .B(n21270), .Z(n21593) );
  NANDN U21799 ( .A(n30482), .B(n21272), .Z(n21274) );
  XOR U21800 ( .A(a[94]), .B(b[11]), .Z(n21589) );
  NANDN U21801 ( .A(n30891), .B(n21589), .Z(n21273) );
  NAND U21802 ( .A(n21274), .B(n21273), .Z(n21592) );
  XOR U21803 ( .A(n21593), .B(n21592), .Z(n21595) );
  XNOR U21804 ( .A(n21594), .B(n21595), .Z(n21637) );
  XNOR U21805 ( .A(n21638), .B(n21637), .Z(n21639) );
  NANDN U21806 ( .A(n21276), .B(n21275), .Z(n21280) );
  OR U21807 ( .A(n21278), .B(n21277), .Z(n21279) );
  NAND U21808 ( .A(n21280), .B(n21279), .Z(n21640) );
  XNOR U21809 ( .A(n21639), .B(n21640), .Z(n21490) );
  XNOR U21810 ( .A(n21491), .B(n21490), .Z(n21492) );
  NANDN U21811 ( .A(n29499), .B(n21281), .Z(n21283) );
  XOR U21812 ( .A(a[98]), .B(b[7]), .Z(n21598) );
  NANDN U21813 ( .A(n29735), .B(n21598), .Z(n21282) );
  AND U21814 ( .A(n21283), .B(n21282), .Z(n21558) );
  NANDN U21815 ( .A(n37857), .B(n21284), .Z(n21286) );
  XOR U21816 ( .A(b[55]), .B(a[50]), .Z(n21601) );
  NANDN U21817 ( .A(n37911), .B(n21601), .Z(n21285) );
  AND U21818 ( .A(n21286), .B(n21285), .Z(n21557) );
  NANDN U21819 ( .A(n35611), .B(n21287), .Z(n21289) );
  XOR U21820 ( .A(b[35]), .B(a[70]), .Z(n21604) );
  NANDN U21821 ( .A(n35801), .B(n21604), .Z(n21288) );
  NAND U21822 ( .A(n21289), .B(n21288), .Z(n21556) );
  XOR U21823 ( .A(n21557), .B(n21556), .Z(n21559) );
  XOR U21824 ( .A(n21558), .B(n21559), .Z(n21632) );
  NANDN U21825 ( .A(n21291), .B(n21290), .Z(n21295) );
  OR U21826 ( .A(n21293), .B(n21292), .Z(n21294) );
  AND U21827 ( .A(n21295), .B(n21294), .Z(n21631) );
  XNOR U21828 ( .A(n21632), .B(n21631), .Z(n21633) );
  NAND U21829 ( .A(n21297), .B(n21296), .Z(n21301) );
  NANDN U21830 ( .A(n21299), .B(n21298), .Z(n21300) );
  NAND U21831 ( .A(n21301), .B(n21300), .Z(n21634) );
  XOR U21832 ( .A(n21633), .B(n21634), .Z(n21493) );
  XNOR U21833 ( .A(n21492), .B(n21493), .Z(n21502) );
  XOR U21834 ( .A(n21503), .B(n21502), .Z(n21505) );
  XOR U21835 ( .A(n21504), .B(n21505), .Z(n21473) );
  NANDN U21836 ( .A(n21303), .B(n21302), .Z(n21307) );
  NANDN U21837 ( .A(n21305), .B(n21304), .Z(n21306) );
  AND U21838 ( .A(n21307), .B(n21306), .Z(n21486) );
  NANDN U21839 ( .A(n21309), .B(n21308), .Z(n21313) );
  NANDN U21840 ( .A(n21311), .B(n21310), .Z(n21312) );
  AND U21841 ( .A(n21313), .B(n21312), .Z(n21485) );
  NANDN U21842 ( .A(n21315), .B(n21314), .Z(n21319) );
  NAND U21843 ( .A(n21317), .B(n21316), .Z(n21318) );
  AND U21844 ( .A(n21319), .B(n21318), .Z(n21484) );
  XOR U21845 ( .A(n21485), .B(n21484), .Z(n21487) );
  XOR U21846 ( .A(n21486), .B(n21487), .Z(n21511) );
  NAND U21847 ( .A(n21321), .B(n21320), .Z(n21325) );
  NANDN U21848 ( .A(n21323), .B(n21322), .Z(n21324) );
  AND U21849 ( .A(n21325), .B(n21324), .Z(n21733) );
  NANDN U21850 ( .A(n21327), .B(n21326), .Z(n21331) );
  OR U21851 ( .A(n21329), .B(n21328), .Z(n21330) );
  AND U21852 ( .A(n21331), .B(n21330), .Z(n21570) );
  NANDN U21853 ( .A(n32996), .B(n21332), .Z(n21334) );
  XOR U21854 ( .A(b[21]), .B(a[84]), .Z(n21643) );
  NANDN U21855 ( .A(n33271), .B(n21643), .Z(n21333) );
  AND U21856 ( .A(n21334), .B(n21333), .Z(n21703) );
  NANDN U21857 ( .A(n33866), .B(n21335), .Z(n21337) );
  XOR U21858 ( .A(b[23]), .B(a[82]), .Z(n21646) );
  NANDN U21859 ( .A(n33644), .B(n21646), .Z(n21336) );
  AND U21860 ( .A(n21337), .B(n21336), .Z(n21701) );
  NANDN U21861 ( .A(n32483), .B(n21338), .Z(n21340) );
  XOR U21862 ( .A(a[86]), .B(b[19]), .Z(n21649) );
  NANDN U21863 ( .A(n32823), .B(n21649), .Z(n21339) );
  NAND U21864 ( .A(n21340), .B(n21339), .Z(n21700) );
  XNOR U21865 ( .A(n21701), .B(n21700), .Z(n21702) );
  XOR U21866 ( .A(n21703), .B(n21702), .Z(n21569) );
  NANDN U21867 ( .A(n34909), .B(n21341), .Z(n21343) );
  XOR U21868 ( .A(b[31]), .B(a[74]), .Z(n21652) );
  NANDN U21869 ( .A(n35145), .B(n21652), .Z(n21342) );
  AND U21870 ( .A(n21343), .B(n21342), .Z(n21610) );
  NANDN U21871 ( .A(n38247), .B(n21344), .Z(n21346) );
  XOR U21872 ( .A(b[61]), .B(a[44]), .Z(n21655) );
  NANDN U21873 ( .A(n38248), .B(n21655), .Z(n21345) );
  AND U21874 ( .A(n21346), .B(n21345), .Z(n21608) );
  AND U21875 ( .A(b[63]), .B(a[40]), .Z(n21607) );
  XNOR U21876 ( .A(n21608), .B(n21607), .Z(n21609) );
  XOR U21877 ( .A(n21610), .B(n21609), .Z(n21568) );
  XNOR U21878 ( .A(n21569), .B(n21568), .Z(n21571) );
  NANDN U21879 ( .A(n21348), .B(n21347), .Z(n21352) );
  OR U21880 ( .A(n21350), .B(n21349), .Z(n21351) );
  AND U21881 ( .A(n21352), .B(n21351), .Z(n21621) );
  NANDN U21882 ( .A(n34223), .B(n21353), .Z(n21355) );
  XOR U21883 ( .A(b[27]), .B(a[78]), .Z(n21664) );
  NANDN U21884 ( .A(n34458), .B(n21664), .Z(n21354) );
  AND U21885 ( .A(n21355), .B(n21354), .Z(n21553) );
  NANDN U21886 ( .A(n34634), .B(n21356), .Z(n21358) );
  XOR U21887 ( .A(b[29]), .B(a[76]), .Z(n21667) );
  NANDN U21888 ( .A(n34722), .B(n21667), .Z(n21357) );
  AND U21889 ( .A(n21358), .B(n21357), .Z(n21551) );
  NANDN U21890 ( .A(n31055), .B(n21359), .Z(n21361) );
  XOR U21891 ( .A(a[92]), .B(b[13]), .Z(n21670) );
  NANDN U21892 ( .A(n31293), .B(n21670), .Z(n21360) );
  NAND U21893 ( .A(n21361), .B(n21360), .Z(n21550) );
  XNOR U21894 ( .A(n21551), .B(n21550), .Z(n21552) );
  XOR U21895 ( .A(n21553), .B(n21552), .Z(n21620) );
  NANDN U21896 ( .A(n28889), .B(n21362), .Z(n21364) );
  XOR U21897 ( .A(a[100]), .B(b[5]), .Z(n21673) );
  NANDN U21898 ( .A(n29138), .B(n21673), .Z(n21363) );
  AND U21899 ( .A(n21364), .B(n21363), .Z(n21697) );
  NANDN U21900 ( .A(n209), .B(n21365), .Z(n21367) );
  XOR U21901 ( .A(a[102]), .B(b[3]), .Z(n21676) );
  NANDN U21902 ( .A(n28941), .B(n21676), .Z(n21366) );
  AND U21903 ( .A(n21367), .B(n21366), .Z(n21695) );
  NANDN U21904 ( .A(n35936), .B(n21368), .Z(n21370) );
  XOR U21905 ( .A(b[37]), .B(a[68]), .Z(n21679) );
  NANDN U21906 ( .A(n36047), .B(n21679), .Z(n21369) );
  NAND U21907 ( .A(n21370), .B(n21369), .Z(n21694) );
  XNOR U21908 ( .A(n21695), .B(n21694), .Z(n21696) );
  XOR U21909 ( .A(n21697), .B(n21696), .Z(n21619) );
  XNOR U21910 ( .A(n21620), .B(n21619), .Z(n21622) );
  XOR U21911 ( .A(n21731), .B(n21730), .Z(n21732) );
  XNOR U21912 ( .A(n21733), .B(n21732), .Z(n21517) );
  NANDN U21913 ( .A(n21372), .B(n21371), .Z(n21376) );
  NANDN U21914 ( .A(n21374), .B(n21373), .Z(n21375) );
  AND U21915 ( .A(n21376), .B(n21375), .Z(n21626) );
  NANDN U21916 ( .A(n21378), .B(n21377), .Z(n21382) );
  OR U21917 ( .A(n21380), .B(n21379), .Z(n21381) );
  NAND U21918 ( .A(n21382), .B(n21381), .Z(n21625) );
  XNOR U21919 ( .A(n21626), .B(n21625), .Z(n21628) );
  NANDN U21920 ( .A(n21384), .B(n21383), .Z(n21388) );
  OR U21921 ( .A(n21386), .B(n21385), .Z(n21387) );
  NAND U21922 ( .A(n21388), .B(n21387), .Z(n21528) );
  NANDN U21923 ( .A(n38278), .B(n21389), .Z(n21391) );
  XOR U21924 ( .A(b[63]), .B(a[42]), .Z(n21709) );
  NANDN U21925 ( .A(n38279), .B(n21709), .Z(n21390) );
  AND U21926 ( .A(n21391), .B(n21390), .Z(n21563) );
  NANDN U21927 ( .A(n35260), .B(n21392), .Z(n21394) );
  XOR U21928 ( .A(b[33]), .B(a[72]), .Z(n21712) );
  NANDN U21929 ( .A(n35456), .B(n21712), .Z(n21393) );
  NAND U21930 ( .A(n21394), .B(n21393), .Z(n21562) );
  XNOR U21931 ( .A(n21563), .B(n21562), .Z(n21564) );
  NAND U21932 ( .A(b[0]), .B(a[104]), .Z(n21395) );
  XNOR U21933 ( .A(b[1]), .B(n21395), .Z(n21397) );
  NANDN U21934 ( .A(b[0]), .B(a[103]), .Z(n21396) );
  NAND U21935 ( .A(n21397), .B(n21396), .Z(n21565) );
  XNOR U21936 ( .A(n21564), .B(n21565), .Z(n21527) );
  NANDN U21937 ( .A(n37974), .B(n21398), .Z(n21400) );
  XOR U21938 ( .A(b[57]), .B(a[48]), .Z(n21715) );
  NANDN U21939 ( .A(n38031), .B(n21715), .Z(n21399) );
  AND U21940 ( .A(n21400), .B(n21399), .Z(n21690) );
  NANDN U21941 ( .A(n38090), .B(n21401), .Z(n21403) );
  XOR U21942 ( .A(b[59]), .B(a[46]), .Z(n21718) );
  NANDN U21943 ( .A(n38130), .B(n21718), .Z(n21402) );
  AND U21944 ( .A(n21403), .B(n21402), .Z(n21689) );
  NANDN U21945 ( .A(n36480), .B(n21404), .Z(n21406) );
  XOR U21946 ( .A(b[41]), .B(a[64]), .Z(n21721) );
  NANDN U21947 ( .A(n36594), .B(n21721), .Z(n21405) );
  NAND U21948 ( .A(n21406), .B(n21405), .Z(n21688) );
  XOR U21949 ( .A(n21689), .B(n21688), .Z(n21691) );
  XOR U21950 ( .A(n21690), .B(n21691), .Z(n21526) );
  XOR U21951 ( .A(n21527), .B(n21526), .Z(n21529) );
  XOR U21952 ( .A(n21528), .B(n21529), .Z(n21627) );
  XOR U21953 ( .A(n21628), .B(n21627), .Z(n21515) );
  NANDN U21954 ( .A(n21408), .B(n21407), .Z(n21412) );
  NAND U21955 ( .A(n21410), .B(n21409), .Z(n21411) );
  NAND U21956 ( .A(n21412), .B(n21411), .Z(n21514) );
  XNOR U21957 ( .A(n21515), .B(n21514), .Z(n21516) );
  XOR U21958 ( .A(n21517), .B(n21516), .Z(n21509) );
  NANDN U21959 ( .A(n21414), .B(n21413), .Z(n21418) );
  NANDN U21960 ( .A(n21416), .B(n21415), .Z(n21417) );
  AND U21961 ( .A(n21418), .B(n21417), .Z(n21508) );
  XNOR U21962 ( .A(n21509), .B(n21508), .Z(n21510) );
  XNOR U21963 ( .A(n21511), .B(n21510), .Z(n21472) );
  XOR U21964 ( .A(n21473), .B(n21472), .Z(n21475) );
  XOR U21965 ( .A(n21474), .B(n21475), .Z(n21736) );
  NANDN U21966 ( .A(n21420), .B(n21419), .Z(n21424) );
  OR U21967 ( .A(n21422), .B(n21421), .Z(n21423) );
  AND U21968 ( .A(n21424), .B(n21423), .Z(n21735) );
  NANDN U21969 ( .A(n21426), .B(n21425), .Z(n21430) );
  OR U21970 ( .A(n21428), .B(n21427), .Z(n21429) );
  AND U21971 ( .A(n21430), .B(n21429), .Z(n21481) );
  NANDN U21972 ( .A(n21432), .B(n21431), .Z(n21436) );
  NANDN U21973 ( .A(n21434), .B(n21433), .Z(n21435) );
  AND U21974 ( .A(n21436), .B(n21435), .Z(n21479) );
  NANDN U21975 ( .A(n21438), .B(n21437), .Z(n21442) );
  OR U21976 ( .A(n21440), .B(n21439), .Z(n21441) );
  AND U21977 ( .A(n21442), .B(n21441), .Z(n21478) );
  XNOR U21978 ( .A(n21479), .B(n21478), .Z(n21480) );
  XNOR U21979 ( .A(n21481), .B(n21480), .Z(n21734) );
  XOR U21980 ( .A(n21735), .B(n21734), .Z(n21737) );
  XOR U21981 ( .A(n21736), .B(n21737), .Z(n21743) );
  NANDN U21982 ( .A(n21444), .B(n21443), .Z(n21448) );
  NANDN U21983 ( .A(n21446), .B(n21445), .Z(n21447) );
  AND U21984 ( .A(n21448), .B(n21447), .Z(n21741) );
  NANDN U21985 ( .A(n21450), .B(n21449), .Z(n21454) );
  NANDN U21986 ( .A(n21452), .B(n21451), .Z(n21453) );
  NAND U21987 ( .A(n21454), .B(n21453), .Z(n21740) );
  XNOR U21988 ( .A(n21741), .B(n21740), .Z(n21742) );
  XNOR U21989 ( .A(n21743), .B(n21742), .Z(n21466) );
  XOR U21990 ( .A(n21467), .B(n21466), .Z(n21469) );
  XNOR U21991 ( .A(n21468), .B(n21469), .Z(n21460) );
  XNOR U21992 ( .A(n21461), .B(n21460), .Z(n21462) );
  XNOR U21993 ( .A(n21463), .B(n21462), .Z(n21746) );
  XNOR U21994 ( .A(sreg[168]), .B(n21746), .Z(n21748) );
  NANDN U21995 ( .A(sreg[167]), .B(n21455), .Z(n21459) );
  NAND U21996 ( .A(n21457), .B(n21456), .Z(n21458) );
  NAND U21997 ( .A(n21459), .B(n21458), .Z(n21747) );
  XNOR U21998 ( .A(n21748), .B(n21747), .Z(c[168]) );
  NANDN U21999 ( .A(n21461), .B(n21460), .Z(n21465) );
  NANDN U22000 ( .A(n21463), .B(n21462), .Z(n21464) );
  AND U22001 ( .A(n21465), .B(n21464), .Z(n21754) );
  NANDN U22002 ( .A(n21467), .B(n21466), .Z(n21471) );
  OR U22003 ( .A(n21469), .B(n21468), .Z(n21470) );
  AND U22004 ( .A(n21471), .B(n21470), .Z(n21751) );
  NANDN U22005 ( .A(n21473), .B(n21472), .Z(n21477) );
  OR U22006 ( .A(n21475), .B(n21474), .Z(n21476) );
  AND U22007 ( .A(n21477), .B(n21476), .Z(n21764) );
  NANDN U22008 ( .A(n21479), .B(n21478), .Z(n21483) );
  NANDN U22009 ( .A(n21481), .B(n21480), .Z(n21482) );
  AND U22010 ( .A(n21483), .B(n21482), .Z(n21763) );
  XNOR U22011 ( .A(n21764), .B(n21763), .Z(n21766) );
  NANDN U22012 ( .A(n21485), .B(n21484), .Z(n21489) );
  OR U22013 ( .A(n21487), .B(n21486), .Z(n21488) );
  AND U22014 ( .A(n21489), .B(n21488), .Z(n22035) );
  NANDN U22015 ( .A(n21491), .B(n21490), .Z(n21495) );
  NANDN U22016 ( .A(n21493), .B(n21492), .Z(n21494) );
  AND U22017 ( .A(n21495), .B(n21494), .Z(n22034) );
  NANDN U22018 ( .A(n21497), .B(n21496), .Z(n21501) );
  OR U22019 ( .A(n21499), .B(n21498), .Z(n21500) );
  AND U22020 ( .A(n21501), .B(n21500), .Z(n22033) );
  XOR U22021 ( .A(n22034), .B(n22033), .Z(n22036) );
  XOR U22022 ( .A(n22035), .B(n22036), .Z(n21770) );
  NANDN U22023 ( .A(n21503), .B(n21502), .Z(n21507) );
  OR U22024 ( .A(n21505), .B(n21504), .Z(n21506) );
  AND U22025 ( .A(n21507), .B(n21506), .Z(n21769) );
  XNOR U22026 ( .A(n21770), .B(n21769), .Z(n21771) );
  NANDN U22027 ( .A(n21509), .B(n21508), .Z(n21513) );
  NANDN U22028 ( .A(n21511), .B(n21510), .Z(n21512) );
  AND U22029 ( .A(n21513), .B(n21512), .Z(n22030) );
  NANDN U22030 ( .A(n21515), .B(n21514), .Z(n21519) );
  NAND U22031 ( .A(n21517), .B(n21516), .Z(n21518) );
  AND U22032 ( .A(n21519), .B(n21518), .Z(n22023) );
  NANDN U22033 ( .A(n21521), .B(n21520), .Z(n21525) );
  NANDN U22034 ( .A(n21523), .B(n21522), .Z(n21524) );
  AND U22035 ( .A(n21525), .B(n21524), .Z(n22011) );
  NAND U22036 ( .A(n21527), .B(n21526), .Z(n21531) );
  NAND U22037 ( .A(n21529), .B(n21528), .Z(n21530) );
  AND U22038 ( .A(n21531), .B(n21530), .Z(n22010) );
  NANDN U22039 ( .A(n33875), .B(n21532), .Z(n21534) );
  XOR U22040 ( .A(b[25]), .B(a[81]), .Z(n21799) );
  NANDN U22041 ( .A(n33994), .B(n21799), .Z(n21533) );
  AND U22042 ( .A(n21534), .B(n21533), .Z(n21969) );
  NANDN U22043 ( .A(n32013), .B(n21535), .Z(n21537) );
  XOR U22044 ( .A(a[89]), .B(b[17]), .Z(n21802) );
  NANDN U22045 ( .A(n32292), .B(n21802), .Z(n21536) );
  AND U22046 ( .A(n21537), .B(n21536), .Z(n21968) );
  NANDN U22047 ( .A(n31536), .B(n21538), .Z(n21540) );
  XOR U22048 ( .A(a[91]), .B(b[15]), .Z(n21805) );
  NANDN U22049 ( .A(n31925), .B(n21805), .Z(n21539) );
  NAND U22050 ( .A(n21540), .B(n21539), .Z(n21967) );
  XOR U22051 ( .A(n21968), .B(n21967), .Z(n21970) );
  XOR U22052 ( .A(n21969), .B(n21970), .Z(n21941) );
  NANDN U22053 ( .A(n37526), .B(n21541), .Z(n21543) );
  XOR U22054 ( .A(b[51]), .B(a[55]), .Z(n21808) );
  NANDN U22055 ( .A(n37605), .B(n21808), .Z(n21542) );
  AND U22056 ( .A(n21543), .B(n21542), .Z(n21993) );
  NANDN U22057 ( .A(n37705), .B(n21544), .Z(n21546) );
  XOR U22058 ( .A(b[53]), .B(a[53]), .Z(n21811) );
  NANDN U22059 ( .A(n37778), .B(n21811), .Z(n21545) );
  AND U22060 ( .A(n21546), .B(n21545), .Z(n21992) );
  NANDN U22061 ( .A(n36210), .B(n21547), .Z(n21549) );
  XOR U22062 ( .A(b[39]), .B(a[67]), .Z(n21814) );
  NANDN U22063 ( .A(n36347), .B(n21814), .Z(n21548) );
  NAND U22064 ( .A(n21549), .B(n21548), .Z(n21991) );
  XOR U22065 ( .A(n21992), .B(n21991), .Z(n21994) );
  XNOR U22066 ( .A(n21993), .B(n21994), .Z(n21940) );
  XNOR U22067 ( .A(n21941), .B(n21940), .Z(n21943) );
  NANDN U22068 ( .A(n21551), .B(n21550), .Z(n21555) );
  NANDN U22069 ( .A(n21553), .B(n21552), .Z(n21554) );
  AND U22070 ( .A(n21555), .B(n21554), .Z(n21942) );
  XOR U22071 ( .A(n21943), .B(n21942), .Z(n21790) );
  NANDN U22072 ( .A(n21557), .B(n21556), .Z(n21561) );
  OR U22073 ( .A(n21559), .B(n21558), .Z(n21560) );
  AND U22074 ( .A(n21561), .B(n21560), .Z(n21788) );
  NANDN U22075 ( .A(n21563), .B(n21562), .Z(n21567) );
  NANDN U22076 ( .A(n21565), .B(n21564), .Z(n21566) );
  NAND U22077 ( .A(n21567), .B(n21566), .Z(n21787) );
  XNOR U22078 ( .A(n21788), .B(n21787), .Z(n21789) );
  XNOR U22079 ( .A(n21790), .B(n21789), .Z(n22009) );
  XOR U22080 ( .A(n22010), .B(n22009), .Z(n22012) );
  XOR U22081 ( .A(n22011), .B(n22012), .Z(n22022) );
  NAND U22082 ( .A(n21569), .B(n21568), .Z(n21573) );
  NANDN U22083 ( .A(n21571), .B(n21570), .Z(n21572) );
  AND U22084 ( .A(n21573), .B(n21572), .Z(n22016) );
  NANDN U22085 ( .A(n211), .B(n21574), .Z(n21576) );
  XOR U22086 ( .A(b[47]), .B(a[59]), .Z(n21841) );
  NANDN U22087 ( .A(n37172), .B(n21841), .Z(n21575) );
  AND U22088 ( .A(n21576), .B(n21575), .Z(n21882) );
  NANDN U22089 ( .A(n210), .B(n21577), .Z(n21579) );
  XOR U22090 ( .A(a[97]), .B(b[9]), .Z(n21844) );
  NANDN U22091 ( .A(n30267), .B(n21844), .Z(n21578) );
  AND U22092 ( .A(n21579), .B(n21578), .Z(n21881) );
  NANDN U22093 ( .A(n212), .B(n21580), .Z(n21582) );
  XOR U22094 ( .A(b[49]), .B(a[57]), .Z(n21847) );
  NANDN U22095 ( .A(n37432), .B(n21847), .Z(n21581) );
  NAND U22096 ( .A(n21582), .B(n21581), .Z(n21880) );
  XOR U22097 ( .A(n21881), .B(n21880), .Z(n21883) );
  XOR U22098 ( .A(n21882), .B(n21883), .Z(n21947) );
  NANDN U22099 ( .A(n36742), .B(n21583), .Z(n21585) );
  XOR U22100 ( .A(b[43]), .B(a[63]), .Z(n21850) );
  NANDN U22101 ( .A(n36891), .B(n21850), .Z(n21584) );
  AND U22102 ( .A(n21585), .B(n21584), .Z(n21861) );
  NANDN U22103 ( .A(n36991), .B(n21586), .Z(n21588) );
  XOR U22104 ( .A(b[45]), .B(a[61]), .Z(n21853) );
  NANDN U22105 ( .A(n37083), .B(n21853), .Z(n21587) );
  AND U22106 ( .A(n21588), .B(n21587), .Z(n21860) );
  NANDN U22107 ( .A(n30482), .B(n21589), .Z(n21591) );
  XOR U22108 ( .A(a[95]), .B(b[11]), .Z(n21856) );
  NANDN U22109 ( .A(n30891), .B(n21856), .Z(n21590) );
  NAND U22110 ( .A(n21591), .B(n21590), .Z(n21859) );
  XOR U22111 ( .A(n21860), .B(n21859), .Z(n21862) );
  XNOR U22112 ( .A(n21861), .B(n21862), .Z(n21946) );
  XNOR U22113 ( .A(n21947), .B(n21946), .Z(n21948) );
  NANDN U22114 ( .A(n21593), .B(n21592), .Z(n21597) );
  OR U22115 ( .A(n21595), .B(n21594), .Z(n21596) );
  NAND U22116 ( .A(n21597), .B(n21596), .Z(n21949) );
  XNOR U22117 ( .A(n21948), .B(n21949), .Z(n22015) );
  XNOR U22118 ( .A(n22016), .B(n22015), .Z(n22017) );
  NANDN U22119 ( .A(n29499), .B(n21598), .Z(n21600) );
  XOR U22120 ( .A(a[99]), .B(b[7]), .Z(n21865) );
  NANDN U22121 ( .A(n29735), .B(n21865), .Z(n21599) );
  AND U22122 ( .A(n21600), .B(n21599), .Z(n21825) );
  NANDN U22123 ( .A(n37857), .B(n21601), .Z(n21603) );
  XOR U22124 ( .A(b[55]), .B(a[51]), .Z(n21868) );
  NANDN U22125 ( .A(n37911), .B(n21868), .Z(n21602) );
  AND U22126 ( .A(n21603), .B(n21602), .Z(n21824) );
  NANDN U22127 ( .A(n35611), .B(n21604), .Z(n21606) );
  XOR U22128 ( .A(b[35]), .B(a[71]), .Z(n21871) );
  NANDN U22129 ( .A(n35801), .B(n21871), .Z(n21605) );
  NAND U22130 ( .A(n21606), .B(n21605), .Z(n21823) );
  XOR U22131 ( .A(n21824), .B(n21823), .Z(n21826) );
  XOR U22132 ( .A(n21825), .B(n21826), .Z(n21887) );
  NANDN U22133 ( .A(n21608), .B(n21607), .Z(n21612) );
  NANDN U22134 ( .A(n21610), .B(n21609), .Z(n21611) );
  AND U22135 ( .A(n21612), .B(n21611), .Z(n21886) );
  XNOR U22136 ( .A(n21887), .B(n21886), .Z(n21888) );
  NANDN U22137 ( .A(n21614), .B(n21613), .Z(n21618) );
  OR U22138 ( .A(n21616), .B(n21615), .Z(n21617) );
  NAND U22139 ( .A(n21618), .B(n21617), .Z(n21889) );
  XOR U22140 ( .A(n21888), .B(n21889), .Z(n22018) );
  XNOR U22141 ( .A(n22017), .B(n22018), .Z(n22021) );
  XOR U22142 ( .A(n22022), .B(n22021), .Z(n22024) );
  XOR U22143 ( .A(n22023), .B(n22024), .Z(n22028) );
  NAND U22144 ( .A(n21620), .B(n21619), .Z(n21624) );
  NANDN U22145 ( .A(n21622), .B(n21621), .Z(n21623) );
  NAND U22146 ( .A(n21624), .B(n21623), .Z(n22003) );
  NANDN U22147 ( .A(n21626), .B(n21625), .Z(n21630) );
  NAND U22148 ( .A(n21628), .B(n21627), .Z(n21629) );
  AND U22149 ( .A(n21630), .B(n21629), .Z(n22004) );
  XOR U22150 ( .A(n22003), .B(n22004), .Z(n22006) );
  NANDN U22151 ( .A(n21632), .B(n21631), .Z(n21636) );
  NANDN U22152 ( .A(n21634), .B(n21633), .Z(n21635) );
  NAND U22153 ( .A(n21636), .B(n21635), .Z(n22005) );
  XOR U22154 ( .A(n22006), .B(n22005), .Z(n21778) );
  NANDN U22155 ( .A(n21638), .B(n21637), .Z(n21642) );
  NANDN U22156 ( .A(n21640), .B(n21639), .Z(n21641) );
  AND U22157 ( .A(n21642), .B(n21641), .Z(n22000) );
  NANDN U22158 ( .A(n32996), .B(n21643), .Z(n21645) );
  XOR U22159 ( .A(b[21]), .B(a[85]), .Z(n21952) );
  NANDN U22160 ( .A(n33271), .B(n21952), .Z(n21644) );
  AND U22161 ( .A(n21645), .B(n21644), .Z(n21918) );
  NANDN U22162 ( .A(n33866), .B(n21646), .Z(n21648) );
  XOR U22163 ( .A(b[23]), .B(a[83]), .Z(n21955) );
  NANDN U22164 ( .A(n33644), .B(n21955), .Z(n21647) );
  AND U22165 ( .A(n21648), .B(n21647), .Z(n21917) );
  NANDN U22166 ( .A(n32483), .B(n21649), .Z(n21651) );
  XOR U22167 ( .A(a[87]), .B(b[19]), .Z(n21958) );
  NANDN U22168 ( .A(n32823), .B(n21958), .Z(n21650) );
  NAND U22169 ( .A(n21651), .B(n21650), .Z(n21916) );
  XOR U22170 ( .A(n21917), .B(n21916), .Z(n21919) );
  XOR U22171 ( .A(n21918), .B(n21919), .Z(n21836) );
  NANDN U22172 ( .A(n34909), .B(n21652), .Z(n21654) );
  XOR U22173 ( .A(b[31]), .B(a[75]), .Z(n21961) );
  NANDN U22174 ( .A(n35145), .B(n21961), .Z(n21653) );
  AND U22175 ( .A(n21654), .B(n21653), .Z(n21876) );
  NANDN U22176 ( .A(n38247), .B(n21655), .Z(n21657) );
  XOR U22177 ( .A(b[61]), .B(a[45]), .Z(n21964) );
  NANDN U22178 ( .A(n38248), .B(n21964), .Z(n21656) );
  AND U22179 ( .A(n21657), .B(n21656), .Z(n21875) );
  AND U22180 ( .A(b[63]), .B(a[41]), .Z(n21874) );
  XOR U22181 ( .A(n21875), .B(n21874), .Z(n21877) );
  XNOR U22182 ( .A(n21876), .B(n21877), .Z(n21835) );
  XNOR U22183 ( .A(n21836), .B(n21835), .Z(n21837) );
  NANDN U22184 ( .A(n21659), .B(n21658), .Z(n21663) );
  OR U22185 ( .A(n21661), .B(n21660), .Z(n21662) );
  NAND U22186 ( .A(n21663), .B(n21662), .Z(n21838) );
  XNOR U22187 ( .A(n21837), .B(n21838), .Z(n21997) );
  NANDN U22188 ( .A(n34223), .B(n21664), .Z(n21666) );
  XOR U22189 ( .A(b[27]), .B(a[79]), .Z(n21973) );
  NANDN U22190 ( .A(n34458), .B(n21973), .Z(n21665) );
  AND U22191 ( .A(n21666), .B(n21665), .Z(n21819) );
  NANDN U22192 ( .A(n34634), .B(n21667), .Z(n21669) );
  XOR U22193 ( .A(b[29]), .B(a[77]), .Z(n21976) );
  NANDN U22194 ( .A(n34722), .B(n21976), .Z(n21668) );
  AND U22195 ( .A(n21669), .B(n21668), .Z(n21818) );
  NANDN U22196 ( .A(n31055), .B(n21670), .Z(n21672) );
  XOR U22197 ( .A(a[93]), .B(b[13]), .Z(n21979) );
  NANDN U22198 ( .A(n31293), .B(n21979), .Z(n21671) );
  NAND U22199 ( .A(n21672), .B(n21671), .Z(n21817) );
  XOR U22200 ( .A(n21818), .B(n21817), .Z(n21820) );
  XOR U22201 ( .A(n21819), .B(n21820), .Z(n21893) );
  NANDN U22202 ( .A(n28889), .B(n21673), .Z(n21675) );
  XOR U22203 ( .A(a[101]), .B(b[5]), .Z(n21982) );
  NANDN U22204 ( .A(n29138), .B(n21982), .Z(n21674) );
  AND U22205 ( .A(n21675), .B(n21674), .Z(n21912) );
  NANDN U22206 ( .A(n209), .B(n21676), .Z(n21678) );
  XOR U22207 ( .A(a[103]), .B(b[3]), .Z(n21985) );
  NANDN U22208 ( .A(n28941), .B(n21985), .Z(n21677) );
  AND U22209 ( .A(n21678), .B(n21677), .Z(n21911) );
  NANDN U22210 ( .A(n35936), .B(n21679), .Z(n21681) );
  XOR U22211 ( .A(b[37]), .B(a[69]), .Z(n21988) );
  NANDN U22212 ( .A(n36047), .B(n21988), .Z(n21680) );
  NAND U22213 ( .A(n21681), .B(n21680), .Z(n21910) );
  XOR U22214 ( .A(n21911), .B(n21910), .Z(n21913) );
  XNOR U22215 ( .A(n21912), .B(n21913), .Z(n21892) );
  XNOR U22216 ( .A(n21893), .B(n21892), .Z(n21894) );
  NANDN U22217 ( .A(n21683), .B(n21682), .Z(n21687) );
  OR U22218 ( .A(n21685), .B(n21684), .Z(n21686) );
  NAND U22219 ( .A(n21687), .B(n21686), .Z(n21895) );
  XOR U22220 ( .A(n21894), .B(n21895), .Z(n21998) );
  XNOR U22221 ( .A(n21997), .B(n21998), .Z(n21999) );
  XNOR U22222 ( .A(n22000), .B(n21999), .Z(n21784) );
  NANDN U22223 ( .A(n21689), .B(n21688), .Z(n21693) );
  OR U22224 ( .A(n21691), .B(n21690), .Z(n21692) );
  AND U22225 ( .A(n21693), .B(n21692), .Z(n21899) );
  NANDN U22226 ( .A(n21695), .B(n21694), .Z(n21699) );
  NANDN U22227 ( .A(n21697), .B(n21696), .Z(n21698) );
  NAND U22228 ( .A(n21699), .B(n21698), .Z(n21898) );
  XNOR U22229 ( .A(n21899), .B(n21898), .Z(n21901) );
  NANDN U22230 ( .A(n21701), .B(n21700), .Z(n21705) );
  NANDN U22231 ( .A(n21703), .B(n21702), .Z(n21704) );
  AND U22232 ( .A(n21705), .B(n21704), .Z(n21796) );
  NAND U22233 ( .A(b[0]), .B(a[105]), .Z(n21706) );
  XNOR U22234 ( .A(b[1]), .B(n21706), .Z(n21708) );
  NANDN U22235 ( .A(b[0]), .B(a[104]), .Z(n21707) );
  NAND U22236 ( .A(n21708), .B(n21707), .Z(n21832) );
  NANDN U22237 ( .A(n38278), .B(n21709), .Z(n21711) );
  XOR U22238 ( .A(b[63]), .B(a[43]), .Z(n21925) );
  NANDN U22239 ( .A(n38279), .B(n21925), .Z(n21710) );
  AND U22240 ( .A(n21711), .B(n21710), .Z(n21830) );
  NANDN U22241 ( .A(n35260), .B(n21712), .Z(n21714) );
  XOR U22242 ( .A(b[33]), .B(a[73]), .Z(n21928) );
  NANDN U22243 ( .A(n35456), .B(n21928), .Z(n21713) );
  NAND U22244 ( .A(n21714), .B(n21713), .Z(n21829) );
  XNOR U22245 ( .A(n21830), .B(n21829), .Z(n21831) );
  XNOR U22246 ( .A(n21832), .B(n21831), .Z(n21793) );
  NANDN U22247 ( .A(n37974), .B(n21715), .Z(n21717) );
  XOR U22248 ( .A(b[57]), .B(a[49]), .Z(n21931) );
  NANDN U22249 ( .A(n38031), .B(n21931), .Z(n21716) );
  AND U22250 ( .A(n21717), .B(n21716), .Z(n21907) );
  NANDN U22251 ( .A(n38090), .B(n21718), .Z(n21720) );
  XOR U22252 ( .A(b[59]), .B(a[47]), .Z(n21934) );
  NANDN U22253 ( .A(n38130), .B(n21934), .Z(n21719) );
  AND U22254 ( .A(n21720), .B(n21719), .Z(n21905) );
  NANDN U22255 ( .A(n36480), .B(n21721), .Z(n21723) );
  XOR U22256 ( .A(b[41]), .B(a[65]), .Z(n21937) );
  NANDN U22257 ( .A(n36594), .B(n21937), .Z(n21722) );
  NAND U22258 ( .A(n21723), .B(n21722), .Z(n21904) );
  XNOR U22259 ( .A(n21905), .B(n21904), .Z(n21906) );
  XOR U22260 ( .A(n21907), .B(n21906), .Z(n21794) );
  XNOR U22261 ( .A(n21793), .B(n21794), .Z(n21795) );
  XNOR U22262 ( .A(n21796), .B(n21795), .Z(n21900) );
  XOR U22263 ( .A(n21901), .B(n21900), .Z(n21782) );
  NANDN U22264 ( .A(n21725), .B(n21724), .Z(n21729) );
  NAND U22265 ( .A(n21727), .B(n21726), .Z(n21728) );
  NAND U22266 ( .A(n21729), .B(n21728), .Z(n21781) );
  XNOR U22267 ( .A(n21782), .B(n21781), .Z(n21783) );
  XOR U22268 ( .A(n21784), .B(n21783), .Z(n21776) );
  XNOR U22269 ( .A(n21776), .B(n21775), .Z(n21777) );
  XNOR U22270 ( .A(n21778), .B(n21777), .Z(n22027) );
  XNOR U22271 ( .A(n22028), .B(n22027), .Z(n22029) );
  XOR U22272 ( .A(n22030), .B(n22029), .Z(n21772) );
  XNOR U22273 ( .A(n21771), .B(n21772), .Z(n21765) );
  XOR U22274 ( .A(n21766), .B(n21765), .Z(n21758) );
  NANDN U22275 ( .A(n21735), .B(n21734), .Z(n21739) );
  OR U22276 ( .A(n21737), .B(n21736), .Z(n21738) );
  NAND U22277 ( .A(n21739), .B(n21738), .Z(n21757) );
  XNOR U22278 ( .A(n21758), .B(n21757), .Z(n21759) );
  NANDN U22279 ( .A(n21741), .B(n21740), .Z(n21745) );
  NANDN U22280 ( .A(n21743), .B(n21742), .Z(n21744) );
  NAND U22281 ( .A(n21745), .B(n21744), .Z(n21760) );
  XOR U22282 ( .A(n21759), .B(n21760), .Z(n21752) );
  XNOR U22283 ( .A(n21751), .B(n21752), .Z(n21753) );
  XNOR U22284 ( .A(n21754), .B(n21753), .Z(n22039) );
  XNOR U22285 ( .A(sreg[169]), .B(n22039), .Z(n22041) );
  NANDN U22286 ( .A(sreg[168]), .B(n21746), .Z(n21750) );
  NAND U22287 ( .A(n21748), .B(n21747), .Z(n21749) );
  NAND U22288 ( .A(n21750), .B(n21749), .Z(n22040) );
  XNOR U22289 ( .A(n22041), .B(n22040), .Z(c[169]) );
  NANDN U22290 ( .A(n21752), .B(n21751), .Z(n21756) );
  NANDN U22291 ( .A(n21754), .B(n21753), .Z(n21755) );
  AND U22292 ( .A(n21756), .B(n21755), .Z(n22047) );
  NANDN U22293 ( .A(n21758), .B(n21757), .Z(n21762) );
  NANDN U22294 ( .A(n21760), .B(n21759), .Z(n21761) );
  AND U22295 ( .A(n21762), .B(n21761), .Z(n22045) );
  NANDN U22296 ( .A(n21764), .B(n21763), .Z(n21768) );
  NAND U22297 ( .A(n21766), .B(n21765), .Z(n21767) );
  AND U22298 ( .A(n21768), .B(n21767), .Z(n22052) );
  NANDN U22299 ( .A(n21770), .B(n21769), .Z(n21774) );
  NANDN U22300 ( .A(n21772), .B(n21771), .Z(n21773) );
  AND U22301 ( .A(n21774), .B(n21773), .Z(n22051) );
  NANDN U22302 ( .A(n21776), .B(n21775), .Z(n21780) );
  NANDN U22303 ( .A(n21778), .B(n21777), .Z(n21779) );
  AND U22304 ( .A(n21780), .B(n21779), .Z(n22058) );
  NANDN U22305 ( .A(n21782), .B(n21781), .Z(n21786) );
  NAND U22306 ( .A(n21784), .B(n21783), .Z(n21785) );
  AND U22307 ( .A(n21786), .B(n21785), .Z(n22088) );
  NANDN U22308 ( .A(n21788), .B(n21787), .Z(n21792) );
  NANDN U22309 ( .A(n21790), .B(n21789), .Z(n21791) );
  AND U22310 ( .A(n21792), .B(n21791), .Z(n22082) );
  NANDN U22311 ( .A(n21794), .B(n21793), .Z(n21798) );
  NANDN U22312 ( .A(n21796), .B(n21795), .Z(n21797) );
  AND U22313 ( .A(n21798), .B(n21797), .Z(n22081) );
  NANDN U22314 ( .A(n33875), .B(n21799), .Z(n21801) );
  XOR U22315 ( .A(b[25]), .B(a[82]), .Z(n22167) );
  NANDN U22316 ( .A(n33994), .B(n22167), .Z(n21800) );
  AND U22317 ( .A(n21801), .B(n21800), .Z(n22286) );
  NANDN U22318 ( .A(n32013), .B(n21802), .Z(n21804) );
  XOR U22319 ( .A(a[90]), .B(b[17]), .Z(n22170) );
  NANDN U22320 ( .A(n32292), .B(n22170), .Z(n21803) );
  AND U22321 ( .A(n21804), .B(n21803), .Z(n22285) );
  NANDN U22322 ( .A(n31536), .B(n21805), .Z(n21807) );
  XOR U22323 ( .A(a[92]), .B(b[15]), .Z(n22173) );
  NANDN U22324 ( .A(n31925), .B(n22173), .Z(n21806) );
  NAND U22325 ( .A(n21807), .B(n21806), .Z(n22284) );
  XOR U22326 ( .A(n22285), .B(n22284), .Z(n22287) );
  XOR U22327 ( .A(n22286), .B(n22287), .Z(n22258) );
  NANDN U22328 ( .A(n37526), .B(n21808), .Z(n21810) );
  XOR U22329 ( .A(b[51]), .B(a[56]), .Z(n22176) );
  NANDN U22330 ( .A(n37605), .B(n22176), .Z(n21809) );
  AND U22331 ( .A(n21810), .B(n21809), .Z(n22310) );
  NANDN U22332 ( .A(n37705), .B(n21811), .Z(n21813) );
  XOR U22333 ( .A(b[53]), .B(a[54]), .Z(n22179) );
  NANDN U22334 ( .A(n37778), .B(n22179), .Z(n21812) );
  AND U22335 ( .A(n21813), .B(n21812), .Z(n22309) );
  NANDN U22336 ( .A(n36210), .B(n21814), .Z(n21816) );
  XOR U22337 ( .A(b[39]), .B(a[68]), .Z(n22182) );
  NANDN U22338 ( .A(n36347), .B(n22182), .Z(n21815) );
  NAND U22339 ( .A(n21816), .B(n21815), .Z(n22308) );
  XOR U22340 ( .A(n22309), .B(n22308), .Z(n22311) );
  XNOR U22341 ( .A(n22310), .B(n22311), .Z(n22257) );
  XNOR U22342 ( .A(n22258), .B(n22257), .Z(n22260) );
  NANDN U22343 ( .A(n21818), .B(n21817), .Z(n21822) );
  OR U22344 ( .A(n21820), .B(n21819), .Z(n21821) );
  AND U22345 ( .A(n21822), .B(n21821), .Z(n22259) );
  XOR U22346 ( .A(n22260), .B(n22259), .Z(n22158) );
  NANDN U22347 ( .A(n21824), .B(n21823), .Z(n21828) );
  OR U22348 ( .A(n21826), .B(n21825), .Z(n21827) );
  AND U22349 ( .A(n21828), .B(n21827), .Z(n22156) );
  NANDN U22350 ( .A(n21830), .B(n21829), .Z(n21834) );
  NANDN U22351 ( .A(n21832), .B(n21831), .Z(n21833) );
  NAND U22352 ( .A(n21834), .B(n21833), .Z(n22155) );
  XNOR U22353 ( .A(n22156), .B(n22155), .Z(n22157) );
  XNOR U22354 ( .A(n22158), .B(n22157), .Z(n22080) );
  XOR U22355 ( .A(n22081), .B(n22080), .Z(n22083) );
  XOR U22356 ( .A(n22082), .B(n22083), .Z(n22087) );
  NANDN U22357 ( .A(n21836), .B(n21835), .Z(n21840) );
  NANDN U22358 ( .A(n21838), .B(n21837), .Z(n21839) );
  AND U22359 ( .A(n21840), .B(n21839), .Z(n22075) );
  NANDN U22360 ( .A(n211), .B(n21841), .Z(n21843) );
  XOR U22361 ( .A(b[47]), .B(a[60]), .Z(n22110) );
  NANDN U22362 ( .A(n37172), .B(n22110), .Z(n21842) );
  AND U22363 ( .A(n21843), .B(n21842), .Z(n22151) );
  NANDN U22364 ( .A(n210), .B(n21844), .Z(n21846) );
  XOR U22365 ( .A(a[98]), .B(b[9]), .Z(n22113) );
  NANDN U22366 ( .A(n30267), .B(n22113), .Z(n21845) );
  AND U22367 ( .A(n21846), .B(n21845), .Z(n22150) );
  NANDN U22368 ( .A(n212), .B(n21847), .Z(n21849) );
  XOR U22369 ( .A(b[49]), .B(a[58]), .Z(n22116) );
  NANDN U22370 ( .A(n37432), .B(n22116), .Z(n21848) );
  NAND U22371 ( .A(n21849), .B(n21848), .Z(n22149) );
  XOR U22372 ( .A(n22150), .B(n22149), .Z(n22152) );
  XOR U22373 ( .A(n22151), .B(n22152), .Z(n22264) );
  NANDN U22374 ( .A(n36742), .B(n21850), .Z(n21852) );
  XOR U22375 ( .A(b[43]), .B(a[64]), .Z(n22119) );
  NANDN U22376 ( .A(n36891), .B(n22119), .Z(n21851) );
  AND U22377 ( .A(n21852), .B(n21851), .Z(n22130) );
  NANDN U22378 ( .A(n36991), .B(n21853), .Z(n21855) );
  XOR U22379 ( .A(b[45]), .B(a[62]), .Z(n22122) );
  NANDN U22380 ( .A(n37083), .B(n22122), .Z(n21854) );
  AND U22381 ( .A(n21855), .B(n21854), .Z(n22129) );
  NANDN U22382 ( .A(n30482), .B(n21856), .Z(n21858) );
  XOR U22383 ( .A(a[96]), .B(b[11]), .Z(n22125) );
  NANDN U22384 ( .A(n30891), .B(n22125), .Z(n21857) );
  NAND U22385 ( .A(n21858), .B(n21857), .Z(n22128) );
  XOR U22386 ( .A(n22129), .B(n22128), .Z(n22131) );
  XNOR U22387 ( .A(n22130), .B(n22131), .Z(n22263) );
  XNOR U22388 ( .A(n22264), .B(n22263), .Z(n22265) );
  NANDN U22389 ( .A(n21860), .B(n21859), .Z(n21864) );
  OR U22390 ( .A(n21862), .B(n21861), .Z(n21863) );
  NAND U22391 ( .A(n21864), .B(n21863), .Z(n22266) );
  XNOR U22392 ( .A(n22265), .B(n22266), .Z(n22074) );
  XNOR U22393 ( .A(n22075), .B(n22074), .Z(n22076) );
  NANDN U22394 ( .A(n29499), .B(n21865), .Z(n21867) );
  XOR U22395 ( .A(a[100]), .B(b[7]), .Z(n22134) );
  NANDN U22396 ( .A(n29735), .B(n22134), .Z(n21866) );
  AND U22397 ( .A(n21867), .B(n21866), .Z(n22193) );
  NANDN U22398 ( .A(n37857), .B(n21868), .Z(n21870) );
  XOR U22399 ( .A(b[55]), .B(a[52]), .Z(n22137) );
  NANDN U22400 ( .A(n37911), .B(n22137), .Z(n21869) );
  AND U22401 ( .A(n21870), .B(n21869), .Z(n22192) );
  NANDN U22402 ( .A(n35611), .B(n21871), .Z(n21873) );
  XOR U22403 ( .A(b[35]), .B(a[72]), .Z(n22140) );
  NANDN U22404 ( .A(n35801), .B(n22140), .Z(n21872) );
  NAND U22405 ( .A(n21873), .B(n21872), .Z(n22191) );
  XOR U22406 ( .A(n22192), .B(n22191), .Z(n22194) );
  XOR U22407 ( .A(n22193), .B(n22194), .Z(n22204) );
  NANDN U22408 ( .A(n21875), .B(n21874), .Z(n21879) );
  OR U22409 ( .A(n21877), .B(n21876), .Z(n21878) );
  AND U22410 ( .A(n21879), .B(n21878), .Z(n22203) );
  XNOR U22411 ( .A(n22204), .B(n22203), .Z(n22205) );
  NANDN U22412 ( .A(n21881), .B(n21880), .Z(n21885) );
  OR U22413 ( .A(n21883), .B(n21882), .Z(n21884) );
  NAND U22414 ( .A(n21885), .B(n21884), .Z(n22206) );
  XOR U22415 ( .A(n22205), .B(n22206), .Z(n22077) );
  XNOR U22416 ( .A(n22076), .B(n22077), .Z(n22086) );
  XOR U22417 ( .A(n22087), .B(n22086), .Z(n22089) );
  XOR U22418 ( .A(n22088), .B(n22089), .Z(n22057) );
  NANDN U22419 ( .A(n21887), .B(n21886), .Z(n21891) );
  NANDN U22420 ( .A(n21889), .B(n21888), .Z(n21890) );
  AND U22421 ( .A(n21891), .B(n21890), .Z(n22070) );
  NANDN U22422 ( .A(n21893), .B(n21892), .Z(n21897) );
  NANDN U22423 ( .A(n21895), .B(n21894), .Z(n21896) );
  AND U22424 ( .A(n21897), .B(n21896), .Z(n22069) );
  NANDN U22425 ( .A(n21899), .B(n21898), .Z(n21903) );
  NAND U22426 ( .A(n21901), .B(n21900), .Z(n21902) );
  AND U22427 ( .A(n21903), .B(n21902), .Z(n22068) );
  XOR U22428 ( .A(n22069), .B(n22068), .Z(n22071) );
  XOR U22429 ( .A(n22070), .B(n22071), .Z(n22095) );
  NANDN U22430 ( .A(n21905), .B(n21904), .Z(n21909) );
  NANDN U22431 ( .A(n21907), .B(n21906), .Z(n21908) );
  AND U22432 ( .A(n21909), .B(n21908), .Z(n22216) );
  NANDN U22433 ( .A(n21911), .B(n21910), .Z(n21915) );
  OR U22434 ( .A(n21913), .B(n21912), .Z(n21914) );
  NAND U22435 ( .A(n21915), .B(n21914), .Z(n22215) );
  XNOR U22436 ( .A(n22216), .B(n22215), .Z(n22218) );
  NANDN U22437 ( .A(n21917), .B(n21916), .Z(n21921) );
  OR U22438 ( .A(n21919), .B(n21918), .Z(n21920) );
  AND U22439 ( .A(n21921), .B(n21920), .Z(n22164) );
  NAND U22440 ( .A(b[0]), .B(a[106]), .Z(n21922) );
  XNOR U22441 ( .A(b[1]), .B(n21922), .Z(n21924) );
  NANDN U22442 ( .A(b[0]), .B(a[105]), .Z(n21923) );
  NAND U22443 ( .A(n21924), .B(n21923), .Z(n22200) );
  NANDN U22444 ( .A(n38278), .B(n21925), .Z(n21927) );
  XOR U22445 ( .A(b[63]), .B(a[44]), .Z(n22242) );
  NANDN U22446 ( .A(n38279), .B(n22242), .Z(n21926) );
  AND U22447 ( .A(n21927), .B(n21926), .Z(n22198) );
  NANDN U22448 ( .A(n35260), .B(n21928), .Z(n21930) );
  XOR U22449 ( .A(b[33]), .B(a[74]), .Z(n22245) );
  NANDN U22450 ( .A(n35456), .B(n22245), .Z(n21929) );
  NAND U22451 ( .A(n21930), .B(n21929), .Z(n22197) );
  XNOR U22452 ( .A(n22198), .B(n22197), .Z(n22199) );
  XNOR U22453 ( .A(n22200), .B(n22199), .Z(n22161) );
  NANDN U22454 ( .A(n37974), .B(n21931), .Z(n21933) );
  XOR U22455 ( .A(b[57]), .B(a[50]), .Z(n22248) );
  NANDN U22456 ( .A(n38031), .B(n22248), .Z(n21932) );
  AND U22457 ( .A(n21933), .B(n21932), .Z(n22224) );
  NANDN U22458 ( .A(n38090), .B(n21934), .Z(n21936) );
  XOR U22459 ( .A(b[59]), .B(a[48]), .Z(n22251) );
  NANDN U22460 ( .A(n38130), .B(n22251), .Z(n21935) );
  AND U22461 ( .A(n21936), .B(n21935), .Z(n22222) );
  NANDN U22462 ( .A(n36480), .B(n21937), .Z(n21939) );
  XOR U22463 ( .A(b[41]), .B(a[66]), .Z(n22254) );
  NANDN U22464 ( .A(n36594), .B(n22254), .Z(n21938) );
  NAND U22465 ( .A(n21939), .B(n21938), .Z(n22221) );
  XNOR U22466 ( .A(n22222), .B(n22221), .Z(n22223) );
  XOR U22467 ( .A(n22224), .B(n22223), .Z(n22162) );
  XNOR U22468 ( .A(n22161), .B(n22162), .Z(n22163) );
  XNOR U22469 ( .A(n22164), .B(n22163), .Z(n22217) );
  XOR U22470 ( .A(n22218), .B(n22217), .Z(n22099) );
  NANDN U22471 ( .A(n21941), .B(n21940), .Z(n21945) );
  NAND U22472 ( .A(n21943), .B(n21942), .Z(n21944) );
  NAND U22473 ( .A(n21945), .B(n21944), .Z(n22098) );
  XNOR U22474 ( .A(n22099), .B(n22098), .Z(n22101) );
  NANDN U22475 ( .A(n21947), .B(n21946), .Z(n21951) );
  NANDN U22476 ( .A(n21949), .B(n21948), .Z(n21950) );
  AND U22477 ( .A(n21951), .B(n21950), .Z(n22317) );
  NANDN U22478 ( .A(n32996), .B(n21952), .Z(n21954) );
  XOR U22479 ( .A(a[86]), .B(b[21]), .Z(n22269) );
  NANDN U22480 ( .A(n33271), .B(n22269), .Z(n21953) );
  AND U22481 ( .A(n21954), .B(n21953), .Z(n22235) );
  NANDN U22482 ( .A(n33866), .B(n21955), .Z(n21957) );
  XOR U22483 ( .A(b[23]), .B(a[84]), .Z(n22272) );
  NANDN U22484 ( .A(n33644), .B(n22272), .Z(n21956) );
  AND U22485 ( .A(n21957), .B(n21956), .Z(n22234) );
  NANDN U22486 ( .A(n32483), .B(n21958), .Z(n21960) );
  XOR U22487 ( .A(a[88]), .B(b[19]), .Z(n22275) );
  NANDN U22488 ( .A(n32823), .B(n22275), .Z(n21959) );
  NAND U22489 ( .A(n21960), .B(n21959), .Z(n22233) );
  XOR U22490 ( .A(n22234), .B(n22233), .Z(n22236) );
  XOR U22491 ( .A(n22235), .B(n22236), .Z(n22105) );
  NANDN U22492 ( .A(n34909), .B(n21961), .Z(n21963) );
  XOR U22493 ( .A(b[31]), .B(a[76]), .Z(n22278) );
  NANDN U22494 ( .A(n35145), .B(n22278), .Z(n21962) );
  AND U22495 ( .A(n21963), .B(n21962), .Z(n22145) );
  NANDN U22496 ( .A(n38247), .B(n21964), .Z(n21966) );
  XOR U22497 ( .A(b[61]), .B(a[46]), .Z(n22281) );
  NANDN U22498 ( .A(n38248), .B(n22281), .Z(n21965) );
  AND U22499 ( .A(n21966), .B(n21965), .Z(n22144) );
  AND U22500 ( .A(b[63]), .B(a[42]), .Z(n22143) );
  XOR U22501 ( .A(n22144), .B(n22143), .Z(n22146) );
  XNOR U22502 ( .A(n22145), .B(n22146), .Z(n22104) );
  XNOR U22503 ( .A(n22105), .B(n22104), .Z(n22106) );
  NANDN U22504 ( .A(n21968), .B(n21967), .Z(n21972) );
  OR U22505 ( .A(n21970), .B(n21969), .Z(n21971) );
  NAND U22506 ( .A(n21972), .B(n21971), .Z(n22107) );
  XNOR U22507 ( .A(n22106), .B(n22107), .Z(n22314) );
  NANDN U22508 ( .A(n34223), .B(n21973), .Z(n21975) );
  XOR U22509 ( .A(b[27]), .B(a[80]), .Z(n22290) );
  NANDN U22510 ( .A(n34458), .B(n22290), .Z(n21974) );
  AND U22511 ( .A(n21975), .B(n21974), .Z(n22187) );
  NANDN U22512 ( .A(n34634), .B(n21976), .Z(n21978) );
  XOR U22513 ( .A(b[29]), .B(a[78]), .Z(n22293) );
  NANDN U22514 ( .A(n34722), .B(n22293), .Z(n21977) );
  AND U22515 ( .A(n21978), .B(n21977), .Z(n22186) );
  NANDN U22516 ( .A(n31055), .B(n21979), .Z(n21981) );
  XOR U22517 ( .A(a[94]), .B(b[13]), .Z(n22296) );
  NANDN U22518 ( .A(n31293), .B(n22296), .Z(n21980) );
  NAND U22519 ( .A(n21981), .B(n21980), .Z(n22185) );
  XOR U22520 ( .A(n22186), .B(n22185), .Z(n22188) );
  XOR U22521 ( .A(n22187), .B(n22188), .Z(n22210) );
  NANDN U22522 ( .A(n28889), .B(n21982), .Z(n21984) );
  XOR U22523 ( .A(a[102]), .B(b[5]), .Z(n22299) );
  NANDN U22524 ( .A(n29138), .B(n22299), .Z(n21983) );
  AND U22525 ( .A(n21984), .B(n21983), .Z(n22229) );
  NANDN U22526 ( .A(n209), .B(n21985), .Z(n21987) );
  XOR U22527 ( .A(a[104]), .B(b[3]), .Z(n22302) );
  NANDN U22528 ( .A(n28941), .B(n22302), .Z(n21986) );
  AND U22529 ( .A(n21987), .B(n21986), .Z(n22228) );
  NANDN U22530 ( .A(n35936), .B(n21988), .Z(n21990) );
  XOR U22531 ( .A(b[37]), .B(a[70]), .Z(n22305) );
  NANDN U22532 ( .A(n36047), .B(n22305), .Z(n21989) );
  NAND U22533 ( .A(n21990), .B(n21989), .Z(n22227) );
  XOR U22534 ( .A(n22228), .B(n22227), .Z(n22230) );
  XNOR U22535 ( .A(n22229), .B(n22230), .Z(n22209) );
  XNOR U22536 ( .A(n22210), .B(n22209), .Z(n22211) );
  NANDN U22537 ( .A(n21992), .B(n21991), .Z(n21996) );
  OR U22538 ( .A(n21994), .B(n21993), .Z(n21995) );
  NAND U22539 ( .A(n21996), .B(n21995), .Z(n22212) );
  XOR U22540 ( .A(n22211), .B(n22212), .Z(n22315) );
  XNOR U22541 ( .A(n22314), .B(n22315), .Z(n22316) );
  XNOR U22542 ( .A(n22317), .B(n22316), .Z(n22100) );
  XOR U22543 ( .A(n22101), .B(n22100), .Z(n22093) );
  NANDN U22544 ( .A(n21998), .B(n21997), .Z(n22002) );
  NANDN U22545 ( .A(n22000), .B(n21999), .Z(n22001) );
  AND U22546 ( .A(n22002), .B(n22001), .Z(n22092) );
  XNOR U22547 ( .A(n22093), .B(n22092), .Z(n22094) );
  XNOR U22548 ( .A(n22095), .B(n22094), .Z(n22056) );
  XOR U22549 ( .A(n22057), .B(n22056), .Z(n22059) );
  XOR U22550 ( .A(n22058), .B(n22059), .Z(n22322) );
  NAND U22551 ( .A(n22004), .B(n22003), .Z(n22008) );
  NAND U22552 ( .A(n22006), .B(n22005), .Z(n22007) );
  AND U22553 ( .A(n22008), .B(n22007), .Z(n22065) );
  NANDN U22554 ( .A(n22010), .B(n22009), .Z(n22014) );
  OR U22555 ( .A(n22012), .B(n22011), .Z(n22013) );
  AND U22556 ( .A(n22014), .B(n22013), .Z(n22063) );
  NANDN U22557 ( .A(n22016), .B(n22015), .Z(n22020) );
  NANDN U22558 ( .A(n22018), .B(n22017), .Z(n22019) );
  AND U22559 ( .A(n22020), .B(n22019), .Z(n22062) );
  XNOR U22560 ( .A(n22063), .B(n22062), .Z(n22064) );
  XOR U22561 ( .A(n22065), .B(n22064), .Z(n22321) );
  NANDN U22562 ( .A(n22022), .B(n22021), .Z(n22026) );
  OR U22563 ( .A(n22024), .B(n22023), .Z(n22025) );
  NAND U22564 ( .A(n22026), .B(n22025), .Z(n22320) );
  XOR U22565 ( .A(n22321), .B(n22320), .Z(n22323) );
  XOR U22566 ( .A(n22322), .B(n22323), .Z(n22329) );
  NANDN U22567 ( .A(n22028), .B(n22027), .Z(n22032) );
  NANDN U22568 ( .A(n22030), .B(n22029), .Z(n22031) );
  AND U22569 ( .A(n22032), .B(n22031), .Z(n22327) );
  NANDN U22570 ( .A(n22034), .B(n22033), .Z(n22038) );
  OR U22571 ( .A(n22036), .B(n22035), .Z(n22037) );
  AND U22572 ( .A(n22038), .B(n22037), .Z(n22326) );
  XNOR U22573 ( .A(n22327), .B(n22326), .Z(n22328) );
  XNOR U22574 ( .A(n22329), .B(n22328), .Z(n22050) );
  XOR U22575 ( .A(n22051), .B(n22050), .Z(n22053) );
  XNOR U22576 ( .A(n22052), .B(n22053), .Z(n22044) );
  XNOR U22577 ( .A(n22045), .B(n22044), .Z(n22046) );
  XNOR U22578 ( .A(n22047), .B(n22046), .Z(n22332) );
  XNOR U22579 ( .A(sreg[170]), .B(n22332), .Z(n22334) );
  NANDN U22580 ( .A(sreg[169]), .B(n22039), .Z(n22043) );
  NAND U22581 ( .A(n22041), .B(n22040), .Z(n22042) );
  NAND U22582 ( .A(n22043), .B(n22042), .Z(n22333) );
  XNOR U22583 ( .A(n22334), .B(n22333), .Z(c[170]) );
  NANDN U22584 ( .A(n22045), .B(n22044), .Z(n22049) );
  NANDN U22585 ( .A(n22047), .B(n22046), .Z(n22048) );
  AND U22586 ( .A(n22049), .B(n22048), .Z(n22340) );
  NANDN U22587 ( .A(n22051), .B(n22050), .Z(n22055) );
  OR U22588 ( .A(n22053), .B(n22052), .Z(n22054) );
  AND U22589 ( .A(n22055), .B(n22054), .Z(n22337) );
  NANDN U22590 ( .A(n22057), .B(n22056), .Z(n22061) );
  OR U22591 ( .A(n22059), .B(n22058), .Z(n22060) );
  AND U22592 ( .A(n22061), .B(n22060), .Z(n22620) );
  NANDN U22593 ( .A(n22063), .B(n22062), .Z(n22067) );
  NAND U22594 ( .A(n22065), .B(n22064), .Z(n22066) );
  NAND U22595 ( .A(n22067), .B(n22066), .Z(n22619) );
  XNOR U22596 ( .A(n22620), .B(n22619), .Z(n22622) );
  NANDN U22597 ( .A(n22069), .B(n22068), .Z(n22073) );
  OR U22598 ( .A(n22071), .B(n22070), .Z(n22072) );
  AND U22599 ( .A(n22073), .B(n22072), .Z(n22357) );
  NANDN U22600 ( .A(n22075), .B(n22074), .Z(n22079) );
  NANDN U22601 ( .A(n22077), .B(n22076), .Z(n22078) );
  AND U22602 ( .A(n22079), .B(n22078), .Z(n22356) );
  NANDN U22603 ( .A(n22081), .B(n22080), .Z(n22085) );
  OR U22604 ( .A(n22083), .B(n22082), .Z(n22084) );
  AND U22605 ( .A(n22085), .B(n22084), .Z(n22355) );
  XOR U22606 ( .A(n22356), .B(n22355), .Z(n22358) );
  XOR U22607 ( .A(n22357), .B(n22358), .Z(n22614) );
  NANDN U22608 ( .A(n22087), .B(n22086), .Z(n22091) );
  OR U22609 ( .A(n22089), .B(n22088), .Z(n22090) );
  AND U22610 ( .A(n22091), .B(n22090), .Z(n22613) );
  XNOR U22611 ( .A(n22614), .B(n22613), .Z(n22615) );
  NANDN U22612 ( .A(n22093), .B(n22092), .Z(n22097) );
  NANDN U22613 ( .A(n22095), .B(n22094), .Z(n22096) );
  AND U22614 ( .A(n22097), .B(n22096), .Z(n22352) );
  NANDN U22615 ( .A(n22099), .B(n22098), .Z(n22103) );
  NAND U22616 ( .A(n22101), .B(n22100), .Z(n22102) );
  AND U22617 ( .A(n22103), .B(n22102), .Z(n22381) );
  NANDN U22618 ( .A(n22105), .B(n22104), .Z(n22109) );
  NANDN U22619 ( .A(n22107), .B(n22106), .Z(n22108) );
  AND U22620 ( .A(n22109), .B(n22108), .Z(n22368) );
  NAND U22621 ( .A(n37294), .B(n22110), .Z(n22112) );
  XNOR U22622 ( .A(b[47]), .B(a[61]), .Z(n22451) );
  NANDN U22623 ( .A(n22451), .B(n37341), .Z(n22111) );
  NAND U22624 ( .A(n22112), .B(n22111), .Z(n22492) );
  NAND U22625 ( .A(n30627), .B(n22113), .Z(n22115) );
  XNOR U22626 ( .A(a[99]), .B(b[9]), .Z(n22454) );
  NANDN U22627 ( .A(n22454), .B(n30628), .Z(n22114) );
  NAND U22628 ( .A(n22115), .B(n22114), .Z(n22491) );
  NAND U22629 ( .A(n37536), .B(n22116), .Z(n22118) );
  XNOR U22630 ( .A(b[49]), .B(a[59]), .Z(n22457) );
  NANDN U22631 ( .A(n22457), .B(n37537), .Z(n22117) );
  NAND U22632 ( .A(n22118), .B(n22117), .Z(n22490) );
  XNOR U22633 ( .A(n22491), .B(n22490), .Z(n22493) );
  NANDN U22634 ( .A(n36742), .B(n22119), .Z(n22121) );
  XOR U22635 ( .A(b[43]), .B(a[65]), .Z(n22460) );
  NANDN U22636 ( .A(n36891), .B(n22460), .Z(n22120) );
  AND U22637 ( .A(n22121), .B(n22120), .Z(n22471) );
  NANDN U22638 ( .A(n36991), .B(n22122), .Z(n22124) );
  XOR U22639 ( .A(b[45]), .B(a[63]), .Z(n22463) );
  NANDN U22640 ( .A(n37083), .B(n22463), .Z(n22123) );
  AND U22641 ( .A(n22124), .B(n22123), .Z(n22470) );
  NANDN U22642 ( .A(n30482), .B(n22125), .Z(n22127) );
  XOR U22643 ( .A(a[97]), .B(b[11]), .Z(n22466) );
  NANDN U22644 ( .A(n30891), .B(n22466), .Z(n22126) );
  NAND U22645 ( .A(n22127), .B(n22126), .Z(n22469) );
  XOR U22646 ( .A(n22470), .B(n22469), .Z(n22472) );
  XNOR U22647 ( .A(n22471), .B(n22472), .Z(n22514) );
  XOR U22648 ( .A(n22515), .B(n22514), .Z(n22516) );
  NANDN U22649 ( .A(n22129), .B(n22128), .Z(n22133) );
  OR U22650 ( .A(n22131), .B(n22130), .Z(n22132) );
  NAND U22651 ( .A(n22133), .B(n22132), .Z(n22517) );
  XNOR U22652 ( .A(n22516), .B(n22517), .Z(n22367) );
  XNOR U22653 ( .A(n22368), .B(n22367), .Z(n22370) );
  NANDN U22654 ( .A(n29499), .B(n22134), .Z(n22136) );
  XOR U22655 ( .A(a[101]), .B(b[7]), .Z(n22475) );
  NANDN U22656 ( .A(n29735), .B(n22475), .Z(n22135) );
  AND U22657 ( .A(n22136), .B(n22135), .Z(n22435) );
  NANDN U22658 ( .A(n37857), .B(n22137), .Z(n22139) );
  XOR U22659 ( .A(b[55]), .B(a[53]), .Z(n22478) );
  NANDN U22660 ( .A(n37911), .B(n22478), .Z(n22138) );
  AND U22661 ( .A(n22139), .B(n22138), .Z(n22434) );
  NANDN U22662 ( .A(n35611), .B(n22140), .Z(n22142) );
  XOR U22663 ( .A(b[35]), .B(a[73]), .Z(n22481) );
  NANDN U22664 ( .A(n35801), .B(n22481), .Z(n22141) );
  NAND U22665 ( .A(n22142), .B(n22141), .Z(n22433) );
  XOR U22666 ( .A(n22434), .B(n22433), .Z(n22436) );
  XOR U22667 ( .A(n22435), .B(n22436), .Z(n22497) );
  NANDN U22668 ( .A(n22144), .B(n22143), .Z(n22148) );
  OR U22669 ( .A(n22146), .B(n22145), .Z(n22147) );
  AND U22670 ( .A(n22148), .B(n22147), .Z(n22496) );
  XNOR U22671 ( .A(n22497), .B(n22496), .Z(n22498) );
  NANDN U22672 ( .A(n22150), .B(n22149), .Z(n22154) );
  OR U22673 ( .A(n22152), .B(n22151), .Z(n22153) );
  NAND U22674 ( .A(n22154), .B(n22153), .Z(n22499) );
  XNOR U22675 ( .A(n22498), .B(n22499), .Z(n22369) );
  XOR U22676 ( .A(n22370), .B(n22369), .Z(n22380) );
  NANDN U22677 ( .A(n22156), .B(n22155), .Z(n22160) );
  NANDN U22678 ( .A(n22158), .B(n22157), .Z(n22159) );
  AND U22679 ( .A(n22160), .B(n22159), .Z(n22376) );
  NANDN U22680 ( .A(n22162), .B(n22161), .Z(n22166) );
  NANDN U22681 ( .A(n22164), .B(n22163), .Z(n22165) );
  AND U22682 ( .A(n22166), .B(n22165), .Z(n22374) );
  NANDN U22683 ( .A(n33875), .B(n22167), .Z(n22169) );
  XOR U22684 ( .A(b[25]), .B(a[83]), .Z(n22409) );
  NANDN U22685 ( .A(n33994), .B(n22409), .Z(n22168) );
  AND U22686 ( .A(n22169), .B(n22168), .Z(n22546) );
  NANDN U22687 ( .A(n32013), .B(n22170), .Z(n22172) );
  XOR U22688 ( .A(a[91]), .B(b[17]), .Z(n22412) );
  NANDN U22689 ( .A(n32292), .B(n22412), .Z(n22171) );
  AND U22690 ( .A(n22172), .B(n22171), .Z(n22545) );
  NANDN U22691 ( .A(n31536), .B(n22173), .Z(n22175) );
  XOR U22692 ( .A(a[93]), .B(b[15]), .Z(n22415) );
  NANDN U22693 ( .A(n31925), .B(n22415), .Z(n22174) );
  NAND U22694 ( .A(n22175), .B(n22174), .Z(n22544) );
  XOR U22695 ( .A(n22545), .B(n22544), .Z(n22547) );
  XOR U22696 ( .A(n22546), .B(n22547), .Z(n22602) );
  NANDN U22697 ( .A(n37526), .B(n22176), .Z(n22178) );
  XOR U22698 ( .A(b[51]), .B(a[57]), .Z(n22418) );
  NANDN U22699 ( .A(n37605), .B(n22418), .Z(n22177) );
  AND U22700 ( .A(n22178), .B(n22177), .Z(n22522) );
  NANDN U22701 ( .A(n37705), .B(n22179), .Z(n22181) );
  XOR U22702 ( .A(b[53]), .B(a[55]), .Z(n22421) );
  NANDN U22703 ( .A(n37778), .B(n22421), .Z(n22180) );
  AND U22704 ( .A(n22181), .B(n22180), .Z(n22521) );
  NANDN U22705 ( .A(n36210), .B(n22182), .Z(n22184) );
  XOR U22706 ( .A(b[39]), .B(a[69]), .Z(n22424) );
  NANDN U22707 ( .A(n36347), .B(n22424), .Z(n22183) );
  NAND U22708 ( .A(n22184), .B(n22183), .Z(n22520) );
  XOR U22709 ( .A(n22521), .B(n22520), .Z(n22523) );
  XNOR U22710 ( .A(n22522), .B(n22523), .Z(n22601) );
  XNOR U22711 ( .A(n22602), .B(n22601), .Z(n22604) );
  NANDN U22712 ( .A(n22186), .B(n22185), .Z(n22190) );
  OR U22713 ( .A(n22188), .B(n22187), .Z(n22189) );
  AND U22714 ( .A(n22190), .B(n22189), .Z(n22603) );
  XOR U22715 ( .A(n22604), .B(n22603), .Z(n22400) );
  NANDN U22716 ( .A(n22192), .B(n22191), .Z(n22196) );
  OR U22717 ( .A(n22194), .B(n22193), .Z(n22195) );
  AND U22718 ( .A(n22196), .B(n22195), .Z(n22398) );
  NANDN U22719 ( .A(n22198), .B(n22197), .Z(n22202) );
  NANDN U22720 ( .A(n22200), .B(n22199), .Z(n22201) );
  NAND U22721 ( .A(n22202), .B(n22201), .Z(n22397) );
  XNOR U22722 ( .A(n22398), .B(n22397), .Z(n22399) );
  XNOR U22723 ( .A(n22400), .B(n22399), .Z(n22373) );
  XNOR U22724 ( .A(n22374), .B(n22373), .Z(n22375) );
  XNOR U22725 ( .A(n22376), .B(n22375), .Z(n22379) );
  XOR U22726 ( .A(n22380), .B(n22379), .Z(n22382) );
  XNOR U22727 ( .A(n22381), .B(n22382), .Z(n22349) );
  NANDN U22728 ( .A(n22204), .B(n22203), .Z(n22208) );
  NANDN U22729 ( .A(n22206), .B(n22205), .Z(n22207) );
  AND U22730 ( .A(n22208), .B(n22207), .Z(n22363) );
  NANDN U22731 ( .A(n22210), .B(n22209), .Z(n22214) );
  NANDN U22732 ( .A(n22212), .B(n22211), .Z(n22213) );
  AND U22733 ( .A(n22214), .B(n22213), .Z(n22362) );
  NANDN U22734 ( .A(n22216), .B(n22215), .Z(n22220) );
  NAND U22735 ( .A(n22218), .B(n22217), .Z(n22219) );
  AND U22736 ( .A(n22220), .B(n22219), .Z(n22361) );
  XOR U22737 ( .A(n22362), .B(n22361), .Z(n22364) );
  XOR U22738 ( .A(n22363), .B(n22364), .Z(n22388) );
  NANDN U22739 ( .A(n22222), .B(n22221), .Z(n22226) );
  NANDN U22740 ( .A(n22224), .B(n22223), .Z(n22225) );
  AND U22741 ( .A(n22226), .B(n22225), .Z(n22509) );
  NANDN U22742 ( .A(n22228), .B(n22227), .Z(n22232) );
  OR U22743 ( .A(n22230), .B(n22229), .Z(n22231) );
  NAND U22744 ( .A(n22232), .B(n22231), .Z(n22508) );
  XNOR U22745 ( .A(n22509), .B(n22508), .Z(n22511) );
  NANDN U22746 ( .A(n22234), .B(n22233), .Z(n22238) );
  OR U22747 ( .A(n22236), .B(n22235), .Z(n22237) );
  AND U22748 ( .A(n22238), .B(n22237), .Z(n22406) );
  NAND U22749 ( .A(b[0]), .B(a[107]), .Z(n22239) );
  XNOR U22750 ( .A(b[1]), .B(n22239), .Z(n22241) );
  NANDN U22751 ( .A(b[0]), .B(a[106]), .Z(n22240) );
  NAND U22752 ( .A(n22241), .B(n22240), .Z(n22442) );
  NANDN U22753 ( .A(n38278), .B(n22242), .Z(n22244) );
  XOR U22754 ( .A(b[63]), .B(a[45]), .Z(n22583) );
  NANDN U22755 ( .A(n38279), .B(n22583), .Z(n22243) );
  AND U22756 ( .A(n22244), .B(n22243), .Z(n22440) );
  NANDN U22757 ( .A(n35260), .B(n22245), .Z(n22247) );
  XOR U22758 ( .A(b[33]), .B(a[75]), .Z(n22586) );
  NANDN U22759 ( .A(n35456), .B(n22586), .Z(n22246) );
  NAND U22760 ( .A(n22247), .B(n22246), .Z(n22439) );
  XNOR U22761 ( .A(n22440), .B(n22439), .Z(n22441) );
  XNOR U22762 ( .A(n22442), .B(n22441), .Z(n22403) );
  NANDN U22763 ( .A(n37974), .B(n22248), .Z(n22250) );
  XOR U22764 ( .A(b[57]), .B(a[51]), .Z(n22592) );
  NANDN U22765 ( .A(n38031), .B(n22592), .Z(n22249) );
  AND U22766 ( .A(n22250), .B(n22249), .Z(n22568) );
  NANDN U22767 ( .A(n38090), .B(n22251), .Z(n22253) );
  XOR U22768 ( .A(b[59]), .B(a[49]), .Z(n22595) );
  NANDN U22769 ( .A(n38130), .B(n22595), .Z(n22252) );
  AND U22770 ( .A(n22253), .B(n22252), .Z(n22566) );
  NANDN U22771 ( .A(n36480), .B(n22254), .Z(n22256) );
  XOR U22772 ( .A(b[41]), .B(a[67]), .Z(n22598) );
  NANDN U22773 ( .A(n36594), .B(n22598), .Z(n22255) );
  NAND U22774 ( .A(n22256), .B(n22255), .Z(n22565) );
  XNOR U22775 ( .A(n22566), .B(n22565), .Z(n22567) );
  XOR U22776 ( .A(n22568), .B(n22567), .Z(n22404) );
  XNOR U22777 ( .A(n22403), .B(n22404), .Z(n22405) );
  XNOR U22778 ( .A(n22406), .B(n22405), .Z(n22510) );
  XOR U22779 ( .A(n22511), .B(n22510), .Z(n22392) );
  NANDN U22780 ( .A(n22258), .B(n22257), .Z(n22262) );
  NAND U22781 ( .A(n22260), .B(n22259), .Z(n22261) );
  NAND U22782 ( .A(n22262), .B(n22261), .Z(n22391) );
  XNOR U22783 ( .A(n22392), .B(n22391), .Z(n22394) );
  NANDN U22784 ( .A(n22264), .B(n22263), .Z(n22268) );
  NANDN U22785 ( .A(n22266), .B(n22265), .Z(n22267) );
  AND U22786 ( .A(n22268), .B(n22267), .Z(n22610) );
  NANDN U22787 ( .A(n32996), .B(n22269), .Z(n22271) );
  XOR U22788 ( .A(b[21]), .B(a[87]), .Z(n22550) );
  NANDN U22789 ( .A(n33271), .B(n22550), .Z(n22270) );
  AND U22790 ( .A(n22271), .B(n22270), .Z(n22579) );
  NANDN U22791 ( .A(n33866), .B(n22272), .Z(n22274) );
  XOR U22792 ( .A(b[23]), .B(a[85]), .Z(n22553) );
  NANDN U22793 ( .A(n33644), .B(n22553), .Z(n22273) );
  AND U22794 ( .A(n22274), .B(n22273), .Z(n22578) );
  NANDN U22795 ( .A(n32483), .B(n22275), .Z(n22277) );
  XOR U22796 ( .A(a[89]), .B(b[19]), .Z(n22556) );
  NANDN U22797 ( .A(n32823), .B(n22556), .Z(n22276) );
  NAND U22798 ( .A(n22277), .B(n22276), .Z(n22577) );
  XOR U22799 ( .A(n22578), .B(n22577), .Z(n22580) );
  XOR U22800 ( .A(n22579), .B(n22580), .Z(n22446) );
  NANDN U22801 ( .A(n34909), .B(n22278), .Z(n22280) );
  XOR U22802 ( .A(b[31]), .B(a[77]), .Z(n22559) );
  NANDN U22803 ( .A(n35145), .B(n22559), .Z(n22279) );
  AND U22804 ( .A(n22280), .B(n22279), .Z(n22486) );
  NANDN U22805 ( .A(n38247), .B(n22281), .Z(n22283) );
  XOR U22806 ( .A(b[61]), .B(a[47]), .Z(n22562) );
  NANDN U22807 ( .A(n38248), .B(n22562), .Z(n22282) );
  AND U22808 ( .A(n22283), .B(n22282), .Z(n22485) );
  AND U22809 ( .A(b[63]), .B(a[43]), .Z(n22484) );
  XOR U22810 ( .A(n22485), .B(n22484), .Z(n22487) );
  XNOR U22811 ( .A(n22486), .B(n22487), .Z(n22445) );
  XNOR U22812 ( .A(n22446), .B(n22445), .Z(n22447) );
  NANDN U22813 ( .A(n22285), .B(n22284), .Z(n22289) );
  OR U22814 ( .A(n22287), .B(n22286), .Z(n22288) );
  NAND U22815 ( .A(n22289), .B(n22288), .Z(n22448) );
  XNOR U22816 ( .A(n22447), .B(n22448), .Z(n22607) );
  NANDN U22817 ( .A(n34223), .B(n22290), .Z(n22292) );
  XOR U22818 ( .A(b[27]), .B(a[81]), .Z(n22526) );
  NANDN U22819 ( .A(n34458), .B(n22526), .Z(n22291) );
  AND U22820 ( .A(n22292), .B(n22291), .Z(n22429) );
  NANDN U22821 ( .A(n34634), .B(n22293), .Z(n22295) );
  XOR U22822 ( .A(b[29]), .B(a[79]), .Z(n22529) );
  NANDN U22823 ( .A(n34722), .B(n22529), .Z(n22294) );
  AND U22824 ( .A(n22295), .B(n22294), .Z(n22428) );
  NANDN U22825 ( .A(n31055), .B(n22296), .Z(n22298) );
  XOR U22826 ( .A(a[95]), .B(b[13]), .Z(n22532) );
  NANDN U22827 ( .A(n31293), .B(n22532), .Z(n22297) );
  NAND U22828 ( .A(n22298), .B(n22297), .Z(n22427) );
  XOR U22829 ( .A(n22428), .B(n22427), .Z(n22430) );
  XOR U22830 ( .A(n22429), .B(n22430), .Z(n22503) );
  NANDN U22831 ( .A(n28889), .B(n22299), .Z(n22301) );
  XOR U22832 ( .A(a[103]), .B(b[5]), .Z(n22535) );
  NANDN U22833 ( .A(n29138), .B(n22535), .Z(n22300) );
  AND U22834 ( .A(n22301), .B(n22300), .Z(n22573) );
  NANDN U22835 ( .A(n209), .B(n22302), .Z(n22304) );
  XOR U22836 ( .A(a[105]), .B(b[3]), .Z(n22538) );
  NANDN U22837 ( .A(n28941), .B(n22538), .Z(n22303) );
  AND U22838 ( .A(n22304), .B(n22303), .Z(n22572) );
  NANDN U22839 ( .A(n35936), .B(n22305), .Z(n22307) );
  XOR U22840 ( .A(b[37]), .B(a[71]), .Z(n22541) );
  NANDN U22841 ( .A(n36047), .B(n22541), .Z(n22306) );
  NAND U22842 ( .A(n22307), .B(n22306), .Z(n22571) );
  XOR U22843 ( .A(n22572), .B(n22571), .Z(n22574) );
  XNOR U22844 ( .A(n22573), .B(n22574), .Z(n22502) );
  XNOR U22845 ( .A(n22503), .B(n22502), .Z(n22504) );
  NANDN U22846 ( .A(n22309), .B(n22308), .Z(n22313) );
  OR U22847 ( .A(n22311), .B(n22310), .Z(n22312) );
  NAND U22848 ( .A(n22313), .B(n22312), .Z(n22505) );
  XOR U22849 ( .A(n22504), .B(n22505), .Z(n22608) );
  XNOR U22850 ( .A(n22607), .B(n22608), .Z(n22609) );
  XNOR U22851 ( .A(n22610), .B(n22609), .Z(n22393) );
  XOR U22852 ( .A(n22394), .B(n22393), .Z(n22386) );
  NANDN U22853 ( .A(n22315), .B(n22314), .Z(n22319) );
  NANDN U22854 ( .A(n22317), .B(n22316), .Z(n22318) );
  AND U22855 ( .A(n22319), .B(n22318), .Z(n22385) );
  XNOR U22856 ( .A(n22386), .B(n22385), .Z(n22387) );
  XOR U22857 ( .A(n22388), .B(n22387), .Z(n22350) );
  XNOR U22858 ( .A(n22349), .B(n22350), .Z(n22351) );
  XOR U22859 ( .A(n22352), .B(n22351), .Z(n22616) );
  XNOR U22860 ( .A(n22615), .B(n22616), .Z(n22621) );
  XOR U22861 ( .A(n22622), .B(n22621), .Z(n22344) );
  NANDN U22862 ( .A(n22321), .B(n22320), .Z(n22325) );
  OR U22863 ( .A(n22323), .B(n22322), .Z(n22324) );
  NAND U22864 ( .A(n22325), .B(n22324), .Z(n22343) );
  XNOR U22865 ( .A(n22344), .B(n22343), .Z(n22345) );
  NANDN U22866 ( .A(n22327), .B(n22326), .Z(n22331) );
  NANDN U22867 ( .A(n22329), .B(n22328), .Z(n22330) );
  NAND U22868 ( .A(n22331), .B(n22330), .Z(n22346) );
  XOR U22869 ( .A(n22345), .B(n22346), .Z(n22338) );
  XNOR U22870 ( .A(n22337), .B(n22338), .Z(n22339) );
  XNOR U22871 ( .A(n22340), .B(n22339), .Z(n22625) );
  XNOR U22872 ( .A(sreg[171]), .B(n22625), .Z(n22627) );
  NANDN U22873 ( .A(sreg[170]), .B(n22332), .Z(n22336) );
  NAND U22874 ( .A(n22334), .B(n22333), .Z(n22335) );
  NAND U22875 ( .A(n22336), .B(n22335), .Z(n22626) );
  XNOR U22876 ( .A(n22627), .B(n22626), .Z(c[171]) );
  NANDN U22877 ( .A(n22338), .B(n22337), .Z(n22342) );
  NANDN U22878 ( .A(n22340), .B(n22339), .Z(n22341) );
  AND U22879 ( .A(n22342), .B(n22341), .Z(n22633) );
  NANDN U22880 ( .A(n22344), .B(n22343), .Z(n22348) );
  NANDN U22881 ( .A(n22346), .B(n22345), .Z(n22347) );
  AND U22882 ( .A(n22348), .B(n22347), .Z(n22631) );
  NANDN U22883 ( .A(n22350), .B(n22349), .Z(n22354) );
  NANDN U22884 ( .A(n22352), .B(n22351), .Z(n22353) );
  AND U22885 ( .A(n22354), .B(n22353), .Z(n22911) );
  NANDN U22886 ( .A(n22356), .B(n22355), .Z(n22360) );
  OR U22887 ( .A(n22358), .B(n22357), .Z(n22359) );
  AND U22888 ( .A(n22360), .B(n22359), .Z(n22910) );
  XNOR U22889 ( .A(n22911), .B(n22910), .Z(n22913) );
  NANDN U22890 ( .A(n22362), .B(n22361), .Z(n22366) );
  OR U22891 ( .A(n22364), .B(n22363), .Z(n22365) );
  AND U22892 ( .A(n22366), .B(n22365), .Z(n22900) );
  NANDN U22893 ( .A(n22368), .B(n22367), .Z(n22372) );
  NAND U22894 ( .A(n22370), .B(n22369), .Z(n22371) );
  AND U22895 ( .A(n22372), .B(n22371), .Z(n22899) );
  NANDN U22896 ( .A(n22374), .B(n22373), .Z(n22378) );
  NANDN U22897 ( .A(n22376), .B(n22375), .Z(n22377) );
  AND U22898 ( .A(n22378), .B(n22377), .Z(n22898) );
  XOR U22899 ( .A(n22899), .B(n22898), .Z(n22901) );
  XOR U22900 ( .A(n22900), .B(n22901), .Z(n22905) );
  NANDN U22901 ( .A(n22380), .B(n22379), .Z(n22384) );
  NANDN U22902 ( .A(n22382), .B(n22381), .Z(n22383) );
  NAND U22903 ( .A(n22384), .B(n22383), .Z(n22904) );
  XNOR U22904 ( .A(n22905), .B(n22904), .Z(n22906) );
  NANDN U22905 ( .A(n22386), .B(n22385), .Z(n22390) );
  NANDN U22906 ( .A(n22388), .B(n22387), .Z(n22389) );
  AND U22907 ( .A(n22390), .B(n22389), .Z(n22895) );
  NANDN U22908 ( .A(n22392), .B(n22391), .Z(n22396) );
  NAND U22909 ( .A(n22394), .B(n22393), .Z(n22395) );
  AND U22910 ( .A(n22396), .B(n22395), .Z(n22870) );
  NANDN U22911 ( .A(n22398), .B(n22397), .Z(n22402) );
  NANDN U22912 ( .A(n22400), .B(n22399), .Z(n22401) );
  AND U22913 ( .A(n22402), .B(n22401), .Z(n22888) );
  NANDN U22914 ( .A(n22404), .B(n22403), .Z(n22408) );
  NANDN U22915 ( .A(n22406), .B(n22405), .Z(n22407) );
  AND U22916 ( .A(n22408), .B(n22407), .Z(n22887) );
  NANDN U22917 ( .A(n33875), .B(n22409), .Z(n22411) );
  XOR U22918 ( .A(b[25]), .B(a[84]), .Z(n22666) );
  NANDN U22919 ( .A(n33994), .B(n22666), .Z(n22410) );
  AND U22920 ( .A(n22411), .B(n22410), .Z(n22836) );
  NANDN U22921 ( .A(n32013), .B(n22412), .Z(n22414) );
  XOR U22922 ( .A(a[92]), .B(b[17]), .Z(n22669) );
  NANDN U22923 ( .A(n32292), .B(n22669), .Z(n22413) );
  AND U22924 ( .A(n22414), .B(n22413), .Z(n22835) );
  NANDN U22925 ( .A(n31536), .B(n22415), .Z(n22417) );
  XOR U22926 ( .A(a[94]), .B(b[15]), .Z(n22672) );
  NANDN U22927 ( .A(n31925), .B(n22672), .Z(n22416) );
  NAND U22928 ( .A(n22417), .B(n22416), .Z(n22834) );
  XOR U22929 ( .A(n22835), .B(n22834), .Z(n22837) );
  XOR U22930 ( .A(n22836), .B(n22837), .Z(n22808) );
  NANDN U22931 ( .A(n37526), .B(n22418), .Z(n22420) );
  XOR U22932 ( .A(b[51]), .B(a[58]), .Z(n22675) );
  NANDN U22933 ( .A(n37605), .B(n22675), .Z(n22419) );
  AND U22934 ( .A(n22420), .B(n22419), .Z(n22860) );
  NANDN U22935 ( .A(n37705), .B(n22421), .Z(n22423) );
  XOR U22936 ( .A(b[53]), .B(a[56]), .Z(n22678) );
  NANDN U22937 ( .A(n37778), .B(n22678), .Z(n22422) );
  AND U22938 ( .A(n22423), .B(n22422), .Z(n22859) );
  NANDN U22939 ( .A(n36210), .B(n22424), .Z(n22426) );
  XOR U22940 ( .A(b[39]), .B(a[70]), .Z(n22681) );
  NANDN U22941 ( .A(n36347), .B(n22681), .Z(n22425) );
  NAND U22942 ( .A(n22426), .B(n22425), .Z(n22858) );
  XOR U22943 ( .A(n22859), .B(n22858), .Z(n22861) );
  XNOR U22944 ( .A(n22860), .B(n22861), .Z(n22807) );
  XNOR U22945 ( .A(n22808), .B(n22807), .Z(n22810) );
  NANDN U22946 ( .A(n22428), .B(n22427), .Z(n22432) );
  OR U22947 ( .A(n22430), .B(n22429), .Z(n22431) );
  AND U22948 ( .A(n22432), .B(n22431), .Z(n22809) );
  XOR U22949 ( .A(n22810), .B(n22809), .Z(n22657) );
  NANDN U22950 ( .A(n22434), .B(n22433), .Z(n22438) );
  OR U22951 ( .A(n22436), .B(n22435), .Z(n22437) );
  AND U22952 ( .A(n22438), .B(n22437), .Z(n22655) );
  NANDN U22953 ( .A(n22440), .B(n22439), .Z(n22444) );
  NANDN U22954 ( .A(n22442), .B(n22441), .Z(n22443) );
  NAND U22955 ( .A(n22444), .B(n22443), .Z(n22654) );
  XNOR U22956 ( .A(n22655), .B(n22654), .Z(n22656) );
  XNOR U22957 ( .A(n22657), .B(n22656), .Z(n22886) );
  XOR U22958 ( .A(n22887), .B(n22886), .Z(n22889) );
  XOR U22959 ( .A(n22888), .B(n22889), .Z(n22869) );
  NANDN U22960 ( .A(n22446), .B(n22445), .Z(n22450) );
  NANDN U22961 ( .A(n22448), .B(n22447), .Z(n22449) );
  AND U22962 ( .A(n22450), .B(n22449), .Z(n22881) );
  NANDN U22963 ( .A(n22451), .B(n37294), .Z(n22453) );
  XOR U22964 ( .A(b[47]), .B(a[62]), .Z(n22729) );
  NANDN U22965 ( .A(n37172), .B(n22729), .Z(n22452) );
  AND U22966 ( .A(n22453), .B(n22452), .Z(n22719) );
  NANDN U22967 ( .A(n22454), .B(n30627), .Z(n22456) );
  XOR U22968 ( .A(a[100]), .B(b[9]), .Z(n22732) );
  NANDN U22969 ( .A(n30267), .B(n22732), .Z(n22455) );
  AND U22970 ( .A(n22456), .B(n22455), .Z(n22718) );
  NANDN U22971 ( .A(n22457), .B(n37536), .Z(n22459) );
  XOR U22972 ( .A(b[49]), .B(a[60]), .Z(n22735) );
  NANDN U22973 ( .A(n37432), .B(n22735), .Z(n22458) );
  NAND U22974 ( .A(n22459), .B(n22458), .Z(n22717) );
  XOR U22975 ( .A(n22718), .B(n22717), .Z(n22720) );
  XOR U22976 ( .A(n22719), .B(n22720), .Z(n22814) );
  NANDN U22977 ( .A(n36742), .B(n22460), .Z(n22462) );
  XOR U22978 ( .A(b[43]), .B(a[66]), .Z(n22738) );
  NANDN U22979 ( .A(n36891), .B(n22738), .Z(n22461) );
  AND U22980 ( .A(n22462), .B(n22461), .Z(n22749) );
  NANDN U22981 ( .A(n36991), .B(n22463), .Z(n22465) );
  XOR U22982 ( .A(b[45]), .B(a[64]), .Z(n22741) );
  NANDN U22983 ( .A(n37083), .B(n22741), .Z(n22464) );
  AND U22984 ( .A(n22465), .B(n22464), .Z(n22748) );
  NANDN U22985 ( .A(n30482), .B(n22466), .Z(n22468) );
  XOR U22986 ( .A(a[98]), .B(b[11]), .Z(n22744) );
  NANDN U22987 ( .A(n30891), .B(n22744), .Z(n22467) );
  NAND U22988 ( .A(n22468), .B(n22467), .Z(n22747) );
  XOR U22989 ( .A(n22748), .B(n22747), .Z(n22750) );
  XNOR U22990 ( .A(n22749), .B(n22750), .Z(n22813) );
  XNOR U22991 ( .A(n22814), .B(n22813), .Z(n22815) );
  NANDN U22992 ( .A(n22470), .B(n22469), .Z(n22474) );
  OR U22993 ( .A(n22472), .B(n22471), .Z(n22473) );
  NAND U22994 ( .A(n22474), .B(n22473), .Z(n22816) );
  XNOR U22995 ( .A(n22815), .B(n22816), .Z(n22880) );
  XNOR U22996 ( .A(n22881), .B(n22880), .Z(n22882) );
  NANDN U22997 ( .A(n29499), .B(n22475), .Z(n22477) );
  XOR U22998 ( .A(a[102]), .B(b[7]), .Z(n22702) );
  NANDN U22999 ( .A(n29735), .B(n22702), .Z(n22476) );
  AND U23000 ( .A(n22477), .B(n22476), .Z(n22692) );
  NANDN U23001 ( .A(n37857), .B(n22478), .Z(n22480) );
  XOR U23002 ( .A(b[55]), .B(a[54]), .Z(n22705) );
  NANDN U23003 ( .A(n37911), .B(n22705), .Z(n22479) );
  AND U23004 ( .A(n22480), .B(n22479), .Z(n22691) );
  NANDN U23005 ( .A(n35611), .B(n22481), .Z(n22483) );
  XOR U23006 ( .A(b[35]), .B(a[74]), .Z(n22708) );
  NANDN U23007 ( .A(n35801), .B(n22708), .Z(n22482) );
  NAND U23008 ( .A(n22483), .B(n22482), .Z(n22690) );
  XOR U23009 ( .A(n22691), .B(n22690), .Z(n22693) );
  XOR U23010 ( .A(n22692), .B(n22693), .Z(n22766) );
  NANDN U23011 ( .A(n22485), .B(n22484), .Z(n22489) );
  OR U23012 ( .A(n22487), .B(n22486), .Z(n22488) );
  AND U23013 ( .A(n22489), .B(n22488), .Z(n22765) );
  XNOR U23014 ( .A(n22766), .B(n22765), .Z(n22767) );
  NAND U23015 ( .A(n22491), .B(n22490), .Z(n22495) );
  NANDN U23016 ( .A(n22493), .B(n22492), .Z(n22494) );
  NAND U23017 ( .A(n22495), .B(n22494), .Z(n22768) );
  XOR U23018 ( .A(n22767), .B(n22768), .Z(n22883) );
  XNOR U23019 ( .A(n22882), .B(n22883), .Z(n22868) );
  XOR U23020 ( .A(n22869), .B(n22868), .Z(n22871) );
  XOR U23021 ( .A(n22870), .B(n22871), .Z(n22893) );
  NANDN U23022 ( .A(n22497), .B(n22496), .Z(n22501) );
  NANDN U23023 ( .A(n22499), .B(n22498), .Z(n22500) );
  AND U23024 ( .A(n22501), .B(n22500), .Z(n22876) );
  NANDN U23025 ( .A(n22503), .B(n22502), .Z(n22507) );
  NANDN U23026 ( .A(n22505), .B(n22504), .Z(n22506) );
  AND U23027 ( .A(n22507), .B(n22506), .Z(n22875) );
  NANDN U23028 ( .A(n22509), .B(n22508), .Z(n22513) );
  NAND U23029 ( .A(n22511), .B(n22510), .Z(n22512) );
  AND U23030 ( .A(n22513), .B(n22512), .Z(n22874) );
  XOR U23031 ( .A(n22875), .B(n22874), .Z(n22877) );
  XOR U23032 ( .A(n22876), .B(n22877), .Z(n22645) );
  NAND U23033 ( .A(n22515), .B(n22514), .Z(n22519) );
  NANDN U23034 ( .A(n22517), .B(n22516), .Z(n22518) );
  AND U23035 ( .A(n22519), .B(n22518), .Z(n22867) );
  NANDN U23036 ( .A(n22521), .B(n22520), .Z(n22525) );
  OR U23037 ( .A(n22523), .B(n22522), .Z(n22524) );
  AND U23038 ( .A(n22525), .B(n22524), .Z(n22755) );
  NANDN U23039 ( .A(n34223), .B(n22526), .Z(n22528) );
  XOR U23040 ( .A(b[27]), .B(a[82]), .Z(n22840) );
  NANDN U23041 ( .A(n34458), .B(n22840), .Z(n22527) );
  AND U23042 ( .A(n22528), .B(n22527), .Z(n22687) );
  NANDN U23043 ( .A(n34634), .B(n22529), .Z(n22531) );
  XOR U23044 ( .A(b[29]), .B(a[80]), .Z(n22843) );
  NANDN U23045 ( .A(n34722), .B(n22843), .Z(n22530) );
  AND U23046 ( .A(n22531), .B(n22530), .Z(n22685) );
  NANDN U23047 ( .A(n31055), .B(n22532), .Z(n22534) );
  XOR U23048 ( .A(a[96]), .B(b[13]), .Z(n22846) );
  NANDN U23049 ( .A(n31293), .B(n22846), .Z(n22533) );
  NAND U23050 ( .A(n22534), .B(n22533), .Z(n22684) );
  XNOR U23051 ( .A(n22685), .B(n22684), .Z(n22686) );
  XOR U23052 ( .A(n22687), .B(n22686), .Z(n22754) );
  NANDN U23053 ( .A(n28889), .B(n22535), .Z(n22537) );
  XOR U23054 ( .A(a[104]), .B(b[5]), .Z(n22849) );
  NANDN U23055 ( .A(n29138), .B(n22849), .Z(n22536) );
  AND U23056 ( .A(n22537), .B(n22536), .Z(n22780) );
  NANDN U23057 ( .A(n209), .B(n22538), .Z(n22540) );
  XOR U23058 ( .A(a[106]), .B(b[3]), .Z(n22852) );
  NANDN U23059 ( .A(n28941), .B(n22852), .Z(n22539) );
  AND U23060 ( .A(n22540), .B(n22539), .Z(n22778) );
  NANDN U23061 ( .A(n35936), .B(n22541), .Z(n22543) );
  XOR U23062 ( .A(b[37]), .B(a[72]), .Z(n22855) );
  NANDN U23063 ( .A(n36047), .B(n22855), .Z(n22542) );
  NAND U23064 ( .A(n22543), .B(n22542), .Z(n22777) );
  XNOR U23065 ( .A(n22778), .B(n22777), .Z(n22779) );
  XOR U23066 ( .A(n22780), .B(n22779), .Z(n22753) );
  XNOR U23067 ( .A(n22754), .B(n22753), .Z(n22756) );
  NANDN U23068 ( .A(n22545), .B(n22544), .Z(n22549) );
  OR U23069 ( .A(n22547), .B(n22546), .Z(n22548) );
  AND U23070 ( .A(n22549), .B(n22548), .Z(n22725) );
  NANDN U23071 ( .A(n32996), .B(n22550), .Z(n22552) );
  XOR U23072 ( .A(a[88]), .B(b[21]), .Z(n22819) );
  NANDN U23073 ( .A(n33271), .B(n22819), .Z(n22551) );
  AND U23074 ( .A(n22552), .B(n22551), .Z(n22786) );
  NANDN U23075 ( .A(n33866), .B(n22553), .Z(n22555) );
  XOR U23076 ( .A(b[23]), .B(a[86]), .Z(n22822) );
  NANDN U23077 ( .A(n33644), .B(n22822), .Z(n22554) );
  AND U23078 ( .A(n22555), .B(n22554), .Z(n22784) );
  NANDN U23079 ( .A(n32483), .B(n22556), .Z(n22558) );
  XOR U23080 ( .A(a[90]), .B(b[19]), .Z(n22825) );
  NANDN U23081 ( .A(n32823), .B(n22825), .Z(n22557) );
  NAND U23082 ( .A(n22558), .B(n22557), .Z(n22783) );
  XNOR U23083 ( .A(n22784), .B(n22783), .Z(n22785) );
  XOR U23084 ( .A(n22786), .B(n22785), .Z(n22724) );
  NANDN U23085 ( .A(n34909), .B(n22559), .Z(n22561) );
  XOR U23086 ( .A(b[31]), .B(a[78]), .Z(n22828) );
  NANDN U23087 ( .A(n35145), .B(n22828), .Z(n22560) );
  AND U23088 ( .A(n22561), .B(n22560), .Z(n22714) );
  NANDN U23089 ( .A(n38247), .B(n22562), .Z(n22564) );
  XOR U23090 ( .A(b[61]), .B(a[48]), .Z(n22831) );
  NANDN U23091 ( .A(n38248), .B(n22831), .Z(n22563) );
  AND U23092 ( .A(n22564), .B(n22563), .Z(n22712) );
  AND U23093 ( .A(b[63]), .B(a[44]), .Z(n22711) );
  XNOR U23094 ( .A(n22712), .B(n22711), .Z(n22713) );
  XOR U23095 ( .A(n22714), .B(n22713), .Z(n22723) );
  XNOR U23096 ( .A(n22724), .B(n22723), .Z(n22726) );
  XOR U23097 ( .A(n22865), .B(n22864), .Z(n22866) );
  XNOR U23098 ( .A(n22867), .B(n22866), .Z(n22651) );
  NANDN U23099 ( .A(n22566), .B(n22565), .Z(n22570) );
  NANDN U23100 ( .A(n22568), .B(n22567), .Z(n22569) );
  AND U23101 ( .A(n22570), .B(n22569), .Z(n22760) );
  NANDN U23102 ( .A(n22572), .B(n22571), .Z(n22576) );
  OR U23103 ( .A(n22574), .B(n22573), .Z(n22575) );
  NAND U23104 ( .A(n22576), .B(n22575), .Z(n22759) );
  XNOR U23105 ( .A(n22760), .B(n22759), .Z(n22762) );
  NANDN U23106 ( .A(n22578), .B(n22577), .Z(n22582) );
  OR U23107 ( .A(n22580), .B(n22579), .Z(n22581) );
  NAND U23108 ( .A(n22582), .B(n22581), .Z(n22662) );
  NANDN U23109 ( .A(n38278), .B(n22583), .Z(n22585) );
  XOR U23110 ( .A(b[63]), .B(a[46]), .Z(n22792) );
  NANDN U23111 ( .A(n38279), .B(n22792), .Z(n22584) );
  AND U23112 ( .A(n22585), .B(n22584), .Z(n22697) );
  NANDN U23113 ( .A(n35260), .B(n22586), .Z(n22588) );
  XOR U23114 ( .A(b[33]), .B(a[76]), .Z(n22795) );
  NANDN U23115 ( .A(n35456), .B(n22795), .Z(n22587) );
  NAND U23116 ( .A(n22588), .B(n22587), .Z(n22696) );
  XNOR U23117 ( .A(n22697), .B(n22696), .Z(n22698) );
  NAND U23118 ( .A(b[0]), .B(a[108]), .Z(n22589) );
  XNOR U23119 ( .A(b[1]), .B(n22589), .Z(n22591) );
  NANDN U23120 ( .A(b[0]), .B(a[107]), .Z(n22590) );
  NAND U23121 ( .A(n22591), .B(n22590), .Z(n22699) );
  XNOR U23122 ( .A(n22698), .B(n22699), .Z(n22661) );
  NANDN U23123 ( .A(n37974), .B(n22592), .Z(n22594) );
  XOR U23124 ( .A(b[57]), .B(a[52]), .Z(n22798) );
  NANDN U23125 ( .A(n38031), .B(n22798), .Z(n22593) );
  AND U23126 ( .A(n22594), .B(n22593), .Z(n22773) );
  NANDN U23127 ( .A(n38090), .B(n22595), .Z(n22597) );
  XOR U23128 ( .A(b[59]), .B(a[50]), .Z(n22801) );
  NANDN U23129 ( .A(n38130), .B(n22801), .Z(n22596) );
  AND U23130 ( .A(n22597), .B(n22596), .Z(n22772) );
  NANDN U23131 ( .A(n36480), .B(n22598), .Z(n22600) );
  XOR U23132 ( .A(b[41]), .B(a[68]), .Z(n22804) );
  NANDN U23133 ( .A(n36594), .B(n22804), .Z(n22599) );
  NAND U23134 ( .A(n22600), .B(n22599), .Z(n22771) );
  XOR U23135 ( .A(n22772), .B(n22771), .Z(n22774) );
  XOR U23136 ( .A(n22773), .B(n22774), .Z(n22660) );
  XOR U23137 ( .A(n22661), .B(n22660), .Z(n22663) );
  XOR U23138 ( .A(n22662), .B(n22663), .Z(n22761) );
  XOR U23139 ( .A(n22762), .B(n22761), .Z(n22649) );
  NANDN U23140 ( .A(n22602), .B(n22601), .Z(n22606) );
  NAND U23141 ( .A(n22604), .B(n22603), .Z(n22605) );
  NAND U23142 ( .A(n22606), .B(n22605), .Z(n22648) );
  XNOR U23143 ( .A(n22649), .B(n22648), .Z(n22650) );
  XOR U23144 ( .A(n22651), .B(n22650), .Z(n22643) );
  NANDN U23145 ( .A(n22608), .B(n22607), .Z(n22612) );
  NANDN U23146 ( .A(n22610), .B(n22609), .Z(n22611) );
  AND U23147 ( .A(n22612), .B(n22611), .Z(n22642) );
  XNOR U23148 ( .A(n22643), .B(n22642), .Z(n22644) );
  XNOR U23149 ( .A(n22645), .B(n22644), .Z(n22892) );
  XNOR U23150 ( .A(n22893), .B(n22892), .Z(n22894) );
  XOR U23151 ( .A(n22895), .B(n22894), .Z(n22907) );
  XNOR U23152 ( .A(n22906), .B(n22907), .Z(n22912) );
  XOR U23153 ( .A(n22913), .B(n22912), .Z(n22637) );
  NANDN U23154 ( .A(n22614), .B(n22613), .Z(n22618) );
  NANDN U23155 ( .A(n22616), .B(n22615), .Z(n22617) );
  AND U23156 ( .A(n22618), .B(n22617), .Z(n22636) );
  XNOR U23157 ( .A(n22637), .B(n22636), .Z(n22638) );
  NANDN U23158 ( .A(n22620), .B(n22619), .Z(n22624) );
  NAND U23159 ( .A(n22622), .B(n22621), .Z(n22623) );
  NAND U23160 ( .A(n22624), .B(n22623), .Z(n22639) );
  XNOR U23161 ( .A(n22638), .B(n22639), .Z(n22630) );
  XNOR U23162 ( .A(n22631), .B(n22630), .Z(n22632) );
  XNOR U23163 ( .A(n22633), .B(n22632), .Z(n22916) );
  XNOR U23164 ( .A(sreg[172]), .B(n22916), .Z(n22918) );
  NANDN U23165 ( .A(sreg[171]), .B(n22625), .Z(n22629) );
  NAND U23166 ( .A(n22627), .B(n22626), .Z(n22628) );
  NAND U23167 ( .A(n22629), .B(n22628), .Z(n22917) );
  XNOR U23168 ( .A(n22918), .B(n22917), .Z(c[172]) );
  NANDN U23169 ( .A(n22631), .B(n22630), .Z(n22635) );
  NANDN U23170 ( .A(n22633), .B(n22632), .Z(n22634) );
  AND U23171 ( .A(n22635), .B(n22634), .Z(n22924) );
  NANDN U23172 ( .A(n22637), .B(n22636), .Z(n22641) );
  NANDN U23173 ( .A(n22639), .B(n22638), .Z(n22640) );
  AND U23174 ( .A(n22641), .B(n22640), .Z(n22922) );
  NANDN U23175 ( .A(n22643), .B(n22642), .Z(n22647) );
  NANDN U23176 ( .A(n22645), .B(n22644), .Z(n22646) );
  AND U23177 ( .A(n22647), .B(n22646), .Z(n23187) );
  NANDN U23178 ( .A(n22649), .B(n22648), .Z(n22653) );
  NAND U23179 ( .A(n22651), .B(n22650), .Z(n22652) );
  AND U23180 ( .A(n22653), .B(n22652), .Z(n22935) );
  NANDN U23181 ( .A(n22655), .B(n22654), .Z(n22659) );
  NANDN U23182 ( .A(n22657), .B(n22656), .Z(n22658) );
  AND U23183 ( .A(n22659), .B(n22658), .Z(n22947) );
  NAND U23184 ( .A(n22661), .B(n22660), .Z(n22665) );
  NAND U23185 ( .A(n22663), .B(n22662), .Z(n22664) );
  AND U23186 ( .A(n22665), .B(n22664), .Z(n22946) );
  NANDN U23187 ( .A(n33875), .B(n22666), .Z(n22668) );
  XOR U23188 ( .A(b[25]), .B(a[85]), .Z(n22981) );
  NANDN U23189 ( .A(n33994), .B(n22981), .Z(n22667) );
  AND U23190 ( .A(n22668), .B(n22667), .Z(n23151) );
  NANDN U23191 ( .A(n32013), .B(n22669), .Z(n22671) );
  XOR U23192 ( .A(a[93]), .B(b[17]), .Z(n22984) );
  NANDN U23193 ( .A(n32292), .B(n22984), .Z(n22670) );
  AND U23194 ( .A(n22671), .B(n22670), .Z(n23150) );
  NANDN U23195 ( .A(n31536), .B(n22672), .Z(n22674) );
  XOR U23196 ( .A(a[95]), .B(b[15]), .Z(n22987) );
  NANDN U23197 ( .A(n31925), .B(n22987), .Z(n22673) );
  NAND U23198 ( .A(n22674), .B(n22673), .Z(n23149) );
  XOR U23199 ( .A(n23150), .B(n23149), .Z(n23152) );
  XOR U23200 ( .A(n23151), .B(n23152), .Z(n23123) );
  NANDN U23201 ( .A(n37526), .B(n22675), .Z(n22677) );
  XOR U23202 ( .A(b[51]), .B(a[59]), .Z(n22990) );
  NANDN U23203 ( .A(n37605), .B(n22990), .Z(n22676) );
  AND U23204 ( .A(n22677), .B(n22676), .Z(n23175) );
  NANDN U23205 ( .A(n37705), .B(n22678), .Z(n22680) );
  XOR U23206 ( .A(b[53]), .B(a[57]), .Z(n22993) );
  NANDN U23207 ( .A(n37778), .B(n22993), .Z(n22679) );
  AND U23208 ( .A(n22680), .B(n22679), .Z(n23174) );
  NANDN U23209 ( .A(n36210), .B(n22681), .Z(n22683) );
  XOR U23210 ( .A(b[39]), .B(a[71]), .Z(n22996) );
  NANDN U23211 ( .A(n36347), .B(n22996), .Z(n22682) );
  NAND U23212 ( .A(n22683), .B(n22682), .Z(n23173) );
  XOR U23213 ( .A(n23174), .B(n23173), .Z(n23176) );
  XNOR U23214 ( .A(n23175), .B(n23176), .Z(n23122) );
  XNOR U23215 ( .A(n23123), .B(n23122), .Z(n23125) );
  NANDN U23216 ( .A(n22685), .B(n22684), .Z(n22689) );
  NANDN U23217 ( .A(n22687), .B(n22686), .Z(n22688) );
  AND U23218 ( .A(n22689), .B(n22688), .Z(n23124) );
  XOR U23219 ( .A(n23125), .B(n23124), .Z(n22972) );
  NANDN U23220 ( .A(n22691), .B(n22690), .Z(n22695) );
  OR U23221 ( .A(n22693), .B(n22692), .Z(n22694) );
  AND U23222 ( .A(n22695), .B(n22694), .Z(n22970) );
  NANDN U23223 ( .A(n22697), .B(n22696), .Z(n22701) );
  NANDN U23224 ( .A(n22699), .B(n22698), .Z(n22700) );
  NAND U23225 ( .A(n22701), .B(n22700), .Z(n22969) );
  XNOR U23226 ( .A(n22970), .B(n22969), .Z(n22971) );
  XNOR U23227 ( .A(n22972), .B(n22971), .Z(n22945) );
  XOR U23228 ( .A(n22946), .B(n22945), .Z(n22948) );
  XOR U23229 ( .A(n22947), .B(n22948), .Z(n22934) );
  NANDN U23230 ( .A(n29499), .B(n22702), .Z(n22704) );
  XOR U23231 ( .A(a[103]), .B(b[7]), .Z(n23017) );
  NANDN U23232 ( .A(n29735), .B(n23017), .Z(n22703) );
  AND U23233 ( .A(n22704), .B(n22703), .Z(n23007) );
  NANDN U23234 ( .A(n37857), .B(n22705), .Z(n22707) );
  XOR U23235 ( .A(b[55]), .B(a[55]), .Z(n23020) );
  NANDN U23236 ( .A(n37911), .B(n23020), .Z(n22706) );
  AND U23237 ( .A(n22707), .B(n22706), .Z(n23006) );
  NANDN U23238 ( .A(n35611), .B(n22708), .Z(n22710) );
  XOR U23239 ( .A(b[35]), .B(a[75]), .Z(n23023) );
  NANDN U23240 ( .A(n35801), .B(n23023), .Z(n22709) );
  NAND U23241 ( .A(n22710), .B(n22709), .Z(n23005) );
  XOR U23242 ( .A(n23006), .B(n23005), .Z(n23008) );
  XOR U23243 ( .A(n23007), .B(n23008), .Z(n23069) );
  NANDN U23244 ( .A(n22712), .B(n22711), .Z(n22716) );
  NANDN U23245 ( .A(n22714), .B(n22713), .Z(n22715) );
  AND U23246 ( .A(n22716), .B(n22715), .Z(n23068) );
  XNOR U23247 ( .A(n23069), .B(n23068), .Z(n23070) );
  NANDN U23248 ( .A(n22718), .B(n22717), .Z(n22722) );
  OR U23249 ( .A(n22720), .B(n22719), .Z(n22721) );
  NAND U23250 ( .A(n22722), .B(n22721), .Z(n23071) );
  XNOR U23251 ( .A(n23070), .B(n23071), .Z(n22953) );
  NAND U23252 ( .A(n22724), .B(n22723), .Z(n22728) );
  NANDN U23253 ( .A(n22726), .B(n22725), .Z(n22727) );
  AND U23254 ( .A(n22728), .B(n22727), .Z(n22952) );
  NANDN U23255 ( .A(n211), .B(n22729), .Z(n22731) );
  XOR U23256 ( .A(b[47]), .B(a[63]), .Z(n23044) );
  NANDN U23257 ( .A(n37172), .B(n23044), .Z(n22730) );
  AND U23258 ( .A(n22731), .B(n22730), .Z(n23034) );
  NANDN U23259 ( .A(n210), .B(n22732), .Z(n22734) );
  XOR U23260 ( .A(a[101]), .B(b[9]), .Z(n23047) );
  NANDN U23261 ( .A(n30267), .B(n23047), .Z(n22733) );
  AND U23262 ( .A(n22734), .B(n22733), .Z(n23033) );
  NANDN U23263 ( .A(n212), .B(n22735), .Z(n22737) );
  XOR U23264 ( .A(b[49]), .B(a[61]), .Z(n23050) );
  NANDN U23265 ( .A(n37432), .B(n23050), .Z(n22736) );
  NAND U23266 ( .A(n22737), .B(n22736), .Z(n23032) );
  XOR U23267 ( .A(n23033), .B(n23032), .Z(n23035) );
  XOR U23268 ( .A(n23034), .B(n23035), .Z(n23129) );
  NANDN U23269 ( .A(n36742), .B(n22738), .Z(n22740) );
  XOR U23270 ( .A(b[43]), .B(a[67]), .Z(n23053) );
  NANDN U23271 ( .A(n36891), .B(n23053), .Z(n22739) );
  AND U23272 ( .A(n22740), .B(n22739), .Z(n23064) );
  NANDN U23273 ( .A(n36991), .B(n22741), .Z(n22743) );
  XOR U23274 ( .A(b[45]), .B(a[65]), .Z(n23056) );
  NANDN U23275 ( .A(n37083), .B(n23056), .Z(n22742) );
  AND U23276 ( .A(n22743), .B(n22742), .Z(n23063) );
  NANDN U23277 ( .A(n30482), .B(n22744), .Z(n22746) );
  XOR U23278 ( .A(a[99]), .B(b[11]), .Z(n23059) );
  NANDN U23279 ( .A(n30891), .B(n23059), .Z(n22745) );
  NAND U23280 ( .A(n22746), .B(n22745), .Z(n23062) );
  XOR U23281 ( .A(n23063), .B(n23062), .Z(n23065) );
  XNOR U23282 ( .A(n23064), .B(n23065), .Z(n23128) );
  XNOR U23283 ( .A(n23129), .B(n23128), .Z(n23130) );
  NANDN U23284 ( .A(n22748), .B(n22747), .Z(n22752) );
  OR U23285 ( .A(n22750), .B(n22749), .Z(n22751) );
  NAND U23286 ( .A(n22752), .B(n22751), .Z(n23131) );
  XNOR U23287 ( .A(n23130), .B(n23131), .Z(n22951) );
  XOR U23288 ( .A(n22952), .B(n22951), .Z(n22954) );
  XNOR U23289 ( .A(n22953), .B(n22954), .Z(n22933) );
  XOR U23290 ( .A(n22934), .B(n22933), .Z(n22936) );
  XOR U23291 ( .A(n22935), .B(n22936), .Z(n23186) );
  NAND U23292 ( .A(n22754), .B(n22753), .Z(n22758) );
  NANDN U23293 ( .A(n22756), .B(n22755), .Z(n22757) );
  NAND U23294 ( .A(n22758), .B(n22757), .Z(n22939) );
  NANDN U23295 ( .A(n22760), .B(n22759), .Z(n22764) );
  NAND U23296 ( .A(n22762), .B(n22761), .Z(n22763) );
  AND U23297 ( .A(n22764), .B(n22763), .Z(n22940) );
  XOR U23298 ( .A(n22939), .B(n22940), .Z(n22942) );
  NANDN U23299 ( .A(n22766), .B(n22765), .Z(n22770) );
  NANDN U23300 ( .A(n22768), .B(n22767), .Z(n22769) );
  NAND U23301 ( .A(n22770), .B(n22769), .Z(n22941) );
  XOR U23302 ( .A(n22942), .B(n22941), .Z(n22960) );
  NANDN U23303 ( .A(n22772), .B(n22771), .Z(n22776) );
  OR U23304 ( .A(n22774), .B(n22773), .Z(n22775) );
  AND U23305 ( .A(n22776), .B(n22775), .Z(n23081) );
  NANDN U23306 ( .A(n22778), .B(n22777), .Z(n22782) );
  NANDN U23307 ( .A(n22780), .B(n22779), .Z(n22781) );
  NAND U23308 ( .A(n22782), .B(n22781), .Z(n23080) );
  XNOR U23309 ( .A(n23081), .B(n23080), .Z(n23083) );
  NANDN U23310 ( .A(n22784), .B(n22783), .Z(n22788) );
  NANDN U23311 ( .A(n22786), .B(n22785), .Z(n22787) );
  AND U23312 ( .A(n22788), .B(n22787), .Z(n22978) );
  NAND U23313 ( .A(b[0]), .B(a[109]), .Z(n22789) );
  XNOR U23314 ( .A(b[1]), .B(n22789), .Z(n22791) );
  NANDN U23315 ( .A(b[0]), .B(a[108]), .Z(n22790) );
  NAND U23316 ( .A(n22791), .B(n22790), .Z(n23014) );
  NANDN U23317 ( .A(n38278), .B(n22792), .Z(n22794) );
  XOR U23318 ( .A(b[63]), .B(a[47]), .Z(n23107) );
  NANDN U23319 ( .A(n38279), .B(n23107), .Z(n22793) );
  AND U23320 ( .A(n22794), .B(n22793), .Z(n23012) );
  NANDN U23321 ( .A(n35260), .B(n22795), .Z(n22797) );
  XOR U23322 ( .A(b[33]), .B(a[77]), .Z(n23110) );
  NANDN U23323 ( .A(n35456), .B(n23110), .Z(n22796) );
  NAND U23324 ( .A(n22797), .B(n22796), .Z(n23011) );
  XNOR U23325 ( .A(n23012), .B(n23011), .Z(n23013) );
  XNOR U23326 ( .A(n23014), .B(n23013), .Z(n22975) );
  NANDN U23327 ( .A(n37974), .B(n22798), .Z(n22800) );
  XOR U23328 ( .A(b[57]), .B(a[53]), .Z(n23113) );
  NANDN U23329 ( .A(n38031), .B(n23113), .Z(n22799) );
  AND U23330 ( .A(n22800), .B(n22799), .Z(n23089) );
  NANDN U23331 ( .A(n38090), .B(n22801), .Z(n22803) );
  XOR U23332 ( .A(b[59]), .B(a[51]), .Z(n23116) );
  NANDN U23333 ( .A(n38130), .B(n23116), .Z(n22802) );
  AND U23334 ( .A(n22803), .B(n22802), .Z(n23087) );
  NANDN U23335 ( .A(n36480), .B(n22804), .Z(n22806) );
  XOR U23336 ( .A(b[41]), .B(a[69]), .Z(n23119) );
  NANDN U23337 ( .A(n36594), .B(n23119), .Z(n22805) );
  NAND U23338 ( .A(n22806), .B(n22805), .Z(n23086) );
  XNOR U23339 ( .A(n23087), .B(n23086), .Z(n23088) );
  XOR U23340 ( .A(n23089), .B(n23088), .Z(n22976) );
  XNOR U23341 ( .A(n22975), .B(n22976), .Z(n22977) );
  XNOR U23342 ( .A(n22978), .B(n22977), .Z(n23082) );
  XOR U23343 ( .A(n23083), .B(n23082), .Z(n22964) );
  NANDN U23344 ( .A(n22808), .B(n22807), .Z(n22812) );
  NAND U23345 ( .A(n22810), .B(n22809), .Z(n22811) );
  NAND U23346 ( .A(n22812), .B(n22811), .Z(n22963) );
  XNOR U23347 ( .A(n22964), .B(n22963), .Z(n22966) );
  NANDN U23348 ( .A(n22814), .B(n22813), .Z(n22818) );
  NANDN U23349 ( .A(n22816), .B(n22815), .Z(n22817) );
  AND U23350 ( .A(n22818), .B(n22817), .Z(n23182) );
  NANDN U23351 ( .A(n32996), .B(n22819), .Z(n22821) );
  XOR U23352 ( .A(a[89]), .B(b[21]), .Z(n23134) );
  NANDN U23353 ( .A(n33271), .B(n23134), .Z(n22820) );
  AND U23354 ( .A(n22821), .B(n22820), .Z(n23100) );
  NANDN U23355 ( .A(n33866), .B(n22822), .Z(n22824) );
  XOR U23356 ( .A(b[23]), .B(a[87]), .Z(n23137) );
  NANDN U23357 ( .A(n33644), .B(n23137), .Z(n22823) );
  AND U23358 ( .A(n22824), .B(n22823), .Z(n23099) );
  NANDN U23359 ( .A(n32483), .B(n22825), .Z(n22827) );
  XOR U23360 ( .A(a[91]), .B(b[19]), .Z(n23140) );
  NANDN U23361 ( .A(n32823), .B(n23140), .Z(n22826) );
  NAND U23362 ( .A(n22827), .B(n22826), .Z(n23098) );
  XOR U23363 ( .A(n23099), .B(n23098), .Z(n23101) );
  XOR U23364 ( .A(n23100), .B(n23101), .Z(n23039) );
  NANDN U23365 ( .A(n34909), .B(n22828), .Z(n22830) );
  XOR U23366 ( .A(b[31]), .B(a[79]), .Z(n23143) );
  NANDN U23367 ( .A(n35145), .B(n23143), .Z(n22829) );
  AND U23368 ( .A(n22830), .B(n22829), .Z(n23028) );
  NANDN U23369 ( .A(n38247), .B(n22831), .Z(n22833) );
  XOR U23370 ( .A(b[61]), .B(a[49]), .Z(n23146) );
  NANDN U23371 ( .A(n38248), .B(n23146), .Z(n22832) );
  AND U23372 ( .A(n22833), .B(n22832), .Z(n23027) );
  AND U23373 ( .A(b[63]), .B(a[45]), .Z(n23026) );
  XOR U23374 ( .A(n23027), .B(n23026), .Z(n23029) );
  XNOR U23375 ( .A(n23028), .B(n23029), .Z(n23038) );
  XNOR U23376 ( .A(n23039), .B(n23038), .Z(n23040) );
  NANDN U23377 ( .A(n22835), .B(n22834), .Z(n22839) );
  OR U23378 ( .A(n22837), .B(n22836), .Z(n22838) );
  NAND U23379 ( .A(n22839), .B(n22838), .Z(n23041) );
  XNOR U23380 ( .A(n23040), .B(n23041), .Z(n23179) );
  NANDN U23381 ( .A(n34223), .B(n22840), .Z(n22842) );
  XOR U23382 ( .A(b[27]), .B(a[83]), .Z(n23155) );
  NANDN U23383 ( .A(n34458), .B(n23155), .Z(n22841) );
  AND U23384 ( .A(n22842), .B(n22841), .Z(n23001) );
  NANDN U23385 ( .A(n34634), .B(n22843), .Z(n22845) );
  XOR U23386 ( .A(b[29]), .B(a[81]), .Z(n23158) );
  NANDN U23387 ( .A(n34722), .B(n23158), .Z(n22844) );
  AND U23388 ( .A(n22845), .B(n22844), .Z(n23000) );
  NANDN U23389 ( .A(n31055), .B(n22846), .Z(n22848) );
  XOR U23390 ( .A(a[97]), .B(b[13]), .Z(n23161) );
  NANDN U23391 ( .A(n31293), .B(n23161), .Z(n22847) );
  NAND U23392 ( .A(n22848), .B(n22847), .Z(n22999) );
  XOR U23393 ( .A(n23000), .B(n22999), .Z(n23002) );
  XOR U23394 ( .A(n23001), .B(n23002), .Z(n23075) );
  NANDN U23395 ( .A(n28889), .B(n22849), .Z(n22851) );
  XOR U23396 ( .A(a[105]), .B(b[5]), .Z(n23164) );
  NANDN U23397 ( .A(n29138), .B(n23164), .Z(n22850) );
  AND U23398 ( .A(n22851), .B(n22850), .Z(n23094) );
  NANDN U23399 ( .A(n209), .B(n22852), .Z(n22854) );
  XOR U23400 ( .A(a[107]), .B(b[3]), .Z(n23167) );
  NANDN U23401 ( .A(n28941), .B(n23167), .Z(n22853) );
  AND U23402 ( .A(n22854), .B(n22853), .Z(n23093) );
  NANDN U23403 ( .A(n35936), .B(n22855), .Z(n22857) );
  XOR U23404 ( .A(b[37]), .B(a[73]), .Z(n23170) );
  NANDN U23405 ( .A(n36047), .B(n23170), .Z(n22856) );
  NAND U23406 ( .A(n22857), .B(n22856), .Z(n23092) );
  XOR U23407 ( .A(n23093), .B(n23092), .Z(n23095) );
  XNOR U23408 ( .A(n23094), .B(n23095), .Z(n23074) );
  XNOR U23409 ( .A(n23075), .B(n23074), .Z(n23076) );
  NANDN U23410 ( .A(n22859), .B(n22858), .Z(n22863) );
  OR U23411 ( .A(n22861), .B(n22860), .Z(n22862) );
  NAND U23412 ( .A(n22863), .B(n22862), .Z(n23077) );
  XOR U23413 ( .A(n23076), .B(n23077), .Z(n23180) );
  XNOR U23414 ( .A(n23179), .B(n23180), .Z(n23181) );
  XNOR U23415 ( .A(n23182), .B(n23181), .Z(n22965) );
  XOR U23416 ( .A(n22966), .B(n22965), .Z(n22958) );
  XNOR U23417 ( .A(n22958), .B(n22957), .Z(n22959) );
  XNOR U23418 ( .A(n22960), .B(n22959), .Z(n23185) );
  XOR U23419 ( .A(n23186), .B(n23185), .Z(n23188) );
  XOR U23420 ( .A(n23187), .B(n23188), .Z(n23199) );
  NANDN U23421 ( .A(n22869), .B(n22868), .Z(n22873) );
  OR U23422 ( .A(n22871), .B(n22870), .Z(n22872) );
  AND U23423 ( .A(n22873), .B(n22872), .Z(n23198) );
  NANDN U23424 ( .A(n22875), .B(n22874), .Z(n22879) );
  OR U23425 ( .A(n22877), .B(n22876), .Z(n22878) );
  AND U23426 ( .A(n22879), .B(n22878), .Z(n23194) );
  NANDN U23427 ( .A(n22881), .B(n22880), .Z(n22885) );
  NANDN U23428 ( .A(n22883), .B(n22882), .Z(n22884) );
  AND U23429 ( .A(n22885), .B(n22884), .Z(n23192) );
  NANDN U23430 ( .A(n22887), .B(n22886), .Z(n22891) );
  OR U23431 ( .A(n22889), .B(n22888), .Z(n22890) );
  AND U23432 ( .A(n22891), .B(n22890), .Z(n23191) );
  XNOR U23433 ( .A(n23192), .B(n23191), .Z(n23193) );
  XNOR U23434 ( .A(n23194), .B(n23193), .Z(n23197) );
  XOR U23435 ( .A(n23198), .B(n23197), .Z(n23200) );
  XOR U23436 ( .A(n23199), .B(n23200), .Z(n23205) );
  NANDN U23437 ( .A(n22893), .B(n22892), .Z(n22897) );
  NANDN U23438 ( .A(n22895), .B(n22894), .Z(n22896) );
  AND U23439 ( .A(n22897), .B(n22896), .Z(n23204) );
  NANDN U23440 ( .A(n22899), .B(n22898), .Z(n22903) );
  OR U23441 ( .A(n22901), .B(n22900), .Z(n22902) );
  AND U23442 ( .A(n22903), .B(n22902), .Z(n23203) );
  XOR U23443 ( .A(n23204), .B(n23203), .Z(n23206) );
  XOR U23444 ( .A(n23205), .B(n23206), .Z(n22928) );
  NANDN U23445 ( .A(n22905), .B(n22904), .Z(n22909) );
  NANDN U23446 ( .A(n22907), .B(n22906), .Z(n22908) );
  AND U23447 ( .A(n22909), .B(n22908), .Z(n22927) );
  XNOR U23448 ( .A(n22928), .B(n22927), .Z(n22929) );
  NANDN U23449 ( .A(n22911), .B(n22910), .Z(n22915) );
  NAND U23450 ( .A(n22913), .B(n22912), .Z(n22914) );
  NAND U23451 ( .A(n22915), .B(n22914), .Z(n22930) );
  XNOR U23452 ( .A(n22929), .B(n22930), .Z(n22921) );
  XNOR U23453 ( .A(n22922), .B(n22921), .Z(n22923) );
  XNOR U23454 ( .A(n22924), .B(n22923), .Z(n23209) );
  XNOR U23455 ( .A(sreg[173]), .B(n23209), .Z(n23211) );
  NANDN U23456 ( .A(sreg[172]), .B(n22916), .Z(n22920) );
  NAND U23457 ( .A(n22918), .B(n22917), .Z(n22919) );
  NAND U23458 ( .A(n22920), .B(n22919), .Z(n23210) );
  XNOR U23459 ( .A(n23211), .B(n23210), .Z(c[173]) );
  NANDN U23460 ( .A(n22922), .B(n22921), .Z(n22926) );
  NANDN U23461 ( .A(n22924), .B(n22923), .Z(n22925) );
  AND U23462 ( .A(n22926), .B(n22925), .Z(n23217) );
  NANDN U23463 ( .A(n22928), .B(n22927), .Z(n22932) );
  NANDN U23464 ( .A(n22930), .B(n22929), .Z(n22931) );
  AND U23465 ( .A(n22932), .B(n22931), .Z(n23215) );
  NANDN U23466 ( .A(n22934), .B(n22933), .Z(n22938) );
  OR U23467 ( .A(n22936), .B(n22935), .Z(n22937) );
  AND U23468 ( .A(n22938), .B(n22937), .Z(n23490) );
  NAND U23469 ( .A(n22940), .B(n22939), .Z(n22944) );
  NAND U23470 ( .A(n22942), .B(n22941), .Z(n22943) );
  AND U23471 ( .A(n22944), .B(n22943), .Z(n23234) );
  NANDN U23472 ( .A(n22946), .B(n22945), .Z(n22950) );
  OR U23473 ( .A(n22948), .B(n22947), .Z(n22949) );
  AND U23474 ( .A(n22950), .B(n22949), .Z(n23233) );
  NANDN U23475 ( .A(n22952), .B(n22951), .Z(n22956) );
  NANDN U23476 ( .A(n22954), .B(n22953), .Z(n22955) );
  AND U23477 ( .A(n22956), .B(n22955), .Z(n23232) );
  XOR U23478 ( .A(n23233), .B(n23232), .Z(n23235) );
  XOR U23479 ( .A(n23234), .B(n23235), .Z(n23491) );
  XNOR U23480 ( .A(n23490), .B(n23491), .Z(n23492) );
  NANDN U23481 ( .A(n22958), .B(n22957), .Z(n22962) );
  NANDN U23482 ( .A(n22960), .B(n22959), .Z(n22961) );
  AND U23483 ( .A(n22962), .B(n22961), .Z(n23229) );
  NANDN U23484 ( .A(n22964), .B(n22963), .Z(n22968) );
  NAND U23485 ( .A(n22966), .B(n22965), .Z(n22967) );
  AND U23486 ( .A(n22968), .B(n22967), .Z(n23258) );
  NANDN U23487 ( .A(n22970), .B(n22969), .Z(n22974) );
  NANDN U23488 ( .A(n22972), .B(n22971), .Z(n22973) );
  AND U23489 ( .A(n22974), .B(n22973), .Z(n23252) );
  NANDN U23490 ( .A(n22976), .B(n22975), .Z(n22980) );
  NANDN U23491 ( .A(n22978), .B(n22977), .Z(n22979) );
  AND U23492 ( .A(n22980), .B(n22979), .Z(n23251) );
  NANDN U23493 ( .A(n33875), .B(n22981), .Z(n22983) );
  XOR U23494 ( .A(b[25]), .B(a[86]), .Z(n23286) );
  NANDN U23495 ( .A(n33994), .B(n23286), .Z(n22982) );
  AND U23496 ( .A(n22983), .B(n22982), .Z(n23480) );
  NANDN U23497 ( .A(n32013), .B(n22984), .Z(n22986) );
  XOR U23498 ( .A(a[94]), .B(b[17]), .Z(n23289) );
  NANDN U23499 ( .A(n32292), .B(n23289), .Z(n22985) );
  AND U23500 ( .A(n22986), .B(n22985), .Z(n23479) );
  NANDN U23501 ( .A(n31536), .B(n22987), .Z(n22989) );
  XOR U23502 ( .A(a[96]), .B(b[15]), .Z(n23292) );
  NANDN U23503 ( .A(n31925), .B(n23292), .Z(n22988) );
  NAND U23504 ( .A(n22989), .B(n22988), .Z(n23478) );
  XOR U23505 ( .A(n23479), .B(n23478), .Z(n23481) );
  XOR U23506 ( .A(n23480), .B(n23481), .Z(n23428) );
  NANDN U23507 ( .A(n37526), .B(n22990), .Z(n22992) );
  XOR U23508 ( .A(b[51]), .B(a[60]), .Z(n23295) );
  NANDN U23509 ( .A(n37605), .B(n23295), .Z(n22991) );
  AND U23510 ( .A(n22992), .B(n22991), .Z(n23459) );
  NANDN U23511 ( .A(n37705), .B(n22993), .Z(n22995) );
  XOR U23512 ( .A(b[53]), .B(a[58]), .Z(n23298) );
  NANDN U23513 ( .A(n37778), .B(n23298), .Z(n22994) );
  AND U23514 ( .A(n22995), .B(n22994), .Z(n23458) );
  NANDN U23515 ( .A(n36210), .B(n22996), .Z(n22998) );
  XOR U23516 ( .A(b[39]), .B(a[72]), .Z(n23301) );
  NANDN U23517 ( .A(n36347), .B(n23301), .Z(n22997) );
  NAND U23518 ( .A(n22998), .B(n22997), .Z(n23457) );
  XOR U23519 ( .A(n23458), .B(n23457), .Z(n23460) );
  XNOR U23520 ( .A(n23459), .B(n23460), .Z(n23427) );
  XNOR U23521 ( .A(n23428), .B(n23427), .Z(n23430) );
  NANDN U23522 ( .A(n23000), .B(n22999), .Z(n23004) );
  OR U23523 ( .A(n23002), .B(n23001), .Z(n23003) );
  AND U23524 ( .A(n23004), .B(n23003), .Z(n23429) );
  XOR U23525 ( .A(n23430), .B(n23429), .Z(n23277) );
  NANDN U23526 ( .A(n23006), .B(n23005), .Z(n23010) );
  OR U23527 ( .A(n23008), .B(n23007), .Z(n23009) );
  AND U23528 ( .A(n23010), .B(n23009), .Z(n23275) );
  NANDN U23529 ( .A(n23012), .B(n23011), .Z(n23016) );
  NANDN U23530 ( .A(n23014), .B(n23013), .Z(n23015) );
  NAND U23531 ( .A(n23016), .B(n23015), .Z(n23274) );
  XNOR U23532 ( .A(n23275), .B(n23274), .Z(n23276) );
  XNOR U23533 ( .A(n23277), .B(n23276), .Z(n23250) );
  XOR U23534 ( .A(n23251), .B(n23250), .Z(n23253) );
  XOR U23535 ( .A(n23252), .B(n23253), .Z(n23257) );
  NANDN U23536 ( .A(n29499), .B(n23017), .Z(n23019) );
  XOR U23537 ( .A(a[104]), .B(b[7]), .Z(n23322) );
  NANDN U23538 ( .A(n29735), .B(n23322), .Z(n23018) );
  AND U23539 ( .A(n23019), .B(n23018), .Z(n23312) );
  NANDN U23540 ( .A(n37857), .B(n23020), .Z(n23022) );
  XOR U23541 ( .A(b[55]), .B(a[56]), .Z(n23325) );
  NANDN U23542 ( .A(n37911), .B(n23325), .Z(n23021) );
  AND U23543 ( .A(n23022), .B(n23021), .Z(n23311) );
  NANDN U23544 ( .A(n35611), .B(n23023), .Z(n23025) );
  XOR U23545 ( .A(b[35]), .B(a[76]), .Z(n23328) );
  NANDN U23546 ( .A(n35801), .B(n23328), .Z(n23024) );
  NAND U23547 ( .A(n23025), .B(n23024), .Z(n23310) );
  XOR U23548 ( .A(n23311), .B(n23310), .Z(n23313) );
  XOR U23549 ( .A(n23312), .B(n23313), .Z(n23374) );
  NANDN U23550 ( .A(n23027), .B(n23026), .Z(n23031) );
  OR U23551 ( .A(n23029), .B(n23028), .Z(n23030) );
  AND U23552 ( .A(n23031), .B(n23030), .Z(n23373) );
  XNOR U23553 ( .A(n23374), .B(n23373), .Z(n23375) );
  NANDN U23554 ( .A(n23033), .B(n23032), .Z(n23037) );
  OR U23555 ( .A(n23035), .B(n23034), .Z(n23036) );
  NAND U23556 ( .A(n23037), .B(n23036), .Z(n23376) );
  XNOR U23557 ( .A(n23375), .B(n23376), .Z(n23246) );
  NANDN U23558 ( .A(n23039), .B(n23038), .Z(n23043) );
  NANDN U23559 ( .A(n23041), .B(n23040), .Z(n23042) );
  AND U23560 ( .A(n23043), .B(n23042), .Z(n23245) );
  NANDN U23561 ( .A(n211), .B(n23044), .Z(n23046) );
  XOR U23562 ( .A(b[47]), .B(a[64]), .Z(n23349) );
  NANDN U23563 ( .A(n37172), .B(n23349), .Z(n23045) );
  AND U23564 ( .A(n23046), .B(n23045), .Z(n23339) );
  NANDN U23565 ( .A(n210), .B(n23047), .Z(n23049) );
  XOR U23566 ( .A(a[102]), .B(b[9]), .Z(n23352) );
  NANDN U23567 ( .A(n30267), .B(n23352), .Z(n23048) );
  AND U23568 ( .A(n23049), .B(n23048), .Z(n23338) );
  NANDN U23569 ( .A(n212), .B(n23050), .Z(n23052) );
  XOR U23570 ( .A(b[49]), .B(a[62]), .Z(n23355) );
  NANDN U23571 ( .A(n37432), .B(n23355), .Z(n23051) );
  NAND U23572 ( .A(n23052), .B(n23051), .Z(n23337) );
  XOR U23573 ( .A(n23338), .B(n23337), .Z(n23340) );
  XOR U23574 ( .A(n23339), .B(n23340), .Z(n23434) );
  NANDN U23575 ( .A(n36742), .B(n23053), .Z(n23055) );
  XOR U23576 ( .A(b[43]), .B(a[68]), .Z(n23358) );
  NANDN U23577 ( .A(n36891), .B(n23358), .Z(n23054) );
  AND U23578 ( .A(n23055), .B(n23054), .Z(n23369) );
  NANDN U23579 ( .A(n36991), .B(n23056), .Z(n23058) );
  XOR U23580 ( .A(b[45]), .B(a[66]), .Z(n23361) );
  NANDN U23581 ( .A(n37083), .B(n23361), .Z(n23057) );
  AND U23582 ( .A(n23058), .B(n23057), .Z(n23368) );
  NANDN U23583 ( .A(n30482), .B(n23059), .Z(n23061) );
  XOR U23584 ( .A(a[100]), .B(b[11]), .Z(n23364) );
  NANDN U23585 ( .A(n30891), .B(n23364), .Z(n23060) );
  NAND U23586 ( .A(n23061), .B(n23060), .Z(n23367) );
  XOR U23587 ( .A(n23368), .B(n23367), .Z(n23370) );
  XNOR U23588 ( .A(n23369), .B(n23370), .Z(n23433) );
  XNOR U23589 ( .A(n23434), .B(n23433), .Z(n23435) );
  NANDN U23590 ( .A(n23063), .B(n23062), .Z(n23067) );
  OR U23591 ( .A(n23065), .B(n23064), .Z(n23066) );
  NAND U23592 ( .A(n23067), .B(n23066), .Z(n23436) );
  XNOR U23593 ( .A(n23435), .B(n23436), .Z(n23244) );
  XOR U23594 ( .A(n23245), .B(n23244), .Z(n23247) );
  XNOR U23595 ( .A(n23246), .B(n23247), .Z(n23256) );
  XOR U23596 ( .A(n23257), .B(n23256), .Z(n23259) );
  XOR U23597 ( .A(n23258), .B(n23259), .Z(n23227) );
  NANDN U23598 ( .A(n23069), .B(n23068), .Z(n23073) );
  NANDN U23599 ( .A(n23071), .B(n23070), .Z(n23072) );
  AND U23600 ( .A(n23073), .B(n23072), .Z(n23240) );
  NANDN U23601 ( .A(n23075), .B(n23074), .Z(n23079) );
  NANDN U23602 ( .A(n23077), .B(n23076), .Z(n23078) );
  AND U23603 ( .A(n23079), .B(n23078), .Z(n23239) );
  NANDN U23604 ( .A(n23081), .B(n23080), .Z(n23085) );
  NAND U23605 ( .A(n23083), .B(n23082), .Z(n23084) );
  AND U23606 ( .A(n23085), .B(n23084), .Z(n23238) );
  XOR U23607 ( .A(n23239), .B(n23238), .Z(n23241) );
  XOR U23608 ( .A(n23240), .B(n23241), .Z(n23265) );
  NANDN U23609 ( .A(n23087), .B(n23086), .Z(n23091) );
  NANDN U23610 ( .A(n23089), .B(n23088), .Z(n23090) );
  AND U23611 ( .A(n23091), .B(n23090), .Z(n23386) );
  NANDN U23612 ( .A(n23093), .B(n23092), .Z(n23097) );
  OR U23613 ( .A(n23095), .B(n23094), .Z(n23096) );
  NAND U23614 ( .A(n23097), .B(n23096), .Z(n23385) );
  XNOR U23615 ( .A(n23386), .B(n23385), .Z(n23388) );
  NANDN U23616 ( .A(n23099), .B(n23098), .Z(n23103) );
  OR U23617 ( .A(n23101), .B(n23100), .Z(n23102) );
  AND U23618 ( .A(n23103), .B(n23102), .Z(n23283) );
  AND U23619 ( .A(a[110]), .B(b[0]), .Z(n23104) );
  XOR U23620 ( .A(b[1]), .B(n23104), .Z(n23106) );
  NANDN U23621 ( .A(b[0]), .B(a[109]), .Z(n23105) );
  AND U23622 ( .A(n23106), .B(n23105), .Z(n23318) );
  NANDN U23623 ( .A(n38278), .B(n23107), .Z(n23109) );
  XOR U23624 ( .A(b[63]), .B(a[48]), .Z(n23412) );
  NANDN U23625 ( .A(n38279), .B(n23412), .Z(n23108) );
  AND U23626 ( .A(n23109), .B(n23108), .Z(n23317) );
  NANDN U23627 ( .A(n35260), .B(n23110), .Z(n23112) );
  XOR U23628 ( .A(b[33]), .B(a[78]), .Z(n23415) );
  NANDN U23629 ( .A(n35456), .B(n23415), .Z(n23111) );
  NAND U23630 ( .A(n23112), .B(n23111), .Z(n23316) );
  XOR U23631 ( .A(n23317), .B(n23316), .Z(n23319) );
  XNOR U23632 ( .A(n23318), .B(n23319), .Z(n23280) );
  NANDN U23633 ( .A(n37974), .B(n23113), .Z(n23115) );
  XOR U23634 ( .A(b[57]), .B(a[54]), .Z(n23418) );
  NANDN U23635 ( .A(n38031), .B(n23418), .Z(n23114) );
  AND U23636 ( .A(n23115), .B(n23114), .Z(n23394) );
  NANDN U23637 ( .A(n38090), .B(n23116), .Z(n23118) );
  XOR U23638 ( .A(b[59]), .B(a[52]), .Z(n23421) );
  NANDN U23639 ( .A(n38130), .B(n23421), .Z(n23117) );
  AND U23640 ( .A(n23118), .B(n23117), .Z(n23392) );
  NANDN U23641 ( .A(n36480), .B(n23119), .Z(n23121) );
  XOR U23642 ( .A(b[41]), .B(a[70]), .Z(n23424) );
  NANDN U23643 ( .A(n36594), .B(n23424), .Z(n23120) );
  NAND U23644 ( .A(n23121), .B(n23120), .Z(n23391) );
  XNOR U23645 ( .A(n23392), .B(n23391), .Z(n23393) );
  XOR U23646 ( .A(n23394), .B(n23393), .Z(n23281) );
  XNOR U23647 ( .A(n23280), .B(n23281), .Z(n23282) );
  XNOR U23648 ( .A(n23283), .B(n23282), .Z(n23387) );
  XOR U23649 ( .A(n23388), .B(n23387), .Z(n23269) );
  NANDN U23650 ( .A(n23123), .B(n23122), .Z(n23127) );
  NAND U23651 ( .A(n23125), .B(n23124), .Z(n23126) );
  NAND U23652 ( .A(n23127), .B(n23126), .Z(n23268) );
  XNOR U23653 ( .A(n23269), .B(n23268), .Z(n23271) );
  NANDN U23654 ( .A(n23129), .B(n23128), .Z(n23133) );
  NANDN U23655 ( .A(n23131), .B(n23130), .Z(n23132) );
  AND U23656 ( .A(n23133), .B(n23132), .Z(n23487) );
  NANDN U23657 ( .A(n32996), .B(n23134), .Z(n23136) );
  XOR U23658 ( .A(a[90]), .B(b[21]), .Z(n23463) );
  NANDN U23659 ( .A(n33271), .B(n23463), .Z(n23135) );
  AND U23660 ( .A(n23136), .B(n23135), .Z(n23405) );
  NANDN U23661 ( .A(n33866), .B(n23137), .Z(n23139) );
  XOR U23662 ( .A(b[23]), .B(a[88]), .Z(n23466) );
  NANDN U23663 ( .A(n33644), .B(n23466), .Z(n23138) );
  AND U23664 ( .A(n23139), .B(n23138), .Z(n23404) );
  NANDN U23665 ( .A(n32483), .B(n23140), .Z(n23142) );
  XOR U23666 ( .A(a[92]), .B(b[19]), .Z(n23469) );
  NANDN U23667 ( .A(n32823), .B(n23469), .Z(n23141) );
  NAND U23668 ( .A(n23142), .B(n23141), .Z(n23403) );
  XOR U23669 ( .A(n23404), .B(n23403), .Z(n23406) );
  XOR U23670 ( .A(n23405), .B(n23406), .Z(n23344) );
  NANDN U23671 ( .A(n34909), .B(n23143), .Z(n23145) );
  XOR U23672 ( .A(b[31]), .B(a[80]), .Z(n23472) );
  NANDN U23673 ( .A(n35145), .B(n23472), .Z(n23144) );
  AND U23674 ( .A(n23145), .B(n23144), .Z(n23333) );
  NANDN U23675 ( .A(n38247), .B(n23146), .Z(n23148) );
  XOR U23676 ( .A(b[61]), .B(a[50]), .Z(n23475) );
  NANDN U23677 ( .A(n38248), .B(n23475), .Z(n23147) );
  AND U23678 ( .A(n23148), .B(n23147), .Z(n23332) );
  AND U23679 ( .A(b[63]), .B(a[46]), .Z(n23331) );
  XOR U23680 ( .A(n23332), .B(n23331), .Z(n23334) );
  XNOR U23681 ( .A(n23333), .B(n23334), .Z(n23343) );
  XNOR U23682 ( .A(n23344), .B(n23343), .Z(n23345) );
  NANDN U23683 ( .A(n23150), .B(n23149), .Z(n23154) );
  OR U23684 ( .A(n23152), .B(n23151), .Z(n23153) );
  NAND U23685 ( .A(n23154), .B(n23153), .Z(n23346) );
  XNOR U23686 ( .A(n23345), .B(n23346), .Z(n23484) );
  NANDN U23687 ( .A(n34223), .B(n23155), .Z(n23157) );
  XOR U23688 ( .A(b[27]), .B(a[84]), .Z(n23439) );
  NANDN U23689 ( .A(n34458), .B(n23439), .Z(n23156) );
  AND U23690 ( .A(n23157), .B(n23156), .Z(n23306) );
  NANDN U23691 ( .A(n34634), .B(n23158), .Z(n23160) );
  XOR U23692 ( .A(b[29]), .B(a[82]), .Z(n23442) );
  NANDN U23693 ( .A(n34722), .B(n23442), .Z(n23159) );
  AND U23694 ( .A(n23160), .B(n23159), .Z(n23305) );
  NANDN U23695 ( .A(n31055), .B(n23161), .Z(n23163) );
  XOR U23696 ( .A(a[98]), .B(b[13]), .Z(n23445) );
  NANDN U23697 ( .A(n31293), .B(n23445), .Z(n23162) );
  NAND U23698 ( .A(n23163), .B(n23162), .Z(n23304) );
  XOR U23699 ( .A(n23305), .B(n23304), .Z(n23307) );
  XOR U23700 ( .A(n23306), .B(n23307), .Z(n23380) );
  NANDN U23701 ( .A(n28889), .B(n23164), .Z(n23166) );
  XOR U23702 ( .A(a[106]), .B(b[5]), .Z(n23448) );
  NANDN U23703 ( .A(n29138), .B(n23448), .Z(n23165) );
  AND U23704 ( .A(n23166), .B(n23165), .Z(n23399) );
  NANDN U23705 ( .A(n209), .B(n23167), .Z(n23169) );
  XOR U23706 ( .A(a[108]), .B(b[3]), .Z(n23451) );
  NANDN U23707 ( .A(n28941), .B(n23451), .Z(n23168) );
  AND U23708 ( .A(n23169), .B(n23168), .Z(n23398) );
  NANDN U23709 ( .A(n35936), .B(n23170), .Z(n23172) );
  XOR U23710 ( .A(b[37]), .B(a[74]), .Z(n23454) );
  NANDN U23711 ( .A(n36047), .B(n23454), .Z(n23171) );
  NAND U23712 ( .A(n23172), .B(n23171), .Z(n23397) );
  XOR U23713 ( .A(n23398), .B(n23397), .Z(n23400) );
  XNOR U23714 ( .A(n23399), .B(n23400), .Z(n23379) );
  XNOR U23715 ( .A(n23380), .B(n23379), .Z(n23381) );
  NANDN U23716 ( .A(n23174), .B(n23173), .Z(n23178) );
  OR U23717 ( .A(n23176), .B(n23175), .Z(n23177) );
  NAND U23718 ( .A(n23178), .B(n23177), .Z(n23382) );
  XOR U23719 ( .A(n23381), .B(n23382), .Z(n23485) );
  XNOR U23720 ( .A(n23484), .B(n23485), .Z(n23486) );
  XNOR U23721 ( .A(n23487), .B(n23486), .Z(n23270) );
  XOR U23722 ( .A(n23271), .B(n23270), .Z(n23263) );
  NANDN U23723 ( .A(n23180), .B(n23179), .Z(n23184) );
  NANDN U23724 ( .A(n23182), .B(n23181), .Z(n23183) );
  AND U23725 ( .A(n23184), .B(n23183), .Z(n23262) );
  XNOR U23726 ( .A(n23263), .B(n23262), .Z(n23264) );
  XNOR U23727 ( .A(n23265), .B(n23264), .Z(n23226) );
  XNOR U23728 ( .A(n23227), .B(n23226), .Z(n23228) );
  XOR U23729 ( .A(n23229), .B(n23228), .Z(n23493) );
  XNOR U23730 ( .A(n23492), .B(n23493), .Z(n23499) );
  NANDN U23731 ( .A(n23186), .B(n23185), .Z(n23190) );
  OR U23732 ( .A(n23188), .B(n23187), .Z(n23189) );
  AND U23733 ( .A(n23190), .B(n23189), .Z(n23497) );
  NANDN U23734 ( .A(n23192), .B(n23191), .Z(n23196) );
  NANDN U23735 ( .A(n23194), .B(n23193), .Z(n23195) );
  AND U23736 ( .A(n23196), .B(n23195), .Z(n23496) );
  XNOR U23737 ( .A(n23497), .B(n23496), .Z(n23498) );
  XOR U23738 ( .A(n23499), .B(n23498), .Z(n23221) );
  NANDN U23739 ( .A(n23198), .B(n23197), .Z(n23202) );
  OR U23740 ( .A(n23200), .B(n23199), .Z(n23201) );
  NAND U23741 ( .A(n23202), .B(n23201), .Z(n23220) );
  XNOR U23742 ( .A(n23221), .B(n23220), .Z(n23222) );
  NANDN U23743 ( .A(n23204), .B(n23203), .Z(n23208) );
  OR U23744 ( .A(n23206), .B(n23205), .Z(n23207) );
  NAND U23745 ( .A(n23208), .B(n23207), .Z(n23223) );
  XNOR U23746 ( .A(n23222), .B(n23223), .Z(n23214) );
  XNOR U23747 ( .A(n23215), .B(n23214), .Z(n23216) );
  XNOR U23748 ( .A(n23217), .B(n23216), .Z(n23502) );
  XNOR U23749 ( .A(sreg[174]), .B(n23502), .Z(n23504) );
  NANDN U23750 ( .A(sreg[173]), .B(n23209), .Z(n23213) );
  NAND U23751 ( .A(n23211), .B(n23210), .Z(n23212) );
  NAND U23752 ( .A(n23213), .B(n23212), .Z(n23503) );
  XNOR U23753 ( .A(n23504), .B(n23503), .Z(c[174]) );
  NANDN U23754 ( .A(n23215), .B(n23214), .Z(n23219) );
  NANDN U23755 ( .A(n23217), .B(n23216), .Z(n23218) );
  AND U23756 ( .A(n23219), .B(n23218), .Z(n23510) );
  NANDN U23757 ( .A(n23221), .B(n23220), .Z(n23225) );
  NANDN U23758 ( .A(n23223), .B(n23222), .Z(n23224) );
  AND U23759 ( .A(n23225), .B(n23224), .Z(n23508) );
  NANDN U23760 ( .A(n23227), .B(n23226), .Z(n23231) );
  NANDN U23761 ( .A(n23229), .B(n23228), .Z(n23230) );
  AND U23762 ( .A(n23231), .B(n23230), .Z(n23790) );
  NANDN U23763 ( .A(n23233), .B(n23232), .Z(n23237) );
  NANDN U23764 ( .A(n23235), .B(n23234), .Z(n23236) );
  NAND U23765 ( .A(n23237), .B(n23236), .Z(n23789) );
  XNOR U23766 ( .A(n23790), .B(n23789), .Z(n23792) );
  NANDN U23767 ( .A(n23239), .B(n23238), .Z(n23243) );
  OR U23768 ( .A(n23241), .B(n23240), .Z(n23242) );
  AND U23769 ( .A(n23243), .B(n23242), .Z(n23527) );
  NANDN U23770 ( .A(n23245), .B(n23244), .Z(n23249) );
  NANDN U23771 ( .A(n23247), .B(n23246), .Z(n23248) );
  AND U23772 ( .A(n23249), .B(n23248), .Z(n23526) );
  NANDN U23773 ( .A(n23251), .B(n23250), .Z(n23255) );
  OR U23774 ( .A(n23253), .B(n23252), .Z(n23254) );
  AND U23775 ( .A(n23255), .B(n23254), .Z(n23525) );
  XOR U23776 ( .A(n23526), .B(n23525), .Z(n23528) );
  XOR U23777 ( .A(n23527), .B(n23528), .Z(n23784) );
  NANDN U23778 ( .A(n23257), .B(n23256), .Z(n23261) );
  OR U23779 ( .A(n23259), .B(n23258), .Z(n23260) );
  AND U23780 ( .A(n23261), .B(n23260), .Z(n23783) );
  XNOR U23781 ( .A(n23784), .B(n23783), .Z(n23785) );
  NANDN U23782 ( .A(n23263), .B(n23262), .Z(n23267) );
  NANDN U23783 ( .A(n23265), .B(n23264), .Z(n23266) );
  AND U23784 ( .A(n23267), .B(n23266), .Z(n23522) );
  NANDN U23785 ( .A(n23269), .B(n23268), .Z(n23273) );
  NAND U23786 ( .A(n23271), .B(n23270), .Z(n23272) );
  AND U23787 ( .A(n23273), .B(n23272), .Z(n23551) );
  NANDN U23788 ( .A(n23275), .B(n23274), .Z(n23279) );
  NANDN U23789 ( .A(n23277), .B(n23276), .Z(n23278) );
  AND U23790 ( .A(n23279), .B(n23278), .Z(n23545) );
  NANDN U23791 ( .A(n23281), .B(n23280), .Z(n23285) );
  NANDN U23792 ( .A(n23283), .B(n23282), .Z(n23284) );
  AND U23793 ( .A(n23285), .B(n23284), .Z(n23544) );
  NANDN U23794 ( .A(n33875), .B(n23286), .Z(n23288) );
  XOR U23795 ( .A(b[25]), .B(a[87]), .Z(n23579) );
  NANDN U23796 ( .A(n33994), .B(n23579), .Z(n23287) );
  AND U23797 ( .A(n23288), .B(n23287), .Z(n23773) );
  NANDN U23798 ( .A(n32013), .B(n23289), .Z(n23291) );
  XOR U23799 ( .A(a[95]), .B(b[17]), .Z(n23582) );
  NANDN U23800 ( .A(n32292), .B(n23582), .Z(n23290) );
  AND U23801 ( .A(n23291), .B(n23290), .Z(n23772) );
  NANDN U23802 ( .A(n31536), .B(n23292), .Z(n23294) );
  XOR U23803 ( .A(a[97]), .B(b[15]), .Z(n23585) );
  NANDN U23804 ( .A(n31925), .B(n23585), .Z(n23293) );
  NAND U23805 ( .A(n23294), .B(n23293), .Z(n23771) );
  XOR U23806 ( .A(n23772), .B(n23771), .Z(n23774) );
  XOR U23807 ( .A(n23773), .B(n23774), .Z(n23721) );
  NANDN U23808 ( .A(n37526), .B(n23295), .Z(n23297) );
  XOR U23809 ( .A(b[51]), .B(a[61]), .Z(n23588) );
  NANDN U23810 ( .A(n37605), .B(n23588), .Z(n23296) );
  AND U23811 ( .A(n23297), .B(n23296), .Z(n23752) );
  NANDN U23812 ( .A(n37705), .B(n23298), .Z(n23300) );
  XOR U23813 ( .A(b[53]), .B(a[59]), .Z(n23591) );
  NANDN U23814 ( .A(n37778), .B(n23591), .Z(n23299) );
  AND U23815 ( .A(n23300), .B(n23299), .Z(n23751) );
  NANDN U23816 ( .A(n36210), .B(n23301), .Z(n23303) );
  XOR U23817 ( .A(b[39]), .B(a[73]), .Z(n23594) );
  NANDN U23818 ( .A(n36347), .B(n23594), .Z(n23302) );
  NAND U23819 ( .A(n23303), .B(n23302), .Z(n23750) );
  XOR U23820 ( .A(n23751), .B(n23750), .Z(n23753) );
  XNOR U23821 ( .A(n23752), .B(n23753), .Z(n23720) );
  XNOR U23822 ( .A(n23721), .B(n23720), .Z(n23723) );
  NANDN U23823 ( .A(n23305), .B(n23304), .Z(n23309) );
  OR U23824 ( .A(n23307), .B(n23306), .Z(n23308) );
  AND U23825 ( .A(n23309), .B(n23308), .Z(n23722) );
  XOR U23826 ( .A(n23723), .B(n23722), .Z(n23570) );
  NANDN U23827 ( .A(n23311), .B(n23310), .Z(n23315) );
  OR U23828 ( .A(n23313), .B(n23312), .Z(n23314) );
  AND U23829 ( .A(n23315), .B(n23314), .Z(n23568) );
  NANDN U23830 ( .A(n23317), .B(n23316), .Z(n23321) );
  NANDN U23831 ( .A(n23319), .B(n23318), .Z(n23320) );
  NAND U23832 ( .A(n23321), .B(n23320), .Z(n23567) );
  XNOR U23833 ( .A(n23568), .B(n23567), .Z(n23569) );
  XNOR U23834 ( .A(n23570), .B(n23569), .Z(n23543) );
  XOR U23835 ( .A(n23544), .B(n23543), .Z(n23546) );
  XOR U23836 ( .A(n23545), .B(n23546), .Z(n23550) );
  NANDN U23837 ( .A(n29499), .B(n23322), .Z(n23324) );
  XOR U23838 ( .A(a[105]), .B(b[7]), .Z(n23645) );
  NANDN U23839 ( .A(n29735), .B(n23645), .Z(n23323) );
  AND U23840 ( .A(n23324), .B(n23323), .Z(n23605) );
  NANDN U23841 ( .A(n37857), .B(n23325), .Z(n23327) );
  XOR U23842 ( .A(b[55]), .B(a[57]), .Z(n23648) );
  NANDN U23843 ( .A(n37911), .B(n23648), .Z(n23326) );
  AND U23844 ( .A(n23327), .B(n23326), .Z(n23604) );
  NANDN U23845 ( .A(n35611), .B(n23328), .Z(n23330) );
  XOR U23846 ( .A(b[35]), .B(a[77]), .Z(n23651) );
  NANDN U23847 ( .A(n35801), .B(n23651), .Z(n23329) );
  NAND U23848 ( .A(n23330), .B(n23329), .Z(n23603) );
  XOR U23849 ( .A(n23604), .B(n23603), .Z(n23606) );
  XOR U23850 ( .A(n23605), .B(n23606), .Z(n23667) );
  NANDN U23851 ( .A(n23332), .B(n23331), .Z(n23336) );
  OR U23852 ( .A(n23334), .B(n23333), .Z(n23335) );
  AND U23853 ( .A(n23336), .B(n23335), .Z(n23666) );
  XNOR U23854 ( .A(n23667), .B(n23666), .Z(n23668) );
  NANDN U23855 ( .A(n23338), .B(n23337), .Z(n23342) );
  OR U23856 ( .A(n23340), .B(n23339), .Z(n23341) );
  NAND U23857 ( .A(n23342), .B(n23341), .Z(n23669) );
  XNOR U23858 ( .A(n23668), .B(n23669), .Z(n23539) );
  NANDN U23859 ( .A(n23344), .B(n23343), .Z(n23348) );
  NANDN U23860 ( .A(n23346), .B(n23345), .Z(n23347) );
  AND U23861 ( .A(n23348), .B(n23347), .Z(n23538) );
  NANDN U23862 ( .A(n211), .B(n23349), .Z(n23351) );
  XOR U23863 ( .A(b[47]), .B(a[65]), .Z(n23621) );
  NANDN U23864 ( .A(n37172), .B(n23621), .Z(n23350) );
  AND U23865 ( .A(n23351), .B(n23350), .Z(n23662) );
  NANDN U23866 ( .A(n210), .B(n23352), .Z(n23354) );
  XOR U23867 ( .A(a[103]), .B(b[9]), .Z(n23624) );
  NANDN U23868 ( .A(n30267), .B(n23624), .Z(n23353) );
  AND U23869 ( .A(n23354), .B(n23353), .Z(n23661) );
  NANDN U23870 ( .A(n212), .B(n23355), .Z(n23357) );
  XOR U23871 ( .A(b[49]), .B(a[63]), .Z(n23627) );
  NANDN U23872 ( .A(n37432), .B(n23627), .Z(n23356) );
  NAND U23873 ( .A(n23357), .B(n23356), .Z(n23660) );
  XOR U23874 ( .A(n23661), .B(n23660), .Z(n23663) );
  XOR U23875 ( .A(n23662), .B(n23663), .Z(n23727) );
  NANDN U23876 ( .A(n36742), .B(n23358), .Z(n23360) );
  XOR U23877 ( .A(b[43]), .B(a[69]), .Z(n23630) );
  NANDN U23878 ( .A(n36891), .B(n23630), .Z(n23359) );
  AND U23879 ( .A(n23360), .B(n23359), .Z(n23641) );
  NANDN U23880 ( .A(n36991), .B(n23361), .Z(n23363) );
  XOR U23881 ( .A(b[45]), .B(a[67]), .Z(n23633) );
  NANDN U23882 ( .A(n37083), .B(n23633), .Z(n23362) );
  AND U23883 ( .A(n23363), .B(n23362), .Z(n23640) );
  NANDN U23884 ( .A(n30482), .B(n23364), .Z(n23366) );
  XOR U23885 ( .A(a[101]), .B(b[11]), .Z(n23636) );
  NANDN U23886 ( .A(n30891), .B(n23636), .Z(n23365) );
  NAND U23887 ( .A(n23366), .B(n23365), .Z(n23639) );
  XOR U23888 ( .A(n23640), .B(n23639), .Z(n23642) );
  XNOR U23889 ( .A(n23641), .B(n23642), .Z(n23726) );
  XNOR U23890 ( .A(n23727), .B(n23726), .Z(n23728) );
  NANDN U23891 ( .A(n23368), .B(n23367), .Z(n23372) );
  OR U23892 ( .A(n23370), .B(n23369), .Z(n23371) );
  NAND U23893 ( .A(n23372), .B(n23371), .Z(n23729) );
  XNOR U23894 ( .A(n23728), .B(n23729), .Z(n23537) );
  XOR U23895 ( .A(n23538), .B(n23537), .Z(n23540) );
  XNOR U23896 ( .A(n23539), .B(n23540), .Z(n23549) );
  XOR U23897 ( .A(n23550), .B(n23549), .Z(n23552) );
  XOR U23898 ( .A(n23551), .B(n23552), .Z(n23520) );
  NANDN U23899 ( .A(n23374), .B(n23373), .Z(n23378) );
  NANDN U23900 ( .A(n23376), .B(n23375), .Z(n23377) );
  AND U23901 ( .A(n23378), .B(n23377), .Z(n23533) );
  NANDN U23902 ( .A(n23380), .B(n23379), .Z(n23384) );
  NANDN U23903 ( .A(n23382), .B(n23381), .Z(n23383) );
  AND U23904 ( .A(n23384), .B(n23383), .Z(n23532) );
  NANDN U23905 ( .A(n23386), .B(n23385), .Z(n23390) );
  NAND U23906 ( .A(n23388), .B(n23387), .Z(n23389) );
  AND U23907 ( .A(n23390), .B(n23389), .Z(n23531) );
  XOR U23908 ( .A(n23532), .B(n23531), .Z(n23534) );
  XOR U23909 ( .A(n23533), .B(n23534), .Z(n23558) );
  NANDN U23910 ( .A(n23392), .B(n23391), .Z(n23396) );
  NANDN U23911 ( .A(n23394), .B(n23393), .Z(n23395) );
  AND U23912 ( .A(n23396), .B(n23395), .Z(n23679) );
  NANDN U23913 ( .A(n23398), .B(n23397), .Z(n23402) );
  OR U23914 ( .A(n23400), .B(n23399), .Z(n23401) );
  NAND U23915 ( .A(n23402), .B(n23401), .Z(n23678) );
  XNOR U23916 ( .A(n23679), .B(n23678), .Z(n23681) );
  NANDN U23917 ( .A(n23404), .B(n23403), .Z(n23408) );
  OR U23918 ( .A(n23406), .B(n23405), .Z(n23407) );
  AND U23919 ( .A(n23408), .B(n23407), .Z(n23576) );
  NAND U23920 ( .A(b[0]), .B(a[111]), .Z(n23409) );
  XNOR U23921 ( .A(b[1]), .B(n23409), .Z(n23411) );
  NANDN U23922 ( .A(b[0]), .B(a[110]), .Z(n23410) );
  NAND U23923 ( .A(n23411), .B(n23410), .Z(n23612) );
  NANDN U23924 ( .A(n38278), .B(n23412), .Z(n23414) );
  XOR U23925 ( .A(b[63]), .B(a[49]), .Z(n23705) );
  NANDN U23926 ( .A(n38279), .B(n23705), .Z(n23413) );
  AND U23927 ( .A(n23414), .B(n23413), .Z(n23610) );
  NANDN U23928 ( .A(n35260), .B(n23415), .Z(n23417) );
  XOR U23929 ( .A(b[33]), .B(a[79]), .Z(n23708) );
  NANDN U23930 ( .A(n35456), .B(n23708), .Z(n23416) );
  NAND U23931 ( .A(n23417), .B(n23416), .Z(n23609) );
  XNOR U23932 ( .A(n23610), .B(n23609), .Z(n23611) );
  XNOR U23933 ( .A(n23612), .B(n23611), .Z(n23573) );
  NANDN U23934 ( .A(n37974), .B(n23418), .Z(n23420) );
  XOR U23935 ( .A(b[57]), .B(a[55]), .Z(n23711) );
  NANDN U23936 ( .A(n38031), .B(n23711), .Z(n23419) );
  AND U23937 ( .A(n23420), .B(n23419), .Z(n23687) );
  NANDN U23938 ( .A(n38090), .B(n23421), .Z(n23423) );
  XOR U23939 ( .A(b[59]), .B(a[53]), .Z(n23714) );
  NANDN U23940 ( .A(n38130), .B(n23714), .Z(n23422) );
  AND U23941 ( .A(n23423), .B(n23422), .Z(n23685) );
  NANDN U23942 ( .A(n36480), .B(n23424), .Z(n23426) );
  XOR U23943 ( .A(b[41]), .B(a[71]), .Z(n23717) );
  NANDN U23944 ( .A(n36594), .B(n23717), .Z(n23425) );
  NAND U23945 ( .A(n23426), .B(n23425), .Z(n23684) );
  XNOR U23946 ( .A(n23685), .B(n23684), .Z(n23686) );
  XOR U23947 ( .A(n23687), .B(n23686), .Z(n23574) );
  XNOR U23948 ( .A(n23573), .B(n23574), .Z(n23575) );
  XNOR U23949 ( .A(n23576), .B(n23575), .Z(n23680) );
  XOR U23950 ( .A(n23681), .B(n23680), .Z(n23562) );
  NANDN U23951 ( .A(n23428), .B(n23427), .Z(n23432) );
  NAND U23952 ( .A(n23430), .B(n23429), .Z(n23431) );
  NAND U23953 ( .A(n23432), .B(n23431), .Z(n23561) );
  XNOR U23954 ( .A(n23562), .B(n23561), .Z(n23564) );
  NANDN U23955 ( .A(n23434), .B(n23433), .Z(n23438) );
  NANDN U23956 ( .A(n23436), .B(n23435), .Z(n23437) );
  AND U23957 ( .A(n23438), .B(n23437), .Z(n23780) );
  NANDN U23958 ( .A(n34223), .B(n23439), .Z(n23441) );
  XOR U23959 ( .A(b[27]), .B(a[85]), .Z(n23732) );
  NANDN U23960 ( .A(n34458), .B(n23732), .Z(n23440) );
  AND U23961 ( .A(n23441), .B(n23440), .Z(n23599) );
  NANDN U23962 ( .A(n34634), .B(n23442), .Z(n23444) );
  XOR U23963 ( .A(b[29]), .B(a[83]), .Z(n23735) );
  NANDN U23964 ( .A(n34722), .B(n23735), .Z(n23443) );
  AND U23965 ( .A(n23444), .B(n23443), .Z(n23598) );
  NANDN U23966 ( .A(n31055), .B(n23445), .Z(n23447) );
  XOR U23967 ( .A(a[99]), .B(b[13]), .Z(n23738) );
  NANDN U23968 ( .A(n31293), .B(n23738), .Z(n23446) );
  NAND U23969 ( .A(n23447), .B(n23446), .Z(n23597) );
  XOR U23970 ( .A(n23598), .B(n23597), .Z(n23600) );
  XOR U23971 ( .A(n23599), .B(n23600), .Z(n23673) );
  NANDN U23972 ( .A(n28889), .B(n23448), .Z(n23450) );
  XOR U23973 ( .A(a[107]), .B(b[5]), .Z(n23741) );
  NANDN U23974 ( .A(n29138), .B(n23741), .Z(n23449) );
  AND U23975 ( .A(n23450), .B(n23449), .Z(n23692) );
  NANDN U23976 ( .A(n209), .B(n23451), .Z(n23453) );
  XOR U23977 ( .A(a[109]), .B(b[3]), .Z(n23744) );
  NANDN U23978 ( .A(n28941), .B(n23744), .Z(n23452) );
  AND U23979 ( .A(n23453), .B(n23452), .Z(n23691) );
  NANDN U23980 ( .A(n35936), .B(n23454), .Z(n23456) );
  XOR U23981 ( .A(b[37]), .B(a[75]), .Z(n23747) );
  NANDN U23982 ( .A(n36047), .B(n23747), .Z(n23455) );
  NAND U23983 ( .A(n23456), .B(n23455), .Z(n23690) );
  XOR U23984 ( .A(n23691), .B(n23690), .Z(n23693) );
  XNOR U23985 ( .A(n23692), .B(n23693), .Z(n23672) );
  XNOR U23986 ( .A(n23673), .B(n23672), .Z(n23674) );
  NANDN U23987 ( .A(n23458), .B(n23457), .Z(n23462) );
  OR U23988 ( .A(n23460), .B(n23459), .Z(n23461) );
  NAND U23989 ( .A(n23462), .B(n23461), .Z(n23675) );
  XNOR U23990 ( .A(n23674), .B(n23675), .Z(n23777) );
  NANDN U23991 ( .A(n32996), .B(n23463), .Z(n23465) );
  XOR U23992 ( .A(a[91]), .B(b[21]), .Z(n23756) );
  NANDN U23993 ( .A(n33271), .B(n23756), .Z(n23464) );
  AND U23994 ( .A(n23465), .B(n23464), .Z(n23698) );
  NANDN U23995 ( .A(n33866), .B(n23466), .Z(n23468) );
  XOR U23996 ( .A(b[23]), .B(a[89]), .Z(n23759) );
  NANDN U23997 ( .A(n33644), .B(n23759), .Z(n23467) );
  AND U23998 ( .A(n23468), .B(n23467), .Z(n23697) );
  NANDN U23999 ( .A(n32483), .B(n23469), .Z(n23471) );
  XOR U24000 ( .A(a[93]), .B(b[19]), .Z(n23762) );
  NANDN U24001 ( .A(n32823), .B(n23762), .Z(n23470) );
  NAND U24002 ( .A(n23471), .B(n23470), .Z(n23696) );
  XOR U24003 ( .A(n23697), .B(n23696), .Z(n23699) );
  XOR U24004 ( .A(n23698), .B(n23699), .Z(n23616) );
  NANDN U24005 ( .A(n34909), .B(n23472), .Z(n23474) );
  XOR U24006 ( .A(b[31]), .B(a[81]), .Z(n23765) );
  NANDN U24007 ( .A(n35145), .B(n23765), .Z(n23473) );
  AND U24008 ( .A(n23474), .B(n23473), .Z(n23656) );
  NANDN U24009 ( .A(n38247), .B(n23475), .Z(n23477) );
  XOR U24010 ( .A(b[61]), .B(a[51]), .Z(n23768) );
  NANDN U24011 ( .A(n38248), .B(n23768), .Z(n23476) );
  AND U24012 ( .A(n23477), .B(n23476), .Z(n23655) );
  AND U24013 ( .A(b[63]), .B(a[47]), .Z(n23654) );
  XOR U24014 ( .A(n23655), .B(n23654), .Z(n23657) );
  XNOR U24015 ( .A(n23656), .B(n23657), .Z(n23615) );
  XNOR U24016 ( .A(n23616), .B(n23615), .Z(n23617) );
  NANDN U24017 ( .A(n23479), .B(n23478), .Z(n23483) );
  OR U24018 ( .A(n23481), .B(n23480), .Z(n23482) );
  NAND U24019 ( .A(n23483), .B(n23482), .Z(n23618) );
  XOR U24020 ( .A(n23617), .B(n23618), .Z(n23778) );
  XNOR U24021 ( .A(n23777), .B(n23778), .Z(n23779) );
  XNOR U24022 ( .A(n23780), .B(n23779), .Z(n23563) );
  XOR U24023 ( .A(n23564), .B(n23563), .Z(n23556) );
  NANDN U24024 ( .A(n23485), .B(n23484), .Z(n23489) );
  NANDN U24025 ( .A(n23487), .B(n23486), .Z(n23488) );
  AND U24026 ( .A(n23489), .B(n23488), .Z(n23555) );
  XNOR U24027 ( .A(n23556), .B(n23555), .Z(n23557) );
  XNOR U24028 ( .A(n23558), .B(n23557), .Z(n23519) );
  XNOR U24029 ( .A(n23520), .B(n23519), .Z(n23521) );
  XOR U24030 ( .A(n23522), .B(n23521), .Z(n23786) );
  XNOR U24031 ( .A(n23785), .B(n23786), .Z(n23791) );
  XOR U24032 ( .A(n23792), .B(n23791), .Z(n23514) );
  NANDN U24033 ( .A(n23491), .B(n23490), .Z(n23495) );
  NANDN U24034 ( .A(n23493), .B(n23492), .Z(n23494) );
  AND U24035 ( .A(n23495), .B(n23494), .Z(n23513) );
  XNOR U24036 ( .A(n23514), .B(n23513), .Z(n23515) );
  NANDN U24037 ( .A(n23497), .B(n23496), .Z(n23501) );
  NAND U24038 ( .A(n23499), .B(n23498), .Z(n23500) );
  NAND U24039 ( .A(n23501), .B(n23500), .Z(n23516) );
  XNOR U24040 ( .A(n23515), .B(n23516), .Z(n23507) );
  XNOR U24041 ( .A(n23508), .B(n23507), .Z(n23509) );
  XNOR U24042 ( .A(n23510), .B(n23509), .Z(n23795) );
  XNOR U24043 ( .A(sreg[175]), .B(n23795), .Z(n23797) );
  NANDN U24044 ( .A(sreg[174]), .B(n23502), .Z(n23506) );
  NAND U24045 ( .A(n23504), .B(n23503), .Z(n23505) );
  NAND U24046 ( .A(n23506), .B(n23505), .Z(n23796) );
  XNOR U24047 ( .A(n23797), .B(n23796), .Z(c[175]) );
  NANDN U24048 ( .A(n23508), .B(n23507), .Z(n23512) );
  NANDN U24049 ( .A(n23510), .B(n23509), .Z(n23511) );
  AND U24050 ( .A(n23512), .B(n23511), .Z(n23803) );
  NANDN U24051 ( .A(n23514), .B(n23513), .Z(n23518) );
  NANDN U24052 ( .A(n23516), .B(n23515), .Z(n23517) );
  AND U24053 ( .A(n23518), .B(n23517), .Z(n23801) );
  NANDN U24054 ( .A(n23520), .B(n23519), .Z(n23524) );
  NANDN U24055 ( .A(n23522), .B(n23521), .Z(n23523) );
  AND U24056 ( .A(n23524), .B(n23523), .Z(n23813) );
  NANDN U24057 ( .A(n23526), .B(n23525), .Z(n23530) );
  OR U24058 ( .A(n23528), .B(n23527), .Z(n23529) );
  AND U24059 ( .A(n23530), .B(n23529), .Z(n23812) );
  XNOR U24060 ( .A(n23813), .B(n23812), .Z(n23815) );
  NANDN U24061 ( .A(n23532), .B(n23531), .Z(n23536) );
  OR U24062 ( .A(n23534), .B(n23533), .Z(n23535) );
  AND U24063 ( .A(n23536), .B(n23535), .Z(n24084) );
  NANDN U24064 ( .A(n23538), .B(n23537), .Z(n23542) );
  NANDN U24065 ( .A(n23540), .B(n23539), .Z(n23541) );
  AND U24066 ( .A(n23542), .B(n23541), .Z(n24083) );
  NANDN U24067 ( .A(n23544), .B(n23543), .Z(n23548) );
  OR U24068 ( .A(n23546), .B(n23545), .Z(n23547) );
  AND U24069 ( .A(n23548), .B(n23547), .Z(n24082) );
  XOR U24070 ( .A(n24083), .B(n24082), .Z(n24085) );
  XOR U24071 ( .A(n24084), .B(n24085), .Z(n23819) );
  NANDN U24072 ( .A(n23550), .B(n23549), .Z(n23554) );
  OR U24073 ( .A(n23552), .B(n23551), .Z(n23553) );
  AND U24074 ( .A(n23554), .B(n23553), .Z(n23818) );
  XNOR U24075 ( .A(n23819), .B(n23818), .Z(n23820) );
  NANDN U24076 ( .A(n23556), .B(n23555), .Z(n23560) );
  NANDN U24077 ( .A(n23558), .B(n23557), .Z(n23559) );
  AND U24078 ( .A(n23560), .B(n23559), .Z(n24079) );
  NANDN U24079 ( .A(n23562), .B(n23561), .Z(n23566) );
  NAND U24080 ( .A(n23564), .B(n23563), .Z(n23565) );
  AND U24081 ( .A(n23566), .B(n23565), .Z(n24054) );
  NANDN U24082 ( .A(n23568), .B(n23567), .Z(n23572) );
  NANDN U24083 ( .A(n23570), .B(n23569), .Z(n23571) );
  AND U24084 ( .A(n23572), .B(n23571), .Z(n24072) );
  NANDN U24085 ( .A(n23574), .B(n23573), .Z(n23578) );
  NANDN U24086 ( .A(n23576), .B(n23575), .Z(n23577) );
  AND U24087 ( .A(n23578), .B(n23577), .Z(n24071) );
  NANDN U24088 ( .A(n33875), .B(n23579), .Z(n23581) );
  XOR U24089 ( .A(b[25]), .B(a[88]), .Z(n23848) );
  NANDN U24090 ( .A(n33994), .B(n23848), .Z(n23580) );
  AND U24091 ( .A(n23581), .B(n23580), .Z(n23976) );
  NANDN U24092 ( .A(n32013), .B(n23582), .Z(n23584) );
  XOR U24093 ( .A(a[96]), .B(b[17]), .Z(n23851) );
  NANDN U24094 ( .A(n32292), .B(n23851), .Z(n23583) );
  AND U24095 ( .A(n23584), .B(n23583), .Z(n23975) );
  NANDN U24096 ( .A(n31536), .B(n23585), .Z(n23587) );
  XOR U24097 ( .A(a[98]), .B(b[15]), .Z(n23854) );
  NANDN U24098 ( .A(n31925), .B(n23854), .Z(n23586) );
  NAND U24099 ( .A(n23587), .B(n23586), .Z(n23974) );
  XOR U24100 ( .A(n23975), .B(n23974), .Z(n23977) );
  XOR U24101 ( .A(n23976), .B(n23977), .Z(n24041) );
  NANDN U24102 ( .A(n37526), .B(n23588), .Z(n23590) );
  XOR U24103 ( .A(b[51]), .B(a[62]), .Z(n23857) );
  NANDN U24104 ( .A(n37605), .B(n23857), .Z(n23589) );
  AND U24105 ( .A(n23590), .B(n23589), .Z(n24000) );
  NANDN U24106 ( .A(n37705), .B(n23591), .Z(n23593) );
  XOR U24107 ( .A(b[53]), .B(a[60]), .Z(n23860) );
  NANDN U24108 ( .A(n37778), .B(n23860), .Z(n23592) );
  AND U24109 ( .A(n23593), .B(n23592), .Z(n23999) );
  NANDN U24110 ( .A(n36210), .B(n23594), .Z(n23596) );
  XOR U24111 ( .A(b[39]), .B(a[74]), .Z(n23863) );
  NANDN U24112 ( .A(n36347), .B(n23863), .Z(n23595) );
  NAND U24113 ( .A(n23596), .B(n23595), .Z(n23998) );
  XOR U24114 ( .A(n23999), .B(n23998), .Z(n24001) );
  XNOR U24115 ( .A(n24000), .B(n24001), .Z(n24040) );
  XNOR U24116 ( .A(n24041), .B(n24040), .Z(n24043) );
  NANDN U24117 ( .A(n23598), .B(n23597), .Z(n23602) );
  OR U24118 ( .A(n23600), .B(n23599), .Z(n23601) );
  AND U24119 ( .A(n23602), .B(n23601), .Z(n24042) );
  XOR U24120 ( .A(n24043), .B(n24042), .Z(n23839) );
  NANDN U24121 ( .A(n23604), .B(n23603), .Z(n23608) );
  OR U24122 ( .A(n23606), .B(n23605), .Z(n23607) );
  AND U24123 ( .A(n23608), .B(n23607), .Z(n23837) );
  NANDN U24124 ( .A(n23610), .B(n23609), .Z(n23614) );
  NANDN U24125 ( .A(n23612), .B(n23611), .Z(n23613) );
  NAND U24126 ( .A(n23614), .B(n23613), .Z(n23836) );
  XNOR U24127 ( .A(n23837), .B(n23836), .Z(n23838) );
  XNOR U24128 ( .A(n23839), .B(n23838), .Z(n24070) );
  XOR U24129 ( .A(n24071), .B(n24070), .Z(n24073) );
  XOR U24130 ( .A(n24072), .B(n24073), .Z(n24053) );
  NANDN U24131 ( .A(n23616), .B(n23615), .Z(n23620) );
  NANDN U24132 ( .A(n23618), .B(n23617), .Z(n23619) );
  AND U24133 ( .A(n23620), .B(n23619), .Z(n24065) );
  NANDN U24134 ( .A(n211), .B(n23621), .Z(n23623) );
  XOR U24135 ( .A(b[47]), .B(a[66]), .Z(n23890) );
  NANDN U24136 ( .A(n37172), .B(n23890), .Z(n23622) );
  AND U24137 ( .A(n23623), .B(n23622), .Z(n23931) );
  NANDN U24138 ( .A(n210), .B(n23624), .Z(n23626) );
  XOR U24139 ( .A(a[104]), .B(b[9]), .Z(n23893) );
  NANDN U24140 ( .A(n30267), .B(n23893), .Z(n23625) );
  AND U24141 ( .A(n23626), .B(n23625), .Z(n23930) );
  NANDN U24142 ( .A(n212), .B(n23627), .Z(n23629) );
  XOR U24143 ( .A(b[49]), .B(a[64]), .Z(n23896) );
  NANDN U24144 ( .A(n37432), .B(n23896), .Z(n23628) );
  NAND U24145 ( .A(n23629), .B(n23628), .Z(n23929) );
  XOR U24146 ( .A(n23930), .B(n23929), .Z(n23932) );
  XOR U24147 ( .A(n23931), .B(n23932), .Z(n23954) );
  NANDN U24148 ( .A(n36742), .B(n23630), .Z(n23632) );
  XOR U24149 ( .A(b[43]), .B(a[70]), .Z(n23899) );
  NANDN U24150 ( .A(n36891), .B(n23899), .Z(n23631) );
  AND U24151 ( .A(n23632), .B(n23631), .Z(n23910) );
  NANDN U24152 ( .A(n36991), .B(n23633), .Z(n23635) );
  XOR U24153 ( .A(b[45]), .B(a[68]), .Z(n23902) );
  NANDN U24154 ( .A(n37083), .B(n23902), .Z(n23634) );
  AND U24155 ( .A(n23635), .B(n23634), .Z(n23909) );
  NANDN U24156 ( .A(n30482), .B(n23636), .Z(n23638) );
  XOR U24157 ( .A(a[102]), .B(b[11]), .Z(n23905) );
  NANDN U24158 ( .A(n30891), .B(n23905), .Z(n23637) );
  NAND U24159 ( .A(n23638), .B(n23637), .Z(n23908) );
  XOR U24160 ( .A(n23909), .B(n23908), .Z(n23911) );
  XNOR U24161 ( .A(n23910), .B(n23911), .Z(n23953) );
  XNOR U24162 ( .A(n23954), .B(n23953), .Z(n23955) );
  NANDN U24163 ( .A(n23640), .B(n23639), .Z(n23644) );
  OR U24164 ( .A(n23642), .B(n23641), .Z(n23643) );
  NAND U24165 ( .A(n23644), .B(n23643), .Z(n23956) );
  XNOR U24166 ( .A(n23955), .B(n23956), .Z(n24064) );
  XNOR U24167 ( .A(n24065), .B(n24064), .Z(n24066) );
  NANDN U24168 ( .A(n29499), .B(n23645), .Z(n23647) );
  XOR U24169 ( .A(a[106]), .B(b[7]), .Z(n23914) );
  NANDN U24170 ( .A(n29735), .B(n23914), .Z(n23646) );
  AND U24171 ( .A(n23647), .B(n23646), .Z(n23874) );
  NANDN U24172 ( .A(n37857), .B(n23648), .Z(n23650) );
  XOR U24173 ( .A(b[55]), .B(a[58]), .Z(n23917) );
  NANDN U24174 ( .A(n37911), .B(n23917), .Z(n23649) );
  AND U24175 ( .A(n23650), .B(n23649), .Z(n23873) );
  NANDN U24176 ( .A(n35611), .B(n23651), .Z(n23653) );
  XOR U24177 ( .A(b[35]), .B(a[78]), .Z(n23920) );
  NANDN U24178 ( .A(n35801), .B(n23920), .Z(n23652) );
  NAND U24179 ( .A(n23653), .B(n23652), .Z(n23872) );
  XOR U24180 ( .A(n23873), .B(n23872), .Z(n23875) );
  XOR U24181 ( .A(n23874), .B(n23875), .Z(n23936) );
  NANDN U24182 ( .A(n23655), .B(n23654), .Z(n23659) );
  OR U24183 ( .A(n23657), .B(n23656), .Z(n23658) );
  AND U24184 ( .A(n23659), .B(n23658), .Z(n23935) );
  XNOR U24185 ( .A(n23936), .B(n23935), .Z(n23937) );
  NANDN U24186 ( .A(n23661), .B(n23660), .Z(n23665) );
  OR U24187 ( .A(n23663), .B(n23662), .Z(n23664) );
  NAND U24188 ( .A(n23665), .B(n23664), .Z(n23938) );
  XOR U24189 ( .A(n23937), .B(n23938), .Z(n24067) );
  XNOR U24190 ( .A(n24066), .B(n24067), .Z(n24052) );
  XOR U24191 ( .A(n24053), .B(n24052), .Z(n24055) );
  XOR U24192 ( .A(n24054), .B(n24055), .Z(n24077) );
  NANDN U24193 ( .A(n23667), .B(n23666), .Z(n23671) );
  NANDN U24194 ( .A(n23669), .B(n23668), .Z(n23670) );
  AND U24195 ( .A(n23671), .B(n23670), .Z(n24060) );
  NANDN U24196 ( .A(n23673), .B(n23672), .Z(n23677) );
  NANDN U24197 ( .A(n23675), .B(n23674), .Z(n23676) );
  AND U24198 ( .A(n23677), .B(n23676), .Z(n24059) );
  NANDN U24199 ( .A(n23679), .B(n23678), .Z(n23683) );
  NAND U24200 ( .A(n23681), .B(n23680), .Z(n23682) );
  AND U24201 ( .A(n23683), .B(n23682), .Z(n24058) );
  XOR U24202 ( .A(n24059), .B(n24058), .Z(n24061) );
  XOR U24203 ( .A(n24060), .B(n24061), .Z(n23827) );
  NANDN U24204 ( .A(n23685), .B(n23684), .Z(n23689) );
  NANDN U24205 ( .A(n23687), .B(n23686), .Z(n23688) );
  AND U24206 ( .A(n23689), .B(n23688), .Z(n23948) );
  NANDN U24207 ( .A(n23691), .B(n23690), .Z(n23695) );
  OR U24208 ( .A(n23693), .B(n23692), .Z(n23694) );
  NAND U24209 ( .A(n23695), .B(n23694), .Z(n23947) );
  XNOR U24210 ( .A(n23948), .B(n23947), .Z(n23950) );
  NANDN U24211 ( .A(n23697), .B(n23696), .Z(n23701) );
  OR U24212 ( .A(n23699), .B(n23698), .Z(n23700) );
  AND U24213 ( .A(n23701), .B(n23700), .Z(n23845) );
  NAND U24214 ( .A(b[0]), .B(a[112]), .Z(n23702) );
  XNOR U24215 ( .A(b[1]), .B(n23702), .Z(n23704) );
  NANDN U24216 ( .A(b[0]), .B(a[111]), .Z(n23703) );
  NAND U24217 ( .A(n23704), .B(n23703), .Z(n23881) );
  NANDN U24218 ( .A(n38278), .B(n23705), .Z(n23707) );
  XOR U24219 ( .A(b[63]), .B(a[50]), .Z(n24025) );
  NANDN U24220 ( .A(n38279), .B(n24025), .Z(n23706) );
  AND U24221 ( .A(n23707), .B(n23706), .Z(n23879) );
  NANDN U24222 ( .A(n35260), .B(n23708), .Z(n23710) );
  XOR U24223 ( .A(b[33]), .B(a[80]), .Z(n24028) );
  NANDN U24224 ( .A(n35456), .B(n24028), .Z(n23709) );
  NAND U24225 ( .A(n23710), .B(n23709), .Z(n23878) );
  XNOR U24226 ( .A(n23879), .B(n23878), .Z(n23880) );
  XNOR U24227 ( .A(n23881), .B(n23880), .Z(n23842) );
  NANDN U24228 ( .A(n37974), .B(n23711), .Z(n23713) );
  XOR U24229 ( .A(b[57]), .B(a[56]), .Z(n24031) );
  NANDN U24230 ( .A(n38031), .B(n24031), .Z(n23712) );
  AND U24231 ( .A(n23713), .B(n23712), .Z(n24007) );
  NANDN U24232 ( .A(n38090), .B(n23714), .Z(n23716) );
  XOR U24233 ( .A(b[59]), .B(a[54]), .Z(n24034) );
  NANDN U24234 ( .A(n38130), .B(n24034), .Z(n23715) );
  AND U24235 ( .A(n23716), .B(n23715), .Z(n24005) );
  NANDN U24236 ( .A(n36480), .B(n23717), .Z(n23719) );
  XOR U24237 ( .A(b[41]), .B(a[72]), .Z(n24037) );
  NANDN U24238 ( .A(n36594), .B(n24037), .Z(n23718) );
  NAND U24239 ( .A(n23719), .B(n23718), .Z(n24004) );
  XNOR U24240 ( .A(n24005), .B(n24004), .Z(n24006) );
  XOR U24241 ( .A(n24007), .B(n24006), .Z(n23843) );
  XNOR U24242 ( .A(n23842), .B(n23843), .Z(n23844) );
  XNOR U24243 ( .A(n23845), .B(n23844), .Z(n23949) );
  XOR U24244 ( .A(n23950), .B(n23949), .Z(n23831) );
  NANDN U24245 ( .A(n23721), .B(n23720), .Z(n23725) );
  NAND U24246 ( .A(n23723), .B(n23722), .Z(n23724) );
  NAND U24247 ( .A(n23725), .B(n23724), .Z(n23830) );
  XNOR U24248 ( .A(n23831), .B(n23830), .Z(n23833) );
  NANDN U24249 ( .A(n23727), .B(n23726), .Z(n23731) );
  NANDN U24250 ( .A(n23729), .B(n23728), .Z(n23730) );
  AND U24251 ( .A(n23731), .B(n23730), .Z(n24049) );
  NANDN U24252 ( .A(n34223), .B(n23732), .Z(n23734) );
  XOR U24253 ( .A(b[27]), .B(a[86]), .Z(n23980) );
  NANDN U24254 ( .A(n34458), .B(n23980), .Z(n23733) );
  AND U24255 ( .A(n23734), .B(n23733), .Z(n23868) );
  NANDN U24256 ( .A(n34634), .B(n23735), .Z(n23737) );
  XOR U24257 ( .A(b[29]), .B(a[84]), .Z(n23983) );
  NANDN U24258 ( .A(n34722), .B(n23983), .Z(n23736) );
  AND U24259 ( .A(n23737), .B(n23736), .Z(n23867) );
  NANDN U24260 ( .A(n31055), .B(n23738), .Z(n23740) );
  XOR U24261 ( .A(a[100]), .B(b[13]), .Z(n23986) );
  NANDN U24262 ( .A(n31293), .B(n23986), .Z(n23739) );
  NAND U24263 ( .A(n23740), .B(n23739), .Z(n23866) );
  XOR U24264 ( .A(n23867), .B(n23866), .Z(n23869) );
  XOR U24265 ( .A(n23868), .B(n23869), .Z(n23942) );
  NANDN U24266 ( .A(n28889), .B(n23741), .Z(n23743) );
  XOR U24267 ( .A(a[108]), .B(b[5]), .Z(n23989) );
  NANDN U24268 ( .A(n29138), .B(n23989), .Z(n23742) );
  AND U24269 ( .A(n23743), .B(n23742), .Z(n24012) );
  NANDN U24270 ( .A(n209), .B(n23744), .Z(n23746) );
  XOR U24271 ( .A(a[110]), .B(b[3]), .Z(n23992) );
  NANDN U24272 ( .A(n28941), .B(n23992), .Z(n23745) );
  AND U24273 ( .A(n23746), .B(n23745), .Z(n24011) );
  NANDN U24274 ( .A(n35936), .B(n23747), .Z(n23749) );
  XOR U24275 ( .A(b[37]), .B(a[76]), .Z(n23995) );
  NANDN U24276 ( .A(n36047), .B(n23995), .Z(n23748) );
  NAND U24277 ( .A(n23749), .B(n23748), .Z(n24010) );
  XOR U24278 ( .A(n24011), .B(n24010), .Z(n24013) );
  XNOR U24279 ( .A(n24012), .B(n24013), .Z(n23941) );
  XNOR U24280 ( .A(n23942), .B(n23941), .Z(n23943) );
  NANDN U24281 ( .A(n23751), .B(n23750), .Z(n23755) );
  OR U24282 ( .A(n23753), .B(n23752), .Z(n23754) );
  NAND U24283 ( .A(n23755), .B(n23754), .Z(n23944) );
  XNOR U24284 ( .A(n23943), .B(n23944), .Z(n24046) );
  NANDN U24285 ( .A(n32996), .B(n23756), .Z(n23758) );
  XOR U24286 ( .A(a[92]), .B(b[21]), .Z(n23959) );
  NANDN U24287 ( .A(n33271), .B(n23959), .Z(n23757) );
  AND U24288 ( .A(n23758), .B(n23757), .Z(n24018) );
  NANDN U24289 ( .A(n33866), .B(n23759), .Z(n23761) );
  XOR U24290 ( .A(a[90]), .B(b[23]), .Z(n23962) );
  NANDN U24291 ( .A(n33644), .B(n23962), .Z(n23760) );
  AND U24292 ( .A(n23761), .B(n23760), .Z(n24017) );
  NANDN U24293 ( .A(n32483), .B(n23762), .Z(n23764) );
  XOR U24294 ( .A(a[94]), .B(b[19]), .Z(n23965) );
  NANDN U24295 ( .A(n32823), .B(n23965), .Z(n23763) );
  NAND U24296 ( .A(n23764), .B(n23763), .Z(n24016) );
  XOR U24297 ( .A(n24017), .B(n24016), .Z(n24019) );
  XOR U24298 ( .A(n24018), .B(n24019), .Z(n23885) );
  NANDN U24299 ( .A(n34909), .B(n23765), .Z(n23767) );
  XOR U24300 ( .A(b[31]), .B(a[82]), .Z(n23968) );
  NANDN U24301 ( .A(n35145), .B(n23968), .Z(n23766) );
  AND U24302 ( .A(n23767), .B(n23766), .Z(n23925) );
  NANDN U24303 ( .A(n38247), .B(n23768), .Z(n23770) );
  XOR U24304 ( .A(b[61]), .B(a[52]), .Z(n23971) );
  NANDN U24305 ( .A(n38248), .B(n23971), .Z(n23769) );
  AND U24306 ( .A(n23770), .B(n23769), .Z(n23924) );
  AND U24307 ( .A(b[63]), .B(a[48]), .Z(n23923) );
  XOR U24308 ( .A(n23924), .B(n23923), .Z(n23926) );
  XNOR U24309 ( .A(n23925), .B(n23926), .Z(n23884) );
  XNOR U24310 ( .A(n23885), .B(n23884), .Z(n23886) );
  NANDN U24311 ( .A(n23772), .B(n23771), .Z(n23776) );
  OR U24312 ( .A(n23774), .B(n23773), .Z(n23775) );
  NAND U24313 ( .A(n23776), .B(n23775), .Z(n23887) );
  XOR U24314 ( .A(n23886), .B(n23887), .Z(n24047) );
  XNOR U24315 ( .A(n24046), .B(n24047), .Z(n24048) );
  XNOR U24316 ( .A(n24049), .B(n24048), .Z(n23832) );
  XOR U24317 ( .A(n23833), .B(n23832), .Z(n23825) );
  NANDN U24318 ( .A(n23778), .B(n23777), .Z(n23782) );
  NANDN U24319 ( .A(n23780), .B(n23779), .Z(n23781) );
  AND U24320 ( .A(n23782), .B(n23781), .Z(n23824) );
  XNOR U24321 ( .A(n23825), .B(n23824), .Z(n23826) );
  XNOR U24322 ( .A(n23827), .B(n23826), .Z(n24076) );
  XNOR U24323 ( .A(n24077), .B(n24076), .Z(n24078) );
  XOR U24324 ( .A(n24079), .B(n24078), .Z(n23821) );
  XNOR U24325 ( .A(n23820), .B(n23821), .Z(n23814) );
  XOR U24326 ( .A(n23815), .B(n23814), .Z(n23807) );
  NANDN U24327 ( .A(n23784), .B(n23783), .Z(n23788) );
  NANDN U24328 ( .A(n23786), .B(n23785), .Z(n23787) );
  AND U24329 ( .A(n23788), .B(n23787), .Z(n23806) );
  XNOR U24330 ( .A(n23807), .B(n23806), .Z(n23808) );
  NANDN U24331 ( .A(n23790), .B(n23789), .Z(n23794) );
  NAND U24332 ( .A(n23792), .B(n23791), .Z(n23793) );
  NAND U24333 ( .A(n23794), .B(n23793), .Z(n23809) );
  XNOR U24334 ( .A(n23808), .B(n23809), .Z(n23800) );
  XNOR U24335 ( .A(n23801), .B(n23800), .Z(n23802) );
  XNOR U24336 ( .A(n23803), .B(n23802), .Z(n24088) );
  XNOR U24337 ( .A(sreg[176]), .B(n24088), .Z(n24090) );
  NANDN U24338 ( .A(sreg[175]), .B(n23795), .Z(n23799) );
  NAND U24339 ( .A(n23797), .B(n23796), .Z(n23798) );
  NAND U24340 ( .A(n23799), .B(n23798), .Z(n24089) );
  XNOR U24341 ( .A(n24090), .B(n24089), .Z(c[176]) );
  NANDN U24342 ( .A(n23801), .B(n23800), .Z(n23805) );
  NANDN U24343 ( .A(n23803), .B(n23802), .Z(n23804) );
  AND U24344 ( .A(n23805), .B(n23804), .Z(n24096) );
  NANDN U24345 ( .A(n23807), .B(n23806), .Z(n23811) );
  NANDN U24346 ( .A(n23809), .B(n23808), .Z(n23810) );
  AND U24347 ( .A(n23811), .B(n23810), .Z(n24094) );
  NANDN U24348 ( .A(n23813), .B(n23812), .Z(n23817) );
  NAND U24349 ( .A(n23815), .B(n23814), .Z(n23816) );
  AND U24350 ( .A(n23817), .B(n23816), .Z(n24377) );
  NANDN U24351 ( .A(n23819), .B(n23818), .Z(n23823) );
  NANDN U24352 ( .A(n23821), .B(n23820), .Z(n23822) );
  AND U24353 ( .A(n23823), .B(n23822), .Z(n24376) );
  NANDN U24354 ( .A(n23825), .B(n23824), .Z(n23829) );
  NANDN U24355 ( .A(n23827), .B(n23826), .Z(n23828) );
  AND U24356 ( .A(n23829), .B(n23828), .Z(n24101) );
  NANDN U24357 ( .A(n23831), .B(n23830), .Z(n23835) );
  NAND U24358 ( .A(n23833), .B(n23832), .Z(n23834) );
  AND U24359 ( .A(n23835), .B(n23834), .Z(n24131) );
  NANDN U24360 ( .A(n23837), .B(n23836), .Z(n23841) );
  NANDN U24361 ( .A(n23839), .B(n23838), .Z(n23840) );
  AND U24362 ( .A(n23841), .B(n23840), .Z(n24125) );
  NANDN U24363 ( .A(n23843), .B(n23842), .Z(n23847) );
  NANDN U24364 ( .A(n23845), .B(n23844), .Z(n23846) );
  AND U24365 ( .A(n23847), .B(n23846), .Z(n24124) );
  NANDN U24366 ( .A(n33875), .B(n23848), .Z(n23850) );
  XOR U24367 ( .A(b[25]), .B(a[89]), .Z(n24159) );
  NANDN U24368 ( .A(n33994), .B(n24159), .Z(n23849) );
  AND U24369 ( .A(n23850), .B(n23849), .Z(n24287) );
  NANDN U24370 ( .A(n32013), .B(n23851), .Z(n23853) );
  XOR U24371 ( .A(a[97]), .B(b[17]), .Z(n24162) );
  NANDN U24372 ( .A(n32292), .B(n24162), .Z(n23852) );
  AND U24373 ( .A(n23853), .B(n23852), .Z(n24286) );
  NANDN U24374 ( .A(n31536), .B(n23854), .Z(n23856) );
  XOR U24375 ( .A(a[99]), .B(b[15]), .Z(n24165) );
  NANDN U24376 ( .A(n31925), .B(n24165), .Z(n23855) );
  NAND U24377 ( .A(n23856), .B(n23855), .Z(n24285) );
  XOR U24378 ( .A(n24286), .B(n24285), .Z(n24288) );
  XOR U24379 ( .A(n24287), .B(n24288), .Z(n24352) );
  NANDN U24380 ( .A(n37526), .B(n23857), .Z(n23859) );
  XOR U24381 ( .A(b[51]), .B(a[63]), .Z(n24168) );
  NANDN U24382 ( .A(n37605), .B(n24168), .Z(n23858) );
  AND U24383 ( .A(n23859), .B(n23858), .Z(n24311) );
  NANDN U24384 ( .A(n37705), .B(n23860), .Z(n23862) );
  XOR U24385 ( .A(b[53]), .B(a[61]), .Z(n24171) );
  NANDN U24386 ( .A(n37778), .B(n24171), .Z(n23861) );
  AND U24387 ( .A(n23862), .B(n23861), .Z(n24310) );
  NANDN U24388 ( .A(n36210), .B(n23863), .Z(n23865) );
  XOR U24389 ( .A(b[39]), .B(a[75]), .Z(n24174) );
  NANDN U24390 ( .A(n36347), .B(n24174), .Z(n23864) );
  NAND U24391 ( .A(n23865), .B(n23864), .Z(n24309) );
  XOR U24392 ( .A(n24310), .B(n24309), .Z(n24312) );
  XNOR U24393 ( .A(n24311), .B(n24312), .Z(n24351) );
  XNOR U24394 ( .A(n24352), .B(n24351), .Z(n24354) );
  NANDN U24395 ( .A(n23867), .B(n23866), .Z(n23871) );
  OR U24396 ( .A(n23869), .B(n23868), .Z(n23870) );
  AND U24397 ( .A(n23871), .B(n23870), .Z(n24353) );
  XOR U24398 ( .A(n24354), .B(n24353), .Z(n24150) );
  NANDN U24399 ( .A(n23873), .B(n23872), .Z(n23877) );
  OR U24400 ( .A(n23875), .B(n23874), .Z(n23876) );
  AND U24401 ( .A(n23877), .B(n23876), .Z(n24148) );
  NANDN U24402 ( .A(n23879), .B(n23878), .Z(n23883) );
  NANDN U24403 ( .A(n23881), .B(n23880), .Z(n23882) );
  NAND U24404 ( .A(n23883), .B(n23882), .Z(n24147) );
  XNOR U24405 ( .A(n24148), .B(n24147), .Z(n24149) );
  XNOR U24406 ( .A(n24150), .B(n24149), .Z(n24123) );
  XOR U24407 ( .A(n24124), .B(n24123), .Z(n24126) );
  XOR U24408 ( .A(n24125), .B(n24126), .Z(n24130) );
  NANDN U24409 ( .A(n23885), .B(n23884), .Z(n23889) );
  NANDN U24410 ( .A(n23887), .B(n23886), .Z(n23888) );
  AND U24411 ( .A(n23889), .B(n23888), .Z(n24118) );
  NANDN U24412 ( .A(n211), .B(n23890), .Z(n23892) );
  XOR U24413 ( .A(b[47]), .B(a[67]), .Z(n24222) );
  NANDN U24414 ( .A(n37172), .B(n24222), .Z(n23891) );
  AND U24415 ( .A(n23892), .B(n23891), .Z(n24212) );
  NANDN U24416 ( .A(n210), .B(n23893), .Z(n23895) );
  XOR U24417 ( .A(a[105]), .B(b[9]), .Z(n24225) );
  NANDN U24418 ( .A(n30267), .B(n24225), .Z(n23894) );
  AND U24419 ( .A(n23895), .B(n23894), .Z(n24211) );
  NANDN U24420 ( .A(n212), .B(n23896), .Z(n23898) );
  XOR U24421 ( .A(b[49]), .B(a[65]), .Z(n24228) );
  NANDN U24422 ( .A(n37432), .B(n24228), .Z(n23897) );
  NAND U24423 ( .A(n23898), .B(n23897), .Z(n24210) );
  XOR U24424 ( .A(n24211), .B(n24210), .Z(n24213) );
  XOR U24425 ( .A(n24212), .B(n24213), .Z(n24265) );
  NANDN U24426 ( .A(n36742), .B(n23899), .Z(n23901) );
  XOR U24427 ( .A(b[43]), .B(a[71]), .Z(n24231) );
  NANDN U24428 ( .A(n36891), .B(n24231), .Z(n23900) );
  AND U24429 ( .A(n23901), .B(n23900), .Z(n24242) );
  NANDN U24430 ( .A(n36991), .B(n23902), .Z(n23904) );
  XOR U24431 ( .A(b[45]), .B(a[69]), .Z(n24234) );
  NANDN U24432 ( .A(n37083), .B(n24234), .Z(n23903) );
  AND U24433 ( .A(n23904), .B(n23903), .Z(n24241) );
  NANDN U24434 ( .A(n30482), .B(n23905), .Z(n23907) );
  XOR U24435 ( .A(a[103]), .B(b[11]), .Z(n24237) );
  NANDN U24436 ( .A(n30891), .B(n24237), .Z(n23906) );
  NAND U24437 ( .A(n23907), .B(n23906), .Z(n24240) );
  XOR U24438 ( .A(n24241), .B(n24240), .Z(n24243) );
  XNOR U24439 ( .A(n24242), .B(n24243), .Z(n24264) );
  XNOR U24440 ( .A(n24265), .B(n24264), .Z(n24266) );
  NANDN U24441 ( .A(n23909), .B(n23908), .Z(n23913) );
  OR U24442 ( .A(n23911), .B(n23910), .Z(n23912) );
  NAND U24443 ( .A(n23913), .B(n23912), .Z(n24267) );
  XNOR U24444 ( .A(n24266), .B(n24267), .Z(n24117) );
  XNOR U24445 ( .A(n24118), .B(n24117), .Z(n24119) );
  NANDN U24446 ( .A(n29499), .B(n23914), .Z(n23916) );
  XOR U24447 ( .A(a[107]), .B(b[7]), .Z(n24195) );
  NANDN U24448 ( .A(n29735), .B(n24195), .Z(n23915) );
  AND U24449 ( .A(n23916), .B(n23915), .Z(n24185) );
  NANDN U24450 ( .A(n37857), .B(n23917), .Z(n23919) );
  XOR U24451 ( .A(b[55]), .B(a[59]), .Z(n24198) );
  NANDN U24452 ( .A(n37911), .B(n24198), .Z(n23918) );
  AND U24453 ( .A(n23919), .B(n23918), .Z(n24184) );
  NANDN U24454 ( .A(n35611), .B(n23920), .Z(n23922) );
  XOR U24455 ( .A(b[35]), .B(a[79]), .Z(n24201) );
  NANDN U24456 ( .A(n35801), .B(n24201), .Z(n23921) );
  NAND U24457 ( .A(n23922), .B(n23921), .Z(n24183) );
  XOR U24458 ( .A(n24184), .B(n24183), .Z(n24186) );
  XOR U24459 ( .A(n24185), .B(n24186), .Z(n24247) );
  NANDN U24460 ( .A(n23924), .B(n23923), .Z(n23928) );
  OR U24461 ( .A(n23926), .B(n23925), .Z(n23927) );
  AND U24462 ( .A(n23928), .B(n23927), .Z(n24246) );
  XNOR U24463 ( .A(n24247), .B(n24246), .Z(n24248) );
  NANDN U24464 ( .A(n23930), .B(n23929), .Z(n23934) );
  OR U24465 ( .A(n23932), .B(n23931), .Z(n23933) );
  NAND U24466 ( .A(n23934), .B(n23933), .Z(n24249) );
  XOR U24467 ( .A(n24248), .B(n24249), .Z(n24120) );
  XNOR U24468 ( .A(n24119), .B(n24120), .Z(n24129) );
  XOR U24469 ( .A(n24130), .B(n24129), .Z(n24132) );
  XOR U24470 ( .A(n24131), .B(n24132), .Z(n24100) );
  NANDN U24471 ( .A(n23936), .B(n23935), .Z(n23940) );
  NANDN U24472 ( .A(n23938), .B(n23937), .Z(n23939) );
  AND U24473 ( .A(n23940), .B(n23939), .Z(n24113) );
  NANDN U24474 ( .A(n23942), .B(n23941), .Z(n23946) );
  NANDN U24475 ( .A(n23944), .B(n23943), .Z(n23945) );
  AND U24476 ( .A(n23946), .B(n23945), .Z(n24112) );
  NANDN U24477 ( .A(n23948), .B(n23947), .Z(n23952) );
  NAND U24478 ( .A(n23950), .B(n23949), .Z(n23951) );
  AND U24479 ( .A(n23952), .B(n23951), .Z(n24111) );
  XOR U24480 ( .A(n24112), .B(n24111), .Z(n24114) );
  XOR U24481 ( .A(n24113), .B(n24114), .Z(n24138) );
  NANDN U24482 ( .A(n23954), .B(n23953), .Z(n23958) );
  NANDN U24483 ( .A(n23956), .B(n23955), .Z(n23957) );
  AND U24484 ( .A(n23958), .B(n23957), .Z(n24360) );
  NANDN U24485 ( .A(n32996), .B(n23959), .Z(n23961) );
  XOR U24486 ( .A(a[93]), .B(b[21]), .Z(n24270) );
  NANDN U24487 ( .A(n33271), .B(n24270), .Z(n23960) );
  AND U24488 ( .A(n23961), .B(n23960), .Z(n24329) );
  NANDN U24489 ( .A(n33866), .B(n23962), .Z(n23964) );
  XOR U24490 ( .A(a[91]), .B(b[23]), .Z(n24273) );
  NANDN U24491 ( .A(n33644), .B(n24273), .Z(n23963) );
  AND U24492 ( .A(n23964), .B(n23963), .Z(n24328) );
  NANDN U24493 ( .A(n32483), .B(n23965), .Z(n23967) );
  XOR U24494 ( .A(a[95]), .B(b[19]), .Z(n24276) );
  NANDN U24495 ( .A(n32823), .B(n24276), .Z(n23966) );
  NAND U24496 ( .A(n23967), .B(n23966), .Z(n24327) );
  XOR U24497 ( .A(n24328), .B(n24327), .Z(n24330) );
  XOR U24498 ( .A(n24329), .B(n24330), .Z(n24217) );
  NANDN U24499 ( .A(n34909), .B(n23968), .Z(n23970) );
  XOR U24500 ( .A(b[31]), .B(a[83]), .Z(n24279) );
  NANDN U24501 ( .A(n35145), .B(n24279), .Z(n23969) );
  AND U24502 ( .A(n23970), .B(n23969), .Z(n24206) );
  NANDN U24503 ( .A(n38247), .B(n23971), .Z(n23973) );
  XOR U24504 ( .A(b[61]), .B(a[53]), .Z(n24282) );
  NANDN U24505 ( .A(n38248), .B(n24282), .Z(n23972) );
  AND U24506 ( .A(n23973), .B(n23972), .Z(n24205) );
  AND U24507 ( .A(b[63]), .B(a[49]), .Z(n24204) );
  XOR U24508 ( .A(n24205), .B(n24204), .Z(n24207) );
  XNOR U24509 ( .A(n24206), .B(n24207), .Z(n24216) );
  XNOR U24510 ( .A(n24217), .B(n24216), .Z(n24218) );
  NANDN U24511 ( .A(n23975), .B(n23974), .Z(n23979) );
  OR U24512 ( .A(n23977), .B(n23976), .Z(n23978) );
  NAND U24513 ( .A(n23979), .B(n23978), .Z(n24219) );
  XNOR U24514 ( .A(n24218), .B(n24219), .Z(n24357) );
  NANDN U24515 ( .A(n34223), .B(n23980), .Z(n23982) );
  XOR U24516 ( .A(b[27]), .B(a[87]), .Z(n24291) );
  NANDN U24517 ( .A(n34458), .B(n24291), .Z(n23981) );
  AND U24518 ( .A(n23982), .B(n23981), .Z(n24179) );
  NANDN U24519 ( .A(n34634), .B(n23983), .Z(n23985) );
  XOR U24520 ( .A(b[29]), .B(a[85]), .Z(n24294) );
  NANDN U24521 ( .A(n34722), .B(n24294), .Z(n23984) );
  AND U24522 ( .A(n23985), .B(n23984), .Z(n24178) );
  NANDN U24523 ( .A(n31055), .B(n23986), .Z(n23988) );
  XOR U24524 ( .A(a[101]), .B(b[13]), .Z(n24297) );
  NANDN U24525 ( .A(n31293), .B(n24297), .Z(n23987) );
  NAND U24526 ( .A(n23988), .B(n23987), .Z(n24177) );
  XOR U24527 ( .A(n24178), .B(n24177), .Z(n24180) );
  XOR U24528 ( .A(n24179), .B(n24180), .Z(n24253) );
  NANDN U24529 ( .A(n28889), .B(n23989), .Z(n23991) );
  XOR U24530 ( .A(a[109]), .B(b[5]), .Z(n24300) );
  NANDN U24531 ( .A(n29138), .B(n24300), .Z(n23990) );
  AND U24532 ( .A(n23991), .B(n23990), .Z(n24323) );
  NANDN U24533 ( .A(n209), .B(n23992), .Z(n23994) );
  XOR U24534 ( .A(a[111]), .B(b[3]), .Z(n24303) );
  NANDN U24535 ( .A(n28941), .B(n24303), .Z(n23993) );
  AND U24536 ( .A(n23994), .B(n23993), .Z(n24322) );
  NANDN U24537 ( .A(n35936), .B(n23995), .Z(n23997) );
  XOR U24538 ( .A(b[37]), .B(a[77]), .Z(n24306) );
  NANDN U24539 ( .A(n36047), .B(n24306), .Z(n23996) );
  NAND U24540 ( .A(n23997), .B(n23996), .Z(n24321) );
  XOR U24541 ( .A(n24322), .B(n24321), .Z(n24324) );
  XNOR U24542 ( .A(n24323), .B(n24324), .Z(n24252) );
  XNOR U24543 ( .A(n24253), .B(n24252), .Z(n24254) );
  NANDN U24544 ( .A(n23999), .B(n23998), .Z(n24003) );
  OR U24545 ( .A(n24001), .B(n24000), .Z(n24002) );
  NAND U24546 ( .A(n24003), .B(n24002), .Z(n24255) );
  XOR U24547 ( .A(n24254), .B(n24255), .Z(n24358) );
  XNOR U24548 ( .A(n24357), .B(n24358), .Z(n24359) );
  XNOR U24549 ( .A(n24360), .B(n24359), .Z(n24144) );
  NANDN U24550 ( .A(n24005), .B(n24004), .Z(n24009) );
  NANDN U24551 ( .A(n24007), .B(n24006), .Z(n24008) );
  AND U24552 ( .A(n24009), .B(n24008), .Z(n24259) );
  NANDN U24553 ( .A(n24011), .B(n24010), .Z(n24015) );
  OR U24554 ( .A(n24013), .B(n24012), .Z(n24014) );
  NAND U24555 ( .A(n24015), .B(n24014), .Z(n24258) );
  XNOR U24556 ( .A(n24259), .B(n24258), .Z(n24261) );
  NANDN U24557 ( .A(n24017), .B(n24016), .Z(n24021) );
  OR U24558 ( .A(n24019), .B(n24018), .Z(n24020) );
  AND U24559 ( .A(n24021), .B(n24020), .Z(n24156) );
  NAND U24560 ( .A(b[0]), .B(a[113]), .Z(n24022) );
  XNOR U24561 ( .A(b[1]), .B(n24022), .Z(n24024) );
  NANDN U24562 ( .A(b[0]), .B(a[112]), .Z(n24023) );
  NAND U24563 ( .A(n24024), .B(n24023), .Z(n24192) );
  NANDN U24564 ( .A(n38278), .B(n24025), .Z(n24027) );
  XOR U24565 ( .A(b[63]), .B(a[51]), .Z(n24336) );
  NANDN U24566 ( .A(n38279), .B(n24336), .Z(n24026) );
  AND U24567 ( .A(n24027), .B(n24026), .Z(n24190) );
  NANDN U24568 ( .A(n35260), .B(n24028), .Z(n24030) );
  XOR U24569 ( .A(b[33]), .B(a[81]), .Z(n24339) );
  NANDN U24570 ( .A(n35456), .B(n24339), .Z(n24029) );
  NAND U24571 ( .A(n24030), .B(n24029), .Z(n24189) );
  XNOR U24572 ( .A(n24190), .B(n24189), .Z(n24191) );
  XNOR U24573 ( .A(n24192), .B(n24191), .Z(n24153) );
  NANDN U24574 ( .A(n37974), .B(n24031), .Z(n24033) );
  XOR U24575 ( .A(b[57]), .B(a[57]), .Z(n24342) );
  NANDN U24576 ( .A(n38031), .B(n24342), .Z(n24032) );
  AND U24577 ( .A(n24033), .B(n24032), .Z(n24318) );
  NANDN U24578 ( .A(n38090), .B(n24034), .Z(n24036) );
  XOR U24579 ( .A(b[59]), .B(a[55]), .Z(n24345) );
  NANDN U24580 ( .A(n38130), .B(n24345), .Z(n24035) );
  AND U24581 ( .A(n24036), .B(n24035), .Z(n24316) );
  NANDN U24582 ( .A(n36480), .B(n24037), .Z(n24039) );
  XOR U24583 ( .A(b[41]), .B(a[73]), .Z(n24348) );
  NANDN U24584 ( .A(n36594), .B(n24348), .Z(n24038) );
  NAND U24585 ( .A(n24039), .B(n24038), .Z(n24315) );
  XNOR U24586 ( .A(n24316), .B(n24315), .Z(n24317) );
  XOR U24587 ( .A(n24318), .B(n24317), .Z(n24154) );
  XNOR U24588 ( .A(n24153), .B(n24154), .Z(n24155) );
  XNOR U24589 ( .A(n24156), .B(n24155), .Z(n24260) );
  XOR U24590 ( .A(n24261), .B(n24260), .Z(n24142) );
  NANDN U24591 ( .A(n24041), .B(n24040), .Z(n24045) );
  NAND U24592 ( .A(n24043), .B(n24042), .Z(n24044) );
  NAND U24593 ( .A(n24045), .B(n24044), .Z(n24141) );
  XNOR U24594 ( .A(n24142), .B(n24141), .Z(n24143) );
  XOR U24595 ( .A(n24144), .B(n24143), .Z(n24136) );
  NANDN U24596 ( .A(n24047), .B(n24046), .Z(n24051) );
  NANDN U24597 ( .A(n24049), .B(n24048), .Z(n24050) );
  AND U24598 ( .A(n24051), .B(n24050), .Z(n24135) );
  XNOR U24599 ( .A(n24136), .B(n24135), .Z(n24137) );
  XNOR U24600 ( .A(n24138), .B(n24137), .Z(n24099) );
  XOR U24601 ( .A(n24100), .B(n24099), .Z(n24102) );
  XOR U24602 ( .A(n24101), .B(n24102), .Z(n24365) );
  NANDN U24603 ( .A(n24053), .B(n24052), .Z(n24057) );
  OR U24604 ( .A(n24055), .B(n24054), .Z(n24056) );
  AND U24605 ( .A(n24057), .B(n24056), .Z(n24364) );
  NANDN U24606 ( .A(n24059), .B(n24058), .Z(n24063) );
  OR U24607 ( .A(n24061), .B(n24060), .Z(n24062) );
  AND U24608 ( .A(n24063), .B(n24062), .Z(n24108) );
  NANDN U24609 ( .A(n24065), .B(n24064), .Z(n24069) );
  NANDN U24610 ( .A(n24067), .B(n24066), .Z(n24068) );
  AND U24611 ( .A(n24069), .B(n24068), .Z(n24106) );
  NANDN U24612 ( .A(n24071), .B(n24070), .Z(n24075) );
  OR U24613 ( .A(n24073), .B(n24072), .Z(n24074) );
  AND U24614 ( .A(n24075), .B(n24074), .Z(n24105) );
  XNOR U24615 ( .A(n24106), .B(n24105), .Z(n24107) );
  XNOR U24616 ( .A(n24108), .B(n24107), .Z(n24363) );
  XOR U24617 ( .A(n24364), .B(n24363), .Z(n24366) );
  XOR U24618 ( .A(n24365), .B(n24366), .Z(n24372) );
  NANDN U24619 ( .A(n24077), .B(n24076), .Z(n24081) );
  NANDN U24620 ( .A(n24079), .B(n24078), .Z(n24080) );
  AND U24621 ( .A(n24081), .B(n24080), .Z(n24370) );
  NANDN U24622 ( .A(n24083), .B(n24082), .Z(n24087) );
  OR U24623 ( .A(n24085), .B(n24084), .Z(n24086) );
  AND U24624 ( .A(n24087), .B(n24086), .Z(n24369) );
  XNOR U24625 ( .A(n24370), .B(n24369), .Z(n24371) );
  XNOR U24626 ( .A(n24372), .B(n24371), .Z(n24375) );
  XOR U24627 ( .A(n24376), .B(n24375), .Z(n24378) );
  XNOR U24628 ( .A(n24377), .B(n24378), .Z(n24093) );
  XNOR U24629 ( .A(n24094), .B(n24093), .Z(n24095) );
  XNOR U24630 ( .A(n24096), .B(n24095), .Z(n24381) );
  XNOR U24631 ( .A(sreg[177]), .B(n24381), .Z(n24383) );
  NANDN U24632 ( .A(sreg[176]), .B(n24088), .Z(n24092) );
  NAND U24633 ( .A(n24090), .B(n24089), .Z(n24091) );
  NAND U24634 ( .A(n24092), .B(n24091), .Z(n24382) );
  XNOR U24635 ( .A(n24383), .B(n24382), .Z(c[177]) );
  NANDN U24636 ( .A(n24094), .B(n24093), .Z(n24098) );
  NANDN U24637 ( .A(n24096), .B(n24095), .Z(n24097) );
  AND U24638 ( .A(n24098), .B(n24097), .Z(n24389) );
  NANDN U24639 ( .A(n24100), .B(n24099), .Z(n24104) );
  OR U24640 ( .A(n24102), .B(n24101), .Z(n24103) );
  AND U24641 ( .A(n24104), .B(n24103), .Z(n24393) );
  NANDN U24642 ( .A(n24106), .B(n24105), .Z(n24110) );
  NANDN U24643 ( .A(n24108), .B(n24107), .Z(n24109) );
  AND U24644 ( .A(n24110), .B(n24109), .Z(n24392) );
  XNOR U24645 ( .A(n24393), .B(n24392), .Z(n24395) );
  NANDN U24646 ( .A(n24112), .B(n24111), .Z(n24116) );
  OR U24647 ( .A(n24114), .B(n24113), .Z(n24115) );
  AND U24648 ( .A(n24116), .B(n24115), .Z(n24664) );
  NANDN U24649 ( .A(n24118), .B(n24117), .Z(n24122) );
  NANDN U24650 ( .A(n24120), .B(n24119), .Z(n24121) );
  AND U24651 ( .A(n24122), .B(n24121), .Z(n24663) );
  NANDN U24652 ( .A(n24124), .B(n24123), .Z(n24128) );
  OR U24653 ( .A(n24126), .B(n24125), .Z(n24127) );
  AND U24654 ( .A(n24128), .B(n24127), .Z(n24662) );
  XOR U24655 ( .A(n24663), .B(n24662), .Z(n24665) );
  XOR U24656 ( .A(n24664), .B(n24665), .Z(n24399) );
  NANDN U24657 ( .A(n24130), .B(n24129), .Z(n24134) );
  OR U24658 ( .A(n24132), .B(n24131), .Z(n24133) );
  AND U24659 ( .A(n24134), .B(n24133), .Z(n24398) );
  XNOR U24660 ( .A(n24399), .B(n24398), .Z(n24400) );
  NANDN U24661 ( .A(n24136), .B(n24135), .Z(n24140) );
  NANDN U24662 ( .A(n24138), .B(n24137), .Z(n24139) );
  AND U24663 ( .A(n24140), .B(n24139), .Z(n24659) );
  NANDN U24664 ( .A(n24142), .B(n24141), .Z(n24146) );
  NAND U24665 ( .A(n24144), .B(n24143), .Z(n24145) );
  AND U24666 ( .A(n24146), .B(n24145), .Z(n24634) );
  NANDN U24667 ( .A(n24148), .B(n24147), .Z(n24152) );
  NANDN U24668 ( .A(n24150), .B(n24149), .Z(n24151) );
  AND U24669 ( .A(n24152), .B(n24151), .Z(n24652) );
  NANDN U24670 ( .A(n24154), .B(n24153), .Z(n24158) );
  NANDN U24671 ( .A(n24156), .B(n24155), .Z(n24157) );
  AND U24672 ( .A(n24158), .B(n24157), .Z(n24651) );
  NANDN U24673 ( .A(n33875), .B(n24159), .Z(n24161) );
  XOR U24674 ( .A(a[90]), .B(b[25]), .Z(n24428) );
  NANDN U24675 ( .A(n33994), .B(n24428), .Z(n24160) );
  AND U24676 ( .A(n24161), .B(n24160), .Z(n24556) );
  NANDN U24677 ( .A(n32013), .B(n24162), .Z(n24164) );
  XOR U24678 ( .A(a[98]), .B(b[17]), .Z(n24431) );
  NANDN U24679 ( .A(n32292), .B(n24431), .Z(n24163) );
  AND U24680 ( .A(n24164), .B(n24163), .Z(n24555) );
  NANDN U24681 ( .A(n31536), .B(n24165), .Z(n24167) );
  XOR U24682 ( .A(a[100]), .B(b[15]), .Z(n24434) );
  NANDN U24683 ( .A(n31925), .B(n24434), .Z(n24166) );
  NAND U24684 ( .A(n24167), .B(n24166), .Z(n24554) );
  XOR U24685 ( .A(n24555), .B(n24554), .Z(n24557) );
  XOR U24686 ( .A(n24556), .B(n24557), .Z(n24621) );
  NANDN U24687 ( .A(n37526), .B(n24168), .Z(n24170) );
  XOR U24688 ( .A(b[51]), .B(a[64]), .Z(n24437) );
  NANDN U24689 ( .A(n37605), .B(n24437), .Z(n24169) );
  AND U24690 ( .A(n24170), .B(n24169), .Z(n24580) );
  NANDN U24691 ( .A(n37705), .B(n24171), .Z(n24173) );
  XOR U24692 ( .A(b[53]), .B(a[62]), .Z(n24440) );
  NANDN U24693 ( .A(n37778), .B(n24440), .Z(n24172) );
  AND U24694 ( .A(n24173), .B(n24172), .Z(n24579) );
  NANDN U24695 ( .A(n36210), .B(n24174), .Z(n24176) );
  XOR U24696 ( .A(b[39]), .B(a[76]), .Z(n24443) );
  NANDN U24697 ( .A(n36347), .B(n24443), .Z(n24175) );
  NAND U24698 ( .A(n24176), .B(n24175), .Z(n24578) );
  XOR U24699 ( .A(n24579), .B(n24578), .Z(n24581) );
  XNOR U24700 ( .A(n24580), .B(n24581), .Z(n24620) );
  XNOR U24701 ( .A(n24621), .B(n24620), .Z(n24623) );
  NANDN U24702 ( .A(n24178), .B(n24177), .Z(n24182) );
  OR U24703 ( .A(n24180), .B(n24179), .Z(n24181) );
  AND U24704 ( .A(n24182), .B(n24181), .Z(n24622) );
  XOR U24705 ( .A(n24623), .B(n24622), .Z(n24419) );
  NANDN U24706 ( .A(n24184), .B(n24183), .Z(n24188) );
  OR U24707 ( .A(n24186), .B(n24185), .Z(n24187) );
  AND U24708 ( .A(n24188), .B(n24187), .Z(n24417) );
  NANDN U24709 ( .A(n24190), .B(n24189), .Z(n24194) );
  NANDN U24710 ( .A(n24192), .B(n24191), .Z(n24193) );
  NAND U24711 ( .A(n24194), .B(n24193), .Z(n24416) );
  XNOR U24712 ( .A(n24417), .B(n24416), .Z(n24418) );
  XNOR U24713 ( .A(n24419), .B(n24418), .Z(n24650) );
  XOR U24714 ( .A(n24651), .B(n24650), .Z(n24653) );
  XOR U24715 ( .A(n24652), .B(n24653), .Z(n24633) );
  NANDN U24716 ( .A(n29499), .B(n24195), .Z(n24197) );
  XOR U24717 ( .A(a[108]), .B(b[7]), .Z(n24494) );
  NANDN U24718 ( .A(n29735), .B(n24494), .Z(n24196) );
  AND U24719 ( .A(n24197), .B(n24196), .Z(n24454) );
  NANDN U24720 ( .A(n37857), .B(n24198), .Z(n24200) );
  XOR U24721 ( .A(b[55]), .B(a[60]), .Z(n24497) );
  NANDN U24722 ( .A(n37911), .B(n24497), .Z(n24199) );
  AND U24723 ( .A(n24200), .B(n24199), .Z(n24453) );
  NANDN U24724 ( .A(n35611), .B(n24201), .Z(n24203) );
  XOR U24725 ( .A(b[35]), .B(a[80]), .Z(n24500) );
  NANDN U24726 ( .A(n35801), .B(n24500), .Z(n24202) );
  NAND U24727 ( .A(n24203), .B(n24202), .Z(n24452) );
  XOR U24728 ( .A(n24453), .B(n24452), .Z(n24455) );
  XOR U24729 ( .A(n24454), .B(n24455), .Z(n24516) );
  NANDN U24730 ( .A(n24205), .B(n24204), .Z(n24209) );
  OR U24731 ( .A(n24207), .B(n24206), .Z(n24208) );
  AND U24732 ( .A(n24209), .B(n24208), .Z(n24515) );
  XNOR U24733 ( .A(n24516), .B(n24515), .Z(n24517) );
  NANDN U24734 ( .A(n24211), .B(n24210), .Z(n24215) );
  OR U24735 ( .A(n24213), .B(n24212), .Z(n24214) );
  NAND U24736 ( .A(n24215), .B(n24214), .Z(n24518) );
  XNOR U24737 ( .A(n24517), .B(n24518), .Z(n24646) );
  NANDN U24738 ( .A(n24217), .B(n24216), .Z(n24221) );
  NANDN U24739 ( .A(n24219), .B(n24218), .Z(n24220) );
  AND U24740 ( .A(n24221), .B(n24220), .Z(n24645) );
  NANDN U24741 ( .A(n211), .B(n24222), .Z(n24224) );
  XOR U24742 ( .A(b[47]), .B(a[68]), .Z(n24470) );
  NANDN U24743 ( .A(n37172), .B(n24470), .Z(n24223) );
  AND U24744 ( .A(n24224), .B(n24223), .Z(n24511) );
  NANDN U24745 ( .A(n210), .B(n24225), .Z(n24227) );
  XOR U24746 ( .A(a[106]), .B(b[9]), .Z(n24473) );
  NANDN U24747 ( .A(n30267), .B(n24473), .Z(n24226) );
  AND U24748 ( .A(n24227), .B(n24226), .Z(n24510) );
  NANDN U24749 ( .A(n212), .B(n24228), .Z(n24230) );
  XOR U24750 ( .A(b[49]), .B(a[66]), .Z(n24476) );
  NANDN U24751 ( .A(n37432), .B(n24476), .Z(n24229) );
  NAND U24752 ( .A(n24230), .B(n24229), .Z(n24509) );
  XOR U24753 ( .A(n24510), .B(n24509), .Z(n24512) );
  XOR U24754 ( .A(n24511), .B(n24512), .Z(n24534) );
  NANDN U24755 ( .A(n36742), .B(n24231), .Z(n24233) );
  XOR U24756 ( .A(b[43]), .B(a[72]), .Z(n24479) );
  NANDN U24757 ( .A(n36891), .B(n24479), .Z(n24232) );
  AND U24758 ( .A(n24233), .B(n24232), .Z(n24490) );
  NANDN U24759 ( .A(n36991), .B(n24234), .Z(n24236) );
  XOR U24760 ( .A(b[45]), .B(a[70]), .Z(n24482) );
  NANDN U24761 ( .A(n37083), .B(n24482), .Z(n24235) );
  AND U24762 ( .A(n24236), .B(n24235), .Z(n24489) );
  NANDN U24763 ( .A(n30482), .B(n24237), .Z(n24239) );
  XOR U24764 ( .A(a[104]), .B(b[11]), .Z(n24485) );
  NANDN U24765 ( .A(n30891), .B(n24485), .Z(n24238) );
  NAND U24766 ( .A(n24239), .B(n24238), .Z(n24488) );
  XOR U24767 ( .A(n24489), .B(n24488), .Z(n24491) );
  XNOR U24768 ( .A(n24490), .B(n24491), .Z(n24533) );
  XNOR U24769 ( .A(n24534), .B(n24533), .Z(n24535) );
  NANDN U24770 ( .A(n24241), .B(n24240), .Z(n24245) );
  OR U24771 ( .A(n24243), .B(n24242), .Z(n24244) );
  NAND U24772 ( .A(n24245), .B(n24244), .Z(n24536) );
  XNOR U24773 ( .A(n24535), .B(n24536), .Z(n24644) );
  XOR U24774 ( .A(n24645), .B(n24644), .Z(n24647) );
  XNOR U24775 ( .A(n24646), .B(n24647), .Z(n24632) );
  XOR U24776 ( .A(n24633), .B(n24632), .Z(n24635) );
  XOR U24777 ( .A(n24634), .B(n24635), .Z(n24657) );
  NANDN U24778 ( .A(n24247), .B(n24246), .Z(n24251) );
  NANDN U24779 ( .A(n24249), .B(n24248), .Z(n24250) );
  AND U24780 ( .A(n24251), .B(n24250), .Z(n24640) );
  NANDN U24781 ( .A(n24253), .B(n24252), .Z(n24257) );
  NANDN U24782 ( .A(n24255), .B(n24254), .Z(n24256) );
  AND U24783 ( .A(n24257), .B(n24256), .Z(n24639) );
  NANDN U24784 ( .A(n24259), .B(n24258), .Z(n24263) );
  NAND U24785 ( .A(n24261), .B(n24260), .Z(n24262) );
  AND U24786 ( .A(n24263), .B(n24262), .Z(n24638) );
  XOR U24787 ( .A(n24639), .B(n24638), .Z(n24641) );
  XOR U24788 ( .A(n24640), .B(n24641), .Z(n24407) );
  NANDN U24789 ( .A(n24265), .B(n24264), .Z(n24269) );
  NANDN U24790 ( .A(n24267), .B(n24266), .Z(n24268) );
  AND U24791 ( .A(n24269), .B(n24268), .Z(n24629) );
  NANDN U24792 ( .A(n32996), .B(n24270), .Z(n24272) );
  XOR U24793 ( .A(a[94]), .B(b[21]), .Z(n24539) );
  NANDN U24794 ( .A(n33271), .B(n24539), .Z(n24271) );
  AND U24795 ( .A(n24272), .B(n24271), .Z(n24598) );
  NANDN U24796 ( .A(n33866), .B(n24273), .Z(n24275) );
  XOR U24797 ( .A(a[92]), .B(b[23]), .Z(n24542) );
  NANDN U24798 ( .A(n33644), .B(n24542), .Z(n24274) );
  AND U24799 ( .A(n24275), .B(n24274), .Z(n24597) );
  NANDN U24800 ( .A(n32483), .B(n24276), .Z(n24278) );
  XOR U24801 ( .A(a[96]), .B(b[19]), .Z(n24545) );
  NANDN U24802 ( .A(n32823), .B(n24545), .Z(n24277) );
  NAND U24803 ( .A(n24278), .B(n24277), .Z(n24596) );
  XOR U24804 ( .A(n24597), .B(n24596), .Z(n24599) );
  XOR U24805 ( .A(n24598), .B(n24599), .Z(n24465) );
  NANDN U24806 ( .A(n34909), .B(n24279), .Z(n24281) );
  XOR U24807 ( .A(b[31]), .B(a[84]), .Z(n24548) );
  NANDN U24808 ( .A(n35145), .B(n24548), .Z(n24280) );
  AND U24809 ( .A(n24281), .B(n24280), .Z(n24505) );
  NANDN U24810 ( .A(n38247), .B(n24282), .Z(n24284) );
  XOR U24811 ( .A(b[61]), .B(a[54]), .Z(n24551) );
  NANDN U24812 ( .A(n38248), .B(n24551), .Z(n24283) );
  AND U24813 ( .A(n24284), .B(n24283), .Z(n24504) );
  AND U24814 ( .A(b[63]), .B(a[50]), .Z(n24503) );
  XOR U24815 ( .A(n24504), .B(n24503), .Z(n24506) );
  XNOR U24816 ( .A(n24505), .B(n24506), .Z(n24464) );
  XNOR U24817 ( .A(n24465), .B(n24464), .Z(n24466) );
  NANDN U24818 ( .A(n24286), .B(n24285), .Z(n24290) );
  OR U24819 ( .A(n24288), .B(n24287), .Z(n24289) );
  NAND U24820 ( .A(n24290), .B(n24289), .Z(n24467) );
  XNOR U24821 ( .A(n24466), .B(n24467), .Z(n24626) );
  NANDN U24822 ( .A(n34223), .B(n24291), .Z(n24293) );
  XOR U24823 ( .A(b[27]), .B(a[88]), .Z(n24560) );
  NANDN U24824 ( .A(n34458), .B(n24560), .Z(n24292) );
  AND U24825 ( .A(n24293), .B(n24292), .Z(n24448) );
  NANDN U24826 ( .A(n34634), .B(n24294), .Z(n24296) );
  XOR U24827 ( .A(b[29]), .B(a[86]), .Z(n24563) );
  NANDN U24828 ( .A(n34722), .B(n24563), .Z(n24295) );
  AND U24829 ( .A(n24296), .B(n24295), .Z(n24447) );
  NANDN U24830 ( .A(n31055), .B(n24297), .Z(n24299) );
  XOR U24831 ( .A(a[102]), .B(b[13]), .Z(n24566) );
  NANDN U24832 ( .A(n31293), .B(n24566), .Z(n24298) );
  NAND U24833 ( .A(n24299), .B(n24298), .Z(n24446) );
  XOR U24834 ( .A(n24447), .B(n24446), .Z(n24449) );
  XOR U24835 ( .A(n24448), .B(n24449), .Z(n24522) );
  NANDN U24836 ( .A(n28889), .B(n24300), .Z(n24302) );
  XOR U24837 ( .A(a[110]), .B(b[5]), .Z(n24569) );
  NANDN U24838 ( .A(n29138), .B(n24569), .Z(n24301) );
  AND U24839 ( .A(n24302), .B(n24301), .Z(n24592) );
  NANDN U24840 ( .A(n209), .B(n24303), .Z(n24305) );
  XOR U24841 ( .A(a[112]), .B(b[3]), .Z(n24572) );
  NANDN U24842 ( .A(n28941), .B(n24572), .Z(n24304) );
  AND U24843 ( .A(n24305), .B(n24304), .Z(n24591) );
  NANDN U24844 ( .A(n35936), .B(n24306), .Z(n24308) );
  XOR U24845 ( .A(b[37]), .B(a[78]), .Z(n24575) );
  NANDN U24846 ( .A(n36047), .B(n24575), .Z(n24307) );
  NAND U24847 ( .A(n24308), .B(n24307), .Z(n24590) );
  XOR U24848 ( .A(n24591), .B(n24590), .Z(n24593) );
  XNOR U24849 ( .A(n24592), .B(n24593), .Z(n24521) );
  XNOR U24850 ( .A(n24522), .B(n24521), .Z(n24523) );
  NANDN U24851 ( .A(n24310), .B(n24309), .Z(n24314) );
  OR U24852 ( .A(n24312), .B(n24311), .Z(n24313) );
  NAND U24853 ( .A(n24314), .B(n24313), .Z(n24524) );
  XOR U24854 ( .A(n24523), .B(n24524), .Z(n24627) );
  XNOR U24855 ( .A(n24626), .B(n24627), .Z(n24628) );
  XNOR U24856 ( .A(n24629), .B(n24628), .Z(n24413) );
  NANDN U24857 ( .A(n24316), .B(n24315), .Z(n24320) );
  NANDN U24858 ( .A(n24318), .B(n24317), .Z(n24319) );
  AND U24859 ( .A(n24320), .B(n24319), .Z(n24528) );
  NANDN U24860 ( .A(n24322), .B(n24321), .Z(n24326) );
  OR U24861 ( .A(n24324), .B(n24323), .Z(n24325) );
  NAND U24862 ( .A(n24326), .B(n24325), .Z(n24527) );
  XNOR U24863 ( .A(n24528), .B(n24527), .Z(n24530) );
  NANDN U24864 ( .A(n24328), .B(n24327), .Z(n24332) );
  OR U24865 ( .A(n24330), .B(n24329), .Z(n24331) );
  AND U24866 ( .A(n24332), .B(n24331), .Z(n24425) );
  NAND U24867 ( .A(b[0]), .B(a[114]), .Z(n24333) );
  XNOR U24868 ( .A(b[1]), .B(n24333), .Z(n24335) );
  NANDN U24869 ( .A(b[0]), .B(a[113]), .Z(n24334) );
  NAND U24870 ( .A(n24335), .B(n24334), .Z(n24461) );
  NANDN U24871 ( .A(n38278), .B(n24336), .Z(n24338) );
  XOR U24872 ( .A(b[63]), .B(a[52]), .Z(n24605) );
  NANDN U24873 ( .A(n38279), .B(n24605), .Z(n24337) );
  AND U24874 ( .A(n24338), .B(n24337), .Z(n24459) );
  NANDN U24875 ( .A(n35260), .B(n24339), .Z(n24341) );
  XOR U24876 ( .A(b[33]), .B(a[82]), .Z(n24608) );
  NANDN U24877 ( .A(n35456), .B(n24608), .Z(n24340) );
  NAND U24878 ( .A(n24341), .B(n24340), .Z(n24458) );
  XNOR U24879 ( .A(n24459), .B(n24458), .Z(n24460) );
  XNOR U24880 ( .A(n24461), .B(n24460), .Z(n24422) );
  NANDN U24881 ( .A(n37974), .B(n24342), .Z(n24344) );
  XOR U24882 ( .A(b[57]), .B(a[58]), .Z(n24611) );
  NANDN U24883 ( .A(n38031), .B(n24611), .Z(n24343) );
  AND U24884 ( .A(n24344), .B(n24343), .Z(n24587) );
  NANDN U24885 ( .A(n38090), .B(n24345), .Z(n24347) );
  XOR U24886 ( .A(b[59]), .B(a[56]), .Z(n24614) );
  NANDN U24887 ( .A(n38130), .B(n24614), .Z(n24346) );
  AND U24888 ( .A(n24347), .B(n24346), .Z(n24585) );
  NANDN U24889 ( .A(n36480), .B(n24348), .Z(n24350) );
  XOR U24890 ( .A(b[41]), .B(a[74]), .Z(n24617) );
  NANDN U24891 ( .A(n36594), .B(n24617), .Z(n24349) );
  NAND U24892 ( .A(n24350), .B(n24349), .Z(n24584) );
  XNOR U24893 ( .A(n24585), .B(n24584), .Z(n24586) );
  XOR U24894 ( .A(n24587), .B(n24586), .Z(n24423) );
  XNOR U24895 ( .A(n24422), .B(n24423), .Z(n24424) );
  XNOR U24896 ( .A(n24425), .B(n24424), .Z(n24529) );
  XOR U24897 ( .A(n24530), .B(n24529), .Z(n24411) );
  NANDN U24898 ( .A(n24352), .B(n24351), .Z(n24356) );
  NAND U24899 ( .A(n24354), .B(n24353), .Z(n24355) );
  NAND U24900 ( .A(n24356), .B(n24355), .Z(n24410) );
  XNOR U24901 ( .A(n24411), .B(n24410), .Z(n24412) );
  XOR U24902 ( .A(n24413), .B(n24412), .Z(n24405) );
  NANDN U24903 ( .A(n24358), .B(n24357), .Z(n24362) );
  NANDN U24904 ( .A(n24360), .B(n24359), .Z(n24361) );
  AND U24905 ( .A(n24362), .B(n24361), .Z(n24404) );
  XNOR U24906 ( .A(n24405), .B(n24404), .Z(n24406) );
  XNOR U24907 ( .A(n24407), .B(n24406), .Z(n24656) );
  XNOR U24908 ( .A(n24657), .B(n24656), .Z(n24658) );
  XOR U24909 ( .A(n24659), .B(n24658), .Z(n24401) );
  XNOR U24910 ( .A(n24400), .B(n24401), .Z(n24394) );
  XOR U24911 ( .A(n24395), .B(n24394), .Z(n24669) );
  NANDN U24912 ( .A(n24364), .B(n24363), .Z(n24368) );
  OR U24913 ( .A(n24366), .B(n24365), .Z(n24367) );
  NAND U24914 ( .A(n24368), .B(n24367), .Z(n24668) );
  XNOR U24915 ( .A(n24669), .B(n24668), .Z(n24670) );
  NANDN U24916 ( .A(n24370), .B(n24369), .Z(n24374) );
  NANDN U24917 ( .A(n24372), .B(n24371), .Z(n24373) );
  NAND U24918 ( .A(n24374), .B(n24373), .Z(n24671) );
  XNOR U24919 ( .A(n24670), .B(n24671), .Z(n24386) );
  NANDN U24920 ( .A(n24376), .B(n24375), .Z(n24380) );
  OR U24921 ( .A(n24378), .B(n24377), .Z(n24379) );
  NAND U24922 ( .A(n24380), .B(n24379), .Z(n24387) );
  XNOR U24923 ( .A(n24386), .B(n24387), .Z(n24388) );
  XNOR U24924 ( .A(n24389), .B(n24388), .Z(n24674) );
  XNOR U24925 ( .A(sreg[178]), .B(n24674), .Z(n24676) );
  NANDN U24926 ( .A(sreg[177]), .B(n24381), .Z(n24385) );
  NAND U24927 ( .A(n24383), .B(n24382), .Z(n24384) );
  NAND U24928 ( .A(n24385), .B(n24384), .Z(n24675) );
  XNOR U24929 ( .A(n24676), .B(n24675), .Z(c[178]) );
  NANDN U24930 ( .A(n24387), .B(n24386), .Z(n24391) );
  NANDN U24931 ( .A(n24389), .B(n24388), .Z(n24390) );
  AND U24932 ( .A(n24391), .B(n24390), .Z(n24682) );
  NANDN U24933 ( .A(n24393), .B(n24392), .Z(n24397) );
  NAND U24934 ( .A(n24395), .B(n24394), .Z(n24396) );
  AND U24935 ( .A(n24397), .B(n24396), .Z(n24963) );
  NANDN U24936 ( .A(n24399), .B(n24398), .Z(n24403) );
  NANDN U24937 ( .A(n24401), .B(n24400), .Z(n24402) );
  AND U24938 ( .A(n24403), .B(n24402), .Z(n24962) );
  NANDN U24939 ( .A(n24405), .B(n24404), .Z(n24409) );
  NANDN U24940 ( .A(n24407), .B(n24406), .Z(n24408) );
  AND U24941 ( .A(n24409), .B(n24408), .Z(n24939) );
  NANDN U24942 ( .A(n24411), .B(n24410), .Z(n24415) );
  NAND U24943 ( .A(n24413), .B(n24412), .Z(n24414) );
  AND U24944 ( .A(n24415), .B(n24414), .Z(n24705) );
  NANDN U24945 ( .A(n24417), .B(n24416), .Z(n24421) );
  NANDN U24946 ( .A(n24419), .B(n24418), .Z(n24420) );
  AND U24947 ( .A(n24421), .B(n24420), .Z(n24699) );
  NANDN U24948 ( .A(n24423), .B(n24422), .Z(n24427) );
  NANDN U24949 ( .A(n24425), .B(n24424), .Z(n24426) );
  AND U24950 ( .A(n24427), .B(n24426), .Z(n24698) );
  NANDN U24951 ( .A(n33875), .B(n24428), .Z(n24430) );
  XOR U24952 ( .A(a[91]), .B(b[25]), .Z(n24778) );
  NANDN U24953 ( .A(n33994), .B(n24778), .Z(n24429) );
  AND U24954 ( .A(n24430), .B(n24429), .Z(n24861) );
  NANDN U24955 ( .A(n32013), .B(n24431), .Z(n24433) );
  XOR U24956 ( .A(a[99]), .B(b[17]), .Z(n24781) );
  NANDN U24957 ( .A(n32292), .B(n24781), .Z(n24432) );
  AND U24958 ( .A(n24433), .B(n24432), .Z(n24860) );
  NANDN U24959 ( .A(n31536), .B(n24434), .Z(n24436) );
  XOR U24960 ( .A(a[101]), .B(b[15]), .Z(n24784) );
  NANDN U24961 ( .A(n31925), .B(n24784), .Z(n24435) );
  NAND U24962 ( .A(n24436), .B(n24435), .Z(n24859) );
  XOR U24963 ( .A(n24860), .B(n24859), .Z(n24862) );
  XOR U24964 ( .A(n24861), .B(n24862), .Z(n24926) );
  NANDN U24965 ( .A(n37526), .B(n24437), .Z(n24439) );
  XOR U24966 ( .A(b[51]), .B(a[65]), .Z(n24787) );
  NANDN U24967 ( .A(n37605), .B(n24787), .Z(n24438) );
  AND U24968 ( .A(n24439), .B(n24438), .Z(n24885) );
  NANDN U24969 ( .A(n37705), .B(n24440), .Z(n24442) );
  XOR U24970 ( .A(b[53]), .B(a[63]), .Z(n24790) );
  NANDN U24971 ( .A(n37778), .B(n24790), .Z(n24441) );
  AND U24972 ( .A(n24442), .B(n24441), .Z(n24884) );
  NANDN U24973 ( .A(n36210), .B(n24443), .Z(n24445) );
  XOR U24974 ( .A(b[39]), .B(a[77]), .Z(n24793) );
  NANDN U24975 ( .A(n36347), .B(n24793), .Z(n24444) );
  NAND U24976 ( .A(n24445), .B(n24444), .Z(n24883) );
  XOR U24977 ( .A(n24884), .B(n24883), .Z(n24886) );
  XNOR U24978 ( .A(n24885), .B(n24886), .Z(n24925) );
  XNOR U24979 ( .A(n24926), .B(n24925), .Z(n24928) );
  NANDN U24980 ( .A(n24447), .B(n24446), .Z(n24451) );
  OR U24981 ( .A(n24449), .B(n24448), .Z(n24450) );
  AND U24982 ( .A(n24451), .B(n24450), .Z(n24927) );
  XOR U24983 ( .A(n24928), .B(n24927), .Z(n24769) );
  NANDN U24984 ( .A(n24453), .B(n24452), .Z(n24457) );
  OR U24985 ( .A(n24455), .B(n24454), .Z(n24456) );
  AND U24986 ( .A(n24457), .B(n24456), .Z(n24767) );
  NANDN U24987 ( .A(n24459), .B(n24458), .Z(n24463) );
  NANDN U24988 ( .A(n24461), .B(n24460), .Z(n24462) );
  NAND U24989 ( .A(n24463), .B(n24462), .Z(n24766) );
  XNOR U24990 ( .A(n24767), .B(n24766), .Z(n24768) );
  XNOR U24991 ( .A(n24769), .B(n24768), .Z(n24697) );
  XOR U24992 ( .A(n24698), .B(n24697), .Z(n24700) );
  XOR U24993 ( .A(n24699), .B(n24700), .Z(n24704) );
  NANDN U24994 ( .A(n24465), .B(n24464), .Z(n24469) );
  NANDN U24995 ( .A(n24467), .B(n24466), .Z(n24468) );
  AND U24996 ( .A(n24469), .B(n24468), .Z(n24692) );
  NANDN U24997 ( .A(n211), .B(n24470), .Z(n24472) );
  XOR U24998 ( .A(b[47]), .B(a[69]), .Z(n24721) );
  NANDN U24999 ( .A(n37172), .B(n24721), .Z(n24471) );
  AND U25000 ( .A(n24472), .B(n24471), .Z(n24762) );
  NANDN U25001 ( .A(n210), .B(n24473), .Z(n24475) );
  XOR U25002 ( .A(a[107]), .B(b[9]), .Z(n24724) );
  NANDN U25003 ( .A(n30267), .B(n24724), .Z(n24474) );
  AND U25004 ( .A(n24475), .B(n24474), .Z(n24761) );
  NANDN U25005 ( .A(n212), .B(n24476), .Z(n24478) );
  XOR U25006 ( .A(b[49]), .B(a[67]), .Z(n24727) );
  NANDN U25007 ( .A(n37432), .B(n24727), .Z(n24477) );
  NAND U25008 ( .A(n24478), .B(n24477), .Z(n24760) );
  XOR U25009 ( .A(n24761), .B(n24760), .Z(n24763) );
  XOR U25010 ( .A(n24762), .B(n24763), .Z(n24839) );
  NANDN U25011 ( .A(n36742), .B(n24479), .Z(n24481) );
  XOR U25012 ( .A(b[43]), .B(a[73]), .Z(n24730) );
  NANDN U25013 ( .A(n36891), .B(n24730), .Z(n24480) );
  AND U25014 ( .A(n24481), .B(n24480), .Z(n24741) );
  NANDN U25015 ( .A(n36991), .B(n24482), .Z(n24484) );
  XOR U25016 ( .A(b[45]), .B(a[71]), .Z(n24733) );
  NANDN U25017 ( .A(n37083), .B(n24733), .Z(n24483) );
  AND U25018 ( .A(n24484), .B(n24483), .Z(n24740) );
  NANDN U25019 ( .A(n30482), .B(n24485), .Z(n24487) );
  XOR U25020 ( .A(a[105]), .B(b[11]), .Z(n24736) );
  NANDN U25021 ( .A(n30891), .B(n24736), .Z(n24486) );
  NAND U25022 ( .A(n24487), .B(n24486), .Z(n24739) );
  XOR U25023 ( .A(n24740), .B(n24739), .Z(n24742) );
  XNOR U25024 ( .A(n24741), .B(n24742), .Z(n24838) );
  XNOR U25025 ( .A(n24839), .B(n24838), .Z(n24840) );
  NANDN U25026 ( .A(n24489), .B(n24488), .Z(n24493) );
  OR U25027 ( .A(n24491), .B(n24490), .Z(n24492) );
  NAND U25028 ( .A(n24493), .B(n24492), .Z(n24841) );
  XNOR U25029 ( .A(n24840), .B(n24841), .Z(n24691) );
  XNOR U25030 ( .A(n24692), .B(n24691), .Z(n24693) );
  NANDN U25031 ( .A(n29499), .B(n24494), .Z(n24496) );
  XOR U25032 ( .A(a[109]), .B(b[7]), .Z(n24745) );
  NANDN U25033 ( .A(n29735), .B(n24745), .Z(n24495) );
  AND U25034 ( .A(n24496), .B(n24495), .Z(n24804) );
  NANDN U25035 ( .A(n37857), .B(n24497), .Z(n24499) );
  XOR U25036 ( .A(b[55]), .B(a[61]), .Z(n24748) );
  NANDN U25037 ( .A(n37911), .B(n24748), .Z(n24498) );
  AND U25038 ( .A(n24499), .B(n24498), .Z(n24803) );
  NANDN U25039 ( .A(n35611), .B(n24500), .Z(n24502) );
  XOR U25040 ( .A(b[35]), .B(a[81]), .Z(n24751) );
  NANDN U25041 ( .A(n35801), .B(n24751), .Z(n24501) );
  NAND U25042 ( .A(n24502), .B(n24501), .Z(n24802) );
  XOR U25043 ( .A(n24803), .B(n24802), .Z(n24805) );
  XOR U25044 ( .A(n24804), .B(n24805), .Z(n24821) );
  NANDN U25045 ( .A(n24504), .B(n24503), .Z(n24508) );
  OR U25046 ( .A(n24506), .B(n24505), .Z(n24507) );
  AND U25047 ( .A(n24508), .B(n24507), .Z(n24820) );
  XNOR U25048 ( .A(n24821), .B(n24820), .Z(n24822) );
  NANDN U25049 ( .A(n24510), .B(n24509), .Z(n24514) );
  OR U25050 ( .A(n24512), .B(n24511), .Z(n24513) );
  NAND U25051 ( .A(n24514), .B(n24513), .Z(n24823) );
  XOR U25052 ( .A(n24822), .B(n24823), .Z(n24694) );
  XNOR U25053 ( .A(n24693), .B(n24694), .Z(n24703) );
  XOR U25054 ( .A(n24704), .B(n24703), .Z(n24706) );
  XOR U25055 ( .A(n24705), .B(n24706), .Z(n24938) );
  NANDN U25056 ( .A(n24516), .B(n24515), .Z(n24520) );
  NANDN U25057 ( .A(n24518), .B(n24517), .Z(n24519) );
  AND U25058 ( .A(n24520), .B(n24519), .Z(n24687) );
  NANDN U25059 ( .A(n24522), .B(n24521), .Z(n24526) );
  NANDN U25060 ( .A(n24524), .B(n24523), .Z(n24525) );
  AND U25061 ( .A(n24526), .B(n24525), .Z(n24686) );
  NANDN U25062 ( .A(n24528), .B(n24527), .Z(n24532) );
  NAND U25063 ( .A(n24530), .B(n24529), .Z(n24531) );
  AND U25064 ( .A(n24532), .B(n24531), .Z(n24685) );
  XOR U25065 ( .A(n24686), .B(n24685), .Z(n24688) );
  XOR U25066 ( .A(n24687), .B(n24688), .Z(n24712) );
  NANDN U25067 ( .A(n24534), .B(n24533), .Z(n24538) );
  NANDN U25068 ( .A(n24536), .B(n24535), .Z(n24537) );
  AND U25069 ( .A(n24538), .B(n24537), .Z(n24934) );
  NANDN U25070 ( .A(n32996), .B(n24539), .Z(n24541) );
  XOR U25071 ( .A(a[95]), .B(b[21]), .Z(n24844) );
  NANDN U25072 ( .A(n33271), .B(n24844), .Z(n24540) );
  AND U25073 ( .A(n24541), .B(n24540), .Z(n24903) );
  NANDN U25074 ( .A(n33866), .B(n24542), .Z(n24544) );
  XOR U25075 ( .A(a[93]), .B(b[23]), .Z(n24847) );
  NANDN U25076 ( .A(n33644), .B(n24847), .Z(n24543) );
  AND U25077 ( .A(n24544), .B(n24543), .Z(n24902) );
  NANDN U25078 ( .A(n32483), .B(n24545), .Z(n24547) );
  XOR U25079 ( .A(a[97]), .B(b[19]), .Z(n24850) );
  NANDN U25080 ( .A(n32823), .B(n24850), .Z(n24546) );
  NAND U25081 ( .A(n24547), .B(n24546), .Z(n24901) );
  XOR U25082 ( .A(n24902), .B(n24901), .Z(n24904) );
  XOR U25083 ( .A(n24903), .B(n24904), .Z(n24716) );
  NANDN U25084 ( .A(n34909), .B(n24548), .Z(n24550) );
  XOR U25085 ( .A(b[31]), .B(a[85]), .Z(n24853) );
  NANDN U25086 ( .A(n35145), .B(n24853), .Z(n24549) );
  AND U25087 ( .A(n24550), .B(n24549), .Z(n24756) );
  NANDN U25088 ( .A(n38247), .B(n24551), .Z(n24553) );
  XOR U25089 ( .A(b[61]), .B(a[55]), .Z(n24856) );
  NANDN U25090 ( .A(n38248), .B(n24856), .Z(n24552) );
  AND U25091 ( .A(n24553), .B(n24552), .Z(n24755) );
  AND U25092 ( .A(b[63]), .B(a[51]), .Z(n24754) );
  XOR U25093 ( .A(n24755), .B(n24754), .Z(n24757) );
  XNOR U25094 ( .A(n24756), .B(n24757), .Z(n24715) );
  XNOR U25095 ( .A(n24716), .B(n24715), .Z(n24717) );
  NANDN U25096 ( .A(n24555), .B(n24554), .Z(n24559) );
  OR U25097 ( .A(n24557), .B(n24556), .Z(n24558) );
  NAND U25098 ( .A(n24559), .B(n24558), .Z(n24718) );
  XNOR U25099 ( .A(n24717), .B(n24718), .Z(n24931) );
  NANDN U25100 ( .A(n34223), .B(n24560), .Z(n24562) );
  XOR U25101 ( .A(b[27]), .B(a[89]), .Z(n24865) );
  NANDN U25102 ( .A(n34458), .B(n24865), .Z(n24561) );
  AND U25103 ( .A(n24562), .B(n24561), .Z(n24798) );
  NANDN U25104 ( .A(n34634), .B(n24563), .Z(n24565) );
  XOR U25105 ( .A(b[29]), .B(a[87]), .Z(n24868) );
  NANDN U25106 ( .A(n34722), .B(n24868), .Z(n24564) );
  AND U25107 ( .A(n24565), .B(n24564), .Z(n24797) );
  NANDN U25108 ( .A(n31055), .B(n24566), .Z(n24568) );
  XOR U25109 ( .A(a[103]), .B(b[13]), .Z(n24871) );
  NANDN U25110 ( .A(n31293), .B(n24871), .Z(n24567) );
  NAND U25111 ( .A(n24568), .B(n24567), .Z(n24796) );
  XOR U25112 ( .A(n24797), .B(n24796), .Z(n24799) );
  XOR U25113 ( .A(n24798), .B(n24799), .Z(n24827) );
  NANDN U25114 ( .A(n28889), .B(n24569), .Z(n24571) );
  XOR U25115 ( .A(a[111]), .B(b[5]), .Z(n24874) );
  NANDN U25116 ( .A(n29138), .B(n24874), .Z(n24570) );
  AND U25117 ( .A(n24571), .B(n24570), .Z(n24897) );
  NANDN U25118 ( .A(n209), .B(n24572), .Z(n24574) );
  XOR U25119 ( .A(a[113]), .B(b[3]), .Z(n24877) );
  NANDN U25120 ( .A(n28941), .B(n24877), .Z(n24573) );
  AND U25121 ( .A(n24574), .B(n24573), .Z(n24896) );
  NANDN U25122 ( .A(n35936), .B(n24575), .Z(n24577) );
  XOR U25123 ( .A(b[37]), .B(a[79]), .Z(n24880) );
  NANDN U25124 ( .A(n36047), .B(n24880), .Z(n24576) );
  NAND U25125 ( .A(n24577), .B(n24576), .Z(n24895) );
  XOR U25126 ( .A(n24896), .B(n24895), .Z(n24898) );
  XNOR U25127 ( .A(n24897), .B(n24898), .Z(n24826) );
  XNOR U25128 ( .A(n24827), .B(n24826), .Z(n24828) );
  NANDN U25129 ( .A(n24579), .B(n24578), .Z(n24583) );
  OR U25130 ( .A(n24581), .B(n24580), .Z(n24582) );
  NAND U25131 ( .A(n24583), .B(n24582), .Z(n24829) );
  XOR U25132 ( .A(n24828), .B(n24829), .Z(n24932) );
  XNOR U25133 ( .A(n24931), .B(n24932), .Z(n24933) );
  XNOR U25134 ( .A(n24934), .B(n24933), .Z(n24817) );
  NANDN U25135 ( .A(n24585), .B(n24584), .Z(n24589) );
  NANDN U25136 ( .A(n24587), .B(n24586), .Z(n24588) );
  AND U25137 ( .A(n24589), .B(n24588), .Z(n24833) );
  NANDN U25138 ( .A(n24591), .B(n24590), .Z(n24595) );
  OR U25139 ( .A(n24593), .B(n24592), .Z(n24594) );
  NAND U25140 ( .A(n24595), .B(n24594), .Z(n24832) );
  XNOR U25141 ( .A(n24833), .B(n24832), .Z(n24835) );
  NANDN U25142 ( .A(n24597), .B(n24596), .Z(n24601) );
  OR U25143 ( .A(n24599), .B(n24598), .Z(n24600) );
  AND U25144 ( .A(n24601), .B(n24600), .Z(n24775) );
  NAND U25145 ( .A(b[0]), .B(a[115]), .Z(n24602) );
  XNOR U25146 ( .A(b[1]), .B(n24602), .Z(n24604) );
  NANDN U25147 ( .A(b[0]), .B(a[114]), .Z(n24603) );
  NAND U25148 ( .A(n24604), .B(n24603), .Z(n24811) );
  NANDN U25149 ( .A(n38278), .B(n24605), .Z(n24607) );
  XOR U25150 ( .A(b[63]), .B(a[53]), .Z(n24910) );
  NANDN U25151 ( .A(n38279), .B(n24910), .Z(n24606) );
  AND U25152 ( .A(n24607), .B(n24606), .Z(n24809) );
  NANDN U25153 ( .A(n35260), .B(n24608), .Z(n24610) );
  XOR U25154 ( .A(b[33]), .B(a[83]), .Z(n24913) );
  NANDN U25155 ( .A(n35456), .B(n24913), .Z(n24609) );
  NAND U25156 ( .A(n24610), .B(n24609), .Z(n24808) );
  XNOR U25157 ( .A(n24809), .B(n24808), .Z(n24810) );
  XNOR U25158 ( .A(n24811), .B(n24810), .Z(n24772) );
  NANDN U25159 ( .A(n37974), .B(n24611), .Z(n24613) );
  XOR U25160 ( .A(b[57]), .B(a[59]), .Z(n24916) );
  NANDN U25161 ( .A(n38031), .B(n24916), .Z(n24612) );
  AND U25162 ( .A(n24613), .B(n24612), .Z(n24892) );
  NANDN U25163 ( .A(n38090), .B(n24614), .Z(n24616) );
  XOR U25164 ( .A(b[59]), .B(a[57]), .Z(n24919) );
  NANDN U25165 ( .A(n38130), .B(n24919), .Z(n24615) );
  AND U25166 ( .A(n24616), .B(n24615), .Z(n24890) );
  NANDN U25167 ( .A(n36480), .B(n24617), .Z(n24619) );
  XOR U25168 ( .A(b[41]), .B(a[75]), .Z(n24922) );
  NANDN U25169 ( .A(n36594), .B(n24922), .Z(n24618) );
  NAND U25170 ( .A(n24619), .B(n24618), .Z(n24889) );
  XNOR U25171 ( .A(n24890), .B(n24889), .Z(n24891) );
  XOR U25172 ( .A(n24892), .B(n24891), .Z(n24773) );
  XNOR U25173 ( .A(n24772), .B(n24773), .Z(n24774) );
  XNOR U25174 ( .A(n24775), .B(n24774), .Z(n24834) );
  XOR U25175 ( .A(n24835), .B(n24834), .Z(n24815) );
  NANDN U25176 ( .A(n24621), .B(n24620), .Z(n24625) );
  NAND U25177 ( .A(n24623), .B(n24622), .Z(n24624) );
  NAND U25178 ( .A(n24625), .B(n24624), .Z(n24814) );
  XNOR U25179 ( .A(n24815), .B(n24814), .Z(n24816) );
  XOR U25180 ( .A(n24817), .B(n24816), .Z(n24710) );
  NANDN U25181 ( .A(n24627), .B(n24626), .Z(n24631) );
  NANDN U25182 ( .A(n24629), .B(n24628), .Z(n24630) );
  AND U25183 ( .A(n24631), .B(n24630), .Z(n24709) );
  XNOR U25184 ( .A(n24710), .B(n24709), .Z(n24711) );
  XNOR U25185 ( .A(n24712), .B(n24711), .Z(n24937) );
  XOR U25186 ( .A(n24938), .B(n24937), .Z(n24940) );
  XOR U25187 ( .A(n24939), .B(n24940), .Z(n24951) );
  NANDN U25188 ( .A(n24633), .B(n24632), .Z(n24637) );
  OR U25189 ( .A(n24635), .B(n24634), .Z(n24636) );
  AND U25190 ( .A(n24637), .B(n24636), .Z(n24950) );
  NANDN U25191 ( .A(n24639), .B(n24638), .Z(n24643) );
  OR U25192 ( .A(n24641), .B(n24640), .Z(n24642) );
  AND U25193 ( .A(n24643), .B(n24642), .Z(n24946) );
  NANDN U25194 ( .A(n24645), .B(n24644), .Z(n24649) );
  NANDN U25195 ( .A(n24647), .B(n24646), .Z(n24648) );
  AND U25196 ( .A(n24649), .B(n24648), .Z(n24944) );
  NANDN U25197 ( .A(n24651), .B(n24650), .Z(n24655) );
  OR U25198 ( .A(n24653), .B(n24652), .Z(n24654) );
  AND U25199 ( .A(n24655), .B(n24654), .Z(n24943) );
  XNOR U25200 ( .A(n24944), .B(n24943), .Z(n24945) );
  XNOR U25201 ( .A(n24946), .B(n24945), .Z(n24949) );
  XOR U25202 ( .A(n24950), .B(n24949), .Z(n24952) );
  XOR U25203 ( .A(n24951), .B(n24952), .Z(n24958) );
  NANDN U25204 ( .A(n24657), .B(n24656), .Z(n24661) );
  NANDN U25205 ( .A(n24659), .B(n24658), .Z(n24660) );
  AND U25206 ( .A(n24661), .B(n24660), .Z(n24956) );
  NANDN U25207 ( .A(n24663), .B(n24662), .Z(n24667) );
  OR U25208 ( .A(n24665), .B(n24664), .Z(n24666) );
  AND U25209 ( .A(n24667), .B(n24666), .Z(n24955) );
  XNOR U25210 ( .A(n24956), .B(n24955), .Z(n24957) );
  XNOR U25211 ( .A(n24958), .B(n24957), .Z(n24961) );
  XOR U25212 ( .A(n24962), .B(n24961), .Z(n24964) );
  XOR U25213 ( .A(n24963), .B(n24964), .Z(n24680) );
  NANDN U25214 ( .A(n24669), .B(n24668), .Z(n24673) );
  NANDN U25215 ( .A(n24671), .B(n24670), .Z(n24672) );
  NAND U25216 ( .A(n24673), .B(n24672), .Z(n24679) );
  XNOR U25217 ( .A(n24680), .B(n24679), .Z(n24681) );
  XNOR U25218 ( .A(n24682), .B(n24681), .Z(n24967) );
  XNOR U25219 ( .A(sreg[179]), .B(n24967), .Z(n24969) );
  NANDN U25220 ( .A(sreg[178]), .B(n24674), .Z(n24678) );
  NAND U25221 ( .A(n24676), .B(n24675), .Z(n24677) );
  NAND U25222 ( .A(n24678), .B(n24677), .Z(n24968) );
  XNOR U25223 ( .A(n24969), .B(n24968), .Z(c[179]) );
  NANDN U25224 ( .A(n24680), .B(n24679), .Z(n24684) );
  NANDN U25225 ( .A(n24682), .B(n24681), .Z(n24683) );
  AND U25226 ( .A(n24684), .B(n24683), .Z(n24975) );
  NANDN U25227 ( .A(n24686), .B(n24685), .Z(n24690) );
  OR U25228 ( .A(n24688), .B(n24687), .Z(n24689) );
  AND U25229 ( .A(n24690), .B(n24689), .Z(n24992) );
  NANDN U25230 ( .A(n24692), .B(n24691), .Z(n24696) );
  NANDN U25231 ( .A(n24694), .B(n24693), .Z(n24695) );
  AND U25232 ( .A(n24696), .B(n24695), .Z(n24991) );
  NANDN U25233 ( .A(n24698), .B(n24697), .Z(n24702) );
  OR U25234 ( .A(n24700), .B(n24699), .Z(n24701) );
  AND U25235 ( .A(n24702), .B(n24701), .Z(n24990) );
  XOR U25236 ( .A(n24991), .B(n24990), .Z(n24993) );
  XOR U25237 ( .A(n24992), .B(n24993), .Z(n25249) );
  NANDN U25238 ( .A(n24704), .B(n24703), .Z(n24708) );
  OR U25239 ( .A(n24706), .B(n24705), .Z(n24707) );
  AND U25240 ( .A(n24708), .B(n24707), .Z(n25248) );
  XNOR U25241 ( .A(n25249), .B(n25248), .Z(n25250) );
  NANDN U25242 ( .A(n24710), .B(n24709), .Z(n24714) );
  NANDN U25243 ( .A(n24712), .B(n24711), .Z(n24713) );
  AND U25244 ( .A(n24714), .B(n24713), .Z(n24987) );
  NANDN U25245 ( .A(n24716), .B(n24715), .Z(n24720) );
  NANDN U25246 ( .A(n24718), .B(n24717), .Z(n24719) );
  AND U25247 ( .A(n24720), .B(n24719), .Z(n25003) );
  NAND U25248 ( .A(n37294), .B(n24721), .Z(n24723) );
  XNOR U25249 ( .A(b[47]), .B(a[70]), .Z(n25086) );
  NANDN U25250 ( .A(n25086), .B(n37341), .Z(n24722) );
  NAND U25251 ( .A(n24723), .B(n24722), .Z(n25127) );
  NAND U25252 ( .A(n30627), .B(n24724), .Z(n24726) );
  XNOR U25253 ( .A(a[108]), .B(b[9]), .Z(n25089) );
  NANDN U25254 ( .A(n25089), .B(n30628), .Z(n24725) );
  NAND U25255 ( .A(n24726), .B(n24725), .Z(n25126) );
  NAND U25256 ( .A(n37536), .B(n24727), .Z(n24729) );
  XNOR U25257 ( .A(b[49]), .B(a[68]), .Z(n25092) );
  NANDN U25258 ( .A(n25092), .B(n37537), .Z(n24728) );
  NAND U25259 ( .A(n24729), .B(n24728), .Z(n25125) );
  XNOR U25260 ( .A(n25126), .B(n25125), .Z(n25128) );
  NANDN U25261 ( .A(n36742), .B(n24730), .Z(n24732) );
  XOR U25262 ( .A(b[43]), .B(a[74]), .Z(n25095) );
  NANDN U25263 ( .A(n36891), .B(n25095), .Z(n24731) );
  AND U25264 ( .A(n24732), .B(n24731), .Z(n25106) );
  NANDN U25265 ( .A(n36991), .B(n24733), .Z(n24735) );
  XOR U25266 ( .A(b[45]), .B(a[72]), .Z(n25098) );
  NANDN U25267 ( .A(n37083), .B(n25098), .Z(n24734) );
  AND U25268 ( .A(n24735), .B(n24734), .Z(n25105) );
  NANDN U25269 ( .A(n30482), .B(n24736), .Z(n24738) );
  XOR U25270 ( .A(a[106]), .B(b[11]), .Z(n25101) );
  NANDN U25271 ( .A(n30891), .B(n25101), .Z(n24737) );
  NAND U25272 ( .A(n24738), .B(n24737), .Z(n25104) );
  XOR U25273 ( .A(n25105), .B(n25104), .Z(n25107) );
  XNOR U25274 ( .A(n25106), .B(n25107), .Z(n25191) );
  XOR U25275 ( .A(n25192), .B(n25191), .Z(n25193) );
  NANDN U25276 ( .A(n24740), .B(n24739), .Z(n24744) );
  OR U25277 ( .A(n24742), .B(n24741), .Z(n24743) );
  NAND U25278 ( .A(n24744), .B(n24743), .Z(n25194) );
  XNOR U25279 ( .A(n25193), .B(n25194), .Z(n25002) );
  XNOR U25280 ( .A(n25003), .B(n25002), .Z(n25005) );
  NANDN U25281 ( .A(n29499), .B(n24745), .Z(n24747) );
  XOR U25282 ( .A(a[110]), .B(b[7]), .Z(n25110) );
  NANDN U25283 ( .A(n29735), .B(n25110), .Z(n24746) );
  AND U25284 ( .A(n24747), .B(n24746), .Z(n25070) );
  NANDN U25285 ( .A(n37857), .B(n24748), .Z(n24750) );
  XOR U25286 ( .A(b[55]), .B(a[62]), .Z(n25113) );
  NANDN U25287 ( .A(n37911), .B(n25113), .Z(n24749) );
  AND U25288 ( .A(n24750), .B(n24749), .Z(n25069) );
  NANDN U25289 ( .A(n35611), .B(n24751), .Z(n24753) );
  XOR U25290 ( .A(b[35]), .B(a[82]), .Z(n25116) );
  NANDN U25291 ( .A(n35801), .B(n25116), .Z(n24752) );
  NAND U25292 ( .A(n24753), .B(n24752), .Z(n25068) );
  XOR U25293 ( .A(n25069), .B(n25068), .Z(n25071) );
  XOR U25294 ( .A(n25070), .B(n25071), .Z(n25132) );
  NANDN U25295 ( .A(n24755), .B(n24754), .Z(n24759) );
  OR U25296 ( .A(n24757), .B(n24756), .Z(n24758) );
  AND U25297 ( .A(n24759), .B(n24758), .Z(n25131) );
  XNOR U25298 ( .A(n25132), .B(n25131), .Z(n25133) );
  NANDN U25299 ( .A(n24761), .B(n24760), .Z(n24765) );
  OR U25300 ( .A(n24763), .B(n24762), .Z(n24764) );
  NAND U25301 ( .A(n24765), .B(n24764), .Z(n25134) );
  XNOR U25302 ( .A(n25133), .B(n25134), .Z(n25004) );
  XOR U25303 ( .A(n25005), .B(n25004), .Z(n25015) );
  NANDN U25304 ( .A(n24767), .B(n24766), .Z(n24771) );
  NANDN U25305 ( .A(n24769), .B(n24768), .Z(n24770) );
  AND U25306 ( .A(n24771), .B(n24770), .Z(n25011) );
  NANDN U25307 ( .A(n24773), .B(n24772), .Z(n24777) );
  NANDN U25308 ( .A(n24775), .B(n24774), .Z(n24776) );
  AND U25309 ( .A(n24777), .B(n24776), .Z(n25009) );
  NANDN U25310 ( .A(n33875), .B(n24778), .Z(n24780) );
  XOR U25311 ( .A(a[92]), .B(b[25]), .Z(n25044) );
  NANDN U25312 ( .A(n33994), .B(n25044), .Z(n24779) );
  AND U25313 ( .A(n24780), .B(n24779), .Z(n25223) );
  NANDN U25314 ( .A(n32013), .B(n24781), .Z(n24783) );
  XOR U25315 ( .A(a[100]), .B(b[17]), .Z(n25047) );
  NANDN U25316 ( .A(n32292), .B(n25047), .Z(n24782) );
  AND U25317 ( .A(n24783), .B(n24782), .Z(n25222) );
  NANDN U25318 ( .A(n31536), .B(n24784), .Z(n24786) );
  XOR U25319 ( .A(a[102]), .B(b[15]), .Z(n25050) );
  NANDN U25320 ( .A(n31925), .B(n25050), .Z(n24785) );
  NAND U25321 ( .A(n24786), .B(n24785), .Z(n25221) );
  XOR U25322 ( .A(n25222), .B(n25221), .Z(n25224) );
  XOR U25323 ( .A(n25223), .B(n25224), .Z(n25186) );
  NANDN U25324 ( .A(n37526), .B(n24787), .Z(n24789) );
  XOR U25325 ( .A(b[51]), .B(a[66]), .Z(n25053) );
  NANDN U25326 ( .A(n37605), .B(n25053), .Z(n24788) );
  AND U25327 ( .A(n24789), .B(n24788), .Z(n25199) );
  NANDN U25328 ( .A(n37705), .B(n24790), .Z(n24792) );
  XOR U25329 ( .A(b[53]), .B(a[64]), .Z(n25056) );
  NANDN U25330 ( .A(n37778), .B(n25056), .Z(n24791) );
  AND U25331 ( .A(n24792), .B(n24791), .Z(n25198) );
  NANDN U25332 ( .A(n36210), .B(n24793), .Z(n24795) );
  XOR U25333 ( .A(b[39]), .B(a[78]), .Z(n25059) );
  NANDN U25334 ( .A(n36347), .B(n25059), .Z(n24794) );
  NAND U25335 ( .A(n24795), .B(n24794), .Z(n25197) );
  XOR U25336 ( .A(n25198), .B(n25197), .Z(n25200) );
  XNOR U25337 ( .A(n25199), .B(n25200), .Z(n25185) );
  XNOR U25338 ( .A(n25186), .B(n25185), .Z(n25188) );
  NANDN U25339 ( .A(n24797), .B(n24796), .Z(n24801) );
  OR U25340 ( .A(n24799), .B(n24798), .Z(n24800) );
  AND U25341 ( .A(n24801), .B(n24800), .Z(n25187) );
  XOR U25342 ( .A(n25188), .B(n25187), .Z(n25035) );
  NANDN U25343 ( .A(n24803), .B(n24802), .Z(n24807) );
  OR U25344 ( .A(n24805), .B(n24804), .Z(n24806) );
  AND U25345 ( .A(n24807), .B(n24806), .Z(n25033) );
  NANDN U25346 ( .A(n24809), .B(n24808), .Z(n24813) );
  NANDN U25347 ( .A(n24811), .B(n24810), .Z(n24812) );
  NAND U25348 ( .A(n24813), .B(n24812), .Z(n25032) );
  XNOR U25349 ( .A(n25033), .B(n25032), .Z(n25034) );
  XNOR U25350 ( .A(n25035), .B(n25034), .Z(n25008) );
  XNOR U25351 ( .A(n25009), .B(n25008), .Z(n25010) );
  XNOR U25352 ( .A(n25011), .B(n25010), .Z(n25014) );
  XNOR U25353 ( .A(n25015), .B(n25014), .Z(n25016) );
  NANDN U25354 ( .A(n24815), .B(n24814), .Z(n24819) );
  NAND U25355 ( .A(n24817), .B(n24816), .Z(n24818) );
  NAND U25356 ( .A(n24819), .B(n24818), .Z(n25017) );
  XNOR U25357 ( .A(n25016), .B(n25017), .Z(n24984) );
  NANDN U25358 ( .A(n24821), .B(n24820), .Z(n24825) );
  NANDN U25359 ( .A(n24823), .B(n24822), .Z(n24824) );
  AND U25360 ( .A(n24825), .B(n24824), .Z(n24998) );
  NANDN U25361 ( .A(n24827), .B(n24826), .Z(n24831) );
  NANDN U25362 ( .A(n24829), .B(n24828), .Z(n24830) );
  AND U25363 ( .A(n24831), .B(n24830), .Z(n24997) );
  NANDN U25364 ( .A(n24833), .B(n24832), .Z(n24837) );
  NAND U25365 ( .A(n24835), .B(n24834), .Z(n24836) );
  AND U25366 ( .A(n24837), .B(n24836), .Z(n24996) );
  XOR U25367 ( .A(n24997), .B(n24996), .Z(n24999) );
  XOR U25368 ( .A(n24998), .B(n24999), .Z(n25023) );
  NANDN U25369 ( .A(n24839), .B(n24838), .Z(n24843) );
  NANDN U25370 ( .A(n24841), .B(n24840), .Z(n24842) );
  AND U25371 ( .A(n24843), .B(n24842), .Z(n25245) );
  NANDN U25372 ( .A(n32996), .B(n24844), .Z(n24846) );
  XOR U25373 ( .A(a[96]), .B(b[21]), .Z(n25227) );
  NANDN U25374 ( .A(n33271), .B(n25227), .Z(n24845) );
  AND U25375 ( .A(n24846), .B(n24845), .Z(n25163) );
  NANDN U25376 ( .A(n33866), .B(n24847), .Z(n24849) );
  XOR U25377 ( .A(a[94]), .B(b[23]), .Z(n25230) );
  NANDN U25378 ( .A(n33644), .B(n25230), .Z(n24848) );
  AND U25379 ( .A(n24849), .B(n24848), .Z(n25162) );
  NANDN U25380 ( .A(n32483), .B(n24850), .Z(n24852) );
  XOR U25381 ( .A(a[98]), .B(b[19]), .Z(n25233) );
  NANDN U25382 ( .A(n32823), .B(n25233), .Z(n24851) );
  NAND U25383 ( .A(n24852), .B(n24851), .Z(n25161) );
  XOR U25384 ( .A(n25162), .B(n25161), .Z(n25164) );
  XOR U25385 ( .A(n25163), .B(n25164), .Z(n25081) );
  NANDN U25386 ( .A(n34909), .B(n24853), .Z(n24855) );
  XOR U25387 ( .A(b[31]), .B(a[86]), .Z(n25236) );
  NANDN U25388 ( .A(n35145), .B(n25236), .Z(n24854) );
  AND U25389 ( .A(n24855), .B(n24854), .Z(n25121) );
  NANDN U25390 ( .A(n38247), .B(n24856), .Z(n24858) );
  XOR U25391 ( .A(b[61]), .B(a[56]), .Z(n25239) );
  NANDN U25392 ( .A(n38248), .B(n25239), .Z(n24857) );
  AND U25393 ( .A(n24858), .B(n24857), .Z(n25120) );
  AND U25394 ( .A(b[63]), .B(a[52]), .Z(n25119) );
  XOR U25395 ( .A(n25120), .B(n25119), .Z(n25122) );
  XNOR U25396 ( .A(n25121), .B(n25122), .Z(n25080) );
  XNOR U25397 ( .A(n25081), .B(n25080), .Z(n25082) );
  NANDN U25398 ( .A(n24860), .B(n24859), .Z(n24864) );
  OR U25399 ( .A(n24862), .B(n24861), .Z(n24863) );
  NAND U25400 ( .A(n24864), .B(n24863), .Z(n25083) );
  XNOR U25401 ( .A(n25082), .B(n25083), .Z(n25242) );
  NANDN U25402 ( .A(n34223), .B(n24865), .Z(n24867) );
  XOR U25403 ( .A(b[27]), .B(a[90]), .Z(n25203) );
  NANDN U25404 ( .A(n34458), .B(n25203), .Z(n24866) );
  AND U25405 ( .A(n24867), .B(n24866), .Z(n25064) );
  NANDN U25406 ( .A(n34634), .B(n24868), .Z(n24870) );
  XOR U25407 ( .A(b[29]), .B(a[88]), .Z(n25206) );
  NANDN U25408 ( .A(n34722), .B(n25206), .Z(n24869) );
  AND U25409 ( .A(n24870), .B(n24869), .Z(n25063) );
  NANDN U25410 ( .A(n31055), .B(n24871), .Z(n24873) );
  XOR U25411 ( .A(a[104]), .B(b[13]), .Z(n25209) );
  NANDN U25412 ( .A(n31293), .B(n25209), .Z(n24872) );
  NAND U25413 ( .A(n24873), .B(n24872), .Z(n25062) );
  XOR U25414 ( .A(n25063), .B(n25062), .Z(n25065) );
  XOR U25415 ( .A(n25064), .B(n25065), .Z(n25138) );
  NANDN U25416 ( .A(n28889), .B(n24874), .Z(n24876) );
  XOR U25417 ( .A(a[112]), .B(b[5]), .Z(n25212) );
  NANDN U25418 ( .A(n29138), .B(n25212), .Z(n24875) );
  AND U25419 ( .A(n24876), .B(n24875), .Z(n25157) );
  NANDN U25420 ( .A(n209), .B(n24877), .Z(n24879) );
  XOR U25421 ( .A(a[114]), .B(b[3]), .Z(n25215) );
  NANDN U25422 ( .A(n28941), .B(n25215), .Z(n24878) );
  AND U25423 ( .A(n24879), .B(n24878), .Z(n25156) );
  NANDN U25424 ( .A(n35936), .B(n24880), .Z(n24882) );
  XOR U25425 ( .A(b[37]), .B(a[80]), .Z(n25218) );
  NANDN U25426 ( .A(n36047), .B(n25218), .Z(n24881) );
  NAND U25427 ( .A(n24882), .B(n24881), .Z(n25155) );
  XOR U25428 ( .A(n25156), .B(n25155), .Z(n25158) );
  XNOR U25429 ( .A(n25157), .B(n25158), .Z(n25137) );
  XNOR U25430 ( .A(n25138), .B(n25137), .Z(n25139) );
  NANDN U25431 ( .A(n24884), .B(n24883), .Z(n24888) );
  OR U25432 ( .A(n24886), .B(n24885), .Z(n24887) );
  NAND U25433 ( .A(n24888), .B(n24887), .Z(n25140) );
  XOR U25434 ( .A(n25139), .B(n25140), .Z(n25243) );
  XNOR U25435 ( .A(n25242), .B(n25243), .Z(n25244) );
  XNOR U25436 ( .A(n25245), .B(n25244), .Z(n25029) );
  NANDN U25437 ( .A(n24890), .B(n24889), .Z(n24894) );
  NANDN U25438 ( .A(n24892), .B(n24891), .Z(n24893) );
  AND U25439 ( .A(n24894), .B(n24893), .Z(n25144) );
  NANDN U25440 ( .A(n24896), .B(n24895), .Z(n24900) );
  OR U25441 ( .A(n24898), .B(n24897), .Z(n24899) );
  NAND U25442 ( .A(n24900), .B(n24899), .Z(n25143) );
  XNOR U25443 ( .A(n25144), .B(n25143), .Z(n25146) );
  NANDN U25444 ( .A(n24902), .B(n24901), .Z(n24906) );
  OR U25445 ( .A(n24904), .B(n24903), .Z(n24905) );
  AND U25446 ( .A(n24906), .B(n24905), .Z(n25041) );
  NAND U25447 ( .A(b[0]), .B(a[116]), .Z(n24907) );
  XNOR U25448 ( .A(b[1]), .B(n24907), .Z(n24909) );
  NANDN U25449 ( .A(b[0]), .B(a[115]), .Z(n24908) );
  NAND U25450 ( .A(n24909), .B(n24908), .Z(n25077) );
  NANDN U25451 ( .A(n38278), .B(n24910), .Z(n24912) );
  XOR U25452 ( .A(b[63]), .B(a[54]), .Z(n25170) );
  NANDN U25453 ( .A(n38279), .B(n25170), .Z(n24911) );
  AND U25454 ( .A(n24912), .B(n24911), .Z(n25075) );
  NANDN U25455 ( .A(n35260), .B(n24913), .Z(n24915) );
  XOR U25456 ( .A(b[33]), .B(a[84]), .Z(n25173) );
  NANDN U25457 ( .A(n35456), .B(n25173), .Z(n24914) );
  NAND U25458 ( .A(n24915), .B(n24914), .Z(n25074) );
  XNOR U25459 ( .A(n25075), .B(n25074), .Z(n25076) );
  XNOR U25460 ( .A(n25077), .B(n25076), .Z(n25038) );
  NANDN U25461 ( .A(n37974), .B(n24916), .Z(n24918) );
  XOR U25462 ( .A(b[57]), .B(a[60]), .Z(n25176) );
  NANDN U25463 ( .A(n38031), .B(n25176), .Z(n24917) );
  AND U25464 ( .A(n24918), .B(n24917), .Z(n25152) );
  NANDN U25465 ( .A(n38090), .B(n24919), .Z(n24921) );
  XOR U25466 ( .A(b[59]), .B(a[58]), .Z(n25179) );
  NANDN U25467 ( .A(n38130), .B(n25179), .Z(n24920) );
  AND U25468 ( .A(n24921), .B(n24920), .Z(n25150) );
  NANDN U25469 ( .A(n36480), .B(n24922), .Z(n24924) );
  XOR U25470 ( .A(b[41]), .B(a[76]), .Z(n25182) );
  NANDN U25471 ( .A(n36594), .B(n25182), .Z(n24923) );
  NAND U25472 ( .A(n24924), .B(n24923), .Z(n25149) );
  XNOR U25473 ( .A(n25150), .B(n25149), .Z(n25151) );
  XOR U25474 ( .A(n25152), .B(n25151), .Z(n25039) );
  XNOR U25475 ( .A(n25038), .B(n25039), .Z(n25040) );
  XNOR U25476 ( .A(n25041), .B(n25040), .Z(n25145) );
  XOR U25477 ( .A(n25146), .B(n25145), .Z(n25027) );
  NANDN U25478 ( .A(n24926), .B(n24925), .Z(n24930) );
  NAND U25479 ( .A(n24928), .B(n24927), .Z(n24929) );
  NAND U25480 ( .A(n24930), .B(n24929), .Z(n25026) );
  XNOR U25481 ( .A(n25027), .B(n25026), .Z(n25028) );
  XOR U25482 ( .A(n25029), .B(n25028), .Z(n25021) );
  NANDN U25483 ( .A(n24932), .B(n24931), .Z(n24936) );
  NANDN U25484 ( .A(n24934), .B(n24933), .Z(n24935) );
  AND U25485 ( .A(n24936), .B(n24935), .Z(n25020) );
  XNOR U25486 ( .A(n25021), .B(n25020), .Z(n25022) );
  XOR U25487 ( .A(n25023), .B(n25022), .Z(n24985) );
  XNOR U25488 ( .A(n24984), .B(n24985), .Z(n24986) );
  XOR U25489 ( .A(n24987), .B(n24986), .Z(n25251) );
  XNOR U25490 ( .A(n25250), .B(n25251), .Z(n25257) );
  NANDN U25491 ( .A(n24938), .B(n24937), .Z(n24942) );
  OR U25492 ( .A(n24940), .B(n24939), .Z(n24941) );
  AND U25493 ( .A(n24942), .B(n24941), .Z(n25255) );
  NANDN U25494 ( .A(n24944), .B(n24943), .Z(n24948) );
  NANDN U25495 ( .A(n24946), .B(n24945), .Z(n24947) );
  AND U25496 ( .A(n24948), .B(n24947), .Z(n25254) );
  XNOR U25497 ( .A(n25255), .B(n25254), .Z(n25256) );
  XOR U25498 ( .A(n25257), .B(n25256), .Z(n24979) );
  NANDN U25499 ( .A(n24950), .B(n24949), .Z(n24954) );
  OR U25500 ( .A(n24952), .B(n24951), .Z(n24953) );
  NAND U25501 ( .A(n24954), .B(n24953), .Z(n24978) );
  XNOR U25502 ( .A(n24979), .B(n24978), .Z(n24980) );
  NANDN U25503 ( .A(n24956), .B(n24955), .Z(n24960) );
  NANDN U25504 ( .A(n24958), .B(n24957), .Z(n24959) );
  NAND U25505 ( .A(n24960), .B(n24959), .Z(n24981) );
  XNOR U25506 ( .A(n24980), .B(n24981), .Z(n24972) );
  NANDN U25507 ( .A(n24962), .B(n24961), .Z(n24966) );
  OR U25508 ( .A(n24964), .B(n24963), .Z(n24965) );
  NAND U25509 ( .A(n24966), .B(n24965), .Z(n24973) );
  XNOR U25510 ( .A(n24972), .B(n24973), .Z(n24974) );
  XNOR U25511 ( .A(n24975), .B(n24974), .Z(n25260) );
  XNOR U25512 ( .A(sreg[180]), .B(n25260), .Z(n25262) );
  NANDN U25513 ( .A(sreg[179]), .B(n24967), .Z(n24971) );
  NAND U25514 ( .A(n24969), .B(n24968), .Z(n24970) );
  NAND U25515 ( .A(n24971), .B(n24970), .Z(n25261) );
  XNOR U25516 ( .A(n25262), .B(n25261), .Z(c[180]) );
  NANDN U25517 ( .A(n24973), .B(n24972), .Z(n24977) );
  NANDN U25518 ( .A(n24975), .B(n24974), .Z(n24976) );
  AND U25519 ( .A(n24977), .B(n24976), .Z(n25268) );
  NANDN U25520 ( .A(n24979), .B(n24978), .Z(n24983) );
  NANDN U25521 ( .A(n24981), .B(n24980), .Z(n24982) );
  AND U25522 ( .A(n24983), .B(n24982), .Z(n25266) );
  NANDN U25523 ( .A(n24985), .B(n24984), .Z(n24989) );
  NANDN U25524 ( .A(n24987), .B(n24986), .Z(n24988) );
  AND U25525 ( .A(n24989), .B(n24988), .Z(n25546) );
  NANDN U25526 ( .A(n24991), .B(n24990), .Z(n24995) );
  OR U25527 ( .A(n24993), .B(n24992), .Z(n24994) );
  AND U25528 ( .A(n24995), .B(n24994), .Z(n25545) );
  XNOR U25529 ( .A(n25546), .B(n25545), .Z(n25548) );
  NANDN U25530 ( .A(n24997), .B(n24996), .Z(n25001) );
  OR U25531 ( .A(n24999), .B(n24998), .Z(n25000) );
  AND U25532 ( .A(n25001), .B(n25000), .Z(n25535) );
  NANDN U25533 ( .A(n25003), .B(n25002), .Z(n25007) );
  NAND U25534 ( .A(n25005), .B(n25004), .Z(n25006) );
  AND U25535 ( .A(n25007), .B(n25006), .Z(n25534) );
  NANDN U25536 ( .A(n25009), .B(n25008), .Z(n25013) );
  NANDN U25537 ( .A(n25011), .B(n25010), .Z(n25012) );
  AND U25538 ( .A(n25013), .B(n25012), .Z(n25533) );
  XOR U25539 ( .A(n25534), .B(n25533), .Z(n25536) );
  XOR U25540 ( .A(n25535), .B(n25536), .Z(n25540) );
  NANDN U25541 ( .A(n25015), .B(n25014), .Z(n25019) );
  NANDN U25542 ( .A(n25017), .B(n25016), .Z(n25018) );
  NAND U25543 ( .A(n25019), .B(n25018), .Z(n25539) );
  XNOR U25544 ( .A(n25540), .B(n25539), .Z(n25541) );
  NANDN U25545 ( .A(n25021), .B(n25020), .Z(n25025) );
  NANDN U25546 ( .A(n25023), .B(n25022), .Z(n25024) );
  AND U25547 ( .A(n25025), .B(n25024), .Z(n25530) );
  NANDN U25548 ( .A(n25027), .B(n25026), .Z(n25031) );
  NAND U25549 ( .A(n25029), .B(n25028), .Z(n25030) );
  AND U25550 ( .A(n25031), .B(n25030), .Z(n25505) );
  NANDN U25551 ( .A(n25033), .B(n25032), .Z(n25037) );
  NANDN U25552 ( .A(n25035), .B(n25034), .Z(n25036) );
  AND U25553 ( .A(n25037), .B(n25036), .Z(n25523) );
  NANDN U25554 ( .A(n25039), .B(n25038), .Z(n25043) );
  NANDN U25555 ( .A(n25041), .B(n25040), .Z(n25042) );
  AND U25556 ( .A(n25043), .B(n25042), .Z(n25522) );
  NANDN U25557 ( .A(n33875), .B(n25044), .Z(n25046) );
  XOR U25558 ( .A(a[93]), .B(b[25]), .Z(n25301) );
  NANDN U25559 ( .A(n33994), .B(n25301), .Z(n25045) );
  AND U25560 ( .A(n25046), .B(n25045), .Z(n25471) );
  NANDN U25561 ( .A(n32013), .B(n25047), .Z(n25049) );
  XOR U25562 ( .A(a[101]), .B(b[17]), .Z(n25304) );
  NANDN U25563 ( .A(n32292), .B(n25304), .Z(n25048) );
  AND U25564 ( .A(n25049), .B(n25048), .Z(n25470) );
  NANDN U25565 ( .A(n31536), .B(n25050), .Z(n25052) );
  XOR U25566 ( .A(a[103]), .B(b[15]), .Z(n25307) );
  NANDN U25567 ( .A(n31925), .B(n25307), .Z(n25051) );
  NAND U25568 ( .A(n25052), .B(n25051), .Z(n25469) );
  XOR U25569 ( .A(n25470), .B(n25469), .Z(n25472) );
  XOR U25570 ( .A(n25471), .B(n25472), .Z(n25443) );
  NANDN U25571 ( .A(n37526), .B(n25053), .Z(n25055) );
  XOR U25572 ( .A(b[51]), .B(a[67]), .Z(n25310) );
  NANDN U25573 ( .A(n37605), .B(n25310), .Z(n25054) );
  AND U25574 ( .A(n25055), .B(n25054), .Z(n25495) );
  NANDN U25575 ( .A(n37705), .B(n25056), .Z(n25058) );
  XOR U25576 ( .A(b[53]), .B(a[65]), .Z(n25313) );
  NANDN U25577 ( .A(n37778), .B(n25313), .Z(n25057) );
  AND U25578 ( .A(n25058), .B(n25057), .Z(n25494) );
  NANDN U25579 ( .A(n36210), .B(n25059), .Z(n25061) );
  XOR U25580 ( .A(b[39]), .B(a[79]), .Z(n25316) );
  NANDN U25581 ( .A(n36347), .B(n25316), .Z(n25060) );
  NAND U25582 ( .A(n25061), .B(n25060), .Z(n25493) );
  XOR U25583 ( .A(n25494), .B(n25493), .Z(n25496) );
  XNOR U25584 ( .A(n25495), .B(n25496), .Z(n25442) );
  XNOR U25585 ( .A(n25443), .B(n25442), .Z(n25445) );
  NANDN U25586 ( .A(n25063), .B(n25062), .Z(n25067) );
  OR U25587 ( .A(n25065), .B(n25064), .Z(n25066) );
  AND U25588 ( .A(n25067), .B(n25066), .Z(n25444) );
  XOR U25589 ( .A(n25445), .B(n25444), .Z(n25292) );
  NANDN U25590 ( .A(n25069), .B(n25068), .Z(n25073) );
  OR U25591 ( .A(n25071), .B(n25070), .Z(n25072) );
  AND U25592 ( .A(n25073), .B(n25072), .Z(n25290) );
  NANDN U25593 ( .A(n25075), .B(n25074), .Z(n25079) );
  NANDN U25594 ( .A(n25077), .B(n25076), .Z(n25078) );
  NAND U25595 ( .A(n25079), .B(n25078), .Z(n25289) );
  XNOR U25596 ( .A(n25290), .B(n25289), .Z(n25291) );
  XNOR U25597 ( .A(n25292), .B(n25291), .Z(n25521) );
  XOR U25598 ( .A(n25522), .B(n25521), .Z(n25524) );
  XOR U25599 ( .A(n25523), .B(n25524), .Z(n25504) );
  NANDN U25600 ( .A(n25081), .B(n25080), .Z(n25085) );
  NANDN U25601 ( .A(n25083), .B(n25082), .Z(n25084) );
  AND U25602 ( .A(n25085), .B(n25084), .Z(n25516) );
  NANDN U25603 ( .A(n25086), .B(n37294), .Z(n25088) );
  XOR U25604 ( .A(b[47]), .B(a[71]), .Z(n25343) );
  NANDN U25605 ( .A(n37172), .B(n25343), .Z(n25087) );
  AND U25606 ( .A(n25088), .B(n25087), .Z(n25384) );
  NANDN U25607 ( .A(n25089), .B(n30627), .Z(n25091) );
  XOR U25608 ( .A(a[109]), .B(b[9]), .Z(n25346) );
  NANDN U25609 ( .A(n30267), .B(n25346), .Z(n25090) );
  AND U25610 ( .A(n25091), .B(n25090), .Z(n25383) );
  NANDN U25611 ( .A(n25092), .B(n37536), .Z(n25094) );
  XOR U25612 ( .A(b[49]), .B(a[69]), .Z(n25349) );
  NANDN U25613 ( .A(n37432), .B(n25349), .Z(n25093) );
  NAND U25614 ( .A(n25094), .B(n25093), .Z(n25382) );
  XOR U25615 ( .A(n25383), .B(n25382), .Z(n25385) );
  XOR U25616 ( .A(n25384), .B(n25385), .Z(n25449) );
  NANDN U25617 ( .A(n36742), .B(n25095), .Z(n25097) );
  XOR U25618 ( .A(b[43]), .B(a[75]), .Z(n25352) );
  NANDN U25619 ( .A(n36891), .B(n25352), .Z(n25096) );
  AND U25620 ( .A(n25097), .B(n25096), .Z(n25363) );
  NANDN U25621 ( .A(n36991), .B(n25098), .Z(n25100) );
  XOR U25622 ( .A(b[45]), .B(a[73]), .Z(n25355) );
  NANDN U25623 ( .A(n37083), .B(n25355), .Z(n25099) );
  AND U25624 ( .A(n25100), .B(n25099), .Z(n25362) );
  NANDN U25625 ( .A(n30482), .B(n25101), .Z(n25103) );
  XOR U25626 ( .A(a[107]), .B(b[11]), .Z(n25358) );
  NANDN U25627 ( .A(n30891), .B(n25358), .Z(n25102) );
  NAND U25628 ( .A(n25103), .B(n25102), .Z(n25361) );
  XOR U25629 ( .A(n25362), .B(n25361), .Z(n25364) );
  XNOR U25630 ( .A(n25363), .B(n25364), .Z(n25448) );
  XNOR U25631 ( .A(n25449), .B(n25448), .Z(n25450) );
  NANDN U25632 ( .A(n25105), .B(n25104), .Z(n25109) );
  OR U25633 ( .A(n25107), .B(n25106), .Z(n25108) );
  NAND U25634 ( .A(n25109), .B(n25108), .Z(n25451) );
  XNOR U25635 ( .A(n25450), .B(n25451), .Z(n25515) );
  XNOR U25636 ( .A(n25516), .B(n25515), .Z(n25517) );
  NANDN U25637 ( .A(n29499), .B(n25110), .Z(n25112) );
  XOR U25638 ( .A(a[111]), .B(b[7]), .Z(n25367) );
  NANDN U25639 ( .A(n29735), .B(n25367), .Z(n25111) );
  AND U25640 ( .A(n25112), .B(n25111), .Z(n25327) );
  NANDN U25641 ( .A(n37857), .B(n25113), .Z(n25115) );
  XOR U25642 ( .A(b[55]), .B(a[63]), .Z(n25370) );
  NANDN U25643 ( .A(n37911), .B(n25370), .Z(n25114) );
  AND U25644 ( .A(n25115), .B(n25114), .Z(n25326) );
  NANDN U25645 ( .A(n35611), .B(n25116), .Z(n25118) );
  XOR U25646 ( .A(b[35]), .B(a[83]), .Z(n25373) );
  NANDN U25647 ( .A(n35801), .B(n25373), .Z(n25117) );
  NAND U25648 ( .A(n25118), .B(n25117), .Z(n25325) );
  XOR U25649 ( .A(n25326), .B(n25325), .Z(n25328) );
  XOR U25650 ( .A(n25327), .B(n25328), .Z(n25401) );
  NANDN U25651 ( .A(n25120), .B(n25119), .Z(n25124) );
  OR U25652 ( .A(n25122), .B(n25121), .Z(n25123) );
  AND U25653 ( .A(n25124), .B(n25123), .Z(n25400) );
  XNOR U25654 ( .A(n25401), .B(n25400), .Z(n25402) );
  NAND U25655 ( .A(n25126), .B(n25125), .Z(n25130) );
  NANDN U25656 ( .A(n25128), .B(n25127), .Z(n25129) );
  NAND U25657 ( .A(n25130), .B(n25129), .Z(n25403) );
  XOR U25658 ( .A(n25402), .B(n25403), .Z(n25518) );
  XNOR U25659 ( .A(n25517), .B(n25518), .Z(n25503) );
  XOR U25660 ( .A(n25504), .B(n25503), .Z(n25506) );
  XOR U25661 ( .A(n25505), .B(n25506), .Z(n25528) );
  NANDN U25662 ( .A(n25132), .B(n25131), .Z(n25136) );
  NANDN U25663 ( .A(n25134), .B(n25133), .Z(n25135) );
  AND U25664 ( .A(n25136), .B(n25135), .Z(n25511) );
  NANDN U25665 ( .A(n25138), .B(n25137), .Z(n25142) );
  NANDN U25666 ( .A(n25140), .B(n25139), .Z(n25141) );
  AND U25667 ( .A(n25142), .B(n25141), .Z(n25510) );
  NANDN U25668 ( .A(n25144), .B(n25143), .Z(n25148) );
  NAND U25669 ( .A(n25146), .B(n25145), .Z(n25147) );
  AND U25670 ( .A(n25148), .B(n25147), .Z(n25509) );
  XOR U25671 ( .A(n25510), .B(n25509), .Z(n25512) );
  XOR U25672 ( .A(n25511), .B(n25512), .Z(n25280) );
  NANDN U25673 ( .A(n25150), .B(n25149), .Z(n25154) );
  NANDN U25674 ( .A(n25152), .B(n25151), .Z(n25153) );
  AND U25675 ( .A(n25154), .B(n25153), .Z(n25395) );
  NANDN U25676 ( .A(n25156), .B(n25155), .Z(n25160) );
  OR U25677 ( .A(n25158), .B(n25157), .Z(n25159) );
  NAND U25678 ( .A(n25160), .B(n25159), .Z(n25394) );
  XNOR U25679 ( .A(n25395), .B(n25394), .Z(n25397) );
  NANDN U25680 ( .A(n25162), .B(n25161), .Z(n25166) );
  OR U25681 ( .A(n25164), .B(n25163), .Z(n25165) );
  NAND U25682 ( .A(n25166), .B(n25165), .Z(n25297) );
  NAND U25683 ( .A(b[0]), .B(a[117]), .Z(n25167) );
  XNOR U25684 ( .A(b[1]), .B(n25167), .Z(n25169) );
  NANDN U25685 ( .A(b[0]), .B(a[116]), .Z(n25168) );
  NAND U25686 ( .A(n25169), .B(n25168), .Z(n25334) );
  NANDN U25687 ( .A(n38278), .B(n25170), .Z(n25172) );
  XOR U25688 ( .A(b[63]), .B(a[55]), .Z(n25427) );
  NANDN U25689 ( .A(n38279), .B(n25427), .Z(n25171) );
  AND U25690 ( .A(n25172), .B(n25171), .Z(n25332) );
  NANDN U25691 ( .A(n35260), .B(n25173), .Z(n25175) );
  XOR U25692 ( .A(b[33]), .B(a[85]), .Z(n25430) );
  NANDN U25693 ( .A(n35456), .B(n25430), .Z(n25174) );
  NAND U25694 ( .A(n25175), .B(n25174), .Z(n25331) );
  XNOR U25695 ( .A(n25332), .B(n25331), .Z(n25333) );
  XNOR U25696 ( .A(n25334), .B(n25333), .Z(n25296) );
  NANDN U25697 ( .A(n37974), .B(n25176), .Z(n25178) );
  XOR U25698 ( .A(b[57]), .B(a[61]), .Z(n25433) );
  NANDN U25699 ( .A(n38031), .B(n25433), .Z(n25177) );
  AND U25700 ( .A(n25178), .B(n25177), .Z(n25408) );
  NANDN U25701 ( .A(n38090), .B(n25179), .Z(n25181) );
  XOR U25702 ( .A(b[59]), .B(a[59]), .Z(n25436) );
  NANDN U25703 ( .A(n38130), .B(n25436), .Z(n25180) );
  AND U25704 ( .A(n25181), .B(n25180), .Z(n25407) );
  NANDN U25705 ( .A(n36480), .B(n25182), .Z(n25184) );
  XOR U25706 ( .A(b[41]), .B(a[77]), .Z(n25439) );
  NANDN U25707 ( .A(n36594), .B(n25439), .Z(n25183) );
  NAND U25708 ( .A(n25184), .B(n25183), .Z(n25406) );
  XOR U25709 ( .A(n25407), .B(n25406), .Z(n25409) );
  XOR U25710 ( .A(n25408), .B(n25409), .Z(n25295) );
  XOR U25711 ( .A(n25296), .B(n25295), .Z(n25298) );
  XOR U25712 ( .A(n25297), .B(n25298), .Z(n25396) );
  XOR U25713 ( .A(n25397), .B(n25396), .Z(n25284) );
  NANDN U25714 ( .A(n25186), .B(n25185), .Z(n25190) );
  NAND U25715 ( .A(n25188), .B(n25187), .Z(n25189) );
  NAND U25716 ( .A(n25190), .B(n25189), .Z(n25283) );
  XNOR U25717 ( .A(n25284), .B(n25283), .Z(n25286) );
  NAND U25718 ( .A(n25192), .B(n25191), .Z(n25196) );
  NANDN U25719 ( .A(n25194), .B(n25193), .Z(n25195) );
  AND U25720 ( .A(n25196), .B(n25195), .Z(n25502) );
  NANDN U25721 ( .A(n25198), .B(n25197), .Z(n25202) );
  OR U25722 ( .A(n25200), .B(n25199), .Z(n25201) );
  AND U25723 ( .A(n25202), .B(n25201), .Z(n25390) );
  NANDN U25724 ( .A(n34223), .B(n25203), .Z(n25205) );
  XOR U25725 ( .A(b[27]), .B(a[91]), .Z(n25475) );
  NANDN U25726 ( .A(n34458), .B(n25475), .Z(n25204) );
  AND U25727 ( .A(n25205), .B(n25204), .Z(n25322) );
  NANDN U25728 ( .A(n34634), .B(n25206), .Z(n25208) );
  XOR U25729 ( .A(b[29]), .B(a[89]), .Z(n25478) );
  NANDN U25730 ( .A(n34722), .B(n25478), .Z(n25207) );
  AND U25731 ( .A(n25208), .B(n25207), .Z(n25320) );
  NANDN U25732 ( .A(n31055), .B(n25209), .Z(n25211) );
  XOR U25733 ( .A(a[105]), .B(b[13]), .Z(n25481) );
  NANDN U25734 ( .A(n31293), .B(n25481), .Z(n25210) );
  NAND U25735 ( .A(n25211), .B(n25210), .Z(n25319) );
  XNOR U25736 ( .A(n25320), .B(n25319), .Z(n25321) );
  XOR U25737 ( .A(n25322), .B(n25321), .Z(n25389) );
  NANDN U25738 ( .A(n28889), .B(n25212), .Z(n25214) );
  XOR U25739 ( .A(a[113]), .B(b[5]), .Z(n25484) );
  NANDN U25740 ( .A(n29138), .B(n25484), .Z(n25213) );
  AND U25741 ( .A(n25214), .B(n25213), .Z(n25415) );
  NANDN U25742 ( .A(n209), .B(n25215), .Z(n25217) );
  XOR U25743 ( .A(a[115]), .B(b[3]), .Z(n25487) );
  NANDN U25744 ( .A(n28941), .B(n25487), .Z(n25216) );
  AND U25745 ( .A(n25217), .B(n25216), .Z(n25413) );
  NANDN U25746 ( .A(n35936), .B(n25218), .Z(n25220) );
  XOR U25747 ( .A(b[37]), .B(a[81]), .Z(n25490) );
  NANDN U25748 ( .A(n36047), .B(n25490), .Z(n25219) );
  NAND U25749 ( .A(n25220), .B(n25219), .Z(n25412) );
  XNOR U25750 ( .A(n25413), .B(n25412), .Z(n25414) );
  XOR U25751 ( .A(n25415), .B(n25414), .Z(n25388) );
  XNOR U25752 ( .A(n25389), .B(n25388), .Z(n25391) );
  NANDN U25753 ( .A(n25222), .B(n25221), .Z(n25226) );
  OR U25754 ( .A(n25224), .B(n25223), .Z(n25225) );
  AND U25755 ( .A(n25226), .B(n25225), .Z(n25339) );
  NANDN U25756 ( .A(n32996), .B(n25227), .Z(n25229) );
  XOR U25757 ( .A(a[97]), .B(b[21]), .Z(n25454) );
  NANDN U25758 ( .A(n33271), .B(n25454), .Z(n25228) );
  AND U25759 ( .A(n25229), .B(n25228), .Z(n25421) );
  NANDN U25760 ( .A(n33866), .B(n25230), .Z(n25232) );
  XOR U25761 ( .A(a[95]), .B(b[23]), .Z(n25457) );
  NANDN U25762 ( .A(n33644), .B(n25457), .Z(n25231) );
  AND U25763 ( .A(n25232), .B(n25231), .Z(n25419) );
  NANDN U25764 ( .A(n32483), .B(n25233), .Z(n25235) );
  XOR U25765 ( .A(a[99]), .B(b[19]), .Z(n25460) );
  NANDN U25766 ( .A(n32823), .B(n25460), .Z(n25234) );
  NAND U25767 ( .A(n25235), .B(n25234), .Z(n25418) );
  XNOR U25768 ( .A(n25419), .B(n25418), .Z(n25420) );
  XOR U25769 ( .A(n25421), .B(n25420), .Z(n25338) );
  NANDN U25770 ( .A(n34909), .B(n25236), .Z(n25238) );
  XOR U25771 ( .A(b[31]), .B(a[87]), .Z(n25463) );
  NANDN U25772 ( .A(n35145), .B(n25463), .Z(n25237) );
  AND U25773 ( .A(n25238), .B(n25237), .Z(n25379) );
  NANDN U25774 ( .A(n38247), .B(n25239), .Z(n25241) );
  XOR U25775 ( .A(b[61]), .B(a[57]), .Z(n25466) );
  NANDN U25776 ( .A(n38248), .B(n25466), .Z(n25240) );
  AND U25777 ( .A(n25241), .B(n25240), .Z(n25377) );
  AND U25778 ( .A(b[63]), .B(a[53]), .Z(n25376) );
  XNOR U25779 ( .A(n25377), .B(n25376), .Z(n25378) );
  XOR U25780 ( .A(n25379), .B(n25378), .Z(n25337) );
  XNOR U25781 ( .A(n25338), .B(n25337), .Z(n25340) );
  XOR U25782 ( .A(n25500), .B(n25499), .Z(n25501) );
  XNOR U25783 ( .A(n25502), .B(n25501), .Z(n25285) );
  XOR U25784 ( .A(n25286), .B(n25285), .Z(n25278) );
  NANDN U25785 ( .A(n25243), .B(n25242), .Z(n25247) );
  NANDN U25786 ( .A(n25245), .B(n25244), .Z(n25246) );
  AND U25787 ( .A(n25247), .B(n25246), .Z(n25277) );
  XNOR U25788 ( .A(n25278), .B(n25277), .Z(n25279) );
  XNOR U25789 ( .A(n25280), .B(n25279), .Z(n25527) );
  XNOR U25790 ( .A(n25528), .B(n25527), .Z(n25529) );
  XOR U25791 ( .A(n25530), .B(n25529), .Z(n25542) );
  XNOR U25792 ( .A(n25541), .B(n25542), .Z(n25547) );
  XOR U25793 ( .A(n25548), .B(n25547), .Z(n25272) );
  NANDN U25794 ( .A(n25249), .B(n25248), .Z(n25253) );
  NANDN U25795 ( .A(n25251), .B(n25250), .Z(n25252) );
  AND U25796 ( .A(n25253), .B(n25252), .Z(n25271) );
  XNOR U25797 ( .A(n25272), .B(n25271), .Z(n25273) );
  NANDN U25798 ( .A(n25255), .B(n25254), .Z(n25259) );
  NAND U25799 ( .A(n25257), .B(n25256), .Z(n25258) );
  NAND U25800 ( .A(n25259), .B(n25258), .Z(n25274) );
  XNOR U25801 ( .A(n25273), .B(n25274), .Z(n25265) );
  XNOR U25802 ( .A(n25266), .B(n25265), .Z(n25267) );
  XNOR U25803 ( .A(n25268), .B(n25267), .Z(n25551) );
  XNOR U25804 ( .A(sreg[181]), .B(n25551), .Z(n25553) );
  NANDN U25805 ( .A(sreg[180]), .B(n25260), .Z(n25264) );
  NAND U25806 ( .A(n25262), .B(n25261), .Z(n25263) );
  NAND U25807 ( .A(n25264), .B(n25263), .Z(n25552) );
  XNOR U25808 ( .A(n25553), .B(n25552), .Z(c[181]) );
  NANDN U25809 ( .A(n25266), .B(n25265), .Z(n25270) );
  NANDN U25810 ( .A(n25268), .B(n25267), .Z(n25269) );
  AND U25811 ( .A(n25270), .B(n25269), .Z(n25559) );
  NANDN U25812 ( .A(n25272), .B(n25271), .Z(n25276) );
  NANDN U25813 ( .A(n25274), .B(n25273), .Z(n25275) );
  AND U25814 ( .A(n25276), .B(n25275), .Z(n25557) );
  NANDN U25815 ( .A(n25278), .B(n25277), .Z(n25282) );
  NANDN U25816 ( .A(n25280), .B(n25279), .Z(n25281) );
  AND U25817 ( .A(n25282), .B(n25281), .Z(n25576) );
  NANDN U25818 ( .A(n25284), .B(n25283), .Z(n25288) );
  NAND U25819 ( .A(n25286), .B(n25285), .Z(n25287) );
  AND U25820 ( .A(n25288), .B(n25287), .Z(n25588) );
  NANDN U25821 ( .A(n25290), .B(n25289), .Z(n25294) );
  NANDN U25822 ( .A(n25292), .B(n25291), .Z(n25293) );
  AND U25823 ( .A(n25294), .B(n25293), .Z(n25600) );
  NAND U25824 ( .A(n25296), .B(n25295), .Z(n25300) );
  NAND U25825 ( .A(n25298), .B(n25297), .Z(n25299) );
  AND U25826 ( .A(n25300), .B(n25299), .Z(n25599) );
  NANDN U25827 ( .A(n33875), .B(n25301), .Z(n25303) );
  XOR U25828 ( .A(a[94]), .B(b[25]), .Z(n25679) );
  NANDN U25829 ( .A(n33994), .B(n25679), .Z(n25302) );
  AND U25830 ( .A(n25303), .B(n25302), .Z(n25804) );
  NANDN U25831 ( .A(n32013), .B(n25304), .Z(n25306) );
  XOR U25832 ( .A(a[102]), .B(b[17]), .Z(n25682) );
  NANDN U25833 ( .A(n32292), .B(n25682), .Z(n25305) );
  AND U25834 ( .A(n25306), .B(n25305), .Z(n25803) );
  NANDN U25835 ( .A(n31536), .B(n25307), .Z(n25309) );
  XOR U25836 ( .A(a[104]), .B(b[15]), .Z(n25685) );
  NANDN U25837 ( .A(n31925), .B(n25685), .Z(n25308) );
  NAND U25838 ( .A(n25309), .B(n25308), .Z(n25802) );
  XOR U25839 ( .A(n25803), .B(n25802), .Z(n25805) );
  XOR U25840 ( .A(n25804), .B(n25805), .Z(n25776) );
  NANDN U25841 ( .A(n37526), .B(n25310), .Z(n25312) );
  XOR U25842 ( .A(b[51]), .B(a[68]), .Z(n25688) );
  NANDN U25843 ( .A(n37605), .B(n25688), .Z(n25311) );
  AND U25844 ( .A(n25312), .B(n25311), .Z(n25828) );
  NANDN U25845 ( .A(n37705), .B(n25313), .Z(n25315) );
  XOR U25846 ( .A(b[53]), .B(a[66]), .Z(n25691) );
  NANDN U25847 ( .A(n37778), .B(n25691), .Z(n25314) );
  AND U25848 ( .A(n25315), .B(n25314), .Z(n25827) );
  NANDN U25849 ( .A(n36210), .B(n25316), .Z(n25318) );
  XOR U25850 ( .A(b[39]), .B(a[80]), .Z(n25694) );
  NANDN U25851 ( .A(n36347), .B(n25694), .Z(n25317) );
  NAND U25852 ( .A(n25318), .B(n25317), .Z(n25826) );
  XOR U25853 ( .A(n25827), .B(n25826), .Z(n25829) );
  XNOR U25854 ( .A(n25828), .B(n25829), .Z(n25775) );
  XNOR U25855 ( .A(n25776), .B(n25775), .Z(n25778) );
  NANDN U25856 ( .A(n25320), .B(n25319), .Z(n25324) );
  NANDN U25857 ( .A(n25322), .B(n25321), .Z(n25323) );
  AND U25858 ( .A(n25324), .B(n25323), .Z(n25777) );
  XOR U25859 ( .A(n25778), .B(n25777), .Z(n25670) );
  NANDN U25860 ( .A(n25326), .B(n25325), .Z(n25330) );
  OR U25861 ( .A(n25328), .B(n25327), .Z(n25329) );
  AND U25862 ( .A(n25330), .B(n25329), .Z(n25668) );
  NANDN U25863 ( .A(n25332), .B(n25331), .Z(n25336) );
  NANDN U25864 ( .A(n25334), .B(n25333), .Z(n25335) );
  NAND U25865 ( .A(n25336), .B(n25335), .Z(n25667) );
  XNOR U25866 ( .A(n25668), .B(n25667), .Z(n25669) );
  XNOR U25867 ( .A(n25670), .B(n25669), .Z(n25598) );
  XOR U25868 ( .A(n25599), .B(n25598), .Z(n25601) );
  XOR U25869 ( .A(n25600), .B(n25601), .Z(n25587) );
  NAND U25870 ( .A(n25338), .B(n25337), .Z(n25342) );
  NANDN U25871 ( .A(n25340), .B(n25339), .Z(n25341) );
  AND U25872 ( .A(n25342), .B(n25341), .Z(n25605) );
  NANDN U25873 ( .A(n211), .B(n25343), .Z(n25345) );
  XOR U25874 ( .A(b[47]), .B(a[72]), .Z(n25643) );
  NANDN U25875 ( .A(n37172), .B(n25643), .Z(n25344) );
  AND U25876 ( .A(n25345), .B(n25344), .Z(n25633) );
  NANDN U25877 ( .A(n210), .B(n25346), .Z(n25348) );
  XOR U25878 ( .A(a[110]), .B(b[9]), .Z(n25646) );
  NANDN U25879 ( .A(n30267), .B(n25646), .Z(n25347) );
  AND U25880 ( .A(n25348), .B(n25347), .Z(n25632) );
  NANDN U25881 ( .A(n212), .B(n25349), .Z(n25351) );
  XOR U25882 ( .A(b[49]), .B(a[70]), .Z(n25649) );
  NANDN U25883 ( .A(n37432), .B(n25649), .Z(n25350) );
  NAND U25884 ( .A(n25351), .B(n25350), .Z(n25631) );
  XOR U25885 ( .A(n25632), .B(n25631), .Z(n25634) );
  XOR U25886 ( .A(n25633), .B(n25634), .Z(n25782) );
  NANDN U25887 ( .A(n36742), .B(n25352), .Z(n25354) );
  XOR U25888 ( .A(b[43]), .B(a[76]), .Z(n25652) );
  NANDN U25889 ( .A(n36891), .B(n25652), .Z(n25353) );
  AND U25890 ( .A(n25354), .B(n25353), .Z(n25663) );
  NANDN U25891 ( .A(n36991), .B(n25355), .Z(n25357) );
  XOR U25892 ( .A(b[45]), .B(a[74]), .Z(n25655) );
  NANDN U25893 ( .A(n37083), .B(n25655), .Z(n25356) );
  AND U25894 ( .A(n25357), .B(n25356), .Z(n25662) );
  NANDN U25895 ( .A(n30482), .B(n25358), .Z(n25360) );
  XOR U25896 ( .A(a[108]), .B(b[11]), .Z(n25658) );
  NANDN U25897 ( .A(n30891), .B(n25658), .Z(n25359) );
  NAND U25898 ( .A(n25360), .B(n25359), .Z(n25661) );
  XOR U25899 ( .A(n25662), .B(n25661), .Z(n25664) );
  XNOR U25900 ( .A(n25663), .B(n25664), .Z(n25781) );
  XNOR U25901 ( .A(n25782), .B(n25781), .Z(n25783) );
  NANDN U25902 ( .A(n25362), .B(n25361), .Z(n25366) );
  OR U25903 ( .A(n25364), .B(n25363), .Z(n25365) );
  NAND U25904 ( .A(n25366), .B(n25365), .Z(n25784) );
  XNOR U25905 ( .A(n25783), .B(n25784), .Z(n25604) );
  XNOR U25906 ( .A(n25605), .B(n25604), .Z(n25606) );
  NANDN U25907 ( .A(n29499), .B(n25367), .Z(n25369) );
  XOR U25908 ( .A(a[112]), .B(b[7]), .Z(n25616) );
  NANDN U25909 ( .A(n29735), .B(n25616), .Z(n25368) );
  AND U25910 ( .A(n25369), .B(n25368), .Z(n25705) );
  NANDN U25911 ( .A(n37857), .B(n25370), .Z(n25372) );
  XOR U25912 ( .A(b[55]), .B(a[64]), .Z(n25619) );
  NANDN U25913 ( .A(n37911), .B(n25619), .Z(n25371) );
  AND U25914 ( .A(n25372), .B(n25371), .Z(n25704) );
  NANDN U25915 ( .A(n35611), .B(n25373), .Z(n25375) );
  XOR U25916 ( .A(b[35]), .B(a[84]), .Z(n25622) );
  NANDN U25917 ( .A(n35801), .B(n25622), .Z(n25374) );
  NAND U25918 ( .A(n25375), .B(n25374), .Z(n25703) );
  XOR U25919 ( .A(n25704), .B(n25703), .Z(n25706) );
  XOR U25920 ( .A(n25705), .B(n25706), .Z(n25722) );
  NANDN U25921 ( .A(n25377), .B(n25376), .Z(n25381) );
  NANDN U25922 ( .A(n25379), .B(n25378), .Z(n25380) );
  AND U25923 ( .A(n25381), .B(n25380), .Z(n25721) );
  XNOR U25924 ( .A(n25722), .B(n25721), .Z(n25723) );
  NANDN U25925 ( .A(n25383), .B(n25382), .Z(n25387) );
  OR U25926 ( .A(n25385), .B(n25384), .Z(n25386) );
  NAND U25927 ( .A(n25387), .B(n25386), .Z(n25724) );
  XOR U25928 ( .A(n25723), .B(n25724), .Z(n25607) );
  XNOR U25929 ( .A(n25606), .B(n25607), .Z(n25586) );
  XOR U25930 ( .A(n25587), .B(n25586), .Z(n25589) );
  XOR U25931 ( .A(n25588), .B(n25589), .Z(n25575) );
  NAND U25932 ( .A(n25389), .B(n25388), .Z(n25393) );
  NANDN U25933 ( .A(n25391), .B(n25390), .Z(n25392) );
  NAND U25934 ( .A(n25393), .B(n25392), .Z(n25592) );
  NANDN U25935 ( .A(n25395), .B(n25394), .Z(n25399) );
  NAND U25936 ( .A(n25397), .B(n25396), .Z(n25398) );
  AND U25937 ( .A(n25399), .B(n25398), .Z(n25593) );
  XOR U25938 ( .A(n25592), .B(n25593), .Z(n25595) );
  NANDN U25939 ( .A(n25401), .B(n25400), .Z(n25405) );
  NANDN U25940 ( .A(n25403), .B(n25402), .Z(n25404) );
  NAND U25941 ( .A(n25405), .B(n25404), .Z(n25594) );
  XOR U25942 ( .A(n25595), .B(n25594), .Z(n25613) );
  NANDN U25943 ( .A(n25407), .B(n25406), .Z(n25411) );
  OR U25944 ( .A(n25409), .B(n25408), .Z(n25410) );
  AND U25945 ( .A(n25411), .B(n25410), .Z(n25734) );
  NANDN U25946 ( .A(n25413), .B(n25412), .Z(n25417) );
  NANDN U25947 ( .A(n25415), .B(n25414), .Z(n25416) );
  NAND U25948 ( .A(n25417), .B(n25416), .Z(n25733) );
  XNOR U25949 ( .A(n25734), .B(n25733), .Z(n25736) );
  NANDN U25950 ( .A(n25419), .B(n25418), .Z(n25423) );
  NANDN U25951 ( .A(n25421), .B(n25420), .Z(n25422) );
  AND U25952 ( .A(n25423), .B(n25422), .Z(n25676) );
  NAND U25953 ( .A(b[0]), .B(a[118]), .Z(n25424) );
  XNOR U25954 ( .A(b[1]), .B(n25424), .Z(n25426) );
  NANDN U25955 ( .A(b[0]), .B(a[117]), .Z(n25425) );
  NAND U25956 ( .A(n25426), .B(n25425), .Z(n25712) );
  NANDN U25957 ( .A(n38278), .B(n25427), .Z(n25429) );
  XOR U25958 ( .A(b[63]), .B(a[56]), .Z(n25757) );
  NANDN U25959 ( .A(n38279), .B(n25757), .Z(n25428) );
  AND U25960 ( .A(n25429), .B(n25428), .Z(n25710) );
  NANDN U25961 ( .A(n35260), .B(n25430), .Z(n25432) );
  XOR U25962 ( .A(b[33]), .B(a[86]), .Z(n25760) );
  NANDN U25963 ( .A(n35456), .B(n25760), .Z(n25431) );
  NAND U25964 ( .A(n25432), .B(n25431), .Z(n25709) );
  XNOR U25965 ( .A(n25710), .B(n25709), .Z(n25711) );
  XNOR U25966 ( .A(n25712), .B(n25711), .Z(n25673) );
  NANDN U25967 ( .A(n37974), .B(n25433), .Z(n25435) );
  XOR U25968 ( .A(b[57]), .B(a[62]), .Z(n25766) );
  NANDN U25969 ( .A(n38031), .B(n25766), .Z(n25434) );
  AND U25970 ( .A(n25435), .B(n25434), .Z(n25742) );
  NANDN U25971 ( .A(n38090), .B(n25436), .Z(n25438) );
  XOR U25972 ( .A(b[59]), .B(a[60]), .Z(n25769) );
  NANDN U25973 ( .A(n38130), .B(n25769), .Z(n25437) );
  AND U25974 ( .A(n25438), .B(n25437), .Z(n25740) );
  NANDN U25975 ( .A(n36480), .B(n25439), .Z(n25441) );
  XOR U25976 ( .A(b[41]), .B(a[78]), .Z(n25772) );
  NANDN U25977 ( .A(n36594), .B(n25772), .Z(n25440) );
  NAND U25978 ( .A(n25441), .B(n25440), .Z(n25739) );
  XNOR U25979 ( .A(n25740), .B(n25739), .Z(n25741) );
  XOR U25980 ( .A(n25742), .B(n25741), .Z(n25674) );
  XNOR U25981 ( .A(n25673), .B(n25674), .Z(n25675) );
  XNOR U25982 ( .A(n25676), .B(n25675), .Z(n25735) );
  XOR U25983 ( .A(n25736), .B(n25735), .Z(n25716) );
  NANDN U25984 ( .A(n25443), .B(n25442), .Z(n25447) );
  NAND U25985 ( .A(n25445), .B(n25444), .Z(n25446) );
  NAND U25986 ( .A(n25447), .B(n25446), .Z(n25715) );
  XNOR U25987 ( .A(n25716), .B(n25715), .Z(n25718) );
  NANDN U25988 ( .A(n25449), .B(n25448), .Z(n25453) );
  NANDN U25989 ( .A(n25451), .B(n25450), .Z(n25452) );
  AND U25990 ( .A(n25453), .B(n25452), .Z(n25835) );
  NANDN U25991 ( .A(n32996), .B(n25454), .Z(n25456) );
  XOR U25992 ( .A(a[98]), .B(b[21]), .Z(n25787) );
  NANDN U25993 ( .A(n33271), .B(n25787), .Z(n25455) );
  AND U25994 ( .A(n25456), .B(n25455), .Z(n25753) );
  NANDN U25995 ( .A(n33866), .B(n25457), .Z(n25459) );
  XOR U25996 ( .A(a[96]), .B(b[23]), .Z(n25790) );
  NANDN U25997 ( .A(n33644), .B(n25790), .Z(n25458) );
  AND U25998 ( .A(n25459), .B(n25458), .Z(n25752) );
  NANDN U25999 ( .A(n32483), .B(n25460), .Z(n25462) );
  XOR U26000 ( .A(a[100]), .B(b[19]), .Z(n25793) );
  NANDN U26001 ( .A(n32823), .B(n25793), .Z(n25461) );
  NAND U26002 ( .A(n25462), .B(n25461), .Z(n25751) );
  XOR U26003 ( .A(n25752), .B(n25751), .Z(n25754) );
  XOR U26004 ( .A(n25753), .B(n25754), .Z(n25638) );
  NANDN U26005 ( .A(n34909), .B(n25463), .Z(n25465) );
  XOR U26006 ( .A(b[31]), .B(a[88]), .Z(n25796) );
  NANDN U26007 ( .A(n35145), .B(n25796), .Z(n25464) );
  AND U26008 ( .A(n25465), .B(n25464), .Z(n25627) );
  NANDN U26009 ( .A(n38247), .B(n25466), .Z(n25468) );
  XOR U26010 ( .A(b[61]), .B(a[58]), .Z(n25799) );
  NANDN U26011 ( .A(n38248), .B(n25799), .Z(n25467) );
  AND U26012 ( .A(n25468), .B(n25467), .Z(n25626) );
  AND U26013 ( .A(b[63]), .B(a[54]), .Z(n25625) );
  XOR U26014 ( .A(n25626), .B(n25625), .Z(n25628) );
  XNOR U26015 ( .A(n25627), .B(n25628), .Z(n25637) );
  XNOR U26016 ( .A(n25638), .B(n25637), .Z(n25639) );
  NANDN U26017 ( .A(n25470), .B(n25469), .Z(n25474) );
  OR U26018 ( .A(n25472), .B(n25471), .Z(n25473) );
  NAND U26019 ( .A(n25474), .B(n25473), .Z(n25640) );
  XNOR U26020 ( .A(n25639), .B(n25640), .Z(n25832) );
  NANDN U26021 ( .A(n34223), .B(n25475), .Z(n25477) );
  XOR U26022 ( .A(b[27]), .B(a[92]), .Z(n25808) );
  NANDN U26023 ( .A(n34458), .B(n25808), .Z(n25476) );
  AND U26024 ( .A(n25477), .B(n25476), .Z(n25699) );
  NANDN U26025 ( .A(n34634), .B(n25478), .Z(n25480) );
  XOR U26026 ( .A(b[29]), .B(a[90]), .Z(n25811) );
  NANDN U26027 ( .A(n34722), .B(n25811), .Z(n25479) );
  AND U26028 ( .A(n25480), .B(n25479), .Z(n25698) );
  NANDN U26029 ( .A(n31055), .B(n25481), .Z(n25483) );
  XOR U26030 ( .A(a[106]), .B(b[13]), .Z(n25814) );
  NANDN U26031 ( .A(n31293), .B(n25814), .Z(n25482) );
  NAND U26032 ( .A(n25483), .B(n25482), .Z(n25697) );
  XOR U26033 ( .A(n25698), .B(n25697), .Z(n25700) );
  XOR U26034 ( .A(n25699), .B(n25700), .Z(n25728) );
  NANDN U26035 ( .A(n28889), .B(n25484), .Z(n25486) );
  XOR U26036 ( .A(a[114]), .B(b[5]), .Z(n25817) );
  NANDN U26037 ( .A(n29138), .B(n25817), .Z(n25485) );
  AND U26038 ( .A(n25486), .B(n25485), .Z(n25747) );
  NANDN U26039 ( .A(n209), .B(n25487), .Z(n25489) );
  XOR U26040 ( .A(a[116]), .B(b[3]), .Z(n25820) );
  NANDN U26041 ( .A(n28941), .B(n25820), .Z(n25488) );
  AND U26042 ( .A(n25489), .B(n25488), .Z(n25746) );
  NANDN U26043 ( .A(n35936), .B(n25490), .Z(n25492) );
  XOR U26044 ( .A(b[37]), .B(a[82]), .Z(n25823) );
  NANDN U26045 ( .A(n36047), .B(n25823), .Z(n25491) );
  NAND U26046 ( .A(n25492), .B(n25491), .Z(n25745) );
  XOR U26047 ( .A(n25746), .B(n25745), .Z(n25748) );
  XNOR U26048 ( .A(n25747), .B(n25748), .Z(n25727) );
  XNOR U26049 ( .A(n25728), .B(n25727), .Z(n25729) );
  NANDN U26050 ( .A(n25494), .B(n25493), .Z(n25498) );
  OR U26051 ( .A(n25496), .B(n25495), .Z(n25497) );
  NAND U26052 ( .A(n25498), .B(n25497), .Z(n25730) );
  XOR U26053 ( .A(n25729), .B(n25730), .Z(n25833) );
  XNOR U26054 ( .A(n25832), .B(n25833), .Z(n25834) );
  XNOR U26055 ( .A(n25835), .B(n25834), .Z(n25717) );
  XOR U26056 ( .A(n25718), .B(n25717), .Z(n25611) );
  XNOR U26057 ( .A(n25611), .B(n25610), .Z(n25612) );
  XNOR U26058 ( .A(n25613), .B(n25612), .Z(n25574) );
  XOR U26059 ( .A(n25575), .B(n25574), .Z(n25577) );
  XOR U26060 ( .A(n25576), .B(n25577), .Z(n25570) );
  NANDN U26061 ( .A(n25504), .B(n25503), .Z(n25508) );
  OR U26062 ( .A(n25506), .B(n25505), .Z(n25507) );
  AND U26063 ( .A(n25508), .B(n25507), .Z(n25569) );
  NANDN U26064 ( .A(n25510), .B(n25509), .Z(n25514) );
  OR U26065 ( .A(n25512), .B(n25511), .Z(n25513) );
  AND U26066 ( .A(n25514), .B(n25513), .Z(n25583) );
  NANDN U26067 ( .A(n25516), .B(n25515), .Z(n25520) );
  NANDN U26068 ( .A(n25518), .B(n25517), .Z(n25519) );
  AND U26069 ( .A(n25520), .B(n25519), .Z(n25581) );
  NANDN U26070 ( .A(n25522), .B(n25521), .Z(n25526) );
  OR U26071 ( .A(n25524), .B(n25523), .Z(n25525) );
  AND U26072 ( .A(n25526), .B(n25525), .Z(n25580) );
  XNOR U26073 ( .A(n25581), .B(n25580), .Z(n25582) );
  XNOR U26074 ( .A(n25583), .B(n25582), .Z(n25568) );
  XOR U26075 ( .A(n25569), .B(n25568), .Z(n25571) );
  XOR U26076 ( .A(n25570), .B(n25571), .Z(n25564) );
  NANDN U26077 ( .A(n25528), .B(n25527), .Z(n25532) );
  NANDN U26078 ( .A(n25530), .B(n25529), .Z(n25531) );
  AND U26079 ( .A(n25532), .B(n25531), .Z(n25563) );
  NANDN U26080 ( .A(n25534), .B(n25533), .Z(n25538) );
  OR U26081 ( .A(n25536), .B(n25535), .Z(n25537) );
  AND U26082 ( .A(n25538), .B(n25537), .Z(n25562) );
  XOR U26083 ( .A(n25563), .B(n25562), .Z(n25565) );
  XOR U26084 ( .A(n25564), .B(n25565), .Z(n25839) );
  NANDN U26085 ( .A(n25540), .B(n25539), .Z(n25544) );
  NANDN U26086 ( .A(n25542), .B(n25541), .Z(n25543) );
  AND U26087 ( .A(n25544), .B(n25543), .Z(n25838) );
  XNOR U26088 ( .A(n25839), .B(n25838), .Z(n25840) );
  NANDN U26089 ( .A(n25546), .B(n25545), .Z(n25550) );
  NAND U26090 ( .A(n25548), .B(n25547), .Z(n25549) );
  NAND U26091 ( .A(n25550), .B(n25549), .Z(n25841) );
  XNOR U26092 ( .A(n25840), .B(n25841), .Z(n25556) );
  XNOR U26093 ( .A(n25557), .B(n25556), .Z(n25558) );
  XNOR U26094 ( .A(n25559), .B(n25558), .Z(n25844) );
  XNOR U26095 ( .A(sreg[182]), .B(n25844), .Z(n25846) );
  NANDN U26096 ( .A(sreg[181]), .B(n25551), .Z(n25555) );
  NAND U26097 ( .A(n25553), .B(n25552), .Z(n25554) );
  NAND U26098 ( .A(n25555), .B(n25554), .Z(n25845) );
  XNOR U26099 ( .A(n25846), .B(n25845), .Z(c[182]) );
  NANDN U26100 ( .A(n25557), .B(n25556), .Z(n25561) );
  NANDN U26101 ( .A(n25559), .B(n25558), .Z(n25560) );
  AND U26102 ( .A(n25561), .B(n25560), .Z(n25852) );
  NANDN U26103 ( .A(n25563), .B(n25562), .Z(n25567) );
  OR U26104 ( .A(n25565), .B(n25564), .Z(n25566) );
  AND U26105 ( .A(n25567), .B(n25566), .Z(n25857) );
  NANDN U26106 ( .A(n25569), .B(n25568), .Z(n25573) );
  OR U26107 ( .A(n25571), .B(n25570), .Z(n25572) );
  AND U26108 ( .A(n25573), .B(n25572), .Z(n25855) );
  NANDN U26109 ( .A(n25575), .B(n25574), .Z(n25579) );
  OR U26110 ( .A(n25577), .B(n25576), .Z(n25578) );
  AND U26111 ( .A(n25579), .B(n25578), .Z(n26132) );
  NANDN U26112 ( .A(n25581), .B(n25580), .Z(n25585) );
  NANDN U26113 ( .A(n25583), .B(n25582), .Z(n25584) );
  AND U26114 ( .A(n25585), .B(n25584), .Z(n26131) );
  XNOR U26115 ( .A(n26132), .B(n26131), .Z(n26133) );
  NANDN U26116 ( .A(n25587), .B(n25586), .Z(n25591) );
  OR U26117 ( .A(n25589), .B(n25588), .Z(n25590) );
  AND U26118 ( .A(n25591), .B(n25590), .Z(n26125) );
  NAND U26119 ( .A(n25593), .B(n25592), .Z(n25597) );
  NAND U26120 ( .A(n25595), .B(n25594), .Z(n25596) );
  AND U26121 ( .A(n25597), .B(n25596), .Z(n25869) );
  NANDN U26122 ( .A(n25599), .B(n25598), .Z(n25603) );
  OR U26123 ( .A(n25601), .B(n25600), .Z(n25602) );
  AND U26124 ( .A(n25603), .B(n25602), .Z(n25868) );
  NANDN U26125 ( .A(n25605), .B(n25604), .Z(n25609) );
  NANDN U26126 ( .A(n25607), .B(n25606), .Z(n25608) );
  AND U26127 ( .A(n25609), .B(n25608), .Z(n25867) );
  XOR U26128 ( .A(n25868), .B(n25867), .Z(n25870) );
  XOR U26129 ( .A(n25869), .B(n25870), .Z(n26126) );
  XNOR U26130 ( .A(n26125), .B(n26126), .Z(n26127) );
  NANDN U26131 ( .A(n25611), .B(n25610), .Z(n25615) );
  NANDN U26132 ( .A(n25613), .B(n25612), .Z(n25614) );
  AND U26133 ( .A(n25615), .B(n25614), .Z(n25864) );
  NANDN U26134 ( .A(n29499), .B(n25616), .Z(n25618) );
  XOR U26135 ( .A(a[113]), .B(b[7]), .Z(n25987) );
  NANDN U26136 ( .A(n29735), .B(n25987), .Z(n25617) );
  AND U26137 ( .A(n25618), .B(n25617), .Z(n25947) );
  NANDN U26138 ( .A(n37857), .B(n25619), .Z(n25621) );
  XOR U26139 ( .A(b[55]), .B(a[65]), .Z(n25990) );
  NANDN U26140 ( .A(n37911), .B(n25990), .Z(n25620) );
  AND U26141 ( .A(n25621), .B(n25620), .Z(n25946) );
  NANDN U26142 ( .A(n35611), .B(n25622), .Z(n25624) );
  XOR U26143 ( .A(b[35]), .B(a[85]), .Z(n25993) );
  NANDN U26144 ( .A(n35801), .B(n25993), .Z(n25623) );
  NAND U26145 ( .A(n25624), .B(n25623), .Z(n25945) );
  XOR U26146 ( .A(n25946), .B(n25945), .Z(n25948) );
  XOR U26147 ( .A(n25947), .B(n25948), .Z(n26009) );
  NANDN U26148 ( .A(n25626), .B(n25625), .Z(n25630) );
  OR U26149 ( .A(n25628), .B(n25627), .Z(n25629) );
  AND U26150 ( .A(n25630), .B(n25629), .Z(n26008) );
  XNOR U26151 ( .A(n26009), .B(n26008), .Z(n26010) );
  NANDN U26152 ( .A(n25632), .B(n25631), .Z(n25636) );
  OR U26153 ( .A(n25634), .B(n25633), .Z(n25635) );
  NAND U26154 ( .A(n25636), .B(n25635), .Z(n26011) );
  XNOR U26155 ( .A(n26010), .B(n26011), .Z(n25882) );
  NANDN U26156 ( .A(n25638), .B(n25637), .Z(n25642) );
  NANDN U26157 ( .A(n25640), .B(n25639), .Z(n25641) );
  AND U26158 ( .A(n25642), .B(n25641), .Z(n25880) );
  NANDN U26159 ( .A(n211), .B(n25643), .Z(n25645) );
  XOR U26160 ( .A(b[47]), .B(a[73]), .Z(n25963) );
  NANDN U26161 ( .A(n37172), .B(n25963), .Z(n25644) );
  AND U26162 ( .A(n25645), .B(n25644), .Z(n26004) );
  NANDN U26163 ( .A(n210), .B(n25646), .Z(n25648) );
  XOR U26164 ( .A(a[111]), .B(b[9]), .Z(n25966) );
  NANDN U26165 ( .A(n30267), .B(n25966), .Z(n25647) );
  AND U26166 ( .A(n25648), .B(n25647), .Z(n26003) );
  NANDN U26167 ( .A(n212), .B(n25649), .Z(n25651) );
  XOR U26168 ( .A(b[49]), .B(a[71]), .Z(n25969) );
  NANDN U26169 ( .A(n37432), .B(n25969), .Z(n25650) );
  NAND U26170 ( .A(n25651), .B(n25650), .Z(n26002) );
  XOR U26171 ( .A(n26003), .B(n26002), .Z(n26005) );
  XOR U26172 ( .A(n26004), .B(n26005), .Z(n26027) );
  NANDN U26173 ( .A(n36742), .B(n25652), .Z(n25654) );
  XOR U26174 ( .A(b[43]), .B(a[77]), .Z(n25972) );
  NANDN U26175 ( .A(n36891), .B(n25972), .Z(n25653) );
  AND U26176 ( .A(n25654), .B(n25653), .Z(n25983) );
  NANDN U26177 ( .A(n36991), .B(n25655), .Z(n25657) );
  XOR U26178 ( .A(b[45]), .B(a[75]), .Z(n25975) );
  NANDN U26179 ( .A(n37083), .B(n25975), .Z(n25656) );
  AND U26180 ( .A(n25657), .B(n25656), .Z(n25982) );
  NANDN U26181 ( .A(n30482), .B(n25658), .Z(n25660) );
  XOR U26182 ( .A(a[109]), .B(b[11]), .Z(n25978) );
  NANDN U26183 ( .A(n30891), .B(n25978), .Z(n25659) );
  NAND U26184 ( .A(n25660), .B(n25659), .Z(n25981) );
  XOR U26185 ( .A(n25982), .B(n25981), .Z(n25984) );
  XNOR U26186 ( .A(n25983), .B(n25984), .Z(n26026) );
  XNOR U26187 ( .A(n26027), .B(n26026), .Z(n26028) );
  NANDN U26188 ( .A(n25662), .B(n25661), .Z(n25666) );
  OR U26189 ( .A(n25664), .B(n25663), .Z(n25665) );
  NAND U26190 ( .A(n25666), .B(n25665), .Z(n26029) );
  XNOR U26191 ( .A(n26028), .B(n26029), .Z(n25879) );
  XNOR U26192 ( .A(n25880), .B(n25879), .Z(n25881) );
  XOR U26193 ( .A(n25882), .B(n25881), .Z(n25892) );
  NANDN U26194 ( .A(n25668), .B(n25667), .Z(n25672) );
  NANDN U26195 ( .A(n25670), .B(n25669), .Z(n25671) );
  AND U26196 ( .A(n25672), .B(n25671), .Z(n25888) );
  NANDN U26197 ( .A(n25674), .B(n25673), .Z(n25678) );
  NANDN U26198 ( .A(n25676), .B(n25675), .Z(n25677) );
  AND U26199 ( .A(n25678), .B(n25677), .Z(n25886) );
  NANDN U26200 ( .A(n33875), .B(n25679), .Z(n25681) );
  XOR U26201 ( .A(a[95]), .B(b[25]), .Z(n25921) );
  NANDN U26202 ( .A(n33994), .B(n25921), .Z(n25680) );
  AND U26203 ( .A(n25681), .B(n25680), .Z(n26049) );
  NANDN U26204 ( .A(n32013), .B(n25682), .Z(n25684) );
  XOR U26205 ( .A(a[103]), .B(b[17]), .Z(n25924) );
  NANDN U26206 ( .A(n32292), .B(n25924), .Z(n25683) );
  AND U26207 ( .A(n25684), .B(n25683), .Z(n26048) );
  NANDN U26208 ( .A(n31536), .B(n25685), .Z(n25687) );
  XOR U26209 ( .A(a[105]), .B(b[15]), .Z(n25927) );
  NANDN U26210 ( .A(n31925), .B(n25927), .Z(n25686) );
  NAND U26211 ( .A(n25687), .B(n25686), .Z(n26047) );
  XOR U26212 ( .A(n26048), .B(n26047), .Z(n26050) );
  XOR U26213 ( .A(n26049), .B(n26050), .Z(n26114) );
  NANDN U26214 ( .A(n37526), .B(n25688), .Z(n25690) );
  XOR U26215 ( .A(b[51]), .B(a[69]), .Z(n25930) );
  NANDN U26216 ( .A(n37605), .B(n25930), .Z(n25689) );
  AND U26217 ( .A(n25690), .B(n25689), .Z(n26073) );
  NANDN U26218 ( .A(n37705), .B(n25691), .Z(n25693) );
  XOR U26219 ( .A(b[53]), .B(a[67]), .Z(n25933) );
  NANDN U26220 ( .A(n37778), .B(n25933), .Z(n25692) );
  AND U26221 ( .A(n25693), .B(n25692), .Z(n26072) );
  NANDN U26222 ( .A(n36210), .B(n25694), .Z(n25696) );
  XOR U26223 ( .A(b[39]), .B(a[81]), .Z(n25936) );
  NANDN U26224 ( .A(n36347), .B(n25936), .Z(n25695) );
  NAND U26225 ( .A(n25696), .B(n25695), .Z(n26071) );
  XOR U26226 ( .A(n26072), .B(n26071), .Z(n26074) );
  XNOR U26227 ( .A(n26073), .B(n26074), .Z(n26113) );
  XNOR U26228 ( .A(n26114), .B(n26113), .Z(n26116) );
  NANDN U26229 ( .A(n25698), .B(n25697), .Z(n25702) );
  OR U26230 ( .A(n25700), .B(n25699), .Z(n25701) );
  AND U26231 ( .A(n25702), .B(n25701), .Z(n26115) );
  XOR U26232 ( .A(n26116), .B(n26115), .Z(n25912) );
  NANDN U26233 ( .A(n25704), .B(n25703), .Z(n25708) );
  OR U26234 ( .A(n25706), .B(n25705), .Z(n25707) );
  AND U26235 ( .A(n25708), .B(n25707), .Z(n25910) );
  NANDN U26236 ( .A(n25710), .B(n25709), .Z(n25714) );
  NANDN U26237 ( .A(n25712), .B(n25711), .Z(n25713) );
  NAND U26238 ( .A(n25714), .B(n25713), .Z(n25909) );
  XNOR U26239 ( .A(n25910), .B(n25909), .Z(n25911) );
  XNOR U26240 ( .A(n25912), .B(n25911), .Z(n25885) );
  XNOR U26241 ( .A(n25886), .B(n25885), .Z(n25887) );
  XNOR U26242 ( .A(n25888), .B(n25887), .Z(n25891) );
  XNOR U26243 ( .A(n25892), .B(n25891), .Z(n25893) );
  NANDN U26244 ( .A(n25716), .B(n25715), .Z(n25720) );
  NAND U26245 ( .A(n25718), .B(n25717), .Z(n25719) );
  NAND U26246 ( .A(n25720), .B(n25719), .Z(n25894) );
  XNOR U26247 ( .A(n25893), .B(n25894), .Z(n25861) );
  NANDN U26248 ( .A(n25722), .B(n25721), .Z(n25726) );
  NANDN U26249 ( .A(n25724), .B(n25723), .Z(n25725) );
  AND U26250 ( .A(n25726), .B(n25725), .Z(n25875) );
  NANDN U26251 ( .A(n25728), .B(n25727), .Z(n25732) );
  NANDN U26252 ( .A(n25730), .B(n25729), .Z(n25731) );
  AND U26253 ( .A(n25732), .B(n25731), .Z(n25874) );
  NANDN U26254 ( .A(n25734), .B(n25733), .Z(n25738) );
  NAND U26255 ( .A(n25736), .B(n25735), .Z(n25737) );
  AND U26256 ( .A(n25738), .B(n25737), .Z(n25873) );
  XOR U26257 ( .A(n25874), .B(n25873), .Z(n25876) );
  XOR U26258 ( .A(n25875), .B(n25876), .Z(n25900) );
  NANDN U26259 ( .A(n25740), .B(n25739), .Z(n25744) );
  NANDN U26260 ( .A(n25742), .B(n25741), .Z(n25743) );
  AND U26261 ( .A(n25744), .B(n25743), .Z(n26021) );
  NANDN U26262 ( .A(n25746), .B(n25745), .Z(n25750) );
  OR U26263 ( .A(n25748), .B(n25747), .Z(n25749) );
  NAND U26264 ( .A(n25750), .B(n25749), .Z(n26020) );
  XNOR U26265 ( .A(n26021), .B(n26020), .Z(n26023) );
  NANDN U26266 ( .A(n25752), .B(n25751), .Z(n25756) );
  OR U26267 ( .A(n25754), .B(n25753), .Z(n25755) );
  AND U26268 ( .A(n25756), .B(n25755), .Z(n25918) );
  NANDN U26269 ( .A(n38278), .B(n25757), .Z(n25759) );
  XOR U26270 ( .A(b[63]), .B(a[57]), .Z(n26098) );
  NANDN U26271 ( .A(n38279), .B(n26098), .Z(n25758) );
  AND U26272 ( .A(n25759), .B(n25758), .Z(n25952) );
  NANDN U26273 ( .A(n35260), .B(n25760), .Z(n25762) );
  XOR U26274 ( .A(b[33]), .B(a[87]), .Z(n26101) );
  NANDN U26275 ( .A(n35456), .B(n26101), .Z(n25761) );
  NAND U26276 ( .A(n25762), .B(n25761), .Z(n25951) );
  XNOR U26277 ( .A(n25952), .B(n25951), .Z(n25953) );
  NAND U26278 ( .A(b[0]), .B(a[119]), .Z(n25763) );
  XNOR U26279 ( .A(b[1]), .B(n25763), .Z(n25765) );
  NANDN U26280 ( .A(b[0]), .B(a[118]), .Z(n25764) );
  NAND U26281 ( .A(n25765), .B(n25764), .Z(n25954) );
  XNOR U26282 ( .A(n25953), .B(n25954), .Z(n25915) );
  NANDN U26283 ( .A(n37974), .B(n25766), .Z(n25768) );
  XOR U26284 ( .A(b[57]), .B(a[63]), .Z(n26104) );
  NANDN U26285 ( .A(n38031), .B(n26104), .Z(n25767) );
  AND U26286 ( .A(n25768), .B(n25767), .Z(n26080) );
  NANDN U26287 ( .A(n38090), .B(n25769), .Z(n25771) );
  XOR U26288 ( .A(b[59]), .B(a[61]), .Z(n26107) );
  NANDN U26289 ( .A(n38130), .B(n26107), .Z(n25770) );
  AND U26290 ( .A(n25771), .B(n25770), .Z(n26078) );
  NANDN U26291 ( .A(n36480), .B(n25772), .Z(n25774) );
  XOR U26292 ( .A(b[41]), .B(a[79]), .Z(n26110) );
  NANDN U26293 ( .A(n36594), .B(n26110), .Z(n25773) );
  NAND U26294 ( .A(n25774), .B(n25773), .Z(n26077) );
  XNOR U26295 ( .A(n26078), .B(n26077), .Z(n26079) );
  XOR U26296 ( .A(n26080), .B(n26079), .Z(n25916) );
  XNOR U26297 ( .A(n25915), .B(n25916), .Z(n25917) );
  XNOR U26298 ( .A(n25918), .B(n25917), .Z(n26022) );
  XOR U26299 ( .A(n26023), .B(n26022), .Z(n25904) );
  NANDN U26300 ( .A(n25776), .B(n25775), .Z(n25780) );
  NAND U26301 ( .A(n25778), .B(n25777), .Z(n25779) );
  NAND U26302 ( .A(n25780), .B(n25779), .Z(n25903) );
  XNOR U26303 ( .A(n25904), .B(n25903), .Z(n25906) );
  NANDN U26304 ( .A(n25782), .B(n25781), .Z(n25786) );
  NANDN U26305 ( .A(n25784), .B(n25783), .Z(n25785) );
  AND U26306 ( .A(n25786), .B(n25785), .Z(n26122) );
  NANDN U26307 ( .A(n32996), .B(n25787), .Z(n25789) );
  XOR U26308 ( .A(a[99]), .B(b[21]), .Z(n26032) );
  NANDN U26309 ( .A(n33271), .B(n26032), .Z(n25788) );
  AND U26310 ( .A(n25789), .B(n25788), .Z(n26091) );
  NANDN U26311 ( .A(n33866), .B(n25790), .Z(n25792) );
  XOR U26312 ( .A(a[97]), .B(b[23]), .Z(n26035) );
  NANDN U26313 ( .A(n33644), .B(n26035), .Z(n25791) );
  AND U26314 ( .A(n25792), .B(n25791), .Z(n26090) );
  NANDN U26315 ( .A(n32483), .B(n25793), .Z(n25795) );
  XOR U26316 ( .A(a[101]), .B(b[19]), .Z(n26038) );
  NANDN U26317 ( .A(n32823), .B(n26038), .Z(n25794) );
  NAND U26318 ( .A(n25795), .B(n25794), .Z(n26089) );
  XOR U26319 ( .A(n26090), .B(n26089), .Z(n26092) );
  XOR U26320 ( .A(n26091), .B(n26092), .Z(n25958) );
  NANDN U26321 ( .A(n34909), .B(n25796), .Z(n25798) );
  XOR U26322 ( .A(b[31]), .B(a[89]), .Z(n26041) );
  NANDN U26323 ( .A(n35145), .B(n26041), .Z(n25797) );
  AND U26324 ( .A(n25798), .B(n25797), .Z(n25998) );
  NANDN U26325 ( .A(n38247), .B(n25799), .Z(n25801) );
  XOR U26326 ( .A(b[61]), .B(a[59]), .Z(n26044) );
  NANDN U26327 ( .A(n38248), .B(n26044), .Z(n25800) );
  AND U26328 ( .A(n25801), .B(n25800), .Z(n25997) );
  AND U26329 ( .A(b[63]), .B(a[55]), .Z(n25996) );
  XOR U26330 ( .A(n25997), .B(n25996), .Z(n25999) );
  XNOR U26331 ( .A(n25998), .B(n25999), .Z(n25957) );
  XNOR U26332 ( .A(n25958), .B(n25957), .Z(n25959) );
  NANDN U26333 ( .A(n25803), .B(n25802), .Z(n25807) );
  OR U26334 ( .A(n25805), .B(n25804), .Z(n25806) );
  NAND U26335 ( .A(n25807), .B(n25806), .Z(n25960) );
  XNOR U26336 ( .A(n25959), .B(n25960), .Z(n26119) );
  NANDN U26337 ( .A(n34223), .B(n25808), .Z(n25810) );
  XOR U26338 ( .A(b[27]), .B(a[93]), .Z(n26053) );
  NANDN U26339 ( .A(n34458), .B(n26053), .Z(n25809) );
  AND U26340 ( .A(n25810), .B(n25809), .Z(n25941) );
  NANDN U26341 ( .A(n34634), .B(n25811), .Z(n25813) );
  XOR U26342 ( .A(b[29]), .B(a[91]), .Z(n26056) );
  NANDN U26343 ( .A(n34722), .B(n26056), .Z(n25812) );
  AND U26344 ( .A(n25813), .B(n25812), .Z(n25940) );
  NANDN U26345 ( .A(n31055), .B(n25814), .Z(n25816) );
  XOR U26346 ( .A(a[107]), .B(b[13]), .Z(n26059) );
  NANDN U26347 ( .A(n31293), .B(n26059), .Z(n25815) );
  NAND U26348 ( .A(n25816), .B(n25815), .Z(n25939) );
  XOR U26349 ( .A(n25940), .B(n25939), .Z(n25942) );
  XOR U26350 ( .A(n25941), .B(n25942), .Z(n26015) );
  NANDN U26351 ( .A(n28889), .B(n25817), .Z(n25819) );
  XOR U26352 ( .A(a[115]), .B(b[5]), .Z(n26062) );
  NANDN U26353 ( .A(n29138), .B(n26062), .Z(n25818) );
  AND U26354 ( .A(n25819), .B(n25818), .Z(n26085) );
  NANDN U26355 ( .A(n209), .B(n25820), .Z(n25822) );
  XOR U26356 ( .A(a[117]), .B(b[3]), .Z(n26065) );
  NANDN U26357 ( .A(n28941), .B(n26065), .Z(n25821) );
  AND U26358 ( .A(n25822), .B(n25821), .Z(n26084) );
  NANDN U26359 ( .A(n35936), .B(n25823), .Z(n25825) );
  XOR U26360 ( .A(b[37]), .B(a[83]), .Z(n26068) );
  NANDN U26361 ( .A(n36047), .B(n26068), .Z(n25824) );
  NAND U26362 ( .A(n25825), .B(n25824), .Z(n26083) );
  XOR U26363 ( .A(n26084), .B(n26083), .Z(n26086) );
  XNOR U26364 ( .A(n26085), .B(n26086), .Z(n26014) );
  XNOR U26365 ( .A(n26015), .B(n26014), .Z(n26016) );
  NANDN U26366 ( .A(n25827), .B(n25826), .Z(n25831) );
  OR U26367 ( .A(n25829), .B(n25828), .Z(n25830) );
  NAND U26368 ( .A(n25831), .B(n25830), .Z(n26017) );
  XOR U26369 ( .A(n26016), .B(n26017), .Z(n26120) );
  XNOR U26370 ( .A(n26119), .B(n26120), .Z(n26121) );
  XNOR U26371 ( .A(n26122), .B(n26121), .Z(n25905) );
  XOR U26372 ( .A(n25906), .B(n25905), .Z(n25898) );
  NANDN U26373 ( .A(n25833), .B(n25832), .Z(n25837) );
  NANDN U26374 ( .A(n25835), .B(n25834), .Z(n25836) );
  AND U26375 ( .A(n25837), .B(n25836), .Z(n25897) );
  XNOR U26376 ( .A(n25898), .B(n25897), .Z(n25899) );
  XOR U26377 ( .A(n25900), .B(n25899), .Z(n25862) );
  XNOR U26378 ( .A(n25861), .B(n25862), .Z(n25863) );
  XOR U26379 ( .A(n25864), .B(n25863), .Z(n26128) );
  XOR U26380 ( .A(n26127), .B(n26128), .Z(n26134) );
  XOR U26381 ( .A(n26133), .B(n26134), .Z(n25856) );
  XOR U26382 ( .A(n25855), .B(n25856), .Z(n25858) );
  XOR U26383 ( .A(n25857), .B(n25858), .Z(n25850) );
  NANDN U26384 ( .A(n25839), .B(n25838), .Z(n25843) );
  NANDN U26385 ( .A(n25841), .B(n25840), .Z(n25842) );
  NAND U26386 ( .A(n25843), .B(n25842), .Z(n25849) );
  XNOR U26387 ( .A(n25850), .B(n25849), .Z(n25851) );
  XNOR U26388 ( .A(n25852), .B(n25851), .Z(n26137) );
  XNOR U26389 ( .A(sreg[183]), .B(n26137), .Z(n26139) );
  NANDN U26390 ( .A(sreg[182]), .B(n25844), .Z(n25848) );
  NAND U26391 ( .A(n25846), .B(n25845), .Z(n25847) );
  NAND U26392 ( .A(n25848), .B(n25847), .Z(n26138) );
  XNOR U26393 ( .A(n26139), .B(n26138), .Z(c[183]) );
  NANDN U26394 ( .A(n25850), .B(n25849), .Z(n25854) );
  NANDN U26395 ( .A(n25852), .B(n25851), .Z(n25853) );
  AND U26396 ( .A(n25854), .B(n25853), .Z(n26145) );
  NANDN U26397 ( .A(n25856), .B(n25855), .Z(n25860) );
  OR U26398 ( .A(n25858), .B(n25857), .Z(n25859) );
  AND U26399 ( .A(n25860), .B(n25859), .Z(n26142) );
  NANDN U26400 ( .A(n25862), .B(n25861), .Z(n25866) );
  NANDN U26401 ( .A(n25864), .B(n25863), .Z(n25865) );
  AND U26402 ( .A(n25866), .B(n25865), .Z(n26425) );
  NANDN U26403 ( .A(n25868), .B(n25867), .Z(n25872) );
  NANDN U26404 ( .A(n25870), .B(n25869), .Z(n25871) );
  NAND U26405 ( .A(n25872), .B(n25871), .Z(n26424) );
  XNOR U26406 ( .A(n26425), .B(n26424), .Z(n26427) );
  NANDN U26407 ( .A(n25874), .B(n25873), .Z(n25878) );
  OR U26408 ( .A(n25876), .B(n25875), .Z(n25877) );
  AND U26409 ( .A(n25878), .B(n25877), .Z(n26162) );
  NANDN U26410 ( .A(n25880), .B(n25879), .Z(n25884) );
  NAND U26411 ( .A(n25882), .B(n25881), .Z(n25883) );
  AND U26412 ( .A(n25884), .B(n25883), .Z(n26161) );
  NANDN U26413 ( .A(n25886), .B(n25885), .Z(n25890) );
  NANDN U26414 ( .A(n25888), .B(n25887), .Z(n25889) );
  AND U26415 ( .A(n25890), .B(n25889), .Z(n26160) );
  XOR U26416 ( .A(n26161), .B(n26160), .Z(n26163) );
  XOR U26417 ( .A(n26162), .B(n26163), .Z(n26419) );
  NANDN U26418 ( .A(n25892), .B(n25891), .Z(n25896) );
  NANDN U26419 ( .A(n25894), .B(n25893), .Z(n25895) );
  NAND U26420 ( .A(n25896), .B(n25895), .Z(n26418) );
  XNOR U26421 ( .A(n26419), .B(n26418), .Z(n26420) );
  NANDN U26422 ( .A(n25898), .B(n25897), .Z(n25902) );
  NANDN U26423 ( .A(n25900), .B(n25899), .Z(n25901) );
  AND U26424 ( .A(n25902), .B(n25901), .Z(n26157) );
  NANDN U26425 ( .A(n25904), .B(n25903), .Z(n25908) );
  NAND U26426 ( .A(n25906), .B(n25905), .Z(n25907) );
  AND U26427 ( .A(n25908), .B(n25907), .Z(n26186) );
  NANDN U26428 ( .A(n25910), .B(n25909), .Z(n25914) );
  NANDN U26429 ( .A(n25912), .B(n25911), .Z(n25913) );
  AND U26430 ( .A(n25914), .B(n25913), .Z(n26180) );
  NANDN U26431 ( .A(n25916), .B(n25915), .Z(n25920) );
  NANDN U26432 ( .A(n25918), .B(n25917), .Z(n25919) );
  AND U26433 ( .A(n25920), .B(n25919), .Z(n26179) );
  NANDN U26434 ( .A(n33875), .B(n25921), .Z(n25923) );
  XOR U26435 ( .A(a[96]), .B(b[25]), .Z(n26214) );
  NANDN U26436 ( .A(n33994), .B(n26214), .Z(n25922) );
  AND U26437 ( .A(n25923), .B(n25922), .Z(n26372) );
  NANDN U26438 ( .A(n32013), .B(n25924), .Z(n25926) );
  XOR U26439 ( .A(a[104]), .B(b[17]), .Z(n26217) );
  NANDN U26440 ( .A(n32292), .B(n26217), .Z(n25925) );
  AND U26441 ( .A(n25926), .B(n25925), .Z(n26371) );
  NANDN U26442 ( .A(n31536), .B(n25927), .Z(n25929) );
  XOR U26443 ( .A(a[106]), .B(b[15]), .Z(n26220) );
  NANDN U26444 ( .A(n31925), .B(n26220), .Z(n25928) );
  NAND U26445 ( .A(n25929), .B(n25928), .Z(n26370) );
  XOR U26446 ( .A(n26371), .B(n26370), .Z(n26373) );
  XOR U26447 ( .A(n26372), .B(n26373), .Z(n26377) );
  NANDN U26448 ( .A(n37526), .B(n25930), .Z(n25932) );
  XOR U26449 ( .A(b[51]), .B(a[70]), .Z(n26223) );
  NANDN U26450 ( .A(n37605), .B(n26223), .Z(n25931) );
  AND U26451 ( .A(n25932), .B(n25931), .Z(n26351) );
  NANDN U26452 ( .A(n37705), .B(n25933), .Z(n25935) );
  XOR U26453 ( .A(b[53]), .B(a[68]), .Z(n26226) );
  NANDN U26454 ( .A(n37778), .B(n26226), .Z(n25934) );
  AND U26455 ( .A(n25935), .B(n25934), .Z(n26350) );
  NANDN U26456 ( .A(n36210), .B(n25936), .Z(n25938) );
  XOR U26457 ( .A(b[39]), .B(a[82]), .Z(n26229) );
  NANDN U26458 ( .A(n36347), .B(n26229), .Z(n25937) );
  NAND U26459 ( .A(n25938), .B(n25937), .Z(n26349) );
  XOR U26460 ( .A(n26350), .B(n26349), .Z(n26352) );
  XNOR U26461 ( .A(n26351), .B(n26352), .Z(n26376) );
  XNOR U26462 ( .A(n26377), .B(n26376), .Z(n26379) );
  NANDN U26463 ( .A(n25940), .B(n25939), .Z(n25944) );
  OR U26464 ( .A(n25942), .B(n25941), .Z(n25943) );
  AND U26465 ( .A(n25944), .B(n25943), .Z(n26378) );
  XOR U26466 ( .A(n26379), .B(n26378), .Z(n26205) );
  NANDN U26467 ( .A(n25946), .B(n25945), .Z(n25950) );
  OR U26468 ( .A(n25948), .B(n25947), .Z(n25949) );
  AND U26469 ( .A(n25950), .B(n25949), .Z(n26203) );
  NANDN U26470 ( .A(n25952), .B(n25951), .Z(n25956) );
  NANDN U26471 ( .A(n25954), .B(n25953), .Z(n25955) );
  NAND U26472 ( .A(n25956), .B(n25955), .Z(n26202) );
  XNOR U26473 ( .A(n26203), .B(n26202), .Z(n26204) );
  XNOR U26474 ( .A(n26205), .B(n26204), .Z(n26178) );
  XOR U26475 ( .A(n26179), .B(n26178), .Z(n26181) );
  XOR U26476 ( .A(n26180), .B(n26181), .Z(n26185) );
  NANDN U26477 ( .A(n25958), .B(n25957), .Z(n25962) );
  NANDN U26478 ( .A(n25960), .B(n25959), .Z(n25961) );
  AND U26479 ( .A(n25962), .B(n25961), .Z(n26173) );
  NANDN U26480 ( .A(n211), .B(n25963), .Z(n25965) );
  XOR U26481 ( .A(b[47]), .B(a[74]), .Z(n26256) );
  NANDN U26482 ( .A(n37172), .B(n26256), .Z(n25964) );
  AND U26483 ( .A(n25965), .B(n25964), .Z(n26297) );
  NANDN U26484 ( .A(n210), .B(n25966), .Z(n25968) );
  XOR U26485 ( .A(a[112]), .B(b[9]), .Z(n26259) );
  NANDN U26486 ( .A(n30267), .B(n26259), .Z(n25967) );
  AND U26487 ( .A(n25968), .B(n25967), .Z(n26296) );
  NANDN U26488 ( .A(n212), .B(n25969), .Z(n25971) );
  XOR U26489 ( .A(b[49]), .B(a[72]), .Z(n26262) );
  NANDN U26490 ( .A(n37432), .B(n26262), .Z(n25970) );
  NAND U26491 ( .A(n25971), .B(n25970), .Z(n26295) );
  XOR U26492 ( .A(n26296), .B(n26295), .Z(n26298) );
  XOR U26493 ( .A(n26297), .B(n26298), .Z(n26326) );
  NANDN U26494 ( .A(n36742), .B(n25972), .Z(n25974) );
  XOR U26495 ( .A(b[43]), .B(a[78]), .Z(n26265) );
  NANDN U26496 ( .A(n36891), .B(n26265), .Z(n25973) );
  AND U26497 ( .A(n25974), .B(n25973), .Z(n26276) );
  NANDN U26498 ( .A(n36991), .B(n25975), .Z(n25977) );
  XOR U26499 ( .A(b[45]), .B(a[76]), .Z(n26268) );
  NANDN U26500 ( .A(n37083), .B(n26268), .Z(n25976) );
  AND U26501 ( .A(n25977), .B(n25976), .Z(n26275) );
  NANDN U26502 ( .A(n30482), .B(n25978), .Z(n25980) );
  XOR U26503 ( .A(a[110]), .B(b[11]), .Z(n26271) );
  NANDN U26504 ( .A(n30891), .B(n26271), .Z(n25979) );
  NAND U26505 ( .A(n25980), .B(n25979), .Z(n26274) );
  XOR U26506 ( .A(n26275), .B(n26274), .Z(n26277) );
  XNOR U26507 ( .A(n26276), .B(n26277), .Z(n26325) );
  XNOR U26508 ( .A(n26326), .B(n26325), .Z(n26327) );
  NANDN U26509 ( .A(n25982), .B(n25981), .Z(n25986) );
  OR U26510 ( .A(n25984), .B(n25983), .Z(n25985) );
  NAND U26511 ( .A(n25986), .B(n25985), .Z(n26328) );
  XNOR U26512 ( .A(n26327), .B(n26328), .Z(n26172) );
  XNOR U26513 ( .A(n26173), .B(n26172), .Z(n26174) );
  NANDN U26514 ( .A(n29499), .B(n25987), .Z(n25989) );
  XOR U26515 ( .A(a[114]), .B(b[7]), .Z(n26280) );
  NANDN U26516 ( .A(n29735), .B(n26280), .Z(n25988) );
  AND U26517 ( .A(n25989), .B(n25988), .Z(n26240) );
  NANDN U26518 ( .A(n37857), .B(n25990), .Z(n25992) );
  XOR U26519 ( .A(b[55]), .B(a[66]), .Z(n26283) );
  NANDN U26520 ( .A(n37911), .B(n26283), .Z(n25991) );
  AND U26521 ( .A(n25992), .B(n25991), .Z(n26239) );
  NANDN U26522 ( .A(n35611), .B(n25993), .Z(n25995) );
  XOR U26523 ( .A(b[35]), .B(a[86]), .Z(n26286) );
  NANDN U26524 ( .A(n35801), .B(n26286), .Z(n25994) );
  NAND U26525 ( .A(n25995), .B(n25994), .Z(n26238) );
  XOR U26526 ( .A(n26239), .B(n26238), .Z(n26241) );
  XOR U26527 ( .A(n26240), .B(n26241), .Z(n26302) );
  NANDN U26528 ( .A(n25997), .B(n25996), .Z(n26001) );
  OR U26529 ( .A(n25999), .B(n25998), .Z(n26000) );
  AND U26530 ( .A(n26001), .B(n26000), .Z(n26301) );
  XNOR U26531 ( .A(n26302), .B(n26301), .Z(n26303) );
  NANDN U26532 ( .A(n26003), .B(n26002), .Z(n26007) );
  OR U26533 ( .A(n26005), .B(n26004), .Z(n26006) );
  NAND U26534 ( .A(n26007), .B(n26006), .Z(n26304) );
  XOR U26535 ( .A(n26303), .B(n26304), .Z(n26175) );
  XNOR U26536 ( .A(n26174), .B(n26175), .Z(n26184) );
  XOR U26537 ( .A(n26185), .B(n26184), .Z(n26187) );
  XOR U26538 ( .A(n26186), .B(n26187), .Z(n26155) );
  NANDN U26539 ( .A(n26009), .B(n26008), .Z(n26013) );
  NANDN U26540 ( .A(n26011), .B(n26010), .Z(n26012) );
  AND U26541 ( .A(n26013), .B(n26012), .Z(n26168) );
  NANDN U26542 ( .A(n26015), .B(n26014), .Z(n26019) );
  NANDN U26543 ( .A(n26017), .B(n26016), .Z(n26018) );
  AND U26544 ( .A(n26019), .B(n26018), .Z(n26167) );
  NANDN U26545 ( .A(n26021), .B(n26020), .Z(n26025) );
  NAND U26546 ( .A(n26023), .B(n26022), .Z(n26024) );
  AND U26547 ( .A(n26025), .B(n26024), .Z(n26166) );
  XOR U26548 ( .A(n26167), .B(n26166), .Z(n26169) );
  XOR U26549 ( .A(n26168), .B(n26169), .Z(n26193) );
  NANDN U26550 ( .A(n26027), .B(n26026), .Z(n26031) );
  NANDN U26551 ( .A(n26029), .B(n26028), .Z(n26030) );
  AND U26552 ( .A(n26031), .B(n26030), .Z(n26322) );
  NANDN U26553 ( .A(n32996), .B(n26032), .Z(n26034) );
  XOR U26554 ( .A(a[100]), .B(b[21]), .Z(n26355) );
  NANDN U26555 ( .A(n33271), .B(n26355), .Z(n26033) );
  AND U26556 ( .A(n26034), .B(n26033), .Z(n26396) );
  NANDN U26557 ( .A(n33866), .B(n26035), .Z(n26037) );
  XOR U26558 ( .A(a[98]), .B(b[23]), .Z(n26358) );
  NANDN U26559 ( .A(n33644), .B(n26358), .Z(n26036) );
  AND U26560 ( .A(n26037), .B(n26036), .Z(n26395) );
  NANDN U26561 ( .A(n32483), .B(n26038), .Z(n26040) );
  XOR U26562 ( .A(a[102]), .B(b[19]), .Z(n26361) );
  NANDN U26563 ( .A(n32823), .B(n26361), .Z(n26039) );
  NAND U26564 ( .A(n26040), .B(n26039), .Z(n26394) );
  XOR U26565 ( .A(n26395), .B(n26394), .Z(n26397) );
  XOR U26566 ( .A(n26396), .B(n26397), .Z(n26251) );
  NANDN U26567 ( .A(n34909), .B(n26041), .Z(n26043) );
  XOR U26568 ( .A(b[31]), .B(a[90]), .Z(n26364) );
  NANDN U26569 ( .A(n35145), .B(n26364), .Z(n26042) );
  AND U26570 ( .A(n26043), .B(n26042), .Z(n26291) );
  NANDN U26571 ( .A(n38247), .B(n26044), .Z(n26046) );
  XOR U26572 ( .A(b[61]), .B(a[60]), .Z(n26367) );
  NANDN U26573 ( .A(n38248), .B(n26367), .Z(n26045) );
  AND U26574 ( .A(n26046), .B(n26045), .Z(n26290) );
  AND U26575 ( .A(b[63]), .B(a[56]), .Z(n26289) );
  XOR U26576 ( .A(n26290), .B(n26289), .Z(n26292) );
  XNOR U26577 ( .A(n26291), .B(n26292), .Z(n26250) );
  XNOR U26578 ( .A(n26251), .B(n26250), .Z(n26252) );
  NANDN U26579 ( .A(n26048), .B(n26047), .Z(n26052) );
  OR U26580 ( .A(n26050), .B(n26049), .Z(n26051) );
  NAND U26581 ( .A(n26052), .B(n26051), .Z(n26253) );
  XNOR U26582 ( .A(n26252), .B(n26253), .Z(n26319) );
  NANDN U26583 ( .A(n34223), .B(n26053), .Z(n26055) );
  XOR U26584 ( .A(a[94]), .B(b[27]), .Z(n26331) );
  NANDN U26585 ( .A(n34458), .B(n26331), .Z(n26054) );
  AND U26586 ( .A(n26055), .B(n26054), .Z(n26234) );
  NANDN U26587 ( .A(n34634), .B(n26056), .Z(n26058) );
  XOR U26588 ( .A(b[29]), .B(a[92]), .Z(n26334) );
  NANDN U26589 ( .A(n34722), .B(n26334), .Z(n26057) );
  AND U26590 ( .A(n26058), .B(n26057), .Z(n26233) );
  NANDN U26591 ( .A(n31055), .B(n26059), .Z(n26061) );
  XOR U26592 ( .A(a[108]), .B(b[13]), .Z(n26337) );
  NANDN U26593 ( .A(n31293), .B(n26337), .Z(n26060) );
  NAND U26594 ( .A(n26061), .B(n26060), .Z(n26232) );
  XOR U26595 ( .A(n26233), .B(n26232), .Z(n26235) );
  XOR U26596 ( .A(n26234), .B(n26235), .Z(n26308) );
  NANDN U26597 ( .A(n28889), .B(n26062), .Z(n26064) );
  XOR U26598 ( .A(a[116]), .B(b[5]), .Z(n26340) );
  NANDN U26599 ( .A(n29138), .B(n26340), .Z(n26063) );
  AND U26600 ( .A(n26064), .B(n26063), .Z(n26390) );
  NANDN U26601 ( .A(n209), .B(n26065), .Z(n26067) );
  XOR U26602 ( .A(a[118]), .B(b[3]), .Z(n26343) );
  NANDN U26603 ( .A(n28941), .B(n26343), .Z(n26066) );
  AND U26604 ( .A(n26067), .B(n26066), .Z(n26389) );
  NANDN U26605 ( .A(n35936), .B(n26068), .Z(n26070) );
  XOR U26606 ( .A(b[37]), .B(a[84]), .Z(n26346) );
  NANDN U26607 ( .A(n36047), .B(n26346), .Z(n26069) );
  NAND U26608 ( .A(n26070), .B(n26069), .Z(n26388) );
  XOR U26609 ( .A(n26389), .B(n26388), .Z(n26391) );
  XNOR U26610 ( .A(n26390), .B(n26391), .Z(n26307) );
  XNOR U26611 ( .A(n26308), .B(n26307), .Z(n26309) );
  NANDN U26612 ( .A(n26072), .B(n26071), .Z(n26076) );
  OR U26613 ( .A(n26074), .B(n26073), .Z(n26075) );
  NAND U26614 ( .A(n26076), .B(n26075), .Z(n26310) );
  XOR U26615 ( .A(n26309), .B(n26310), .Z(n26320) );
  XNOR U26616 ( .A(n26319), .B(n26320), .Z(n26321) );
  XNOR U26617 ( .A(n26322), .B(n26321), .Z(n26199) );
  NANDN U26618 ( .A(n26078), .B(n26077), .Z(n26082) );
  NANDN U26619 ( .A(n26080), .B(n26079), .Z(n26081) );
  AND U26620 ( .A(n26082), .B(n26081), .Z(n26314) );
  NANDN U26621 ( .A(n26084), .B(n26083), .Z(n26088) );
  OR U26622 ( .A(n26086), .B(n26085), .Z(n26087) );
  NAND U26623 ( .A(n26088), .B(n26087), .Z(n26313) );
  XNOR U26624 ( .A(n26314), .B(n26313), .Z(n26316) );
  NANDN U26625 ( .A(n26090), .B(n26089), .Z(n26094) );
  OR U26626 ( .A(n26092), .B(n26091), .Z(n26093) );
  AND U26627 ( .A(n26094), .B(n26093), .Z(n26211) );
  NAND U26628 ( .A(b[0]), .B(a[120]), .Z(n26095) );
  XNOR U26629 ( .A(b[1]), .B(n26095), .Z(n26097) );
  NANDN U26630 ( .A(b[0]), .B(a[119]), .Z(n26096) );
  NAND U26631 ( .A(n26097), .B(n26096), .Z(n26247) );
  NANDN U26632 ( .A(n38278), .B(n26098), .Z(n26100) );
  XOR U26633 ( .A(b[63]), .B(a[58]), .Z(n26403) );
  NANDN U26634 ( .A(n38279), .B(n26403), .Z(n26099) );
  AND U26635 ( .A(n26100), .B(n26099), .Z(n26245) );
  NANDN U26636 ( .A(n35260), .B(n26101), .Z(n26103) );
  XOR U26637 ( .A(b[33]), .B(a[88]), .Z(n26406) );
  NANDN U26638 ( .A(n35456), .B(n26406), .Z(n26102) );
  NAND U26639 ( .A(n26103), .B(n26102), .Z(n26244) );
  XNOR U26640 ( .A(n26245), .B(n26244), .Z(n26246) );
  XNOR U26641 ( .A(n26247), .B(n26246), .Z(n26208) );
  NANDN U26642 ( .A(n37974), .B(n26104), .Z(n26106) );
  XOR U26643 ( .A(b[57]), .B(a[64]), .Z(n26409) );
  NANDN U26644 ( .A(n38031), .B(n26409), .Z(n26105) );
  AND U26645 ( .A(n26106), .B(n26105), .Z(n26385) );
  NANDN U26646 ( .A(n38090), .B(n26107), .Z(n26109) );
  XOR U26647 ( .A(b[59]), .B(a[62]), .Z(n26412) );
  NANDN U26648 ( .A(n38130), .B(n26412), .Z(n26108) );
  AND U26649 ( .A(n26109), .B(n26108), .Z(n26383) );
  NANDN U26650 ( .A(n36480), .B(n26110), .Z(n26112) );
  XOR U26651 ( .A(b[41]), .B(a[80]), .Z(n26415) );
  NANDN U26652 ( .A(n36594), .B(n26415), .Z(n26111) );
  NAND U26653 ( .A(n26112), .B(n26111), .Z(n26382) );
  XNOR U26654 ( .A(n26383), .B(n26382), .Z(n26384) );
  XOR U26655 ( .A(n26385), .B(n26384), .Z(n26209) );
  XNOR U26656 ( .A(n26208), .B(n26209), .Z(n26210) );
  XNOR U26657 ( .A(n26211), .B(n26210), .Z(n26315) );
  XOR U26658 ( .A(n26316), .B(n26315), .Z(n26197) );
  NANDN U26659 ( .A(n26114), .B(n26113), .Z(n26118) );
  NAND U26660 ( .A(n26116), .B(n26115), .Z(n26117) );
  NAND U26661 ( .A(n26118), .B(n26117), .Z(n26196) );
  XNOR U26662 ( .A(n26197), .B(n26196), .Z(n26198) );
  XOR U26663 ( .A(n26199), .B(n26198), .Z(n26191) );
  NANDN U26664 ( .A(n26120), .B(n26119), .Z(n26124) );
  NANDN U26665 ( .A(n26122), .B(n26121), .Z(n26123) );
  AND U26666 ( .A(n26124), .B(n26123), .Z(n26190) );
  XNOR U26667 ( .A(n26191), .B(n26190), .Z(n26192) );
  XNOR U26668 ( .A(n26193), .B(n26192), .Z(n26154) );
  XNOR U26669 ( .A(n26155), .B(n26154), .Z(n26156) );
  XOR U26670 ( .A(n26157), .B(n26156), .Z(n26421) );
  XNOR U26671 ( .A(n26420), .B(n26421), .Z(n26426) );
  XOR U26672 ( .A(n26427), .B(n26426), .Z(n26149) );
  NANDN U26673 ( .A(n26126), .B(n26125), .Z(n26130) );
  NANDN U26674 ( .A(n26128), .B(n26127), .Z(n26129) );
  AND U26675 ( .A(n26130), .B(n26129), .Z(n26148) );
  XNOR U26676 ( .A(n26149), .B(n26148), .Z(n26150) );
  NANDN U26677 ( .A(n26132), .B(n26131), .Z(n26136) );
  NANDN U26678 ( .A(n26134), .B(n26133), .Z(n26135) );
  NAND U26679 ( .A(n26136), .B(n26135), .Z(n26151) );
  XOR U26680 ( .A(n26150), .B(n26151), .Z(n26143) );
  XNOR U26681 ( .A(n26142), .B(n26143), .Z(n26144) );
  XNOR U26682 ( .A(n26145), .B(n26144), .Z(n26430) );
  XNOR U26683 ( .A(sreg[184]), .B(n26430), .Z(n26432) );
  NANDN U26684 ( .A(sreg[183]), .B(n26137), .Z(n26141) );
  NAND U26685 ( .A(n26139), .B(n26138), .Z(n26140) );
  NAND U26686 ( .A(n26141), .B(n26140), .Z(n26431) );
  XNOR U26687 ( .A(n26432), .B(n26431), .Z(c[184]) );
  NANDN U26688 ( .A(n26143), .B(n26142), .Z(n26147) );
  NANDN U26689 ( .A(n26145), .B(n26144), .Z(n26146) );
  AND U26690 ( .A(n26147), .B(n26146), .Z(n26438) );
  NANDN U26691 ( .A(n26149), .B(n26148), .Z(n26153) );
  NANDN U26692 ( .A(n26151), .B(n26150), .Z(n26152) );
  AND U26693 ( .A(n26153), .B(n26152), .Z(n26436) );
  NANDN U26694 ( .A(n26155), .B(n26154), .Z(n26159) );
  NANDN U26695 ( .A(n26157), .B(n26156), .Z(n26158) );
  AND U26696 ( .A(n26159), .B(n26158), .Z(n26718) );
  NANDN U26697 ( .A(n26161), .B(n26160), .Z(n26165) );
  OR U26698 ( .A(n26163), .B(n26162), .Z(n26164) );
  AND U26699 ( .A(n26165), .B(n26164), .Z(n26717) );
  XNOR U26700 ( .A(n26718), .B(n26717), .Z(n26720) );
  NANDN U26701 ( .A(n26167), .B(n26166), .Z(n26171) );
  OR U26702 ( .A(n26169), .B(n26168), .Z(n26170) );
  AND U26703 ( .A(n26171), .B(n26170), .Z(n26455) );
  NANDN U26704 ( .A(n26173), .B(n26172), .Z(n26177) );
  NANDN U26705 ( .A(n26175), .B(n26174), .Z(n26176) );
  AND U26706 ( .A(n26177), .B(n26176), .Z(n26454) );
  NANDN U26707 ( .A(n26179), .B(n26178), .Z(n26183) );
  OR U26708 ( .A(n26181), .B(n26180), .Z(n26182) );
  AND U26709 ( .A(n26183), .B(n26182), .Z(n26453) );
  XOR U26710 ( .A(n26454), .B(n26453), .Z(n26456) );
  XOR U26711 ( .A(n26455), .B(n26456), .Z(n26712) );
  NANDN U26712 ( .A(n26185), .B(n26184), .Z(n26189) );
  OR U26713 ( .A(n26187), .B(n26186), .Z(n26188) );
  AND U26714 ( .A(n26189), .B(n26188), .Z(n26711) );
  XNOR U26715 ( .A(n26712), .B(n26711), .Z(n26713) );
  NANDN U26716 ( .A(n26191), .B(n26190), .Z(n26195) );
  NANDN U26717 ( .A(n26193), .B(n26192), .Z(n26194) );
  AND U26718 ( .A(n26195), .B(n26194), .Z(n26450) );
  NANDN U26719 ( .A(n26197), .B(n26196), .Z(n26201) );
  NAND U26720 ( .A(n26199), .B(n26198), .Z(n26200) );
  AND U26721 ( .A(n26201), .B(n26200), .Z(n26479) );
  NANDN U26722 ( .A(n26203), .B(n26202), .Z(n26207) );
  NANDN U26723 ( .A(n26205), .B(n26204), .Z(n26206) );
  AND U26724 ( .A(n26207), .B(n26206), .Z(n26473) );
  NANDN U26725 ( .A(n26209), .B(n26208), .Z(n26213) );
  NANDN U26726 ( .A(n26211), .B(n26210), .Z(n26212) );
  AND U26727 ( .A(n26213), .B(n26212), .Z(n26472) );
  NANDN U26728 ( .A(n33875), .B(n26214), .Z(n26216) );
  XOR U26729 ( .A(a[97]), .B(b[25]), .Z(n26507) );
  NANDN U26730 ( .A(n33994), .B(n26507), .Z(n26215) );
  AND U26731 ( .A(n26216), .B(n26215), .Z(n26635) );
  NANDN U26732 ( .A(n32013), .B(n26217), .Z(n26219) );
  XOR U26733 ( .A(a[105]), .B(b[17]), .Z(n26510) );
  NANDN U26734 ( .A(n32292), .B(n26510), .Z(n26218) );
  AND U26735 ( .A(n26219), .B(n26218), .Z(n26634) );
  NANDN U26736 ( .A(n31536), .B(n26220), .Z(n26222) );
  XOR U26737 ( .A(a[107]), .B(b[15]), .Z(n26513) );
  NANDN U26738 ( .A(n31925), .B(n26513), .Z(n26221) );
  NAND U26739 ( .A(n26222), .B(n26221), .Z(n26633) );
  XOR U26740 ( .A(n26634), .B(n26633), .Z(n26636) );
  XOR U26741 ( .A(n26635), .B(n26636), .Z(n26700) );
  NANDN U26742 ( .A(n37526), .B(n26223), .Z(n26225) );
  XOR U26743 ( .A(b[51]), .B(a[71]), .Z(n26516) );
  NANDN U26744 ( .A(n37605), .B(n26516), .Z(n26224) );
  AND U26745 ( .A(n26225), .B(n26224), .Z(n26659) );
  NANDN U26746 ( .A(n37705), .B(n26226), .Z(n26228) );
  XOR U26747 ( .A(b[53]), .B(a[69]), .Z(n26519) );
  NANDN U26748 ( .A(n37778), .B(n26519), .Z(n26227) );
  AND U26749 ( .A(n26228), .B(n26227), .Z(n26658) );
  NANDN U26750 ( .A(n36210), .B(n26229), .Z(n26231) );
  XOR U26751 ( .A(b[39]), .B(a[83]), .Z(n26522) );
  NANDN U26752 ( .A(n36347), .B(n26522), .Z(n26230) );
  NAND U26753 ( .A(n26231), .B(n26230), .Z(n26657) );
  XOR U26754 ( .A(n26658), .B(n26657), .Z(n26660) );
  XNOR U26755 ( .A(n26659), .B(n26660), .Z(n26699) );
  XNOR U26756 ( .A(n26700), .B(n26699), .Z(n26702) );
  NANDN U26757 ( .A(n26233), .B(n26232), .Z(n26237) );
  OR U26758 ( .A(n26235), .B(n26234), .Z(n26236) );
  AND U26759 ( .A(n26237), .B(n26236), .Z(n26701) );
  XOR U26760 ( .A(n26702), .B(n26701), .Z(n26498) );
  NANDN U26761 ( .A(n26239), .B(n26238), .Z(n26243) );
  OR U26762 ( .A(n26241), .B(n26240), .Z(n26242) );
  AND U26763 ( .A(n26243), .B(n26242), .Z(n26496) );
  NANDN U26764 ( .A(n26245), .B(n26244), .Z(n26249) );
  NANDN U26765 ( .A(n26247), .B(n26246), .Z(n26248) );
  NAND U26766 ( .A(n26249), .B(n26248), .Z(n26495) );
  XNOR U26767 ( .A(n26496), .B(n26495), .Z(n26497) );
  XNOR U26768 ( .A(n26498), .B(n26497), .Z(n26471) );
  XOR U26769 ( .A(n26472), .B(n26471), .Z(n26474) );
  XOR U26770 ( .A(n26473), .B(n26474), .Z(n26478) );
  NANDN U26771 ( .A(n26251), .B(n26250), .Z(n26255) );
  NANDN U26772 ( .A(n26253), .B(n26252), .Z(n26254) );
  AND U26773 ( .A(n26255), .B(n26254), .Z(n26466) );
  NANDN U26774 ( .A(n211), .B(n26256), .Z(n26258) );
  XOR U26775 ( .A(b[47]), .B(a[75]), .Z(n26549) );
  NANDN U26776 ( .A(n37172), .B(n26549), .Z(n26257) );
  AND U26777 ( .A(n26258), .B(n26257), .Z(n26590) );
  NANDN U26778 ( .A(n210), .B(n26259), .Z(n26261) );
  XOR U26779 ( .A(a[113]), .B(b[9]), .Z(n26552) );
  NANDN U26780 ( .A(n30267), .B(n26552), .Z(n26260) );
  AND U26781 ( .A(n26261), .B(n26260), .Z(n26589) );
  NANDN U26782 ( .A(n212), .B(n26262), .Z(n26264) );
  XOR U26783 ( .A(b[49]), .B(a[73]), .Z(n26555) );
  NANDN U26784 ( .A(n37432), .B(n26555), .Z(n26263) );
  NAND U26785 ( .A(n26264), .B(n26263), .Z(n26588) );
  XOR U26786 ( .A(n26589), .B(n26588), .Z(n26591) );
  XOR U26787 ( .A(n26590), .B(n26591), .Z(n26613) );
  NANDN U26788 ( .A(n36742), .B(n26265), .Z(n26267) );
  XOR U26789 ( .A(b[43]), .B(a[79]), .Z(n26558) );
  NANDN U26790 ( .A(n36891), .B(n26558), .Z(n26266) );
  AND U26791 ( .A(n26267), .B(n26266), .Z(n26569) );
  NANDN U26792 ( .A(n36991), .B(n26268), .Z(n26270) );
  XOR U26793 ( .A(b[45]), .B(a[77]), .Z(n26561) );
  NANDN U26794 ( .A(n37083), .B(n26561), .Z(n26269) );
  AND U26795 ( .A(n26270), .B(n26269), .Z(n26568) );
  NANDN U26796 ( .A(n30482), .B(n26271), .Z(n26273) );
  XOR U26797 ( .A(a[111]), .B(b[11]), .Z(n26564) );
  NANDN U26798 ( .A(n30891), .B(n26564), .Z(n26272) );
  NAND U26799 ( .A(n26273), .B(n26272), .Z(n26567) );
  XOR U26800 ( .A(n26568), .B(n26567), .Z(n26570) );
  XNOR U26801 ( .A(n26569), .B(n26570), .Z(n26612) );
  XNOR U26802 ( .A(n26613), .B(n26612), .Z(n26614) );
  NANDN U26803 ( .A(n26275), .B(n26274), .Z(n26279) );
  OR U26804 ( .A(n26277), .B(n26276), .Z(n26278) );
  NAND U26805 ( .A(n26279), .B(n26278), .Z(n26615) );
  XNOR U26806 ( .A(n26614), .B(n26615), .Z(n26465) );
  XNOR U26807 ( .A(n26466), .B(n26465), .Z(n26467) );
  NANDN U26808 ( .A(n29499), .B(n26280), .Z(n26282) );
  XOR U26809 ( .A(a[115]), .B(b[7]), .Z(n26573) );
  NANDN U26810 ( .A(n29735), .B(n26573), .Z(n26281) );
  AND U26811 ( .A(n26282), .B(n26281), .Z(n26533) );
  NANDN U26812 ( .A(n37857), .B(n26283), .Z(n26285) );
  XOR U26813 ( .A(b[55]), .B(a[67]), .Z(n26576) );
  NANDN U26814 ( .A(n37911), .B(n26576), .Z(n26284) );
  AND U26815 ( .A(n26285), .B(n26284), .Z(n26532) );
  NANDN U26816 ( .A(n35611), .B(n26286), .Z(n26288) );
  XOR U26817 ( .A(b[35]), .B(a[87]), .Z(n26579) );
  NANDN U26818 ( .A(n35801), .B(n26579), .Z(n26287) );
  NAND U26819 ( .A(n26288), .B(n26287), .Z(n26531) );
  XOR U26820 ( .A(n26532), .B(n26531), .Z(n26534) );
  XOR U26821 ( .A(n26533), .B(n26534), .Z(n26595) );
  NANDN U26822 ( .A(n26290), .B(n26289), .Z(n26294) );
  OR U26823 ( .A(n26292), .B(n26291), .Z(n26293) );
  AND U26824 ( .A(n26294), .B(n26293), .Z(n26594) );
  XNOR U26825 ( .A(n26595), .B(n26594), .Z(n26596) );
  NANDN U26826 ( .A(n26296), .B(n26295), .Z(n26300) );
  OR U26827 ( .A(n26298), .B(n26297), .Z(n26299) );
  NAND U26828 ( .A(n26300), .B(n26299), .Z(n26597) );
  XOR U26829 ( .A(n26596), .B(n26597), .Z(n26468) );
  XNOR U26830 ( .A(n26467), .B(n26468), .Z(n26477) );
  XOR U26831 ( .A(n26478), .B(n26477), .Z(n26480) );
  XOR U26832 ( .A(n26479), .B(n26480), .Z(n26448) );
  NANDN U26833 ( .A(n26302), .B(n26301), .Z(n26306) );
  NANDN U26834 ( .A(n26304), .B(n26303), .Z(n26305) );
  AND U26835 ( .A(n26306), .B(n26305), .Z(n26461) );
  NANDN U26836 ( .A(n26308), .B(n26307), .Z(n26312) );
  NANDN U26837 ( .A(n26310), .B(n26309), .Z(n26311) );
  AND U26838 ( .A(n26312), .B(n26311), .Z(n26460) );
  NANDN U26839 ( .A(n26314), .B(n26313), .Z(n26318) );
  NAND U26840 ( .A(n26316), .B(n26315), .Z(n26317) );
  AND U26841 ( .A(n26318), .B(n26317), .Z(n26459) );
  XOR U26842 ( .A(n26460), .B(n26459), .Z(n26462) );
  XOR U26843 ( .A(n26461), .B(n26462), .Z(n26486) );
  NANDN U26844 ( .A(n26320), .B(n26319), .Z(n26324) );
  NANDN U26845 ( .A(n26322), .B(n26321), .Z(n26323) );
  AND U26846 ( .A(n26324), .B(n26323), .Z(n26483) );
  NANDN U26847 ( .A(n26326), .B(n26325), .Z(n26330) );
  NANDN U26848 ( .A(n26328), .B(n26327), .Z(n26329) );
  AND U26849 ( .A(n26330), .B(n26329), .Z(n26707) );
  NANDN U26850 ( .A(n34223), .B(n26331), .Z(n26333) );
  XOR U26851 ( .A(a[95]), .B(b[27]), .Z(n26639) );
  NANDN U26852 ( .A(n34458), .B(n26639), .Z(n26332) );
  AND U26853 ( .A(n26333), .B(n26332), .Z(n26527) );
  NANDN U26854 ( .A(n34634), .B(n26334), .Z(n26336) );
  XOR U26855 ( .A(b[29]), .B(a[93]), .Z(n26642) );
  NANDN U26856 ( .A(n34722), .B(n26642), .Z(n26335) );
  AND U26857 ( .A(n26336), .B(n26335), .Z(n26526) );
  NANDN U26858 ( .A(n31055), .B(n26337), .Z(n26339) );
  XOR U26859 ( .A(a[109]), .B(b[13]), .Z(n26645) );
  NANDN U26860 ( .A(n31293), .B(n26645), .Z(n26338) );
  NAND U26861 ( .A(n26339), .B(n26338), .Z(n26525) );
  XOR U26862 ( .A(n26526), .B(n26525), .Z(n26528) );
  XOR U26863 ( .A(n26527), .B(n26528), .Z(n26601) );
  NANDN U26864 ( .A(n28889), .B(n26340), .Z(n26342) );
  XOR U26865 ( .A(a[117]), .B(b[5]), .Z(n26648) );
  NANDN U26866 ( .A(n29138), .B(n26648), .Z(n26341) );
  AND U26867 ( .A(n26342), .B(n26341), .Z(n26671) );
  NANDN U26868 ( .A(n209), .B(n26343), .Z(n26345) );
  XOR U26869 ( .A(a[119]), .B(b[3]), .Z(n26651) );
  NANDN U26870 ( .A(n28941), .B(n26651), .Z(n26344) );
  AND U26871 ( .A(n26345), .B(n26344), .Z(n26670) );
  NANDN U26872 ( .A(n35936), .B(n26346), .Z(n26348) );
  XOR U26873 ( .A(b[37]), .B(a[85]), .Z(n26654) );
  NANDN U26874 ( .A(n36047), .B(n26654), .Z(n26347) );
  NAND U26875 ( .A(n26348), .B(n26347), .Z(n26669) );
  XOR U26876 ( .A(n26670), .B(n26669), .Z(n26672) );
  XNOR U26877 ( .A(n26671), .B(n26672), .Z(n26600) );
  XNOR U26878 ( .A(n26601), .B(n26600), .Z(n26602) );
  NANDN U26879 ( .A(n26350), .B(n26349), .Z(n26354) );
  OR U26880 ( .A(n26352), .B(n26351), .Z(n26353) );
  NAND U26881 ( .A(n26354), .B(n26353), .Z(n26603) );
  XNOR U26882 ( .A(n26602), .B(n26603), .Z(n26705) );
  NANDN U26883 ( .A(n32996), .B(n26355), .Z(n26357) );
  XOR U26884 ( .A(a[101]), .B(b[21]), .Z(n26618) );
  NANDN U26885 ( .A(n33271), .B(n26618), .Z(n26356) );
  AND U26886 ( .A(n26357), .B(n26356), .Z(n26677) );
  NANDN U26887 ( .A(n33866), .B(n26358), .Z(n26360) );
  XOR U26888 ( .A(a[99]), .B(b[23]), .Z(n26621) );
  NANDN U26889 ( .A(n33644), .B(n26621), .Z(n26359) );
  AND U26890 ( .A(n26360), .B(n26359), .Z(n26676) );
  NANDN U26891 ( .A(n32483), .B(n26361), .Z(n26363) );
  XOR U26892 ( .A(a[103]), .B(b[19]), .Z(n26624) );
  NANDN U26893 ( .A(n32823), .B(n26624), .Z(n26362) );
  NAND U26894 ( .A(n26363), .B(n26362), .Z(n26675) );
  XOR U26895 ( .A(n26676), .B(n26675), .Z(n26678) );
  XOR U26896 ( .A(n26677), .B(n26678), .Z(n26544) );
  NANDN U26897 ( .A(n34909), .B(n26364), .Z(n26366) );
  XOR U26898 ( .A(b[31]), .B(a[91]), .Z(n26627) );
  NANDN U26899 ( .A(n35145), .B(n26627), .Z(n26365) );
  AND U26900 ( .A(n26366), .B(n26365), .Z(n26584) );
  NANDN U26901 ( .A(n38247), .B(n26367), .Z(n26369) );
  XOR U26902 ( .A(b[61]), .B(a[61]), .Z(n26630) );
  NANDN U26903 ( .A(n38248), .B(n26630), .Z(n26368) );
  AND U26904 ( .A(n26369), .B(n26368), .Z(n26583) );
  AND U26905 ( .A(b[63]), .B(a[57]), .Z(n26582) );
  XOR U26906 ( .A(n26583), .B(n26582), .Z(n26585) );
  XNOR U26907 ( .A(n26584), .B(n26585), .Z(n26543) );
  XNOR U26908 ( .A(n26544), .B(n26543), .Z(n26545) );
  NANDN U26909 ( .A(n26371), .B(n26370), .Z(n26375) );
  OR U26910 ( .A(n26373), .B(n26372), .Z(n26374) );
  NAND U26911 ( .A(n26375), .B(n26374), .Z(n26546) );
  XOR U26912 ( .A(n26545), .B(n26546), .Z(n26706) );
  XOR U26913 ( .A(n26705), .B(n26706), .Z(n26708) );
  XOR U26914 ( .A(n26707), .B(n26708), .Z(n26492) );
  NANDN U26915 ( .A(n26377), .B(n26376), .Z(n26381) );
  NAND U26916 ( .A(n26379), .B(n26378), .Z(n26380) );
  AND U26917 ( .A(n26381), .B(n26380), .Z(n26489) );
  NANDN U26918 ( .A(n26383), .B(n26382), .Z(n26387) );
  NANDN U26919 ( .A(n26385), .B(n26384), .Z(n26386) );
  AND U26920 ( .A(n26387), .B(n26386), .Z(n26607) );
  NANDN U26921 ( .A(n26389), .B(n26388), .Z(n26393) );
  OR U26922 ( .A(n26391), .B(n26390), .Z(n26392) );
  NAND U26923 ( .A(n26393), .B(n26392), .Z(n26606) );
  XNOR U26924 ( .A(n26607), .B(n26606), .Z(n26608) );
  NANDN U26925 ( .A(n26395), .B(n26394), .Z(n26399) );
  OR U26926 ( .A(n26397), .B(n26396), .Z(n26398) );
  AND U26927 ( .A(n26399), .B(n26398), .Z(n26504) );
  NAND U26928 ( .A(b[0]), .B(a[121]), .Z(n26400) );
  XNOR U26929 ( .A(b[1]), .B(n26400), .Z(n26402) );
  NANDN U26930 ( .A(b[0]), .B(a[120]), .Z(n26401) );
  NAND U26931 ( .A(n26402), .B(n26401), .Z(n26540) );
  NANDN U26932 ( .A(n38278), .B(n26403), .Z(n26405) );
  XOR U26933 ( .A(b[63]), .B(a[59]), .Z(n26684) );
  NANDN U26934 ( .A(n38279), .B(n26684), .Z(n26404) );
  AND U26935 ( .A(n26405), .B(n26404), .Z(n26538) );
  NANDN U26936 ( .A(n35260), .B(n26406), .Z(n26408) );
  XOR U26937 ( .A(b[33]), .B(a[89]), .Z(n26687) );
  NANDN U26938 ( .A(n35456), .B(n26687), .Z(n26407) );
  NAND U26939 ( .A(n26408), .B(n26407), .Z(n26537) );
  XNOR U26940 ( .A(n26538), .B(n26537), .Z(n26539) );
  XNOR U26941 ( .A(n26540), .B(n26539), .Z(n26501) );
  NANDN U26942 ( .A(n37974), .B(n26409), .Z(n26411) );
  XOR U26943 ( .A(b[57]), .B(a[65]), .Z(n26690) );
  NANDN U26944 ( .A(n38031), .B(n26690), .Z(n26410) );
  AND U26945 ( .A(n26411), .B(n26410), .Z(n26666) );
  NANDN U26946 ( .A(n38090), .B(n26412), .Z(n26414) );
  XOR U26947 ( .A(b[59]), .B(a[63]), .Z(n26693) );
  NANDN U26948 ( .A(n38130), .B(n26693), .Z(n26413) );
  AND U26949 ( .A(n26414), .B(n26413), .Z(n26664) );
  NANDN U26950 ( .A(n36480), .B(n26415), .Z(n26417) );
  XOR U26951 ( .A(b[41]), .B(a[81]), .Z(n26696) );
  NANDN U26952 ( .A(n36594), .B(n26696), .Z(n26416) );
  NAND U26953 ( .A(n26417), .B(n26416), .Z(n26663) );
  XNOR U26954 ( .A(n26664), .B(n26663), .Z(n26665) );
  XOR U26955 ( .A(n26666), .B(n26665), .Z(n26502) );
  XNOR U26956 ( .A(n26501), .B(n26502), .Z(n26503) );
  XOR U26957 ( .A(n26504), .B(n26503), .Z(n26609) );
  XOR U26958 ( .A(n26608), .B(n26609), .Z(n26490) );
  XNOR U26959 ( .A(n26489), .B(n26490), .Z(n26491) );
  XOR U26960 ( .A(n26492), .B(n26491), .Z(n26484) );
  XNOR U26961 ( .A(n26483), .B(n26484), .Z(n26485) );
  XNOR U26962 ( .A(n26486), .B(n26485), .Z(n26447) );
  XNOR U26963 ( .A(n26448), .B(n26447), .Z(n26449) );
  XOR U26964 ( .A(n26450), .B(n26449), .Z(n26714) );
  XNOR U26965 ( .A(n26713), .B(n26714), .Z(n26719) );
  XOR U26966 ( .A(n26720), .B(n26719), .Z(n26442) );
  NANDN U26967 ( .A(n26419), .B(n26418), .Z(n26423) );
  NANDN U26968 ( .A(n26421), .B(n26420), .Z(n26422) );
  AND U26969 ( .A(n26423), .B(n26422), .Z(n26441) );
  XNOR U26970 ( .A(n26442), .B(n26441), .Z(n26443) );
  NANDN U26971 ( .A(n26425), .B(n26424), .Z(n26429) );
  NAND U26972 ( .A(n26427), .B(n26426), .Z(n26428) );
  NAND U26973 ( .A(n26429), .B(n26428), .Z(n26444) );
  XNOR U26974 ( .A(n26443), .B(n26444), .Z(n26435) );
  XNOR U26975 ( .A(n26436), .B(n26435), .Z(n26437) );
  XNOR U26976 ( .A(n26438), .B(n26437), .Z(n26723) );
  XNOR U26977 ( .A(sreg[185]), .B(n26723), .Z(n26725) );
  NANDN U26978 ( .A(sreg[184]), .B(n26430), .Z(n26434) );
  NAND U26979 ( .A(n26432), .B(n26431), .Z(n26433) );
  NAND U26980 ( .A(n26434), .B(n26433), .Z(n26724) );
  XNOR U26981 ( .A(n26725), .B(n26724), .Z(c[185]) );
  NANDN U26982 ( .A(n26436), .B(n26435), .Z(n26440) );
  NANDN U26983 ( .A(n26438), .B(n26437), .Z(n26439) );
  AND U26984 ( .A(n26440), .B(n26439), .Z(n26731) );
  NANDN U26985 ( .A(n26442), .B(n26441), .Z(n26446) );
  NANDN U26986 ( .A(n26444), .B(n26443), .Z(n26445) );
  AND U26987 ( .A(n26446), .B(n26445), .Z(n26729) );
  NANDN U26988 ( .A(n26448), .B(n26447), .Z(n26452) );
  NANDN U26989 ( .A(n26450), .B(n26449), .Z(n26451) );
  AND U26990 ( .A(n26452), .B(n26451), .Z(n27011) );
  NANDN U26991 ( .A(n26454), .B(n26453), .Z(n26458) );
  OR U26992 ( .A(n26456), .B(n26455), .Z(n26457) );
  AND U26993 ( .A(n26458), .B(n26457), .Z(n27010) );
  XNOR U26994 ( .A(n27011), .B(n27010), .Z(n27013) );
  NANDN U26995 ( .A(n26460), .B(n26459), .Z(n26464) );
  OR U26996 ( .A(n26462), .B(n26461), .Z(n26463) );
  AND U26997 ( .A(n26464), .B(n26463), .Z(n27000) );
  NANDN U26998 ( .A(n26466), .B(n26465), .Z(n26470) );
  NANDN U26999 ( .A(n26468), .B(n26467), .Z(n26469) );
  AND U27000 ( .A(n26470), .B(n26469), .Z(n26999) );
  NANDN U27001 ( .A(n26472), .B(n26471), .Z(n26476) );
  OR U27002 ( .A(n26474), .B(n26473), .Z(n26475) );
  AND U27003 ( .A(n26476), .B(n26475), .Z(n26998) );
  XOR U27004 ( .A(n26999), .B(n26998), .Z(n27001) );
  XOR U27005 ( .A(n27000), .B(n27001), .Z(n27005) );
  NANDN U27006 ( .A(n26478), .B(n26477), .Z(n26482) );
  OR U27007 ( .A(n26480), .B(n26479), .Z(n26481) );
  AND U27008 ( .A(n26482), .B(n26481), .Z(n27004) );
  XNOR U27009 ( .A(n27005), .B(n27004), .Z(n27006) );
  NANDN U27010 ( .A(n26484), .B(n26483), .Z(n26488) );
  NANDN U27011 ( .A(n26486), .B(n26485), .Z(n26487) );
  AND U27012 ( .A(n26488), .B(n26487), .Z(n26995) );
  NANDN U27013 ( .A(n26490), .B(n26489), .Z(n26494) );
  NANDN U27014 ( .A(n26492), .B(n26491), .Z(n26493) );
  AND U27015 ( .A(n26494), .B(n26493), .Z(n26971) );
  NANDN U27016 ( .A(n26496), .B(n26495), .Z(n26500) );
  NANDN U27017 ( .A(n26498), .B(n26497), .Z(n26499) );
  AND U27018 ( .A(n26500), .B(n26499), .Z(n26988) );
  NANDN U27019 ( .A(n26502), .B(n26501), .Z(n26506) );
  NANDN U27020 ( .A(n26504), .B(n26503), .Z(n26505) );
  AND U27021 ( .A(n26506), .B(n26505), .Z(n26987) );
  NANDN U27022 ( .A(n33875), .B(n26507), .Z(n26509) );
  XOR U27023 ( .A(a[98]), .B(b[25]), .Z(n26764) );
  NANDN U27024 ( .A(n33994), .B(n26764), .Z(n26508) );
  AND U27025 ( .A(n26509), .B(n26508), .Z(n26898) );
  NANDN U27026 ( .A(n32013), .B(n26510), .Z(n26512) );
  XOR U27027 ( .A(a[106]), .B(b[17]), .Z(n26767) );
  NANDN U27028 ( .A(n32292), .B(n26767), .Z(n26511) );
  AND U27029 ( .A(n26512), .B(n26511), .Z(n26897) );
  NANDN U27030 ( .A(n31536), .B(n26513), .Z(n26515) );
  XOR U27031 ( .A(a[108]), .B(b[15]), .Z(n26770) );
  NANDN U27032 ( .A(n31925), .B(n26770), .Z(n26514) );
  NAND U27033 ( .A(n26515), .B(n26514), .Z(n26896) );
  XOR U27034 ( .A(n26897), .B(n26896), .Z(n26899) );
  XOR U27035 ( .A(n26898), .B(n26899), .Z(n26927) );
  NANDN U27036 ( .A(n37526), .B(n26516), .Z(n26518) );
  XOR U27037 ( .A(b[51]), .B(a[72]), .Z(n26773) );
  NANDN U27038 ( .A(n37605), .B(n26773), .Z(n26517) );
  AND U27039 ( .A(n26518), .B(n26517), .Z(n26922) );
  NANDN U27040 ( .A(n37705), .B(n26519), .Z(n26521) );
  XOR U27041 ( .A(b[53]), .B(a[70]), .Z(n26776) );
  NANDN U27042 ( .A(n37778), .B(n26776), .Z(n26520) );
  AND U27043 ( .A(n26521), .B(n26520), .Z(n26921) );
  NANDN U27044 ( .A(n36210), .B(n26522), .Z(n26524) );
  XOR U27045 ( .A(b[39]), .B(a[84]), .Z(n26779) );
  NANDN U27046 ( .A(n36347), .B(n26779), .Z(n26523) );
  NAND U27047 ( .A(n26524), .B(n26523), .Z(n26920) );
  XOR U27048 ( .A(n26921), .B(n26920), .Z(n26923) );
  XNOR U27049 ( .A(n26922), .B(n26923), .Z(n26926) );
  XNOR U27050 ( .A(n26927), .B(n26926), .Z(n26929) );
  NANDN U27051 ( .A(n26526), .B(n26525), .Z(n26530) );
  OR U27052 ( .A(n26528), .B(n26527), .Z(n26529) );
  AND U27053 ( .A(n26530), .B(n26529), .Z(n26928) );
  XOR U27054 ( .A(n26929), .B(n26928), .Z(n26755) );
  NANDN U27055 ( .A(n26532), .B(n26531), .Z(n26536) );
  OR U27056 ( .A(n26534), .B(n26533), .Z(n26535) );
  AND U27057 ( .A(n26536), .B(n26535), .Z(n26753) );
  NANDN U27058 ( .A(n26538), .B(n26537), .Z(n26542) );
  NANDN U27059 ( .A(n26540), .B(n26539), .Z(n26541) );
  NAND U27060 ( .A(n26542), .B(n26541), .Z(n26752) );
  XNOR U27061 ( .A(n26753), .B(n26752), .Z(n26754) );
  XNOR U27062 ( .A(n26755), .B(n26754), .Z(n26986) );
  XOR U27063 ( .A(n26987), .B(n26986), .Z(n26989) );
  XOR U27064 ( .A(n26988), .B(n26989), .Z(n26969) );
  NANDN U27065 ( .A(n26544), .B(n26543), .Z(n26548) );
  NANDN U27066 ( .A(n26546), .B(n26545), .Z(n26547) );
  AND U27067 ( .A(n26548), .B(n26547), .Z(n26981) );
  NANDN U27068 ( .A(n211), .B(n26549), .Z(n26551) );
  XOR U27069 ( .A(b[47]), .B(a[76]), .Z(n26806) );
  NANDN U27070 ( .A(n37172), .B(n26806), .Z(n26550) );
  AND U27071 ( .A(n26551), .B(n26550), .Z(n26847) );
  NANDN U27072 ( .A(n210), .B(n26552), .Z(n26554) );
  XOR U27073 ( .A(a[114]), .B(b[9]), .Z(n26809) );
  NANDN U27074 ( .A(n30267), .B(n26809), .Z(n26553) );
  AND U27075 ( .A(n26554), .B(n26553), .Z(n26846) );
  NANDN U27076 ( .A(n212), .B(n26555), .Z(n26557) );
  XOR U27077 ( .A(b[49]), .B(a[74]), .Z(n26812) );
  NANDN U27078 ( .A(n37432), .B(n26812), .Z(n26556) );
  NAND U27079 ( .A(n26557), .B(n26556), .Z(n26845) );
  XOR U27080 ( .A(n26846), .B(n26845), .Z(n26848) );
  XOR U27081 ( .A(n26847), .B(n26848), .Z(n26876) );
  NANDN U27082 ( .A(n36742), .B(n26558), .Z(n26560) );
  XOR U27083 ( .A(b[43]), .B(a[80]), .Z(n26815) );
  NANDN U27084 ( .A(n36891), .B(n26815), .Z(n26559) );
  AND U27085 ( .A(n26560), .B(n26559), .Z(n26826) );
  NANDN U27086 ( .A(n36991), .B(n26561), .Z(n26563) );
  XOR U27087 ( .A(b[45]), .B(a[78]), .Z(n26818) );
  NANDN U27088 ( .A(n37083), .B(n26818), .Z(n26562) );
  AND U27089 ( .A(n26563), .B(n26562), .Z(n26825) );
  NANDN U27090 ( .A(n30482), .B(n26564), .Z(n26566) );
  XOR U27091 ( .A(a[112]), .B(b[11]), .Z(n26821) );
  NANDN U27092 ( .A(n30891), .B(n26821), .Z(n26565) );
  NAND U27093 ( .A(n26566), .B(n26565), .Z(n26824) );
  XOR U27094 ( .A(n26825), .B(n26824), .Z(n26827) );
  XNOR U27095 ( .A(n26826), .B(n26827), .Z(n26875) );
  XNOR U27096 ( .A(n26876), .B(n26875), .Z(n26877) );
  NANDN U27097 ( .A(n26568), .B(n26567), .Z(n26572) );
  OR U27098 ( .A(n26570), .B(n26569), .Z(n26571) );
  NAND U27099 ( .A(n26572), .B(n26571), .Z(n26878) );
  XNOR U27100 ( .A(n26877), .B(n26878), .Z(n26980) );
  XNOR U27101 ( .A(n26981), .B(n26980), .Z(n26982) );
  NANDN U27102 ( .A(n29499), .B(n26573), .Z(n26575) );
  XOR U27103 ( .A(a[116]), .B(b[7]), .Z(n26830) );
  NANDN U27104 ( .A(n29735), .B(n26830), .Z(n26574) );
  AND U27105 ( .A(n26575), .B(n26574), .Z(n26790) );
  NANDN U27106 ( .A(n37857), .B(n26576), .Z(n26578) );
  XOR U27107 ( .A(b[55]), .B(a[68]), .Z(n26833) );
  NANDN U27108 ( .A(n37911), .B(n26833), .Z(n26577) );
  AND U27109 ( .A(n26578), .B(n26577), .Z(n26789) );
  NANDN U27110 ( .A(n35611), .B(n26579), .Z(n26581) );
  XOR U27111 ( .A(b[35]), .B(a[88]), .Z(n26836) );
  NANDN U27112 ( .A(n35801), .B(n26836), .Z(n26580) );
  NAND U27113 ( .A(n26581), .B(n26580), .Z(n26788) );
  XOR U27114 ( .A(n26789), .B(n26788), .Z(n26791) );
  XOR U27115 ( .A(n26790), .B(n26791), .Z(n26852) );
  NANDN U27116 ( .A(n26583), .B(n26582), .Z(n26587) );
  OR U27117 ( .A(n26585), .B(n26584), .Z(n26586) );
  AND U27118 ( .A(n26587), .B(n26586), .Z(n26851) );
  XNOR U27119 ( .A(n26852), .B(n26851), .Z(n26853) );
  NANDN U27120 ( .A(n26589), .B(n26588), .Z(n26593) );
  OR U27121 ( .A(n26591), .B(n26590), .Z(n26592) );
  NAND U27122 ( .A(n26593), .B(n26592), .Z(n26854) );
  XOR U27123 ( .A(n26853), .B(n26854), .Z(n26983) );
  XNOR U27124 ( .A(n26982), .B(n26983), .Z(n26968) );
  XNOR U27125 ( .A(n26969), .B(n26968), .Z(n26970) );
  XOR U27126 ( .A(n26971), .B(n26970), .Z(n26993) );
  NANDN U27127 ( .A(n26595), .B(n26594), .Z(n26599) );
  NANDN U27128 ( .A(n26597), .B(n26596), .Z(n26598) );
  AND U27129 ( .A(n26599), .B(n26598), .Z(n26976) );
  NANDN U27130 ( .A(n26601), .B(n26600), .Z(n26605) );
  NANDN U27131 ( .A(n26603), .B(n26602), .Z(n26604) );
  AND U27132 ( .A(n26605), .B(n26604), .Z(n26975) );
  NANDN U27133 ( .A(n26607), .B(n26606), .Z(n26611) );
  NANDN U27134 ( .A(n26609), .B(n26608), .Z(n26610) );
  AND U27135 ( .A(n26611), .B(n26610), .Z(n26974) );
  XOR U27136 ( .A(n26975), .B(n26974), .Z(n26977) );
  XOR U27137 ( .A(n26976), .B(n26977), .Z(n26743) );
  NANDN U27138 ( .A(n26613), .B(n26612), .Z(n26617) );
  NANDN U27139 ( .A(n26615), .B(n26614), .Z(n26616) );
  AND U27140 ( .A(n26617), .B(n26616), .Z(n26872) );
  NANDN U27141 ( .A(n32996), .B(n26618), .Z(n26620) );
  XOR U27142 ( .A(a[102]), .B(b[21]), .Z(n26881) );
  NANDN U27143 ( .A(n33271), .B(n26881), .Z(n26619) );
  AND U27144 ( .A(n26620), .B(n26619), .Z(n26946) );
  NANDN U27145 ( .A(n33866), .B(n26621), .Z(n26623) );
  XOR U27146 ( .A(a[100]), .B(b[23]), .Z(n26884) );
  NANDN U27147 ( .A(n33644), .B(n26884), .Z(n26622) );
  AND U27148 ( .A(n26623), .B(n26622), .Z(n26945) );
  NANDN U27149 ( .A(n32483), .B(n26624), .Z(n26626) );
  XOR U27150 ( .A(a[104]), .B(b[19]), .Z(n26887) );
  NANDN U27151 ( .A(n32823), .B(n26887), .Z(n26625) );
  NAND U27152 ( .A(n26626), .B(n26625), .Z(n26944) );
  XOR U27153 ( .A(n26945), .B(n26944), .Z(n26947) );
  XOR U27154 ( .A(n26946), .B(n26947), .Z(n26801) );
  NANDN U27155 ( .A(n34909), .B(n26627), .Z(n26629) );
  XOR U27156 ( .A(b[31]), .B(a[92]), .Z(n26890) );
  NANDN U27157 ( .A(n35145), .B(n26890), .Z(n26628) );
  AND U27158 ( .A(n26629), .B(n26628), .Z(n26841) );
  NANDN U27159 ( .A(n38247), .B(n26630), .Z(n26632) );
  XOR U27160 ( .A(b[61]), .B(a[62]), .Z(n26893) );
  NANDN U27161 ( .A(n38248), .B(n26893), .Z(n26631) );
  AND U27162 ( .A(n26632), .B(n26631), .Z(n26840) );
  AND U27163 ( .A(b[63]), .B(a[58]), .Z(n26839) );
  XOR U27164 ( .A(n26840), .B(n26839), .Z(n26842) );
  XNOR U27165 ( .A(n26841), .B(n26842), .Z(n26800) );
  XNOR U27166 ( .A(n26801), .B(n26800), .Z(n26802) );
  NANDN U27167 ( .A(n26634), .B(n26633), .Z(n26638) );
  OR U27168 ( .A(n26636), .B(n26635), .Z(n26637) );
  NAND U27169 ( .A(n26638), .B(n26637), .Z(n26803) );
  XNOR U27170 ( .A(n26802), .B(n26803), .Z(n26869) );
  NANDN U27171 ( .A(n34223), .B(n26639), .Z(n26641) );
  XOR U27172 ( .A(a[96]), .B(b[27]), .Z(n26902) );
  NANDN U27173 ( .A(n34458), .B(n26902), .Z(n26640) );
  AND U27174 ( .A(n26641), .B(n26640), .Z(n26784) );
  NANDN U27175 ( .A(n34634), .B(n26642), .Z(n26644) );
  XOR U27176 ( .A(b[29]), .B(a[94]), .Z(n26905) );
  NANDN U27177 ( .A(n34722), .B(n26905), .Z(n26643) );
  AND U27178 ( .A(n26644), .B(n26643), .Z(n26783) );
  NANDN U27179 ( .A(n31055), .B(n26645), .Z(n26647) );
  XOR U27180 ( .A(a[110]), .B(b[13]), .Z(n26908) );
  NANDN U27181 ( .A(n31293), .B(n26908), .Z(n26646) );
  NAND U27182 ( .A(n26647), .B(n26646), .Z(n26782) );
  XOR U27183 ( .A(n26783), .B(n26782), .Z(n26785) );
  XOR U27184 ( .A(n26784), .B(n26785), .Z(n26858) );
  NANDN U27185 ( .A(n28889), .B(n26648), .Z(n26650) );
  XOR U27186 ( .A(a[118]), .B(b[5]), .Z(n26911) );
  NANDN U27187 ( .A(n29138), .B(n26911), .Z(n26649) );
  AND U27188 ( .A(n26650), .B(n26649), .Z(n26940) );
  NANDN U27189 ( .A(n209), .B(n26651), .Z(n26653) );
  XOR U27190 ( .A(a[120]), .B(b[3]), .Z(n26914) );
  NANDN U27191 ( .A(n28941), .B(n26914), .Z(n26652) );
  AND U27192 ( .A(n26653), .B(n26652), .Z(n26939) );
  NANDN U27193 ( .A(n35936), .B(n26654), .Z(n26656) );
  XOR U27194 ( .A(b[37]), .B(a[86]), .Z(n26917) );
  NANDN U27195 ( .A(n36047), .B(n26917), .Z(n26655) );
  NAND U27196 ( .A(n26656), .B(n26655), .Z(n26938) );
  XOR U27197 ( .A(n26939), .B(n26938), .Z(n26941) );
  XNOR U27198 ( .A(n26940), .B(n26941), .Z(n26857) );
  XNOR U27199 ( .A(n26858), .B(n26857), .Z(n26859) );
  NANDN U27200 ( .A(n26658), .B(n26657), .Z(n26662) );
  OR U27201 ( .A(n26660), .B(n26659), .Z(n26661) );
  NAND U27202 ( .A(n26662), .B(n26661), .Z(n26860) );
  XOR U27203 ( .A(n26859), .B(n26860), .Z(n26870) );
  XNOR U27204 ( .A(n26869), .B(n26870), .Z(n26871) );
  XNOR U27205 ( .A(n26872), .B(n26871), .Z(n26749) );
  NANDN U27206 ( .A(n26664), .B(n26663), .Z(n26668) );
  NANDN U27207 ( .A(n26666), .B(n26665), .Z(n26667) );
  AND U27208 ( .A(n26668), .B(n26667), .Z(n26864) );
  NANDN U27209 ( .A(n26670), .B(n26669), .Z(n26674) );
  OR U27210 ( .A(n26672), .B(n26671), .Z(n26673) );
  NAND U27211 ( .A(n26674), .B(n26673), .Z(n26863) );
  XNOR U27212 ( .A(n26864), .B(n26863), .Z(n26866) );
  NANDN U27213 ( .A(n26676), .B(n26675), .Z(n26680) );
  OR U27214 ( .A(n26678), .B(n26677), .Z(n26679) );
  AND U27215 ( .A(n26680), .B(n26679), .Z(n26761) );
  NAND U27216 ( .A(b[0]), .B(a[122]), .Z(n26681) );
  XNOR U27217 ( .A(b[1]), .B(n26681), .Z(n26683) );
  NANDN U27218 ( .A(b[0]), .B(a[121]), .Z(n26682) );
  NAND U27219 ( .A(n26683), .B(n26682), .Z(n26797) );
  NANDN U27220 ( .A(n38278), .B(n26684), .Z(n26686) );
  XOR U27221 ( .A(b[63]), .B(a[60]), .Z(n26953) );
  NANDN U27222 ( .A(n38279), .B(n26953), .Z(n26685) );
  AND U27223 ( .A(n26686), .B(n26685), .Z(n26795) );
  NANDN U27224 ( .A(n35260), .B(n26687), .Z(n26689) );
  XOR U27225 ( .A(b[33]), .B(a[90]), .Z(n26956) );
  NANDN U27226 ( .A(n35456), .B(n26956), .Z(n26688) );
  NAND U27227 ( .A(n26689), .B(n26688), .Z(n26794) );
  XNOR U27228 ( .A(n26795), .B(n26794), .Z(n26796) );
  XNOR U27229 ( .A(n26797), .B(n26796), .Z(n26758) );
  NANDN U27230 ( .A(n37974), .B(n26690), .Z(n26692) );
  XOR U27231 ( .A(b[57]), .B(a[66]), .Z(n26959) );
  NANDN U27232 ( .A(n38031), .B(n26959), .Z(n26691) );
  AND U27233 ( .A(n26692), .B(n26691), .Z(n26935) );
  NANDN U27234 ( .A(n38090), .B(n26693), .Z(n26695) );
  XOR U27235 ( .A(b[59]), .B(a[64]), .Z(n26962) );
  NANDN U27236 ( .A(n38130), .B(n26962), .Z(n26694) );
  AND U27237 ( .A(n26695), .B(n26694), .Z(n26933) );
  NANDN U27238 ( .A(n36480), .B(n26696), .Z(n26698) );
  XOR U27239 ( .A(b[41]), .B(a[82]), .Z(n26965) );
  NANDN U27240 ( .A(n36594), .B(n26965), .Z(n26697) );
  NAND U27241 ( .A(n26698), .B(n26697), .Z(n26932) );
  XNOR U27242 ( .A(n26933), .B(n26932), .Z(n26934) );
  XOR U27243 ( .A(n26935), .B(n26934), .Z(n26759) );
  XNOR U27244 ( .A(n26758), .B(n26759), .Z(n26760) );
  XNOR U27245 ( .A(n26761), .B(n26760), .Z(n26865) );
  XOR U27246 ( .A(n26866), .B(n26865), .Z(n26747) );
  NANDN U27247 ( .A(n26700), .B(n26699), .Z(n26704) );
  NAND U27248 ( .A(n26702), .B(n26701), .Z(n26703) );
  NAND U27249 ( .A(n26704), .B(n26703), .Z(n26746) );
  XNOR U27250 ( .A(n26747), .B(n26746), .Z(n26748) );
  XOR U27251 ( .A(n26749), .B(n26748), .Z(n26741) );
  NANDN U27252 ( .A(n26706), .B(n26705), .Z(n26710) );
  OR U27253 ( .A(n26708), .B(n26707), .Z(n26709) );
  AND U27254 ( .A(n26710), .B(n26709), .Z(n26740) );
  XNOR U27255 ( .A(n26741), .B(n26740), .Z(n26742) );
  XNOR U27256 ( .A(n26743), .B(n26742), .Z(n26992) );
  XNOR U27257 ( .A(n26993), .B(n26992), .Z(n26994) );
  XOR U27258 ( .A(n26995), .B(n26994), .Z(n27007) );
  XNOR U27259 ( .A(n27006), .B(n27007), .Z(n27012) );
  XOR U27260 ( .A(n27013), .B(n27012), .Z(n26735) );
  NANDN U27261 ( .A(n26712), .B(n26711), .Z(n26716) );
  NANDN U27262 ( .A(n26714), .B(n26713), .Z(n26715) );
  AND U27263 ( .A(n26716), .B(n26715), .Z(n26734) );
  XNOR U27264 ( .A(n26735), .B(n26734), .Z(n26736) );
  NANDN U27265 ( .A(n26718), .B(n26717), .Z(n26722) );
  NAND U27266 ( .A(n26720), .B(n26719), .Z(n26721) );
  NAND U27267 ( .A(n26722), .B(n26721), .Z(n26737) );
  XNOR U27268 ( .A(n26736), .B(n26737), .Z(n26728) );
  XNOR U27269 ( .A(n26729), .B(n26728), .Z(n26730) );
  XNOR U27270 ( .A(n26731), .B(n26730), .Z(n27016) );
  XNOR U27271 ( .A(sreg[186]), .B(n27016), .Z(n27018) );
  NANDN U27272 ( .A(sreg[185]), .B(n26723), .Z(n26727) );
  NAND U27273 ( .A(n26725), .B(n26724), .Z(n26726) );
  NAND U27274 ( .A(n26727), .B(n26726), .Z(n27017) );
  XNOR U27275 ( .A(n27018), .B(n27017), .Z(c[186]) );
  NANDN U27276 ( .A(n26729), .B(n26728), .Z(n26733) );
  NANDN U27277 ( .A(n26731), .B(n26730), .Z(n26732) );
  AND U27278 ( .A(n26733), .B(n26732), .Z(n27024) );
  NANDN U27279 ( .A(n26735), .B(n26734), .Z(n26739) );
  NANDN U27280 ( .A(n26737), .B(n26736), .Z(n26738) );
  AND U27281 ( .A(n26739), .B(n26738), .Z(n27022) );
  NANDN U27282 ( .A(n26741), .B(n26740), .Z(n26745) );
  NANDN U27283 ( .A(n26743), .B(n26742), .Z(n26744) );
  AND U27284 ( .A(n26745), .B(n26744), .Z(n27299) );
  NANDN U27285 ( .A(n26747), .B(n26746), .Z(n26751) );
  NAND U27286 ( .A(n26749), .B(n26748), .Z(n26750) );
  AND U27287 ( .A(n26751), .B(n26750), .Z(n27275) );
  NANDN U27288 ( .A(n26753), .B(n26752), .Z(n26757) );
  NANDN U27289 ( .A(n26755), .B(n26754), .Z(n26756) );
  AND U27290 ( .A(n26757), .B(n26756), .Z(n27293) );
  NANDN U27291 ( .A(n26759), .B(n26758), .Z(n26763) );
  NANDN U27292 ( .A(n26761), .B(n26760), .Z(n26762) );
  AND U27293 ( .A(n26763), .B(n26762), .Z(n27292) );
  NANDN U27294 ( .A(n33875), .B(n26764), .Z(n26766) );
  XOR U27295 ( .A(a[99]), .B(b[25]), .Z(n27120) );
  NANDN U27296 ( .A(n33994), .B(n27120), .Z(n26765) );
  AND U27297 ( .A(n26766), .B(n26765), .Z(n27224) );
  NANDN U27298 ( .A(n32013), .B(n26767), .Z(n26769) );
  XOR U27299 ( .A(a[107]), .B(b[17]), .Z(n27123) );
  NANDN U27300 ( .A(n32292), .B(n27123), .Z(n26768) );
  AND U27301 ( .A(n26769), .B(n26768), .Z(n27223) );
  NANDN U27302 ( .A(n31536), .B(n26770), .Z(n26772) );
  XOR U27303 ( .A(a[109]), .B(b[15]), .Z(n27126) );
  NANDN U27304 ( .A(n31925), .B(n27126), .Z(n26771) );
  NAND U27305 ( .A(n26772), .B(n26771), .Z(n27222) );
  XOR U27306 ( .A(n27223), .B(n27222), .Z(n27225) );
  XOR U27307 ( .A(n27224), .B(n27225), .Z(n27211) );
  NANDN U27308 ( .A(n37526), .B(n26773), .Z(n26775) );
  XOR U27309 ( .A(b[51]), .B(a[73]), .Z(n27129) );
  NANDN U27310 ( .A(n37605), .B(n27129), .Z(n26774) );
  AND U27311 ( .A(n26775), .B(n26774), .Z(n27245) );
  NANDN U27312 ( .A(n37705), .B(n26776), .Z(n26778) );
  XOR U27313 ( .A(b[53]), .B(a[71]), .Z(n27132) );
  NANDN U27314 ( .A(n37778), .B(n27132), .Z(n26777) );
  AND U27315 ( .A(n26778), .B(n26777), .Z(n27244) );
  NANDN U27316 ( .A(n36210), .B(n26779), .Z(n26781) );
  XOR U27317 ( .A(b[39]), .B(a[85]), .Z(n27135) );
  NANDN U27318 ( .A(n36347), .B(n27135), .Z(n26780) );
  NAND U27319 ( .A(n26781), .B(n26780), .Z(n27243) );
  XOR U27320 ( .A(n27244), .B(n27243), .Z(n27246) );
  XNOR U27321 ( .A(n27245), .B(n27246), .Z(n27210) );
  XNOR U27322 ( .A(n27211), .B(n27210), .Z(n27213) );
  NANDN U27323 ( .A(n26783), .B(n26782), .Z(n26787) );
  OR U27324 ( .A(n26785), .B(n26784), .Z(n26786) );
  AND U27325 ( .A(n26787), .B(n26786), .Z(n27212) );
  XOR U27326 ( .A(n27213), .B(n27212), .Z(n27111) );
  NANDN U27327 ( .A(n26789), .B(n26788), .Z(n26793) );
  OR U27328 ( .A(n26791), .B(n26790), .Z(n26792) );
  AND U27329 ( .A(n26793), .B(n26792), .Z(n27109) );
  NANDN U27330 ( .A(n26795), .B(n26794), .Z(n26799) );
  NANDN U27331 ( .A(n26797), .B(n26796), .Z(n26798) );
  NAND U27332 ( .A(n26799), .B(n26798), .Z(n27108) );
  XNOR U27333 ( .A(n27109), .B(n27108), .Z(n27110) );
  XNOR U27334 ( .A(n27111), .B(n27110), .Z(n27291) );
  XOR U27335 ( .A(n27292), .B(n27291), .Z(n27294) );
  XOR U27336 ( .A(n27293), .B(n27294), .Z(n27274) );
  NANDN U27337 ( .A(n26801), .B(n26800), .Z(n26805) );
  NANDN U27338 ( .A(n26803), .B(n26802), .Z(n26804) );
  AND U27339 ( .A(n26805), .B(n26804), .Z(n27286) );
  NANDN U27340 ( .A(n211), .B(n26806), .Z(n26808) );
  XOR U27341 ( .A(b[47]), .B(a[77]), .Z(n27084) );
  NANDN U27342 ( .A(n37172), .B(n27084), .Z(n26807) );
  AND U27343 ( .A(n26808), .B(n26807), .Z(n27074) );
  NANDN U27344 ( .A(n210), .B(n26809), .Z(n26811) );
  XOR U27345 ( .A(a[115]), .B(b[9]), .Z(n27087) );
  NANDN U27346 ( .A(n30267), .B(n27087), .Z(n26810) );
  AND U27347 ( .A(n26811), .B(n26810), .Z(n27073) );
  NANDN U27348 ( .A(n212), .B(n26812), .Z(n26814) );
  XOR U27349 ( .A(b[49]), .B(a[75]), .Z(n27090) );
  NANDN U27350 ( .A(n37432), .B(n27090), .Z(n26813) );
  NAND U27351 ( .A(n26814), .B(n26813), .Z(n27072) );
  XOR U27352 ( .A(n27073), .B(n27072), .Z(n27075) );
  XOR U27353 ( .A(n27074), .B(n27075), .Z(n27217) );
  NANDN U27354 ( .A(n36742), .B(n26815), .Z(n26817) );
  XOR U27355 ( .A(b[43]), .B(a[81]), .Z(n27093) );
  NANDN U27356 ( .A(n36891), .B(n27093), .Z(n26816) );
  AND U27357 ( .A(n26817), .B(n26816), .Z(n27104) );
  NANDN U27358 ( .A(n36991), .B(n26818), .Z(n26820) );
  XOR U27359 ( .A(b[45]), .B(a[79]), .Z(n27096) );
  NANDN U27360 ( .A(n37083), .B(n27096), .Z(n26819) );
  AND U27361 ( .A(n26820), .B(n26819), .Z(n27103) );
  NANDN U27362 ( .A(n30482), .B(n26821), .Z(n26823) );
  XOR U27363 ( .A(a[113]), .B(b[11]), .Z(n27099) );
  NANDN U27364 ( .A(n30891), .B(n27099), .Z(n26822) );
  NAND U27365 ( .A(n26823), .B(n26822), .Z(n27102) );
  XOR U27366 ( .A(n27103), .B(n27102), .Z(n27105) );
  XNOR U27367 ( .A(n27104), .B(n27105), .Z(n27216) );
  XNOR U27368 ( .A(n27217), .B(n27216), .Z(n27218) );
  NANDN U27369 ( .A(n26825), .B(n26824), .Z(n26829) );
  OR U27370 ( .A(n26827), .B(n26826), .Z(n26828) );
  NAND U27371 ( .A(n26829), .B(n26828), .Z(n27219) );
  XNOR U27372 ( .A(n27218), .B(n27219), .Z(n27285) );
  XNOR U27373 ( .A(n27286), .B(n27285), .Z(n27287) );
  NANDN U27374 ( .A(n29499), .B(n26830), .Z(n26832) );
  XOR U27375 ( .A(a[117]), .B(b[7]), .Z(n27057) );
  NANDN U27376 ( .A(n29735), .B(n27057), .Z(n26831) );
  AND U27377 ( .A(n26832), .B(n26831), .Z(n27146) );
  NANDN U27378 ( .A(n37857), .B(n26833), .Z(n26835) );
  XOR U27379 ( .A(b[55]), .B(a[69]), .Z(n27060) );
  NANDN U27380 ( .A(n37911), .B(n27060), .Z(n26834) );
  AND U27381 ( .A(n26835), .B(n26834), .Z(n27145) );
  NANDN U27382 ( .A(n35611), .B(n26836), .Z(n26838) );
  XOR U27383 ( .A(b[35]), .B(a[89]), .Z(n27063) );
  NANDN U27384 ( .A(n35801), .B(n27063), .Z(n26837) );
  NAND U27385 ( .A(n26838), .B(n26837), .Z(n27144) );
  XOR U27386 ( .A(n27145), .B(n27144), .Z(n27147) );
  XOR U27387 ( .A(n27146), .B(n27147), .Z(n27157) );
  NANDN U27388 ( .A(n26840), .B(n26839), .Z(n26844) );
  OR U27389 ( .A(n26842), .B(n26841), .Z(n26843) );
  AND U27390 ( .A(n26844), .B(n26843), .Z(n27156) );
  XNOR U27391 ( .A(n27157), .B(n27156), .Z(n27158) );
  NANDN U27392 ( .A(n26846), .B(n26845), .Z(n26850) );
  OR U27393 ( .A(n26848), .B(n26847), .Z(n26849) );
  NAND U27394 ( .A(n26850), .B(n26849), .Z(n27159) );
  XOR U27395 ( .A(n27158), .B(n27159), .Z(n27288) );
  XNOR U27396 ( .A(n27287), .B(n27288), .Z(n27273) );
  XOR U27397 ( .A(n27274), .B(n27273), .Z(n27276) );
  XOR U27398 ( .A(n27275), .B(n27276), .Z(n27298) );
  NANDN U27399 ( .A(n26852), .B(n26851), .Z(n26856) );
  NANDN U27400 ( .A(n26854), .B(n26853), .Z(n26855) );
  AND U27401 ( .A(n26856), .B(n26855), .Z(n27281) );
  NANDN U27402 ( .A(n26858), .B(n26857), .Z(n26862) );
  NANDN U27403 ( .A(n26860), .B(n26859), .Z(n26861) );
  AND U27404 ( .A(n26862), .B(n26861), .Z(n27280) );
  NANDN U27405 ( .A(n26864), .B(n26863), .Z(n26868) );
  NAND U27406 ( .A(n26866), .B(n26865), .Z(n26867) );
  AND U27407 ( .A(n26868), .B(n26867), .Z(n27279) );
  XOR U27408 ( .A(n27280), .B(n27279), .Z(n27282) );
  XOR U27409 ( .A(n27281), .B(n27282), .Z(n27048) );
  NANDN U27410 ( .A(n26870), .B(n26869), .Z(n26874) );
  NANDN U27411 ( .A(n26872), .B(n26871), .Z(n26873) );
  AND U27412 ( .A(n26874), .B(n26873), .Z(n27045) );
  NANDN U27413 ( .A(n26876), .B(n26875), .Z(n26880) );
  NANDN U27414 ( .A(n26878), .B(n26877), .Z(n26879) );
  AND U27415 ( .A(n26880), .B(n26879), .Z(n27269) );
  NANDN U27416 ( .A(n32996), .B(n26881), .Z(n26883) );
  XOR U27417 ( .A(a[103]), .B(b[21]), .Z(n27228) );
  NANDN U27418 ( .A(n33271), .B(n27228), .Z(n26882) );
  AND U27419 ( .A(n26883), .B(n26882), .Z(n27188) );
  NANDN U27420 ( .A(n33866), .B(n26884), .Z(n26886) );
  XOR U27421 ( .A(a[101]), .B(b[23]), .Z(n27231) );
  NANDN U27422 ( .A(n33644), .B(n27231), .Z(n26885) );
  AND U27423 ( .A(n26886), .B(n26885), .Z(n27187) );
  NANDN U27424 ( .A(n32483), .B(n26887), .Z(n26889) );
  XOR U27425 ( .A(a[105]), .B(b[19]), .Z(n27234) );
  NANDN U27426 ( .A(n32823), .B(n27234), .Z(n26888) );
  NAND U27427 ( .A(n26889), .B(n26888), .Z(n27186) );
  XOR U27428 ( .A(n27187), .B(n27186), .Z(n27189) );
  XOR U27429 ( .A(n27188), .B(n27189), .Z(n27079) );
  NANDN U27430 ( .A(n34909), .B(n26890), .Z(n26892) );
  XOR U27431 ( .A(b[31]), .B(a[93]), .Z(n27237) );
  NANDN U27432 ( .A(n35145), .B(n27237), .Z(n26891) );
  AND U27433 ( .A(n26892), .B(n26891), .Z(n27068) );
  NANDN U27434 ( .A(n38247), .B(n26893), .Z(n26895) );
  XOR U27435 ( .A(b[61]), .B(a[63]), .Z(n27240) );
  NANDN U27436 ( .A(n38248), .B(n27240), .Z(n26894) );
  AND U27437 ( .A(n26895), .B(n26894), .Z(n27067) );
  AND U27438 ( .A(b[63]), .B(a[59]), .Z(n27066) );
  XOR U27439 ( .A(n27067), .B(n27066), .Z(n27069) );
  XNOR U27440 ( .A(n27068), .B(n27069), .Z(n27078) );
  XNOR U27441 ( .A(n27079), .B(n27078), .Z(n27080) );
  NANDN U27442 ( .A(n26897), .B(n26896), .Z(n26901) );
  OR U27443 ( .A(n26899), .B(n26898), .Z(n26900) );
  NAND U27444 ( .A(n26901), .B(n26900), .Z(n27081) );
  XNOR U27445 ( .A(n27080), .B(n27081), .Z(n27267) );
  NANDN U27446 ( .A(n34223), .B(n26902), .Z(n26904) );
  XOR U27447 ( .A(a[97]), .B(b[27]), .Z(n27249) );
  NANDN U27448 ( .A(n34458), .B(n27249), .Z(n26903) );
  AND U27449 ( .A(n26904), .B(n26903), .Z(n27140) );
  NANDN U27450 ( .A(n34634), .B(n26905), .Z(n26907) );
  XOR U27451 ( .A(b[29]), .B(a[95]), .Z(n27252) );
  NANDN U27452 ( .A(n34722), .B(n27252), .Z(n26906) );
  AND U27453 ( .A(n26907), .B(n26906), .Z(n27139) );
  NANDN U27454 ( .A(n31055), .B(n26908), .Z(n26910) );
  XOR U27455 ( .A(a[111]), .B(b[13]), .Z(n27255) );
  NANDN U27456 ( .A(n31293), .B(n27255), .Z(n26909) );
  NAND U27457 ( .A(n26910), .B(n26909), .Z(n27138) );
  XOR U27458 ( .A(n27139), .B(n27138), .Z(n27141) );
  XOR U27459 ( .A(n27140), .B(n27141), .Z(n27163) );
  NANDN U27460 ( .A(n28889), .B(n26911), .Z(n26913) );
  XOR U27461 ( .A(a[119]), .B(b[5]), .Z(n27258) );
  NANDN U27462 ( .A(n29138), .B(n27258), .Z(n26912) );
  AND U27463 ( .A(n26913), .B(n26912), .Z(n27182) );
  NANDN U27464 ( .A(n209), .B(n26914), .Z(n26916) );
  XOR U27465 ( .A(a[121]), .B(b[3]), .Z(n27261) );
  NANDN U27466 ( .A(n28941), .B(n27261), .Z(n26915) );
  AND U27467 ( .A(n26916), .B(n26915), .Z(n27181) );
  NANDN U27468 ( .A(n35936), .B(n26917), .Z(n26919) );
  XOR U27469 ( .A(b[37]), .B(a[87]), .Z(n27264) );
  NANDN U27470 ( .A(n36047), .B(n27264), .Z(n26918) );
  NAND U27471 ( .A(n26919), .B(n26918), .Z(n27180) );
  XOR U27472 ( .A(n27181), .B(n27180), .Z(n27183) );
  XNOR U27473 ( .A(n27182), .B(n27183), .Z(n27162) );
  XNOR U27474 ( .A(n27163), .B(n27162), .Z(n27164) );
  NANDN U27475 ( .A(n26921), .B(n26920), .Z(n26925) );
  OR U27476 ( .A(n26923), .B(n26922), .Z(n26924) );
  NAND U27477 ( .A(n26925), .B(n26924), .Z(n27165) );
  XOR U27478 ( .A(n27164), .B(n27165), .Z(n27268) );
  XOR U27479 ( .A(n27267), .B(n27268), .Z(n27270) );
  XOR U27480 ( .A(n27269), .B(n27270), .Z(n27054) );
  NANDN U27481 ( .A(n26927), .B(n26926), .Z(n26931) );
  NAND U27482 ( .A(n26929), .B(n26928), .Z(n26930) );
  AND U27483 ( .A(n26931), .B(n26930), .Z(n27051) );
  NANDN U27484 ( .A(n26933), .B(n26932), .Z(n26937) );
  NANDN U27485 ( .A(n26935), .B(n26934), .Z(n26936) );
  AND U27486 ( .A(n26937), .B(n26936), .Z(n27169) );
  NANDN U27487 ( .A(n26939), .B(n26938), .Z(n26943) );
  OR U27488 ( .A(n26941), .B(n26940), .Z(n26942) );
  NAND U27489 ( .A(n26943), .B(n26942), .Z(n27168) );
  XNOR U27490 ( .A(n27169), .B(n27168), .Z(n27170) );
  NANDN U27491 ( .A(n26945), .B(n26944), .Z(n26949) );
  OR U27492 ( .A(n26947), .B(n26946), .Z(n26948) );
  AND U27493 ( .A(n26949), .B(n26948), .Z(n27117) );
  NAND U27494 ( .A(b[0]), .B(a[123]), .Z(n26950) );
  XNOR U27495 ( .A(b[1]), .B(n26950), .Z(n26952) );
  NANDN U27496 ( .A(b[0]), .B(a[122]), .Z(n26951) );
  NAND U27497 ( .A(n26952), .B(n26951), .Z(n27153) );
  NANDN U27498 ( .A(n38278), .B(n26953), .Z(n26955) );
  XOR U27499 ( .A(b[63]), .B(a[61]), .Z(n27192) );
  NANDN U27500 ( .A(n38279), .B(n27192), .Z(n26954) );
  AND U27501 ( .A(n26955), .B(n26954), .Z(n27151) );
  NANDN U27502 ( .A(n35260), .B(n26956), .Z(n26958) );
  XOR U27503 ( .A(b[33]), .B(a[91]), .Z(n27195) );
  NANDN U27504 ( .A(n35456), .B(n27195), .Z(n26957) );
  NAND U27505 ( .A(n26958), .B(n26957), .Z(n27150) );
  XNOR U27506 ( .A(n27151), .B(n27150), .Z(n27152) );
  XNOR U27507 ( .A(n27153), .B(n27152), .Z(n27114) );
  NANDN U27508 ( .A(n37974), .B(n26959), .Z(n26961) );
  XOR U27509 ( .A(b[57]), .B(a[67]), .Z(n27201) );
  NANDN U27510 ( .A(n38031), .B(n27201), .Z(n26960) );
  AND U27511 ( .A(n26961), .B(n26960), .Z(n27177) );
  NANDN U27512 ( .A(n38090), .B(n26962), .Z(n26964) );
  XOR U27513 ( .A(b[59]), .B(a[65]), .Z(n27204) );
  NANDN U27514 ( .A(n38130), .B(n27204), .Z(n26963) );
  AND U27515 ( .A(n26964), .B(n26963), .Z(n27175) );
  NANDN U27516 ( .A(n36480), .B(n26965), .Z(n26967) );
  XOR U27517 ( .A(b[41]), .B(a[83]), .Z(n27207) );
  NANDN U27518 ( .A(n36594), .B(n27207), .Z(n26966) );
  NAND U27519 ( .A(n26967), .B(n26966), .Z(n27174) );
  XNOR U27520 ( .A(n27175), .B(n27174), .Z(n27176) );
  XOR U27521 ( .A(n27177), .B(n27176), .Z(n27115) );
  XNOR U27522 ( .A(n27114), .B(n27115), .Z(n27116) );
  XOR U27523 ( .A(n27117), .B(n27116), .Z(n27171) );
  XOR U27524 ( .A(n27170), .B(n27171), .Z(n27052) );
  XNOR U27525 ( .A(n27051), .B(n27052), .Z(n27053) );
  XOR U27526 ( .A(n27054), .B(n27053), .Z(n27046) );
  XNOR U27527 ( .A(n27045), .B(n27046), .Z(n27047) );
  XNOR U27528 ( .A(n27048), .B(n27047), .Z(n27297) );
  XOR U27529 ( .A(n27298), .B(n27297), .Z(n27300) );
  XOR U27530 ( .A(n27299), .B(n27300), .Z(n27041) );
  NANDN U27531 ( .A(n26969), .B(n26968), .Z(n26973) );
  NAND U27532 ( .A(n26971), .B(n26970), .Z(n26972) );
  AND U27533 ( .A(n26973), .B(n26972), .Z(n27040) );
  NANDN U27534 ( .A(n26975), .B(n26974), .Z(n26979) );
  OR U27535 ( .A(n26977), .B(n26976), .Z(n26978) );
  AND U27536 ( .A(n26979), .B(n26978), .Z(n27306) );
  NANDN U27537 ( .A(n26981), .B(n26980), .Z(n26985) );
  NANDN U27538 ( .A(n26983), .B(n26982), .Z(n26984) );
  AND U27539 ( .A(n26985), .B(n26984), .Z(n27304) );
  NANDN U27540 ( .A(n26987), .B(n26986), .Z(n26991) );
  OR U27541 ( .A(n26989), .B(n26988), .Z(n26990) );
  AND U27542 ( .A(n26991), .B(n26990), .Z(n27303) );
  XNOR U27543 ( .A(n27304), .B(n27303), .Z(n27305) );
  XNOR U27544 ( .A(n27306), .B(n27305), .Z(n27039) );
  XOR U27545 ( .A(n27040), .B(n27039), .Z(n27042) );
  XOR U27546 ( .A(n27041), .B(n27042), .Z(n27035) );
  NANDN U27547 ( .A(n26993), .B(n26992), .Z(n26997) );
  NANDN U27548 ( .A(n26995), .B(n26994), .Z(n26996) );
  AND U27549 ( .A(n26997), .B(n26996), .Z(n27034) );
  NANDN U27550 ( .A(n26999), .B(n26998), .Z(n27003) );
  OR U27551 ( .A(n27001), .B(n27000), .Z(n27002) );
  AND U27552 ( .A(n27003), .B(n27002), .Z(n27033) );
  XOR U27553 ( .A(n27034), .B(n27033), .Z(n27036) );
  XOR U27554 ( .A(n27035), .B(n27036), .Z(n27028) );
  NANDN U27555 ( .A(n27005), .B(n27004), .Z(n27009) );
  NANDN U27556 ( .A(n27007), .B(n27006), .Z(n27008) );
  AND U27557 ( .A(n27009), .B(n27008), .Z(n27027) );
  XNOR U27558 ( .A(n27028), .B(n27027), .Z(n27029) );
  NANDN U27559 ( .A(n27011), .B(n27010), .Z(n27015) );
  NAND U27560 ( .A(n27013), .B(n27012), .Z(n27014) );
  NAND U27561 ( .A(n27015), .B(n27014), .Z(n27030) );
  XNOR U27562 ( .A(n27029), .B(n27030), .Z(n27021) );
  XNOR U27563 ( .A(n27022), .B(n27021), .Z(n27023) );
  XNOR U27564 ( .A(n27024), .B(n27023), .Z(n27309) );
  XNOR U27565 ( .A(sreg[187]), .B(n27309), .Z(n27311) );
  NANDN U27566 ( .A(sreg[186]), .B(n27016), .Z(n27020) );
  NAND U27567 ( .A(n27018), .B(n27017), .Z(n27019) );
  NAND U27568 ( .A(n27020), .B(n27019), .Z(n27310) );
  XNOR U27569 ( .A(n27311), .B(n27310), .Z(c[187]) );
  NANDN U27570 ( .A(n27022), .B(n27021), .Z(n27026) );
  NANDN U27571 ( .A(n27024), .B(n27023), .Z(n27025) );
  AND U27572 ( .A(n27026), .B(n27025), .Z(n27317) );
  NANDN U27573 ( .A(n27028), .B(n27027), .Z(n27032) );
  NANDN U27574 ( .A(n27030), .B(n27029), .Z(n27031) );
  AND U27575 ( .A(n27032), .B(n27031), .Z(n27315) );
  NANDN U27576 ( .A(n27034), .B(n27033), .Z(n27038) );
  OR U27577 ( .A(n27036), .B(n27035), .Z(n27037) );
  AND U27578 ( .A(n27038), .B(n27037), .Z(n27322) );
  NANDN U27579 ( .A(n27040), .B(n27039), .Z(n27044) );
  OR U27580 ( .A(n27042), .B(n27041), .Z(n27043) );
  AND U27581 ( .A(n27044), .B(n27043), .Z(n27320) );
  NANDN U27582 ( .A(n27046), .B(n27045), .Z(n27050) );
  NANDN U27583 ( .A(n27048), .B(n27047), .Z(n27049) );
  AND U27584 ( .A(n27050), .B(n27049), .Z(n27580) );
  NANDN U27585 ( .A(n27052), .B(n27051), .Z(n27056) );
  NANDN U27586 ( .A(n27054), .B(n27053), .Z(n27055) );
  AND U27587 ( .A(n27056), .B(n27055), .Z(n27347) );
  NANDN U27588 ( .A(n29499), .B(n27057), .Z(n27059) );
  XOR U27589 ( .A(a[118]), .B(b[7]), .Z(n27440) );
  NANDN U27590 ( .A(n29735), .B(n27440), .Z(n27058) );
  AND U27591 ( .A(n27059), .B(n27058), .Z(n27400) );
  NANDN U27592 ( .A(n37857), .B(n27060), .Z(n27062) );
  XOR U27593 ( .A(b[55]), .B(a[70]), .Z(n27443) );
  NANDN U27594 ( .A(n37911), .B(n27443), .Z(n27061) );
  AND U27595 ( .A(n27062), .B(n27061), .Z(n27399) );
  NANDN U27596 ( .A(n35611), .B(n27063), .Z(n27065) );
  XOR U27597 ( .A(b[35]), .B(a[90]), .Z(n27446) );
  NANDN U27598 ( .A(n35801), .B(n27446), .Z(n27064) );
  NAND U27599 ( .A(n27065), .B(n27064), .Z(n27398) );
  XOR U27600 ( .A(n27399), .B(n27398), .Z(n27401) );
  XOR U27601 ( .A(n27400), .B(n27401), .Z(n27474) );
  NANDN U27602 ( .A(n27067), .B(n27066), .Z(n27071) );
  OR U27603 ( .A(n27069), .B(n27068), .Z(n27070) );
  AND U27604 ( .A(n27071), .B(n27070), .Z(n27473) );
  XNOR U27605 ( .A(n27474), .B(n27473), .Z(n27475) );
  NANDN U27606 ( .A(n27073), .B(n27072), .Z(n27077) );
  OR U27607 ( .A(n27075), .B(n27074), .Z(n27076) );
  NAND U27608 ( .A(n27077), .B(n27076), .Z(n27476) );
  XNOR U27609 ( .A(n27475), .B(n27476), .Z(n27335) );
  NANDN U27610 ( .A(n27079), .B(n27078), .Z(n27083) );
  NANDN U27611 ( .A(n27081), .B(n27080), .Z(n27082) );
  AND U27612 ( .A(n27083), .B(n27082), .Z(n27333) );
  NAND U27613 ( .A(n37294), .B(n27084), .Z(n27086) );
  XNOR U27614 ( .A(b[47]), .B(a[78]), .Z(n27416) );
  NANDN U27615 ( .A(n27416), .B(n37341), .Z(n27085) );
  NAND U27616 ( .A(n27086), .B(n27085), .Z(n27457) );
  NAND U27617 ( .A(n30627), .B(n27087), .Z(n27089) );
  XNOR U27618 ( .A(a[116]), .B(b[9]), .Z(n27419) );
  NANDN U27619 ( .A(n27419), .B(n30628), .Z(n27088) );
  NAND U27620 ( .A(n27089), .B(n27088), .Z(n27456) );
  NAND U27621 ( .A(n37536), .B(n27090), .Z(n27092) );
  XNOR U27622 ( .A(b[49]), .B(a[76]), .Z(n27422) );
  NANDN U27623 ( .A(n27422), .B(n37537), .Z(n27091) );
  NAND U27624 ( .A(n27092), .B(n27091), .Z(n27455) );
  XOR U27625 ( .A(n27456), .B(n27455), .Z(n27458) );
  XNOR U27626 ( .A(n27457), .B(n27458), .Z(n27486) );
  NANDN U27627 ( .A(n36742), .B(n27093), .Z(n27095) );
  XOR U27628 ( .A(b[43]), .B(a[82]), .Z(n27425) );
  NANDN U27629 ( .A(n36891), .B(n27425), .Z(n27094) );
  AND U27630 ( .A(n27095), .B(n27094), .Z(n27436) );
  NANDN U27631 ( .A(n36991), .B(n27096), .Z(n27098) );
  XOR U27632 ( .A(b[45]), .B(a[80]), .Z(n27428) );
  NANDN U27633 ( .A(n37083), .B(n27428), .Z(n27097) );
  AND U27634 ( .A(n27098), .B(n27097), .Z(n27435) );
  NANDN U27635 ( .A(n30482), .B(n27099), .Z(n27101) );
  XOR U27636 ( .A(a[114]), .B(b[11]), .Z(n27431) );
  NANDN U27637 ( .A(n30891), .B(n27431), .Z(n27100) );
  NAND U27638 ( .A(n27101), .B(n27100), .Z(n27434) );
  XOR U27639 ( .A(n27435), .B(n27434), .Z(n27437) );
  XNOR U27640 ( .A(n27436), .B(n27437), .Z(n27485) );
  XOR U27641 ( .A(n27486), .B(n27485), .Z(n27487) );
  NANDN U27642 ( .A(n27103), .B(n27102), .Z(n27107) );
  OR U27643 ( .A(n27105), .B(n27104), .Z(n27106) );
  NAND U27644 ( .A(n27107), .B(n27106), .Z(n27488) );
  XNOR U27645 ( .A(n27487), .B(n27488), .Z(n27332) );
  XNOR U27646 ( .A(n27333), .B(n27332), .Z(n27334) );
  XOR U27647 ( .A(n27335), .B(n27334), .Z(n27345) );
  NANDN U27648 ( .A(n27109), .B(n27108), .Z(n27113) );
  NANDN U27649 ( .A(n27111), .B(n27110), .Z(n27112) );
  AND U27650 ( .A(n27113), .B(n27112), .Z(n27341) );
  NANDN U27651 ( .A(n27115), .B(n27114), .Z(n27119) );
  NANDN U27652 ( .A(n27117), .B(n27116), .Z(n27118) );
  AND U27653 ( .A(n27119), .B(n27118), .Z(n27339) );
  NANDN U27654 ( .A(n33875), .B(n27120), .Z(n27122) );
  XOR U27655 ( .A(a[100]), .B(b[25]), .Z(n27374) );
  NANDN U27656 ( .A(n33994), .B(n27374), .Z(n27121) );
  AND U27657 ( .A(n27122), .B(n27121), .Z(n27517) );
  NANDN U27658 ( .A(n32013), .B(n27123), .Z(n27125) );
  XOR U27659 ( .A(a[108]), .B(b[17]), .Z(n27377) );
  NANDN U27660 ( .A(n32292), .B(n27377), .Z(n27124) );
  AND U27661 ( .A(n27125), .B(n27124), .Z(n27516) );
  NANDN U27662 ( .A(n31536), .B(n27126), .Z(n27128) );
  XOR U27663 ( .A(a[110]), .B(b[15]), .Z(n27380) );
  NANDN U27664 ( .A(n31925), .B(n27380), .Z(n27127) );
  NAND U27665 ( .A(n27128), .B(n27127), .Z(n27515) );
  XOR U27666 ( .A(n27516), .B(n27515), .Z(n27518) );
  XOR U27667 ( .A(n27517), .B(n27518), .Z(n27537) );
  NANDN U27668 ( .A(n37526), .B(n27129), .Z(n27131) );
  XOR U27669 ( .A(b[51]), .B(a[74]), .Z(n27383) );
  NANDN U27670 ( .A(n37605), .B(n27383), .Z(n27130) );
  AND U27671 ( .A(n27131), .B(n27130), .Z(n27511) );
  NANDN U27672 ( .A(n37705), .B(n27132), .Z(n27134) );
  XOR U27673 ( .A(b[53]), .B(a[72]), .Z(n27386) );
  NANDN U27674 ( .A(n37778), .B(n27386), .Z(n27133) );
  AND U27675 ( .A(n27134), .B(n27133), .Z(n27510) );
  NANDN U27676 ( .A(n36210), .B(n27135), .Z(n27137) );
  XOR U27677 ( .A(b[39]), .B(a[86]), .Z(n27389) );
  NANDN U27678 ( .A(n36347), .B(n27389), .Z(n27136) );
  NAND U27679 ( .A(n27137), .B(n27136), .Z(n27509) );
  XOR U27680 ( .A(n27510), .B(n27509), .Z(n27512) );
  XNOR U27681 ( .A(n27511), .B(n27512), .Z(n27536) );
  XNOR U27682 ( .A(n27537), .B(n27536), .Z(n27539) );
  NANDN U27683 ( .A(n27139), .B(n27138), .Z(n27143) );
  OR U27684 ( .A(n27141), .B(n27140), .Z(n27142) );
  AND U27685 ( .A(n27143), .B(n27142), .Z(n27538) );
  XOR U27686 ( .A(n27539), .B(n27538), .Z(n27365) );
  NANDN U27687 ( .A(n27145), .B(n27144), .Z(n27149) );
  OR U27688 ( .A(n27147), .B(n27146), .Z(n27148) );
  AND U27689 ( .A(n27149), .B(n27148), .Z(n27363) );
  NANDN U27690 ( .A(n27151), .B(n27150), .Z(n27155) );
  NANDN U27691 ( .A(n27153), .B(n27152), .Z(n27154) );
  NAND U27692 ( .A(n27155), .B(n27154), .Z(n27362) );
  XNOR U27693 ( .A(n27363), .B(n27362), .Z(n27364) );
  XNOR U27694 ( .A(n27365), .B(n27364), .Z(n27338) );
  XNOR U27695 ( .A(n27339), .B(n27338), .Z(n27340) );
  XNOR U27696 ( .A(n27341), .B(n27340), .Z(n27344) );
  XNOR U27697 ( .A(n27345), .B(n27344), .Z(n27346) );
  XNOR U27698 ( .A(n27347), .B(n27346), .Z(n27578) );
  NANDN U27699 ( .A(n27157), .B(n27156), .Z(n27161) );
  NANDN U27700 ( .A(n27159), .B(n27158), .Z(n27160) );
  AND U27701 ( .A(n27161), .B(n27160), .Z(n27328) );
  NANDN U27702 ( .A(n27163), .B(n27162), .Z(n27167) );
  NANDN U27703 ( .A(n27165), .B(n27164), .Z(n27166) );
  AND U27704 ( .A(n27167), .B(n27166), .Z(n27327) );
  NANDN U27705 ( .A(n27169), .B(n27168), .Z(n27173) );
  NANDN U27706 ( .A(n27171), .B(n27170), .Z(n27172) );
  AND U27707 ( .A(n27173), .B(n27172), .Z(n27326) );
  XOR U27708 ( .A(n27327), .B(n27326), .Z(n27329) );
  XOR U27709 ( .A(n27328), .B(n27329), .Z(n27353) );
  NANDN U27710 ( .A(n27175), .B(n27174), .Z(n27179) );
  NANDN U27711 ( .A(n27177), .B(n27176), .Z(n27178) );
  AND U27712 ( .A(n27179), .B(n27178), .Z(n27468) );
  NANDN U27713 ( .A(n27181), .B(n27180), .Z(n27185) );
  OR U27714 ( .A(n27183), .B(n27182), .Z(n27184) );
  NAND U27715 ( .A(n27185), .B(n27184), .Z(n27467) );
  XNOR U27716 ( .A(n27468), .B(n27467), .Z(n27470) );
  NANDN U27717 ( .A(n27187), .B(n27186), .Z(n27191) );
  OR U27718 ( .A(n27189), .B(n27188), .Z(n27190) );
  AND U27719 ( .A(n27191), .B(n27190), .Z(n27371) );
  NANDN U27720 ( .A(n38278), .B(n27192), .Z(n27194) );
  XOR U27721 ( .A(b[63]), .B(a[62]), .Z(n27563) );
  NANDN U27722 ( .A(n38279), .B(n27563), .Z(n27193) );
  AND U27723 ( .A(n27194), .B(n27193), .Z(n27405) );
  NANDN U27724 ( .A(n35260), .B(n27195), .Z(n27197) );
  XOR U27725 ( .A(b[33]), .B(a[92]), .Z(n27566) );
  NANDN U27726 ( .A(n35456), .B(n27566), .Z(n27196) );
  NAND U27727 ( .A(n27197), .B(n27196), .Z(n27404) );
  XNOR U27728 ( .A(n27405), .B(n27404), .Z(n27406) );
  NAND U27729 ( .A(b[0]), .B(a[124]), .Z(n27198) );
  XNOR U27730 ( .A(b[1]), .B(n27198), .Z(n27200) );
  NANDN U27731 ( .A(b[0]), .B(a[123]), .Z(n27199) );
  NAND U27732 ( .A(n27200), .B(n27199), .Z(n27407) );
  XNOR U27733 ( .A(n27406), .B(n27407), .Z(n27368) );
  NANDN U27734 ( .A(n37974), .B(n27201), .Z(n27203) );
  XOR U27735 ( .A(b[57]), .B(a[68]), .Z(n27569) );
  NANDN U27736 ( .A(n38031), .B(n27569), .Z(n27202) );
  AND U27737 ( .A(n27203), .B(n27202), .Z(n27545) );
  NANDN U27738 ( .A(n38090), .B(n27204), .Z(n27206) );
  XOR U27739 ( .A(b[59]), .B(a[66]), .Z(n27572) );
  NANDN U27740 ( .A(n38130), .B(n27572), .Z(n27205) );
  AND U27741 ( .A(n27206), .B(n27205), .Z(n27543) );
  NANDN U27742 ( .A(n36480), .B(n27207), .Z(n27209) );
  XOR U27743 ( .A(b[41]), .B(a[84]), .Z(n27575) );
  NANDN U27744 ( .A(n36594), .B(n27575), .Z(n27208) );
  NAND U27745 ( .A(n27209), .B(n27208), .Z(n27542) );
  XNOR U27746 ( .A(n27543), .B(n27542), .Z(n27544) );
  XOR U27747 ( .A(n27545), .B(n27544), .Z(n27369) );
  XNOR U27748 ( .A(n27368), .B(n27369), .Z(n27370) );
  XNOR U27749 ( .A(n27371), .B(n27370), .Z(n27469) );
  XOR U27750 ( .A(n27470), .B(n27469), .Z(n27357) );
  NANDN U27751 ( .A(n27211), .B(n27210), .Z(n27215) );
  NAND U27752 ( .A(n27213), .B(n27212), .Z(n27214) );
  NAND U27753 ( .A(n27215), .B(n27214), .Z(n27356) );
  XNOR U27754 ( .A(n27357), .B(n27356), .Z(n27359) );
  NANDN U27755 ( .A(n27217), .B(n27216), .Z(n27221) );
  NANDN U27756 ( .A(n27219), .B(n27218), .Z(n27220) );
  AND U27757 ( .A(n27221), .B(n27220), .Z(n27482) );
  NANDN U27758 ( .A(n27223), .B(n27222), .Z(n27227) );
  OR U27759 ( .A(n27225), .B(n27224), .Z(n27226) );
  AND U27760 ( .A(n27227), .B(n27226), .Z(n27412) );
  NANDN U27761 ( .A(n32996), .B(n27228), .Z(n27230) );
  XOR U27762 ( .A(a[104]), .B(b[21]), .Z(n27521) );
  NANDN U27763 ( .A(n33271), .B(n27521), .Z(n27229) );
  AND U27764 ( .A(n27230), .B(n27229), .Z(n27556) );
  NANDN U27765 ( .A(n33866), .B(n27231), .Z(n27233) );
  XOR U27766 ( .A(a[102]), .B(b[23]), .Z(n27524) );
  NANDN U27767 ( .A(n33644), .B(n27524), .Z(n27232) );
  AND U27768 ( .A(n27233), .B(n27232), .Z(n27555) );
  NANDN U27769 ( .A(n32483), .B(n27234), .Z(n27236) );
  XOR U27770 ( .A(a[106]), .B(b[19]), .Z(n27527) );
  NANDN U27771 ( .A(n32823), .B(n27527), .Z(n27235) );
  NAND U27772 ( .A(n27236), .B(n27235), .Z(n27554) );
  XOR U27773 ( .A(n27555), .B(n27554), .Z(n27557) );
  XOR U27774 ( .A(n27556), .B(n27557), .Z(n27411) );
  NANDN U27775 ( .A(n34909), .B(n27237), .Z(n27239) );
  XOR U27776 ( .A(b[31]), .B(a[94]), .Z(n27530) );
  NANDN U27777 ( .A(n35145), .B(n27530), .Z(n27238) );
  AND U27778 ( .A(n27239), .B(n27238), .Z(n27451) );
  NANDN U27779 ( .A(n38247), .B(n27240), .Z(n27242) );
  XOR U27780 ( .A(b[61]), .B(a[64]), .Z(n27533) );
  NANDN U27781 ( .A(n38248), .B(n27533), .Z(n27241) );
  AND U27782 ( .A(n27242), .B(n27241), .Z(n27450) );
  AND U27783 ( .A(b[63]), .B(a[60]), .Z(n27449) );
  XOR U27784 ( .A(n27450), .B(n27449), .Z(n27452) );
  XNOR U27785 ( .A(n27451), .B(n27452), .Z(n27410) );
  XOR U27786 ( .A(n27411), .B(n27410), .Z(n27413) );
  XNOR U27787 ( .A(n27412), .B(n27413), .Z(n27479) );
  NANDN U27788 ( .A(n27244), .B(n27243), .Z(n27248) );
  OR U27789 ( .A(n27246), .B(n27245), .Z(n27247) );
  AND U27790 ( .A(n27248), .B(n27247), .Z(n27463) );
  NANDN U27791 ( .A(n34223), .B(n27249), .Z(n27251) );
  XOR U27792 ( .A(a[98]), .B(b[27]), .Z(n27491) );
  NANDN U27793 ( .A(n34458), .B(n27491), .Z(n27250) );
  AND U27794 ( .A(n27251), .B(n27250), .Z(n27394) );
  NANDN U27795 ( .A(n34634), .B(n27252), .Z(n27254) );
  XOR U27796 ( .A(a[96]), .B(b[29]), .Z(n27494) );
  NANDN U27797 ( .A(n34722), .B(n27494), .Z(n27253) );
  AND U27798 ( .A(n27254), .B(n27253), .Z(n27393) );
  NANDN U27799 ( .A(n31055), .B(n27255), .Z(n27257) );
  XOR U27800 ( .A(a[112]), .B(b[13]), .Z(n27497) );
  NANDN U27801 ( .A(n31293), .B(n27497), .Z(n27256) );
  NAND U27802 ( .A(n27257), .B(n27256), .Z(n27392) );
  XOR U27803 ( .A(n27393), .B(n27392), .Z(n27395) );
  XOR U27804 ( .A(n27394), .B(n27395), .Z(n27462) );
  NANDN U27805 ( .A(n28889), .B(n27258), .Z(n27260) );
  XOR U27806 ( .A(a[120]), .B(b[5]), .Z(n27500) );
  NANDN U27807 ( .A(n29138), .B(n27500), .Z(n27259) );
  AND U27808 ( .A(n27260), .B(n27259), .Z(n27550) );
  NANDN U27809 ( .A(n209), .B(n27261), .Z(n27263) );
  XOR U27810 ( .A(a[122]), .B(b[3]), .Z(n27503) );
  NANDN U27811 ( .A(n28941), .B(n27503), .Z(n27262) );
  AND U27812 ( .A(n27263), .B(n27262), .Z(n27549) );
  NANDN U27813 ( .A(n35936), .B(n27264), .Z(n27266) );
  XOR U27814 ( .A(b[37]), .B(a[88]), .Z(n27506) );
  NANDN U27815 ( .A(n36047), .B(n27506), .Z(n27265) );
  NAND U27816 ( .A(n27266), .B(n27265), .Z(n27548) );
  XOR U27817 ( .A(n27549), .B(n27548), .Z(n27551) );
  XNOR U27818 ( .A(n27550), .B(n27551), .Z(n27461) );
  XOR U27819 ( .A(n27462), .B(n27461), .Z(n27464) );
  XOR U27820 ( .A(n27463), .B(n27464), .Z(n27480) );
  XNOR U27821 ( .A(n27479), .B(n27480), .Z(n27481) );
  XNOR U27822 ( .A(n27482), .B(n27481), .Z(n27358) );
  XOR U27823 ( .A(n27359), .B(n27358), .Z(n27351) );
  NANDN U27824 ( .A(n27268), .B(n27267), .Z(n27272) );
  OR U27825 ( .A(n27270), .B(n27269), .Z(n27271) );
  AND U27826 ( .A(n27272), .B(n27271), .Z(n27350) );
  XNOR U27827 ( .A(n27351), .B(n27350), .Z(n27352) );
  XOR U27828 ( .A(n27353), .B(n27352), .Z(n27579) );
  XOR U27829 ( .A(n27578), .B(n27579), .Z(n27581) );
  XOR U27830 ( .A(n27580), .B(n27581), .Z(n27592) );
  NANDN U27831 ( .A(n27274), .B(n27273), .Z(n27278) );
  OR U27832 ( .A(n27276), .B(n27275), .Z(n27277) );
  AND U27833 ( .A(n27278), .B(n27277), .Z(n27591) );
  NANDN U27834 ( .A(n27280), .B(n27279), .Z(n27284) );
  OR U27835 ( .A(n27282), .B(n27281), .Z(n27283) );
  AND U27836 ( .A(n27284), .B(n27283), .Z(n27587) );
  NANDN U27837 ( .A(n27286), .B(n27285), .Z(n27290) );
  NANDN U27838 ( .A(n27288), .B(n27287), .Z(n27289) );
  AND U27839 ( .A(n27290), .B(n27289), .Z(n27585) );
  NANDN U27840 ( .A(n27292), .B(n27291), .Z(n27296) );
  OR U27841 ( .A(n27294), .B(n27293), .Z(n27295) );
  AND U27842 ( .A(n27296), .B(n27295), .Z(n27584) );
  XNOR U27843 ( .A(n27585), .B(n27584), .Z(n27586) );
  XNOR U27844 ( .A(n27587), .B(n27586), .Z(n27590) );
  XOR U27845 ( .A(n27591), .B(n27590), .Z(n27593) );
  XOR U27846 ( .A(n27592), .B(n27593), .Z(n27599) );
  NANDN U27847 ( .A(n27298), .B(n27297), .Z(n27302) );
  OR U27848 ( .A(n27300), .B(n27299), .Z(n27301) );
  AND U27849 ( .A(n27302), .B(n27301), .Z(n27597) );
  NANDN U27850 ( .A(n27304), .B(n27303), .Z(n27308) );
  NANDN U27851 ( .A(n27306), .B(n27305), .Z(n27307) );
  AND U27852 ( .A(n27308), .B(n27307), .Z(n27596) );
  XNOR U27853 ( .A(n27597), .B(n27596), .Z(n27598) );
  XOR U27854 ( .A(n27599), .B(n27598), .Z(n27321) );
  XOR U27855 ( .A(n27320), .B(n27321), .Z(n27323) );
  XNOR U27856 ( .A(n27322), .B(n27323), .Z(n27314) );
  XNOR U27857 ( .A(n27315), .B(n27314), .Z(n27316) );
  XNOR U27858 ( .A(n27317), .B(n27316), .Z(n27602) );
  XNOR U27859 ( .A(sreg[188]), .B(n27602), .Z(n27604) );
  NANDN U27860 ( .A(sreg[187]), .B(n27309), .Z(n27313) );
  NAND U27861 ( .A(n27311), .B(n27310), .Z(n27312) );
  NAND U27862 ( .A(n27313), .B(n27312), .Z(n27603) );
  XNOR U27863 ( .A(n27604), .B(n27603), .Z(c[188]) );
  NANDN U27864 ( .A(n27315), .B(n27314), .Z(n27319) );
  NANDN U27865 ( .A(n27317), .B(n27316), .Z(n27318) );
  AND U27866 ( .A(n27319), .B(n27318), .Z(n27610) );
  NANDN U27867 ( .A(n27321), .B(n27320), .Z(n27325) );
  OR U27868 ( .A(n27323), .B(n27322), .Z(n27324) );
  AND U27869 ( .A(n27325), .B(n27324), .Z(n27607) );
  NANDN U27870 ( .A(n27327), .B(n27326), .Z(n27331) );
  OR U27871 ( .A(n27329), .B(n27328), .Z(n27330) );
  AND U27872 ( .A(n27331), .B(n27330), .Z(n27633) );
  NANDN U27873 ( .A(n27333), .B(n27332), .Z(n27337) );
  NAND U27874 ( .A(n27335), .B(n27334), .Z(n27336) );
  AND U27875 ( .A(n27337), .B(n27336), .Z(n27632) );
  NANDN U27876 ( .A(n27339), .B(n27338), .Z(n27343) );
  NANDN U27877 ( .A(n27341), .B(n27340), .Z(n27342) );
  AND U27878 ( .A(n27343), .B(n27342), .Z(n27631) );
  XOR U27879 ( .A(n27632), .B(n27631), .Z(n27634) );
  XOR U27880 ( .A(n27633), .B(n27634), .Z(n27620) );
  NANDN U27881 ( .A(n27345), .B(n27344), .Z(n27349) );
  NANDN U27882 ( .A(n27347), .B(n27346), .Z(n27348) );
  NAND U27883 ( .A(n27349), .B(n27348), .Z(n27619) );
  XNOR U27884 ( .A(n27620), .B(n27619), .Z(n27621) );
  NANDN U27885 ( .A(n27351), .B(n27350), .Z(n27355) );
  NANDN U27886 ( .A(n27353), .B(n27352), .Z(n27354) );
  AND U27887 ( .A(n27355), .B(n27354), .Z(n27628) );
  NANDN U27888 ( .A(n27357), .B(n27356), .Z(n27361) );
  NAND U27889 ( .A(n27359), .B(n27358), .Z(n27360) );
  AND U27890 ( .A(n27361), .B(n27360), .Z(n27657) );
  NANDN U27891 ( .A(n27363), .B(n27362), .Z(n27367) );
  NANDN U27892 ( .A(n27365), .B(n27364), .Z(n27366) );
  AND U27893 ( .A(n27367), .B(n27366), .Z(n27651) );
  NANDN U27894 ( .A(n27369), .B(n27368), .Z(n27373) );
  NANDN U27895 ( .A(n27371), .B(n27370), .Z(n27372) );
  AND U27896 ( .A(n27373), .B(n27372), .Z(n27650) );
  NANDN U27897 ( .A(n33875), .B(n27374), .Z(n27376) );
  XOR U27898 ( .A(a[101]), .B(b[25]), .Z(n27732) );
  NANDN U27899 ( .A(n33994), .B(n27732), .Z(n27375) );
  AND U27900 ( .A(n27376), .B(n27375), .Z(n27820) );
  NANDN U27901 ( .A(n32013), .B(n27377), .Z(n27379) );
  XOR U27902 ( .A(a[109]), .B(b[17]), .Z(n27735) );
  NANDN U27903 ( .A(n32292), .B(n27735), .Z(n27378) );
  AND U27904 ( .A(n27379), .B(n27378), .Z(n27819) );
  NANDN U27905 ( .A(n31536), .B(n27380), .Z(n27382) );
  XOR U27906 ( .A(a[111]), .B(b[15]), .Z(n27738) );
  NANDN U27907 ( .A(n31925), .B(n27738), .Z(n27381) );
  NAND U27908 ( .A(n27382), .B(n27381), .Z(n27818) );
  XOR U27909 ( .A(n27819), .B(n27818), .Z(n27821) );
  XOR U27910 ( .A(n27820), .B(n27821), .Z(n27840) );
  NANDN U27911 ( .A(n37526), .B(n27383), .Z(n27385) );
  XOR U27912 ( .A(b[51]), .B(a[75]), .Z(n27741) );
  NANDN U27913 ( .A(n37605), .B(n27741), .Z(n27384) );
  AND U27914 ( .A(n27385), .B(n27384), .Z(n27796) );
  NANDN U27915 ( .A(n37705), .B(n27386), .Z(n27388) );
  XOR U27916 ( .A(b[53]), .B(a[73]), .Z(n27744) );
  NANDN U27917 ( .A(n37778), .B(n27744), .Z(n27387) );
  AND U27918 ( .A(n27388), .B(n27387), .Z(n27795) );
  NANDN U27919 ( .A(n36210), .B(n27389), .Z(n27391) );
  XOR U27920 ( .A(b[39]), .B(a[87]), .Z(n27747) );
  NANDN U27921 ( .A(n36347), .B(n27747), .Z(n27390) );
  NAND U27922 ( .A(n27391), .B(n27390), .Z(n27794) );
  XOR U27923 ( .A(n27795), .B(n27794), .Z(n27797) );
  XNOR U27924 ( .A(n27796), .B(n27797), .Z(n27839) );
  XNOR U27925 ( .A(n27840), .B(n27839), .Z(n27842) );
  NANDN U27926 ( .A(n27393), .B(n27392), .Z(n27397) );
  OR U27927 ( .A(n27395), .B(n27394), .Z(n27396) );
  AND U27928 ( .A(n27397), .B(n27396), .Z(n27841) );
  XOR U27929 ( .A(n27842), .B(n27841), .Z(n27723) );
  NANDN U27930 ( .A(n27399), .B(n27398), .Z(n27403) );
  OR U27931 ( .A(n27401), .B(n27400), .Z(n27402) );
  AND U27932 ( .A(n27403), .B(n27402), .Z(n27721) );
  NANDN U27933 ( .A(n27405), .B(n27404), .Z(n27409) );
  NANDN U27934 ( .A(n27407), .B(n27406), .Z(n27408) );
  NAND U27935 ( .A(n27409), .B(n27408), .Z(n27720) );
  XNOR U27936 ( .A(n27721), .B(n27720), .Z(n27722) );
  XNOR U27937 ( .A(n27723), .B(n27722), .Z(n27649) );
  XOR U27938 ( .A(n27650), .B(n27649), .Z(n27652) );
  XOR U27939 ( .A(n27651), .B(n27652), .Z(n27656) );
  NANDN U27940 ( .A(n27411), .B(n27410), .Z(n27415) );
  NANDN U27941 ( .A(n27413), .B(n27412), .Z(n27414) );
  AND U27942 ( .A(n27415), .B(n27414), .Z(n27644) );
  NANDN U27943 ( .A(n27416), .B(n37294), .Z(n27418) );
  XOR U27944 ( .A(b[47]), .B(a[79]), .Z(n27675) );
  NANDN U27945 ( .A(n37172), .B(n27675), .Z(n27417) );
  AND U27946 ( .A(n27418), .B(n27417), .Z(n27716) );
  NANDN U27947 ( .A(n27419), .B(n30627), .Z(n27421) );
  XOR U27948 ( .A(a[117]), .B(b[9]), .Z(n27678) );
  NANDN U27949 ( .A(n30267), .B(n27678), .Z(n27420) );
  AND U27950 ( .A(n27421), .B(n27420), .Z(n27715) );
  NANDN U27951 ( .A(n27422), .B(n37536), .Z(n27424) );
  XOR U27952 ( .A(b[49]), .B(a[77]), .Z(n27681) );
  NANDN U27953 ( .A(n37432), .B(n27681), .Z(n27423) );
  NAND U27954 ( .A(n27424), .B(n27423), .Z(n27714) );
  XOR U27955 ( .A(n27715), .B(n27714), .Z(n27717) );
  XOR U27956 ( .A(n27716), .B(n27717), .Z(n27789) );
  NANDN U27957 ( .A(n36742), .B(n27425), .Z(n27427) );
  XOR U27958 ( .A(b[43]), .B(a[83]), .Z(n27684) );
  NANDN U27959 ( .A(n36891), .B(n27684), .Z(n27426) );
  AND U27960 ( .A(n27427), .B(n27426), .Z(n27695) );
  NANDN U27961 ( .A(n36991), .B(n27428), .Z(n27430) );
  XOR U27962 ( .A(b[45]), .B(a[81]), .Z(n27687) );
  NANDN U27963 ( .A(n37083), .B(n27687), .Z(n27429) );
  AND U27964 ( .A(n27430), .B(n27429), .Z(n27694) );
  NANDN U27965 ( .A(n30482), .B(n27431), .Z(n27433) );
  XOR U27966 ( .A(a[115]), .B(b[11]), .Z(n27690) );
  NANDN U27967 ( .A(n30891), .B(n27690), .Z(n27432) );
  NAND U27968 ( .A(n27433), .B(n27432), .Z(n27693) );
  XOR U27969 ( .A(n27694), .B(n27693), .Z(n27696) );
  XNOR U27970 ( .A(n27695), .B(n27696), .Z(n27788) );
  XNOR U27971 ( .A(n27789), .B(n27788), .Z(n27790) );
  NANDN U27972 ( .A(n27435), .B(n27434), .Z(n27439) );
  OR U27973 ( .A(n27437), .B(n27436), .Z(n27438) );
  NAND U27974 ( .A(n27439), .B(n27438), .Z(n27791) );
  XNOR U27975 ( .A(n27790), .B(n27791), .Z(n27643) );
  XNOR U27976 ( .A(n27644), .B(n27643), .Z(n27645) );
  NANDN U27977 ( .A(n29499), .B(n27440), .Z(n27442) );
  XOR U27978 ( .A(a[119]), .B(b[7]), .Z(n27699) );
  NANDN U27979 ( .A(n29735), .B(n27699), .Z(n27441) );
  AND U27980 ( .A(n27442), .B(n27441), .Z(n27758) );
  NANDN U27981 ( .A(n37857), .B(n27443), .Z(n27445) );
  XOR U27982 ( .A(b[55]), .B(a[71]), .Z(n27702) );
  NANDN U27983 ( .A(n37911), .B(n27702), .Z(n27444) );
  AND U27984 ( .A(n27445), .B(n27444), .Z(n27757) );
  NANDN U27985 ( .A(n35611), .B(n27446), .Z(n27448) );
  XOR U27986 ( .A(b[35]), .B(a[91]), .Z(n27705) );
  NANDN U27987 ( .A(n35801), .B(n27705), .Z(n27447) );
  NAND U27988 ( .A(n27448), .B(n27447), .Z(n27756) );
  XOR U27989 ( .A(n27757), .B(n27756), .Z(n27759) );
  XOR U27990 ( .A(n27758), .B(n27759), .Z(n27769) );
  NANDN U27991 ( .A(n27450), .B(n27449), .Z(n27454) );
  OR U27992 ( .A(n27452), .B(n27451), .Z(n27453) );
  AND U27993 ( .A(n27454), .B(n27453), .Z(n27768) );
  XNOR U27994 ( .A(n27769), .B(n27768), .Z(n27770) );
  NAND U27995 ( .A(n27456), .B(n27455), .Z(n27460) );
  NAND U27996 ( .A(n27458), .B(n27457), .Z(n27459) );
  NAND U27997 ( .A(n27460), .B(n27459), .Z(n27771) );
  XOR U27998 ( .A(n27770), .B(n27771), .Z(n27646) );
  XNOR U27999 ( .A(n27645), .B(n27646), .Z(n27655) );
  XOR U28000 ( .A(n27656), .B(n27655), .Z(n27658) );
  XOR U28001 ( .A(n27657), .B(n27658), .Z(n27626) );
  NANDN U28002 ( .A(n27462), .B(n27461), .Z(n27466) );
  NANDN U28003 ( .A(n27464), .B(n27463), .Z(n27465) );
  AND U28004 ( .A(n27466), .B(n27465), .Z(n27638) );
  NANDN U28005 ( .A(n27468), .B(n27467), .Z(n27472) );
  NAND U28006 ( .A(n27470), .B(n27469), .Z(n27471) );
  AND U28007 ( .A(n27472), .B(n27471), .Z(n27637) );
  XNOR U28008 ( .A(n27638), .B(n27637), .Z(n27640) );
  NANDN U28009 ( .A(n27474), .B(n27473), .Z(n27478) );
  NANDN U28010 ( .A(n27476), .B(n27475), .Z(n27477) );
  NAND U28011 ( .A(n27478), .B(n27477), .Z(n27639) );
  XOR U28012 ( .A(n27640), .B(n27639), .Z(n27664) );
  NANDN U28013 ( .A(n27480), .B(n27479), .Z(n27484) );
  NANDN U28014 ( .A(n27482), .B(n27481), .Z(n27483) );
  AND U28015 ( .A(n27484), .B(n27483), .Z(n27662) );
  NAND U28016 ( .A(n27486), .B(n27485), .Z(n27490) );
  NANDN U28017 ( .A(n27488), .B(n27487), .Z(n27489) );
  AND U28018 ( .A(n27490), .B(n27489), .Z(n27787) );
  NANDN U28019 ( .A(n34223), .B(n27491), .Z(n27493) );
  XOR U28020 ( .A(a[99]), .B(b[27]), .Z(n27800) );
  NANDN U28021 ( .A(n34458), .B(n27800), .Z(n27492) );
  AND U28022 ( .A(n27493), .B(n27492), .Z(n27753) );
  NANDN U28023 ( .A(n34634), .B(n27494), .Z(n27496) );
  XOR U28024 ( .A(a[97]), .B(b[29]), .Z(n27803) );
  NANDN U28025 ( .A(n34722), .B(n27803), .Z(n27495) );
  AND U28026 ( .A(n27496), .B(n27495), .Z(n27751) );
  NANDN U28027 ( .A(n31055), .B(n27497), .Z(n27499) );
  XOR U28028 ( .A(a[113]), .B(b[13]), .Z(n27806) );
  NANDN U28029 ( .A(n31293), .B(n27806), .Z(n27498) );
  NAND U28030 ( .A(n27499), .B(n27498), .Z(n27750) );
  XNOR U28031 ( .A(n27751), .B(n27750), .Z(n27752) );
  XOR U28032 ( .A(n27753), .B(n27752), .Z(n27775) );
  NANDN U28033 ( .A(n28889), .B(n27500), .Z(n27502) );
  XOR U28034 ( .A(a[121]), .B(b[5]), .Z(n27809) );
  NANDN U28035 ( .A(n29138), .B(n27809), .Z(n27501) );
  AND U28036 ( .A(n27502), .B(n27501), .Z(n27853) );
  NANDN U28037 ( .A(n209), .B(n27503), .Z(n27505) );
  XOR U28038 ( .A(a[123]), .B(b[3]), .Z(n27812) );
  NANDN U28039 ( .A(n28941), .B(n27812), .Z(n27504) );
  AND U28040 ( .A(n27505), .B(n27504), .Z(n27852) );
  NANDN U28041 ( .A(n35936), .B(n27506), .Z(n27508) );
  XOR U28042 ( .A(b[37]), .B(a[89]), .Z(n27815) );
  NANDN U28043 ( .A(n36047), .B(n27815), .Z(n27507) );
  NAND U28044 ( .A(n27508), .B(n27507), .Z(n27851) );
  XOR U28045 ( .A(n27852), .B(n27851), .Z(n27854) );
  XNOR U28046 ( .A(n27853), .B(n27854), .Z(n27774) );
  XOR U28047 ( .A(n27775), .B(n27774), .Z(n27777) );
  NANDN U28048 ( .A(n27510), .B(n27509), .Z(n27514) );
  OR U28049 ( .A(n27512), .B(n27511), .Z(n27513) );
  AND U28050 ( .A(n27514), .B(n27513), .Z(n27776) );
  XOR U28051 ( .A(n27777), .B(n27776), .Z(n27785) );
  NANDN U28052 ( .A(n27516), .B(n27515), .Z(n27520) );
  OR U28053 ( .A(n27518), .B(n27517), .Z(n27519) );
  AND U28054 ( .A(n27520), .B(n27519), .Z(n27671) );
  NANDN U28055 ( .A(n32996), .B(n27521), .Z(n27523) );
  XOR U28056 ( .A(a[105]), .B(b[21]), .Z(n27824) );
  NANDN U28057 ( .A(n33271), .B(n27824), .Z(n27522) );
  AND U28058 ( .A(n27523), .B(n27522), .Z(n27860) );
  NANDN U28059 ( .A(n33866), .B(n27524), .Z(n27526) );
  XOR U28060 ( .A(a[103]), .B(b[23]), .Z(n27827) );
  NANDN U28061 ( .A(n33644), .B(n27827), .Z(n27525) );
  AND U28062 ( .A(n27526), .B(n27525), .Z(n27858) );
  NANDN U28063 ( .A(n32483), .B(n27527), .Z(n27529) );
  XOR U28064 ( .A(a[107]), .B(b[19]), .Z(n27830) );
  NANDN U28065 ( .A(n32823), .B(n27830), .Z(n27528) );
  NAND U28066 ( .A(n27529), .B(n27528), .Z(n27857) );
  XNOR U28067 ( .A(n27858), .B(n27857), .Z(n27859) );
  XOR U28068 ( .A(n27860), .B(n27859), .Z(n27670) );
  NANDN U28069 ( .A(n34909), .B(n27530), .Z(n27532) );
  XOR U28070 ( .A(b[31]), .B(a[95]), .Z(n27833) );
  NANDN U28071 ( .A(n35145), .B(n27833), .Z(n27531) );
  AND U28072 ( .A(n27532), .B(n27531), .Z(n27711) );
  NANDN U28073 ( .A(n38247), .B(n27533), .Z(n27535) );
  XOR U28074 ( .A(b[61]), .B(a[65]), .Z(n27836) );
  NANDN U28075 ( .A(n38248), .B(n27836), .Z(n27534) );
  AND U28076 ( .A(n27535), .B(n27534), .Z(n27709) );
  AND U28077 ( .A(b[63]), .B(a[61]), .Z(n27708) );
  XNOR U28078 ( .A(n27709), .B(n27708), .Z(n27710) );
  XOR U28079 ( .A(n27711), .B(n27710), .Z(n27669) );
  XOR U28080 ( .A(n27670), .B(n27669), .Z(n27672) );
  XOR U28081 ( .A(n27671), .B(n27672), .Z(n27784) );
  XOR U28082 ( .A(n27785), .B(n27784), .Z(n27786) );
  XOR U28083 ( .A(n27787), .B(n27786), .Z(n27667) );
  NANDN U28084 ( .A(n27537), .B(n27536), .Z(n27541) );
  NAND U28085 ( .A(n27539), .B(n27538), .Z(n27540) );
  AND U28086 ( .A(n27541), .B(n27540), .Z(n27666) );
  NANDN U28087 ( .A(n27543), .B(n27542), .Z(n27547) );
  NANDN U28088 ( .A(n27545), .B(n27544), .Z(n27546) );
  AND U28089 ( .A(n27547), .B(n27546), .Z(n27781) );
  NANDN U28090 ( .A(n27549), .B(n27548), .Z(n27553) );
  OR U28091 ( .A(n27551), .B(n27550), .Z(n27552) );
  NAND U28092 ( .A(n27553), .B(n27552), .Z(n27780) );
  XNOR U28093 ( .A(n27781), .B(n27780), .Z(n27783) );
  NANDN U28094 ( .A(n27555), .B(n27554), .Z(n27559) );
  OR U28095 ( .A(n27557), .B(n27556), .Z(n27558) );
  NAND U28096 ( .A(n27559), .B(n27558), .Z(n27728) );
  NAND U28097 ( .A(b[0]), .B(a[125]), .Z(n27560) );
  XNOR U28098 ( .A(b[1]), .B(n27560), .Z(n27562) );
  NANDN U28099 ( .A(b[0]), .B(a[124]), .Z(n27561) );
  NAND U28100 ( .A(n27562), .B(n27561), .Z(n27765) );
  NANDN U28101 ( .A(n38278), .B(n27563), .Z(n27565) );
  XOR U28102 ( .A(b[63]), .B(a[63]), .Z(n27863) );
  NANDN U28103 ( .A(n38279), .B(n27863), .Z(n27564) );
  AND U28104 ( .A(n27565), .B(n27564), .Z(n27763) );
  NANDN U28105 ( .A(n35260), .B(n27566), .Z(n27568) );
  XOR U28106 ( .A(b[33]), .B(a[93]), .Z(n27866) );
  NANDN U28107 ( .A(n35456), .B(n27866), .Z(n27567) );
  NAND U28108 ( .A(n27568), .B(n27567), .Z(n27762) );
  XNOR U28109 ( .A(n27763), .B(n27762), .Z(n27764) );
  XNOR U28110 ( .A(n27765), .B(n27764), .Z(n27727) );
  NANDN U28111 ( .A(n37974), .B(n27569), .Z(n27571) );
  XOR U28112 ( .A(b[57]), .B(a[69]), .Z(n27872) );
  NANDN U28113 ( .A(n38031), .B(n27872), .Z(n27570) );
  AND U28114 ( .A(n27571), .B(n27570), .Z(n27847) );
  NANDN U28115 ( .A(n38090), .B(n27572), .Z(n27574) );
  XOR U28116 ( .A(b[59]), .B(a[67]), .Z(n27875) );
  NANDN U28117 ( .A(n38130), .B(n27875), .Z(n27573) );
  AND U28118 ( .A(n27574), .B(n27573), .Z(n27846) );
  NANDN U28119 ( .A(n36480), .B(n27575), .Z(n27577) );
  XOR U28120 ( .A(b[41]), .B(a[85]), .Z(n27878) );
  NANDN U28121 ( .A(n36594), .B(n27878), .Z(n27576) );
  NAND U28122 ( .A(n27577), .B(n27576), .Z(n27845) );
  XOR U28123 ( .A(n27846), .B(n27845), .Z(n27848) );
  XOR U28124 ( .A(n27847), .B(n27848), .Z(n27726) );
  XOR U28125 ( .A(n27727), .B(n27726), .Z(n27729) );
  XOR U28126 ( .A(n27728), .B(n27729), .Z(n27782) );
  XOR U28127 ( .A(n27783), .B(n27782), .Z(n27665) );
  XOR U28128 ( .A(n27666), .B(n27665), .Z(n27668) );
  XOR U28129 ( .A(n27667), .B(n27668), .Z(n27661) );
  XOR U28130 ( .A(n27662), .B(n27661), .Z(n27663) );
  XNOR U28131 ( .A(n27664), .B(n27663), .Z(n27625) );
  XNOR U28132 ( .A(n27626), .B(n27625), .Z(n27627) );
  XOR U28133 ( .A(n27628), .B(n27627), .Z(n27622) );
  XNOR U28134 ( .A(n27621), .B(n27622), .Z(n27616) );
  NANDN U28135 ( .A(n27579), .B(n27578), .Z(n27583) );
  OR U28136 ( .A(n27581), .B(n27580), .Z(n27582) );
  AND U28137 ( .A(n27583), .B(n27582), .Z(n27614) );
  NANDN U28138 ( .A(n27585), .B(n27584), .Z(n27589) );
  NANDN U28139 ( .A(n27587), .B(n27586), .Z(n27588) );
  AND U28140 ( .A(n27589), .B(n27588), .Z(n27613) );
  XNOR U28141 ( .A(n27614), .B(n27613), .Z(n27615) );
  XOR U28142 ( .A(n27616), .B(n27615), .Z(n27882) );
  NANDN U28143 ( .A(n27591), .B(n27590), .Z(n27595) );
  OR U28144 ( .A(n27593), .B(n27592), .Z(n27594) );
  NAND U28145 ( .A(n27595), .B(n27594), .Z(n27881) );
  XNOR U28146 ( .A(n27882), .B(n27881), .Z(n27883) );
  NANDN U28147 ( .A(n27597), .B(n27596), .Z(n27601) );
  NANDN U28148 ( .A(n27599), .B(n27598), .Z(n27600) );
  NAND U28149 ( .A(n27601), .B(n27600), .Z(n27884) );
  XOR U28150 ( .A(n27883), .B(n27884), .Z(n27608) );
  XNOR U28151 ( .A(n27607), .B(n27608), .Z(n27609) );
  XNOR U28152 ( .A(n27610), .B(n27609), .Z(n27887) );
  XNOR U28153 ( .A(sreg[189]), .B(n27887), .Z(n27889) );
  NANDN U28154 ( .A(sreg[188]), .B(n27602), .Z(n27606) );
  NAND U28155 ( .A(n27604), .B(n27603), .Z(n27605) );
  NAND U28156 ( .A(n27606), .B(n27605), .Z(n27888) );
  XNOR U28157 ( .A(n27889), .B(n27888), .Z(c[189]) );
  NANDN U28158 ( .A(n27608), .B(n27607), .Z(n27612) );
  NANDN U28159 ( .A(n27610), .B(n27609), .Z(n27611) );
  AND U28160 ( .A(n27612), .B(n27611), .Z(n27895) );
  NANDN U28161 ( .A(n27614), .B(n27613), .Z(n27618) );
  NAND U28162 ( .A(n27616), .B(n27615), .Z(n27617) );
  AND U28163 ( .A(n27618), .B(n27617), .Z(n28174) );
  NANDN U28164 ( .A(n27620), .B(n27619), .Z(n27624) );
  NANDN U28165 ( .A(n27622), .B(n27621), .Z(n27623) );
  AND U28166 ( .A(n27624), .B(n27623), .Z(n28173) );
  NANDN U28167 ( .A(n27626), .B(n27625), .Z(n27630) );
  NANDN U28168 ( .A(n27628), .B(n27627), .Z(n27629) );
  AND U28169 ( .A(n27630), .B(n27629), .Z(n27899) );
  NANDN U28170 ( .A(n27632), .B(n27631), .Z(n27636) );
  OR U28171 ( .A(n27634), .B(n27633), .Z(n27635) );
  AND U28172 ( .A(n27636), .B(n27635), .Z(n27898) );
  XNOR U28173 ( .A(n27899), .B(n27898), .Z(n27900) );
  NANDN U28174 ( .A(n27638), .B(n27637), .Z(n27642) );
  NAND U28175 ( .A(n27640), .B(n27639), .Z(n27641) );
  AND U28176 ( .A(n27642), .B(n27641), .Z(n28168) );
  NANDN U28177 ( .A(n27644), .B(n27643), .Z(n27648) );
  NANDN U28178 ( .A(n27646), .B(n27645), .Z(n27647) );
  AND U28179 ( .A(n27648), .B(n27647), .Z(n28167) );
  NANDN U28180 ( .A(n27650), .B(n27649), .Z(n27654) );
  OR U28181 ( .A(n27652), .B(n27651), .Z(n27653) );
  AND U28182 ( .A(n27654), .B(n27653), .Z(n28166) );
  XOR U28183 ( .A(n28167), .B(n28166), .Z(n28169) );
  XOR U28184 ( .A(n28168), .B(n28169), .Z(n27905) );
  NANDN U28185 ( .A(n27656), .B(n27655), .Z(n27660) );
  OR U28186 ( .A(n27658), .B(n27657), .Z(n27659) );
  AND U28187 ( .A(n27660), .B(n27659), .Z(n27904) );
  XNOR U28188 ( .A(n27905), .B(n27904), .Z(n27906) );
  NAND U28189 ( .A(n27670), .B(n27669), .Z(n27674) );
  NAND U28190 ( .A(n27672), .B(n27671), .Z(n27673) );
  AND U28191 ( .A(n27674), .B(n27673), .Z(n28145) );
  NANDN U28192 ( .A(n211), .B(n27675), .Z(n27677) );
  XOR U28193 ( .A(b[47]), .B(a[80]), .Z(n27979) );
  NANDN U28194 ( .A(n37172), .B(n27979), .Z(n27676) );
  AND U28195 ( .A(n27677), .B(n27676), .Z(n27975) );
  NANDN U28196 ( .A(n210), .B(n27678), .Z(n27680) );
  XOR U28197 ( .A(a[118]), .B(b[9]), .Z(n27982) );
  NANDN U28198 ( .A(n30267), .B(n27982), .Z(n27679) );
  AND U28199 ( .A(n27680), .B(n27679), .Z(n27974) );
  NANDN U28200 ( .A(n212), .B(n27681), .Z(n27683) );
  XOR U28201 ( .A(b[49]), .B(a[78]), .Z(n27985) );
  NANDN U28202 ( .A(n37432), .B(n27985), .Z(n27682) );
  NAND U28203 ( .A(n27683), .B(n27682), .Z(n27973) );
  XOR U28204 ( .A(n27974), .B(n27973), .Z(n27976) );
  XOR U28205 ( .A(n27975), .B(n27976), .Z(n28082) );
  NANDN U28206 ( .A(n36742), .B(n27684), .Z(n27686) );
  XOR U28207 ( .A(b[43]), .B(a[84]), .Z(n27988) );
  NANDN U28208 ( .A(n36891), .B(n27988), .Z(n27685) );
  AND U28209 ( .A(n27686), .B(n27685), .Z(n27999) );
  NANDN U28210 ( .A(n36991), .B(n27687), .Z(n27689) );
  XOR U28211 ( .A(b[45]), .B(a[82]), .Z(n27991) );
  NANDN U28212 ( .A(n37083), .B(n27991), .Z(n27688) );
  AND U28213 ( .A(n27689), .B(n27688), .Z(n27998) );
  NANDN U28214 ( .A(n30482), .B(n27690), .Z(n27692) );
  XOR U28215 ( .A(a[116]), .B(b[11]), .Z(n27994) );
  NANDN U28216 ( .A(n30891), .B(n27994), .Z(n27691) );
  NAND U28217 ( .A(n27692), .B(n27691), .Z(n27997) );
  XOR U28218 ( .A(n27998), .B(n27997), .Z(n28000) );
  XNOR U28219 ( .A(n27999), .B(n28000), .Z(n28081) );
  XNOR U28220 ( .A(n28082), .B(n28081), .Z(n28083) );
  NANDN U28221 ( .A(n27694), .B(n27693), .Z(n27698) );
  OR U28222 ( .A(n27696), .B(n27695), .Z(n27697) );
  NAND U28223 ( .A(n27698), .B(n27697), .Z(n28084) );
  XNOR U28224 ( .A(n28083), .B(n28084), .Z(n28144) );
  XNOR U28225 ( .A(n28145), .B(n28144), .Z(n28147) );
  NANDN U28226 ( .A(n29499), .B(n27699), .Z(n27701) );
  XOR U28227 ( .A(a[120]), .B(b[7]), .Z(n27958) );
  NANDN U28228 ( .A(n29735), .B(n27958), .Z(n27700) );
  AND U28229 ( .A(n27701), .B(n27700), .Z(n27948) );
  NANDN U28230 ( .A(n37857), .B(n27702), .Z(n27704) );
  XOR U28231 ( .A(b[55]), .B(a[72]), .Z(n27961) );
  NANDN U28232 ( .A(n37911), .B(n27961), .Z(n27703) );
  AND U28233 ( .A(n27704), .B(n27703), .Z(n27947) );
  NANDN U28234 ( .A(n35611), .B(n27705), .Z(n27707) );
  XOR U28235 ( .A(b[35]), .B(a[92]), .Z(n27964) );
  NANDN U28236 ( .A(n35801), .B(n27964), .Z(n27706) );
  NAND U28237 ( .A(n27707), .B(n27706), .Z(n27946) );
  XOR U28238 ( .A(n27947), .B(n27946), .Z(n27949) );
  XOR U28239 ( .A(n27948), .B(n27949), .Z(n28016) );
  NANDN U28240 ( .A(n27709), .B(n27708), .Z(n27713) );
  NANDN U28241 ( .A(n27711), .B(n27710), .Z(n27712) );
  AND U28242 ( .A(n27713), .B(n27712), .Z(n28015) );
  XNOR U28243 ( .A(n28016), .B(n28015), .Z(n28017) );
  NANDN U28244 ( .A(n27715), .B(n27714), .Z(n27719) );
  OR U28245 ( .A(n27717), .B(n27716), .Z(n27718) );
  NAND U28246 ( .A(n27719), .B(n27718), .Z(n28018) );
  XNOR U28247 ( .A(n28017), .B(n28018), .Z(n28146) );
  XOR U28248 ( .A(n28147), .B(n28146), .Z(n28139) );
  NANDN U28249 ( .A(n27721), .B(n27720), .Z(n27725) );
  NANDN U28250 ( .A(n27723), .B(n27722), .Z(n27724) );
  AND U28251 ( .A(n27725), .B(n27724), .Z(n28159) );
  NAND U28252 ( .A(n27727), .B(n27726), .Z(n27731) );
  NAND U28253 ( .A(n27729), .B(n27728), .Z(n27730) );
  AND U28254 ( .A(n27731), .B(n27730), .Z(n28157) );
  NANDN U28255 ( .A(n33875), .B(n27732), .Z(n27734) );
  XOR U28256 ( .A(a[102]), .B(b[25]), .Z(n27922) );
  NANDN U28257 ( .A(n33994), .B(n27922), .Z(n27733) );
  AND U28258 ( .A(n27734), .B(n27733), .Z(n28113) );
  NANDN U28259 ( .A(n32013), .B(n27735), .Z(n27737) );
  XOR U28260 ( .A(a[110]), .B(b[17]), .Z(n27925) );
  NANDN U28261 ( .A(n32292), .B(n27925), .Z(n27736) );
  AND U28262 ( .A(n27737), .B(n27736), .Z(n28112) );
  NANDN U28263 ( .A(n31536), .B(n27738), .Z(n27740) );
  XOR U28264 ( .A(a[112]), .B(b[15]), .Z(n27928) );
  NANDN U28265 ( .A(n31925), .B(n27928), .Z(n27739) );
  NAND U28266 ( .A(n27740), .B(n27739), .Z(n28111) );
  XOR U28267 ( .A(n28112), .B(n28111), .Z(n28114) );
  XOR U28268 ( .A(n28113), .B(n28114), .Z(n28076) );
  NANDN U28269 ( .A(n37526), .B(n27741), .Z(n27743) );
  XOR U28270 ( .A(b[51]), .B(a[76]), .Z(n27931) );
  NANDN U28271 ( .A(n37605), .B(n27931), .Z(n27742) );
  AND U28272 ( .A(n27743), .B(n27742), .Z(n28107) );
  NANDN U28273 ( .A(n37705), .B(n27744), .Z(n27746) );
  XOR U28274 ( .A(b[53]), .B(a[74]), .Z(n27934) );
  NANDN U28275 ( .A(n37778), .B(n27934), .Z(n27745) );
  AND U28276 ( .A(n27746), .B(n27745), .Z(n28106) );
  NANDN U28277 ( .A(n36210), .B(n27747), .Z(n27749) );
  XOR U28278 ( .A(b[39]), .B(a[88]), .Z(n27937) );
  NANDN U28279 ( .A(n36347), .B(n27937), .Z(n27748) );
  NAND U28280 ( .A(n27749), .B(n27748), .Z(n28105) );
  XOR U28281 ( .A(n28106), .B(n28105), .Z(n28108) );
  XNOR U28282 ( .A(n28107), .B(n28108), .Z(n28075) );
  XNOR U28283 ( .A(n28076), .B(n28075), .Z(n28078) );
  NANDN U28284 ( .A(n27751), .B(n27750), .Z(n27755) );
  NANDN U28285 ( .A(n27753), .B(n27752), .Z(n27754) );
  AND U28286 ( .A(n27755), .B(n27754), .Z(n28077) );
  XOR U28287 ( .A(n28078), .B(n28077), .Z(n27913) );
  NANDN U28288 ( .A(n27757), .B(n27756), .Z(n27761) );
  OR U28289 ( .A(n27759), .B(n27758), .Z(n27760) );
  AND U28290 ( .A(n27761), .B(n27760), .Z(n27911) );
  NANDN U28291 ( .A(n27763), .B(n27762), .Z(n27767) );
  NANDN U28292 ( .A(n27765), .B(n27764), .Z(n27766) );
  NAND U28293 ( .A(n27767), .B(n27766), .Z(n27910) );
  XNOR U28294 ( .A(n27911), .B(n27910), .Z(n27912) );
  XNOR U28295 ( .A(n27913), .B(n27912), .Z(n28156) );
  XNOR U28296 ( .A(n28157), .B(n28156), .Z(n28158) );
  XNOR U28297 ( .A(n28159), .B(n28158), .Z(n28138) );
  XNOR U28298 ( .A(n28139), .B(n28138), .Z(n28140) );
  XNOR U28299 ( .A(n28141), .B(n28140), .Z(n28163) );
  NANDN U28300 ( .A(n27769), .B(n27768), .Z(n27773) );
  NANDN U28301 ( .A(n27771), .B(n27770), .Z(n27772) );
  NAND U28302 ( .A(n27773), .B(n27772), .Z(n28152) );
  NAND U28303 ( .A(n27775), .B(n27774), .Z(n27779) );
  NAND U28304 ( .A(n27777), .B(n27776), .Z(n27778) );
  NAND U28305 ( .A(n27779), .B(n27778), .Z(n28150) );
  XOR U28306 ( .A(n28150), .B(n28151), .Z(n28153) );
  XNOR U28307 ( .A(n28152), .B(n28153), .Z(n28135) );
  NANDN U28308 ( .A(n27789), .B(n27788), .Z(n27793) );
  NANDN U28309 ( .A(n27791), .B(n27790), .Z(n27792) );
  AND U28310 ( .A(n27793), .B(n27792), .Z(n28035) );
  NANDN U28311 ( .A(n27795), .B(n27794), .Z(n27799) );
  OR U28312 ( .A(n27797), .B(n27796), .Z(n27798) );
  AND U28313 ( .A(n27799), .B(n27798), .Z(n28023) );
  NANDN U28314 ( .A(n34223), .B(n27800), .Z(n27802) );
  XOR U28315 ( .A(a[100]), .B(b[27]), .Z(n28087) );
  NANDN U28316 ( .A(n34458), .B(n28087), .Z(n27801) );
  AND U28317 ( .A(n27802), .B(n27801), .Z(n27942) );
  NANDN U28318 ( .A(n34634), .B(n27803), .Z(n27805) );
  XOR U28319 ( .A(a[98]), .B(b[29]), .Z(n28090) );
  NANDN U28320 ( .A(n34722), .B(n28090), .Z(n27804) );
  AND U28321 ( .A(n27805), .B(n27804), .Z(n27941) );
  NANDN U28322 ( .A(n31055), .B(n27806), .Z(n27808) );
  XOR U28323 ( .A(a[114]), .B(b[13]), .Z(n28093) );
  NANDN U28324 ( .A(n31293), .B(n28093), .Z(n27807) );
  NAND U28325 ( .A(n27808), .B(n27807), .Z(n27940) );
  XOR U28326 ( .A(n27941), .B(n27940), .Z(n27943) );
  XOR U28327 ( .A(n27942), .B(n27943), .Z(n28022) );
  NANDN U28328 ( .A(n28889), .B(n27809), .Z(n27811) );
  XOR U28329 ( .A(a[122]), .B(b[5]), .Z(n28096) );
  NANDN U28330 ( .A(n29138), .B(n28096), .Z(n27810) );
  AND U28331 ( .A(n27811), .B(n27810), .Z(n28047) );
  NANDN U28332 ( .A(n209), .B(n27812), .Z(n27814) );
  XOR U28333 ( .A(a[124]), .B(b[3]), .Z(n28099) );
  NANDN U28334 ( .A(n28941), .B(n28099), .Z(n27813) );
  AND U28335 ( .A(n27814), .B(n27813), .Z(n28046) );
  NANDN U28336 ( .A(n35936), .B(n27815), .Z(n27817) );
  XOR U28337 ( .A(b[37]), .B(a[90]), .Z(n28102) );
  NANDN U28338 ( .A(n36047), .B(n28102), .Z(n27816) );
  NAND U28339 ( .A(n27817), .B(n27816), .Z(n28045) );
  XOR U28340 ( .A(n28046), .B(n28045), .Z(n28048) );
  XNOR U28341 ( .A(n28047), .B(n28048), .Z(n28021) );
  XOR U28342 ( .A(n28022), .B(n28021), .Z(n28024) );
  XNOR U28343 ( .A(n28023), .B(n28024), .Z(n28033) );
  NANDN U28344 ( .A(n27819), .B(n27818), .Z(n27823) );
  OR U28345 ( .A(n27821), .B(n27820), .Z(n27822) );
  AND U28346 ( .A(n27823), .B(n27822), .Z(n28005) );
  NANDN U28347 ( .A(n32996), .B(n27824), .Z(n27826) );
  XOR U28348 ( .A(a[106]), .B(b[21]), .Z(n28117) );
  NANDN U28349 ( .A(n33271), .B(n28117), .Z(n27825) );
  AND U28350 ( .A(n27826), .B(n27825), .Z(n28053) );
  NANDN U28351 ( .A(n33866), .B(n27827), .Z(n27829) );
  XOR U28352 ( .A(a[104]), .B(b[23]), .Z(n28120) );
  NANDN U28353 ( .A(n33644), .B(n28120), .Z(n27828) );
  AND U28354 ( .A(n27829), .B(n27828), .Z(n28052) );
  NANDN U28355 ( .A(n32483), .B(n27830), .Z(n27832) );
  XOR U28356 ( .A(a[108]), .B(b[19]), .Z(n28123) );
  NANDN U28357 ( .A(n32823), .B(n28123), .Z(n27831) );
  NAND U28358 ( .A(n27832), .B(n27831), .Z(n28051) );
  XOR U28359 ( .A(n28052), .B(n28051), .Z(n28054) );
  XOR U28360 ( .A(n28053), .B(n28054), .Z(n28004) );
  NANDN U28361 ( .A(n34909), .B(n27833), .Z(n27835) );
  XOR U28362 ( .A(b[31]), .B(a[96]), .Z(n28126) );
  NANDN U28363 ( .A(n35145), .B(n28126), .Z(n27834) );
  AND U28364 ( .A(n27835), .B(n27834), .Z(n27969) );
  NANDN U28365 ( .A(n38247), .B(n27836), .Z(n27838) );
  XOR U28366 ( .A(b[61]), .B(a[66]), .Z(n28129) );
  NANDN U28367 ( .A(n38248), .B(n28129), .Z(n27837) );
  AND U28368 ( .A(n27838), .B(n27837), .Z(n27968) );
  AND U28369 ( .A(b[63]), .B(a[62]), .Z(n27967) );
  XOR U28370 ( .A(n27968), .B(n27967), .Z(n27970) );
  XNOR U28371 ( .A(n27969), .B(n27970), .Z(n28003) );
  XOR U28372 ( .A(n28004), .B(n28003), .Z(n28006) );
  XOR U28373 ( .A(n28005), .B(n28006), .Z(n28034) );
  XOR U28374 ( .A(n28033), .B(n28034), .Z(n28036) );
  XOR U28375 ( .A(n28035), .B(n28036), .Z(n28012) );
  NANDN U28376 ( .A(n27840), .B(n27839), .Z(n27844) );
  NAND U28377 ( .A(n27842), .B(n27841), .Z(n27843) );
  AND U28378 ( .A(n27844), .B(n27843), .Z(n28009) );
  NANDN U28379 ( .A(n27846), .B(n27845), .Z(n27850) );
  OR U28380 ( .A(n27848), .B(n27847), .Z(n27849) );
  AND U28381 ( .A(n27850), .B(n27849), .Z(n28028) );
  NANDN U28382 ( .A(n27852), .B(n27851), .Z(n27856) );
  OR U28383 ( .A(n27854), .B(n27853), .Z(n27855) );
  NAND U28384 ( .A(n27856), .B(n27855), .Z(n28027) );
  XNOR U28385 ( .A(n28028), .B(n28027), .Z(n28029) );
  NANDN U28386 ( .A(n27858), .B(n27857), .Z(n27862) );
  NANDN U28387 ( .A(n27860), .B(n27859), .Z(n27861) );
  AND U28388 ( .A(n27862), .B(n27861), .Z(n27919) );
  NANDN U28389 ( .A(n38278), .B(n27863), .Z(n27865) );
  XOR U28390 ( .A(b[63]), .B(a[64]), .Z(n28057) );
  NANDN U28391 ( .A(n38279), .B(n28057), .Z(n27864) );
  AND U28392 ( .A(n27865), .B(n27864), .Z(n27953) );
  NANDN U28393 ( .A(n35260), .B(n27866), .Z(n27868) );
  XOR U28394 ( .A(b[33]), .B(a[94]), .Z(n28060) );
  NANDN U28395 ( .A(n35456), .B(n28060), .Z(n27867) );
  NAND U28396 ( .A(n27868), .B(n27867), .Z(n27952) );
  XNOR U28397 ( .A(n27953), .B(n27952), .Z(n27954) );
  NAND U28398 ( .A(b[0]), .B(a[126]), .Z(n27869) );
  XNOR U28399 ( .A(b[1]), .B(n27869), .Z(n27871) );
  NANDN U28400 ( .A(b[0]), .B(a[125]), .Z(n27870) );
  NAND U28401 ( .A(n27871), .B(n27870), .Z(n27955) );
  XNOR U28402 ( .A(n27954), .B(n27955), .Z(n27916) );
  NANDN U28403 ( .A(n37974), .B(n27872), .Z(n27874) );
  XOR U28404 ( .A(b[57]), .B(a[70]), .Z(n28066) );
  NANDN U28405 ( .A(n38031), .B(n28066), .Z(n27873) );
  AND U28406 ( .A(n27874), .B(n27873), .Z(n28042) );
  NANDN U28407 ( .A(n38090), .B(n27875), .Z(n27877) );
  XOR U28408 ( .A(b[59]), .B(a[68]), .Z(n28069) );
  NANDN U28409 ( .A(n38130), .B(n28069), .Z(n27876) );
  AND U28410 ( .A(n27877), .B(n27876), .Z(n28040) );
  NANDN U28411 ( .A(n36480), .B(n27878), .Z(n27880) );
  XOR U28412 ( .A(b[41]), .B(a[86]), .Z(n28072) );
  NANDN U28413 ( .A(n36594), .B(n28072), .Z(n27879) );
  NAND U28414 ( .A(n27880), .B(n27879), .Z(n28039) );
  XNOR U28415 ( .A(n28040), .B(n28039), .Z(n28041) );
  XOR U28416 ( .A(n28042), .B(n28041), .Z(n27917) );
  XNOR U28417 ( .A(n27916), .B(n27917), .Z(n27918) );
  XOR U28418 ( .A(n27919), .B(n27918), .Z(n28030) );
  XOR U28419 ( .A(n28029), .B(n28030), .Z(n28010) );
  XNOR U28420 ( .A(n28009), .B(n28010), .Z(n28011) );
  XOR U28421 ( .A(n28012), .B(n28011), .Z(n28133) );
  XNOR U28422 ( .A(n28132), .B(n28133), .Z(n28134) );
  XOR U28423 ( .A(n28135), .B(n28134), .Z(n28162) );
  XOR U28424 ( .A(n28163), .B(n28162), .Z(n28164) );
  XOR U28425 ( .A(n28165), .B(n28164), .Z(n27907) );
  XOR U28426 ( .A(n27906), .B(n27907), .Z(n27901) );
  XNOR U28427 ( .A(n27900), .B(n27901), .Z(n28172) );
  XOR U28428 ( .A(n28173), .B(n28172), .Z(n28175) );
  XOR U28429 ( .A(n28174), .B(n28175), .Z(n27893) );
  NANDN U28430 ( .A(n27882), .B(n27881), .Z(n27886) );
  NANDN U28431 ( .A(n27884), .B(n27883), .Z(n27885) );
  NAND U28432 ( .A(n27886), .B(n27885), .Z(n27892) );
  XNOR U28433 ( .A(n27893), .B(n27892), .Z(n27894) );
  XNOR U28434 ( .A(n27895), .B(n27894), .Z(n28178) );
  XNOR U28435 ( .A(sreg[190]), .B(n28178), .Z(n28180) );
  NANDN U28436 ( .A(sreg[189]), .B(n27887), .Z(n27891) );
  NAND U28437 ( .A(n27889), .B(n27888), .Z(n27890) );
  NAND U28438 ( .A(n27891), .B(n27890), .Z(n28179) );
  XNOR U28439 ( .A(n28180), .B(n28179), .Z(c[190]) );
  NANDN U28440 ( .A(n27893), .B(n27892), .Z(n27897) );
  NANDN U28441 ( .A(n27895), .B(n27894), .Z(n27896) );
  AND U28442 ( .A(n27897), .B(n27896), .Z(n28191) );
  NANDN U28443 ( .A(n27899), .B(n27898), .Z(n27903) );
  NANDN U28444 ( .A(n27901), .B(n27900), .Z(n27902) );
  AND U28445 ( .A(n27903), .B(n27902), .Z(n28469) );
  NANDN U28446 ( .A(n27905), .B(n27904), .Z(n27909) );
  NANDN U28447 ( .A(n27907), .B(n27906), .Z(n27908) );
  AND U28448 ( .A(n27909), .B(n27908), .Z(n28468) );
  NANDN U28449 ( .A(n27911), .B(n27910), .Z(n27915) );
  NANDN U28450 ( .A(n27913), .B(n27912), .Z(n27914) );
  AND U28451 ( .A(n27915), .B(n27914), .Z(n28439) );
  NANDN U28452 ( .A(n27917), .B(n27916), .Z(n27921) );
  NANDN U28453 ( .A(n27919), .B(n27918), .Z(n27920) );
  AND U28454 ( .A(n27921), .B(n27920), .Z(n28438) );
  NANDN U28455 ( .A(n33875), .B(n27922), .Z(n27924) );
  XOR U28456 ( .A(a[103]), .B(b[25]), .Z(n28389) );
  NANDN U28457 ( .A(n33994), .B(n28389), .Z(n27923) );
  AND U28458 ( .A(n27924), .B(n27923), .Z(n28301) );
  NANDN U28459 ( .A(n32013), .B(n27925), .Z(n27927) );
  XOR U28460 ( .A(a[111]), .B(b[17]), .Z(n28392) );
  NANDN U28461 ( .A(n32292), .B(n28392), .Z(n27926) );
  AND U28462 ( .A(n27927), .B(n27926), .Z(n28300) );
  NANDN U28463 ( .A(n31536), .B(n27928), .Z(n27930) );
  XOR U28464 ( .A(a[113]), .B(b[15]), .Z(n28395) );
  NANDN U28465 ( .A(n31925), .B(n28395), .Z(n27929) );
  NAND U28466 ( .A(n27930), .B(n27929), .Z(n28299) );
  XOR U28467 ( .A(n28300), .B(n28299), .Z(n28302) );
  XOR U28468 ( .A(n28301), .B(n28302), .Z(n28264) );
  NANDN U28469 ( .A(n37526), .B(n27931), .Z(n27933) );
  XOR U28470 ( .A(b[51]), .B(a[77]), .Z(n28398) );
  NANDN U28471 ( .A(n37605), .B(n28398), .Z(n27932) );
  AND U28472 ( .A(n27933), .B(n27932), .Z(n28295) );
  NANDN U28473 ( .A(n37705), .B(n27934), .Z(n27936) );
  XOR U28474 ( .A(b[53]), .B(a[75]), .Z(n28401) );
  NANDN U28475 ( .A(n37778), .B(n28401), .Z(n27935) );
  AND U28476 ( .A(n27936), .B(n27935), .Z(n28294) );
  NANDN U28477 ( .A(n36210), .B(n27937), .Z(n27939) );
  XOR U28478 ( .A(b[39]), .B(a[89]), .Z(n28404) );
  NANDN U28479 ( .A(n36347), .B(n28404), .Z(n27938) );
  NAND U28480 ( .A(n27939), .B(n27938), .Z(n28293) );
  XOR U28481 ( .A(n28294), .B(n28293), .Z(n28296) );
  XNOR U28482 ( .A(n28295), .B(n28296), .Z(n28263) );
  XNOR U28483 ( .A(n28264), .B(n28263), .Z(n28266) );
  NANDN U28484 ( .A(n27941), .B(n27940), .Z(n27945) );
  OR U28485 ( .A(n27943), .B(n27942), .Z(n27944) );
  AND U28486 ( .A(n27945), .B(n27944), .Z(n28265) );
  XOR U28487 ( .A(n28266), .B(n28265), .Z(n28380) );
  NANDN U28488 ( .A(n27947), .B(n27946), .Z(n27951) );
  OR U28489 ( .A(n27949), .B(n27948), .Z(n27950) );
  AND U28490 ( .A(n27951), .B(n27950), .Z(n28378) );
  NANDN U28491 ( .A(n27953), .B(n27952), .Z(n27957) );
  NANDN U28492 ( .A(n27955), .B(n27954), .Z(n27956) );
  NAND U28493 ( .A(n27957), .B(n27956), .Z(n28377) );
  XNOR U28494 ( .A(n28378), .B(n28377), .Z(n28379) );
  XNOR U28495 ( .A(n28380), .B(n28379), .Z(n28437) );
  XOR U28496 ( .A(n28438), .B(n28437), .Z(n28440) );
  XOR U28497 ( .A(n28439), .B(n28440), .Z(n28432) );
  NANDN U28498 ( .A(n29499), .B(n27958), .Z(n27960) );
  XOR U28499 ( .A(a[121]), .B(b[7]), .Z(n28356) );
  NANDN U28500 ( .A(n29735), .B(n28356), .Z(n27959) );
  AND U28501 ( .A(n27960), .B(n27959), .Z(n28415) );
  NANDN U28502 ( .A(n37857), .B(n27961), .Z(n27963) );
  XOR U28503 ( .A(b[55]), .B(a[73]), .Z(n28359) );
  NANDN U28504 ( .A(n37911), .B(n28359), .Z(n27962) );
  AND U28505 ( .A(n27963), .B(n27962), .Z(n28414) );
  NANDN U28506 ( .A(n35611), .B(n27964), .Z(n27966) );
  XOR U28507 ( .A(b[35]), .B(a[93]), .Z(n28362) );
  NANDN U28508 ( .A(n35801), .B(n28362), .Z(n27965) );
  NAND U28509 ( .A(n27966), .B(n27965), .Z(n28413) );
  XOR U28510 ( .A(n28414), .B(n28413), .Z(n28416) );
  XOR U28511 ( .A(n28415), .B(n28416), .Z(n28207) );
  NANDN U28512 ( .A(n27968), .B(n27967), .Z(n27972) );
  OR U28513 ( .A(n27970), .B(n27969), .Z(n27971) );
  AND U28514 ( .A(n27972), .B(n27971), .Z(n28206) );
  XNOR U28515 ( .A(n28207), .B(n28206), .Z(n28209) );
  NANDN U28516 ( .A(n27974), .B(n27973), .Z(n27978) );
  OR U28517 ( .A(n27976), .B(n27975), .Z(n27977) );
  AND U28518 ( .A(n27978), .B(n27977), .Z(n28208) );
  XOR U28519 ( .A(n28209), .B(n28208), .Z(n28445) );
  NANDN U28520 ( .A(n211), .B(n27979), .Z(n27981) );
  XOR U28521 ( .A(b[47]), .B(a[81]), .Z(n28332) );
  NANDN U28522 ( .A(n37172), .B(n28332), .Z(n27980) );
  AND U28523 ( .A(n27981), .B(n27980), .Z(n28373) );
  NANDN U28524 ( .A(n210), .B(n27982), .Z(n27984) );
  XOR U28525 ( .A(a[119]), .B(b[9]), .Z(n28335) );
  NANDN U28526 ( .A(n30267), .B(n28335), .Z(n27983) );
  AND U28527 ( .A(n27984), .B(n27983), .Z(n28372) );
  NANDN U28528 ( .A(n212), .B(n27985), .Z(n27987) );
  XOR U28529 ( .A(b[49]), .B(a[79]), .Z(n28338) );
  NANDN U28530 ( .A(n37432), .B(n28338), .Z(n27986) );
  NAND U28531 ( .A(n27987), .B(n27986), .Z(n28371) );
  XOR U28532 ( .A(n28372), .B(n28371), .Z(n28374) );
  XOR U28533 ( .A(n28373), .B(n28374), .Z(n28270) );
  NANDN U28534 ( .A(n36742), .B(n27988), .Z(n27990) );
  XOR U28535 ( .A(b[43]), .B(a[85]), .Z(n28341) );
  NANDN U28536 ( .A(n36891), .B(n28341), .Z(n27989) );
  AND U28537 ( .A(n27990), .B(n27989), .Z(n28352) );
  NANDN U28538 ( .A(n36991), .B(n27991), .Z(n27993) );
  XOR U28539 ( .A(b[45]), .B(a[83]), .Z(n28344) );
  NANDN U28540 ( .A(n37083), .B(n28344), .Z(n27992) );
  AND U28541 ( .A(n27993), .B(n27992), .Z(n28351) );
  NANDN U28542 ( .A(n30482), .B(n27994), .Z(n27996) );
  XOR U28543 ( .A(a[117]), .B(b[11]), .Z(n28347) );
  NANDN U28544 ( .A(n30891), .B(n28347), .Z(n27995) );
  NAND U28545 ( .A(n27996), .B(n27995), .Z(n28350) );
  XOR U28546 ( .A(n28351), .B(n28350), .Z(n28353) );
  XNOR U28547 ( .A(n28352), .B(n28353), .Z(n28269) );
  XNOR U28548 ( .A(n28270), .B(n28269), .Z(n28272) );
  NANDN U28549 ( .A(n27998), .B(n27997), .Z(n28002) );
  OR U28550 ( .A(n28000), .B(n27999), .Z(n28001) );
  AND U28551 ( .A(n28002), .B(n28001), .Z(n28271) );
  XOR U28552 ( .A(n28272), .B(n28271), .Z(n28444) );
  NANDN U28553 ( .A(n28004), .B(n28003), .Z(n28008) );
  NANDN U28554 ( .A(n28006), .B(n28005), .Z(n28007) );
  AND U28555 ( .A(n28008), .B(n28007), .Z(n28443) );
  XOR U28556 ( .A(n28444), .B(n28443), .Z(n28446) );
  XNOR U28557 ( .A(n28445), .B(n28446), .Z(n28431) );
  XNOR U28558 ( .A(n28432), .B(n28431), .Z(n28433) );
  NANDN U28559 ( .A(n28010), .B(n28009), .Z(n28014) );
  NANDN U28560 ( .A(n28012), .B(n28011), .Z(n28013) );
  NAND U28561 ( .A(n28014), .B(n28013), .Z(n28434) );
  XNOR U28562 ( .A(n28433), .B(n28434), .Z(n28455) );
  NANDN U28563 ( .A(n28016), .B(n28015), .Z(n28020) );
  NANDN U28564 ( .A(n28018), .B(n28017), .Z(n28019) );
  AND U28565 ( .A(n28020), .B(n28019), .Z(n28452) );
  NANDN U28566 ( .A(n28022), .B(n28021), .Z(n28026) );
  NANDN U28567 ( .A(n28024), .B(n28023), .Z(n28025) );
  AND U28568 ( .A(n28026), .B(n28025), .Z(n28450) );
  NANDN U28569 ( .A(n28028), .B(n28027), .Z(n28032) );
  NANDN U28570 ( .A(n28030), .B(n28029), .Z(n28031) );
  AND U28571 ( .A(n28032), .B(n28031), .Z(n28449) );
  XNOR U28572 ( .A(n28450), .B(n28449), .Z(n28451) );
  XNOR U28573 ( .A(n28452), .B(n28451), .Z(n28427) );
  NANDN U28574 ( .A(n28034), .B(n28033), .Z(n28038) );
  OR U28575 ( .A(n28036), .B(n28035), .Z(n28037) );
  AND U28576 ( .A(n28038), .B(n28037), .Z(n28426) );
  NANDN U28577 ( .A(n28040), .B(n28039), .Z(n28044) );
  NANDN U28578 ( .A(n28042), .B(n28041), .Z(n28043) );
  AND U28579 ( .A(n28044), .B(n28043), .Z(n28219) );
  NANDN U28580 ( .A(n28046), .B(n28045), .Z(n28050) );
  OR U28581 ( .A(n28048), .B(n28047), .Z(n28049) );
  NAND U28582 ( .A(n28050), .B(n28049), .Z(n28218) );
  XNOR U28583 ( .A(n28219), .B(n28218), .Z(n28221) );
  NANDN U28584 ( .A(n28052), .B(n28051), .Z(n28056) );
  OR U28585 ( .A(n28054), .B(n28053), .Z(n28055) );
  AND U28586 ( .A(n28056), .B(n28055), .Z(n28386) );
  NANDN U28587 ( .A(n38278), .B(n28057), .Z(n28059) );
  XOR U28588 ( .A(b[63]), .B(a[65]), .Z(n28248) );
  NANDN U28589 ( .A(n38279), .B(n28248), .Z(n28058) );
  AND U28590 ( .A(n28059), .B(n28058), .Z(n28420) );
  NANDN U28591 ( .A(n35260), .B(n28060), .Z(n28062) );
  XOR U28592 ( .A(b[33]), .B(a[95]), .Z(n28251) );
  NANDN U28593 ( .A(n35456), .B(n28251), .Z(n28061) );
  NAND U28594 ( .A(n28062), .B(n28061), .Z(n28419) );
  XNOR U28595 ( .A(n28420), .B(n28419), .Z(n28421) );
  NAND U28596 ( .A(b[0]), .B(a[127]), .Z(n28063) );
  XNOR U28597 ( .A(b[1]), .B(n28063), .Z(n28065) );
  NANDN U28598 ( .A(b[0]), .B(a[126]), .Z(n28064) );
  NAND U28599 ( .A(n28065), .B(n28064), .Z(n28422) );
  XNOR U28600 ( .A(n28421), .B(n28422), .Z(n28383) );
  NANDN U28601 ( .A(n37974), .B(n28066), .Z(n28068) );
  XOR U28602 ( .A(b[57]), .B(a[71]), .Z(n28254) );
  NANDN U28603 ( .A(n38031), .B(n28254), .Z(n28067) );
  AND U28604 ( .A(n28068), .B(n28067), .Z(n28233) );
  NANDN U28605 ( .A(n38090), .B(n28069), .Z(n28071) );
  XOR U28606 ( .A(b[59]), .B(a[69]), .Z(n28257) );
  NANDN U28607 ( .A(n38130), .B(n28257), .Z(n28070) );
  AND U28608 ( .A(n28071), .B(n28070), .Z(n28231) );
  NANDN U28609 ( .A(n36480), .B(n28072), .Z(n28074) );
  XOR U28610 ( .A(b[41]), .B(a[87]), .Z(n28260) );
  NANDN U28611 ( .A(n36594), .B(n28260), .Z(n28073) );
  NAND U28612 ( .A(n28074), .B(n28073), .Z(n28230) );
  XNOR U28613 ( .A(n28231), .B(n28230), .Z(n28232) );
  XOR U28614 ( .A(n28233), .B(n28232), .Z(n28384) );
  XNOR U28615 ( .A(n28383), .B(n28384), .Z(n28385) );
  XNOR U28616 ( .A(n28386), .B(n28385), .Z(n28220) );
  XOR U28617 ( .A(n28221), .B(n28220), .Z(n28321) );
  NANDN U28618 ( .A(n28076), .B(n28075), .Z(n28080) );
  NAND U28619 ( .A(n28078), .B(n28077), .Z(n28079) );
  NAND U28620 ( .A(n28080), .B(n28079), .Z(n28320) );
  XNOR U28621 ( .A(n28321), .B(n28320), .Z(n28322) );
  NANDN U28622 ( .A(n28082), .B(n28081), .Z(n28086) );
  NANDN U28623 ( .A(n28084), .B(n28083), .Z(n28085) );
  AND U28624 ( .A(n28086), .B(n28085), .Z(n28227) );
  NANDN U28625 ( .A(n34223), .B(n28087), .Z(n28089) );
  XOR U28626 ( .A(a[101]), .B(b[27]), .Z(n28275) );
  NANDN U28627 ( .A(n34458), .B(n28275), .Z(n28088) );
  AND U28628 ( .A(n28089), .B(n28088), .Z(n28409) );
  NANDN U28629 ( .A(n34634), .B(n28090), .Z(n28092) );
  XOR U28630 ( .A(a[99]), .B(b[29]), .Z(n28278) );
  NANDN U28631 ( .A(n34722), .B(n28278), .Z(n28091) );
  AND U28632 ( .A(n28092), .B(n28091), .Z(n28408) );
  NANDN U28633 ( .A(n31055), .B(n28093), .Z(n28095) );
  XOR U28634 ( .A(a[115]), .B(b[13]), .Z(n28281) );
  NANDN U28635 ( .A(n31293), .B(n28281), .Z(n28094) );
  NAND U28636 ( .A(n28095), .B(n28094), .Z(n28407) );
  XOR U28637 ( .A(n28408), .B(n28407), .Z(n28410) );
  XOR U28638 ( .A(n28409), .B(n28410), .Z(n28213) );
  NANDN U28639 ( .A(n28889), .B(n28096), .Z(n28098) );
  XOR U28640 ( .A(a[123]), .B(b[5]), .Z(n28284) );
  NANDN U28641 ( .A(n29138), .B(n28284), .Z(n28097) );
  AND U28642 ( .A(n28098), .B(n28097), .Z(n28238) );
  NANDN U28643 ( .A(n209), .B(n28099), .Z(n28101) );
  XOR U28644 ( .A(a[125]), .B(b[3]), .Z(n28287) );
  NANDN U28645 ( .A(n28941), .B(n28287), .Z(n28100) );
  AND U28646 ( .A(n28101), .B(n28100), .Z(n28237) );
  NANDN U28647 ( .A(n35936), .B(n28102), .Z(n28104) );
  XOR U28648 ( .A(b[37]), .B(a[91]), .Z(n28290) );
  NANDN U28649 ( .A(n36047), .B(n28290), .Z(n28103) );
  NAND U28650 ( .A(n28104), .B(n28103), .Z(n28236) );
  XOR U28651 ( .A(n28237), .B(n28236), .Z(n28239) );
  XNOR U28652 ( .A(n28238), .B(n28239), .Z(n28212) );
  XNOR U28653 ( .A(n28213), .B(n28212), .Z(n28214) );
  NANDN U28654 ( .A(n28106), .B(n28105), .Z(n28110) );
  OR U28655 ( .A(n28108), .B(n28107), .Z(n28109) );
  NAND U28656 ( .A(n28110), .B(n28109), .Z(n28215) );
  XNOR U28657 ( .A(n28214), .B(n28215), .Z(n28224) );
  NANDN U28658 ( .A(n28112), .B(n28111), .Z(n28116) );
  OR U28659 ( .A(n28114), .B(n28113), .Z(n28115) );
  AND U28660 ( .A(n28116), .B(n28115), .Z(n28328) );
  NANDN U28661 ( .A(n32996), .B(n28117), .Z(n28119) );
  XOR U28662 ( .A(a[107]), .B(b[21]), .Z(n28305) );
  NANDN U28663 ( .A(n33271), .B(n28305), .Z(n28118) );
  AND U28664 ( .A(n28119), .B(n28118), .Z(n28244) );
  NANDN U28665 ( .A(n33866), .B(n28120), .Z(n28122) );
  XOR U28666 ( .A(a[105]), .B(b[23]), .Z(n28308) );
  NANDN U28667 ( .A(n33644), .B(n28308), .Z(n28121) );
  AND U28668 ( .A(n28122), .B(n28121), .Z(n28243) );
  NANDN U28669 ( .A(n32483), .B(n28123), .Z(n28125) );
  XOR U28670 ( .A(a[109]), .B(b[19]), .Z(n28311) );
  NANDN U28671 ( .A(n32823), .B(n28311), .Z(n28124) );
  NAND U28672 ( .A(n28125), .B(n28124), .Z(n28242) );
  XOR U28673 ( .A(n28243), .B(n28242), .Z(n28245) );
  XOR U28674 ( .A(n28244), .B(n28245), .Z(n28327) );
  NANDN U28675 ( .A(n34909), .B(n28126), .Z(n28128) );
  XOR U28676 ( .A(b[31]), .B(a[97]), .Z(n28314) );
  NANDN U28677 ( .A(n35145), .B(n28314), .Z(n28127) );
  AND U28678 ( .A(n28128), .B(n28127), .Z(n28367) );
  NANDN U28679 ( .A(n38247), .B(n28129), .Z(n28131) );
  XOR U28680 ( .A(b[61]), .B(a[67]), .Z(n28317) );
  NANDN U28681 ( .A(n38248), .B(n28317), .Z(n28130) );
  AND U28682 ( .A(n28131), .B(n28130), .Z(n28366) );
  AND U28683 ( .A(b[63]), .B(a[63]), .Z(n28365) );
  XOR U28684 ( .A(n28366), .B(n28365), .Z(n28368) );
  XNOR U28685 ( .A(n28367), .B(n28368), .Z(n28326) );
  XOR U28686 ( .A(n28327), .B(n28326), .Z(n28329) );
  XOR U28687 ( .A(n28328), .B(n28329), .Z(n28225) );
  XNOR U28688 ( .A(n28224), .B(n28225), .Z(n28226) );
  XOR U28689 ( .A(n28227), .B(n28226), .Z(n28323) );
  XNOR U28690 ( .A(n28322), .B(n28323), .Z(n28425) );
  XOR U28691 ( .A(n28426), .B(n28425), .Z(n28428) );
  XOR U28692 ( .A(n28427), .B(n28428), .Z(n28456) );
  XNOR U28693 ( .A(n28455), .B(n28456), .Z(n28457) );
  NANDN U28694 ( .A(n28133), .B(n28132), .Z(n28137) );
  NAND U28695 ( .A(n28135), .B(n28134), .Z(n28136) );
  NAND U28696 ( .A(n28137), .B(n28136), .Z(n28458) );
  XNOR U28697 ( .A(n28457), .B(n28458), .Z(n28203) );
  NANDN U28698 ( .A(n28139), .B(n28138), .Z(n28143) );
  NANDN U28699 ( .A(n28141), .B(n28140), .Z(n28142) );
  AND U28700 ( .A(n28143), .B(n28142), .Z(n28200) );
  NANDN U28701 ( .A(n28145), .B(n28144), .Z(n28149) );
  NAND U28702 ( .A(n28147), .B(n28146), .Z(n28148) );
  AND U28703 ( .A(n28149), .B(n28148), .Z(n28464) );
  NAND U28704 ( .A(n28151), .B(n28150), .Z(n28155) );
  NAND U28705 ( .A(n28153), .B(n28152), .Z(n28154) );
  AND U28706 ( .A(n28155), .B(n28154), .Z(n28462) );
  NANDN U28707 ( .A(n28157), .B(n28156), .Z(n28161) );
  NANDN U28708 ( .A(n28159), .B(n28158), .Z(n28160) );
  AND U28709 ( .A(n28161), .B(n28160), .Z(n28461) );
  XNOR U28710 ( .A(n28462), .B(n28461), .Z(n28463) );
  XOR U28711 ( .A(n28464), .B(n28463), .Z(n28201) );
  XNOR U28712 ( .A(n28200), .B(n28201), .Z(n28202) );
  XOR U28713 ( .A(n28203), .B(n28202), .Z(n28197) );
  NANDN U28714 ( .A(n28167), .B(n28166), .Z(n28171) );
  OR U28715 ( .A(n28169), .B(n28168), .Z(n28170) );
  AND U28716 ( .A(n28171), .B(n28170), .Z(n28194) );
  XNOR U28717 ( .A(n28195), .B(n28194), .Z(n28196) );
  XNOR U28718 ( .A(n28197), .B(n28196), .Z(n28467) );
  XOR U28719 ( .A(n28468), .B(n28467), .Z(n28470) );
  XOR U28720 ( .A(n28469), .B(n28470), .Z(n28189) );
  NANDN U28721 ( .A(n28173), .B(n28172), .Z(n28177) );
  OR U28722 ( .A(n28175), .B(n28174), .Z(n28176) );
  AND U28723 ( .A(n28177), .B(n28176), .Z(n28188) );
  XNOR U28724 ( .A(n28189), .B(n28188), .Z(n28190) );
  XNOR U28725 ( .A(n28191), .B(n28190), .Z(n28183) );
  XNOR U28726 ( .A(sreg[191]), .B(n28183), .Z(n28185) );
  NANDN U28727 ( .A(sreg[190]), .B(n28178), .Z(n28182) );
  NAND U28728 ( .A(n28180), .B(n28179), .Z(n28181) );
  NAND U28729 ( .A(n28182), .B(n28181), .Z(n28184) );
  XNOR U28730 ( .A(n28185), .B(n28184), .Z(c[191]) );
  NANDN U28731 ( .A(sreg[191]), .B(n28183), .Z(n28187) );
  NAND U28732 ( .A(n28185), .B(n28184), .Z(n28186) );
  AND U28733 ( .A(n28187), .B(n28186), .Z(n28474) );
  NANDN U28734 ( .A(n28189), .B(n28188), .Z(n28193) );
  NANDN U28735 ( .A(n28191), .B(n28190), .Z(n28192) );
  AND U28736 ( .A(n28193), .B(n28192), .Z(n28477) );
  NANDN U28737 ( .A(n28195), .B(n28194), .Z(n28199) );
  NANDN U28738 ( .A(n28197), .B(n28196), .Z(n28198) );
  AND U28739 ( .A(n28199), .B(n28198), .Z(n28483) );
  NANDN U28740 ( .A(n28201), .B(n28200), .Z(n28205) );
  NAND U28741 ( .A(n28203), .B(n28202), .Z(n28204) );
  AND U28742 ( .A(n28205), .B(n28204), .Z(n28481) );
  NANDN U28743 ( .A(n28207), .B(n28206), .Z(n28211) );
  NAND U28744 ( .A(n28209), .B(n28208), .Z(n28210) );
  AND U28745 ( .A(n28211), .B(n28210), .Z(n28502) );
  NANDN U28746 ( .A(n28213), .B(n28212), .Z(n28217) );
  NANDN U28747 ( .A(n28215), .B(n28214), .Z(n28216) );
  AND U28748 ( .A(n28217), .B(n28216), .Z(n28500) );
  NANDN U28749 ( .A(n28219), .B(n28218), .Z(n28223) );
  NAND U28750 ( .A(n28221), .B(n28220), .Z(n28222) );
  AND U28751 ( .A(n28223), .B(n28222), .Z(n28499) );
  XNOR U28752 ( .A(n28500), .B(n28499), .Z(n28501) );
  XNOR U28753 ( .A(n28502), .B(n28501), .Z(n28526) );
  NANDN U28754 ( .A(n28225), .B(n28224), .Z(n28229) );
  NANDN U28755 ( .A(n28227), .B(n28226), .Z(n28228) );
  AND U28756 ( .A(n28229), .B(n28228), .Z(n28524) );
  NANDN U28757 ( .A(n28231), .B(n28230), .Z(n28235) );
  NANDN U28758 ( .A(n28233), .B(n28232), .Z(n28234) );
  AND U28759 ( .A(n28235), .B(n28234), .Z(n28647) );
  NANDN U28760 ( .A(n28237), .B(n28236), .Z(n28241) );
  OR U28761 ( .A(n28239), .B(n28238), .Z(n28240) );
  NAND U28762 ( .A(n28241), .B(n28240), .Z(n28646) );
  XNOR U28763 ( .A(n28647), .B(n28646), .Z(n28649) );
  NANDN U28764 ( .A(n28243), .B(n28242), .Z(n28247) );
  OR U28765 ( .A(n28245), .B(n28244), .Z(n28246) );
  NAND U28766 ( .A(n28247), .B(n28246), .Z(n28543) );
  NANDN U28767 ( .A(n38278), .B(n28248), .Z(n28250) );
  XOR U28768 ( .A(b[63]), .B(a[66]), .Z(n28725) );
  NANDN U28769 ( .A(n38279), .B(n28725), .Z(n28249) );
  AND U28770 ( .A(n28250), .B(n28249), .Z(n28572) );
  NANDN U28771 ( .A(n35260), .B(n28251), .Z(n28253) );
  XOR U28772 ( .A(b[33]), .B(a[96]), .Z(n28728) );
  NANDN U28773 ( .A(n35456), .B(n28728), .Z(n28252) );
  NAND U28774 ( .A(n28253), .B(n28252), .Z(n28571) );
  XNOR U28775 ( .A(n28572), .B(n28571), .Z(n28573) );
  XNOR U28776 ( .A(n28574), .B(n28573), .Z(n28542) );
  NANDN U28777 ( .A(n37974), .B(n28254), .Z(n28256) );
  XOR U28778 ( .A(b[57]), .B(a[72]), .Z(n28713) );
  NANDN U28779 ( .A(n38031), .B(n28713), .Z(n28255) );
  AND U28780 ( .A(n28256), .B(n28255), .Z(n28733) );
  NANDN U28781 ( .A(n38090), .B(n28257), .Z(n28259) );
  XOR U28782 ( .A(b[59]), .B(a[70]), .Z(n28716) );
  NANDN U28783 ( .A(n38130), .B(n28716), .Z(n28258) );
  AND U28784 ( .A(n28259), .B(n28258), .Z(n28732) );
  NANDN U28785 ( .A(n36480), .B(n28260), .Z(n28262) );
  XOR U28786 ( .A(b[41]), .B(a[88]), .Z(n28719) );
  NANDN U28787 ( .A(n36594), .B(n28719), .Z(n28261) );
  NAND U28788 ( .A(n28262), .B(n28261), .Z(n28731) );
  XOR U28789 ( .A(n28732), .B(n28731), .Z(n28734) );
  XOR U28790 ( .A(n28733), .B(n28734), .Z(n28541) );
  XOR U28791 ( .A(n28542), .B(n28541), .Z(n28544) );
  XOR U28792 ( .A(n28543), .B(n28544), .Z(n28648) );
  XOR U28793 ( .A(n28649), .B(n28648), .Z(n28530) );
  NANDN U28794 ( .A(n28264), .B(n28263), .Z(n28268) );
  NAND U28795 ( .A(n28266), .B(n28265), .Z(n28267) );
  NAND U28796 ( .A(n28268), .B(n28267), .Z(n28529) );
  XNOR U28797 ( .A(n28530), .B(n28529), .Z(n28531) );
  NANDN U28798 ( .A(n28270), .B(n28269), .Z(n28274) );
  NAND U28799 ( .A(n28272), .B(n28271), .Z(n28273) );
  AND U28800 ( .A(n28274), .B(n28273), .Z(n28746) );
  NANDN U28801 ( .A(n34223), .B(n28275), .Z(n28277) );
  XOR U28802 ( .A(a[102]), .B(b[27]), .Z(n28547) );
  NANDN U28803 ( .A(n34458), .B(n28547), .Z(n28276) );
  AND U28804 ( .A(n28277), .B(n28276), .Z(n28567) );
  NANDN U28805 ( .A(n34634), .B(n28278), .Z(n28280) );
  XOR U28806 ( .A(a[100]), .B(b[29]), .Z(n28677) );
  NANDN U28807 ( .A(n34722), .B(n28677), .Z(n28279) );
  AND U28808 ( .A(n28280), .B(n28279), .Z(n28566) );
  NANDN U28809 ( .A(n31055), .B(n28281), .Z(n28283) );
  XOR U28810 ( .A(a[116]), .B(b[13]), .Z(n28604) );
  NANDN U28811 ( .A(n31293), .B(n28604), .Z(n28282) );
  NAND U28812 ( .A(n28283), .B(n28282), .Z(n28565) );
  XOR U28813 ( .A(n28566), .B(n28565), .Z(n28568) );
  XOR U28814 ( .A(n28567), .B(n28568), .Z(n28641) );
  NANDN U28815 ( .A(n28889), .B(n28284), .Z(n28286) );
  XOR U28816 ( .A(a[124]), .B(b[5]), .Z(n28689) );
  NANDN U28817 ( .A(n29138), .B(n28689), .Z(n28285) );
  AND U28818 ( .A(n28286), .B(n28285), .Z(n28739) );
  NANDN U28819 ( .A(n209), .B(n28287), .Z(n28289) );
  XOR U28820 ( .A(a[126]), .B(b[3]), .Z(n28722) );
  NANDN U28821 ( .A(n28941), .B(n28722), .Z(n28288) );
  AND U28822 ( .A(n28289), .B(n28288), .Z(n28738) );
  NANDN U28823 ( .A(n35936), .B(n28290), .Z(n28292) );
  XOR U28824 ( .A(b[37]), .B(a[92]), .Z(n28692) );
  NANDN U28825 ( .A(n36047), .B(n28692), .Z(n28291) );
  NAND U28826 ( .A(n28292), .B(n28291), .Z(n28737) );
  XOR U28827 ( .A(n28738), .B(n28737), .Z(n28740) );
  XNOR U28828 ( .A(n28739), .B(n28740), .Z(n28640) );
  XNOR U28829 ( .A(n28641), .B(n28640), .Z(n28642) );
  NANDN U28830 ( .A(n28294), .B(n28293), .Z(n28298) );
  OR U28831 ( .A(n28296), .B(n28295), .Z(n28297) );
  NAND U28832 ( .A(n28298), .B(n28297), .Z(n28643) );
  XNOR U28833 ( .A(n28642), .B(n28643), .Z(n28743) );
  NANDN U28834 ( .A(n28300), .B(n28299), .Z(n28304) );
  OR U28835 ( .A(n28302), .B(n28301), .Z(n28303) );
  AND U28836 ( .A(n28304), .B(n28303), .Z(n28585) );
  NANDN U28837 ( .A(n32996), .B(n28305), .Z(n28307) );
  XOR U28838 ( .A(a[108]), .B(b[21]), .Z(n28664) );
  NANDN U28839 ( .A(n33271), .B(n28664), .Z(n28306) );
  AND U28840 ( .A(n28307), .B(n28306), .Z(n28709) );
  NANDN U28841 ( .A(n33866), .B(n28308), .Z(n28310) );
  XOR U28842 ( .A(a[106]), .B(b[23]), .Z(n28658) );
  NANDN U28843 ( .A(n33644), .B(n28658), .Z(n28309) );
  AND U28844 ( .A(n28310), .B(n28309), .Z(n28708) );
  NANDN U28845 ( .A(n32483), .B(n28311), .Z(n28313) );
  XOR U28846 ( .A(a[110]), .B(b[19]), .Z(n28550) );
  NANDN U28847 ( .A(n32823), .B(n28550), .Z(n28312) );
  NAND U28848 ( .A(n28313), .B(n28312), .Z(n28707) );
  XOR U28849 ( .A(n28708), .B(n28707), .Z(n28710) );
  XOR U28850 ( .A(n28709), .B(n28710), .Z(n28584) );
  NANDN U28851 ( .A(n34909), .B(n28314), .Z(n28316) );
  XOR U28852 ( .A(a[98]), .B(b[31]), .Z(n28680) );
  NANDN U28853 ( .A(n35145), .B(n28680), .Z(n28315) );
  AND U28854 ( .A(n28316), .B(n28315), .Z(n28624) );
  NANDN U28855 ( .A(n38247), .B(n28317), .Z(n28319) );
  XOR U28856 ( .A(b[61]), .B(a[68]), .Z(n28667) );
  NANDN U28857 ( .A(n38248), .B(n28667), .Z(n28318) );
  AND U28858 ( .A(n28319), .B(n28318), .Z(n28623) );
  AND U28859 ( .A(b[63]), .B(a[64]), .Z(n28622) );
  XOR U28860 ( .A(n28623), .B(n28622), .Z(n28625) );
  XNOR U28861 ( .A(n28624), .B(n28625), .Z(n28583) );
  XOR U28862 ( .A(n28584), .B(n28583), .Z(n28586) );
  XOR U28863 ( .A(n28585), .B(n28586), .Z(n28744) );
  XNOR U28864 ( .A(n28743), .B(n28744), .Z(n28745) );
  XOR U28865 ( .A(n28746), .B(n28745), .Z(n28532) );
  XNOR U28866 ( .A(n28531), .B(n28532), .Z(n28523) );
  XNOR U28867 ( .A(n28524), .B(n28523), .Z(n28525) );
  XOR U28868 ( .A(n28526), .B(n28525), .Z(n28494) );
  NANDN U28869 ( .A(n28321), .B(n28320), .Z(n28325) );
  NANDN U28870 ( .A(n28323), .B(n28322), .Z(n28324) );
  AND U28871 ( .A(n28325), .B(n28324), .Z(n28519) );
  NANDN U28872 ( .A(n28327), .B(n28326), .Z(n28331) );
  NANDN U28873 ( .A(n28329), .B(n28328), .Z(n28330) );
  AND U28874 ( .A(n28331), .B(n28330), .Z(n28506) );
  NANDN U28875 ( .A(n211), .B(n28332), .Z(n28334) );
  XOR U28876 ( .A(b[47]), .B(a[82]), .Z(n28589) );
  NANDN U28877 ( .A(n37172), .B(n28589), .Z(n28333) );
  AND U28878 ( .A(n28334), .B(n28333), .Z(n28630) );
  NANDN U28879 ( .A(n210), .B(n28335), .Z(n28337) );
  XOR U28880 ( .A(a[120]), .B(b[9]), .Z(n28613) );
  NANDN U28881 ( .A(n30267), .B(n28613), .Z(n28336) );
  AND U28882 ( .A(n28337), .B(n28336), .Z(n28629) );
  NANDN U28883 ( .A(n212), .B(n28338), .Z(n28340) );
  XOR U28884 ( .A(b[49]), .B(a[80]), .Z(n28595) );
  NANDN U28885 ( .A(n37432), .B(n28595), .Z(n28339) );
  NAND U28886 ( .A(n28340), .B(n28339), .Z(n28628) );
  XOR U28887 ( .A(n28629), .B(n28628), .Z(n28631) );
  XOR U28888 ( .A(n28630), .B(n28631), .Z(n28653) );
  NANDN U28889 ( .A(n36742), .B(n28341), .Z(n28343) );
  XOR U28890 ( .A(b[43]), .B(a[86]), .Z(n28598) );
  NANDN U28891 ( .A(n36891), .B(n28598), .Z(n28342) );
  AND U28892 ( .A(n28343), .B(n28342), .Z(n28609) );
  NANDN U28893 ( .A(n36991), .B(n28344), .Z(n28346) );
  XOR U28894 ( .A(b[45]), .B(a[84]), .Z(n28601) );
  NANDN U28895 ( .A(n37083), .B(n28601), .Z(n28345) );
  AND U28896 ( .A(n28346), .B(n28345), .Z(n28608) );
  NANDN U28897 ( .A(n30482), .B(n28347), .Z(n28349) );
  XOR U28898 ( .A(a[118]), .B(b[11]), .Z(n28592) );
  NANDN U28899 ( .A(n30891), .B(n28592), .Z(n28348) );
  NAND U28900 ( .A(n28349), .B(n28348), .Z(n28607) );
  XOR U28901 ( .A(n28608), .B(n28607), .Z(n28610) );
  XNOR U28902 ( .A(n28609), .B(n28610), .Z(n28652) );
  XNOR U28903 ( .A(n28653), .B(n28652), .Z(n28654) );
  NANDN U28904 ( .A(n28351), .B(n28350), .Z(n28355) );
  OR U28905 ( .A(n28353), .B(n28352), .Z(n28354) );
  NAND U28906 ( .A(n28355), .B(n28354), .Z(n28655) );
  XNOR U28907 ( .A(n28654), .B(n28655), .Z(n28505) );
  XNOR U28908 ( .A(n28506), .B(n28505), .Z(n28508) );
  NANDN U28909 ( .A(n29499), .B(n28356), .Z(n28358) );
  XOR U28910 ( .A(a[122]), .B(b[7]), .Z(n28686) );
  NANDN U28911 ( .A(n29735), .B(n28686), .Z(n28357) );
  AND U28912 ( .A(n28358), .B(n28357), .Z(n28579) );
  NANDN U28913 ( .A(n37857), .B(n28359), .Z(n28361) );
  XOR U28914 ( .A(b[55]), .B(a[74]), .Z(n28616) );
  NANDN U28915 ( .A(n37911), .B(n28616), .Z(n28360) );
  AND U28916 ( .A(n28361), .B(n28360), .Z(n28578) );
  NANDN U28917 ( .A(n35611), .B(n28362), .Z(n28364) );
  XOR U28918 ( .A(b[35]), .B(a[94]), .Z(n28619) );
  NANDN U28919 ( .A(n35801), .B(n28619), .Z(n28363) );
  NAND U28920 ( .A(n28364), .B(n28363), .Z(n28577) );
  XOR U28921 ( .A(n28578), .B(n28577), .Z(n28580) );
  XOR U28922 ( .A(n28579), .B(n28580), .Z(n28635) );
  NANDN U28923 ( .A(n28366), .B(n28365), .Z(n28370) );
  OR U28924 ( .A(n28368), .B(n28367), .Z(n28369) );
  AND U28925 ( .A(n28370), .B(n28369), .Z(n28634) );
  XNOR U28926 ( .A(n28635), .B(n28634), .Z(n28636) );
  NANDN U28927 ( .A(n28372), .B(n28371), .Z(n28376) );
  OR U28928 ( .A(n28374), .B(n28373), .Z(n28375) );
  NAND U28929 ( .A(n28376), .B(n28375), .Z(n28637) );
  XNOR U28930 ( .A(n28636), .B(n28637), .Z(n28507) );
  XOR U28931 ( .A(n28508), .B(n28507), .Z(n28518) );
  NANDN U28932 ( .A(n28378), .B(n28377), .Z(n28382) );
  NANDN U28933 ( .A(n28380), .B(n28379), .Z(n28381) );
  AND U28934 ( .A(n28382), .B(n28381), .Z(n28514) );
  NANDN U28935 ( .A(n28384), .B(n28383), .Z(n28388) );
  NANDN U28936 ( .A(n28386), .B(n28385), .Z(n28387) );
  AND U28937 ( .A(n28388), .B(n28387), .Z(n28512) );
  NANDN U28938 ( .A(n33875), .B(n28389), .Z(n28391) );
  XOR U28939 ( .A(a[104]), .B(b[25]), .Z(n28661) );
  NANDN U28940 ( .A(n33994), .B(n28661), .Z(n28390) );
  AND U28941 ( .A(n28391), .B(n28390), .Z(n28673) );
  NANDN U28942 ( .A(n32013), .B(n28392), .Z(n28394) );
  XOR U28943 ( .A(a[112]), .B(b[17]), .Z(n28553) );
  NANDN U28944 ( .A(n32292), .B(n28553), .Z(n28393) );
  AND U28945 ( .A(n28394), .B(n28393), .Z(n28672) );
  NANDN U28946 ( .A(n31536), .B(n28395), .Z(n28397) );
  XOR U28947 ( .A(a[114]), .B(b[15]), .Z(n28683) );
  NANDN U28948 ( .A(n31925), .B(n28683), .Z(n28396) );
  NAND U28949 ( .A(n28397), .B(n28396), .Z(n28671) );
  XOR U28950 ( .A(n28672), .B(n28671), .Z(n28674) );
  XOR U28951 ( .A(n28673), .B(n28674), .Z(n28702) );
  NANDN U28952 ( .A(n37526), .B(n28398), .Z(n28400) );
  XOR U28953 ( .A(b[51]), .B(a[78]), .Z(n28556) );
  NANDN U28954 ( .A(n37605), .B(n28556), .Z(n28399) );
  AND U28955 ( .A(n28400), .B(n28399), .Z(n28697) );
  NANDN U28956 ( .A(n37705), .B(n28401), .Z(n28403) );
  XOR U28957 ( .A(b[53]), .B(a[76]), .Z(n28559) );
  NANDN U28958 ( .A(n37778), .B(n28559), .Z(n28402) );
  AND U28959 ( .A(n28403), .B(n28402), .Z(n28696) );
  NANDN U28960 ( .A(n36210), .B(n28404), .Z(n28406) );
  XOR U28961 ( .A(b[39]), .B(a[90]), .Z(n28562) );
  NANDN U28962 ( .A(n36347), .B(n28562), .Z(n28405) );
  NAND U28963 ( .A(n28406), .B(n28405), .Z(n28695) );
  XOR U28964 ( .A(n28696), .B(n28695), .Z(n28698) );
  XNOR U28965 ( .A(n28697), .B(n28698), .Z(n28701) );
  XNOR U28966 ( .A(n28702), .B(n28701), .Z(n28704) );
  NANDN U28967 ( .A(n28408), .B(n28407), .Z(n28412) );
  OR U28968 ( .A(n28410), .B(n28409), .Z(n28411) );
  AND U28969 ( .A(n28412), .B(n28411), .Z(n28703) );
  XOR U28970 ( .A(n28704), .B(n28703), .Z(n28538) );
  NANDN U28971 ( .A(n28414), .B(n28413), .Z(n28418) );
  OR U28972 ( .A(n28416), .B(n28415), .Z(n28417) );
  AND U28973 ( .A(n28418), .B(n28417), .Z(n28536) );
  NANDN U28974 ( .A(n28420), .B(n28419), .Z(n28424) );
  NANDN U28975 ( .A(n28422), .B(n28421), .Z(n28423) );
  NAND U28976 ( .A(n28424), .B(n28423), .Z(n28535) );
  XNOR U28977 ( .A(n28536), .B(n28535), .Z(n28537) );
  XNOR U28978 ( .A(n28538), .B(n28537), .Z(n28511) );
  XNOR U28979 ( .A(n28512), .B(n28511), .Z(n28513) );
  XNOR U28980 ( .A(n28514), .B(n28513), .Z(n28517) );
  XOR U28981 ( .A(n28518), .B(n28517), .Z(n28520) );
  XNOR U28982 ( .A(n28519), .B(n28520), .Z(n28493) );
  XNOR U28983 ( .A(n28494), .B(n28493), .Z(n28496) );
  NANDN U28984 ( .A(n28426), .B(n28425), .Z(n28430) );
  NANDN U28985 ( .A(n28428), .B(n28427), .Z(n28429) );
  AND U28986 ( .A(n28430), .B(n28429), .Z(n28495) );
  XOR U28987 ( .A(n28496), .B(n28495), .Z(n28751) );
  NANDN U28988 ( .A(n28432), .B(n28431), .Z(n28436) );
  NANDN U28989 ( .A(n28434), .B(n28433), .Z(n28435) );
  AND U28990 ( .A(n28436), .B(n28435), .Z(n28750) );
  NANDN U28991 ( .A(n28438), .B(n28437), .Z(n28442) );
  OR U28992 ( .A(n28440), .B(n28439), .Z(n28441) );
  AND U28993 ( .A(n28442), .B(n28441), .Z(n28488) );
  NANDN U28994 ( .A(n28444), .B(n28443), .Z(n28448) );
  OR U28995 ( .A(n28446), .B(n28445), .Z(n28447) );
  NAND U28996 ( .A(n28448), .B(n28447), .Z(n28487) );
  XNOR U28997 ( .A(n28488), .B(n28487), .Z(n28490) );
  NANDN U28998 ( .A(n28450), .B(n28449), .Z(n28454) );
  NANDN U28999 ( .A(n28452), .B(n28451), .Z(n28453) );
  AND U29000 ( .A(n28454), .B(n28453), .Z(n28489) );
  XNOR U29001 ( .A(n28490), .B(n28489), .Z(n28749) );
  XOR U29002 ( .A(n28750), .B(n28749), .Z(n28752) );
  XOR U29003 ( .A(n28751), .B(n28752), .Z(n28758) );
  NANDN U29004 ( .A(n28456), .B(n28455), .Z(n28460) );
  NANDN U29005 ( .A(n28458), .B(n28457), .Z(n28459) );
  AND U29006 ( .A(n28460), .B(n28459), .Z(n28755) );
  NANDN U29007 ( .A(n28462), .B(n28461), .Z(n28466) );
  NANDN U29008 ( .A(n28464), .B(n28463), .Z(n28465) );
  NAND U29009 ( .A(n28466), .B(n28465), .Z(n28756) );
  XNOR U29010 ( .A(n28755), .B(n28756), .Z(n28757) );
  XOR U29011 ( .A(n28758), .B(n28757), .Z(n28482) );
  XOR U29012 ( .A(n28481), .B(n28482), .Z(n28484) );
  XOR U29013 ( .A(n28483), .B(n28484), .Z(n28476) );
  NANDN U29014 ( .A(n28468), .B(n28467), .Z(n28472) );
  OR U29015 ( .A(n28470), .B(n28469), .Z(n28471) );
  AND U29016 ( .A(n28472), .B(n28471), .Z(n28475) );
  XOR U29017 ( .A(n28476), .B(n28475), .Z(n28478) );
  XNOR U29018 ( .A(n28477), .B(n28478), .Z(n28473) );
  XOR U29019 ( .A(n28474), .B(n28473), .Z(c[192]) );
  AND U29020 ( .A(n28474), .B(n28473), .Z(n28762) );
  NANDN U29021 ( .A(n28476), .B(n28475), .Z(n28480) );
  OR U29022 ( .A(n28478), .B(n28477), .Z(n28479) );
  AND U29023 ( .A(n28480), .B(n28479), .Z(n28765) );
  NANDN U29024 ( .A(n28482), .B(n28481), .Z(n28486) );
  OR U29025 ( .A(n28484), .B(n28483), .Z(n28485) );
  AND U29026 ( .A(n28486), .B(n28485), .Z(n28763) );
  NANDN U29027 ( .A(n28488), .B(n28487), .Z(n28492) );
  NAND U29028 ( .A(n28490), .B(n28489), .Z(n28491) );
  AND U29029 ( .A(n28492), .B(n28491), .Z(n28776) );
  NANDN U29030 ( .A(n28494), .B(n28493), .Z(n28498) );
  NAND U29031 ( .A(n28496), .B(n28495), .Z(n28497) );
  NAND U29032 ( .A(n28498), .B(n28497), .Z(n28775) );
  XNOR U29033 ( .A(n28776), .B(n28775), .Z(n28778) );
  NANDN U29034 ( .A(n28500), .B(n28499), .Z(n28504) );
  NANDN U29035 ( .A(n28502), .B(n28501), .Z(n28503) );
  AND U29036 ( .A(n28504), .B(n28503), .Z(n28789) );
  NANDN U29037 ( .A(n28506), .B(n28505), .Z(n28510) );
  NAND U29038 ( .A(n28508), .B(n28507), .Z(n28509) );
  AND U29039 ( .A(n28510), .B(n28509), .Z(n28788) );
  NANDN U29040 ( .A(n28512), .B(n28511), .Z(n28516) );
  NANDN U29041 ( .A(n28514), .B(n28513), .Z(n28515) );
  AND U29042 ( .A(n28516), .B(n28515), .Z(n28787) );
  XOR U29043 ( .A(n28788), .B(n28787), .Z(n28790) );
  XOR U29044 ( .A(n28789), .B(n28790), .Z(n29038) );
  NANDN U29045 ( .A(n28518), .B(n28517), .Z(n28522) );
  NANDN U29046 ( .A(n28520), .B(n28519), .Z(n28521) );
  NAND U29047 ( .A(n28522), .B(n28521), .Z(n29037) );
  XNOR U29048 ( .A(n29038), .B(n29037), .Z(n29039) );
  NANDN U29049 ( .A(n28524), .B(n28523), .Z(n28528) );
  NAND U29050 ( .A(n28526), .B(n28525), .Z(n28527) );
  AND U29051 ( .A(n28528), .B(n28527), .Z(n28783) );
  NANDN U29052 ( .A(n28530), .B(n28529), .Z(n28534) );
  NANDN U29053 ( .A(n28532), .B(n28531), .Z(n28533) );
  AND U29054 ( .A(n28534), .B(n28533), .Z(n28872) );
  NANDN U29055 ( .A(n28536), .B(n28535), .Z(n28540) );
  NANDN U29056 ( .A(n28538), .B(n28537), .Z(n28539) );
  AND U29057 ( .A(n28540), .B(n28539), .Z(n29027) );
  NAND U29058 ( .A(n28542), .B(n28541), .Z(n28546) );
  NAND U29059 ( .A(n28544), .B(n28543), .Z(n28545) );
  AND U29060 ( .A(n28546), .B(n28545), .Z(n29026) );
  NANDN U29061 ( .A(n34223), .B(n28547), .Z(n28549) );
  XOR U29062 ( .A(a[103]), .B(b[27]), .Z(n28895) );
  NANDN U29063 ( .A(n34458), .B(n28895), .Z(n28548) );
  AND U29064 ( .A(n28549), .B(n28548), .Z(n28933) );
  NANDN U29065 ( .A(n32483), .B(n28550), .Z(n28552) );
  XOR U29066 ( .A(a[111]), .B(b[19]), .Z(n28971) );
  NANDN U29067 ( .A(n32823), .B(n28971), .Z(n28551) );
  AND U29068 ( .A(n28552), .B(n28551), .Z(n28932) );
  NANDN U29069 ( .A(n32013), .B(n28553), .Z(n28555) );
  XOR U29070 ( .A(a[113]), .B(b[17]), .Z(n28980) );
  NANDN U29071 ( .A(n32292), .B(n28980), .Z(n28554) );
  NAND U29072 ( .A(n28555), .B(n28554), .Z(n28931) );
  XOR U29073 ( .A(n28932), .B(n28931), .Z(n28934) );
  XOR U29074 ( .A(n28933), .B(n28934), .Z(n28984) );
  NANDN U29075 ( .A(n37526), .B(n28556), .Z(n28558) );
  XOR U29076 ( .A(b[51]), .B(a[79]), .Z(n28892) );
  NANDN U29077 ( .A(n37605), .B(n28892), .Z(n28557) );
  AND U29078 ( .A(n28558), .B(n28557), .Z(n28915) );
  NANDN U29079 ( .A(n37705), .B(n28559), .Z(n28561) );
  XOR U29080 ( .A(b[53]), .B(a[77]), .Z(n28947) );
  NANDN U29081 ( .A(n37778), .B(n28947), .Z(n28560) );
  AND U29082 ( .A(n28561), .B(n28560), .Z(n28914) );
  NANDN U29083 ( .A(n36210), .B(n28562), .Z(n28564) );
  XOR U29084 ( .A(b[39]), .B(a[91]), .Z(n28953) );
  NANDN U29085 ( .A(n36347), .B(n28953), .Z(n28563) );
  NAND U29086 ( .A(n28564), .B(n28563), .Z(n28913) );
  XOR U29087 ( .A(n28914), .B(n28913), .Z(n28916) );
  XNOR U29088 ( .A(n28915), .B(n28916), .Z(n28983) );
  XNOR U29089 ( .A(n28984), .B(n28983), .Z(n28985) );
  NANDN U29090 ( .A(n28566), .B(n28565), .Z(n28570) );
  OR U29091 ( .A(n28568), .B(n28567), .Z(n28569) );
  NAND U29092 ( .A(n28570), .B(n28569), .Z(n28986) );
  XNOR U29093 ( .A(n28985), .B(n28986), .Z(n28885) );
  NANDN U29094 ( .A(n28572), .B(n28571), .Z(n28576) );
  NANDN U29095 ( .A(n28574), .B(n28573), .Z(n28575) );
  AND U29096 ( .A(n28576), .B(n28575), .Z(n28882) );
  NANDN U29097 ( .A(n28578), .B(n28577), .Z(n28582) );
  OR U29098 ( .A(n28580), .B(n28579), .Z(n28581) );
  NAND U29099 ( .A(n28582), .B(n28581), .Z(n28883) );
  XNOR U29100 ( .A(n28882), .B(n28883), .Z(n28884) );
  XNOR U29101 ( .A(n28885), .B(n28884), .Z(n29025) );
  XOR U29102 ( .A(n29026), .B(n29025), .Z(n29028) );
  XOR U29103 ( .A(n29027), .B(n29028), .Z(n28871) );
  NANDN U29104 ( .A(n28584), .B(n28583), .Z(n28588) );
  NANDN U29105 ( .A(n28586), .B(n28585), .Z(n28587) );
  AND U29106 ( .A(n28588), .B(n28587), .Z(n28798) );
  NANDN U29107 ( .A(n211), .B(n28589), .Z(n28591) );
  XOR U29108 ( .A(b[47]), .B(a[83]), .Z(n28998) );
  NANDN U29109 ( .A(n37172), .B(n28998), .Z(n28590) );
  AND U29110 ( .A(n28591), .B(n28590), .Z(n28836) );
  NANDN U29111 ( .A(n30482), .B(n28592), .Z(n28594) );
  XOR U29112 ( .A(a[119]), .B(b[11]), .Z(n28904) );
  NANDN U29113 ( .A(n30891), .B(n28904), .Z(n28593) );
  AND U29114 ( .A(n28594), .B(n28593), .Z(n28835) );
  NANDN U29115 ( .A(n212), .B(n28595), .Z(n28597) );
  XOR U29116 ( .A(b[49]), .B(a[81]), .Z(n29001) );
  NANDN U29117 ( .A(n37432), .B(n29001), .Z(n28596) );
  NAND U29118 ( .A(n28597), .B(n28596), .Z(n28834) );
  XOR U29119 ( .A(n28835), .B(n28834), .Z(n28837) );
  XOR U29120 ( .A(n28836), .B(n28837), .Z(n28810) );
  NANDN U29121 ( .A(n36742), .B(n28598), .Z(n28600) );
  XOR U29122 ( .A(b[43]), .B(a[87]), .Z(n28898) );
  NANDN U29123 ( .A(n36891), .B(n28898), .Z(n28599) );
  AND U29124 ( .A(n28600), .B(n28599), .Z(n28909) );
  NANDN U29125 ( .A(n36991), .B(n28601), .Z(n28603) );
  XOR U29126 ( .A(b[45]), .B(a[85]), .Z(n28901) );
  NANDN U29127 ( .A(n37083), .B(n28901), .Z(n28602) );
  AND U29128 ( .A(n28603), .B(n28602), .Z(n28908) );
  NANDN U29129 ( .A(n31055), .B(n28604), .Z(n28606) );
  XOR U29130 ( .A(a[117]), .B(b[13]), .Z(n28968) );
  NANDN U29131 ( .A(n31293), .B(n28968), .Z(n28605) );
  NAND U29132 ( .A(n28606), .B(n28605), .Z(n28907) );
  XOR U29133 ( .A(n28908), .B(n28907), .Z(n28910) );
  XNOR U29134 ( .A(n28909), .B(n28910), .Z(n28809) );
  XNOR U29135 ( .A(n28810), .B(n28809), .Z(n28811) );
  NANDN U29136 ( .A(n28608), .B(n28607), .Z(n28612) );
  OR U29137 ( .A(n28610), .B(n28609), .Z(n28611) );
  NAND U29138 ( .A(n28612), .B(n28611), .Z(n28812) );
  XNOR U29139 ( .A(n28811), .B(n28812), .Z(n28797) );
  XNOR U29140 ( .A(n28798), .B(n28797), .Z(n28799) );
  NANDN U29141 ( .A(n210), .B(n28613), .Z(n28615) );
  XOR U29142 ( .A(a[121]), .B(b[9]), .Z(n28989) );
  NANDN U29143 ( .A(n30267), .B(n28989), .Z(n28614) );
  AND U29144 ( .A(n28615), .B(n28614), .Z(n29015) );
  NANDN U29145 ( .A(n37857), .B(n28616), .Z(n28618) );
  XOR U29146 ( .A(b[55]), .B(a[75]), .Z(n28950) );
  NANDN U29147 ( .A(n37911), .B(n28950), .Z(n28617) );
  AND U29148 ( .A(n28618), .B(n28617), .Z(n29014) );
  NANDN U29149 ( .A(n35611), .B(n28619), .Z(n28621) );
  XOR U29150 ( .A(b[35]), .B(a[95]), .Z(n28858) );
  NANDN U29151 ( .A(n35801), .B(n28858), .Z(n28620) );
  NAND U29152 ( .A(n28621), .B(n28620), .Z(n29013) );
  XOR U29153 ( .A(n29014), .B(n29013), .Z(n29016) );
  XOR U29154 ( .A(n29015), .B(n29016), .Z(n28822) );
  NANDN U29155 ( .A(n28623), .B(n28622), .Z(n28627) );
  OR U29156 ( .A(n28625), .B(n28624), .Z(n28626) );
  AND U29157 ( .A(n28627), .B(n28626), .Z(n28821) );
  XNOR U29158 ( .A(n28822), .B(n28821), .Z(n28823) );
  NANDN U29159 ( .A(n28629), .B(n28628), .Z(n28633) );
  OR U29160 ( .A(n28631), .B(n28630), .Z(n28632) );
  NAND U29161 ( .A(n28633), .B(n28632), .Z(n28824) );
  XOR U29162 ( .A(n28823), .B(n28824), .Z(n28800) );
  XNOR U29163 ( .A(n28799), .B(n28800), .Z(n28870) );
  XOR U29164 ( .A(n28871), .B(n28870), .Z(n28873) );
  XOR U29165 ( .A(n28872), .B(n28873), .Z(n28782) );
  NANDN U29166 ( .A(n28635), .B(n28634), .Z(n28639) );
  NANDN U29167 ( .A(n28637), .B(n28636), .Z(n28638) );
  AND U29168 ( .A(n28639), .B(n28638), .Z(n28867) );
  NANDN U29169 ( .A(n28641), .B(n28640), .Z(n28645) );
  NANDN U29170 ( .A(n28643), .B(n28642), .Z(n28644) );
  AND U29171 ( .A(n28645), .B(n28644), .Z(n28865) );
  NANDN U29172 ( .A(n28647), .B(n28646), .Z(n28651) );
  NAND U29173 ( .A(n28649), .B(n28648), .Z(n28650) );
  AND U29174 ( .A(n28651), .B(n28650), .Z(n28864) );
  XNOR U29175 ( .A(n28865), .B(n28864), .Z(n28866) );
  XNOR U29176 ( .A(n28867), .B(n28866), .Z(n28796) );
  NANDN U29177 ( .A(n28653), .B(n28652), .Z(n28657) );
  NANDN U29178 ( .A(n28655), .B(n28654), .Z(n28656) );
  NAND U29179 ( .A(n28657), .B(n28656), .Z(n29033) );
  NANDN U29180 ( .A(n33866), .B(n28658), .Z(n28660) );
  XOR U29181 ( .A(a[107]), .B(b[23]), .Z(n28977) );
  NANDN U29182 ( .A(n33644), .B(n28977), .Z(n28659) );
  AND U29183 ( .A(n28660), .B(n28659), .Z(n28842) );
  NANDN U29184 ( .A(n33875), .B(n28661), .Z(n28663) );
  XOR U29185 ( .A(a[105]), .B(b[25]), .Z(n28974) );
  NANDN U29186 ( .A(n33994), .B(n28974), .Z(n28662) );
  AND U29187 ( .A(n28663), .B(n28662), .Z(n28841) );
  NANDN U29188 ( .A(n32996), .B(n28664), .Z(n28666) );
  XOR U29189 ( .A(a[109]), .B(b[21]), .Z(n29004) );
  NANDN U29190 ( .A(n33271), .B(n29004), .Z(n28665) );
  NAND U29191 ( .A(n28666), .B(n28665), .Z(n28840) );
  XOR U29192 ( .A(n28841), .B(n28840), .Z(n28843) );
  XOR U29193 ( .A(n28842), .B(n28843), .Z(n28828) );
  NANDN U29194 ( .A(n38247), .B(n28667), .Z(n28669) );
  XOR U29195 ( .A(b[61]), .B(a[69]), .Z(n28849) );
  NANDN U29196 ( .A(n38248), .B(n28849), .Z(n28668) );
  AND U29197 ( .A(n28669), .B(n28668), .Z(n28833) );
  NAND U29198 ( .A(b[63]), .B(a[65]), .Z(n29147) );
  XOR U29199 ( .A(b[1]), .B(n29147), .Z(n28670) );
  XNOR U29200 ( .A(n28833), .B(n28670), .Z(n28827) );
  XNOR U29201 ( .A(n28828), .B(n28827), .Z(n28829) );
  NANDN U29202 ( .A(n28672), .B(n28671), .Z(n28676) );
  OR U29203 ( .A(n28674), .B(n28673), .Z(n28675) );
  NAND U29204 ( .A(n28676), .B(n28675), .Z(n28830) );
  XNOR U29205 ( .A(n28829), .B(n28830), .Z(n29032) );
  NANDN U29206 ( .A(n34634), .B(n28677), .Z(n28679) );
  XOR U29207 ( .A(a[101]), .B(b[29]), .Z(n28995) );
  NANDN U29208 ( .A(n34722), .B(n28995), .Z(n28678) );
  AND U29209 ( .A(n28679), .B(n28678), .Z(n29009) );
  NANDN U29210 ( .A(n34909), .B(n28680), .Z(n28682) );
  XOR U29211 ( .A(a[99]), .B(b[31]), .Z(n28944) );
  NANDN U29212 ( .A(n35145), .B(n28944), .Z(n28681) );
  AND U29213 ( .A(n28682), .B(n28681), .Z(n29008) );
  NANDN U29214 ( .A(n31536), .B(n28683), .Z(n28685) );
  XOR U29215 ( .A(a[115]), .B(b[15]), .Z(n28962) );
  NANDN U29216 ( .A(n31925), .B(n28962), .Z(n28684) );
  NAND U29217 ( .A(n28685), .B(n28684), .Z(n29007) );
  XOR U29218 ( .A(n29008), .B(n29007), .Z(n29010) );
  XOR U29219 ( .A(n29009), .B(n29010), .Z(n28804) );
  NANDN U29220 ( .A(n29499), .B(n28686), .Z(n28688) );
  XOR U29221 ( .A(a[123]), .B(b[7]), .Z(n28992) );
  NANDN U29222 ( .A(n29735), .B(n28992), .Z(n28687) );
  AND U29223 ( .A(n28688), .B(n28687), .Z(n29021) );
  NANDN U29224 ( .A(n28889), .B(n28689), .Z(n28691) );
  XOR U29225 ( .A(a[125]), .B(b[5]), .Z(n28888) );
  NANDN U29226 ( .A(n29138), .B(n28888), .Z(n28690) );
  AND U29227 ( .A(n28691), .B(n28690), .Z(n29020) );
  NANDN U29228 ( .A(n35936), .B(n28692), .Z(n28694) );
  XOR U29229 ( .A(b[37]), .B(a[93]), .Z(n28852) );
  NANDN U29230 ( .A(n36047), .B(n28852), .Z(n28693) );
  NAND U29231 ( .A(n28694), .B(n28693), .Z(n29019) );
  XOR U29232 ( .A(n29020), .B(n29019), .Z(n29022) );
  XNOR U29233 ( .A(n29021), .B(n29022), .Z(n28803) );
  XNOR U29234 ( .A(n28804), .B(n28803), .Z(n28805) );
  NANDN U29235 ( .A(n28696), .B(n28695), .Z(n28700) );
  OR U29236 ( .A(n28698), .B(n28697), .Z(n28699) );
  NAND U29237 ( .A(n28700), .B(n28699), .Z(n28806) );
  XNOR U29238 ( .A(n28805), .B(n28806), .Z(n29031) );
  XOR U29239 ( .A(n29032), .B(n29031), .Z(n29034) );
  XNOR U29240 ( .A(n29033), .B(n29034), .Z(n28878) );
  NANDN U29241 ( .A(n28702), .B(n28701), .Z(n28706) );
  NAND U29242 ( .A(n28704), .B(n28703), .Z(n28705) );
  AND U29243 ( .A(n28706), .B(n28705), .Z(n28876) );
  NANDN U29244 ( .A(n28708), .B(n28707), .Z(n28712) );
  OR U29245 ( .A(n28710), .B(n28709), .Z(n28711) );
  AND U29246 ( .A(n28712), .B(n28711), .Z(n28928) );
  NANDN U29247 ( .A(n37974), .B(n28713), .Z(n28715) );
  XOR U29248 ( .A(b[57]), .B(a[73]), .Z(n28937) );
  NANDN U29249 ( .A(n38031), .B(n28937), .Z(n28714) );
  AND U29250 ( .A(n28715), .B(n28714), .Z(n28958) );
  NANDN U29251 ( .A(n38090), .B(n28716), .Z(n28718) );
  XOR U29252 ( .A(b[59]), .B(a[71]), .Z(n28846) );
  NANDN U29253 ( .A(n38130), .B(n28846), .Z(n28717) );
  AND U29254 ( .A(n28718), .B(n28717), .Z(n28957) );
  NANDN U29255 ( .A(n36480), .B(n28719), .Z(n28721) );
  XOR U29256 ( .A(b[41]), .B(a[89]), .Z(n28965) );
  NANDN U29257 ( .A(n36594), .B(n28965), .Z(n28720) );
  NAND U29258 ( .A(n28721), .B(n28720), .Z(n28956) );
  XOR U29259 ( .A(n28957), .B(n28956), .Z(n28959) );
  XOR U29260 ( .A(n28958), .B(n28959), .Z(n28926) );
  NANDN U29261 ( .A(n209), .B(n28722), .Z(n28724) );
  XOR U29262 ( .A(a[127]), .B(b[3]), .Z(n28940) );
  NANDN U29263 ( .A(n28941), .B(n28940), .Z(n28723) );
  AND U29264 ( .A(n28724), .B(n28723), .Z(n28921) );
  NANDN U29265 ( .A(n38278), .B(n28725), .Z(n28727) );
  XOR U29266 ( .A(b[63]), .B(a[67]), .Z(n28855) );
  NANDN U29267 ( .A(n38279), .B(n28855), .Z(n28726) );
  AND U29268 ( .A(n28727), .B(n28726), .Z(n28920) );
  NANDN U29269 ( .A(n35260), .B(n28728), .Z(n28730) );
  XOR U29270 ( .A(b[33]), .B(a[97]), .Z(n28861) );
  NANDN U29271 ( .A(n35456), .B(n28861), .Z(n28729) );
  NAND U29272 ( .A(n28730), .B(n28729), .Z(n28919) );
  XOR U29273 ( .A(n28920), .B(n28919), .Z(n28922) );
  XNOR U29274 ( .A(n28921), .B(n28922), .Z(n28925) );
  XNOR U29275 ( .A(n28926), .B(n28925), .Z(n28927) );
  XOR U29276 ( .A(n28928), .B(n28927), .Z(n28818) );
  NANDN U29277 ( .A(n28732), .B(n28731), .Z(n28736) );
  OR U29278 ( .A(n28734), .B(n28733), .Z(n28735) );
  AND U29279 ( .A(n28736), .B(n28735), .Z(n28816) );
  NANDN U29280 ( .A(n28738), .B(n28737), .Z(n28742) );
  OR U29281 ( .A(n28740), .B(n28739), .Z(n28741) );
  NAND U29282 ( .A(n28742), .B(n28741), .Z(n28815) );
  XNOR U29283 ( .A(n28816), .B(n28815), .Z(n28817) );
  XOR U29284 ( .A(n28818), .B(n28817), .Z(n28877) );
  XOR U29285 ( .A(n28876), .B(n28877), .Z(n28879) );
  XOR U29286 ( .A(n28878), .B(n28879), .Z(n28793) );
  NANDN U29287 ( .A(n28744), .B(n28743), .Z(n28748) );
  NANDN U29288 ( .A(n28746), .B(n28745), .Z(n28747) );
  NAND U29289 ( .A(n28748), .B(n28747), .Z(n28794) );
  XOR U29290 ( .A(n28793), .B(n28794), .Z(n28795) );
  XNOR U29291 ( .A(n28796), .B(n28795), .Z(n28781) );
  XOR U29292 ( .A(n28782), .B(n28781), .Z(n28784) );
  XOR U29293 ( .A(n28783), .B(n28784), .Z(n29040) );
  XNOR U29294 ( .A(n29039), .B(n29040), .Z(n28777) );
  XOR U29295 ( .A(n28778), .B(n28777), .Z(n28770) );
  NANDN U29296 ( .A(n28750), .B(n28749), .Z(n28754) );
  OR U29297 ( .A(n28752), .B(n28751), .Z(n28753) );
  NAND U29298 ( .A(n28754), .B(n28753), .Z(n28769) );
  XNOR U29299 ( .A(n28770), .B(n28769), .Z(n28771) );
  NANDN U29300 ( .A(n28756), .B(n28755), .Z(n28760) );
  NANDN U29301 ( .A(n28758), .B(n28757), .Z(n28759) );
  NAND U29302 ( .A(n28760), .B(n28759), .Z(n28772) );
  XOR U29303 ( .A(n28771), .B(n28772), .Z(n28764) );
  XOR U29304 ( .A(n28763), .B(n28764), .Z(n28766) );
  XNOR U29305 ( .A(n28765), .B(n28766), .Z(n28761) );
  XOR U29306 ( .A(n28762), .B(n28761), .Z(c[193]) );
  AND U29307 ( .A(n28762), .B(n28761), .Z(n29044) );
  NANDN U29308 ( .A(n28764), .B(n28763), .Z(n28768) );
  OR U29309 ( .A(n28766), .B(n28765), .Z(n28767) );
  AND U29310 ( .A(n28768), .B(n28767), .Z(n29047) );
  NANDN U29311 ( .A(n28770), .B(n28769), .Z(n28774) );
  NANDN U29312 ( .A(n28772), .B(n28771), .Z(n28773) );
  AND U29313 ( .A(n28774), .B(n28773), .Z(n29046) );
  NANDN U29314 ( .A(n28776), .B(n28775), .Z(n28780) );
  NAND U29315 ( .A(n28778), .B(n28777), .Z(n28779) );
  AND U29316 ( .A(n28780), .B(n28779), .Z(n29053) );
  NANDN U29317 ( .A(n28782), .B(n28781), .Z(n28786) );
  NANDN U29318 ( .A(n28784), .B(n28783), .Z(n28785) );
  AND U29319 ( .A(n28786), .B(n28785), .Z(n29058) );
  NANDN U29320 ( .A(n28788), .B(n28787), .Z(n28792) );
  OR U29321 ( .A(n28790), .B(n28789), .Z(n28791) );
  AND U29322 ( .A(n28792), .B(n28791), .Z(n29057) );
  XNOR U29323 ( .A(n29058), .B(n29057), .Z(n29060) );
  NANDN U29324 ( .A(n28798), .B(n28797), .Z(n28802) );
  NANDN U29325 ( .A(n28800), .B(n28799), .Z(n28801) );
  AND U29326 ( .A(n28802), .B(n28801), .Z(n29312) );
  NANDN U29327 ( .A(n28804), .B(n28803), .Z(n28808) );
  NANDN U29328 ( .A(n28806), .B(n28805), .Z(n28807) );
  AND U29329 ( .A(n28808), .B(n28807), .Z(n29170) );
  NANDN U29330 ( .A(n28810), .B(n28809), .Z(n28814) );
  NANDN U29331 ( .A(n28812), .B(n28811), .Z(n28813) );
  NAND U29332 ( .A(n28814), .B(n28813), .Z(n29169) );
  XNOR U29333 ( .A(n29170), .B(n29169), .Z(n29171) );
  NANDN U29334 ( .A(n28816), .B(n28815), .Z(n28820) );
  NANDN U29335 ( .A(n28818), .B(n28817), .Z(n28819) );
  NAND U29336 ( .A(n28820), .B(n28819), .Z(n29172) );
  XNOR U29337 ( .A(n29171), .B(n29172), .Z(n29310) );
  NANDN U29338 ( .A(n28822), .B(n28821), .Z(n28826) );
  NANDN U29339 ( .A(n28824), .B(n28823), .Z(n28825) );
  AND U29340 ( .A(n28826), .B(n28825), .Z(n29178) );
  NANDN U29341 ( .A(n28828), .B(n28827), .Z(n28832) );
  NANDN U29342 ( .A(n28830), .B(n28829), .Z(n28831) );
  AND U29343 ( .A(n28832), .B(n28831), .Z(n29176) );
  NANDN U29344 ( .A(n28835), .B(n28834), .Z(n28839) );
  OR U29345 ( .A(n28837), .B(n28836), .Z(n28838) );
  NAND U29346 ( .A(n28839), .B(n28838), .Z(n29188) );
  XNOR U29347 ( .A(n29187), .B(n29188), .Z(n29189) );
  NANDN U29348 ( .A(n28841), .B(n28840), .Z(n28845) );
  OR U29349 ( .A(n28843), .B(n28842), .Z(n28844) );
  AND U29350 ( .A(n28845), .B(n28844), .Z(n29201) );
  NANDN U29351 ( .A(n38090), .B(n28846), .Z(n28848) );
  XOR U29352 ( .A(b[59]), .B(a[72]), .Z(n29247) );
  NANDN U29353 ( .A(n38130), .B(n29247), .Z(n28847) );
  AND U29354 ( .A(n28848), .B(n28847), .Z(n29288) );
  NANDN U29355 ( .A(n38247), .B(n28849), .Z(n28851) );
  XOR U29356 ( .A(b[61]), .B(a[70]), .Z(n29250) );
  NANDN U29357 ( .A(n38248), .B(n29250), .Z(n28850) );
  AND U29358 ( .A(n28851), .B(n28850), .Z(n29287) );
  NANDN U29359 ( .A(n35936), .B(n28852), .Z(n28854) );
  XOR U29360 ( .A(b[37]), .B(a[94]), .Z(n29142) );
  NANDN U29361 ( .A(n36047), .B(n29142), .Z(n28853) );
  NAND U29362 ( .A(n28854), .B(n28853), .Z(n29286) );
  XOR U29363 ( .A(n29287), .B(n29286), .Z(n29289) );
  XOR U29364 ( .A(n29288), .B(n29289), .Z(n29200) );
  NANDN U29365 ( .A(n38278), .B(n28855), .Z(n28857) );
  XOR U29366 ( .A(b[63]), .B(a[68]), .Z(n29105) );
  NANDN U29367 ( .A(n38279), .B(n29105), .Z(n28856) );
  AND U29368 ( .A(n28857), .B(n28856), .Z(n29242) );
  NANDN U29369 ( .A(n35611), .B(n28858), .Z(n28860) );
  XOR U29370 ( .A(b[35]), .B(a[96]), .Z(n29271) );
  NANDN U29371 ( .A(n35801), .B(n29271), .Z(n28859) );
  NAND U29372 ( .A(n28860), .B(n28859), .Z(n29241) );
  XNOR U29373 ( .A(n29242), .B(n29241), .Z(n29244) );
  NAND U29374 ( .A(n35654), .B(n28861), .Z(n28863) );
  XNOR U29375 ( .A(a[98]), .B(b[33]), .Z(n29220) );
  NANDN U29376 ( .A(n29220), .B(n35655), .Z(n28862) );
  NAND U29377 ( .A(n28863), .B(n28862), .Z(n29145) );
  AND U29378 ( .A(b[63]), .B(a[66]), .Z(n29146) );
  XOR U29379 ( .A(n29145), .B(n29146), .Z(n29148) );
  XOR U29380 ( .A(n29147), .B(n29148), .Z(n29243) );
  XNOR U29381 ( .A(n29244), .B(n29243), .Z(n29199) );
  XOR U29382 ( .A(n29200), .B(n29199), .Z(n29202) );
  XOR U29383 ( .A(n29201), .B(n29202), .Z(n29190) );
  XNOR U29384 ( .A(n29189), .B(n29190), .Z(n29175) );
  XNOR U29385 ( .A(n29176), .B(n29175), .Z(n29177) );
  XOR U29386 ( .A(n29178), .B(n29177), .Z(n29311) );
  XOR U29387 ( .A(n29310), .B(n29311), .Z(n29313) );
  XOR U29388 ( .A(n29312), .B(n29313), .Z(n29317) );
  NANDN U29389 ( .A(n28865), .B(n28864), .Z(n28869) );
  NANDN U29390 ( .A(n28867), .B(n28866), .Z(n28868) );
  AND U29391 ( .A(n28869), .B(n28868), .Z(n29316) );
  XOR U29392 ( .A(n29317), .B(n29316), .Z(n29319) );
  XNOR U29393 ( .A(n29318), .B(n29319), .Z(n29065) );
  NANDN U29394 ( .A(n28871), .B(n28870), .Z(n28875) );
  OR U29395 ( .A(n28873), .B(n28872), .Z(n28874) );
  AND U29396 ( .A(n28875), .B(n28874), .Z(n29063) );
  NANDN U29397 ( .A(n28877), .B(n28876), .Z(n28881) );
  NANDN U29398 ( .A(n28879), .B(n28878), .Z(n28880) );
  AND U29399 ( .A(n28881), .B(n28880), .Z(n29307) );
  NANDN U29400 ( .A(n28883), .B(n28882), .Z(n28887) );
  NAND U29401 ( .A(n28885), .B(n28884), .Z(n28886) );
  AND U29402 ( .A(n28887), .B(n28886), .Z(n29183) );
  NANDN U29403 ( .A(n28889), .B(n28888), .Z(n28891) );
  XOR U29404 ( .A(a[126]), .B(b[5]), .Z(n29139) );
  NANDN U29405 ( .A(n29138), .B(n29139), .Z(n28890) );
  AND U29406 ( .A(n28891), .B(n28890), .Z(n29282) );
  NANDN U29407 ( .A(n37526), .B(n28892), .Z(n28894) );
  XOR U29408 ( .A(b[51]), .B(a[80]), .Z(n29217) );
  NANDN U29409 ( .A(n37605), .B(n29217), .Z(n28893) );
  AND U29410 ( .A(n28894), .B(n28893), .Z(n29281) );
  NANDN U29411 ( .A(n34223), .B(n28895), .Z(n28897) );
  XOR U29412 ( .A(a[104]), .B(b[27]), .Z(n29111) );
  NANDN U29413 ( .A(n34458), .B(n29111), .Z(n28896) );
  NAND U29414 ( .A(n28897), .B(n28896), .Z(n29280) );
  XOR U29415 ( .A(n29281), .B(n29280), .Z(n29283) );
  XOR U29416 ( .A(n29282), .B(n29283), .Z(n29164) );
  NANDN U29417 ( .A(n36742), .B(n28898), .Z(n28900) );
  XOR U29418 ( .A(b[43]), .B(a[88]), .Z(n29256) );
  NANDN U29419 ( .A(n36891), .B(n29256), .Z(n28899) );
  AND U29420 ( .A(n28900), .B(n28899), .Z(n29225) );
  NANDN U29421 ( .A(n36991), .B(n28901), .Z(n28903) );
  XOR U29422 ( .A(b[45]), .B(a[86]), .Z(n29259) );
  NANDN U29423 ( .A(n37083), .B(n29259), .Z(n28902) );
  AND U29424 ( .A(n28903), .B(n28902), .Z(n29224) );
  NANDN U29425 ( .A(n30482), .B(n28904), .Z(n28906) );
  XOR U29426 ( .A(a[120]), .B(b[11]), .Z(n29214) );
  NANDN U29427 ( .A(n30891), .B(n29214), .Z(n28905) );
  NAND U29428 ( .A(n28906), .B(n28905), .Z(n29223) );
  XOR U29429 ( .A(n29224), .B(n29223), .Z(n29226) );
  XNOR U29430 ( .A(n29225), .B(n29226), .Z(n29163) );
  XNOR U29431 ( .A(n29164), .B(n29163), .Z(n29166) );
  NANDN U29432 ( .A(n28908), .B(n28907), .Z(n28912) );
  OR U29433 ( .A(n28910), .B(n28909), .Z(n28911) );
  AND U29434 ( .A(n28912), .B(n28911), .Z(n29165) );
  XOR U29435 ( .A(n29166), .B(n29165), .Z(n29300) );
  NANDN U29436 ( .A(n28914), .B(n28913), .Z(n28918) );
  OR U29437 ( .A(n28916), .B(n28915), .Z(n28917) );
  AND U29438 ( .A(n28918), .B(n28917), .Z(n29299) );
  NANDN U29439 ( .A(n28920), .B(n28919), .Z(n28924) );
  OR U29440 ( .A(n28922), .B(n28921), .Z(n28923) );
  NAND U29441 ( .A(n28924), .B(n28923), .Z(n29298) );
  XOR U29442 ( .A(n29299), .B(n29298), .Z(n29301) );
  XOR U29443 ( .A(n29300), .B(n29301), .Z(n29182) );
  NANDN U29444 ( .A(n28926), .B(n28925), .Z(n28930) );
  NAND U29445 ( .A(n28928), .B(n28927), .Z(n28929) );
  NAND U29446 ( .A(n28930), .B(n28929), .Z(n29181) );
  XOR U29447 ( .A(n29182), .B(n29181), .Z(n29184) );
  XOR U29448 ( .A(n29183), .B(n29184), .Z(n29305) );
  NANDN U29449 ( .A(n28932), .B(n28931), .Z(n28936) );
  OR U29450 ( .A(n28934), .B(n28933), .Z(n28935) );
  AND U29451 ( .A(n28936), .B(n28935), .Z(n29294) );
  NANDN U29452 ( .A(n37974), .B(n28937), .Z(n28939) );
  XOR U29453 ( .A(b[57]), .B(a[74]), .Z(n29268) );
  NANDN U29454 ( .A(n38031), .B(n29268), .Z(n28938) );
  AND U29455 ( .A(n28939), .B(n28938), .Z(n29159) );
  NANDN U29456 ( .A(n209), .B(n28940), .Z(n28943) );
  NANDN U29457 ( .A(n28941), .B(b[3]), .Z(n28942) );
  AND U29458 ( .A(n28943), .B(n28942), .Z(n29158) );
  NANDN U29459 ( .A(n34909), .B(n28944), .Z(n28946) );
  XOR U29460 ( .A(a[100]), .B(b[31]), .Z(n29211) );
  NANDN U29461 ( .A(n35145), .B(n29211), .Z(n28945) );
  NAND U29462 ( .A(n28946), .B(n28945), .Z(n29157) );
  XOR U29463 ( .A(n29158), .B(n29157), .Z(n29160) );
  XOR U29464 ( .A(n29159), .B(n29160), .Z(n29293) );
  NANDN U29465 ( .A(n37705), .B(n28947), .Z(n28949) );
  XOR U29466 ( .A(b[53]), .B(a[78]), .Z(n29205) );
  NANDN U29467 ( .A(n37778), .B(n29205), .Z(n28948) );
  AND U29468 ( .A(n28949), .B(n28948), .Z(n29153) );
  NANDN U29469 ( .A(n37857), .B(n28950), .Z(n28952) );
  XOR U29470 ( .A(b[55]), .B(a[76]), .Z(n29265) );
  NANDN U29471 ( .A(n37911), .B(n29265), .Z(n28951) );
  AND U29472 ( .A(n28952), .B(n28951), .Z(n29152) );
  NANDN U29473 ( .A(n36210), .B(n28953), .Z(n28955) );
  XOR U29474 ( .A(b[39]), .B(a[92]), .Z(n29108) );
  NANDN U29475 ( .A(n36347), .B(n29108), .Z(n28954) );
  NAND U29476 ( .A(n28955), .B(n28954), .Z(n29151) );
  XOR U29477 ( .A(n29152), .B(n29151), .Z(n29154) );
  XNOR U29478 ( .A(n29153), .B(n29154), .Z(n29292) );
  XOR U29479 ( .A(n29293), .B(n29292), .Z(n29295) );
  XNOR U29480 ( .A(n29294), .B(n29295), .Z(n29075) );
  NANDN U29481 ( .A(n28957), .B(n28956), .Z(n28961) );
  OR U29482 ( .A(n28959), .B(n28958), .Z(n28960) );
  NAND U29483 ( .A(n28961), .B(n28960), .Z(n29076) );
  XNOR U29484 ( .A(n29075), .B(n29076), .Z(n29078) );
  NANDN U29485 ( .A(n31536), .B(n28962), .Z(n28964) );
  XOR U29486 ( .A(a[116]), .B(b[15]), .Z(n29117) );
  NANDN U29487 ( .A(n31925), .B(n29117), .Z(n28963) );
  AND U29488 ( .A(n28964), .B(n28963), .Z(n29276) );
  NANDN U29489 ( .A(n36480), .B(n28965), .Z(n28967) );
  XOR U29490 ( .A(b[41]), .B(a[90]), .Z(n29253) );
  NANDN U29491 ( .A(n36594), .B(n29253), .Z(n28966) );
  AND U29492 ( .A(n28967), .B(n28966), .Z(n29275) );
  NANDN U29493 ( .A(n31055), .B(n28968), .Z(n28970) );
  XOR U29494 ( .A(a[118]), .B(b[13]), .Z(n29262) );
  NANDN U29495 ( .A(n31293), .B(n29262), .Z(n28969) );
  NAND U29496 ( .A(n28970), .B(n28969), .Z(n29274) );
  XOR U29497 ( .A(n29275), .B(n29274), .Z(n29277) );
  XOR U29498 ( .A(n29276), .B(n29277), .Z(n29232) );
  NANDN U29499 ( .A(n32483), .B(n28971), .Z(n28973) );
  XOR U29500 ( .A(a[112]), .B(b[19]), .Z(n29120) );
  NANDN U29501 ( .A(n32823), .B(n29120), .Z(n28972) );
  AND U29502 ( .A(n28973), .B(n28972), .Z(n29134) );
  NANDN U29503 ( .A(n33875), .B(n28974), .Z(n28976) );
  XOR U29504 ( .A(a[106]), .B(b[25]), .Z(n29123) );
  NANDN U29505 ( .A(n33994), .B(n29123), .Z(n28975) );
  AND U29506 ( .A(n28976), .B(n28975), .Z(n29133) );
  NANDN U29507 ( .A(n33866), .B(n28977), .Z(n28979) );
  XOR U29508 ( .A(a[108]), .B(b[23]), .Z(n29099) );
  NANDN U29509 ( .A(n33644), .B(n29099), .Z(n28978) );
  NAND U29510 ( .A(n28979), .B(n28978), .Z(n29132) );
  XOR U29511 ( .A(n29133), .B(n29132), .Z(n29135) );
  XOR U29512 ( .A(n29134), .B(n29135), .Z(n29230) );
  NAND U29513 ( .A(n32544), .B(n28980), .Z(n28982) );
  XNOR U29514 ( .A(a[114]), .B(b[17]), .Z(n29129) );
  NANDN U29515 ( .A(n29129), .B(n32545), .Z(n28981) );
  AND U29516 ( .A(n28982), .B(n28981), .Z(n29229) );
  XNOR U29517 ( .A(n29230), .B(n29229), .Z(n29231) );
  XNOR U29518 ( .A(n29232), .B(n29231), .Z(n29077) );
  XOR U29519 ( .A(n29078), .B(n29077), .Z(n29072) );
  NANDN U29520 ( .A(n28984), .B(n28983), .Z(n28988) );
  NANDN U29521 ( .A(n28986), .B(n28985), .Z(n28987) );
  AND U29522 ( .A(n28988), .B(n28987), .Z(n29069) );
  NANDN U29523 ( .A(n210), .B(n28989), .Z(n28991) );
  XOR U29524 ( .A(a[122]), .B(b[9]), .Z(n29208) );
  NANDN U29525 ( .A(n30267), .B(n29208), .Z(n28990) );
  AND U29526 ( .A(n28991), .B(n28990), .Z(n29089) );
  NANDN U29527 ( .A(n29499), .B(n28992), .Z(n28994) );
  XOR U29528 ( .A(a[124]), .B(b[7]), .Z(n29102) );
  NANDN U29529 ( .A(n29735), .B(n29102), .Z(n28993) );
  AND U29530 ( .A(n28994), .B(n28993), .Z(n29088) );
  NANDN U29531 ( .A(n34634), .B(n28995), .Z(n28997) );
  XOR U29532 ( .A(a[102]), .B(b[29]), .Z(n29114) );
  NANDN U29533 ( .A(n34722), .B(n29114), .Z(n28996) );
  NAND U29534 ( .A(n28997), .B(n28996), .Z(n29087) );
  XOR U29535 ( .A(n29088), .B(n29087), .Z(n29090) );
  XOR U29536 ( .A(n29089), .B(n29090), .Z(n29082) );
  NAND U29537 ( .A(n37294), .B(n28998), .Z(n29000) );
  XNOR U29538 ( .A(b[47]), .B(a[84]), .Z(n29093) );
  NANDN U29539 ( .A(n29093), .B(n37341), .Z(n28999) );
  NAND U29540 ( .A(n29000), .B(n28999), .Z(n29237) );
  NAND U29541 ( .A(n37536), .B(n29001), .Z(n29003) );
  XNOR U29542 ( .A(b[49]), .B(a[82]), .Z(n29096) );
  NANDN U29543 ( .A(n29096), .B(n37537), .Z(n29002) );
  NAND U29544 ( .A(n29003), .B(n29002), .Z(n29236) );
  NAND U29545 ( .A(n33413), .B(n29004), .Z(n29006) );
  XNOR U29546 ( .A(a[110]), .B(b[21]), .Z(n29126) );
  NANDN U29547 ( .A(n29126), .B(n33414), .Z(n29005) );
  NAND U29548 ( .A(n29006), .B(n29005), .Z(n29235) );
  XNOR U29549 ( .A(n29236), .B(n29235), .Z(n29238) );
  XOR U29550 ( .A(n29237), .B(n29238), .Z(n29081) );
  XNOR U29551 ( .A(n29082), .B(n29081), .Z(n29084) );
  NANDN U29552 ( .A(n29008), .B(n29007), .Z(n29012) );
  OR U29553 ( .A(n29010), .B(n29009), .Z(n29011) );
  AND U29554 ( .A(n29012), .B(n29011), .Z(n29083) );
  XOR U29555 ( .A(n29084), .B(n29083), .Z(n29196) );
  NANDN U29556 ( .A(n29014), .B(n29013), .Z(n29018) );
  OR U29557 ( .A(n29016), .B(n29015), .Z(n29017) );
  AND U29558 ( .A(n29018), .B(n29017), .Z(n29194) );
  NANDN U29559 ( .A(n29020), .B(n29019), .Z(n29024) );
  OR U29560 ( .A(n29022), .B(n29021), .Z(n29023) );
  NAND U29561 ( .A(n29024), .B(n29023), .Z(n29193) );
  XNOR U29562 ( .A(n29194), .B(n29193), .Z(n29195) );
  XOR U29563 ( .A(n29196), .B(n29195), .Z(n29070) );
  XNOR U29564 ( .A(n29069), .B(n29070), .Z(n29071) );
  XNOR U29565 ( .A(n29072), .B(n29071), .Z(n29304) );
  XNOR U29566 ( .A(n29305), .B(n29304), .Z(n29306) );
  XNOR U29567 ( .A(n29307), .B(n29306), .Z(n29324) );
  NANDN U29568 ( .A(n29026), .B(n29025), .Z(n29030) );
  OR U29569 ( .A(n29028), .B(n29027), .Z(n29029) );
  AND U29570 ( .A(n29030), .B(n29029), .Z(n29323) );
  NAND U29571 ( .A(n29032), .B(n29031), .Z(n29036) );
  NAND U29572 ( .A(n29034), .B(n29033), .Z(n29035) );
  AND U29573 ( .A(n29036), .B(n29035), .Z(n29322) );
  XOR U29574 ( .A(n29323), .B(n29322), .Z(n29325) );
  XOR U29575 ( .A(n29324), .B(n29325), .Z(n29064) );
  XOR U29576 ( .A(n29063), .B(n29064), .Z(n29066) );
  XNOR U29577 ( .A(n29065), .B(n29066), .Z(n29059) );
  XOR U29578 ( .A(n29060), .B(n29059), .Z(n29052) );
  NANDN U29579 ( .A(n29038), .B(n29037), .Z(n29042) );
  NANDN U29580 ( .A(n29040), .B(n29039), .Z(n29041) );
  AND U29581 ( .A(n29042), .B(n29041), .Z(n29051) );
  XOR U29582 ( .A(n29052), .B(n29051), .Z(n29054) );
  XNOR U29583 ( .A(n29053), .B(n29054), .Z(n29045) );
  XOR U29584 ( .A(n29046), .B(n29045), .Z(n29048) );
  XNOR U29585 ( .A(n29047), .B(n29048), .Z(n29043) );
  XOR U29586 ( .A(n29044), .B(n29043), .Z(c[194]) );
  AND U29587 ( .A(n29044), .B(n29043), .Z(n29329) );
  NANDN U29588 ( .A(n29046), .B(n29045), .Z(n29050) );
  OR U29589 ( .A(n29048), .B(n29047), .Z(n29049) );
  AND U29590 ( .A(n29050), .B(n29049), .Z(n29332) );
  NANDN U29591 ( .A(n29052), .B(n29051), .Z(n29056) );
  NANDN U29592 ( .A(n29054), .B(n29053), .Z(n29055) );
  AND U29593 ( .A(n29056), .B(n29055), .Z(n29331) );
  NANDN U29594 ( .A(n29058), .B(n29057), .Z(n29062) );
  NAND U29595 ( .A(n29060), .B(n29059), .Z(n29061) );
  AND U29596 ( .A(n29062), .B(n29061), .Z(n29339) );
  NANDN U29597 ( .A(n29064), .B(n29063), .Z(n29068) );
  NANDN U29598 ( .A(n29066), .B(n29065), .Z(n29067) );
  AND U29599 ( .A(n29068), .B(n29067), .Z(n29337) );
  NANDN U29600 ( .A(n29070), .B(n29069), .Z(n29074) );
  NANDN U29601 ( .A(n29072), .B(n29071), .Z(n29073) );
  AND U29602 ( .A(n29074), .B(n29073), .Z(n29575) );
  NANDN U29603 ( .A(n29076), .B(n29075), .Z(n29080) );
  NAND U29604 ( .A(n29078), .B(n29077), .Z(n29079) );
  AND U29605 ( .A(n29080), .B(n29079), .Z(n29574) );
  NANDN U29606 ( .A(n29082), .B(n29081), .Z(n29086) );
  NAND U29607 ( .A(n29084), .B(n29083), .Z(n29085) );
  AND U29608 ( .A(n29086), .B(n29085), .Z(n29480) );
  NANDN U29609 ( .A(n29088), .B(n29087), .Z(n29092) );
  OR U29610 ( .A(n29090), .B(n29089), .Z(n29091) );
  AND U29611 ( .A(n29092), .B(n29091), .Z(n29468) );
  NANDN U29612 ( .A(n29093), .B(n37294), .Z(n29095) );
  XOR U29613 ( .A(b[47]), .B(a[85]), .Z(n29492) );
  NANDN U29614 ( .A(n37172), .B(n29492), .Z(n29094) );
  AND U29615 ( .A(n29095), .B(n29094), .Z(n29378) );
  NANDN U29616 ( .A(n29096), .B(n37536), .Z(n29098) );
  XOR U29617 ( .A(b[49]), .B(a[83]), .Z(n29393) );
  NANDN U29618 ( .A(n37432), .B(n29393), .Z(n29097) );
  AND U29619 ( .A(n29098), .B(n29097), .Z(n29376) );
  NANDN U29620 ( .A(n33866), .B(n29099), .Z(n29101) );
  XOR U29621 ( .A(a[109]), .B(b[23]), .Z(n29495) );
  NANDN U29622 ( .A(n33644), .B(n29495), .Z(n29100) );
  NAND U29623 ( .A(n29101), .B(n29100), .Z(n29375) );
  XNOR U29624 ( .A(n29376), .B(n29375), .Z(n29377) );
  XOR U29625 ( .A(n29378), .B(n29377), .Z(n29466) );
  NANDN U29626 ( .A(n29499), .B(n29102), .Z(n29104) );
  XOR U29627 ( .A(a[125]), .B(b[7]), .Z(n29498) );
  NANDN U29628 ( .A(n29735), .B(n29498), .Z(n29103) );
  AND U29629 ( .A(n29104), .B(n29103), .Z(n29443) );
  NANDN U29630 ( .A(n38278), .B(n29105), .Z(n29107) );
  XOR U29631 ( .A(b[63]), .B(a[69]), .Z(n29547) );
  NANDN U29632 ( .A(n38279), .B(n29547), .Z(n29106) );
  AND U29633 ( .A(n29107), .B(n29106), .Z(n29442) );
  NANDN U29634 ( .A(n36210), .B(n29108), .Z(n29110) );
  XOR U29635 ( .A(b[39]), .B(a[93]), .Z(n29368) );
  NANDN U29636 ( .A(n36347), .B(n29368), .Z(n29109) );
  NAND U29637 ( .A(n29110), .B(n29109), .Z(n29441) );
  XOR U29638 ( .A(n29442), .B(n29441), .Z(n29444) );
  XNOR U29639 ( .A(n29443), .B(n29444), .Z(n29465) );
  XOR U29640 ( .A(n29466), .B(n29465), .Z(n29467) );
  XOR U29641 ( .A(n29468), .B(n29467), .Z(n29478) );
  NANDN U29642 ( .A(n34223), .B(n29111), .Z(n29113) );
  XOR U29643 ( .A(a[105]), .B(b[27]), .Z(n29514) );
  NANDN U29644 ( .A(n34458), .B(n29514), .Z(n29112) );
  AND U29645 ( .A(n29113), .B(n29112), .Z(n29432) );
  NANDN U29646 ( .A(n34634), .B(n29114), .Z(n29116) );
  XOR U29647 ( .A(a[103]), .B(b[29]), .Z(n29517) );
  NANDN U29648 ( .A(n34722), .B(n29517), .Z(n29115) );
  AND U29649 ( .A(n29116), .B(n29115), .Z(n29430) );
  NANDN U29650 ( .A(n31536), .B(n29117), .Z(n29119) );
  XOR U29651 ( .A(a[117]), .B(b[15]), .Z(n29520) );
  NANDN U29652 ( .A(n31925), .B(n29520), .Z(n29118) );
  NAND U29653 ( .A(n29119), .B(n29118), .Z(n29429) );
  XNOR U29654 ( .A(n29430), .B(n29429), .Z(n29431) );
  XOR U29655 ( .A(n29432), .B(n29431), .Z(n29407) );
  NANDN U29656 ( .A(n32483), .B(n29120), .Z(n29122) );
  XOR U29657 ( .A(a[113]), .B(b[19]), .Z(n29523) );
  NANDN U29658 ( .A(n32823), .B(n29523), .Z(n29121) );
  AND U29659 ( .A(n29122), .B(n29121), .Z(n29564) );
  NANDN U29660 ( .A(n33875), .B(n29123), .Z(n29125) );
  XOR U29661 ( .A(a[107]), .B(b[25]), .Z(n29526) );
  NANDN U29662 ( .A(n33994), .B(n29526), .Z(n29124) );
  AND U29663 ( .A(n29125), .B(n29124), .Z(n29562) );
  NANDN U29664 ( .A(n29126), .B(n33413), .Z(n29128) );
  XOR U29665 ( .A(a[111]), .B(b[21]), .Z(n29529) );
  NANDN U29666 ( .A(n33271), .B(n29529), .Z(n29127) );
  NAND U29667 ( .A(n29128), .B(n29127), .Z(n29561) );
  XNOR U29668 ( .A(n29562), .B(n29561), .Z(n29563) );
  XOR U29669 ( .A(n29564), .B(n29563), .Z(n29405) );
  NANDN U29670 ( .A(n29129), .B(n32544), .Z(n29131) );
  XOR U29671 ( .A(a[115]), .B(b[17]), .Z(n29532) );
  NANDN U29672 ( .A(n32292), .B(n29532), .Z(n29130) );
  AND U29673 ( .A(n29131), .B(n29130), .Z(n29406) );
  XNOR U29674 ( .A(n29405), .B(n29406), .Z(n29408) );
  XOR U29675 ( .A(n29407), .B(n29408), .Z(n29477) );
  XNOR U29676 ( .A(n29478), .B(n29477), .Z(n29479) );
  XOR U29677 ( .A(n29480), .B(n29479), .Z(n29359) );
  NANDN U29678 ( .A(n29133), .B(n29132), .Z(n29137) );
  OR U29679 ( .A(n29135), .B(n29134), .Z(n29136) );
  AND U29680 ( .A(n29137), .B(n29136), .Z(n29450) );
  XNOR U29681 ( .A(a[127]), .B(b[5]), .Z(n29550) );
  OR U29682 ( .A(n29550), .B(n29138), .Z(n29141) );
  NAND U29683 ( .A(n29551), .B(n29139), .Z(n29140) );
  AND U29684 ( .A(n29141), .B(n29140), .Z(n29372) );
  NANDN U29685 ( .A(n35936), .B(n29142), .Z(n29144) );
  XOR U29686 ( .A(b[37]), .B(a[95]), .Z(n29505) );
  NANDN U29687 ( .A(n36047), .B(n29505), .Z(n29143) );
  NAND U29688 ( .A(n29144), .B(n29143), .Z(n29371) );
  XNOR U29689 ( .A(n29372), .B(n29371), .Z(n29374) );
  AND U29690 ( .A(b[63]), .B(a[67]), .Z(n29555) );
  XOR U29691 ( .A(n29556), .B(n29555), .Z(n29558) );
  XOR U29692 ( .A(n29147), .B(n29558), .Z(n29373) );
  XOR U29693 ( .A(n29374), .B(n29373), .Z(n29448) );
  NAND U29694 ( .A(n29146), .B(n29145), .Z(n29150) );
  IV U29695 ( .A(n29147), .Z(n29557) );
  NANDN U29696 ( .A(n29557), .B(n29148), .Z(n29149) );
  AND U29697 ( .A(n29150), .B(n29149), .Z(n29447) );
  XOR U29698 ( .A(n29450), .B(n29449), .Z(n29473) );
  NANDN U29699 ( .A(n29152), .B(n29151), .Z(n29156) );
  OR U29700 ( .A(n29154), .B(n29153), .Z(n29155) );
  AND U29701 ( .A(n29156), .B(n29155), .Z(n29472) );
  NANDN U29702 ( .A(n29158), .B(n29157), .Z(n29162) );
  OR U29703 ( .A(n29160), .B(n29159), .Z(n29161) );
  NAND U29704 ( .A(n29162), .B(n29161), .Z(n29471) );
  XOR U29705 ( .A(n29472), .B(n29471), .Z(n29474) );
  XOR U29706 ( .A(n29473), .B(n29474), .Z(n29357) );
  NANDN U29707 ( .A(n29164), .B(n29163), .Z(n29168) );
  NAND U29708 ( .A(n29166), .B(n29165), .Z(n29167) );
  NAND U29709 ( .A(n29168), .B(n29167), .Z(n29356) );
  XNOR U29710 ( .A(n29357), .B(n29356), .Z(n29358) );
  XNOR U29711 ( .A(n29359), .B(n29358), .Z(n29573) );
  XOR U29712 ( .A(n29574), .B(n29573), .Z(n29576) );
  XOR U29713 ( .A(n29575), .B(n29576), .Z(n29346) );
  NANDN U29714 ( .A(n29170), .B(n29169), .Z(n29174) );
  NANDN U29715 ( .A(n29172), .B(n29171), .Z(n29173) );
  AND U29716 ( .A(n29174), .B(n29173), .Z(n29345) );
  NANDN U29717 ( .A(n29176), .B(n29175), .Z(n29180) );
  NANDN U29718 ( .A(n29178), .B(n29177), .Z(n29179) );
  AND U29719 ( .A(n29180), .B(n29179), .Z(n29344) );
  XOR U29720 ( .A(n29345), .B(n29344), .Z(n29347) );
  XNOR U29721 ( .A(n29346), .B(n29347), .Z(n29352) );
  NANDN U29722 ( .A(n29182), .B(n29181), .Z(n29186) );
  OR U29723 ( .A(n29184), .B(n29183), .Z(n29185) );
  AND U29724 ( .A(n29186), .B(n29185), .Z(n29351) );
  NANDN U29725 ( .A(n29188), .B(n29187), .Z(n29192) );
  NANDN U29726 ( .A(n29190), .B(n29189), .Z(n29191) );
  AND U29727 ( .A(n29192), .B(n29191), .Z(n29594) );
  NANDN U29728 ( .A(n29194), .B(n29193), .Z(n29198) );
  NANDN U29729 ( .A(n29196), .B(n29195), .Z(n29197) );
  AND U29730 ( .A(n29198), .B(n29197), .Z(n29592) );
  NANDN U29731 ( .A(n29200), .B(n29199), .Z(n29204) );
  NANDN U29732 ( .A(n29202), .B(n29201), .Z(n29203) );
  AND U29733 ( .A(n29204), .B(n29203), .Z(n29591) );
  XNOR U29734 ( .A(n29592), .B(n29591), .Z(n29593) );
  XOR U29735 ( .A(n29594), .B(n29593), .Z(n29600) );
  NANDN U29736 ( .A(n37705), .B(n29205), .Z(n29207) );
  XOR U29737 ( .A(b[53]), .B(a[79]), .Z(n29420) );
  NANDN U29738 ( .A(n37778), .B(n29420), .Z(n29206) );
  AND U29739 ( .A(n29207), .B(n29206), .Z(n29437) );
  NANDN U29740 ( .A(n210), .B(n29208), .Z(n29210) );
  XOR U29741 ( .A(a[123]), .B(b[9]), .Z(n29384) );
  NANDN U29742 ( .A(n30267), .B(n29384), .Z(n29209) );
  AND U29743 ( .A(n29210), .B(n29209), .Z(n29436) );
  NANDN U29744 ( .A(n34909), .B(n29211), .Z(n29213) );
  XOR U29745 ( .A(a[101]), .B(b[31]), .Z(n29387) );
  NANDN U29746 ( .A(n35145), .B(n29387), .Z(n29212) );
  NAND U29747 ( .A(n29213), .B(n29212), .Z(n29435) );
  XOR U29748 ( .A(n29436), .B(n29435), .Z(n29438) );
  XOR U29749 ( .A(n29437), .B(n29438), .Z(n29484) );
  NANDN U29750 ( .A(n30482), .B(n29214), .Z(n29216) );
  XOR U29751 ( .A(a[121]), .B(b[11]), .Z(n29390) );
  NANDN U29752 ( .A(n30891), .B(n29390), .Z(n29215) );
  AND U29753 ( .A(n29216), .B(n29215), .Z(n29510) );
  NANDN U29754 ( .A(n37526), .B(n29217), .Z(n29219) );
  XOR U29755 ( .A(b[51]), .B(a[81]), .Z(n29381) );
  NANDN U29756 ( .A(n37605), .B(n29381), .Z(n29218) );
  AND U29757 ( .A(n29219), .B(n29218), .Z(n29509) );
  NANDN U29758 ( .A(n29220), .B(n35654), .Z(n29222) );
  XOR U29759 ( .A(a[99]), .B(b[33]), .Z(n29396) );
  NANDN U29760 ( .A(n35456), .B(n29396), .Z(n29221) );
  NAND U29761 ( .A(n29222), .B(n29221), .Z(n29508) );
  XOR U29762 ( .A(n29509), .B(n29508), .Z(n29511) );
  XNOR U29763 ( .A(n29510), .B(n29511), .Z(n29483) );
  XNOR U29764 ( .A(n29484), .B(n29483), .Z(n29486) );
  NANDN U29765 ( .A(n29224), .B(n29223), .Z(n29228) );
  OR U29766 ( .A(n29226), .B(n29225), .Z(n29227) );
  AND U29767 ( .A(n29228), .B(n29227), .Z(n29485) );
  XOR U29768 ( .A(n29486), .B(n29485), .Z(n29586) );
  NANDN U29769 ( .A(n29230), .B(n29229), .Z(n29234) );
  NANDN U29770 ( .A(n29232), .B(n29231), .Z(n29233) );
  AND U29771 ( .A(n29234), .B(n29233), .Z(n29585) );
  XNOR U29772 ( .A(n29586), .B(n29585), .Z(n29588) );
  NAND U29773 ( .A(n29236), .B(n29235), .Z(n29240) );
  NANDN U29774 ( .A(n29238), .B(n29237), .Z(n29239) );
  AND U29775 ( .A(n29240), .B(n29239), .Z(n29462) );
  NANDN U29776 ( .A(n29242), .B(n29241), .Z(n29246) );
  NAND U29777 ( .A(n29244), .B(n29243), .Z(n29245) );
  AND U29778 ( .A(n29246), .B(n29245), .Z(n29460) );
  NANDN U29779 ( .A(n38090), .B(n29247), .Z(n29249) );
  XOR U29780 ( .A(b[59]), .B(a[73]), .Z(n29365) );
  NANDN U29781 ( .A(n38130), .B(n29365), .Z(n29248) );
  AND U29782 ( .A(n29249), .B(n29248), .Z(n29544) );
  NANDN U29783 ( .A(n38247), .B(n29250), .Z(n29252) );
  XOR U29784 ( .A(b[61]), .B(a[71]), .Z(n29502) );
  NANDN U29785 ( .A(n38248), .B(n29502), .Z(n29251) );
  AND U29786 ( .A(n29252), .B(n29251), .Z(n29542) );
  NANDN U29787 ( .A(n36480), .B(n29253), .Z(n29255) );
  XOR U29788 ( .A(b[41]), .B(a[91]), .Z(n29411) );
  NANDN U29789 ( .A(n36594), .B(n29411), .Z(n29254) );
  NAND U29790 ( .A(n29255), .B(n29254), .Z(n29541) );
  XNOR U29791 ( .A(n29542), .B(n29541), .Z(n29543) );
  XNOR U29792 ( .A(n29544), .B(n29543), .Z(n29459) );
  XNOR U29793 ( .A(n29460), .B(n29459), .Z(n29461) );
  XNOR U29794 ( .A(n29462), .B(n29461), .Z(n29587) );
  XOR U29795 ( .A(n29588), .B(n29587), .Z(n29598) );
  NANDN U29796 ( .A(n36742), .B(n29256), .Z(n29258) );
  XOR U29797 ( .A(b[43]), .B(a[89]), .Z(n29414) );
  NANDN U29798 ( .A(n36891), .B(n29414), .Z(n29257) );
  AND U29799 ( .A(n29258), .B(n29257), .Z(n29401) );
  NANDN U29800 ( .A(n36991), .B(n29259), .Z(n29261) );
  XOR U29801 ( .A(b[45]), .B(a[87]), .Z(n29489) );
  NANDN U29802 ( .A(n37083), .B(n29489), .Z(n29260) );
  AND U29803 ( .A(n29261), .B(n29260), .Z(n29400) );
  NANDN U29804 ( .A(n31055), .B(n29262), .Z(n29264) );
  XOR U29805 ( .A(a[119]), .B(b[13]), .Z(n29417) );
  NANDN U29806 ( .A(n31293), .B(n29417), .Z(n29263) );
  NAND U29807 ( .A(n29264), .B(n29263), .Z(n29399) );
  XOR U29808 ( .A(n29400), .B(n29399), .Z(n29402) );
  XOR U29809 ( .A(n29401), .B(n29402), .Z(n29568) );
  NANDN U29810 ( .A(n37857), .B(n29265), .Z(n29267) );
  XOR U29811 ( .A(b[55]), .B(a[77]), .Z(n29423) );
  NANDN U29812 ( .A(n37911), .B(n29423), .Z(n29266) );
  AND U29813 ( .A(n29267), .B(n29266), .Z(n29537) );
  NANDN U29814 ( .A(n37974), .B(n29268), .Z(n29270) );
  XOR U29815 ( .A(b[57]), .B(a[75]), .Z(n29362) );
  NANDN U29816 ( .A(n38031), .B(n29362), .Z(n29269) );
  AND U29817 ( .A(n29270), .B(n29269), .Z(n29536) );
  NANDN U29818 ( .A(n35611), .B(n29271), .Z(n29273) );
  XOR U29819 ( .A(b[35]), .B(a[97]), .Z(n29426) );
  NANDN U29820 ( .A(n35801), .B(n29426), .Z(n29272) );
  NAND U29821 ( .A(n29273), .B(n29272), .Z(n29535) );
  XOR U29822 ( .A(n29536), .B(n29535), .Z(n29538) );
  XNOR U29823 ( .A(n29537), .B(n29538), .Z(n29567) );
  XNOR U29824 ( .A(n29568), .B(n29567), .Z(n29570) );
  NANDN U29825 ( .A(n29275), .B(n29274), .Z(n29279) );
  OR U29826 ( .A(n29277), .B(n29276), .Z(n29278) );
  AND U29827 ( .A(n29279), .B(n29278), .Z(n29569) );
  XOR U29828 ( .A(n29570), .B(n29569), .Z(n29455) );
  NANDN U29829 ( .A(n29281), .B(n29280), .Z(n29285) );
  OR U29830 ( .A(n29283), .B(n29282), .Z(n29284) );
  AND U29831 ( .A(n29285), .B(n29284), .Z(n29454) );
  NANDN U29832 ( .A(n29287), .B(n29286), .Z(n29291) );
  OR U29833 ( .A(n29289), .B(n29288), .Z(n29290) );
  NAND U29834 ( .A(n29291), .B(n29290), .Z(n29453) );
  XOR U29835 ( .A(n29454), .B(n29453), .Z(n29456) );
  XOR U29836 ( .A(n29455), .B(n29456), .Z(n29580) );
  NANDN U29837 ( .A(n29293), .B(n29292), .Z(n29297) );
  NANDN U29838 ( .A(n29295), .B(n29294), .Z(n29296) );
  NAND U29839 ( .A(n29297), .B(n29296), .Z(n29579) );
  XNOR U29840 ( .A(n29580), .B(n29579), .Z(n29581) );
  NANDN U29841 ( .A(n29299), .B(n29298), .Z(n29303) );
  OR U29842 ( .A(n29301), .B(n29300), .Z(n29302) );
  NAND U29843 ( .A(n29303), .B(n29302), .Z(n29582) );
  XNOR U29844 ( .A(n29581), .B(n29582), .Z(n29597) );
  XNOR U29845 ( .A(n29598), .B(n29597), .Z(n29599) );
  XNOR U29846 ( .A(n29600), .B(n29599), .Z(n29350) );
  XOR U29847 ( .A(n29351), .B(n29350), .Z(n29353) );
  XOR U29848 ( .A(n29352), .B(n29353), .Z(n29605) );
  NANDN U29849 ( .A(n29305), .B(n29304), .Z(n29309) );
  NANDN U29850 ( .A(n29307), .B(n29306), .Z(n29308) );
  AND U29851 ( .A(n29309), .B(n29308), .Z(n29604) );
  NANDN U29852 ( .A(n29311), .B(n29310), .Z(n29315) );
  OR U29853 ( .A(n29313), .B(n29312), .Z(n29314) );
  AND U29854 ( .A(n29315), .B(n29314), .Z(n29603) );
  XOR U29855 ( .A(n29604), .B(n29603), .Z(n29606) );
  XOR U29856 ( .A(n29605), .B(n29606), .Z(n29342) );
  NANDN U29857 ( .A(n29317), .B(n29316), .Z(n29321) );
  NANDN U29858 ( .A(n29319), .B(n29318), .Z(n29320) );
  AND U29859 ( .A(n29321), .B(n29320), .Z(n29340) );
  NANDN U29860 ( .A(n29323), .B(n29322), .Z(n29327) );
  NANDN U29861 ( .A(n29325), .B(n29324), .Z(n29326) );
  NAND U29862 ( .A(n29327), .B(n29326), .Z(n29341) );
  XNOR U29863 ( .A(n29340), .B(n29341), .Z(n29343) );
  XOR U29864 ( .A(n29342), .B(n29343), .Z(n29336) );
  XOR U29865 ( .A(n29337), .B(n29336), .Z(n29338) );
  XOR U29866 ( .A(n29339), .B(n29338), .Z(n29330) );
  XOR U29867 ( .A(n29331), .B(n29330), .Z(n29333) );
  XNOR U29868 ( .A(n29332), .B(n29333), .Z(n29328) );
  XOR U29869 ( .A(n29329), .B(n29328), .Z(c[195]) );
  AND U29870 ( .A(n29329), .B(n29328), .Z(n29610) );
  NANDN U29871 ( .A(n29331), .B(n29330), .Z(n29335) );
  OR U29872 ( .A(n29333), .B(n29332), .Z(n29334) );
  AND U29873 ( .A(n29335), .B(n29334), .Z(n29613) );
  NAND U29874 ( .A(n29345), .B(n29344), .Z(n29349) );
  NAND U29875 ( .A(n29347), .B(n29346), .Z(n29348) );
  AND U29876 ( .A(n29349), .B(n29348), .Z(n29624) );
  NANDN U29877 ( .A(n29351), .B(n29350), .Z(n29355) );
  NANDN U29878 ( .A(n29353), .B(n29352), .Z(n29354) );
  AND U29879 ( .A(n29355), .B(n29354), .Z(n29623) );
  XNOR U29880 ( .A(n29624), .B(n29623), .Z(n29626) );
  NANDN U29881 ( .A(n29357), .B(n29356), .Z(n29361) );
  NANDN U29882 ( .A(n29359), .B(n29358), .Z(n29360) );
  AND U29883 ( .A(n29361), .B(n29360), .Z(n29631) );
  NANDN U29884 ( .A(n37974), .B(n29362), .Z(n29364) );
  XOR U29885 ( .A(b[57]), .B(a[76]), .Z(n29802) );
  NANDN U29886 ( .A(n38031), .B(n29802), .Z(n29363) );
  AND U29887 ( .A(n29364), .B(n29363), .Z(n29750) );
  NANDN U29888 ( .A(n38090), .B(n29365), .Z(n29367) );
  XOR U29889 ( .A(b[59]), .B(a[74]), .Z(n29732) );
  NANDN U29890 ( .A(n38130), .B(n29732), .Z(n29366) );
  AND U29891 ( .A(n29367), .B(n29366), .Z(n29749) );
  NANDN U29892 ( .A(n36210), .B(n29368), .Z(n29370) );
  XOR U29893 ( .A(b[39]), .B(a[94]), .Z(n29729) );
  NANDN U29894 ( .A(n36347), .B(n29729), .Z(n29369) );
  NAND U29895 ( .A(n29370), .B(n29369), .Z(n29748) );
  XOR U29896 ( .A(n29749), .B(n29748), .Z(n29751) );
  XOR U29897 ( .A(n29750), .B(n29751), .Z(n29821) );
  XNOR U29898 ( .A(n29821), .B(n29820), .Z(n29823) );
  NANDN U29899 ( .A(n29376), .B(n29375), .Z(n29380) );
  NANDN U29900 ( .A(n29378), .B(n29377), .Z(n29379) );
  AND U29901 ( .A(n29380), .B(n29379), .Z(n29822) );
  XOR U29902 ( .A(n29823), .B(n29822), .Z(n29649) );
  NANDN U29903 ( .A(n37526), .B(n29381), .Z(n29383) );
  XOR U29904 ( .A(b[51]), .B(a[82]), .Z(n29693) );
  NANDN U29905 ( .A(n37605), .B(n29693), .Z(n29382) );
  AND U29906 ( .A(n29383), .B(n29382), .Z(n29682) );
  NANDN U29907 ( .A(n210), .B(n29384), .Z(n29386) );
  XOR U29908 ( .A(a[124]), .B(b[9]), .Z(n29799) );
  NANDN U29909 ( .A(n30267), .B(n29799), .Z(n29385) );
  AND U29910 ( .A(n29386), .B(n29385), .Z(n29681) );
  NANDN U29911 ( .A(n34909), .B(n29387), .Z(n29389) );
  XOR U29912 ( .A(a[102]), .B(b[31]), .Z(n29760) );
  NANDN U29913 ( .A(n35145), .B(n29760), .Z(n29388) );
  NAND U29914 ( .A(n29389), .B(n29388), .Z(n29680) );
  XOR U29915 ( .A(n29681), .B(n29680), .Z(n29683) );
  XOR U29916 ( .A(n29682), .B(n29683), .Z(n29827) );
  NANDN U29917 ( .A(n30482), .B(n29390), .Z(n29392) );
  XOR U29918 ( .A(a[122]), .B(b[11]), .Z(n29757) );
  NANDN U29919 ( .A(n30891), .B(n29757), .Z(n29391) );
  AND U29920 ( .A(n29392), .B(n29391), .Z(n29713) );
  NANDN U29921 ( .A(n212), .B(n29393), .Z(n29395) );
  XOR U29922 ( .A(b[49]), .B(a[84]), .Z(n29705) );
  NANDN U29923 ( .A(n37432), .B(n29705), .Z(n29394) );
  AND U29924 ( .A(n29395), .B(n29394), .Z(n29712) );
  NANDN U29925 ( .A(n35260), .B(n29396), .Z(n29398) );
  XOR U29926 ( .A(a[100]), .B(b[33]), .Z(n29739) );
  NANDN U29927 ( .A(n35456), .B(n29739), .Z(n29397) );
  NAND U29928 ( .A(n29398), .B(n29397), .Z(n29711) );
  XOR U29929 ( .A(n29712), .B(n29711), .Z(n29714) );
  XNOR U29930 ( .A(n29713), .B(n29714), .Z(n29826) );
  XNOR U29931 ( .A(n29827), .B(n29826), .Z(n29829) );
  NANDN U29932 ( .A(n29400), .B(n29399), .Z(n29404) );
  OR U29933 ( .A(n29402), .B(n29401), .Z(n29403) );
  AND U29934 ( .A(n29404), .B(n29403), .Z(n29828) );
  XOR U29935 ( .A(n29829), .B(n29828), .Z(n29648) );
  NAND U29936 ( .A(n29406), .B(n29405), .Z(n29410) );
  NANDN U29937 ( .A(n29408), .B(n29407), .Z(n29409) );
  AND U29938 ( .A(n29410), .B(n29409), .Z(n29647) );
  XOR U29939 ( .A(n29648), .B(n29647), .Z(n29650) );
  XOR U29940 ( .A(n29649), .B(n29650), .Z(n29630) );
  NANDN U29941 ( .A(n36480), .B(n29411), .Z(n29413) );
  XOR U29942 ( .A(b[41]), .B(a[92]), .Z(n29805) );
  NANDN U29943 ( .A(n36594), .B(n29805), .Z(n29412) );
  AND U29944 ( .A(n29413), .B(n29412), .Z(n29744) );
  NANDN U29945 ( .A(n36742), .B(n29414), .Z(n29416) );
  XOR U29946 ( .A(b[43]), .B(a[90]), .Z(n29662) );
  NANDN U29947 ( .A(n36891), .B(n29662), .Z(n29415) );
  AND U29948 ( .A(n29416), .B(n29415), .Z(n29743) );
  NANDN U29949 ( .A(n31055), .B(n29417), .Z(n29419) );
  XOR U29950 ( .A(a[120]), .B(b[13]), .Z(n29754) );
  NANDN U29951 ( .A(n31293), .B(n29754), .Z(n29418) );
  NAND U29952 ( .A(n29419), .B(n29418), .Z(n29742) );
  XOR U29953 ( .A(n29743), .B(n29742), .Z(n29745) );
  XOR U29954 ( .A(n29744), .B(n29745), .Z(n29851) );
  NANDN U29955 ( .A(n37705), .B(n29420), .Z(n29422) );
  XOR U29956 ( .A(b[53]), .B(a[80]), .Z(n29769) );
  NANDN U29957 ( .A(n37778), .B(n29769), .Z(n29421) );
  AND U29958 ( .A(n29422), .B(n29421), .Z(n29810) );
  NANDN U29959 ( .A(n37857), .B(n29423), .Z(n29425) );
  XOR U29960 ( .A(b[55]), .B(a[78]), .Z(n29696) );
  NANDN U29961 ( .A(n37911), .B(n29696), .Z(n29424) );
  AND U29962 ( .A(n29425), .B(n29424), .Z(n29809) );
  NANDN U29963 ( .A(n35611), .B(n29426), .Z(n29428) );
  XOR U29964 ( .A(b[35]), .B(a[98]), .Z(n29671) );
  NANDN U29965 ( .A(n35801), .B(n29671), .Z(n29427) );
  NAND U29966 ( .A(n29428), .B(n29427), .Z(n29808) );
  XOR U29967 ( .A(n29809), .B(n29808), .Z(n29811) );
  XNOR U29968 ( .A(n29810), .B(n29811), .Z(n29850) );
  XNOR U29969 ( .A(n29851), .B(n29850), .Z(n29853) );
  NANDN U29970 ( .A(n29430), .B(n29429), .Z(n29434) );
  NANDN U29971 ( .A(n29432), .B(n29431), .Z(n29433) );
  AND U29972 ( .A(n29434), .B(n29433), .Z(n29852) );
  XOR U29973 ( .A(n29853), .B(n29852), .Z(n29834) );
  NANDN U29974 ( .A(n29436), .B(n29435), .Z(n29440) );
  OR U29975 ( .A(n29438), .B(n29437), .Z(n29439) );
  AND U29976 ( .A(n29440), .B(n29439), .Z(n29833) );
  NANDN U29977 ( .A(n29442), .B(n29441), .Z(n29446) );
  OR U29978 ( .A(n29444), .B(n29443), .Z(n29445) );
  NAND U29979 ( .A(n29446), .B(n29445), .Z(n29832) );
  XOR U29980 ( .A(n29833), .B(n29832), .Z(n29835) );
  XOR U29981 ( .A(n29834), .B(n29835), .Z(n29642) );
  NANDN U29982 ( .A(n29448), .B(n29447), .Z(n29452) );
  NAND U29983 ( .A(n29450), .B(n29449), .Z(n29451) );
  NAND U29984 ( .A(n29452), .B(n29451), .Z(n29641) );
  XNOR U29985 ( .A(n29642), .B(n29641), .Z(n29643) );
  NANDN U29986 ( .A(n29454), .B(n29453), .Z(n29458) );
  OR U29987 ( .A(n29456), .B(n29455), .Z(n29457) );
  NAND U29988 ( .A(n29458), .B(n29457), .Z(n29644) );
  XNOR U29989 ( .A(n29643), .B(n29644), .Z(n29629) );
  XOR U29990 ( .A(n29630), .B(n29629), .Z(n29632) );
  XOR U29991 ( .A(n29631), .B(n29632), .Z(n29869) );
  NANDN U29992 ( .A(n29460), .B(n29459), .Z(n29464) );
  NANDN U29993 ( .A(n29462), .B(n29461), .Z(n29463) );
  AND U29994 ( .A(n29464), .B(n29463), .Z(n29638) );
  NAND U29995 ( .A(n29466), .B(n29465), .Z(n29470) );
  NAND U29996 ( .A(n29468), .B(n29467), .Z(n29469) );
  NAND U29997 ( .A(n29470), .B(n29469), .Z(n29635) );
  NANDN U29998 ( .A(n29472), .B(n29471), .Z(n29476) );
  OR U29999 ( .A(n29474), .B(n29473), .Z(n29475) );
  AND U30000 ( .A(n29476), .B(n29475), .Z(n29636) );
  XOR U30001 ( .A(n29635), .B(n29636), .Z(n29637) );
  XOR U30002 ( .A(n29638), .B(n29637), .Z(n29865) );
  NANDN U30003 ( .A(n29478), .B(n29477), .Z(n29482) );
  NAND U30004 ( .A(n29480), .B(n29479), .Z(n29481) );
  AND U30005 ( .A(n29482), .B(n29481), .Z(n29863) );
  NANDN U30006 ( .A(n29484), .B(n29483), .Z(n29488) );
  NAND U30007 ( .A(n29486), .B(n29485), .Z(n29487) );
  AND U30008 ( .A(n29488), .B(n29487), .Z(n29841) );
  NANDN U30009 ( .A(n36991), .B(n29489), .Z(n29491) );
  XOR U30010 ( .A(b[45]), .B(a[88]), .Z(n29790) );
  NANDN U30011 ( .A(n37083), .B(n29790), .Z(n29490) );
  AND U30012 ( .A(n29491), .B(n29490), .Z(n29774) );
  NANDN U30013 ( .A(n211), .B(n29492), .Z(n29494) );
  XOR U30014 ( .A(b[47]), .B(a[86]), .Z(n29702) );
  NANDN U30015 ( .A(n37172), .B(n29702), .Z(n29493) );
  AND U30016 ( .A(n29494), .B(n29493), .Z(n29773) );
  NANDN U30017 ( .A(n33866), .B(n29495), .Z(n29497) );
  XOR U30018 ( .A(a[110]), .B(b[23]), .Z(n29796) );
  NANDN U30019 ( .A(n33644), .B(n29796), .Z(n29496) );
  NAND U30020 ( .A(n29497), .B(n29496), .Z(n29772) );
  XOR U30021 ( .A(n29773), .B(n29772), .Z(n29775) );
  XOR U30022 ( .A(n29774), .B(n29775), .Z(n29845) );
  NANDN U30023 ( .A(n29499), .B(n29498), .Z(n29501) );
  XOR U30024 ( .A(a[126]), .B(b[7]), .Z(n29736) );
  NANDN U30025 ( .A(n29735), .B(n29736), .Z(n29500) );
  AND U30026 ( .A(n29501), .B(n29500), .Z(n29816) );
  NANDN U30027 ( .A(n38247), .B(n29502), .Z(n29504) );
  XOR U30028 ( .A(b[61]), .B(a[72]), .Z(n29723) );
  NANDN U30029 ( .A(n38248), .B(n29723), .Z(n29503) );
  AND U30030 ( .A(n29504), .B(n29503), .Z(n29815) );
  NANDN U30031 ( .A(n35936), .B(n29505), .Z(n29507) );
  XOR U30032 ( .A(b[37]), .B(a[96]), .Z(n29668) );
  NANDN U30033 ( .A(n36047), .B(n29668), .Z(n29506) );
  NAND U30034 ( .A(n29507), .B(n29506), .Z(n29814) );
  XOR U30035 ( .A(n29815), .B(n29814), .Z(n29817) );
  XNOR U30036 ( .A(n29816), .B(n29817), .Z(n29844) );
  XNOR U30037 ( .A(n29845), .B(n29844), .Z(n29847) );
  NANDN U30038 ( .A(n29509), .B(n29508), .Z(n29513) );
  OR U30039 ( .A(n29511), .B(n29510), .Z(n29512) );
  AND U30040 ( .A(n29513), .B(n29512), .Z(n29846) );
  XOR U30041 ( .A(n29847), .B(n29846), .Z(n29839) );
  NANDN U30042 ( .A(n34223), .B(n29514), .Z(n29516) );
  XOR U30043 ( .A(a[106]), .B(b[27]), .Z(n29665) );
  NANDN U30044 ( .A(n34458), .B(n29665), .Z(n29515) );
  AND U30045 ( .A(n29516), .B(n29515), .Z(n29676) );
  NANDN U30046 ( .A(n34634), .B(n29517), .Z(n29519) );
  XOR U30047 ( .A(a[104]), .B(b[29]), .Z(n29659) );
  NANDN U30048 ( .A(n34722), .B(n29659), .Z(n29518) );
  AND U30049 ( .A(n29519), .B(n29518), .Z(n29675) );
  NANDN U30050 ( .A(n31536), .B(n29520), .Z(n29522) );
  XOR U30051 ( .A(a[118]), .B(b[15]), .Z(n29766) );
  NANDN U30052 ( .A(n31925), .B(n29766), .Z(n29521) );
  NAND U30053 ( .A(n29522), .B(n29521), .Z(n29674) );
  XOR U30054 ( .A(n29675), .B(n29674), .Z(n29677) );
  XOR U30055 ( .A(n29676), .B(n29677), .Z(n29719) );
  NANDN U30056 ( .A(n32483), .B(n29523), .Z(n29525) );
  XOR U30057 ( .A(a[114]), .B(b[19]), .Z(n29699) );
  NANDN U30058 ( .A(n32823), .B(n29699), .Z(n29524) );
  AND U30059 ( .A(n29525), .B(n29524), .Z(n29786) );
  NANDN U30060 ( .A(n33875), .B(n29526), .Z(n29528) );
  XOR U30061 ( .A(a[108]), .B(b[25]), .Z(n29793) );
  NANDN U30062 ( .A(n33994), .B(n29793), .Z(n29527) );
  AND U30063 ( .A(n29528), .B(n29527), .Z(n29785) );
  NANDN U30064 ( .A(n32996), .B(n29529), .Z(n29531) );
  XOR U30065 ( .A(a[112]), .B(b[21]), .Z(n29708) );
  NANDN U30066 ( .A(n33271), .B(n29708), .Z(n29530) );
  NAND U30067 ( .A(n29531), .B(n29530), .Z(n29784) );
  XOR U30068 ( .A(n29785), .B(n29784), .Z(n29787) );
  XOR U30069 ( .A(n29786), .B(n29787), .Z(n29718) );
  NAND U30070 ( .A(n32544), .B(n29532), .Z(n29534) );
  XNOR U30071 ( .A(a[116]), .B(b[17]), .Z(n29763) );
  NANDN U30072 ( .A(n29763), .B(n32545), .Z(n29533) );
  AND U30073 ( .A(n29534), .B(n29533), .Z(n29717) );
  XOR U30074 ( .A(n29718), .B(n29717), .Z(n29720) );
  XNOR U30075 ( .A(n29719), .B(n29720), .Z(n29838) );
  XNOR U30076 ( .A(n29839), .B(n29838), .Z(n29840) );
  XOR U30077 ( .A(n29841), .B(n29840), .Z(n29655) );
  NANDN U30078 ( .A(n29536), .B(n29535), .Z(n29540) );
  OR U30079 ( .A(n29538), .B(n29537), .Z(n29539) );
  AND U30080 ( .A(n29540), .B(n29539), .Z(n29857) );
  NANDN U30081 ( .A(n29542), .B(n29541), .Z(n29546) );
  NANDN U30082 ( .A(n29544), .B(n29543), .Z(n29545) );
  NAND U30083 ( .A(n29546), .B(n29545), .Z(n29856) );
  XNOR U30084 ( .A(n29857), .B(n29856), .Z(n29859) );
  NANDN U30085 ( .A(n38278), .B(n29547), .Z(n29549) );
  XOR U30086 ( .A(b[63]), .B(a[70]), .Z(n29726) );
  NANDN U30087 ( .A(n38279), .B(n29726), .Z(n29548) );
  AND U30088 ( .A(n29549), .B(n29548), .Z(n29689) );
  NAND U30089 ( .A(b[63]), .B(a[68]), .Z(n30085) );
  ANDN U30090 ( .B(n29551), .A(n29550), .Z(n29554) );
  NAND U30091 ( .A(b[5]), .B(n29552), .Z(n29553) );
  NANDN U30092 ( .A(n29554), .B(n29553), .Z(n29686) );
  XOR U30093 ( .A(n30085), .B(n29686), .Z(n29688) );
  XNOR U30094 ( .A(n29689), .B(n29688), .Z(n29779) );
  NANDN U30095 ( .A(n29556), .B(n29555), .Z(n29560) );
  NANDN U30096 ( .A(n29558), .B(n29557), .Z(n29559) );
  NAND U30097 ( .A(n29560), .B(n29559), .Z(n29778) );
  XOR U30098 ( .A(n29779), .B(n29778), .Z(n29781) );
  NANDN U30099 ( .A(n29562), .B(n29561), .Z(n29566) );
  NANDN U30100 ( .A(n29564), .B(n29563), .Z(n29565) );
  NAND U30101 ( .A(n29566), .B(n29565), .Z(n29780) );
  XOR U30102 ( .A(n29781), .B(n29780), .Z(n29858) );
  XOR U30103 ( .A(n29859), .B(n29858), .Z(n29654) );
  NANDN U30104 ( .A(n29568), .B(n29567), .Z(n29572) );
  NAND U30105 ( .A(n29570), .B(n29569), .Z(n29571) );
  NAND U30106 ( .A(n29572), .B(n29571), .Z(n29653) );
  XOR U30107 ( .A(n29654), .B(n29653), .Z(n29656) );
  XNOR U30108 ( .A(n29655), .B(n29656), .Z(n29862) );
  XNOR U30109 ( .A(n29863), .B(n29862), .Z(n29864) );
  XNOR U30110 ( .A(n29865), .B(n29864), .Z(n29868) );
  XNOR U30111 ( .A(n29869), .B(n29868), .Z(n29870) );
  NANDN U30112 ( .A(n29574), .B(n29573), .Z(n29578) );
  NANDN U30113 ( .A(n29576), .B(n29575), .Z(n29577) );
  NAND U30114 ( .A(n29578), .B(n29577), .Z(n29871) );
  XNOR U30115 ( .A(n29870), .B(n29871), .Z(n29882) );
  NANDN U30116 ( .A(n29580), .B(n29579), .Z(n29584) );
  NANDN U30117 ( .A(n29582), .B(n29581), .Z(n29583) );
  AND U30118 ( .A(n29584), .B(n29583), .Z(n29875) );
  NANDN U30119 ( .A(n29586), .B(n29585), .Z(n29590) );
  NAND U30120 ( .A(n29588), .B(n29587), .Z(n29589) );
  AND U30121 ( .A(n29590), .B(n29589), .Z(n29874) );
  XNOR U30122 ( .A(n29875), .B(n29874), .Z(n29877) );
  NANDN U30123 ( .A(n29592), .B(n29591), .Z(n29596) );
  NAND U30124 ( .A(n29594), .B(n29593), .Z(n29595) );
  AND U30125 ( .A(n29596), .B(n29595), .Z(n29876) );
  XOR U30126 ( .A(n29877), .B(n29876), .Z(n29881) );
  NANDN U30127 ( .A(n29598), .B(n29597), .Z(n29602) );
  NANDN U30128 ( .A(n29600), .B(n29599), .Z(n29601) );
  AND U30129 ( .A(n29602), .B(n29601), .Z(n29880) );
  XOR U30130 ( .A(n29881), .B(n29880), .Z(n29883) );
  XNOR U30131 ( .A(n29882), .B(n29883), .Z(n29625) );
  XOR U30132 ( .A(n29626), .B(n29625), .Z(n29618) );
  NANDN U30133 ( .A(n29604), .B(n29603), .Z(n29608) );
  NANDN U30134 ( .A(n29606), .B(n29605), .Z(n29607) );
  AND U30135 ( .A(n29608), .B(n29607), .Z(n29617) );
  XNOR U30136 ( .A(n29618), .B(n29617), .Z(n29619) );
  XNOR U30137 ( .A(n29620), .B(n29619), .Z(n29611) );
  XOR U30138 ( .A(n29612), .B(n29611), .Z(n29614) );
  XNOR U30139 ( .A(n29613), .B(n29614), .Z(n29609) );
  XOR U30140 ( .A(n29610), .B(n29609), .Z(c[196]) );
  AND U30141 ( .A(n29610), .B(n29609), .Z(n29887) );
  NANDN U30142 ( .A(n29612), .B(n29611), .Z(n29616) );
  OR U30143 ( .A(n29614), .B(n29613), .Z(n29615) );
  AND U30144 ( .A(n29616), .B(n29615), .Z(n29890) );
  NANDN U30145 ( .A(n29618), .B(n29617), .Z(n29622) );
  NANDN U30146 ( .A(n29620), .B(n29619), .Z(n29621) );
  AND U30147 ( .A(n29622), .B(n29621), .Z(n29889) );
  NANDN U30148 ( .A(n29624), .B(n29623), .Z(n29628) );
  NAND U30149 ( .A(n29626), .B(n29625), .Z(n29627) );
  AND U30150 ( .A(n29628), .B(n29627), .Z(n29896) );
  NANDN U30151 ( .A(n29630), .B(n29629), .Z(n29634) );
  OR U30152 ( .A(n29632), .B(n29631), .Z(n29633) );
  AND U30153 ( .A(n29634), .B(n29633), .Z(n29907) );
  NAND U30154 ( .A(n29636), .B(n29635), .Z(n29640) );
  NAND U30155 ( .A(n29638), .B(n29637), .Z(n29639) );
  AND U30156 ( .A(n29640), .B(n29639), .Z(n30155) );
  NANDN U30157 ( .A(n29642), .B(n29641), .Z(n29646) );
  NANDN U30158 ( .A(n29644), .B(n29643), .Z(n29645) );
  AND U30159 ( .A(n29646), .B(n29645), .Z(n30153) );
  NANDN U30160 ( .A(n29648), .B(n29647), .Z(n29652) );
  OR U30161 ( .A(n29650), .B(n29649), .Z(n29651) );
  AND U30162 ( .A(n29652), .B(n29651), .Z(n30152) );
  XNOR U30163 ( .A(n30153), .B(n30152), .Z(n30154) );
  XNOR U30164 ( .A(n30155), .B(n30154), .Z(n29906) );
  XNOR U30165 ( .A(n29907), .B(n29906), .Z(n29909) );
  NANDN U30166 ( .A(n29654), .B(n29653), .Z(n29658) );
  OR U30167 ( .A(n29656), .B(n29655), .Z(n29657) );
  AND U30168 ( .A(n29658), .B(n29657), .Z(n30143) );
  NANDN U30169 ( .A(n34634), .B(n29659), .Z(n29661) );
  XOR U30170 ( .A(a[105]), .B(b[29]), .Z(n29990) );
  NANDN U30171 ( .A(n34722), .B(n29990), .Z(n29660) );
  AND U30172 ( .A(n29661), .B(n29660), .Z(n30091) );
  NANDN U30173 ( .A(n36742), .B(n29662), .Z(n29664) );
  XOR U30174 ( .A(b[43]), .B(a[91]), .Z(n30055) );
  NANDN U30175 ( .A(n36891), .B(n30055), .Z(n29663) );
  AND U30176 ( .A(n29664), .B(n29663), .Z(n30089) );
  NANDN U30177 ( .A(n34223), .B(n29665), .Z(n29667) );
  XOR U30178 ( .A(a[107]), .B(b[27]), .Z(n29996) );
  NANDN U30179 ( .A(n34458), .B(n29996), .Z(n29666) );
  NAND U30180 ( .A(n29667), .B(n29666), .Z(n30088) );
  XNOR U30181 ( .A(n30089), .B(n30088), .Z(n30090) );
  XOR U30182 ( .A(n30091), .B(n30090), .Z(n29985) );
  NANDN U30183 ( .A(n35936), .B(n29668), .Z(n29670) );
  XOR U30184 ( .A(b[37]), .B(a[97]), .Z(n29957) );
  NANDN U30185 ( .A(n36047), .B(n29957), .Z(n29669) );
  NAND U30186 ( .A(n29670), .B(n29669), .Z(n30103) );
  XNOR U30187 ( .A(n30104), .B(n30103), .Z(n30106) );
  IV U30188 ( .A(n30085), .Z(n29687) );
  AND U30189 ( .A(b[63]), .B(a[69]), .Z(n30083) );
  NANDN U30190 ( .A(n35611), .B(n29671), .Z(n29673) );
  XOR U30191 ( .A(b[35]), .B(a[99]), .Z(n29942) );
  NANDN U30192 ( .A(n35801), .B(n29942), .Z(n29672) );
  NAND U30193 ( .A(n29673), .B(n29672), .Z(n30082) );
  XOR U30194 ( .A(n30083), .B(n30082), .Z(n30084) );
  XOR U30195 ( .A(n29687), .B(n30084), .Z(n30105) );
  XNOR U30196 ( .A(n30106), .B(n30105), .Z(n29984) );
  XOR U30197 ( .A(n29985), .B(n29984), .Z(n29987) );
  NANDN U30198 ( .A(n29675), .B(n29674), .Z(n29679) );
  OR U30199 ( .A(n29677), .B(n29676), .Z(n29678) );
  AND U30200 ( .A(n29679), .B(n29678), .Z(n29986) );
  XOR U30201 ( .A(n29987), .B(n29986), .Z(n30117) );
  NANDN U30202 ( .A(n29681), .B(n29680), .Z(n29685) );
  OR U30203 ( .A(n29683), .B(n29682), .Z(n29684) );
  AND U30204 ( .A(n29685), .B(n29684), .Z(n30116) );
  NANDN U30205 ( .A(n29687), .B(n29686), .Z(n29691) );
  NANDN U30206 ( .A(n29689), .B(n29688), .Z(n29690) );
  NAND U30207 ( .A(n29691), .B(n29690), .Z(n30115) );
  XOR U30208 ( .A(n30116), .B(n30115), .Z(n29692) );
  XOR U30209 ( .A(n30117), .B(n29692), .Z(n30138) );
  NANDN U30210 ( .A(n37526), .B(n29693), .Z(n29695) );
  XOR U30211 ( .A(b[51]), .B(a[83]), .Z(n29924) );
  NANDN U30212 ( .A(n37605), .B(n29924), .Z(n29694) );
  AND U30213 ( .A(n29695), .B(n29694), .Z(n30009) );
  NANDN U30214 ( .A(n37857), .B(n29696), .Z(n29698) );
  XOR U30215 ( .A(b[55]), .B(a[79]), .Z(n30061) );
  NANDN U30216 ( .A(n37911), .B(n30061), .Z(n29697) );
  AND U30217 ( .A(n29698), .B(n29697), .Z(n30008) );
  NANDN U30218 ( .A(n32483), .B(n29699), .Z(n29701) );
  XOR U30219 ( .A(a[115]), .B(b[19]), .Z(n30076) );
  NANDN U30220 ( .A(n32823), .B(n30076), .Z(n29700) );
  NAND U30221 ( .A(n29701), .B(n29700), .Z(n30007) );
  XOR U30222 ( .A(n30008), .B(n30007), .Z(n30010) );
  XOR U30223 ( .A(n30009), .B(n30010), .Z(n30044) );
  NANDN U30224 ( .A(n211), .B(n29702), .Z(n29704) );
  XOR U30225 ( .A(b[47]), .B(a[87]), .Z(n30079) );
  NANDN U30226 ( .A(n37172), .B(n30079), .Z(n29703) );
  AND U30227 ( .A(n29704), .B(n29703), .Z(n29932) );
  NANDN U30228 ( .A(n212), .B(n29705), .Z(n29707) );
  XOR U30229 ( .A(b[49]), .B(a[85]), .Z(n29921) );
  NANDN U30230 ( .A(n37432), .B(n29921), .Z(n29706) );
  AND U30231 ( .A(n29707), .B(n29706), .Z(n29931) );
  NANDN U30232 ( .A(n32996), .B(n29708), .Z(n29710) );
  XOR U30233 ( .A(a[113]), .B(b[21]), .Z(n30073) );
  NANDN U30234 ( .A(n33271), .B(n30073), .Z(n29709) );
  NAND U30235 ( .A(n29710), .B(n29709), .Z(n29930) );
  XOR U30236 ( .A(n29931), .B(n29930), .Z(n29933) );
  XNOR U30237 ( .A(n29932), .B(n29933), .Z(n30043) );
  XNOR U30238 ( .A(n30044), .B(n30043), .Z(n30046) );
  NANDN U30239 ( .A(n29712), .B(n29711), .Z(n29716) );
  OR U30240 ( .A(n29714), .B(n29713), .Z(n29715) );
  AND U30241 ( .A(n29716), .B(n29715), .Z(n30045) );
  XOR U30242 ( .A(n30046), .B(n30045), .Z(n30137) );
  NANDN U30243 ( .A(n29718), .B(n29717), .Z(n29722) );
  OR U30244 ( .A(n29720), .B(n29719), .Z(n29721) );
  AND U30245 ( .A(n29722), .B(n29721), .Z(n30136) );
  XNOR U30246 ( .A(n30137), .B(n30136), .Z(n30139) );
  XOR U30247 ( .A(n30138), .B(n30139), .Z(n30140) );
  NANDN U30248 ( .A(n38247), .B(n29723), .Z(n29725) );
  XOR U30249 ( .A(b[61]), .B(a[73]), .Z(n30094) );
  NANDN U30250 ( .A(n38248), .B(n30094), .Z(n29724) );
  AND U30251 ( .A(n29725), .B(n29724), .Z(n30022) );
  NANDN U30252 ( .A(n38278), .B(n29726), .Z(n29728) );
  XOR U30253 ( .A(b[63]), .B(a[71]), .Z(n30097) );
  NANDN U30254 ( .A(n38279), .B(n30097), .Z(n29727) );
  AND U30255 ( .A(n29728), .B(n29727), .Z(n30020) );
  NANDN U30256 ( .A(n36210), .B(n29729), .Z(n29731) );
  XOR U30257 ( .A(b[39]), .B(a[95]), .Z(n29918) );
  NANDN U30258 ( .A(n36347), .B(n29918), .Z(n29730) );
  NAND U30259 ( .A(n29731), .B(n29730), .Z(n30019) );
  XNOR U30260 ( .A(n30020), .B(n30019), .Z(n30021) );
  XOR U30261 ( .A(n30022), .B(n30021), .Z(n29967) );
  NANDN U30262 ( .A(n38090), .B(n29732), .Z(n29734) );
  XOR U30263 ( .A(b[59]), .B(a[75]), .Z(n29912) );
  NANDN U30264 ( .A(n38130), .B(n29912), .Z(n29733) );
  AND U30265 ( .A(n29734), .B(n29733), .Z(n29938) );
  XNOR U30266 ( .A(a[127]), .B(b[7]), .Z(n30002) );
  OR U30267 ( .A(n30002), .B(n29735), .Z(n29738) );
  NAND U30268 ( .A(n30003), .B(n29736), .Z(n29737) );
  AND U30269 ( .A(n29738), .B(n29737), .Z(n29937) );
  NANDN U30270 ( .A(n35260), .B(n29739), .Z(n29741) );
  XOR U30271 ( .A(a[101]), .B(b[33]), .Z(n30064) );
  NANDN U30272 ( .A(n35456), .B(n30064), .Z(n29740) );
  NAND U30273 ( .A(n29741), .B(n29740), .Z(n29936) );
  XOR U30274 ( .A(n29937), .B(n29936), .Z(n29939) );
  XNOR U30275 ( .A(n29938), .B(n29939), .Z(n29966) );
  XOR U30276 ( .A(n29967), .B(n29966), .Z(n29969) );
  NANDN U30277 ( .A(n29743), .B(n29742), .Z(n29747) );
  OR U30278 ( .A(n29745), .B(n29744), .Z(n29746) );
  AND U30279 ( .A(n29747), .B(n29746), .Z(n29968) );
  XOR U30280 ( .A(n29969), .B(n29968), .Z(n30031) );
  NANDN U30281 ( .A(n29749), .B(n29748), .Z(n29753) );
  OR U30282 ( .A(n29751), .B(n29750), .Z(n29752) );
  NAND U30283 ( .A(n29753), .B(n29752), .Z(n30032) );
  XNOR U30284 ( .A(n30031), .B(n30032), .Z(n30034) );
  NANDN U30285 ( .A(n31055), .B(n29754), .Z(n29756) );
  XOR U30286 ( .A(a[121]), .B(b[13]), .Z(n29954) );
  NANDN U30287 ( .A(n31293), .B(n29954), .Z(n29755) );
  AND U30288 ( .A(n29756), .B(n29755), .Z(n30111) );
  NANDN U30289 ( .A(n30482), .B(n29757), .Z(n29759) );
  XOR U30290 ( .A(a[123]), .B(b[11]), .Z(n29915) );
  NANDN U30291 ( .A(n30891), .B(n29915), .Z(n29758) );
  AND U30292 ( .A(n29759), .B(n29758), .Z(n30110) );
  NANDN U30293 ( .A(n34909), .B(n29760), .Z(n29762) );
  XOR U30294 ( .A(a[103]), .B(b[31]), .Z(n29993) );
  NANDN U30295 ( .A(n35145), .B(n29993), .Z(n29761) );
  NAND U30296 ( .A(n29762), .B(n29761), .Z(n30109) );
  XOR U30297 ( .A(n30110), .B(n30109), .Z(n30112) );
  XOR U30298 ( .A(n30111), .B(n30112), .Z(n30038) );
  NANDN U30299 ( .A(n29763), .B(n32544), .Z(n29765) );
  XOR U30300 ( .A(a[117]), .B(b[17]), .Z(n30049) );
  NANDN U30301 ( .A(n32292), .B(n30049), .Z(n29764) );
  AND U30302 ( .A(n29765), .B(n29764), .Z(n30069) );
  NANDN U30303 ( .A(n31536), .B(n29766), .Z(n29768) );
  XOR U30304 ( .A(a[119]), .B(b[15]), .Z(n30052) );
  NANDN U30305 ( .A(n31925), .B(n30052), .Z(n29767) );
  AND U30306 ( .A(n29768), .B(n29767), .Z(n30068) );
  NANDN U30307 ( .A(n37705), .B(n29769), .Z(n29771) );
  XOR U30308 ( .A(b[53]), .B(a[81]), .Z(n30058) );
  NANDN U30309 ( .A(n37778), .B(n30058), .Z(n29770) );
  NAND U30310 ( .A(n29771), .B(n29770), .Z(n30067) );
  XOR U30311 ( .A(n30068), .B(n30067), .Z(n30070) );
  XNOR U30312 ( .A(n30069), .B(n30070), .Z(n30037) );
  XNOR U30313 ( .A(n30038), .B(n30037), .Z(n30039) );
  NANDN U30314 ( .A(n29773), .B(n29772), .Z(n29777) );
  OR U30315 ( .A(n29775), .B(n29774), .Z(n29776) );
  NAND U30316 ( .A(n29777), .B(n29776), .Z(n30040) );
  XNOR U30317 ( .A(n30039), .B(n30040), .Z(n30033) );
  XOR U30318 ( .A(n30034), .B(n30033), .Z(n30133) );
  NAND U30319 ( .A(n29779), .B(n29778), .Z(n29783) );
  NAND U30320 ( .A(n29781), .B(n29780), .Z(n29782) );
  AND U30321 ( .A(n29783), .B(n29782), .Z(n30131) );
  NANDN U30322 ( .A(n29785), .B(n29784), .Z(n29789) );
  OR U30323 ( .A(n29787), .B(n29786), .Z(n29788) );
  AND U30324 ( .A(n29789), .B(n29788), .Z(n29975) );
  NANDN U30325 ( .A(n36991), .B(n29790), .Z(n29792) );
  XOR U30326 ( .A(b[45]), .B(a[89]), .Z(n29945) );
  NANDN U30327 ( .A(n37083), .B(n29945), .Z(n29791) );
  AND U30328 ( .A(n29792), .B(n29791), .Z(n29963) );
  NANDN U30329 ( .A(n33875), .B(n29793), .Z(n29795) );
  XOR U30330 ( .A(a[109]), .B(b[25]), .Z(n29948) );
  NANDN U30331 ( .A(n33994), .B(n29948), .Z(n29794) );
  AND U30332 ( .A(n29795), .B(n29794), .Z(n29961) );
  NANDN U30333 ( .A(n33866), .B(n29796), .Z(n29798) );
  XOR U30334 ( .A(a[111]), .B(b[23]), .Z(n29927) );
  NANDN U30335 ( .A(n33644), .B(n29927), .Z(n29797) );
  NAND U30336 ( .A(n29798), .B(n29797), .Z(n29960) );
  XNOR U30337 ( .A(n29961), .B(n29960), .Z(n29962) );
  XOR U30338 ( .A(n29963), .B(n29962), .Z(n29973) );
  NANDN U30339 ( .A(n210), .B(n29799), .Z(n29801) );
  XOR U30340 ( .A(a[125]), .B(b[9]), .Z(n29999) );
  NANDN U30341 ( .A(n30267), .B(n29999), .Z(n29800) );
  AND U30342 ( .A(n29801), .B(n29800), .Z(n30015) );
  NANDN U30343 ( .A(n37974), .B(n29802), .Z(n29804) );
  XOR U30344 ( .A(b[57]), .B(a[77]), .Z(n29951) );
  NANDN U30345 ( .A(n38031), .B(n29951), .Z(n29803) );
  AND U30346 ( .A(n29804), .B(n29803), .Z(n30014) );
  NANDN U30347 ( .A(n36480), .B(n29805), .Z(n29807) );
  XOR U30348 ( .A(b[41]), .B(a[93]), .Z(n30100) );
  NANDN U30349 ( .A(n36594), .B(n30100), .Z(n29806) );
  NAND U30350 ( .A(n29807), .B(n29806), .Z(n30013) );
  XOR U30351 ( .A(n30014), .B(n30013), .Z(n30016) );
  XNOR U30352 ( .A(n30015), .B(n30016), .Z(n29972) );
  XOR U30353 ( .A(n29973), .B(n29972), .Z(n29974) );
  XOR U30354 ( .A(n29975), .B(n29974), .Z(n29981) );
  NANDN U30355 ( .A(n29809), .B(n29808), .Z(n29813) );
  OR U30356 ( .A(n29811), .B(n29810), .Z(n29812) );
  AND U30357 ( .A(n29813), .B(n29812), .Z(n29979) );
  NANDN U30358 ( .A(n29815), .B(n29814), .Z(n29819) );
  OR U30359 ( .A(n29817), .B(n29816), .Z(n29818) );
  NAND U30360 ( .A(n29819), .B(n29818), .Z(n29978) );
  XNOR U30361 ( .A(n29979), .B(n29978), .Z(n29980) );
  XNOR U30362 ( .A(n29981), .B(n29980), .Z(n30130) );
  XNOR U30363 ( .A(n30131), .B(n30130), .Z(n30132) );
  XOR U30364 ( .A(n30133), .B(n30132), .Z(n30141) );
  XNOR U30365 ( .A(n30140), .B(n30141), .Z(n30142) );
  XOR U30366 ( .A(n30143), .B(n30142), .Z(n30147) );
  NANDN U30367 ( .A(n29821), .B(n29820), .Z(n29825) );
  NAND U30368 ( .A(n29823), .B(n29822), .Z(n29824) );
  AND U30369 ( .A(n29825), .B(n29824), .Z(n30126) );
  NANDN U30370 ( .A(n29827), .B(n29826), .Z(n29831) );
  NAND U30371 ( .A(n29829), .B(n29828), .Z(n29830) );
  AND U30372 ( .A(n29831), .B(n29830), .Z(n30125) );
  NANDN U30373 ( .A(n29833), .B(n29832), .Z(n29837) );
  OR U30374 ( .A(n29835), .B(n29834), .Z(n29836) );
  AND U30375 ( .A(n29837), .B(n29836), .Z(n30124) );
  XOR U30376 ( .A(n30125), .B(n30124), .Z(n30127) );
  XOR U30377 ( .A(n30126), .B(n30127), .Z(n30120) );
  NANDN U30378 ( .A(n29839), .B(n29838), .Z(n29843) );
  NAND U30379 ( .A(n29841), .B(n29840), .Z(n29842) );
  AND U30380 ( .A(n29843), .B(n29842), .Z(n30119) );
  NANDN U30381 ( .A(n29845), .B(n29844), .Z(n29849) );
  NAND U30382 ( .A(n29847), .B(n29846), .Z(n29848) );
  AND U30383 ( .A(n29849), .B(n29848), .Z(n30026) );
  NANDN U30384 ( .A(n29851), .B(n29850), .Z(n29855) );
  NAND U30385 ( .A(n29853), .B(n29852), .Z(n29854) );
  NAND U30386 ( .A(n29855), .B(n29854), .Z(n30025) );
  XNOR U30387 ( .A(n30026), .B(n30025), .Z(n30028) );
  NANDN U30388 ( .A(n29857), .B(n29856), .Z(n29861) );
  NAND U30389 ( .A(n29859), .B(n29858), .Z(n29860) );
  AND U30390 ( .A(n29861), .B(n29860), .Z(n30027) );
  XNOR U30391 ( .A(n30028), .B(n30027), .Z(n30118) );
  XOR U30392 ( .A(n30119), .B(n30118), .Z(n30121) );
  XNOR U30393 ( .A(n30120), .B(n30121), .Z(n30146) );
  XNOR U30394 ( .A(n30147), .B(n30146), .Z(n30148) );
  NANDN U30395 ( .A(n29863), .B(n29862), .Z(n29867) );
  NANDN U30396 ( .A(n29865), .B(n29864), .Z(n29866) );
  NAND U30397 ( .A(n29867), .B(n29866), .Z(n30149) );
  XNOR U30398 ( .A(n30148), .B(n30149), .Z(n29908) );
  XOR U30399 ( .A(n29909), .B(n29908), .Z(n29902) );
  NANDN U30400 ( .A(n29869), .B(n29868), .Z(n29873) );
  NANDN U30401 ( .A(n29871), .B(n29870), .Z(n29872) );
  AND U30402 ( .A(n29873), .B(n29872), .Z(n29901) );
  NANDN U30403 ( .A(n29875), .B(n29874), .Z(n29879) );
  NAND U30404 ( .A(n29877), .B(n29876), .Z(n29878) );
  AND U30405 ( .A(n29879), .B(n29878), .Z(n29900) );
  XOR U30406 ( .A(n29901), .B(n29900), .Z(n29903) );
  XOR U30407 ( .A(n29902), .B(n29903), .Z(n29895) );
  NANDN U30408 ( .A(n29881), .B(n29880), .Z(n29885) );
  NANDN U30409 ( .A(n29883), .B(n29882), .Z(n29884) );
  AND U30410 ( .A(n29885), .B(n29884), .Z(n29894) );
  XOR U30411 ( .A(n29895), .B(n29894), .Z(n29897) );
  XNOR U30412 ( .A(n29896), .B(n29897), .Z(n29888) );
  XOR U30413 ( .A(n29889), .B(n29888), .Z(n29891) );
  XNOR U30414 ( .A(n29890), .B(n29891), .Z(n29886) );
  XOR U30415 ( .A(n29887), .B(n29886), .Z(c[197]) );
  AND U30416 ( .A(n29887), .B(n29886), .Z(n30159) );
  NANDN U30417 ( .A(n29889), .B(n29888), .Z(n29893) );
  OR U30418 ( .A(n29891), .B(n29890), .Z(n29892) );
  AND U30419 ( .A(n29893), .B(n29892), .Z(n30162) );
  NANDN U30420 ( .A(n29895), .B(n29894), .Z(n29899) );
  NANDN U30421 ( .A(n29897), .B(n29896), .Z(n29898) );
  AND U30422 ( .A(n29899), .B(n29898), .Z(n30161) );
  NANDN U30423 ( .A(n29901), .B(n29900), .Z(n29905) );
  OR U30424 ( .A(n29903), .B(n29902), .Z(n29904) );
  AND U30425 ( .A(n29905), .B(n29904), .Z(n30168) );
  NANDN U30426 ( .A(n29907), .B(n29906), .Z(n29911) );
  NAND U30427 ( .A(n29909), .B(n29908), .Z(n29910) );
  AND U30428 ( .A(n29911), .B(n29910), .Z(n30167) );
  NANDN U30429 ( .A(n38090), .B(n29912), .Z(n29914) );
  XOR U30430 ( .A(b[59]), .B(a[76]), .Z(n30264) );
  NANDN U30431 ( .A(n38130), .B(n30264), .Z(n29913) );
  AND U30432 ( .A(n29914), .B(n29913), .Z(n30367) );
  NANDN U30433 ( .A(n30482), .B(n29915), .Z(n29917) );
  XOR U30434 ( .A(a[124]), .B(b[11]), .Z(n30347) );
  NANDN U30435 ( .A(n30891), .B(n30347), .Z(n29916) );
  AND U30436 ( .A(n29917), .B(n29916), .Z(n30366) );
  NANDN U30437 ( .A(n36210), .B(n29918), .Z(n29920) );
  XOR U30438 ( .A(b[39]), .B(a[96]), .Z(n30313) );
  NANDN U30439 ( .A(n36347), .B(n30313), .Z(n29919) );
  NAND U30440 ( .A(n29920), .B(n29919), .Z(n30365) );
  XOR U30441 ( .A(n30366), .B(n30365), .Z(n30368) );
  XOR U30442 ( .A(n30367), .B(n30368), .Z(n30185) );
  NANDN U30443 ( .A(n212), .B(n29921), .Z(n29923) );
  XOR U30444 ( .A(b[49]), .B(a[86]), .Z(n30277) );
  NANDN U30445 ( .A(n37432), .B(n30277), .Z(n29922) );
  AND U30446 ( .A(n29923), .B(n29922), .Z(n30340) );
  NANDN U30447 ( .A(n37526), .B(n29924), .Z(n29926) );
  XOR U30448 ( .A(b[51]), .B(a[84]), .Z(n30241) );
  NANDN U30449 ( .A(n37605), .B(n30241), .Z(n29925) );
  AND U30450 ( .A(n29926), .B(n29925), .Z(n30339) );
  NANDN U30451 ( .A(n33866), .B(n29927), .Z(n29929) );
  XOR U30452 ( .A(a[112]), .B(b[23]), .Z(n30220) );
  NANDN U30453 ( .A(n33644), .B(n30220), .Z(n29928) );
  NAND U30454 ( .A(n29929), .B(n29928), .Z(n30338) );
  XOR U30455 ( .A(n30339), .B(n30338), .Z(n30341) );
  XNOR U30456 ( .A(n30340), .B(n30341), .Z(n30184) );
  XNOR U30457 ( .A(n30185), .B(n30184), .Z(n30186) );
  NANDN U30458 ( .A(n29931), .B(n29930), .Z(n29935) );
  OR U30459 ( .A(n29933), .B(n29932), .Z(n29934) );
  NAND U30460 ( .A(n29935), .B(n29934), .Z(n30187) );
  XNOR U30461 ( .A(n30186), .B(n30187), .Z(n30202) );
  NANDN U30462 ( .A(n29937), .B(n29936), .Z(n29941) );
  OR U30463 ( .A(n29939), .B(n29938), .Z(n29940) );
  NAND U30464 ( .A(n29941), .B(n29940), .Z(n30203) );
  XNOR U30465 ( .A(n30202), .B(n30203), .Z(n30204) );
  NANDN U30466 ( .A(n35611), .B(n29942), .Z(n29944) );
  XOR U30467 ( .A(b[35]), .B(a[100]), .Z(n30356) );
  NANDN U30468 ( .A(n35801), .B(n30356), .Z(n29943) );
  AND U30469 ( .A(n29944), .B(n29943), .Z(n30285) );
  NANDN U30470 ( .A(n36991), .B(n29945), .Z(n29947) );
  XOR U30471 ( .A(b[45]), .B(a[90]), .Z(n30304) );
  NANDN U30472 ( .A(n37083), .B(n30304), .Z(n29946) );
  AND U30473 ( .A(n29947), .B(n29946), .Z(n30284) );
  NANDN U30474 ( .A(n33875), .B(n29948), .Z(n29950) );
  XOR U30475 ( .A(a[110]), .B(b[25]), .Z(n30232) );
  NANDN U30476 ( .A(n33994), .B(n30232), .Z(n29949) );
  NAND U30477 ( .A(n29950), .B(n29949), .Z(n30283) );
  XOR U30478 ( .A(n30284), .B(n30283), .Z(n30286) );
  XOR U30479 ( .A(n30285), .B(n30286), .Z(n30333) );
  NANDN U30480 ( .A(n37974), .B(n29951), .Z(n29953) );
  XOR U30481 ( .A(b[57]), .B(a[78]), .Z(n30344) );
  NANDN U30482 ( .A(n38031), .B(n30344), .Z(n29952) );
  AND U30483 ( .A(n29953), .B(n29952), .Z(n30328) );
  NANDN U30484 ( .A(n31055), .B(n29954), .Z(n29956) );
  XOR U30485 ( .A(a[122]), .B(b[13]), .Z(n30238) );
  NANDN U30486 ( .A(n31293), .B(n30238), .Z(n29955) );
  AND U30487 ( .A(n29956), .B(n29955), .Z(n30327) );
  NANDN U30488 ( .A(n35936), .B(n29957), .Z(n29959) );
  XOR U30489 ( .A(b[37]), .B(a[98]), .Z(n30316) );
  NANDN U30490 ( .A(n36047), .B(n30316), .Z(n29958) );
  NAND U30491 ( .A(n29959), .B(n29958), .Z(n30326) );
  XOR U30492 ( .A(n30327), .B(n30326), .Z(n30329) );
  XNOR U30493 ( .A(n30328), .B(n30329), .Z(n30332) );
  XNOR U30494 ( .A(n30333), .B(n30332), .Z(n30334) );
  NANDN U30495 ( .A(n29961), .B(n29960), .Z(n29965) );
  NANDN U30496 ( .A(n29963), .B(n29962), .Z(n29964) );
  NAND U30497 ( .A(n29965), .B(n29964), .Z(n30335) );
  XOR U30498 ( .A(n30334), .B(n30335), .Z(n30205) );
  XNOR U30499 ( .A(n30204), .B(n30205), .Z(n30386) );
  NAND U30500 ( .A(n29967), .B(n29966), .Z(n29971) );
  NAND U30501 ( .A(n29969), .B(n29968), .Z(n29970) );
  AND U30502 ( .A(n29971), .B(n29970), .Z(n30384) );
  NAND U30503 ( .A(n29973), .B(n29972), .Z(n29977) );
  NAND U30504 ( .A(n29975), .B(n29974), .Z(n29976) );
  NAND U30505 ( .A(n29977), .B(n29976), .Z(n30383) );
  XNOR U30506 ( .A(n30384), .B(n30383), .Z(n30385) );
  XOR U30507 ( .A(n30386), .B(n30385), .Z(n30378) );
  NANDN U30508 ( .A(n29979), .B(n29978), .Z(n29983) );
  NANDN U30509 ( .A(n29981), .B(n29980), .Z(n29982) );
  AND U30510 ( .A(n29983), .B(n29982), .Z(n30392) );
  NAND U30511 ( .A(n29985), .B(n29984), .Z(n29989) );
  NAND U30512 ( .A(n29987), .B(n29986), .Z(n29988) );
  AND U30513 ( .A(n29989), .B(n29988), .Z(n30389) );
  NANDN U30514 ( .A(n34634), .B(n29990), .Z(n29992) );
  XOR U30515 ( .A(a[106]), .B(b[29]), .Z(n30229) );
  NANDN U30516 ( .A(n34722), .B(n30229), .Z(n29991) );
  AND U30517 ( .A(n29992), .B(n29991), .Z(n30256) );
  NANDN U30518 ( .A(n34909), .B(n29993), .Z(n29995) );
  XOR U30519 ( .A(a[104]), .B(b[31]), .Z(n30301) );
  NANDN U30520 ( .A(n35145), .B(n30301), .Z(n29994) );
  AND U30521 ( .A(n29995), .B(n29994), .Z(n30254) );
  NANDN U30522 ( .A(n34223), .B(n29996), .Z(n29998) );
  XOR U30523 ( .A(a[108]), .B(b[27]), .Z(n30226) );
  NANDN U30524 ( .A(n34458), .B(n30226), .Z(n29997) );
  NAND U30525 ( .A(n29998), .B(n29997), .Z(n30253) );
  XNOR U30526 ( .A(n30254), .B(n30253), .Z(n30255) );
  XOR U30527 ( .A(n30256), .B(n30255), .Z(n30215) );
  NANDN U30528 ( .A(n210), .B(n29999), .Z(n30001) );
  XOR U30529 ( .A(a[126]), .B(b[9]), .Z(n30268) );
  NANDN U30530 ( .A(n30267), .B(n30268), .Z(n30000) );
  AND U30531 ( .A(n30001), .B(n30000), .Z(n30261) );
  NAND U30532 ( .A(b[63]), .B(a[70]), .Z(n30319) );
  ANDN U30533 ( .B(n30003), .A(n30002), .Z(n30006) );
  NAND U30534 ( .A(b[7]), .B(n30004), .Z(n30005) );
  NANDN U30535 ( .A(n30006), .B(n30005), .Z(n30259) );
  XOR U30536 ( .A(n30319), .B(n30259), .Z(n30260) );
  XOR U30537 ( .A(n30261), .B(n30260), .Z(n30214) );
  XOR U30538 ( .A(n30215), .B(n30214), .Z(n30217) );
  NANDN U30539 ( .A(n30008), .B(n30007), .Z(n30012) );
  OR U30540 ( .A(n30010), .B(n30009), .Z(n30011) );
  AND U30541 ( .A(n30012), .B(n30011), .Z(n30216) );
  XOR U30542 ( .A(n30217), .B(n30216), .Z(n30199) );
  NANDN U30543 ( .A(n30014), .B(n30013), .Z(n30018) );
  OR U30544 ( .A(n30016), .B(n30015), .Z(n30017) );
  AND U30545 ( .A(n30018), .B(n30017), .Z(n30197) );
  NANDN U30546 ( .A(n30020), .B(n30019), .Z(n30024) );
  NANDN U30547 ( .A(n30022), .B(n30021), .Z(n30023) );
  NAND U30548 ( .A(n30024), .B(n30023), .Z(n30196) );
  XNOR U30549 ( .A(n30197), .B(n30196), .Z(n30198) );
  XOR U30550 ( .A(n30199), .B(n30198), .Z(n30390) );
  XNOR U30551 ( .A(n30389), .B(n30390), .Z(n30391) );
  XNOR U30552 ( .A(n30392), .B(n30391), .Z(n30377) );
  XNOR U30553 ( .A(n30378), .B(n30377), .Z(n30380) );
  NANDN U30554 ( .A(n30026), .B(n30025), .Z(n30030) );
  NAND U30555 ( .A(n30028), .B(n30027), .Z(n30029) );
  AND U30556 ( .A(n30030), .B(n30029), .Z(n30379) );
  XOR U30557 ( .A(n30380), .B(n30379), .Z(n30402) );
  NANDN U30558 ( .A(n30032), .B(n30031), .Z(n30036) );
  NAND U30559 ( .A(n30034), .B(n30033), .Z(n30035) );
  AND U30560 ( .A(n30036), .B(n30035), .Z(n30175) );
  NANDN U30561 ( .A(n30038), .B(n30037), .Z(n30042) );
  NANDN U30562 ( .A(n30040), .B(n30039), .Z(n30041) );
  AND U30563 ( .A(n30042), .B(n30041), .Z(n30178) );
  NANDN U30564 ( .A(n30044), .B(n30043), .Z(n30048) );
  NAND U30565 ( .A(n30046), .B(n30045), .Z(n30047) );
  NAND U30566 ( .A(n30048), .B(n30047), .Z(n30179) );
  XNOR U30567 ( .A(n30178), .B(n30179), .Z(n30181) );
  NANDN U30568 ( .A(n32013), .B(n30049), .Z(n30051) );
  XOR U30569 ( .A(a[118]), .B(b[17]), .Z(n30280) );
  NANDN U30570 ( .A(n32292), .B(n30280), .Z(n30050) );
  AND U30571 ( .A(n30051), .B(n30050), .Z(n30361) );
  NANDN U30572 ( .A(n31536), .B(n30052), .Z(n30054) );
  XOR U30573 ( .A(a[120]), .B(b[15]), .Z(n30235) );
  NANDN U30574 ( .A(n31925), .B(n30235), .Z(n30053) );
  AND U30575 ( .A(n30054), .B(n30053), .Z(n30360) );
  NANDN U30576 ( .A(n36742), .B(n30055), .Z(n30057) );
  XOR U30577 ( .A(b[43]), .B(a[92]), .Z(n30250) );
  NANDN U30578 ( .A(n36891), .B(n30250), .Z(n30056) );
  NAND U30579 ( .A(n30057), .B(n30056), .Z(n30359) );
  XOR U30580 ( .A(n30360), .B(n30359), .Z(n30362) );
  XOR U30581 ( .A(n30361), .B(n30362), .Z(n30191) );
  NANDN U30582 ( .A(n37705), .B(n30058), .Z(n30060) );
  XOR U30583 ( .A(b[53]), .B(a[82]), .Z(n30244) );
  NANDN U30584 ( .A(n37778), .B(n30244), .Z(n30059) );
  AND U30585 ( .A(n30060), .B(n30059), .Z(n30322) );
  NANDN U30586 ( .A(n37857), .B(n30061), .Z(n30063) );
  XOR U30587 ( .A(b[55]), .B(a[80]), .Z(n30247) );
  NANDN U30588 ( .A(n37911), .B(n30247), .Z(n30062) );
  AND U30589 ( .A(n30063), .B(n30062), .Z(n30321) );
  NANDN U30590 ( .A(n35260), .B(n30064), .Z(n30066) );
  XOR U30591 ( .A(a[102]), .B(b[33]), .Z(n30350) );
  NANDN U30592 ( .A(n35456), .B(n30350), .Z(n30065) );
  NAND U30593 ( .A(n30066), .B(n30065), .Z(n30320) );
  XOR U30594 ( .A(n30321), .B(n30320), .Z(n30323) );
  XNOR U30595 ( .A(n30322), .B(n30323), .Z(n30190) );
  XNOR U30596 ( .A(n30191), .B(n30190), .Z(n30192) );
  NANDN U30597 ( .A(n30068), .B(n30067), .Z(n30072) );
  OR U30598 ( .A(n30070), .B(n30069), .Z(n30071) );
  NAND U30599 ( .A(n30072), .B(n30071), .Z(n30193) );
  XOR U30600 ( .A(n30192), .B(n30193), .Z(n30396) );
  NANDN U30601 ( .A(n32996), .B(n30073), .Z(n30075) );
  XOR U30602 ( .A(a[114]), .B(b[21]), .Z(n30223) );
  NANDN U30603 ( .A(n33271), .B(n30223), .Z(n30074) );
  AND U30604 ( .A(n30075), .B(n30074), .Z(n30291) );
  NANDN U30605 ( .A(n32483), .B(n30076), .Z(n30078) );
  XOR U30606 ( .A(a[116]), .B(b[19]), .Z(n30307) );
  NANDN U30607 ( .A(n32823), .B(n30307), .Z(n30077) );
  AND U30608 ( .A(n30078), .B(n30077), .Z(n30290) );
  NANDN U30609 ( .A(n211), .B(n30079), .Z(n30081) );
  XOR U30610 ( .A(b[47]), .B(a[88]), .Z(n30274) );
  NANDN U30611 ( .A(n37172), .B(n30274), .Z(n30080) );
  NAND U30612 ( .A(n30081), .B(n30080), .Z(n30289) );
  XOR U30613 ( .A(n30290), .B(n30289), .Z(n30292) );
  XOR U30614 ( .A(n30291), .B(n30292), .Z(n30372) );
  NAND U30615 ( .A(n30083), .B(n30082), .Z(n30087) );
  NANDN U30616 ( .A(n30085), .B(n30084), .Z(n30086) );
  AND U30617 ( .A(n30087), .B(n30086), .Z(n30371) );
  XNOR U30618 ( .A(n30372), .B(n30371), .Z(n30374) );
  NANDN U30619 ( .A(n30089), .B(n30088), .Z(n30093) );
  NANDN U30620 ( .A(n30091), .B(n30090), .Z(n30092) );
  AND U30621 ( .A(n30093), .B(n30092), .Z(n30373) );
  XNOR U30622 ( .A(n30374), .B(n30373), .Z(n30395) );
  XOR U30623 ( .A(n30396), .B(n30395), .Z(n30398) );
  NANDN U30624 ( .A(n38247), .B(n30094), .Z(n30096) );
  XOR U30625 ( .A(b[61]), .B(a[74]), .Z(n30353) );
  NANDN U30626 ( .A(n38248), .B(n30353), .Z(n30095) );
  AND U30627 ( .A(n30096), .B(n30095), .Z(n30297) );
  NANDN U30628 ( .A(n38278), .B(n30097), .Z(n30099) );
  XOR U30629 ( .A(b[63]), .B(a[72]), .Z(n30310) );
  NANDN U30630 ( .A(n38279), .B(n30310), .Z(n30098) );
  AND U30631 ( .A(n30099), .B(n30098), .Z(n30296) );
  NANDN U30632 ( .A(n36480), .B(n30100), .Z(n30102) );
  XOR U30633 ( .A(b[41]), .B(a[94]), .Z(n30271) );
  NANDN U30634 ( .A(n36594), .B(n30271), .Z(n30101) );
  NAND U30635 ( .A(n30102), .B(n30101), .Z(n30295) );
  XOR U30636 ( .A(n30296), .B(n30295), .Z(n30298) );
  XOR U30637 ( .A(n30297), .B(n30298), .Z(n30209) );
  NANDN U30638 ( .A(n30104), .B(n30103), .Z(n30108) );
  NAND U30639 ( .A(n30106), .B(n30105), .Z(n30107) );
  AND U30640 ( .A(n30108), .B(n30107), .Z(n30208) );
  XNOR U30641 ( .A(n30209), .B(n30208), .Z(n30210) );
  NANDN U30642 ( .A(n30110), .B(n30109), .Z(n30114) );
  OR U30643 ( .A(n30112), .B(n30111), .Z(n30113) );
  NAND U30644 ( .A(n30114), .B(n30113), .Z(n30211) );
  XOR U30645 ( .A(n30210), .B(n30211), .Z(n30397) );
  XOR U30646 ( .A(n30398), .B(n30397), .Z(n30180) );
  XOR U30647 ( .A(n30181), .B(n30180), .Z(n30173) );
  XNOR U30648 ( .A(n30173), .B(n30172), .Z(n30174) );
  XNOR U30649 ( .A(n30175), .B(n30174), .Z(n30401) );
  XNOR U30650 ( .A(n30402), .B(n30401), .Z(n30403) );
  NANDN U30651 ( .A(n30119), .B(n30118), .Z(n30123) );
  OR U30652 ( .A(n30121), .B(n30120), .Z(n30122) );
  NAND U30653 ( .A(n30123), .B(n30122), .Z(n30404) );
  XNOR U30654 ( .A(n30403), .B(n30404), .Z(n30415) );
  NANDN U30655 ( .A(n30125), .B(n30124), .Z(n30129) );
  OR U30656 ( .A(n30127), .B(n30126), .Z(n30128) );
  AND U30657 ( .A(n30129), .B(n30128), .Z(n30410) );
  NANDN U30658 ( .A(n30131), .B(n30130), .Z(n30135) );
  NANDN U30659 ( .A(n30133), .B(n30132), .Z(n30134) );
  AND U30660 ( .A(n30135), .B(n30134), .Z(n30408) );
  XNOR U30661 ( .A(n30408), .B(n30407), .Z(n30409) );
  XOR U30662 ( .A(n30410), .B(n30409), .Z(n30414) );
  NANDN U30663 ( .A(n30141), .B(n30140), .Z(n30145) );
  NAND U30664 ( .A(n30143), .B(n30142), .Z(n30144) );
  AND U30665 ( .A(n30145), .B(n30144), .Z(n30413) );
  XOR U30666 ( .A(n30414), .B(n30413), .Z(n30416) );
  XNOR U30667 ( .A(n30415), .B(n30416), .Z(n30421) );
  NANDN U30668 ( .A(n30147), .B(n30146), .Z(n30151) );
  NANDN U30669 ( .A(n30149), .B(n30148), .Z(n30150) );
  AND U30670 ( .A(n30151), .B(n30150), .Z(n30420) );
  NANDN U30671 ( .A(n30153), .B(n30152), .Z(n30157) );
  NANDN U30672 ( .A(n30155), .B(n30154), .Z(n30156) );
  NAND U30673 ( .A(n30157), .B(n30156), .Z(n30419) );
  XOR U30674 ( .A(n30420), .B(n30419), .Z(n30422) );
  XNOR U30675 ( .A(n30421), .B(n30422), .Z(n30166) );
  XOR U30676 ( .A(n30167), .B(n30166), .Z(n30169) );
  XNOR U30677 ( .A(n30168), .B(n30169), .Z(n30160) );
  XOR U30678 ( .A(n30161), .B(n30160), .Z(n30163) );
  XNOR U30679 ( .A(n30162), .B(n30163), .Z(n30158) );
  XOR U30680 ( .A(n30159), .B(n30158), .Z(c[198]) );
  AND U30681 ( .A(n30159), .B(n30158), .Z(n30426) );
  NANDN U30682 ( .A(n30161), .B(n30160), .Z(n30165) );
  OR U30683 ( .A(n30163), .B(n30162), .Z(n30164) );
  AND U30684 ( .A(n30165), .B(n30164), .Z(n30429) );
  NANDN U30685 ( .A(n30167), .B(n30166), .Z(n30171) );
  NANDN U30686 ( .A(n30169), .B(n30168), .Z(n30170) );
  AND U30687 ( .A(n30171), .B(n30170), .Z(n30428) );
  NANDN U30688 ( .A(n30173), .B(n30172), .Z(n30177) );
  NANDN U30689 ( .A(n30175), .B(n30174), .Z(n30176) );
  AND U30690 ( .A(n30177), .B(n30176), .Z(n30453) );
  NANDN U30691 ( .A(n30179), .B(n30178), .Z(n30183) );
  NAND U30692 ( .A(n30181), .B(n30180), .Z(n30182) );
  AND U30693 ( .A(n30183), .B(n30182), .Z(n30465) );
  NANDN U30694 ( .A(n30185), .B(n30184), .Z(n30189) );
  NANDN U30695 ( .A(n30187), .B(n30186), .Z(n30188) );
  AND U30696 ( .A(n30189), .B(n30188), .Z(n30476) );
  NANDN U30697 ( .A(n30191), .B(n30190), .Z(n30195) );
  NANDN U30698 ( .A(n30193), .B(n30192), .Z(n30194) );
  NAND U30699 ( .A(n30195), .B(n30194), .Z(n30475) );
  XNOR U30700 ( .A(n30476), .B(n30475), .Z(n30478) );
  NANDN U30701 ( .A(n30197), .B(n30196), .Z(n30201) );
  NANDN U30702 ( .A(n30199), .B(n30198), .Z(n30200) );
  AND U30703 ( .A(n30201), .B(n30200), .Z(n30477) );
  XOR U30704 ( .A(n30478), .B(n30477), .Z(n30464) );
  NANDN U30705 ( .A(n30203), .B(n30202), .Z(n30207) );
  NANDN U30706 ( .A(n30205), .B(n30204), .Z(n30206) );
  AND U30707 ( .A(n30207), .B(n30206), .Z(n30463) );
  XOR U30708 ( .A(n30464), .B(n30463), .Z(n30466) );
  XOR U30709 ( .A(n30465), .B(n30466), .Z(n30452) );
  NANDN U30710 ( .A(n30209), .B(n30208), .Z(n30213) );
  NANDN U30711 ( .A(n30211), .B(n30210), .Z(n30212) );
  AND U30712 ( .A(n30213), .B(n30212), .Z(n30471) );
  NAND U30713 ( .A(n30215), .B(n30214), .Z(n30219) );
  NAND U30714 ( .A(n30217), .B(n30216), .Z(n30218) );
  AND U30715 ( .A(n30219), .B(n30218), .Z(n30470) );
  NANDN U30716 ( .A(n33866), .B(n30220), .Z(n30222) );
  XOR U30717 ( .A(a[113]), .B(b[23]), .Z(n30494) );
  NANDN U30718 ( .A(n33644), .B(n30494), .Z(n30221) );
  AND U30719 ( .A(n30222), .B(n30221), .Z(n30544) );
  NANDN U30720 ( .A(n32996), .B(n30223), .Z(n30225) );
  XOR U30721 ( .A(a[115]), .B(b[21]), .Z(n30590) );
  NANDN U30722 ( .A(n33271), .B(n30590), .Z(n30224) );
  AND U30723 ( .A(n30225), .B(n30224), .Z(n30543) );
  NANDN U30724 ( .A(n34223), .B(n30226), .Z(n30228) );
  XOR U30725 ( .A(a[109]), .B(b[27]), .Z(n30664) );
  NANDN U30726 ( .A(n34458), .B(n30664), .Z(n30227) );
  AND U30727 ( .A(n30228), .B(n30227), .Z(n30655) );
  NANDN U30728 ( .A(n34634), .B(n30229), .Z(n30231) );
  XOR U30729 ( .A(a[107]), .B(b[29]), .Z(n30566) );
  NANDN U30730 ( .A(n34722), .B(n30566), .Z(n30230) );
  AND U30731 ( .A(n30231), .B(n30230), .Z(n30653) );
  NANDN U30732 ( .A(n33875), .B(n30232), .Z(n30234) );
  XOR U30733 ( .A(a[111]), .B(b[25]), .Z(n30491) );
  NANDN U30734 ( .A(n33994), .B(n30491), .Z(n30233) );
  NAND U30735 ( .A(n30234), .B(n30233), .Z(n30652) );
  XNOR U30736 ( .A(n30653), .B(n30652), .Z(n30654) );
  XNOR U30737 ( .A(n30655), .B(n30654), .Z(n30542) );
  XOR U30738 ( .A(n30543), .B(n30542), .Z(n30545) );
  XOR U30739 ( .A(n30544), .B(n30545), .Z(n30613) );
  NANDN U30740 ( .A(n31536), .B(n30235), .Z(n30237) );
  XOR U30741 ( .A(a[121]), .B(b[15]), .Z(n30670) );
  NANDN U30742 ( .A(n31925), .B(n30670), .Z(n30236) );
  AND U30743 ( .A(n30237), .B(n30236), .Z(n30502) );
  NANDN U30744 ( .A(n31055), .B(n30238), .Z(n30240) );
  XOR U30745 ( .A(a[123]), .B(b[13]), .Z(n30584) );
  NANDN U30746 ( .A(n31293), .B(n30584), .Z(n30239) );
  AND U30747 ( .A(n30240), .B(n30239), .Z(n30501) );
  NANDN U30748 ( .A(n37526), .B(n30241), .Z(n30243) );
  XOR U30749 ( .A(b[51]), .B(a[85]), .Z(n30563) );
  NANDN U30750 ( .A(n37605), .B(n30563), .Z(n30242) );
  NAND U30751 ( .A(n30243), .B(n30242), .Z(n30500) );
  XOR U30752 ( .A(n30501), .B(n30500), .Z(n30503) );
  XOR U30753 ( .A(n30502), .B(n30503), .Z(n30612) );
  NANDN U30754 ( .A(n37705), .B(n30244), .Z(n30246) );
  XOR U30755 ( .A(b[53]), .B(a[83]), .Z(n30658) );
  NANDN U30756 ( .A(n37778), .B(n30658), .Z(n30245) );
  AND U30757 ( .A(n30246), .B(n30245), .Z(n30508) );
  NANDN U30758 ( .A(n37857), .B(n30247), .Z(n30249) );
  XOR U30759 ( .A(b[55]), .B(a[81]), .Z(n30661) );
  NANDN U30760 ( .A(n37911), .B(n30661), .Z(n30248) );
  AND U30761 ( .A(n30249), .B(n30248), .Z(n30507) );
  NANDN U30762 ( .A(n36742), .B(n30250), .Z(n30252) );
  XOR U30763 ( .A(b[43]), .B(a[93]), .Z(n30673) );
  NANDN U30764 ( .A(n36891), .B(n30673), .Z(n30251) );
  NAND U30765 ( .A(n30252), .B(n30251), .Z(n30506) );
  XOR U30766 ( .A(n30507), .B(n30506), .Z(n30509) );
  XNOR U30767 ( .A(n30508), .B(n30509), .Z(n30611) );
  XOR U30768 ( .A(n30612), .B(n30611), .Z(n30614) );
  XOR U30769 ( .A(n30613), .B(n30614), .Z(n30684) );
  NANDN U30770 ( .A(n30254), .B(n30253), .Z(n30258) );
  NANDN U30771 ( .A(n30256), .B(n30255), .Z(n30257) );
  AND U30772 ( .A(n30258), .B(n30257), .Z(n30683) );
  IV U30773 ( .A(n30319), .Z(n30571) );
  NANDN U30774 ( .A(n30571), .B(n30259), .Z(n30263) );
  NANDN U30775 ( .A(n30261), .B(n30260), .Z(n30262) );
  NAND U30776 ( .A(n30263), .B(n30262), .Z(n30682) );
  XOR U30777 ( .A(n30683), .B(n30682), .Z(n30685) );
  XNOR U30778 ( .A(n30684), .B(n30685), .Z(n30469) );
  XOR U30779 ( .A(n30470), .B(n30469), .Z(n30472) );
  XOR U30780 ( .A(n30471), .B(n30472), .Z(n30459) );
  NANDN U30781 ( .A(n38090), .B(n30264), .Z(n30266) );
  XOR U30782 ( .A(b[59]), .B(a[77]), .Z(n30581) );
  NANDN U30783 ( .A(n38130), .B(n30581), .Z(n30265) );
  AND U30784 ( .A(n30266), .B(n30265), .Z(n30556) );
  XNOR U30785 ( .A(a[127]), .B(b[9]), .Z(n30626) );
  OR U30786 ( .A(n30626), .B(n30267), .Z(n30270) );
  NAND U30787 ( .A(n30627), .B(n30268), .Z(n30269) );
  AND U30788 ( .A(n30270), .B(n30269), .Z(n30555) );
  NANDN U30789 ( .A(n36480), .B(n30271), .Z(n30273) );
  XOR U30790 ( .A(b[41]), .B(a[95]), .Z(n30587) );
  NANDN U30791 ( .A(n36594), .B(n30587), .Z(n30272) );
  NAND U30792 ( .A(n30273), .B(n30272), .Z(n30554) );
  XOR U30793 ( .A(n30555), .B(n30554), .Z(n30557) );
  XOR U30794 ( .A(n30556), .B(n30557), .Z(n30519) );
  NANDN U30795 ( .A(n211), .B(n30274), .Z(n30276) );
  XOR U30796 ( .A(b[47]), .B(a[89]), .Z(n30643) );
  NANDN U30797 ( .A(n37172), .B(n30643), .Z(n30275) );
  AND U30798 ( .A(n30276), .B(n30275), .Z(n30577) );
  NANDN U30799 ( .A(n212), .B(n30277), .Z(n30279) );
  XOR U30800 ( .A(b[49]), .B(a[87]), .Z(n30560) );
  NANDN U30801 ( .A(n37432), .B(n30560), .Z(n30278) );
  AND U30802 ( .A(n30279), .B(n30278), .Z(n30576) );
  NANDN U30803 ( .A(n32013), .B(n30280), .Z(n30282) );
  XOR U30804 ( .A(a[119]), .B(b[17]), .Z(n30667) );
  NANDN U30805 ( .A(n32292), .B(n30667), .Z(n30281) );
  NAND U30806 ( .A(n30282), .B(n30281), .Z(n30575) );
  XOR U30807 ( .A(n30576), .B(n30575), .Z(n30578) );
  XNOR U30808 ( .A(n30577), .B(n30578), .Z(n30518) );
  XNOR U30809 ( .A(n30519), .B(n30518), .Z(n30521) );
  NANDN U30810 ( .A(n30284), .B(n30283), .Z(n30288) );
  OR U30811 ( .A(n30286), .B(n30285), .Z(n30287) );
  AND U30812 ( .A(n30288), .B(n30287), .Z(n30520) );
  XOR U30813 ( .A(n30521), .B(n30520), .Z(n30678) );
  NANDN U30814 ( .A(n30290), .B(n30289), .Z(n30294) );
  OR U30815 ( .A(n30292), .B(n30291), .Z(n30293) );
  AND U30816 ( .A(n30294), .B(n30293), .Z(n30677) );
  NANDN U30817 ( .A(n30296), .B(n30295), .Z(n30300) );
  OR U30818 ( .A(n30298), .B(n30297), .Z(n30299) );
  NAND U30819 ( .A(n30300), .B(n30299), .Z(n30676) );
  XOR U30820 ( .A(n30677), .B(n30676), .Z(n30679) );
  XOR U30821 ( .A(n30678), .B(n30679), .Z(n30538) );
  NANDN U30822 ( .A(n34909), .B(n30301), .Z(n30303) );
  XOR U30823 ( .A(a[105]), .B(b[31]), .Z(n30640) );
  NANDN U30824 ( .A(n35145), .B(n30640), .Z(n30302) );
  AND U30825 ( .A(n30303), .B(n30302), .Z(n30601) );
  NANDN U30826 ( .A(n36991), .B(n30304), .Z(n30306) );
  XOR U30827 ( .A(b[45]), .B(a[91]), .Z(n30596) );
  NANDN U30828 ( .A(n37083), .B(n30596), .Z(n30305) );
  AND U30829 ( .A(n30306), .B(n30305), .Z(n30600) );
  NANDN U30830 ( .A(n32483), .B(n30307), .Z(n30309) );
  XOR U30831 ( .A(a[117]), .B(b[19]), .Z(n30593) );
  NANDN U30832 ( .A(n32823), .B(n30593), .Z(n30308) );
  NAND U30833 ( .A(n30309), .B(n30308), .Z(n30599) );
  XOR U30834 ( .A(n30600), .B(n30599), .Z(n30602) );
  XOR U30835 ( .A(n30601), .B(n30602), .Z(n30647) );
  NANDN U30836 ( .A(n38278), .B(n30310), .Z(n30312) );
  XOR U30837 ( .A(b[63]), .B(a[73]), .Z(n30623) );
  NANDN U30838 ( .A(n38279), .B(n30623), .Z(n30311) );
  AND U30839 ( .A(n30312), .B(n30311), .Z(n30618) );
  NANDN U30840 ( .A(n36210), .B(n30313), .Z(n30315) );
  XOR U30841 ( .A(b[39]), .B(a[97]), .Z(n30488) );
  NANDN U30842 ( .A(n36347), .B(n30488), .Z(n30314) );
  NAND U30843 ( .A(n30315), .B(n30314), .Z(n30617) );
  XNOR U30844 ( .A(n30618), .B(n30617), .Z(n30620) );
  NAND U30845 ( .A(n36238), .B(n30316), .Z(n30318) );
  XNOR U30846 ( .A(b[37]), .B(a[99]), .Z(n30637) );
  NANDN U30847 ( .A(n30637), .B(n36239), .Z(n30317) );
  NAND U30848 ( .A(n30318), .B(n30317), .Z(n30569) );
  AND U30849 ( .A(b[63]), .B(a[71]), .Z(n30570) );
  XNOR U30850 ( .A(n30569), .B(n30570), .Z(n30572) );
  XOR U30851 ( .A(n30319), .B(n30572), .Z(n30619) );
  XNOR U30852 ( .A(n30620), .B(n30619), .Z(n30646) );
  XNOR U30853 ( .A(n30647), .B(n30646), .Z(n30648) );
  NANDN U30854 ( .A(n30321), .B(n30320), .Z(n30325) );
  OR U30855 ( .A(n30323), .B(n30322), .Z(n30324) );
  NAND U30856 ( .A(n30325), .B(n30324), .Z(n30649) );
  XNOR U30857 ( .A(n30648), .B(n30649), .Z(n30536) );
  NANDN U30858 ( .A(n30327), .B(n30326), .Z(n30331) );
  OR U30859 ( .A(n30329), .B(n30328), .Z(n30330) );
  NAND U30860 ( .A(n30331), .B(n30330), .Z(n30537) );
  XOR U30861 ( .A(n30536), .B(n30537), .Z(n30539) );
  XOR U30862 ( .A(n30538), .B(n30539), .Z(n30533) );
  NANDN U30863 ( .A(n30333), .B(n30332), .Z(n30337) );
  NANDN U30864 ( .A(n30335), .B(n30334), .Z(n30336) );
  AND U30865 ( .A(n30337), .B(n30336), .Z(n30530) );
  NANDN U30866 ( .A(n30339), .B(n30338), .Z(n30343) );
  OR U30867 ( .A(n30341), .B(n30340), .Z(n30342) );
  AND U30868 ( .A(n30343), .B(n30342), .Z(n30608) );
  NANDN U30869 ( .A(n37974), .B(n30344), .Z(n30346) );
  XOR U30870 ( .A(b[57]), .B(a[79]), .Z(n30497) );
  NANDN U30871 ( .A(n38031), .B(n30497), .Z(n30345) );
  AND U30872 ( .A(n30346), .B(n30345), .Z(n30550) );
  NANDN U30873 ( .A(n30482), .B(n30347), .Z(n30349) );
  XOR U30874 ( .A(a[125]), .B(b[11]), .Z(n30481) );
  NANDN U30875 ( .A(n30891), .B(n30481), .Z(n30348) );
  AND U30876 ( .A(n30349), .B(n30348), .Z(n30549) );
  NANDN U30877 ( .A(n35260), .B(n30350), .Z(n30352) );
  XOR U30878 ( .A(a[103]), .B(b[33]), .Z(n30634) );
  NANDN U30879 ( .A(n35456), .B(n30634), .Z(n30351) );
  NAND U30880 ( .A(n30352), .B(n30351), .Z(n30548) );
  XOR U30881 ( .A(n30549), .B(n30548), .Z(n30551) );
  XOR U30882 ( .A(n30550), .B(n30551), .Z(n30606) );
  NANDN U30883 ( .A(n38247), .B(n30353), .Z(n30355) );
  XOR U30884 ( .A(b[61]), .B(a[75]), .Z(n30485) );
  NANDN U30885 ( .A(n38248), .B(n30485), .Z(n30354) );
  AND U30886 ( .A(n30355), .B(n30354), .Z(n30513) );
  NANDN U30887 ( .A(n35611), .B(n30356), .Z(n30358) );
  XOR U30888 ( .A(b[35]), .B(a[101]), .Z(n30631) );
  NANDN U30889 ( .A(n35801), .B(n30631), .Z(n30357) );
  NAND U30890 ( .A(n30358), .B(n30357), .Z(n30512) );
  XOR U30891 ( .A(n30513), .B(n30512), .Z(n30515) );
  XNOR U30892 ( .A(n30514), .B(n30515), .Z(n30605) );
  XNOR U30893 ( .A(n30606), .B(n30605), .Z(n30607) );
  XOR U30894 ( .A(n30608), .B(n30607), .Z(n30527) );
  NANDN U30895 ( .A(n30360), .B(n30359), .Z(n30364) );
  OR U30896 ( .A(n30362), .B(n30361), .Z(n30363) );
  AND U30897 ( .A(n30364), .B(n30363), .Z(n30525) );
  NANDN U30898 ( .A(n30366), .B(n30365), .Z(n30370) );
  OR U30899 ( .A(n30368), .B(n30367), .Z(n30369) );
  NAND U30900 ( .A(n30370), .B(n30369), .Z(n30524) );
  XNOR U30901 ( .A(n30525), .B(n30524), .Z(n30526) );
  XOR U30902 ( .A(n30527), .B(n30526), .Z(n30531) );
  XNOR U30903 ( .A(n30530), .B(n30531), .Z(n30532) );
  XNOR U30904 ( .A(n30533), .B(n30532), .Z(n30457) );
  NANDN U30905 ( .A(n30372), .B(n30371), .Z(n30376) );
  NAND U30906 ( .A(n30374), .B(n30373), .Z(n30375) );
  NAND U30907 ( .A(n30376), .B(n30375), .Z(n30458) );
  XOR U30908 ( .A(n30457), .B(n30458), .Z(n30460) );
  XNOR U30909 ( .A(n30459), .B(n30460), .Z(n30451) );
  XOR U30910 ( .A(n30452), .B(n30451), .Z(n30454) );
  XOR U30911 ( .A(n30453), .B(n30454), .Z(n30690) );
  NANDN U30912 ( .A(n30378), .B(n30377), .Z(n30382) );
  NAND U30913 ( .A(n30380), .B(n30379), .Z(n30381) );
  AND U30914 ( .A(n30382), .B(n30381), .Z(n30689) );
  NANDN U30915 ( .A(n30384), .B(n30383), .Z(n30388) );
  NAND U30916 ( .A(n30386), .B(n30385), .Z(n30387) );
  AND U30917 ( .A(n30388), .B(n30387), .Z(n30447) );
  NANDN U30918 ( .A(n30390), .B(n30389), .Z(n30394) );
  NANDN U30919 ( .A(n30392), .B(n30391), .Z(n30393) );
  AND U30920 ( .A(n30394), .B(n30393), .Z(n30446) );
  NAND U30921 ( .A(n30396), .B(n30395), .Z(n30400) );
  NAND U30922 ( .A(n30398), .B(n30397), .Z(n30399) );
  NAND U30923 ( .A(n30400), .B(n30399), .Z(n30445) );
  XOR U30924 ( .A(n30446), .B(n30445), .Z(n30448) );
  XNOR U30925 ( .A(n30447), .B(n30448), .Z(n30688) );
  XOR U30926 ( .A(n30689), .B(n30688), .Z(n30691) );
  XOR U30927 ( .A(n30690), .B(n30691), .Z(n30441) );
  NANDN U30928 ( .A(n30402), .B(n30401), .Z(n30406) );
  NANDN U30929 ( .A(n30404), .B(n30403), .Z(n30405) );
  AND U30930 ( .A(n30406), .B(n30405), .Z(n30440) );
  NANDN U30931 ( .A(n30408), .B(n30407), .Z(n30412) );
  NAND U30932 ( .A(n30410), .B(n30409), .Z(n30411) );
  AND U30933 ( .A(n30412), .B(n30411), .Z(n30439) );
  XOR U30934 ( .A(n30440), .B(n30439), .Z(n30442) );
  XOR U30935 ( .A(n30441), .B(n30442), .Z(n30434) );
  NANDN U30936 ( .A(n30414), .B(n30413), .Z(n30418) );
  NANDN U30937 ( .A(n30416), .B(n30415), .Z(n30417) );
  AND U30938 ( .A(n30418), .B(n30417), .Z(n30433) );
  XNOR U30939 ( .A(n30434), .B(n30433), .Z(n30436) );
  NANDN U30940 ( .A(n30420), .B(n30419), .Z(n30424) );
  NANDN U30941 ( .A(n30422), .B(n30421), .Z(n30423) );
  AND U30942 ( .A(n30424), .B(n30423), .Z(n30435) );
  XNOR U30943 ( .A(n30436), .B(n30435), .Z(n30427) );
  XOR U30944 ( .A(n30428), .B(n30427), .Z(n30430) );
  XNOR U30945 ( .A(n30429), .B(n30430), .Z(n30425) );
  XOR U30946 ( .A(n30426), .B(n30425), .Z(c[199]) );
  AND U30947 ( .A(n30426), .B(n30425), .Z(n30695) );
  NANDN U30948 ( .A(n30428), .B(n30427), .Z(n30432) );
  OR U30949 ( .A(n30430), .B(n30429), .Z(n30431) );
  AND U30950 ( .A(n30432), .B(n30431), .Z(n30698) );
  NANDN U30951 ( .A(n30434), .B(n30433), .Z(n30438) );
  NAND U30952 ( .A(n30436), .B(n30435), .Z(n30437) );
  AND U30953 ( .A(n30438), .B(n30437), .Z(n30696) );
  NANDN U30954 ( .A(n30440), .B(n30439), .Z(n30444) );
  OR U30955 ( .A(n30442), .B(n30441), .Z(n30443) );
  AND U30956 ( .A(n30444), .B(n30443), .Z(n30705) );
  NANDN U30957 ( .A(n30446), .B(n30445), .Z(n30450) );
  NANDN U30958 ( .A(n30448), .B(n30447), .Z(n30449) );
  AND U30959 ( .A(n30450), .B(n30449), .Z(n30709) );
  NANDN U30960 ( .A(n30452), .B(n30451), .Z(n30456) );
  OR U30961 ( .A(n30454), .B(n30453), .Z(n30455) );
  AND U30962 ( .A(n30456), .B(n30455), .Z(n30708) );
  XNOR U30963 ( .A(n30709), .B(n30708), .Z(n30711) );
  NANDN U30964 ( .A(n30458), .B(n30457), .Z(n30462) );
  OR U30965 ( .A(n30460), .B(n30459), .Z(n30461) );
  AND U30966 ( .A(n30462), .B(n30461), .Z(n30948) );
  NANDN U30967 ( .A(n30464), .B(n30463), .Z(n30468) );
  OR U30968 ( .A(n30466), .B(n30465), .Z(n30467) );
  NAND U30969 ( .A(n30468), .B(n30467), .Z(n30947) );
  XNOR U30970 ( .A(n30948), .B(n30947), .Z(n30949) );
  NANDN U30971 ( .A(n30470), .B(n30469), .Z(n30474) );
  OR U30972 ( .A(n30472), .B(n30471), .Z(n30473) );
  AND U30973 ( .A(n30474), .B(n30473), .Z(n30722) );
  NANDN U30974 ( .A(n30476), .B(n30475), .Z(n30480) );
  NAND U30975 ( .A(n30478), .B(n30477), .Z(n30479) );
  AND U30976 ( .A(n30480), .B(n30479), .Z(n30721) );
  NANDN U30977 ( .A(n30482), .B(n30481), .Z(n30484) );
  XOR U30978 ( .A(a[126]), .B(b[11]), .Z(n30892) );
  NANDN U30979 ( .A(n30891), .B(n30892), .Z(n30483) );
  AND U30980 ( .A(n30484), .B(n30483), .Z(n30789) );
  NANDN U30981 ( .A(n38247), .B(n30485), .Z(n30487) );
  XOR U30982 ( .A(b[61]), .B(a[76]), .Z(n30762) );
  NANDN U30983 ( .A(n38248), .B(n30762), .Z(n30486) );
  AND U30984 ( .A(n30487), .B(n30486), .Z(n30787) );
  NANDN U30985 ( .A(n36210), .B(n30488), .Z(n30490) );
  XOR U30986 ( .A(b[39]), .B(a[98]), .Z(n30895) );
  NANDN U30987 ( .A(n36347), .B(n30895), .Z(n30489) );
  NAND U30988 ( .A(n30490), .B(n30489), .Z(n30786) );
  XNOR U30989 ( .A(n30787), .B(n30786), .Z(n30788) );
  XOR U30990 ( .A(n30789), .B(n30788), .Z(n30874) );
  NANDN U30991 ( .A(n33875), .B(n30491), .Z(n30493) );
  XOR U30992 ( .A(a[112]), .B(b[25]), .Z(n30846) );
  NANDN U30993 ( .A(n33994), .B(n30846), .Z(n30492) );
  AND U30994 ( .A(n30493), .B(n30492), .Z(n30869) );
  NANDN U30995 ( .A(n33866), .B(n30494), .Z(n30496) );
  XOR U30996 ( .A(a[114]), .B(b[23]), .Z(n30840) );
  NANDN U30997 ( .A(n33644), .B(n30840), .Z(n30495) );
  AND U30998 ( .A(n30496), .B(n30495), .Z(n30868) );
  NANDN U30999 ( .A(n37974), .B(n30497), .Z(n30499) );
  XOR U31000 ( .A(b[57]), .B(a[80]), .Z(n30849) );
  NANDN U31001 ( .A(n38031), .B(n30849), .Z(n30498) );
  NAND U31002 ( .A(n30499), .B(n30498), .Z(n30867) );
  XOR U31003 ( .A(n30868), .B(n30867), .Z(n30870) );
  XNOR U31004 ( .A(n30869), .B(n30870), .Z(n30873) );
  XOR U31005 ( .A(n30874), .B(n30873), .Z(n30876) );
  NANDN U31006 ( .A(n30501), .B(n30500), .Z(n30505) );
  OR U31007 ( .A(n30503), .B(n30502), .Z(n30504) );
  AND U31008 ( .A(n30505), .B(n30504), .Z(n30875) );
  XOR U31009 ( .A(n30876), .B(n30875), .Z(n30937) );
  NANDN U31010 ( .A(n30507), .B(n30506), .Z(n30511) );
  OR U31011 ( .A(n30509), .B(n30508), .Z(n30510) );
  AND U31012 ( .A(n30511), .B(n30510), .Z(n30936) );
  NANDN U31013 ( .A(n30513), .B(n30512), .Z(n30517) );
  OR U31014 ( .A(n30515), .B(n30514), .Z(n30516) );
  NAND U31015 ( .A(n30517), .B(n30516), .Z(n30935) );
  XOR U31016 ( .A(n30936), .B(n30935), .Z(n30938) );
  XOR U31017 ( .A(n30937), .B(n30938), .Z(n30799) );
  NANDN U31018 ( .A(n30519), .B(n30518), .Z(n30523) );
  NAND U31019 ( .A(n30521), .B(n30520), .Z(n30522) );
  NAND U31020 ( .A(n30523), .B(n30522), .Z(n30798) );
  XNOR U31021 ( .A(n30799), .B(n30798), .Z(n30800) );
  NANDN U31022 ( .A(n30525), .B(n30524), .Z(n30529) );
  NANDN U31023 ( .A(n30527), .B(n30526), .Z(n30528) );
  NAND U31024 ( .A(n30529), .B(n30528), .Z(n30801) );
  XNOR U31025 ( .A(n30800), .B(n30801), .Z(n30720) );
  XOR U31026 ( .A(n30721), .B(n30720), .Z(n30723) );
  XOR U31027 ( .A(n30722), .B(n30723), .Z(n30717) );
  NANDN U31028 ( .A(n30531), .B(n30530), .Z(n30535) );
  NANDN U31029 ( .A(n30533), .B(n30532), .Z(n30534) );
  AND U31030 ( .A(n30535), .B(n30534), .Z(n30715) );
  NANDN U31031 ( .A(n30537), .B(n30536), .Z(n30541) );
  OR U31032 ( .A(n30539), .B(n30538), .Z(n30540) );
  AND U31033 ( .A(n30541), .B(n30540), .Z(n30726) );
  NANDN U31034 ( .A(n30543), .B(n30542), .Z(n30547) );
  OR U31035 ( .A(n30545), .B(n30544), .Z(n30546) );
  AND U31036 ( .A(n30547), .B(n30546), .Z(n30746) );
  NANDN U31037 ( .A(n30549), .B(n30548), .Z(n30553) );
  OR U31038 ( .A(n30551), .B(n30550), .Z(n30552) );
  AND U31039 ( .A(n30553), .B(n30552), .Z(n30745) );
  NANDN U31040 ( .A(n30555), .B(n30554), .Z(n30559) );
  OR U31041 ( .A(n30557), .B(n30556), .Z(n30558) );
  NAND U31042 ( .A(n30559), .B(n30558), .Z(n30744) );
  XOR U31043 ( .A(n30745), .B(n30744), .Z(n30747) );
  XOR U31044 ( .A(n30746), .B(n30747), .Z(n30806) );
  NANDN U31045 ( .A(n212), .B(n30560), .Z(n30562) );
  XOR U31046 ( .A(b[49]), .B(a[88]), .Z(n30861) );
  NANDN U31047 ( .A(n37432), .B(n30861), .Z(n30561) );
  AND U31048 ( .A(n30562), .B(n30561), .Z(n30931) );
  NANDN U31049 ( .A(n37526), .B(n30563), .Z(n30565) );
  XOR U31050 ( .A(b[51]), .B(a[86]), .Z(n30864) );
  NANDN U31051 ( .A(n37605), .B(n30864), .Z(n30564) );
  AND U31052 ( .A(n30565), .B(n30564), .Z(n30930) );
  NANDN U31053 ( .A(n34634), .B(n30566), .Z(n30568) );
  XOR U31054 ( .A(a[108]), .B(b[29]), .Z(n30828) );
  NANDN U31055 ( .A(n34722), .B(n30828), .Z(n30567) );
  NAND U31056 ( .A(n30568), .B(n30567), .Z(n30929) );
  XOR U31057 ( .A(n30930), .B(n30929), .Z(n30932) );
  XOR U31058 ( .A(n30931), .B(n30932), .Z(n30906) );
  NAND U31059 ( .A(n30570), .B(n30569), .Z(n30574) );
  NANDN U31060 ( .A(n30572), .B(n30571), .Z(n30573) );
  AND U31061 ( .A(n30574), .B(n30573), .Z(n30905) );
  XNOR U31062 ( .A(n30906), .B(n30905), .Z(n30907) );
  NANDN U31063 ( .A(n30576), .B(n30575), .Z(n30580) );
  OR U31064 ( .A(n30578), .B(n30577), .Z(n30579) );
  NAND U31065 ( .A(n30580), .B(n30579), .Z(n30908) );
  XNOR U31066 ( .A(n30907), .B(n30908), .Z(n30804) );
  NANDN U31067 ( .A(n38090), .B(n30581), .Z(n30583) );
  XOR U31068 ( .A(b[59]), .B(a[78]), .Z(n30852) );
  NANDN U31069 ( .A(n38130), .B(n30852), .Z(n30582) );
  AND U31070 ( .A(n30583), .B(n30582), .Z(n30824) );
  NANDN U31071 ( .A(n31055), .B(n30584), .Z(n30586) );
  XOR U31072 ( .A(a[124]), .B(b[13]), .Z(n30911) );
  NANDN U31073 ( .A(n31293), .B(n30911), .Z(n30585) );
  AND U31074 ( .A(n30586), .B(n30585), .Z(n30823) );
  NANDN U31075 ( .A(n36480), .B(n30587), .Z(n30589) );
  XOR U31076 ( .A(b[41]), .B(a[96]), .Z(n30917) );
  NANDN U31077 ( .A(n36594), .B(n30917), .Z(n30588) );
  NAND U31078 ( .A(n30589), .B(n30588), .Z(n30822) );
  XOR U31079 ( .A(n30823), .B(n30822), .Z(n30825) );
  XOR U31080 ( .A(n30824), .B(n30825), .Z(n30880) );
  NANDN U31081 ( .A(n32996), .B(n30590), .Z(n30592) );
  XOR U31082 ( .A(a[116]), .B(b[21]), .Z(n30843) );
  NANDN U31083 ( .A(n33271), .B(n30843), .Z(n30591) );
  AND U31084 ( .A(n30592), .B(n30591), .Z(n30782) );
  NANDN U31085 ( .A(n32483), .B(n30593), .Z(n30595) );
  XOR U31086 ( .A(a[118]), .B(b[19]), .Z(n30834) );
  NANDN U31087 ( .A(n32823), .B(n30834), .Z(n30594) );
  AND U31088 ( .A(n30595), .B(n30594), .Z(n30781) );
  NANDN U31089 ( .A(n36991), .B(n30596), .Z(n30598) );
  XOR U31090 ( .A(b[45]), .B(a[92]), .Z(n30926) );
  NANDN U31091 ( .A(n37083), .B(n30926), .Z(n30597) );
  NAND U31092 ( .A(n30598), .B(n30597), .Z(n30780) );
  XOR U31093 ( .A(n30781), .B(n30780), .Z(n30783) );
  XNOR U31094 ( .A(n30782), .B(n30783), .Z(n30879) );
  XNOR U31095 ( .A(n30880), .B(n30879), .Z(n30881) );
  NANDN U31096 ( .A(n30600), .B(n30599), .Z(n30604) );
  OR U31097 ( .A(n30602), .B(n30601), .Z(n30603) );
  NAND U31098 ( .A(n30604), .B(n30603), .Z(n30882) );
  XOR U31099 ( .A(n30881), .B(n30882), .Z(n30805) );
  XOR U31100 ( .A(n30804), .B(n30805), .Z(n30807) );
  XOR U31101 ( .A(n30806), .B(n30807), .Z(n30741) );
  NANDN U31102 ( .A(n30606), .B(n30605), .Z(n30610) );
  NAND U31103 ( .A(n30608), .B(n30607), .Z(n30609) );
  AND U31104 ( .A(n30610), .B(n30609), .Z(n30738) );
  NANDN U31105 ( .A(n30612), .B(n30611), .Z(n30616) );
  OR U31106 ( .A(n30614), .B(n30613), .Z(n30615) );
  NAND U31107 ( .A(n30616), .B(n30615), .Z(n30739) );
  XNOR U31108 ( .A(n30738), .B(n30739), .Z(n30740) );
  XOR U31109 ( .A(n30741), .B(n30740), .Z(n30727) );
  XNOR U31110 ( .A(n30726), .B(n30727), .Z(n30728) );
  NANDN U31111 ( .A(n30618), .B(n30617), .Z(n30622) );
  NAND U31112 ( .A(n30620), .B(n30619), .Z(n30621) );
  AND U31113 ( .A(n30622), .B(n30621), .Z(n30942) );
  NANDN U31114 ( .A(n38278), .B(n30623), .Z(n30625) );
  XOR U31115 ( .A(b[63]), .B(a[74]), .Z(n30914) );
  NANDN U31116 ( .A(n38279), .B(n30914), .Z(n30624) );
  AND U31117 ( .A(n30625), .B(n30624), .Z(n30902) );
  NAND U31118 ( .A(b[63]), .B(a[72]), .Z(n30899) );
  ANDN U31119 ( .B(n30627), .A(n30626), .Z(n30630) );
  NAND U31120 ( .A(b[9]), .B(n30628), .Z(n30629) );
  NANDN U31121 ( .A(n30630), .B(n30629), .Z(n30900) );
  XOR U31122 ( .A(n30899), .B(n30900), .Z(n30901) );
  XNOR U31123 ( .A(n30902), .B(n30901), .Z(n30941) );
  XNOR U31124 ( .A(n30942), .B(n30941), .Z(n30944) );
  NANDN U31125 ( .A(n35611), .B(n30631), .Z(n30633) );
  XOR U31126 ( .A(a[102]), .B(b[35]), .Z(n30774) );
  NANDN U31127 ( .A(n35801), .B(n30774), .Z(n30632) );
  AND U31128 ( .A(n30633), .B(n30632), .Z(n30813) );
  NANDN U31129 ( .A(n35260), .B(n30634), .Z(n30636) );
  XOR U31130 ( .A(a[104]), .B(b[33]), .Z(n30771) );
  NANDN U31131 ( .A(n35456), .B(n30771), .Z(n30635) );
  AND U31132 ( .A(n30636), .B(n30635), .Z(n30811) );
  NANDN U31133 ( .A(n30637), .B(n36238), .Z(n30639) );
  XNOR U31134 ( .A(b[37]), .B(a[100]), .Z(n30855) );
  NANDN U31135 ( .A(n30855), .B(n36239), .Z(n30638) );
  NAND U31136 ( .A(n30639), .B(n30638), .Z(n30887) );
  NAND U31137 ( .A(n35309), .B(n30640), .Z(n30642) );
  XNOR U31138 ( .A(a[106]), .B(b[31]), .Z(n30831) );
  NANDN U31139 ( .A(n30831), .B(n35310), .Z(n30641) );
  NAND U31140 ( .A(n30642), .B(n30641), .Z(n30886) );
  NANDN U31141 ( .A(n211), .B(n30643), .Z(n30645) );
  XOR U31142 ( .A(b[47]), .B(a[90]), .Z(n30858) );
  NANDN U31143 ( .A(n37172), .B(n30858), .Z(n30644) );
  NAND U31144 ( .A(n30645), .B(n30644), .Z(n30885) );
  XOR U31145 ( .A(n30886), .B(n30885), .Z(n30888) );
  XOR U31146 ( .A(n30887), .B(n30888), .Z(n30810) );
  XNOR U31147 ( .A(n30811), .B(n30810), .Z(n30812) );
  XNOR U31148 ( .A(n30813), .B(n30812), .Z(n30943) );
  XOR U31149 ( .A(n30944), .B(n30943), .Z(n30734) );
  NANDN U31150 ( .A(n30647), .B(n30646), .Z(n30651) );
  NANDN U31151 ( .A(n30649), .B(n30648), .Z(n30650) );
  AND U31152 ( .A(n30651), .B(n30650), .Z(n30733) );
  NANDN U31153 ( .A(n30653), .B(n30652), .Z(n30657) );
  NANDN U31154 ( .A(n30655), .B(n30654), .Z(n30656) );
  AND U31155 ( .A(n30657), .B(n30656), .Z(n30752) );
  NANDN U31156 ( .A(n37705), .B(n30658), .Z(n30660) );
  XOR U31157 ( .A(b[53]), .B(a[84]), .Z(n30920) );
  NANDN U31158 ( .A(n37778), .B(n30920), .Z(n30659) );
  AND U31159 ( .A(n30660), .B(n30659), .Z(n30758) );
  NANDN U31160 ( .A(n37857), .B(n30661), .Z(n30663) );
  XOR U31161 ( .A(b[55]), .B(a[82]), .Z(n30923) );
  NANDN U31162 ( .A(n37911), .B(n30923), .Z(n30662) );
  AND U31163 ( .A(n30663), .B(n30662), .Z(n30757) );
  NANDN U31164 ( .A(n34223), .B(n30664), .Z(n30666) );
  XOR U31165 ( .A(a[110]), .B(b[27]), .Z(n30837) );
  NANDN U31166 ( .A(n34458), .B(n30837), .Z(n30665) );
  NAND U31167 ( .A(n30666), .B(n30665), .Z(n30756) );
  XOR U31168 ( .A(n30757), .B(n30756), .Z(n30759) );
  XOR U31169 ( .A(n30758), .B(n30759), .Z(n30751) );
  NANDN U31170 ( .A(n32013), .B(n30667), .Z(n30669) );
  XOR U31171 ( .A(a[120]), .B(b[17]), .Z(n30777) );
  NANDN U31172 ( .A(n32292), .B(n30777), .Z(n30668) );
  AND U31173 ( .A(n30669), .B(n30668), .Z(n30818) );
  NANDN U31174 ( .A(n31536), .B(n30670), .Z(n30672) );
  XOR U31175 ( .A(a[122]), .B(b[15]), .Z(n30765) );
  NANDN U31176 ( .A(n31925), .B(n30765), .Z(n30671) );
  AND U31177 ( .A(n30672), .B(n30671), .Z(n30817) );
  NANDN U31178 ( .A(n36742), .B(n30673), .Z(n30675) );
  XOR U31179 ( .A(b[43]), .B(a[94]), .Z(n30768) );
  NANDN U31180 ( .A(n36891), .B(n30768), .Z(n30674) );
  NAND U31181 ( .A(n30675), .B(n30674), .Z(n30816) );
  XOR U31182 ( .A(n30817), .B(n30816), .Z(n30819) );
  XNOR U31183 ( .A(n30818), .B(n30819), .Z(n30750) );
  XOR U31184 ( .A(n30751), .B(n30750), .Z(n30753) );
  XNOR U31185 ( .A(n30752), .B(n30753), .Z(n30732) );
  XOR U31186 ( .A(n30733), .B(n30732), .Z(n30735) );
  XOR U31187 ( .A(n30734), .B(n30735), .Z(n30795) );
  NANDN U31188 ( .A(n30677), .B(n30676), .Z(n30681) );
  OR U31189 ( .A(n30679), .B(n30678), .Z(n30680) );
  AND U31190 ( .A(n30681), .B(n30680), .Z(n30793) );
  NANDN U31191 ( .A(n30683), .B(n30682), .Z(n30687) );
  OR U31192 ( .A(n30685), .B(n30684), .Z(n30686) );
  NAND U31193 ( .A(n30687), .B(n30686), .Z(n30792) );
  XNOR U31194 ( .A(n30793), .B(n30792), .Z(n30794) );
  XOR U31195 ( .A(n30795), .B(n30794), .Z(n30729) );
  XNOR U31196 ( .A(n30728), .B(n30729), .Z(n30714) );
  XNOR U31197 ( .A(n30715), .B(n30714), .Z(n30716) );
  XOR U31198 ( .A(n30717), .B(n30716), .Z(n30950) );
  XNOR U31199 ( .A(n30949), .B(n30950), .Z(n30710) );
  XOR U31200 ( .A(n30711), .B(n30710), .Z(n30703) );
  NANDN U31201 ( .A(n30689), .B(n30688), .Z(n30693) );
  OR U31202 ( .A(n30691), .B(n30690), .Z(n30692) );
  AND U31203 ( .A(n30693), .B(n30692), .Z(n30702) );
  XNOR U31204 ( .A(n30703), .B(n30702), .Z(n30704) );
  XOR U31205 ( .A(n30705), .B(n30704), .Z(n30697) );
  XOR U31206 ( .A(n30696), .B(n30697), .Z(n30699) );
  XNOR U31207 ( .A(n30698), .B(n30699), .Z(n30694) );
  XOR U31208 ( .A(n30695), .B(n30694), .Z(c[200]) );
  AND U31209 ( .A(n30695), .B(n30694), .Z(n30954) );
  NANDN U31210 ( .A(n30697), .B(n30696), .Z(n30701) );
  OR U31211 ( .A(n30699), .B(n30698), .Z(n30700) );
  AND U31212 ( .A(n30701), .B(n30700), .Z(n30957) );
  NANDN U31213 ( .A(n30703), .B(n30702), .Z(n30707) );
  NANDN U31214 ( .A(n30705), .B(n30704), .Z(n30706) );
  AND U31215 ( .A(n30707), .B(n30706), .Z(n30956) );
  NANDN U31216 ( .A(n30709), .B(n30708), .Z(n30713) );
  NAND U31217 ( .A(n30711), .B(n30710), .Z(n30712) );
  AND U31218 ( .A(n30713), .B(n30712), .Z(n30963) );
  NANDN U31219 ( .A(n30715), .B(n30714), .Z(n30719) );
  NANDN U31220 ( .A(n30717), .B(n30716), .Z(n30718) );
  AND U31221 ( .A(n30719), .B(n30718), .Z(n30968) );
  NANDN U31222 ( .A(n30721), .B(n30720), .Z(n30725) );
  OR U31223 ( .A(n30723), .B(n30722), .Z(n30724) );
  AND U31224 ( .A(n30725), .B(n30724), .Z(n30967) );
  XNOR U31225 ( .A(n30968), .B(n30967), .Z(n30970) );
  NANDN U31226 ( .A(n30727), .B(n30726), .Z(n30731) );
  NANDN U31227 ( .A(n30729), .B(n30728), .Z(n30730) );
  AND U31228 ( .A(n30731), .B(n30730), .Z(n30974) );
  NANDN U31229 ( .A(n30733), .B(n30732), .Z(n30737) );
  OR U31230 ( .A(n30735), .B(n30734), .Z(n30736) );
  AND U31231 ( .A(n30737), .B(n30736), .Z(n31203) );
  NANDN U31232 ( .A(n30739), .B(n30738), .Z(n30743) );
  NANDN U31233 ( .A(n30741), .B(n30740), .Z(n30742) );
  AND U31234 ( .A(n30743), .B(n30742), .Z(n31202) );
  NANDN U31235 ( .A(n30745), .B(n30744), .Z(n30749) );
  OR U31236 ( .A(n30747), .B(n30746), .Z(n30748) );
  AND U31237 ( .A(n30749), .B(n30748), .Z(n31051) );
  NANDN U31238 ( .A(n30751), .B(n30750), .Z(n30755) );
  NANDN U31239 ( .A(n30753), .B(n30752), .Z(n30754) );
  AND U31240 ( .A(n30755), .B(n30754), .Z(n31048) );
  NANDN U31241 ( .A(n30757), .B(n30756), .Z(n30761) );
  OR U31242 ( .A(n30759), .B(n30758), .Z(n30760) );
  AND U31243 ( .A(n30761), .B(n30760), .Z(n31117) );
  NANDN U31244 ( .A(n38247), .B(n30762), .Z(n30764) );
  XOR U31245 ( .A(b[61]), .B(a[77]), .Z(n31063) );
  NANDN U31246 ( .A(n38248), .B(n31063), .Z(n30763) );
  AND U31247 ( .A(n30764), .B(n30763), .Z(n31006) );
  NANDN U31248 ( .A(n31536), .B(n30765), .Z(n30767) );
  XOR U31249 ( .A(a[123]), .B(b[15]), .Z(n31087) );
  NANDN U31250 ( .A(n31925), .B(n31087), .Z(n30766) );
  AND U31251 ( .A(n30767), .B(n30766), .Z(n31004) );
  NANDN U31252 ( .A(n36742), .B(n30768), .Z(n30770) );
  XOR U31253 ( .A(b[43]), .B(a[95]), .Z(n31099) );
  NANDN U31254 ( .A(n36891), .B(n31099), .Z(n30769) );
  NAND U31255 ( .A(n30770), .B(n30769), .Z(n31003) );
  XNOR U31256 ( .A(n31004), .B(n31003), .Z(n31005) );
  XOR U31257 ( .A(n31006), .B(n31005), .Z(n31115) );
  NANDN U31258 ( .A(n35260), .B(n30771), .Z(n30773) );
  XOR U31259 ( .A(a[105]), .B(b[33]), .Z(n31186) );
  NANDN U31260 ( .A(n35456), .B(n31186), .Z(n30772) );
  AND U31261 ( .A(n30773), .B(n30772), .Z(n31104) );
  NANDN U31262 ( .A(n35611), .B(n30774), .Z(n30776) );
  XOR U31263 ( .A(a[103]), .B(b[35]), .Z(n31189) );
  NANDN U31264 ( .A(n35801), .B(n31189), .Z(n30775) );
  AND U31265 ( .A(n30776), .B(n30775), .Z(n31103) );
  NANDN U31266 ( .A(n32013), .B(n30777), .Z(n30779) );
  XOR U31267 ( .A(a[121]), .B(b[17]), .Z(n31192) );
  NANDN U31268 ( .A(n32292), .B(n31192), .Z(n30778) );
  NAND U31269 ( .A(n30779), .B(n30778), .Z(n31102) );
  XOR U31270 ( .A(n31103), .B(n31102), .Z(n31105) );
  XNOR U31271 ( .A(n31104), .B(n31105), .Z(n31114) );
  XOR U31272 ( .A(n31115), .B(n31114), .Z(n31116) );
  XOR U31273 ( .A(n31117), .B(n31116), .Z(n31129) );
  NANDN U31274 ( .A(n30781), .B(n30780), .Z(n30785) );
  OR U31275 ( .A(n30783), .B(n30782), .Z(n30784) );
  AND U31276 ( .A(n30785), .B(n30784), .Z(n31127) );
  NANDN U31277 ( .A(n30787), .B(n30786), .Z(n30791) );
  NANDN U31278 ( .A(n30789), .B(n30788), .Z(n30790) );
  NAND U31279 ( .A(n30791), .B(n30790), .Z(n31126) );
  XNOR U31280 ( .A(n31127), .B(n31126), .Z(n31128) );
  XOR U31281 ( .A(n31129), .B(n31128), .Z(n31049) );
  XNOR U31282 ( .A(n31048), .B(n31049), .Z(n31050) );
  XNOR U31283 ( .A(n31051), .B(n31050), .Z(n31201) );
  XOR U31284 ( .A(n31202), .B(n31201), .Z(n31204) );
  XNOR U31285 ( .A(n31203), .B(n31204), .Z(n30973) );
  XNOR U31286 ( .A(n30974), .B(n30973), .Z(n30975) );
  NANDN U31287 ( .A(n30793), .B(n30792), .Z(n30797) );
  NANDN U31288 ( .A(n30795), .B(n30794), .Z(n30796) );
  AND U31289 ( .A(n30797), .B(n30796), .Z(n31210) );
  NANDN U31290 ( .A(n30799), .B(n30798), .Z(n30803) );
  NANDN U31291 ( .A(n30801), .B(n30800), .Z(n30802) );
  AND U31292 ( .A(n30803), .B(n30802), .Z(n31207) );
  NANDN U31293 ( .A(n30805), .B(n30804), .Z(n30809) );
  OR U31294 ( .A(n30807), .B(n30806), .Z(n30808) );
  AND U31295 ( .A(n30809), .B(n30808), .Z(n30979) );
  NANDN U31296 ( .A(n30811), .B(n30810), .Z(n30815) );
  NANDN U31297 ( .A(n30813), .B(n30812), .Z(n30814) );
  AND U31298 ( .A(n30815), .B(n30814), .Z(n30993) );
  NANDN U31299 ( .A(n30817), .B(n30816), .Z(n30821) );
  OR U31300 ( .A(n30819), .B(n30818), .Z(n30820) );
  AND U31301 ( .A(n30821), .B(n30820), .Z(n30992) );
  NANDN U31302 ( .A(n30823), .B(n30822), .Z(n30827) );
  OR U31303 ( .A(n30825), .B(n30824), .Z(n30826) );
  NAND U31304 ( .A(n30827), .B(n30826), .Z(n30991) );
  XOR U31305 ( .A(n30992), .B(n30991), .Z(n30994) );
  XOR U31306 ( .A(n30993), .B(n30994), .Z(n31122) );
  NANDN U31307 ( .A(n34634), .B(n30828), .Z(n30830) );
  XOR U31308 ( .A(a[109]), .B(b[29]), .Z(n31138) );
  NANDN U31309 ( .A(n34722), .B(n31138), .Z(n30829) );
  AND U31310 ( .A(n30830), .B(n30829), .Z(n31074) );
  NANDN U31311 ( .A(n30831), .B(n35309), .Z(n30833) );
  XOR U31312 ( .A(a[107]), .B(b[31]), .Z(n31141) );
  NANDN U31313 ( .A(n35145), .B(n31141), .Z(n30832) );
  AND U31314 ( .A(n30833), .B(n30832), .Z(n31073) );
  NANDN U31315 ( .A(n32483), .B(n30834), .Z(n30836) );
  XOR U31316 ( .A(a[119]), .B(b[19]), .Z(n31144) );
  NANDN U31317 ( .A(n32823), .B(n31144), .Z(n30835) );
  NAND U31318 ( .A(n30836), .B(n30835), .Z(n31072) );
  XOR U31319 ( .A(n31073), .B(n31072), .Z(n31075) );
  XOR U31320 ( .A(n31074), .B(n31075), .Z(n31174) );
  NANDN U31321 ( .A(n34223), .B(n30837), .Z(n30839) );
  XOR U31322 ( .A(a[111]), .B(b[27]), .Z(n31156) );
  NANDN U31323 ( .A(n34458), .B(n31156), .Z(n30838) );
  AND U31324 ( .A(n30839), .B(n30838), .Z(n31017) );
  NANDN U31325 ( .A(n33866), .B(n30840), .Z(n30842) );
  XOR U31326 ( .A(a[115]), .B(b[23]), .Z(n31150) );
  NANDN U31327 ( .A(n33644), .B(n31150), .Z(n30841) );
  AND U31328 ( .A(n30842), .B(n30841), .Z(n31016) );
  NANDN U31329 ( .A(n32996), .B(n30843), .Z(n30845) );
  XOR U31330 ( .A(a[117]), .B(b[21]), .Z(n31153) );
  NANDN U31331 ( .A(n33271), .B(n31153), .Z(n30844) );
  NAND U31332 ( .A(n30845), .B(n30844), .Z(n31015) );
  XOR U31333 ( .A(n31016), .B(n31015), .Z(n31018) );
  XOR U31334 ( .A(n31017), .B(n31018), .Z(n31172) );
  NAND U31335 ( .A(n34297), .B(n30846), .Z(n30848) );
  XNOR U31336 ( .A(a[113]), .B(b[25]), .Z(n31147) );
  NANDN U31337 ( .A(n31147), .B(n34298), .Z(n30847) );
  AND U31338 ( .A(n30848), .B(n30847), .Z(n31171) );
  XNOR U31339 ( .A(n31172), .B(n31171), .Z(n31173) );
  XNOR U31340 ( .A(n31174), .B(n31173), .Z(n31120) );
  NANDN U31341 ( .A(n37974), .B(n30849), .Z(n30851) );
  XOR U31342 ( .A(b[57]), .B(a[81]), .Z(n31027) );
  NANDN U31343 ( .A(n38031), .B(n31027), .Z(n30850) );
  AND U31344 ( .A(n30851), .B(n30850), .Z(n31080) );
  NANDN U31345 ( .A(n38090), .B(n30852), .Z(n30854) );
  XOR U31346 ( .A(b[59]), .B(a[79]), .Z(n31030) );
  NANDN U31347 ( .A(n38130), .B(n31030), .Z(n30853) );
  AND U31348 ( .A(n30854), .B(n30853), .Z(n31079) );
  NANDN U31349 ( .A(n30855), .B(n36238), .Z(n30857) );
  XOR U31350 ( .A(b[37]), .B(a[101]), .Z(n31090) );
  NANDN U31351 ( .A(n36047), .B(n31090), .Z(n30856) );
  NAND U31352 ( .A(n30857), .B(n30856), .Z(n31078) );
  XOR U31353 ( .A(n31079), .B(n31078), .Z(n31081) );
  XOR U31354 ( .A(n31080), .B(n31081), .Z(n31109) );
  NANDN U31355 ( .A(n211), .B(n30858), .Z(n30860) );
  XOR U31356 ( .A(b[47]), .B(a[91]), .Z(n31180) );
  NANDN U31357 ( .A(n37172), .B(n31180), .Z(n30859) );
  AND U31358 ( .A(n30860), .B(n30859), .Z(n31197) );
  NANDN U31359 ( .A(n212), .B(n30861), .Z(n30863) );
  XOR U31360 ( .A(b[49]), .B(a[89]), .Z(n31183) );
  NANDN U31361 ( .A(n37432), .B(n31183), .Z(n30862) );
  AND U31362 ( .A(n30863), .B(n30862), .Z(n31196) );
  NANDN U31363 ( .A(n37526), .B(n30864), .Z(n30866) );
  XOR U31364 ( .A(b[51]), .B(a[87]), .Z(n31093) );
  NANDN U31365 ( .A(n37605), .B(n31093), .Z(n30865) );
  NAND U31366 ( .A(n30866), .B(n30865), .Z(n31195) );
  XOR U31367 ( .A(n31196), .B(n31195), .Z(n31198) );
  XNOR U31368 ( .A(n31197), .B(n31198), .Z(n31108) );
  XNOR U31369 ( .A(n31109), .B(n31108), .Z(n31110) );
  NANDN U31370 ( .A(n30868), .B(n30867), .Z(n30872) );
  OR U31371 ( .A(n30870), .B(n30869), .Z(n30871) );
  NAND U31372 ( .A(n30872), .B(n30871), .Z(n31111) );
  XOR U31373 ( .A(n31110), .B(n31111), .Z(n31121) );
  XOR U31374 ( .A(n31120), .B(n31121), .Z(n31123) );
  XOR U31375 ( .A(n31122), .B(n31123), .Z(n31039) );
  NAND U31376 ( .A(n30874), .B(n30873), .Z(n30878) );
  NAND U31377 ( .A(n30876), .B(n30875), .Z(n30877) );
  AND U31378 ( .A(n30878), .B(n30877), .Z(n31036) );
  NANDN U31379 ( .A(n30880), .B(n30879), .Z(n30884) );
  NANDN U31380 ( .A(n30882), .B(n30881), .Z(n30883) );
  NAND U31381 ( .A(n30884), .B(n30883), .Z(n31037) );
  XNOR U31382 ( .A(n31036), .B(n31037), .Z(n31038) );
  XOR U31383 ( .A(n31039), .B(n31038), .Z(n30980) );
  XNOR U31384 ( .A(n30979), .B(n30980), .Z(n30981) );
  NAND U31385 ( .A(n30886), .B(n30885), .Z(n30890) );
  NAND U31386 ( .A(n30888), .B(n30887), .Z(n30889) );
  AND U31387 ( .A(n30890), .B(n30889), .Z(n31134) );
  XNOR U31388 ( .A(a[127]), .B(b[11]), .Z(n31058) );
  OR U31389 ( .A(n31058), .B(n30891), .Z(n30894) );
  NAND U31390 ( .A(n31059), .B(n30892), .Z(n30893) );
  AND U31391 ( .A(n30894), .B(n30893), .Z(n31166) );
  NANDN U31392 ( .A(n36210), .B(n30895), .Z(n30897) );
  XOR U31393 ( .A(b[39]), .B(a[99]), .Z(n31033) );
  NANDN U31394 ( .A(n36347), .B(n31033), .Z(n30896) );
  NAND U31395 ( .A(n30897), .B(n30896), .Z(n31165) );
  XNOR U31396 ( .A(n31166), .B(n31165), .Z(n31168) );
  IV U31397 ( .A(n30898), .Z(n31022) );
  AND U31398 ( .A(b[63]), .B(a[73]), .Z(n31021) );
  XOR U31399 ( .A(n31022), .B(n31021), .Z(n31023) );
  XOR U31400 ( .A(n30899), .B(n31023), .Z(n31167) );
  XOR U31401 ( .A(n31168), .B(n31167), .Z(n31133) );
  IV U31402 ( .A(n30899), .Z(n31024) );
  NANDN U31403 ( .A(n31024), .B(n30900), .Z(n30904) );
  NANDN U31404 ( .A(n30902), .B(n30901), .Z(n30903) );
  AND U31405 ( .A(n30904), .B(n30903), .Z(n31132) );
  XOR U31406 ( .A(n31133), .B(n31132), .Z(n31135) );
  XNOR U31407 ( .A(n31134), .B(n31135), .Z(n30988) );
  NANDN U31408 ( .A(n30906), .B(n30905), .Z(n30910) );
  NANDN U31409 ( .A(n30908), .B(n30907), .Z(n30909) );
  NAND U31410 ( .A(n30910), .B(n30909), .Z(n30985) );
  NANDN U31411 ( .A(n31055), .B(n30911), .Z(n30913) );
  XOR U31412 ( .A(a[125]), .B(b[13]), .Z(n31054) );
  NANDN U31413 ( .A(n31293), .B(n31054), .Z(n30912) );
  AND U31414 ( .A(n30913), .B(n30912), .Z(n31011) );
  NANDN U31415 ( .A(n38278), .B(n30914), .Z(n30916) );
  XOR U31416 ( .A(b[63]), .B(a[75]), .Z(n31066) );
  NANDN U31417 ( .A(n38279), .B(n31066), .Z(n30915) );
  AND U31418 ( .A(n30916), .B(n30915), .Z(n31010) );
  NANDN U31419 ( .A(n36480), .B(n30917), .Z(n30919) );
  XOR U31420 ( .A(b[41]), .B(a[97]), .Z(n31069) );
  NANDN U31421 ( .A(n36594), .B(n31069), .Z(n30918) );
  NAND U31422 ( .A(n30919), .B(n30918), .Z(n31009) );
  XOR U31423 ( .A(n31010), .B(n31009), .Z(n31012) );
  XOR U31424 ( .A(n31011), .B(n31012), .Z(n30998) );
  NANDN U31425 ( .A(n37705), .B(n30920), .Z(n30922) );
  XOR U31426 ( .A(b[53]), .B(a[85]), .Z(n31096) );
  NANDN U31427 ( .A(n37778), .B(n31096), .Z(n30921) );
  AND U31428 ( .A(n30922), .B(n30921), .Z(n31161) );
  NANDN U31429 ( .A(n37857), .B(n30923), .Z(n30925) );
  XOR U31430 ( .A(b[55]), .B(a[83]), .Z(n31084) );
  NANDN U31431 ( .A(n37911), .B(n31084), .Z(n30924) );
  AND U31432 ( .A(n30925), .B(n30924), .Z(n31160) );
  NANDN U31433 ( .A(n36991), .B(n30926), .Z(n30928) );
  XOR U31434 ( .A(b[45]), .B(a[93]), .Z(n31177) );
  NANDN U31435 ( .A(n37083), .B(n31177), .Z(n30927) );
  NAND U31436 ( .A(n30928), .B(n30927), .Z(n31159) );
  XOR U31437 ( .A(n31160), .B(n31159), .Z(n31162) );
  XNOR U31438 ( .A(n31161), .B(n31162), .Z(n30997) );
  XNOR U31439 ( .A(n30998), .B(n30997), .Z(n30999) );
  NANDN U31440 ( .A(n30930), .B(n30929), .Z(n30934) );
  OR U31441 ( .A(n30932), .B(n30931), .Z(n30933) );
  NAND U31442 ( .A(n30934), .B(n30933), .Z(n31000) );
  XNOR U31443 ( .A(n30999), .B(n31000), .Z(n30986) );
  XOR U31444 ( .A(n30985), .B(n30986), .Z(n30987) );
  XOR U31445 ( .A(n30988), .B(n30987), .Z(n31045) );
  NANDN U31446 ( .A(n30936), .B(n30935), .Z(n30940) );
  OR U31447 ( .A(n30938), .B(n30937), .Z(n30939) );
  AND U31448 ( .A(n30940), .B(n30939), .Z(n31043) );
  NANDN U31449 ( .A(n30942), .B(n30941), .Z(n30946) );
  NAND U31450 ( .A(n30944), .B(n30943), .Z(n30945) );
  NAND U31451 ( .A(n30946), .B(n30945), .Z(n31042) );
  XNOR U31452 ( .A(n31043), .B(n31042), .Z(n31044) );
  XOR U31453 ( .A(n31045), .B(n31044), .Z(n30982) );
  XOR U31454 ( .A(n30981), .B(n30982), .Z(n31208) );
  XNOR U31455 ( .A(n31207), .B(n31208), .Z(n31209) );
  XOR U31456 ( .A(n31210), .B(n31209), .Z(n30976) );
  XNOR U31457 ( .A(n30975), .B(n30976), .Z(n30969) );
  XOR U31458 ( .A(n30970), .B(n30969), .Z(n30962) );
  NANDN U31459 ( .A(n30948), .B(n30947), .Z(n30952) );
  NANDN U31460 ( .A(n30950), .B(n30949), .Z(n30951) );
  AND U31461 ( .A(n30952), .B(n30951), .Z(n30961) );
  XOR U31462 ( .A(n30962), .B(n30961), .Z(n30964) );
  XNOR U31463 ( .A(n30963), .B(n30964), .Z(n30955) );
  XOR U31464 ( .A(n30956), .B(n30955), .Z(n30958) );
  XNOR U31465 ( .A(n30957), .B(n30958), .Z(n30953) );
  XOR U31466 ( .A(n30954), .B(n30953), .Z(c[201]) );
  AND U31467 ( .A(n30954), .B(n30953), .Z(n31214) );
  NANDN U31468 ( .A(n30956), .B(n30955), .Z(n30960) );
  OR U31469 ( .A(n30958), .B(n30957), .Z(n30959) );
  AND U31470 ( .A(n30960), .B(n30959), .Z(n31217) );
  NANDN U31471 ( .A(n30962), .B(n30961), .Z(n30966) );
  NANDN U31472 ( .A(n30964), .B(n30963), .Z(n30965) );
  AND U31473 ( .A(n30966), .B(n30965), .Z(n31216) );
  NANDN U31474 ( .A(n30968), .B(n30967), .Z(n30972) );
  NAND U31475 ( .A(n30970), .B(n30969), .Z(n30971) );
  AND U31476 ( .A(n30972), .B(n30971), .Z(n31223) );
  NANDN U31477 ( .A(n30974), .B(n30973), .Z(n30978) );
  NANDN U31478 ( .A(n30976), .B(n30975), .Z(n30977) );
  AND U31479 ( .A(n30978), .B(n30977), .Z(n31221) );
  NANDN U31480 ( .A(n30980), .B(n30979), .Z(n30984) );
  NANDN U31481 ( .A(n30982), .B(n30981), .Z(n30983) );
  AND U31482 ( .A(n30984), .B(n30983), .Z(n31234) );
  NAND U31483 ( .A(n30986), .B(n30985), .Z(n30990) );
  NAND U31484 ( .A(n30988), .B(n30987), .Z(n30989) );
  AND U31485 ( .A(n30990), .B(n30989), .Z(n31446) );
  NANDN U31486 ( .A(n30992), .B(n30991), .Z(n30996) );
  OR U31487 ( .A(n30994), .B(n30993), .Z(n30995) );
  AND U31488 ( .A(n30996), .B(n30995), .Z(n31369) );
  NANDN U31489 ( .A(n30998), .B(n30997), .Z(n31002) );
  NANDN U31490 ( .A(n31000), .B(n30999), .Z(n31001) );
  AND U31491 ( .A(n31002), .B(n31001), .Z(n31367) );
  NANDN U31492 ( .A(n31004), .B(n31003), .Z(n31008) );
  NANDN U31493 ( .A(n31006), .B(n31005), .Z(n31007) );
  AND U31494 ( .A(n31008), .B(n31007), .Z(n31282) );
  NANDN U31495 ( .A(n31010), .B(n31009), .Z(n31014) );
  OR U31496 ( .A(n31012), .B(n31011), .Z(n31013) );
  NAND U31497 ( .A(n31014), .B(n31013), .Z(n31281) );
  XNOR U31498 ( .A(n31282), .B(n31281), .Z(n31283) );
  NANDN U31499 ( .A(n31016), .B(n31015), .Z(n31020) );
  OR U31500 ( .A(n31018), .B(n31017), .Z(n31019) );
  AND U31501 ( .A(n31020), .B(n31019), .Z(n31278) );
  NANDN U31502 ( .A(n31022), .B(n31021), .Z(n31026) );
  ANDN U31503 ( .B(n31024), .A(n31023), .Z(n31025) );
  ANDN U31504 ( .B(n31026), .A(n31025), .Z(n31276) );
  NANDN U31505 ( .A(n37974), .B(n31027), .Z(n31029) );
  XOR U31506 ( .A(b[57]), .B(a[82]), .Z(n31414) );
  NANDN U31507 ( .A(n38031), .B(n31414), .Z(n31028) );
  AND U31508 ( .A(n31029), .B(n31028), .Z(n31318) );
  NANDN U31509 ( .A(n38090), .B(n31030), .Z(n31032) );
  XOR U31510 ( .A(b[59]), .B(a[80]), .Z(n31330) );
  NANDN U31511 ( .A(n38130), .B(n31330), .Z(n31031) );
  AND U31512 ( .A(n31032), .B(n31031), .Z(n31316) );
  NANDN U31513 ( .A(n36210), .B(n31033), .Z(n31035) );
  XOR U31514 ( .A(b[39]), .B(a[100]), .Z(n31251) );
  NANDN U31515 ( .A(n36347), .B(n31251), .Z(n31034) );
  NAND U31516 ( .A(n31035), .B(n31034), .Z(n31315) );
  XNOR U31517 ( .A(n31316), .B(n31315), .Z(n31317) );
  XNOR U31518 ( .A(n31318), .B(n31317), .Z(n31275) );
  XNOR U31519 ( .A(n31276), .B(n31275), .Z(n31277) );
  XOR U31520 ( .A(n31278), .B(n31277), .Z(n31284) );
  XOR U31521 ( .A(n31283), .B(n31284), .Z(n31368) );
  XOR U31522 ( .A(n31367), .B(n31368), .Z(n31370) );
  XOR U31523 ( .A(n31369), .B(n31370), .Z(n31445) );
  NANDN U31524 ( .A(n31037), .B(n31036), .Z(n31041) );
  NANDN U31525 ( .A(n31039), .B(n31038), .Z(n31040) );
  AND U31526 ( .A(n31041), .B(n31040), .Z(n31444) );
  XOR U31527 ( .A(n31445), .B(n31444), .Z(n31447) );
  XNOR U31528 ( .A(n31446), .B(n31447), .Z(n31233) );
  XNOR U31529 ( .A(n31234), .B(n31233), .Z(n31236) );
  NANDN U31530 ( .A(n31043), .B(n31042), .Z(n31047) );
  NANDN U31531 ( .A(n31045), .B(n31044), .Z(n31046) );
  AND U31532 ( .A(n31047), .B(n31046), .Z(n31453) );
  NANDN U31533 ( .A(n31049), .B(n31048), .Z(n31053) );
  NANDN U31534 ( .A(n31051), .B(n31050), .Z(n31052) );
  AND U31535 ( .A(n31053), .B(n31052), .Z(n31451) );
  NANDN U31536 ( .A(n31055), .B(n31054), .Z(n31057) );
  XOR U31537 ( .A(a[126]), .B(b[13]), .Z(n31294) );
  NANDN U31538 ( .A(n31293), .B(n31294), .Z(n31056) );
  AND U31539 ( .A(n31057), .B(n31056), .Z(n31399) );
  NAND U31540 ( .A(b[63]), .B(a[74]), .Z(n31396) );
  ANDN U31541 ( .B(n31059), .A(n31058), .Z(n31062) );
  NAND U31542 ( .A(b[11]), .B(n31060), .Z(n31061) );
  NANDN U31543 ( .A(n31062), .B(n31061), .Z(n31397) );
  XOR U31544 ( .A(n31396), .B(n31397), .Z(n31398) );
  XOR U31545 ( .A(n31399), .B(n31398), .Z(n31345) );
  NANDN U31546 ( .A(n38247), .B(n31063), .Z(n31065) );
  XOR U31547 ( .A(b[61]), .B(a[78]), .Z(n31303) );
  NANDN U31548 ( .A(n38248), .B(n31303), .Z(n31064) );
  AND U31549 ( .A(n31065), .B(n31064), .Z(n31265) );
  NANDN U31550 ( .A(n38278), .B(n31066), .Z(n31068) );
  XOR U31551 ( .A(b[63]), .B(a[76]), .Z(n31248) );
  NANDN U31552 ( .A(n38279), .B(n31248), .Z(n31067) );
  AND U31553 ( .A(n31068), .B(n31067), .Z(n31264) );
  NANDN U31554 ( .A(n36480), .B(n31069), .Z(n31071) );
  XOR U31555 ( .A(b[41]), .B(a[98]), .Z(n31245) );
  NANDN U31556 ( .A(n36594), .B(n31245), .Z(n31070) );
  NAND U31557 ( .A(n31071), .B(n31070), .Z(n31263) );
  XOR U31558 ( .A(n31264), .B(n31263), .Z(n31266) );
  XNOR U31559 ( .A(n31265), .B(n31266), .Z(n31346) );
  XOR U31560 ( .A(n31345), .B(n31346), .Z(n31347) );
  NANDN U31561 ( .A(n31073), .B(n31072), .Z(n31077) );
  OR U31562 ( .A(n31075), .B(n31074), .Z(n31076) );
  NAND U31563 ( .A(n31077), .B(n31076), .Z(n31348) );
  XNOR U31564 ( .A(n31347), .B(n31348), .Z(n31287) );
  NANDN U31565 ( .A(n31079), .B(n31078), .Z(n31083) );
  OR U31566 ( .A(n31081), .B(n31080), .Z(n31082) );
  NAND U31567 ( .A(n31083), .B(n31082), .Z(n31288) );
  XNOR U31568 ( .A(n31287), .B(n31288), .Z(n31289) );
  NANDN U31569 ( .A(n37857), .B(n31084), .Z(n31086) );
  XOR U31570 ( .A(b[55]), .B(a[84]), .Z(n31390) );
  NANDN U31571 ( .A(n37911), .B(n31390), .Z(n31085) );
  AND U31572 ( .A(n31086), .B(n31085), .Z(n31271) );
  NANDN U31573 ( .A(n31536), .B(n31087), .Z(n31089) );
  XOR U31574 ( .A(a[124]), .B(b[15]), .Z(n31300) );
  NANDN U31575 ( .A(n31925), .B(n31300), .Z(n31088) );
  AND U31576 ( .A(n31089), .B(n31088), .Z(n31270) );
  NANDN U31577 ( .A(n35936), .B(n31090), .Z(n31092) );
  XOR U31578 ( .A(b[37]), .B(a[102]), .Z(n31254) );
  NANDN U31579 ( .A(n36047), .B(n31254), .Z(n31091) );
  NAND U31580 ( .A(n31092), .B(n31091), .Z(n31269) );
  XOR U31581 ( .A(n31270), .B(n31269), .Z(n31272) );
  XOR U31582 ( .A(n31271), .B(n31272), .Z(n31350) );
  NANDN U31583 ( .A(n37526), .B(n31093), .Z(n31095) );
  XOR U31584 ( .A(b[51]), .B(a[88]), .Z(n31420) );
  NANDN U31585 ( .A(n37605), .B(n31420), .Z(n31094) );
  AND U31586 ( .A(n31095), .B(n31094), .Z(n31311) );
  NANDN U31587 ( .A(n37705), .B(n31096), .Z(n31098) );
  XOR U31588 ( .A(b[53]), .B(a[86]), .Z(n31387) );
  NANDN U31589 ( .A(n37778), .B(n31387), .Z(n31097) );
  AND U31590 ( .A(n31098), .B(n31097), .Z(n31310) );
  NANDN U31591 ( .A(n36742), .B(n31099), .Z(n31101) );
  XOR U31592 ( .A(b[43]), .B(a[96]), .Z(n31306) );
  NANDN U31593 ( .A(n36891), .B(n31306), .Z(n31100) );
  NAND U31594 ( .A(n31101), .B(n31100), .Z(n31309) );
  XOR U31595 ( .A(n31310), .B(n31309), .Z(n31312) );
  XNOR U31596 ( .A(n31311), .B(n31312), .Z(n31349) );
  XNOR U31597 ( .A(n31350), .B(n31349), .Z(n31351) );
  NANDN U31598 ( .A(n31103), .B(n31102), .Z(n31107) );
  OR U31599 ( .A(n31105), .B(n31104), .Z(n31106) );
  NAND U31600 ( .A(n31107), .B(n31106), .Z(n31352) );
  XOR U31601 ( .A(n31351), .B(n31352), .Z(n31290) );
  XNOR U31602 ( .A(n31289), .B(n31290), .Z(n31441) );
  NANDN U31603 ( .A(n31109), .B(n31108), .Z(n31113) );
  NANDN U31604 ( .A(n31111), .B(n31110), .Z(n31112) );
  AND U31605 ( .A(n31113), .B(n31112), .Z(n31439) );
  NAND U31606 ( .A(n31115), .B(n31114), .Z(n31119) );
  NAND U31607 ( .A(n31117), .B(n31116), .Z(n31118) );
  NAND U31608 ( .A(n31119), .B(n31118), .Z(n31438) );
  XNOR U31609 ( .A(n31439), .B(n31438), .Z(n31440) );
  XOR U31610 ( .A(n31441), .B(n31440), .Z(n31378) );
  NANDN U31611 ( .A(n31121), .B(n31120), .Z(n31125) );
  OR U31612 ( .A(n31123), .B(n31122), .Z(n31124) );
  AND U31613 ( .A(n31125), .B(n31124), .Z(n31377) );
  XNOR U31614 ( .A(n31378), .B(n31377), .Z(n31380) );
  NANDN U31615 ( .A(n31127), .B(n31126), .Z(n31131) );
  NANDN U31616 ( .A(n31129), .B(n31128), .Z(n31130) );
  AND U31617 ( .A(n31131), .B(n31130), .Z(n31374) );
  NANDN U31618 ( .A(n31133), .B(n31132), .Z(n31137) );
  NANDN U31619 ( .A(n31135), .B(n31134), .Z(n31136) );
  AND U31620 ( .A(n31137), .B(n31136), .Z(n31373) );
  XNOR U31621 ( .A(n31374), .B(n31373), .Z(n31376) );
  NANDN U31622 ( .A(n34634), .B(n31138), .Z(n31140) );
  XOR U31623 ( .A(a[110]), .B(b[29]), .Z(n31423) );
  NANDN U31624 ( .A(n34722), .B(n31423), .Z(n31139) );
  AND U31625 ( .A(n31140), .B(n31139), .Z(n31259) );
  NANDN U31626 ( .A(n34909), .B(n31141), .Z(n31143) );
  XOR U31627 ( .A(a[108]), .B(b[31]), .Z(n31239) );
  NANDN U31628 ( .A(n35145), .B(n31239), .Z(n31142) );
  AND U31629 ( .A(n31143), .B(n31142), .Z(n31258) );
  NANDN U31630 ( .A(n32483), .B(n31144), .Z(n31146) );
  XOR U31631 ( .A(a[120]), .B(b[19]), .Z(n31321) );
  NANDN U31632 ( .A(n32823), .B(n31321), .Z(n31145) );
  NAND U31633 ( .A(n31146), .B(n31145), .Z(n31257) );
  XOR U31634 ( .A(n31258), .B(n31257), .Z(n31260) );
  XOR U31635 ( .A(n31259), .B(n31260), .Z(n31434) );
  NANDN U31636 ( .A(n31147), .B(n34297), .Z(n31149) );
  XOR U31637 ( .A(a[114]), .B(b[25]), .Z(n31408) );
  NANDN U31638 ( .A(n33994), .B(n31408), .Z(n31148) );
  AND U31639 ( .A(n31149), .B(n31148), .Z(n31341) );
  NANDN U31640 ( .A(n33866), .B(n31150), .Z(n31152) );
  XOR U31641 ( .A(a[116]), .B(b[23]), .Z(n31411) );
  NANDN U31642 ( .A(n33644), .B(n31411), .Z(n31151) );
  AND U31643 ( .A(n31152), .B(n31151), .Z(n31340) );
  NANDN U31644 ( .A(n32996), .B(n31153), .Z(n31155) );
  XOR U31645 ( .A(a[118]), .B(b[21]), .Z(n31333) );
  NANDN U31646 ( .A(n33271), .B(n31333), .Z(n31154) );
  NAND U31647 ( .A(n31155), .B(n31154), .Z(n31339) );
  XOR U31648 ( .A(n31340), .B(n31339), .Z(n31342) );
  XOR U31649 ( .A(n31341), .B(n31342), .Z(n31433) );
  NAND U31650 ( .A(n34647), .B(n31156), .Z(n31158) );
  XNOR U31651 ( .A(a[112]), .B(b[27]), .Z(n31393) );
  NANDN U31652 ( .A(n31393), .B(n34648), .Z(n31157) );
  AND U31653 ( .A(n31158), .B(n31157), .Z(n31432) );
  XOR U31654 ( .A(n31433), .B(n31432), .Z(n31435) );
  XOR U31655 ( .A(n31434), .B(n31435), .Z(n31358) );
  NANDN U31656 ( .A(n31160), .B(n31159), .Z(n31164) );
  OR U31657 ( .A(n31162), .B(n31161), .Z(n31163) );
  AND U31658 ( .A(n31164), .B(n31163), .Z(n31356) );
  NANDN U31659 ( .A(n31166), .B(n31165), .Z(n31170) );
  NAND U31660 ( .A(n31168), .B(n31167), .Z(n31169) );
  NAND U31661 ( .A(n31170), .B(n31169), .Z(n31355) );
  XNOR U31662 ( .A(n31356), .B(n31355), .Z(n31357) );
  XNOR U31663 ( .A(n31358), .B(n31357), .Z(n31384) );
  NANDN U31664 ( .A(n31172), .B(n31171), .Z(n31176) );
  NANDN U31665 ( .A(n31174), .B(n31173), .Z(n31175) );
  AND U31666 ( .A(n31176), .B(n31175), .Z(n31382) );
  NANDN U31667 ( .A(n36991), .B(n31177), .Z(n31179) );
  XOR U31668 ( .A(b[45]), .B(a[94]), .Z(n31327) );
  NANDN U31669 ( .A(n37083), .B(n31327), .Z(n31178) );
  AND U31670 ( .A(n31179), .B(n31178), .Z(n31428) );
  NANDN U31671 ( .A(n211), .B(n31180), .Z(n31182) );
  XOR U31672 ( .A(b[47]), .B(a[92]), .Z(n31417) );
  NANDN U31673 ( .A(n37172), .B(n31417), .Z(n31181) );
  AND U31674 ( .A(n31182), .B(n31181), .Z(n31427) );
  NANDN U31675 ( .A(n212), .B(n31183), .Z(n31185) );
  XOR U31676 ( .A(b[49]), .B(a[90]), .Z(n31336) );
  NANDN U31677 ( .A(n37432), .B(n31336), .Z(n31184) );
  NAND U31678 ( .A(n31185), .B(n31184), .Z(n31426) );
  XOR U31679 ( .A(n31427), .B(n31426), .Z(n31429) );
  XOR U31680 ( .A(n31428), .B(n31429), .Z(n31362) );
  NANDN U31681 ( .A(n35260), .B(n31186), .Z(n31188) );
  XOR U31682 ( .A(a[106]), .B(b[33]), .Z(n31242) );
  NANDN U31683 ( .A(n35456), .B(n31242), .Z(n31187) );
  AND U31684 ( .A(n31188), .B(n31187), .Z(n31404) );
  NANDN U31685 ( .A(n35611), .B(n31189), .Z(n31191) );
  XOR U31686 ( .A(a[104]), .B(b[35]), .Z(n31297) );
  NANDN U31687 ( .A(n35801), .B(n31297), .Z(n31190) );
  AND U31688 ( .A(n31191), .B(n31190), .Z(n31403) );
  NANDN U31689 ( .A(n32013), .B(n31192), .Z(n31194) );
  XOR U31690 ( .A(a[122]), .B(b[17]), .Z(n31324) );
  NANDN U31691 ( .A(n32292), .B(n31324), .Z(n31193) );
  NAND U31692 ( .A(n31194), .B(n31193), .Z(n31402) );
  XOR U31693 ( .A(n31403), .B(n31402), .Z(n31405) );
  XNOR U31694 ( .A(n31404), .B(n31405), .Z(n31361) );
  XNOR U31695 ( .A(n31362), .B(n31361), .Z(n31364) );
  NANDN U31696 ( .A(n31196), .B(n31195), .Z(n31200) );
  OR U31697 ( .A(n31198), .B(n31197), .Z(n31199) );
  AND U31698 ( .A(n31200), .B(n31199), .Z(n31363) );
  XNOR U31699 ( .A(n31364), .B(n31363), .Z(n31381) );
  XOR U31700 ( .A(n31382), .B(n31381), .Z(n31383) );
  XOR U31701 ( .A(n31384), .B(n31383), .Z(n31375) );
  XOR U31702 ( .A(n31376), .B(n31375), .Z(n31379) );
  XOR U31703 ( .A(n31380), .B(n31379), .Z(n31450) );
  XNOR U31704 ( .A(n31451), .B(n31450), .Z(n31452) );
  XNOR U31705 ( .A(n31453), .B(n31452), .Z(n31235) );
  XOR U31706 ( .A(n31236), .B(n31235), .Z(n31230) );
  NANDN U31707 ( .A(n31202), .B(n31201), .Z(n31206) );
  NANDN U31708 ( .A(n31204), .B(n31203), .Z(n31205) );
  AND U31709 ( .A(n31206), .B(n31205), .Z(n31227) );
  NANDN U31710 ( .A(n31208), .B(n31207), .Z(n31212) );
  NANDN U31711 ( .A(n31210), .B(n31209), .Z(n31211) );
  NAND U31712 ( .A(n31212), .B(n31211), .Z(n31228) );
  XNOR U31713 ( .A(n31227), .B(n31228), .Z(n31229) );
  XOR U31714 ( .A(n31230), .B(n31229), .Z(n31222) );
  XOR U31715 ( .A(n31221), .B(n31222), .Z(n31224) );
  XNOR U31716 ( .A(n31223), .B(n31224), .Z(n31215) );
  XOR U31717 ( .A(n31216), .B(n31215), .Z(n31218) );
  XNOR U31718 ( .A(n31217), .B(n31218), .Z(n31213) );
  XOR U31719 ( .A(n31214), .B(n31213), .Z(c[202]) );
  AND U31720 ( .A(n31214), .B(n31213), .Z(n31457) );
  NANDN U31721 ( .A(n31216), .B(n31215), .Z(n31220) );
  OR U31722 ( .A(n31218), .B(n31217), .Z(n31219) );
  AND U31723 ( .A(n31220), .B(n31219), .Z(n31460) );
  NANDN U31724 ( .A(n31222), .B(n31221), .Z(n31226) );
  NANDN U31725 ( .A(n31224), .B(n31223), .Z(n31225) );
  AND U31726 ( .A(n31226), .B(n31225), .Z(n31459) );
  NANDN U31727 ( .A(n31228), .B(n31227), .Z(n31232) );
  NANDN U31728 ( .A(n31230), .B(n31229), .Z(n31231) );
  AND U31729 ( .A(n31232), .B(n31231), .Z(n31467) );
  NANDN U31730 ( .A(n31234), .B(n31233), .Z(n31238) );
  NAND U31731 ( .A(n31236), .B(n31235), .Z(n31237) );
  AND U31732 ( .A(n31238), .B(n31237), .Z(n31464) );
  NANDN U31733 ( .A(n34909), .B(n31239), .Z(n31241) );
  XOR U31734 ( .A(a[109]), .B(b[31]), .Z(n31500) );
  NANDN U31735 ( .A(n35145), .B(n31500), .Z(n31240) );
  AND U31736 ( .A(n31241), .B(n31240), .Z(n31490) );
  NANDN U31737 ( .A(n35260), .B(n31242), .Z(n31244) );
  XOR U31738 ( .A(a[107]), .B(b[33]), .Z(n31581) );
  NANDN U31739 ( .A(n35456), .B(n31581), .Z(n31243) );
  AND U31740 ( .A(n31244), .B(n31243), .Z(n31489) );
  NANDN U31741 ( .A(n36480), .B(n31245), .Z(n31247) );
  XOR U31742 ( .A(b[41]), .B(a[99]), .Z(n31539) );
  NANDN U31743 ( .A(n36594), .B(n31539), .Z(n31246) );
  NAND U31744 ( .A(n31247), .B(n31246), .Z(n31488) );
  XOR U31745 ( .A(n31489), .B(n31488), .Z(n31491) );
  XOR U31746 ( .A(n31490), .B(n31491), .Z(n31654) );
  NANDN U31747 ( .A(n38278), .B(n31248), .Z(n31250) );
  XOR U31748 ( .A(b[63]), .B(a[77]), .Z(n31503) );
  NANDN U31749 ( .A(n38279), .B(n31503), .Z(n31249) );
  AND U31750 ( .A(n31250), .B(n31249), .Z(n31606) );
  NANDN U31751 ( .A(n36210), .B(n31251), .Z(n31253) );
  XOR U31752 ( .A(b[39]), .B(a[101]), .Z(n31584) );
  NANDN U31753 ( .A(n36347), .B(n31584), .Z(n31252) );
  NAND U31754 ( .A(n31253), .B(n31252), .Z(n31605) );
  XNOR U31755 ( .A(n31606), .B(n31605), .Z(n31608) );
  NANDN U31756 ( .A(n35936), .B(n31254), .Z(n31256) );
  XOR U31757 ( .A(b[37]), .B(a[103]), .Z(n31554) );
  NANDN U31758 ( .A(n36047), .B(n31554), .Z(n31255) );
  AND U31759 ( .A(n31256), .B(n31255), .Z(n31588) );
  AND U31760 ( .A(b[63]), .B(a[75]), .Z(n31587) );
  XOR U31761 ( .A(n31588), .B(n31587), .Z(n31590) );
  XOR U31762 ( .A(n31396), .B(n31590), .Z(n31607) );
  XNOR U31763 ( .A(n31608), .B(n31607), .Z(n31653) );
  XNOR U31764 ( .A(n31654), .B(n31653), .Z(n31655) );
  NANDN U31765 ( .A(n31258), .B(n31257), .Z(n31262) );
  OR U31766 ( .A(n31260), .B(n31259), .Z(n31261) );
  NAND U31767 ( .A(n31262), .B(n31261), .Z(n31656) );
  XNOR U31768 ( .A(n31655), .B(n31656), .Z(n31613) );
  NANDN U31769 ( .A(n31264), .B(n31263), .Z(n31268) );
  OR U31770 ( .A(n31266), .B(n31265), .Z(n31267) );
  AND U31771 ( .A(n31268), .B(n31267), .Z(n31611) );
  NANDN U31772 ( .A(n31270), .B(n31269), .Z(n31274) );
  OR U31773 ( .A(n31272), .B(n31271), .Z(n31273) );
  NAND U31774 ( .A(n31274), .B(n31273), .Z(n31612) );
  XOR U31775 ( .A(n31611), .B(n31612), .Z(n31614) );
  XNOR U31776 ( .A(n31613), .B(n31614), .Z(n31629) );
  NANDN U31777 ( .A(n31276), .B(n31275), .Z(n31280) );
  NANDN U31778 ( .A(n31278), .B(n31277), .Z(n31279) );
  NAND U31779 ( .A(n31280), .B(n31279), .Z(n31630) );
  XNOR U31780 ( .A(n31629), .B(n31630), .Z(n31632) );
  NANDN U31781 ( .A(n31282), .B(n31281), .Z(n31286) );
  NANDN U31782 ( .A(n31284), .B(n31283), .Z(n31285) );
  AND U31783 ( .A(n31286), .B(n31285), .Z(n31631) );
  XOR U31784 ( .A(n31632), .B(n31631), .Z(n31642) );
  NANDN U31785 ( .A(n31288), .B(n31287), .Z(n31292) );
  NANDN U31786 ( .A(n31290), .B(n31289), .Z(n31291) );
  AND U31787 ( .A(n31292), .B(n31291), .Z(n31641) );
  XNOR U31788 ( .A(n31642), .B(n31641), .Z(n31644) );
  XNOR U31789 ( .A(a[127]), .B(b[13]), .Z(n31506) );
  OR U31790 ( .A(n31506), .B(n31293), .Z(n31296) );
  NAND U31791 ( .A(n31507), .B(n31294), .Z(n31295) );
  AND U31792 ( .A(n31296), .B(n31295), .Z(n31513) );
  NANDN U31793 ( .A(n35611), .B(n31297), .Z(n31299) );
  XOR U31794 ( .A(a[105]), .B(b[35]), .Z(n31578) );
  NANDN U31795 ( .A(n35801), .B(n31578), .Z(n31298) );
  NAND U31796 ( .A(n31299), .B(n31298), .Z(n31511) );
  XOR U31797 ( .A(n31512), .B(n31511), .Z(n31514) );
  XOR U31798 ( .A(n31513), .B(n31514), .Z(n31618) );
  NANDN U31799 ( .A(n31536), .B(n31300), .Z(n31302) );
  XOR U31800 ( .A(a[125]), .B(b[15]), .Z(n31535) );
  NANDN U31801 ( .A(n31925), .B(n31535), .Z(n31301) );
  AND U31802 ( .A(n31302), .B(n31301), .Z(n31519) );
  NANDN U31803 ( .A(n38247), .B(n31303), .Z(n31305) );
  XOR U31804 ( .A(b[61]), .B(a[79]), .Z(n31526) );
  NANDN U31805 ( .A(n38248), .B(n31526), .Z(n31304) );
  AND U31806 ( .A(n31305), .B(n31304), .Z(n31518) );
  NANDN U31807 ( .A(n36742), .B(n31306), .Z(n31308) );
  XOR U31808 ( .A(b[43]), .B(a[97]), .Z(n31494) );
  NANDN U31809 ( .A(n36891), .B(n31494), .Z(n31307) );
  NAND U31810 ( .A(n31308), .B(n31307), .Z(n31517) );
  XOR U31811 ( .A(n31518), .B(n31517), .Z(n31520) );
  XNOR U31812 ( .A(n31519), .B(n31520), .Z(n31617) );
  XNOR U31813 ( .A(n31618), .B(n31617), .Z(n31619) );
  NANDN U31814 ( .A(n31310), .B(n31309), .Z(n31314) );
  OR U31815 ( .A(n31312), .B(n31311), .Z(n31313) );
  NAND U31816 ( .A(n31314), .B(n31313), .Z(n31620) );
  XNOR U31817 ( .A(n31619), .B(n31620), .Z(n31482) );
  NANDN U31818 ( .A(n31316), .B(n31315), .Z(n31320) );
  NANDN U31819 ( .A(n31318), .B(n31317), .Z(n31319) );
  NAND U31820 ( .A(n31320), .B(n31319), .Z(n31483) );
  XNOR U31821 ( .A(n31482), .B(n31483), .Z(n31484) );
  NANDN U31822 ( .A(n32483), .B(n31321), .Z(n31323) );
  XOR U31823 ( .A(a[121]), .B(b[19]), .Z(n31523) );
  NANDN U31824 ( .A(n32823), .B(n31523), .Z(n31322) );
  AND U31825 ( .A(n31323), .B(n31322), .Z(n31601) );
  NANDN U31826 ( .A(n32013), .B(n31324), .Z(n31326) );
  XOR U31827 ( .A(a[123]), .B(b[17]), .Z(n31532) );
  NANDN U31828 ( .A(n32292), .B(n31532), .Z(n31325) );
  AND U31829 ( .A(n31326), .B(n31325), .Z(n31600) );
  NANDN U31830 ( .A(n36991), .B(n31327), .Z(n31329) );
  XOR U31831 ( .A(b[45]), .B(a[95]), .Z(n31529) );
  NANDN U31832 ( .A(n37083), .B(n31529), .Z(n31328) );
  NAND U31833 ( .A(n31329), .B(n31328), .Z(n31599) );
  XOR U31834 ( .A(n31600), .B(n31599), .Z(n31602) );
  XOR U31835 ( .A(n31601), .B(n31602), .Z(n31660) );
  NANDN U31836 ( .A(n38090), .B(n31330), .Z(n31332) );
  XOR U31837 ( .A(b[59]), .B(a[81]), .Z(n31674) );
  NANDN U31838 ( .A(n38130), .B(n31674), .Z(n31331) );
  AND U31839 ( .A(n31332), .B(n31331), .Z(n31568) );
  NANDN U31840 ( .A(n32996), .B(n31333), .Z(n31335) );
  XOR U31841 ( .A(a[119]), .B(b[21]), .Z(n31560) );
  NANDN U31842 ( .A(n33271), .B(n31560), .Z(n31334) );
  AND U31843 ( .A(n31335), .B(n31334), .Z(n31567) );
  NANDN U31844 ( .A(n212), .B(n31336), .Z(n31338) );
  XOR U31845 ( .A(b[49]), .B(a[91]), .Z(n31497) );
  NANDN U31846 ( .A(n37432), .B(n31497), .Z(n31337) );
  NAND U31847 ( .A(n31338), .B(n31337), .Z(n31566) );
  XOR U31848 ( .A(n31567), .B(n31566), .Z(n31569) );
  XNOR U31849 ( .A(n31568), .B(n31569), .Z(n31659) );
  XNOR U31850 ( .A(n31660), .B(n31659), .Z(n31661) );
  NANDN U31851 ( .A(n31340), .B(n31339), .Z(n31344) );
  OR U31852 ( .A(n31342), .B(n31341), .Z(n31343) );
  NAND U31853 ( .A(n31344), .B(n31343), .Z(n31662) );
  XOR U31854 ( .A(n31661), .B(n31662), .Z(n31485) );
  XNOR U31855 ( .A(n31484), .B(n31485), .Z(n31650) );
  NANDN U31856 ( .A(n31350), .B(n31349), .Z(n31354) );
  NANDN U31857 ( .A(n31352), .B(n31351), .Z(n31353) );
  NAND U31858 ( .A(n31354), .B(n31353), .Z(n31647) );
  XNOR U31859 ( .A(n31648), .B(n31647), .Z(n31649) );
  XOR U31860 ( .A(n31650), .B(n31649), .Z(n31638) );
  NANDN U31861 ( .A(n31356), .B(n31355), .Z(n31360) );
  NANDN U31862 ( .A(n31358), .B(n31357), .Z(n31359) );
  AND U31863 ( .A(n31360), .B(n31359), .Z(n31636) );
  NANDN U31864 ( .A(n31362), .B(n31361), .Z(n31366) );
  NAND U31865 ( .A(n31364), .B(n31363), .Z(n31365) );
  AND U31866 ( .A(n31366), .B(n31365), .Z(n31635) );
  XNOR U31867 ( .A(n31636), .B(n31635), .Z(n31637) );
  XNOR U31868 ( .A(n31638), .B(n31637), .Z(n31643) );
  XOR U31869 ( .A(n31644), .B(n31643), .Z(n31696) );
  NANDN U31870 ( .A(n31368), .B(n31367), .Z(n31372) );
  OR U31871 ( .A(n31370), .B(n31369), .Z(n31371) );
  AND U31872 ( .A(n31372), .B(n31371), .Z(n31695) );
  XNOR U31873 ( .A(n31696), .B(n31695), .Z(n31698) );
  XOR U31874 ( .A(n31698), .B(n31697), .Z(n31478) );
  NAND U31875 ( .A(n31382), .B(n31381), .Z(n31386) );
  NAND U31876 ( .A(n31384), .B(n31383), .Z(n31385) );
  AND U31877 ( .A(n31386), .B(n31385), .Z(n31704) );
  NANDN U31878 ( .A(n37705), .B(n31387), .Z(n31389) );
  XOR U31879 ( .A(b[53]), .B(a[87]), .Z(n31665) );
  NANDN U31880 ( .A(n37778), .B(n31665), .Z(n31388) );
  AND U31881 ( .A(n31389), .B(n31388), .Z(n31685) );
  NANDN U31882 ( .A(n37857), .B(n31390), .Z(n31392) );
  XOR U31883 ( .A(b[55]), .B(a[85]), .Z(n31668) );
  NANDN U31884 ( .A(n37911), .B(n31668), .Z(n31391) );
  AND U31885 ( .A(n31392), .B(n31391), .Z(n31684) );
  NANDN U31886 ( .A(n31393), .B(n34647), .Z(n31395) );
  XOR U31887 ( .A(a[113]), .B(b[27]), .Z(n31551) );
  NANDN U31888 ( .A(n34458), .B(n31551), .Z(n31394) );
  NAND U31889 ( .A(n31395), .B(n31394), .Z(n31683) );
  XOR U31890 ( .A(n31684), .B(n31683), .Z(n31686) );
  XOR U31891 ( .A(n31685), .B(n31686), .Z(n31624) );
  IV U31892 ( .A(n31396), .Z(n31589) );
  NANDN U31893 ( .A(n31589), .B(n31397), .Z(n31401) );
  NANDN U31894 ( .A(n31399), .B(n31398), .Z(n31400) );
  AND U31895 ( .A(n31401), .B(n31400), .Z(n31623) );
  XNOR U31896 ( .A(n31624), .B(n31623), .Z(n31626) );
  NANDN U31897 ( .A(n31403), .B(n31402), .Z(n31407) );
  OR U31898 ( .A(n31405), .B(n31404), .Z(n31406) );
  AND U31899 ( .A(n31407), .B(n31406), .Z(n31625) );
  XOR U31900 ( .A(n31626), .B(n31625), .Z(n31691) );
  NANDN U31901 ( .A(n33875), .B(n31408), .Z(n31410) );
  XOR U31902 ( .A(a[115]), .B(b[25]), .Z(n31677) );
  NANDN U31903 ( .A(n33994), .B(n31677), .Z(n31409) );
  AND U31904 ( .A(n31410), .B(n31409), .Z(n31544) );
  NANDN U31905 ( .A(n33866), .B(n31411), .Z(n31413) );
  XOR U31906 ( .A(a[117]), .B(b[23]), .Z(n31557) );
  NANDN U31907 ( .A(n33644), .B(n31557), .Z(n31412) );
  AND U31908 ( .A(n31413), .B(n31412), .Z(n31543) );
  NANDN U31909 ( .A(n37974), .B(n31414), .Z(n31416) );
  XOR U31910 ( .A(b[57]), .B(a[83]), .Z(n31548) );
  NANDN U31911 ( .A(n38031), .B(n31548), .Z(n31415) );
  NAND U31912 ( .A(n31416), .B(n31415), .Z(n31542) );
  XOR U31913 ( .A(n31543), .B(n31542), .Z(n31545) );
  XOR U31914 ( .A(n31544), .B(n31545), .Z(n31573) );
  NANDN U31915 ( .A(n211), .B(n31417), .Z(n31419) );
  XOR U31916 ( .A(b[47]), .B(a[93]), .Z(n31563) );
  NANDN U31917 ( .A(n37172), .B(n31563), .Z(n31418) );
  AND U31918 ( .A(n31419), .B(n31418), .Z(n31595) );
  NANDN U31919 ( .A(n37526), .B(n31420), .Z(n31422) );
  XOR U31920 ( .A(b[51]), .B(a[89]), .Z(n31680) );
  NANDN U31921 ( .A(n37605), .B(n31680), .Z(n31421) );
  AND U31922 ( .A(n31422), .B(n31421), .Z(n31594) );
  NANDN U31923 ( .A(n34634), .B(n31423), .Z(n31425) );
  XOR U31924 ( .A(a[111]), .B(b[29]), .Z(n31671) );
  NANDN U31925 ( .A(n34722), .B(n31671), .Z(n31424) );
  NAND U31926 ( .A(n31425), .B(n31424), .Z(n31593) );
  XOR U31927 ( .A(n31594), .B(n31593), .Z(n31596) );
  XNOR U31928 ( .A(n31595), .B(n31596), .Z(n31572) );
  XNOR U31929 ( .A(n31573), .B(n31572), .Z(n31575) );
  NANDN U31930 ( .A(n31427), .B(n31426), .Z(n31431) );
  OR U31931 ( .A(n31429), .B(n31428), .Z(n31430) );
  AND U31932 ( .A(n31431), .B(n31430), .Z(n31574) );
  XOR U31933 ( .A(n31575), .B(n31574), .Z(n31690) );
  NANDN U31934 ( .A(n31433), .B(n31432), .Z(n31437) );
  OR U31935 ( .A(n31435), .B(n31434), .Z(n31436) );
  AND U31936 ( .A(n31437), .B(n31436), .Z(n31689) );
  XOR U31937 ( .A(n31690), .B(n31689), .Z(n31692) );
  XOR U31938 ( .A(n31691), .B(n31692), .Z(n31702) );
  NANDN U31939 ( .A(n31439), .B(n31438), .Z(n31443) );
  NAND U31940 ( .A(n31441), .B(n31440), .Z(n31442) );
  NAND U31941 ( .A(n31443), .B(n31442), .Z(n31701) );
  XNOR U31942 ( .A(n31702), .B(n31701), .Z(n31703) );
  XNOR U31943 ( .A(n31704), .B(n31703), .Z(n31476) );
  XOR U31944 ( .A(n31477), .B(n31476), .Z(n31479) );
  XOR U31945 ( .A(n31478), .B(n31479), .Z(n31473) );
  NANDN U31946 ( .A(n31445), .B(n31444), .Z(n31449) );
  OR U31947 ( .A(n31447), .B(n31446), .Z(n31448) );
  AND U31948 ( .A(n31449), .B(n31448), .Z(n31471) );
  NANDN U31949 ( .A(n31451), .B(n31450), .Z(n31455) );
  NANDN U31950 ( .A(n31453), .B(n31452), .Z(n31454) );
  AND U31951 ( .A(n31455), .B(n31454), .Z(n31470) );
  XNOR U31952 ( .A(n31471), .B(n31470), .Z(n31472) );
  XOR U31953 ( .A(n31473), .B(n31472), .Z(n31465) );
  XNOR U31954 ( .A(n31464), .B(n31465), .Z(n31466) );
  XNOR U31955 ( .A(n31467), .B(n31466), .Z(n31458) );
  XOR U31956 ( .A(n31459), .B(n31458), .Z(n31461) );
  XNOR U31957 ( .A(n31460), .B(n31461), .Z(n31456) );
  XOR U31958 ( .A(n31457), .B(n31456), .Z(c[203]) );
  AND U31959 ( .A(n31457), .B(n31456), .Z(n31708) );
  NANDN U31960 ( .A(n31459), .B(n31458), .Z(n31463) );
  OR U31961 ( .A(n31461), .B(n31460), .Z(n31462) );
  AND U31962 ( .A(n31463), .B(n31462), .Z(n31711) );
  NANDN U31963 ( .A(n31465), .B(n31464), .Z(n31469) );
  NANDN U31964 ( .A(n31467), .B(n31466), .Z(n31468) );
  AND U31965 ( .A(n31469), .B(n31468), .Z(n31710) );
  NANDN U31966 ( .A(n31471), .B(n31470), .Z(n31475) );
  NANDN U31967 ( .A(n31473), .B(n31472), .Z(n31474) );
  AND U31968 ( .A(n31475), .B(n31474), .Z(n31718) );
  NANDN U31969 ( .A(n31477), .B(n31476), .Z(n31481) );
  OR U31970 ( .A(n31479), .B(n31478), .Z(n31480) );
  AND U31971 ( .A(n31481), .B(n31480), .Z(n31715) );
  NANDN U31972 ( .A(n31483), .B(n31482), .Z(n31487) );
  NANDN U31973 ( .A(n31485), .B(n31484), .Z(n31486) );
  AND U31974 ( .A(n31487), .B(n31486), .Z(n31733) );
  NANDN U31975 ( .A(n31489), .B(n31488), .Z(n31493) );
  OR U31976 ( .A(n31491), .B(n31490), .Z(n31492) );
  AND U31977 ( .A(n31493), .B(n31492), .Z(n31775) );
  NANDN U31978 ( .A(n36742), .B(n31494), .Z(n31496) );
  XOR U31979 ( .A(b[43]), .B(a[98]), .Z(n31932) );
  NANDN U31980 ( .A(n36891), .B(n31932), .Z(n31495) );
  AND U31981 ( .A(n31496), .B(n31495), .Z(n31829) );
  NANDN U31982 ( .A(n212), .B(n31497), .Z(n31499) );
  XOR U31983 ( .A(b[49]), .B(a[92]), .Z(n31790) );
  NANDN U31984 ( .A(n37432), .B(n31790), .Z(n31498) );
  AND U31985 ( .A(n31499), .B(n31498), .Z(n31827) );
  NANDN U31986 ( .A(n34909), .B(n31500), .Z(n31502) );
  XOR U31987 ( .A(a[110]), .B(b[31]), .Z(n31913) );
  NANDN U31988 ( .A(n35145), .B(n31913), .Z(n31501) );
  NAND U31989 ( .A(n31502), .B(n31501), .Z(n31826) );
  XNOR U31990 ( .A(n31827), .B(n31826), .Z(n31828) );
  XOR U31991 ( .A(n31829), .B(n31828), .Z(n31773) );
  NANDN U31992 ( .A(n38278), .B(n31503), .Z(n31505) );
  XOR U31993 ( .A(b[63]), .B(a[78]), .Z(n31929) );
  NANDN U31994 ( .A(n38279), .B(n31929), .Z(n31504) );
  AND U31995 ( .A(n31505), .B(n31504), .Z(n31938) );
  NAND U31996 ( .A(b[63]), .B(a[76]), .Z(n31935) );
  ANDN U31997 ( .B(n31507), .A(n31506), .Z(n31510) );
  NAND U31998 ( .A(b[13]), .B(n31508), .Z(n31509) );
  NANDN U31999 ( .A(n31510), .B(n31509), .Z(n31936) );
  XOR U32000 ( .A(n31935), .B(n31936), .Z(n31937) );
  XOR U32001 ( .A(n31938), .B(n31937), .Z(n31772) );
  XOR U32002 ( .A(n31773), .B(n31772), .Z(n31774) );
  XOR U32003 ( .A(n31775), .B(n31774), .Z(n31858) );
  NANDN U32004 ( .A(n31512), .B(n31511), .Z(n31516) );
  OR U32005 ( .A(n31514), .B(n31513), .Z(n31515) );
  AND U32006 ( .A(n31516), .B(n31515), .Z(n31857) );
  NANDN U32007 ( .A(n31518), .B(n31517), .Z(n31522) );
  OR U32008 ( .A(n31520), .B(n31519), .Z(n31521) );
  NAND U32009 ( .A(n31522), .B(n31521), .Z(n31856) );
  XOR U32010 ( .A(n31857), .B(n31856), .Z(n31859) );
  XOR U32011 ( .A(n31858), .B(n31859), .Z(n31943) );
  NANDN U32012 ( .A(n32483), .B(n31523), .Z(n31525) );
  XOR U32013 ( .A(a[122]), .B(b[19]), .Z(n31808) );
  NANDN U32014 ( .A(n32823), .B(n31808), .Z(n31524) );
  AND U32015 ( .A(n31525), .B(n31524), .Z(n31741) );
  NANDN U32016 ( .A(n38247), .B(n31526), .Z(n31528) );
  XOR U32017 ( .A(b[61]), .B(a[80]), .Z(n31784) );
  NANDN U32018 ( .A(n38248), .B(n31784), .Z(n31527) );
  AND U32019 ( .A(n31528), .B(n31527), .Z(n31740) );
  NANDN U32020 ( .A(n36991), .B(n31529), .Z(n31531) );
  XOR U32021 ( .A(b[45]), .B(a[96]), .Z(n31814) );
  NANDN U32022 ( .A(n37083), .B(n31814), .Z(n31530) );
  NAND U32023 ( .A(n31531), .B(n31530), .Z(n31739) );
  XOR U32024 ( .A(n31740), .B(n31739), .Z(n31742) );
  XOR U32025 ( .A(n31741), .B(n31742), .Z(n31851) );
  NANDN U32026 ( .A(n32013), .B(n31532), .Z(n31534) );
  XOR U32027 ( .A(a[124]), .B(b[17]), .Z(n31811) );
  NANDN U32028 ( .A(n32292), .B(n31811), .Z(n31533) );
  AND U32029 ( .A(n31534), .B(n31533), .Z(n31840) );
  NANDN U32030 ( .A(n31536), .B(n31535), .Z(n31538) );
  XOR U32031 ( .A(a[126]), .B(b[15]), .Z(n31926) );
  NANDN U32032 ( .A(n31925), .B(n31926), .Z(n31537) );
  AND U32033 ( .A(n31538), .B(n31537), .Z(n31839) );
  NANDN U32034 ( .A(n36480), .B(n31539), .Z(n31541) );
  XOR U32035 ( .A(b[41]), .B(a[100]), .Z(n31760) );
  NANDN U32036 ( .A(n36594), .B(n31760), .Z(n31540) );
  NAND U32037 ( .A(n31541), .B(n31540), .Z(n31838) );
  XOR U32038 ( .A(n31839), .B(n31838), .Z(n31841) );
  XNOR U32039 ( .A(n31840), .B(n31841), .Z(n31850) );
  XNOR U32040 ( .A(n31851), .B(n31850), .Z(n31852) );
  NANDN U32041 ( .A(n31543), .B(n31542), .Z(n31547) );
  OR U32042 ( .A(n31545), .B(n31544), .Z(n31546) );
  NAND U32043 ( .A(n31547), .B(n31546), .Z(n31853) );
  XNOR U32044 ( .A(n31852), .B(n31853), .Z(n31941) );
  NANDN U32045 ( .A(n37974), .B(n31548), .Z(n31550) );
  XOR U32046 ( .A(b[57]), .B(a[84]), .Z(n31820) );
  NANDN U32047 ( .A(n38031), .B(n31820), .Z(n31549) );
  AND U32048 ( .A(n31550), .B(n31549), .Z(n31747) );
  NANDN U32049 ( .A(n34223), .B(n31551), .Z(n31553) );
  XOR U32050 ( .A(a[114]), .B(b[27]), .Z(n31922) );
  NANDN U32051 ( .A(n34458), .B(n31922), .Z(n31552) );
  AND U32052 ( .A(n31553), .B(n31552), .Z(n31746) );
  NANDN U32053 ( .A(n35936), .B(n31554), .Z(n31556) );
  XOR U32054 ( .A(a[104]), .B(b[37]), .Z(n31919) );
  NANDN U32055 ( .A(n36047), .B(n31919), .Z(n31555) );
  NAND U32056 ( .A(n31556), .B(n31555), .Z(n31745) );
  XOR U32057 ( .A(n31746), .B(n31745), .Z(n31748) );
  XOR U32058 ( .A(n31747), .B(n31748), .Z(n31845) );
  NANDN U32059 ( .A(n33866), .B(n31557), .Z(n31559) );
  XOR U32060 ( .A(a[118]), .B(b[23]), .Z(n31793) );
  NANDN U32061 ( .A(n33644), .B(n31793), .Z(n31558) );
  AND U32062 ( .A(n31559), .B(n31558), .Z(n31768) );
  NANDN U32063 ( .A(n32996), .B(n31560), .Z(n31562) );
  XOR U32064 ( .A(a[120]), .B(b[21]), .Z(n31787) );
  NANDN U32065 ( .A(n33271), .B(n31787), .Z(n31561) );
  AND U32066 ( .A(n31562), .B(n31561), .Z(n31767) );
  NANDN U32067 ( .A(n211), .B(n31563), .Z(n31565) );
  XOR U32068 ( .A(b[47]), .B(a[94]), .Z(n31751) );
  NANDN U32069 ( .A(n37172), .B(n31751), .Z(n31564) );
  NAND U32070 ( .A(n31565), .B(n31564), .Z(n31766) );
  XOR U32071 ( .A(n31767), .B(n31766), .Z(n31769) );
  XNOR U32072 ( .A(n31768), .B(n31769), .Z(n31844) );
  XNOR U32073 ( .A(n31845), .B(n31844), .Z(n31846) );
  NANDN U32074 ( .A(n31567), .B(n31566), .Z(n31571) );
  OR U32075 ( .A(n31569), .B(n31568), .Z(n31570) );
  NAND U32076 ( .A(n31571), .B(n31570), .Z(n31847) );
  XOR U32077 ( .A(n31846), .B(n31847), .Z(n31942) );
  XOR U32078 ( .A(n31941), .B(n31942), .Z(n31944) );
  XOR U32079 ( .A(n31943), .B(n31944), .Z(n31889) );
  NANDN U32080 ( .A(n31573), .B(n31572), .Z(n31577) );
  NAND U32081 ( .A(n31575), .B(n31574), .Z(n31576) );
  AND U32082 ( .A(n31577), .B(n31576), .Z(n31886) );
  NANDN U32083 ( .A(n35611), .B(n31578), .Z(n31580) );
  XOR U32084 ( .A(a[106]), .B(b[35]), .Z(n31823) );
  NANDN U32085 ( .A(n35801), .B(n31823), .Z(n31579) );
  AND U32086 ( .A(n31580), .B(n31579), .Z(n31834) );
  NANDN U32087 ( .A(n35260), .B(n31581), .Z(n31583) );
  XOR U32088 ( .A(a[108]), .B(b[33]), .Z(n31910) );
  NANDN U32089 ( .A(n35456), .B(n31910), .Z(n31582) );
  AND U32090 ( .A(n31583), .B(n31582), .Z(n31833) );
  NANDN U32091 ( .A(n36210), .B(n31584), .Z(n31586) );
  XOR U32092 ( .A(b[39]), .B(a[102]), .Z(n31763) );
  NANDN U32093 ( .A(n36347), .B(n31763), .Z(n31585) );
  NAND U32094 ( .A(n31586), .B(n31585), .Z(n31832) );
  XOR U32095 ( .A(n31833), .B(n31832), .Z(n31835) );
  XOR U32096 ( .A(n31834), .B(n31835), .Z(n31905) );
  NANDN U32097 ( .A(n31588), .B(n31587), .Z(n31592) );
  NANDN U32098 ( .A(n31590), .B(n31589), .Z(n31591) );
  AND U32099 ( .A(n31592), .B(n31591), .Z(n31904) );
  XNOR U32100 ( .A(n31905), .B(n31904), .Z(n31907) );
  NANDN U32101 ( .A(n31594), .B(n31593), .Z(n31598) );
  OR U32102 ( .A(n31596), .B(n31595), .Z(n31597) );
  AND U32103 ( .A(n31598), .B(n31597), .Z(n31906) );
  XOR U32104 ( .A(n31907), .B(n31906), .Z(n31901) );
  NANDN U32105 ( .A(n31600), .B(n31599), .Z(n31604) );
  OR U32106 ( .A(n31602), .B(n31601), .Z(n31603) );
  AND U32107 ( .A(n31604), .B(n31603), .Z(n31899) );
  NANDN U32108 ( .A(n31606), .B(n31605), .Z(n31610) );
  NAND U32109 ( .A(n31608), .B(n31607), .Z(n31609) );
  NAND U32110 ( .A(n31610), .B(n31609), .Z(n31898) );
  XNOR U32111 ( .A(n31899), .B(n31898), .Z(n31900) );
  XOR U32112 ( .A(n31901), .B(n31900), .Z(n31887) );
  XNOR U32113 ( .A(n31886), .B(n31887), .Z(n31888) );
  XOR U32114 ( .A(n31889), .B(n31888), .Z(n31734) );
  XNOR U32115 ( .A(n31733), .B(n31734), .Z(n31736) );
  NANDN U32116 ( .A(n31612), .B(n31611), .Z(n31616) );
  NANDN U32117 ( .A(n31614), .B(n31613), .Z(n31615) );
  AND U32118 ( .A(n31616), .B(n31615), .Z(n31882) );
  NANDN U32119 ( .A(n31618), .B(n31617), .Z(n31622) );
  NANDN U32120 ( .A(n31620), .B(n31619), .Z(n31621) );
  AND U32121 ( .A(n31622), .B(n31621), .Z(n31880) );
  NANDN U32122 ( .A(n31624), .B(n31623), .Z(n31628) );
  NAND U32123 ( .A(n31626), .B(n31625), .Z(n31627) );
  NAND U32124 ( .A(n31628), .B(n31627), .Z(n31881) );
  XOR U32125 ( .A(n31880), .B(n31881), .Z(n31883) );
  XNOR U32126 ( .A(n31882), .B(n31883), .Z(n31735) );
  XOR U32127 ( .A(n31736), .B(n31735), .Z(n31875) );
  NANDN U32128 ( .A(n31630), .B(n31629), .Z(n31634) );
  NAND U32129 ( .A(n31632), .B(n31631), .Z(n31633) );
  NAND U32130 ( .A(n31634), .B(n31633), .Z(n31874) );
  XNOR U32131 ( .A(n31875), .B(n31874), .Z(n31877) );
  NANDN U32132 ( .A(n31636), .B(n31635), .Z(n31640) );
  NANDN U32133 ( .A(n31638), .B(n31637), .Z(n31639) );
  AND U32134 ( .A(n31640), .B(n31639), .Z(n31876) );
  XOR U32135 ( .A(n31877), .B(n31876), .Z(n31729) );
  NANDN U32136 ( .A(n31642), .B(n31641), .Z(n31646) );
  NAND U32137 ( .A(n31644), .B(n31643), .Z(n31645) );
  AND U32138 ( .A(n31646), .B(n31645), .Z(n31728) );
  NANDN U32139 ( .A(n31648), .B(n31647), .Z(n31652) );
  NAND U32140 ( .A(n31650), .B(n31649), .Z(n31651) );
  AND U32141 ( .A(n31652), .B(n31651), .Z(n31869) );
  NANDN U32142 ( .A(n31654), .B(n31653), .Z(n31658) );
  NANDN U32143 ( .A(n31656), .B(n31655), .Z(n31657) );
  AND U32144 ( .A(n31658), .B(n31657), .Z(n31895) );
  NANDN U32145 ( .A(n31660), .B(n31659), .Z(n31664) );
  NANDN U32146 ( .A(n31662), .B(n31661), .Z(n31663) );
  AND U32147 ( .A(n31664), .B(n31663), .Z(n31893) );
  NANDN U32148 ( .A(n37705), .B(n31665), .Z(n31667) );
  XOR U32149 ( .A(b[53]), .B(a[88]), .Z(n31754) );
  NANDN U32150 ( .A(n37778), .B(n31754), .Z(n31666) );
  AND U32151 ( .A(n31667), .B(n31666), .Z(n31805) );
  NANDN U32152 ( .A(n37857), .B(n31668), .Z(n31670) );
  XOR U32153 ( .A(b[55]), .B(a[86]), .Z(n31817) );
  NANDN U32154 ( .A(n37911), .B(n31817), .Z(n31669) );
  AND U32155 ( .A(n31670), .B(n31669), .Z(n31803) );
  NANDN U32156 ( .A(n34634), .B(n31671), .Z(n31673) );
  XOR U32157 ( .A(a[112]), .B(b[29]), .Z(n31916) );
  NANDN U32158 ( .A(n34722), .B(n31916), .Z(n31672) );
  NAND U32159 ( .A(n31673), .B(n31672), .Z(n31802) );
  XNOR U32160 ( .A(n31803), .B(n31802), .Z(n31804) );
  XOR U32161 ( .A(n31805), .B(n31804), .Z(n31863) );
  NANDN U32162 ( .A(n38090), .B(n31674), .Z(n31676) );
  XOR U32163 ( .A(b[59]), .B(a[82]), .Z(n31796) );
  NANDN U32164 ( .A(n38130), .B(n31796), .Z(n31675) );
  AND U32165 ( .A(n31676), .B(n31675), .Z(n31780) );
  NANDN U32166 ( .A(n33875), .B(n31677), .Z(n31679) );
  XOR U32167 ( .A(a[116]), .B(b[25]), .Z(n31757) );
  NANDN U32168 ( .A(n33994), .B(n31757), .Z(n31678) );
  AND U32169 ( .A(n31679), .B(n31678), .Z(n31779) );
  NANDN U32170 ( .A(n37526), .B(n31680), .Z(n31682) );
  XOR U32171 ( .A(b[51]), .B(a[90]), .Z(n31799) );
  NANDN U32172 ( .A(n37605), .B(n31799), .Z(n31681) );
  NAND U32173 ( .A(n31682), .B(n31681), .Z(n31778) );
  XOR U32174 ( .A(n31779), .B(n31778), .Z(n31781) );
  XNOR U32175 ( .A(n31780), .B(n31781), .Z(n31862) );
  XOR U32176 ( .A(n31863), .B(n31862), .Z(n31865) );
  NANDN U32177 ( .A(n31684), .B(n31683), .Z(n31688) );
  OR U32178 ( .A(n31686), .B(n31685), .Z(n31687) );
  AND U32179 ( .A(n31688), .B(n31687), .Z(n31864) );
  XOR U32180 ( .A(n31865), .B(n31864), .Z(n31892) );
  XNOR U32181 ( .A(n31893), .B(n31892), .Z(n31894) );
  XNOR U32182 ( .A(n31895), .B(n31894), .Z(n31868) );
  XNOR U32183 ( .A(n31869), .B(n31868), .Z(n31871) );
  NANDN U32184 ( .A(n31690), .B(n31689), .Z(n31694) );
  OR U32185 ( .A(n31692), .B(n31691), .Z(n31693) );
  AND U32186 ( .A(n31694), .B(n31693), .Z(n31870) );
  XNOR U32187 ( .A(n31871), .B(n31870), .Z(n31727) );
  XOR U32188 ( .A(n31728), .B(n31727), .Z(n31730) );
  XOR U32189 ( .A(n31729), .B(n31730), .Z(n31724) );
  NANDN U32190 ( .A(n31696), .B(n31695), .Z(n31700) );
  NAND U32191 ( .A(n31698), .B(n31697), .Z(n31699) );
  AND U32192 ( .A(n31700), .B(n31699), .Z(n31722) );
  NANDN U32193 ( .A(n31702), .B(n31701), .Z(n31706) );
  NAND U32194 ( .A(n31704), .B(n31703), .Z(n31705) );
  NAND U32195 ( .A(n31706), .B(n31705), .Z(n31721) );
  XNOR U32196 ( .A(n31722), .B(n31721), .Z(n31723) );
  XOR U32197 ( .A(n31724), .B(n31723), .Z(n31716) );
  XNOR U32198 ( .A(n31715), .B(n31716), .Z(n31717) );
  XNOR U32199 ( .A(n31718), .B(n31717), .Z(n31709) );
  XOR U32200 ( .A(n31710), .B(n31709), .Z(n31712) );
  XNOR U32201 ( .A(n31711), .B(n31712), .Z(n31707) );
  XOR U32202 ( .A(n31708), .B(n31707), .Z(c[204]) );
  AND U32203 ( .A(n31708), .B(n31707), .Z(n31948) );
  NANDN U32204 ( .A(n31710), .B(n31709), .Z(n31714) );
  OR U32205 ( .A(n31712), .B(n31711), .Z(n31713) );
  AND U32206 ( .A(n31714), .B(n31713), .Z(n31951) );
  NANDN U32207 ( .A(n31716), .B(n31715), .Z(n31720) );
  NANDN U32208 ( .A(n31718), .B(n31717), .Z(n31719) );
  AND U32209 ( .A(n31720), .B(n31719), .Z(n31950) );
  NANDN U32210 ( .A(n31722), .B(n31721), .Z(n31726) );
  NANDN U32211 ( .A(n31724), .B(n31723), .Z(n31725) );
  AND U32212 ( .A(n31726), .B(n31725), .Z(n31958) );
  NANDN U32213 ( .A(n31728), .B(n31727), .Z(n31732) );
  OR U32214 ( .A(n31730), .B(n31729), .Z(n31731) );
  AND U32215 ( .A(n31732), .B(n31731), .Z(n31955) );
  NANDN U32216 ( .A(n31734), .B(n31733), .Z(n31738) );
  NAND U32217 ( .A(n31736), .B(n31735), .Z(n31737) );
  AND U32218 ( .A(n31738), .B(n31737), .Z(n32178) );
  NANDN U32219 ( .A(n31740), .B(n31739), .Z(n31744) );
  OR U32220 ( .A(n31742), .B(n31741), .Z(n31743) );
  AND U32221 ( .A(n31744), .B(n31743), .Z(n32159) );
  NANDN U32222 ( .A(n31746), .B(n31745), .Z(n31750) );
  OR U32223 ( .A(n31748), .B(n31747), .Z(n31749) );
  NAND U32224 ( .A(n31750), .B(n31749), .Z(n32160) );
  XNOR U32225 ( .A(n32159), .B(n32160), .Z(n32162) );
  NANDN U32226 ( .A(n211), .B(n31751), .Z(n31753) );
  XOR U32227 ( .A(b[47]), .B(a[95]), .Z(n32051) );
  NANDN U32228 ( .A(n37172), .B(n32051), .Z(n31752) );
  AND U32229 ( .A(n31753), .B(n31752), .Z(n32068) );
  NANDN U32230 ( .A(n37705), .B(n31754), .Z(n31756) );
  XOR U32231 ( .A(b[53]), .B(a[89]), .Z(n32054) );
  NANDN U32232 ( .A(n37778), .B(n32054), .Z(n31755) );
  AND U32233 ( .A(n31756), .B(n31755), .Z(n32067) );
  NANDN U32234 ( .A(n33875), .B(n31757), .Z(n31759) );
  XOR U32235 ( .A(a[117]), .B(b[25]), .Z(n31976) );
  NANDN U32236 ( .A(n33994), .B(n31976), .Z(n31758) );
  NAND U32237 ( .A(n31759), .B(n31758), .Z(n32066) );
  XOR U32238 ( .A(n32067), .B(n32066), .Z(n32069) );
  XOR U32239 ( .A(n32068), .B(n32069), .Z(n32073) );
  NANDN U32240 ( .A(n36480), .B(n31760), .Z(n31762) );
  XOR U32241 ( .A(b[41]), .B(a[101]), .Z(n32016) );
  NANDN U32242 ( .A(n36594), .B(n32016), .Z(n31761) );
  NAND U32243 ( .A(n31762), .B(n31761), .Z(n32141) );
  XNOR U32244 ( .A(n32142), .B(n32141), .Z(n32144) );
  NANDN U32245 ( .A(n36210), .B(n31763), .Z(n31765) );
  XOR U32246 ( .A(b[39]), .B(a[103]), .Z(n31973) );
  NANDN U32247 ( .A(n36347), .B(n31973), .Z(n31764) );
  AND U32248 ( .A(n31765), .B(n31764), .Z(n32061) );
  AND U32249 ( .A(b[63]), .B(a[77]), .Z(n32060) );
  XOR U32250 ( .A(n32061), .B(n32060), .Z(n32063) );
  XOR U32251 ( .A(n31935), .B(n32063), .Z(n32143) );
  XNOR U32252 ( .A(n32144), .B(n32143), .Z(n32072) );
  XNOR U32253 ( .A(n32073), .B(n32072), .Z(n32074) );
  NANDN U32254 ( .A(n31767), .B(n31766), .Z(n31771) );
  OR U32255 ( .A(n31769), .B(n31768), .Z(n31770) );
  NAND U32256 ( .A(n31771), .B(n31770), .Z(n32075) );
  XNOR U32257 ( .A(n32074), .B(n32075), .Z(n32161) );
  XOR U32258 ( .A(n32162), .B(n32161), .Z(n32085) );
  NAND U32259 ( .A(n31773), .B(n31772), .Z(n31777) );
  NAND U32260 ( .A(n31775), .B(n31774), .Z(n31776) );
  AND U32261 ( .A(n31777), .B(n31776), .Z(n32084) );
  XNOR U32262 ( .A(n32085), .B(n32084), .Z(n32086) );
  NANDN U32263 ( .A(n31779), .B(n31778), .Z(n31783) );
  OR U32264 ( .A(n31781), .B(n31780), .Z(n31782) );
  AND U32265 ( .A(n31783), .B(n31782), .Z(n32097) );
  NANDN U32266 ( .A(n38247), .B(n31784), .Z(n31786) );
  XOR U32267 ( .A(b[61]), .B(a[81]), .Z(n31979) );
  NANDN U32268 ( .A(n38248), .B(n31979), .Z(n31785) );
  AND U32269 ( .A(n31786), .B(n31785), .Z(n32035) );
  NANDN U32270 ( .A(n32996), .B(n31787), .Z(n31789) );
  XOR U32271 ( .A(a[121]), .B(b[21]), .Z(n32135) );
  NANDN U32272 ( .A(n33271), .B(n32135), .Z(n31788) );
  AND U32273 ( .A(n31789), .B(n31788), .Z(n32034) );
  NANDN U32274 ( .A(n212), .B(n31790), .Z(n31792) );
  XOR U32275 ( .A(b[49]), .B(a[93]), .Z(n31982) );
  NANDN U32276 ( .A(n37432), .B(n31982), .Z(n31791) );
  NAND U32277 ( .A(n31792), .B(n31791), .Z(n32033) );
  XOR U32278 ( .A(n32034), .B(n32033), .Z(n32036) );
  XOR U32279 ( .A(n32035), .B(n32036), .Z(n32154) );
  NANDN U32280 ( .A(n33866), .B(n31793), .Z(n31795) );
  XOR U32281 ( .A(a[119]), .B(b[23]), .Z(n32132) );
  NANDN U32282 ( .A(n33644), .B(n32132), .Z(n31794) );
  AND U32283 ( .A(n31795), .B(n31794), .Z(n32149) );
  NANDN U32284 ( .A(n38090), .B(n31796), .Z(n31798) );
  XOR U32285 ( .A(b[59]), .B(a[83]), .Z(n32126) );
  NANDN U32286 ( .A(n38130), .B(n32126), .Z(n31797) );
  AND U32287 ( .A(n31798), .B(n31797), .Z(n32148) );
  NANDN U32288 ( .A(n37526), .B(n31799), .Z(n31801) );
  XOR U32289 ( .A(b[51]), .B(a[91]), .Z(n32129) );
  NANDN U32290 ( .A(n37605), .B(n32129), .Z(n31800) );
  NAND U32291 ( .A(n31801), .B(n31800), .Z(n32147) );
  XOR U32292 ( .A(n32148), .B(n32147), .Z(n32150) );
  XNOR U32293 ( .A(n32149), .B(n32150), .Z(n32153) );
  XNOR U32294 ( .A(n32154), .B(n32153), .Z(n32156) );
  NANDN U32295 ( .A(n31803), .B(n31802), .Z(n31807) );
  NANDN U32296 ( .A(n31805), .B(n31804), .Z(n31806) );
  AND U32297 ( .A(n31807), .B(n31806), .Z(n32155) );
  XNOR U32298 ( .A(n32156), .B(n32155), .Z(n32096) );
  XNOR U32299 ( .A(n32097), .B(n32096), .Z(n32098) );
  NANDN U32300 ( .A(n32483), .B(n31808), .Z(n31810) );
  XOR U32301 ( .A(a[123]), .B(b[19]), .Z(n32009) );
  NANDN U32302 ( .A(n32823), .B(n32009), .Z(n31809) );
  AND U32303 ( .A(n31810), .B(n31809), .Z(n31993) );
  NANDN U32304 ( .A(n32013), .B(n31811), .Z(n31813) );
  XOR U32305 ( .A(a[125]), .B(b[17]), .Z(n32012) );
  NANDN U32306 ( .A(n32292), .B(n32012), .Z(n31812) );
  AND U32307 ( .A(n31813), .B(n31812), .Z(n31992) );
  NANDN U32308 ( .A(n36991), .B(n31814), .Z(n31816) );
  XOR U32309 ( .A(b[45]), .B(a[97]), .Z(n32138) );
  NANDN U32310 ( .A(n37083), .B(n32138), .Z(n31815) );
  NAND U32311 ( .A(n31816), .B(n31815), .Z(n31991) );
  XOR U32312 ( .A(n31992), .B(n31991), .Z(n31994) );
  XOR U32313 ( .A(n31993), .B(n31994), .Z(n32079) );
  NANDN U32314 ( .A(n37857), .B(n31817), .Z(n31819) );
  XOR U32315 ( .A(b[55]), .B(a[87]), .Z(n31967) );
  NANDN U32316 ( .A(n37911), .B(n31967), .Z(n31818) );
  AND U32317 ( .A(n31819), .B(n31818), .Z(n31987) );
  NANDN U32318 ( .A(n37974), .B(n31820), .Z(n31822) );
  XOR U32319 ( .A(b[57]), .B(a[85]), .Z(n31970) );
  NANDN U32320 ( .A(n38031), .B(n31970), .Z(n31821) );
  AND U32321 ( .A(n31822), .B(n31821), .Z(n31986) );
  NANDN U32322 ( .A(n35611), .B(n31823), .Z(n31825) );
  XOR U32323 ( .A(a[107]), .B(b[35]), .Z(n32108) );
  NANDN U32324 ( .A(n35801), .B(n32108), .Z(n31824) );
  NAND U32325 ( .A(n31825), .B(n31824), .Z(n31985) );
  XOR U32326 ( .A(n31986), .B(n31985), .Z(n31988) );
  XNOR U32327 ( .A(n31987), .B(n31988), .Z(n32078) );
  XNOR U32328 ( .A(n32079), .B(n32078), .Z(n32081) );
  NANDN U32329 ( .A(n31827), .B(n31826), .Z(n31831) );
  NANDN U32330 ( .A(n31829), .B(n31828), .Z(n31830) );
  AND U32331 ( .A(n31831), .B(n31830), .Z(n32080) );
  XOR U32332 ( .A(n32081), .B(n32080), .Z(n32105) );
  NANDN U32333 ( .A(n31833), .B(n31832), .Z(n31837) );
  OR U32334 ( .A(n31835), .B(n31834), .Z(n31836) );
  AND U32335 ( .A(n31837), .B(n31836), .Z(n32103) );
  NANDN U32336 ( .A(n31839), .B(n31838), .Z(n31843) );
  OR U32337 ( .A(n31841), .B(n31840), .Z(n31842) );
  NAND U32338 ( .A(n31843), .B(n31842), .Z(n32102) );
  XNOR U32339 ( .A(n32103), .B(n32102), .Z(n32104) );
  XOR U32340 ( .A(n32105), .B(n32104), .Z(n32099) );
  XOR U32341 ( .A(n32098), .B(n32099), .Z(n32087) );
  XNOR U32342 ( .A(n32086), .B(n32087), .Z(n32173) );
  NANDN U32343 ( .A(n31845), .B(n31844), .Z(n31849) );
  NANDN U32344 ( .A(n31847), .B(n31846), .Z(n31848) );
  AND U32345 ( .A(n31849), .B(n31848), .Z(n32091) );
  NANDN U32346 ( .A(n31851), .B(n31850), .Z(n31855) );
  NANDN U32347 ( .A(n31853), .B(n31852), .Z(n31854) );
  NAND U32348 ( .A(n31855), .B(n31854), .Z(n32090) );
  XNOR U32349 ( .A(n32091), .B(n32090), .Z(n32093) );
  NANDN U32350 ( .A(n31857), .B(n31856), .Z(n31861) );
  OR U32351 ( .A(n31859), .B(n31858), .Z(n31860) );
  AND U32352 ( .A(n31861), .B(n31860), .Z(n32092) );
  XOR U32353 ( .A(n32093), .B(n32092), .Z(n32172) );
  NAND U32354 ( .A(n31863), .B(n31862), .Z(n31867) );
  NAND U32355 ( .A(n31865), .B(n31864), .Z(n31866) );
  AND U32356 ( .A(n31867), .B(n31866), .Z(n32171) );
  XOR U32357 ( .A(n32172), .B(n32171), .Z(n32174) );
  XNOR U32358 ( .A(n32173), .B(n32174), .Z(n32177) );
  XNOR U32359 ( .A(n32178), .B(n32177), .Z(n32180) );
  NANDN U32360 ( .A(n31869), .B(n31868), .Z(n31873) );
  NAND U32361 ( .A(n31871), .B(n31870), .Z(n31872) );
  AND U32362 ( .A(n31873), .B(n31872), .Z(n32179) );
  XOR U32363 ( .A(n32180), .B(n32179), .Z(n32186) );
  NANDN U32364 ( .A(n31875), .B(n31874), .Z(n31879) );
  NAND U32365 ( .A(n31877), .B(n31876), .Z(n31878) );
  AND U32366 ( .A(n31879), .B(n31878), .Z(n32184) );
  NANDN U32367 ( .A(n31881), .B(n31880), .Z(n31885) );
  NANDN U32368 ( .A(n31883), .B(n31882), .Z(n31884) );
  AND U32369 ( .A(n31885), .B(n31884), .Z(n32167) );
  NANDN U32370 ( .A(n31887), .B(n31886), .Z(n31891) );
  NANDN U32371 ( .A(n31889), .B(n31888), .Z(n31890) );
  AND U32372 ( .A(n31891), .B(n31890), .Z(n32166) );
  NANDN U32373 ( .A(n31893), .B(n31892), .Z(n31897) );
  NANDN U32374 ( .A(n31895), .B(n31894), .Z(n31896) );
  AND U32375 ( .A(n31897), .B(n31896), .Z(n31963) );
  NANDN U32376 ( .A(n31899), .B(n31898), .Z(n31903) );
  NANDN U32377 ( .A(n31901), .B(n31900), .Z(n31902) );
  AND U32378 ( .A(n31903), .B(n31902), .Z(n32048) );
  NANDN U32379 ( .A(n31905), .B(n31904), .Z(n31909) );
  NAND U32380 ( .A(n31907), .B(n31906), .Z(n31908) );
  AND U32381 ( .A(n31909), .B(n31908), .Z(n32046) );
  NANDN U32382 ( .A(n35260), .B(n31910), .Z(n31912) );
  XOR U32383 ( .A(a[109]), .B(b[33]), .Z(n32114) );
  NANDN U32384 ( .A(n35456), .B(n32114), .Z(n31911) );
  AND U32385 ( .A(n31912), .B(n31911), .Z(n31999) );
  NANDN U32386 ( .A(n34909), .B(n31913), .Z(n31915) );
  XOR U32387 ( .A(a[111]), .B(b[31]), .Z(n32120) );
  NANDN U32388 ( .A(n35145), .B(n32120), .Z(n31914) );
  AND U32389 ( .A(n31915), .B(n31914), .Z(n31998) );
  NANDN U32390 ( .A(n34634), .B(n31916), .Z(n31918) );
  XOR U32391 ( .A(a[113]), .B(b[29]), .Z(n32057) );
  NANDN U32392 ( .A(n34722), .B(n32057), .Z(n31917) );
  AND U32393 ( .A(n31918), .B(n31917), .Z(n32030) );
  NANDN U32394 ( .A(n35936), .B(n31919), .Z(n31921) );
  XOR U32395 ( .A(a[105]), .B(b[37]), .Z(n32111) );
  NANDN U32396 ( .A(n36047), .B(n32111), .Z(n31920) );
  AND U32397 ( .A(n31921), .B(n31920), .Z(n32028) );
  NANDN U32398 ( .A(n34223), .B(n31922), .Z(n31924) );
  XOR U32399 ( .A(a[115]), .B(b[27]), .Z(n32123) );
  NANDN U32400 ( .A(n34458), .B(n32123), .Z(n31923) );
  NAND U32401 ( .A(n31924), .B(n31923), .Z(n32027) );
  XNOR U32402 ( .A(n32028), .B(n32027), .Z(n32029) );
  XNOR U32403 ( .A(n32030), .B(n32029), .Z(n31997) );
  XOR U32404 ( .A(n31998), .B(n31997), .Z(n32000) );
  XOR U32405 ( .A(n31999), .B(n32000), .Z(n32006) );
  XNOR U32406 ( .A(a[127]), .B(b[15]), .Z(n32022) );
  OR U32407 ( .A(n32022), .B(n31925), .Z(n31928) );
  NAND U32408 ( .A(n32023), .B(n31926), .Z(n31927) );
  AND U32409 ( .A(n31928), .B(n31927), .Z(n32041) );
  NANDN U32410 ( .A(n38278), .B(n31929), .Z(n31931) );
  XOR U32411 ( .A(b[63]), .B(a[79]), .Z(n32019) );
  NANDN U32412 ( .A(n38279), .B(n32019), .Z(n31930) );
  AND U32413 ( .A(n31931), .B(n31930), .Z(n32040) );
  NANDN U32414 ( .A(n36742), .B(n31932), .Z(n31934) );
  XOR U32415 ( .A(b[43]), .B(a[99]), .Z(n32117) );
  NANDN U32416 ( .A(n36891), .B(n32117), .Z(n31933) );
  NAND U32417 ( .A(n31934), .B(n31933), .Z(n32039) );
  XOR U32418 ( .A(n32040), .B(n32039), .Z(n32042) );
  XOR U32419 ( .A(n32041), .B(n32042), .Z(n32004) );
  IV U32420 ( .A(n31935), .Z(n32062) );
  NANDN U32421 ( .A(n32062), .B(n31936), .Z(n31940) );
  NANDN U32422 ( .A(n31938), .B(n31937), .Z(n31939) );
  AND U32423 ( .A(n31940), .B(n31939), .Z(n32003) );
  XNOR U32424 ( .A(n32004), .B(n32003), .Z(n32005) );
  XNOR U32425 ( .A(n32006), .B(n32005), .Z(n32045) );
  XNOR U32426 ( .A(n32046), .B(n32045), .Z(n32047) );
  XOR U32427 ( .A(n32048), .B(n32047), .Z(n31962) );
  NANDN U32428 ( .A(n31942), .B(n31941), .Z(n31946) );
  OR U32429 ( .A(n31944), .B(n31943), .Z(n31945) );
  AND U32430 ( .A(n31946), .B(n31945), .Z(n31961) );
  XOR U32431 ( .A(n31962), .B(n31961), .Z(n31964) );
  XNOR U32432 ( .A(n31963), .B(n31964), .Z(n32165) );
  XOR U32433 ( .A(n32166), .B(n32165), .Z(n32168) );
  XNOR U32434 ( .A(n32167), .B(n32168), .Z(n32183) );
  XNOR U32435 ( .A(n32184), .B(n32183), .Z(n32185) );
  XOR U32436 ( .A(n32186), .B(n32185), .Z(n31956) );
  XNOR U32437 ( .A(n31955), .B(n31956), .Z(n31957) );
  XNOR U32438 ( .A(n31958), .B(n31957), .Z(n31949) );
  XOR U32439 ( .A(n31950), .B(n31949), .Z(n31952) );
  XNOR U32440 ( .A(n31951), .B(n31952), .Z(n31947) );
  XOR U32441 ( .A(n31948), .B(n31947), .Z(c[205]) );
  AND U32442 ( .A(n31948), .B(n31947), .Z(n32190) );
  NANDN U32443 ( .A(n31950), .B(n31949), .Z(n31954) );
  OR U32444 ( .A(n31952), .B(n31951), .Z(n31953) );
  AND U32445 ( .A(n31954), .B(n31953), .Z(n32193) );
  NANDN U32446 ( .A(n31956), .B(n31955), .Z(n31960) );
  NANDN U32447 ( .A(n31958), .B(n31957), .Z(n31959) );
  AND U32448 ( .A(n31960), .B(n31959), .Z(n32192) );
  NANDN U32449 ( .A(n31962), .B(n31961), .Z(n31966) );
  NANDN U32450 ( .A(n31964), .B(n31963), .Z(n31965) );
  AND U32451 ( .A(n31966), .B(n31965), .Z(n32211) );
  NANDN U32452 ( .A(n37857), .B(n31967), .Z(n31969) );
  XOR U32453 ( .A(b[55]), .B(a[88]), .Z(n32384) );
  NANDN U32454 ( .A(n37911), .B(n32384), .Z(n31968) );
  AND U32455 ( .A(n31969), .B(n31968), .Z(n32356) );
  NANDN U32456 ( .A(n37974), .B(n31970), .Z(n31972) );
  XOR U32457 ( .A(b[57]), .B(a[86]), .Z(n32345) );
  NANDN U32458 ( .A(n38031), .B(n32345), .Z(n31971) );
  AND U32459 ( .A(n31972), .B(n31971), .Z(n32355) );
  NANDN U32460 ( .A(n36210), .B(n31973), .Z(n31975) );
  XOR U32461 ( .A(a[104]), .B(b[39]), .Z(n32318) );
  NANDN U32462 ( .A(n36347), .B(n32318), .Z(n31974) );
  NAND U32463 ( .A(n31975), .B(n31974), .Z(n32354) );
  XOR U32464 ( .A(n32355), .B(n32354), .Z(n32357) );
  XOR U32465 ( .A(n32356), .B(n32357), .Z(n32252) );
  NANDN U32466 ( .A(n33875), .B(n31976), .Z(n31978) );
  XOR U32467 ( .A(a[118]), .B(b[25]), .Z(n32306) );
  NANDN U32468 ( .A(n33994), .B(n32306), .Z(n31977) );
  AND U32469 ( .A(n31978), .B(n31977), .Z(n32398) );
  NANDN U32470 ( .A(n38247), .B(n31979), .Z(n31981) );
  XOR U32471 ( .A(b[61]), .B(a[82]), .Z(n32339) );
  NANDN U32472 ( .A(n38248), .B(n32339), .Z(n31980) );
  AND U32473 ( .A(n31981), .B(n31980), .Z(n32397) );
  NANDN U32474 ( .A(n212), .B(n31982), .Z(n31984) );
  XOR U32475 ( .A(b[49]), .B(a[94]), .Z(n32300) );
  NANDN U32476 ( .A(n37432), .B(n32300), .Z(n31983) );
  NAND U32477 ( .A(n31984), .B(n31983), .Z(n32396) );
  XOR U32478 ( .A(n32397), .B(n32396), .Z(n32399) );
  XNOR U32479 ( .A(n32398), .B(n32399), .Z(n32251) );
  XNOR U32480 ( .A(n32252), .B(n32251), .Z(n32253) );
  NANDN U32481 ( .A(n31986), .B(n31985), .Z(n31990) );
  OR U32482 ( .A(n31988), .B(n31987), .Z(n31989) );
  NAND U32483 ( .A(n31990), .B(n31989), .Z(n32254) );
  XNOR U32484 ( .A(n32253), .B(n32254), .Z(n32227) );
  NANDN U32485 ( .A(n31992), .B(n31991), .Z(n31996) );
  OR U32486 ( .A(n31994), .B(n31993), .Z(n31995) );
  NAND U32487 ( .A(n31996), .B(n31995), .Z(n32228) );
  XNOR U32488 ( .A(n32227), .B(n32228), .Z(n32230) );
  NANDN U32489 ( .A(n31998), .B(n31997), .Z(n32002) );
  OR U32490 ( .A(n32000), .B(n31999), .Z(n32001) );
  AND U32491 ( .A(n32002), .B(n32001), .Z(n32229) );
  XOR U32492 ( .A(n32230), .B(n32229), .Z(n32259) );
  NANDN U32493 ( .A(n32004), .B(n32003), .Z(n32008) );
  NANDN U32494 ( .A(n32006), .B(n32005), .Z(n32007) );
  AND U32495 ( .A(n32008), .B(n32007), .Z(n32257) );
  NANDN U32496 ( .A(n32483), .B(n32009), .Z(n32011) );
  XOR U32497 ( .A(a[124]), .B(b[19]), .Z(n32372) );
  NANDN U32498 ( .A(n32823), .B(n32372), .Z(n32010) );
  AND U32499 ( .A(n32011), .B(n32010), .Z(n32404) );
  NANDN U32500 ( .A(n32013), .B(n32012), .Z(n32015) );
  XOR U32501 ( .A(a[126]), .B(b[17]), .Z(n32293) );
  NANDN U32502 ( .A(n32292), .B(n32293), .Z(n32014) );
  AND U32503 ( .A(n32015), .B(n32014), .Z(n32403) );
  NANDN U32504 ( .A(n36480), .B(n32016), .Z(n32018) );
  XOR U32505 ( .A(b[41]), .B(a[102]), .Z(n32296) );
  NANDN U32506 ( .A(n36594), .B(n32296), .Z(n32017) );
  NAND U32507 ( .A(n32018), .B(n32017), .Z(n32402) );
  XOR U32508 ( .A(n32403), .B(n32402), .Z(n32405) );
  XOR U32509 ( .A(n32404), .B(n32405), .Z(n32409) );
  NANDN U32510 ( .A(n38278), .B(n32019), .Z(n32021) );
  XOR U32511 ( .A(b[63]), .B(a[80]), .Z(n32375) );
  NANDN U32512 ( .A(n38279), .B(n32375), .Z(n32020) );
  AND U32513 ( .A(n32021), .B(n32020), .Z(n32283) );
  NAND U32514 ( .A(b[63]), .B(a[78]), .Z(n32299) );
  ANDN U32515 ( .B(n32023), .A(n32022), .Z(n32026) );
  NAND U32516 ( .A(b[15]), .B(n32024), .Z(n32025) );
  NANDN U32517 ( .A(n32026), .B(n32025), .Z(n32281) );
  XOR U32518 ( .A(n32299), .B(n32281), .Z(n32282) );
  XOR U32519 ( .A(n32283), .B(n32282), .Z(n32408) );
  XNOR U32520 ( .A(n32409), .B(n32408), .Z(n32411) );
  NANDN U32521 ( .A(n32028), .B(n32027), .Z(n32032) );
  NANDN U32522 ( .A(n32030), .B(n32029), .Z(n32031) );
  AND U32523 ( .A(n32032), .B(n32031), .Z(n32410) );
  XOR U32524 ( .A(n32411), .B(n32410), .Z(n32242) );
  NANDN U32525 ( .A(n32034), .B(n32033), .Z(n32038) );
  OR U32526 ( .A(n32036), .B(n32035), .Z(n32037) );
  AND U32527 ( .A(n32038), .B(n32037), .Z(n32240) );
  NANDN U32528 ( .A(n32040), .B(n32039), .Z(n32044) );
  OR U32529 ( .A(n32042), .B(n32041), .Z(n32043) );
  NAND U32530 ( .A(n32044), .B(n32043), .Z(n32239) );
  XNOR U32531 ( .A(n32240), .B(n32239), .Z(n32241) );
  XOR U32532 ( .A(n32242), .B(n32241), .Z(n32258) );
  XOR U32533 ( .A(n32257), .B(n32258), .Z(n32260) );
  XOR U32534 ( .A(n32259), .B(n32260), .Z(n32217) );
  NANDN U32535 ( .A(n32046), .B(n32045), .Z(n32050) );
  NAND U32536 ( .A(n32048), .B(n32047), .Z(n32049) );
  AND U32537 ( .A(n32050), .B(n32049), .Z(n32216) );
  NANDN U32538 ( .A(n211), .B(n32051), .Z(n32053) );
  XOR U32539 ( .A(b[47]), .B(a[96]), .Z(n32351) );
  NANDN U32540 ( .A(n37172), .B(n32351), .Z(n32052) );
  AND U32541 ( .A(n32053), .B(n32052), .Z(n32392) );
  NANDN U32542 ( .A(n37705), .B(n32054), .Z(n32056) );
  XOR U32543 ( .A(b[53]), .B(a[90]), .Z(n32387) );
  NANDN U32544 ( .A(n37778), .B(n32387), .Z(n32055) );
  AND U32545 ( .A(n32056), .B(n32055), .Z(n32391) );
  NANDN U32546 ( .A(n34634), .B(n32057), .Z(n32059) );
  XNOR U32547 ( .A(a[114]), .B(b[29]), .Z(n32333) );
  NANDN U32548 ( .A(n32333), .B(n35002), .Z(n32058) );
  NAND U32549 ( .A(n32059), .B(n32058), .Z(n32390) );
  XOR U32550 ( .A(n32391), .B(n32390), .Z(n32393) );
  XOR U32551 ( .A(n32392), .B(n32393), .Z(n32310) );
  NANDN U32552 ( .A(n32061), .B(n32060), .Z(n32065) );
  NANDN U32553 ( .A(n32063), .B(n32062), .Z(n32064) );
  AND U32554 ( .A(n32065), .B(n32064), .Z(n32309) );
  XNOR U32555 ( .A(n32310), .B(n32309), .Z(n32312) );
  NANDN U32556 ( .A(n32067), .B(n32066), .Z(n32071) );
  OR U32557 ( .A(n32069), .B(n32068), .Z(n32070) );
  AND U32558 ( .A(n32071), .B(n32070), .Z(n32311) );
  XOR U32559 ( .A(n32312), .B(n32311), .Z(n32270) );
  NANDN U32560 ( .A(n32073), .B(n32072), .Z(n32077) );
  NANDN U32561 ( .A(n32075), .B(n32074), .Z(n32076) );
  AND U32562 ( .A(n32077), .B(n32076), .Z(n32269) );
  XNOR U32563 ( .A(n32270), .B(n32269), .Z(n32272) );
  NANDN U32564 ( .A(n32079), .B(n32078), .Z(n32083) );
  NAND U32565 ( .A(n32081), .B(n32080), .Z(n32082) );
  AND U32566 ( .A(n32083), .B(n32082), .Z(n32271) );
  XNOR U32567 ( .A(n32272), .B(n32271), .Z(n32215) );
  XOR U32568 ( .A(n32216), .B(n32215), .Z(n32218) );
  XOR U32569 ( .A(n32217), .B(n32218), .Z(n32210) );
  NANDN U32570 ( .A(n32085), .B(n32084), .Z(n32089) );
  NANDN U32571 ( .A(n32087), .B(n32086), .Z(n32088) );
  AND U32572 ( .A(n32089), .B(n32088), .Z(n32415) );
  NANDN U32573 ( .A(n32091), .B(n32090), .Z(n32095) );
  NAND U32574 ( .A(n32093), .B(n32092), .Z(n32094) );
  AND U32575 ( .A(n32095), .B(n32094), .Z(n32414) );
  XNOR U32576 ( .A(n32415), .B(n32414), .Z(n32416) );
  NANDN U32577 ( .A(n32097), .B(n32096), .Z(n32101) );
  NANDN U32578 ( .A(n32099), .B(n32098), .Z(n32100) );
  AND U32579 ( .A(n32101), .B(n32100), .Z(n32224) );
  NANDN U32580 ( .A(n32103), .B(n32102), .Z(n32107) );
  NANDN U32581 ( .A(n32105), .B(n32104), .Z(n32106) );
  AND U32582 ( .A(n32107), .B(n32106), .Z(n32222) );
  NANDN U32583 ( .A(n35611), .B(n32108), .Z(n32110) );
  XOR U32584 ( .A(a[108]), .B(b[35]), .Z(n32327) );
  NANDN U32585 ( .A(n35801), .B(n32327), .Z(n32109) );
  AND U32586 ( .A(n32110), .B(n32109), .Z(n32368) );
  NANDN U32587 ( .A(n35936), .B(n32111), .Z(n32113) );
  XOR U32588 ( .A(a[106]), .B(b[37]), .Z(n32315) );
  NANDN U32589 ( .A(n36047), .B(n32315), .Z(n32112) );
  AND U32590 ( .A(n32113), .B(n32112), .Z(n32367) );
  NANDN U32591 ( .A(n35260), .B(n32114), .Z(n32116) );
  XOR U32592 ( .A(a[110]), .B(b[33]), .Z(n32330) );
  NANDN U32593 ( .A(n35456), .B(n32330), .Z(n32115) );
  AND U32594 ( .A(n32116), .B(n32115), .Z(n32289) );
  NANDN U32595 ( .A(n36742), .B(n32117), .Z(n32119) );
  XOR U32596 ( .A(b[43]), .B(a[100]), .Z(n32378) );
  NANDN U32597 ( .A(n36891), .B(n32378), .Z(n32118) );
  AND U32598 ( .A(n32119), .B(n32118), .Z(n32287) );
  NANDN U32599 ( .A(n34909), .B(n32120), .Z(n32122) );
  XOR U32600 ( .A(a[112]), .B(b[31]), .Z(n32324) );
  NANDN U32601 ( .A(n35145), .B(n32324), .Z(n32121) );
  NAND U32602 ( .A(n32122), .B(n32121), .Z(n32286) );
  XNOR U32603 ( .A(n32287), .B(n32286), .Z(n32288) );
  XNOR U32604 ( .A(n32289), .B(n32288), .Z(n32366) );
  XOR U32605 ( .A(n32367), .B(n32366), .Z(n32369) );
  XOR U32606 ( .A(n32368), .B(n32369), .Z(n32248) );
  NANDN U32607 ( .A(n34223), .B(n32123), .Z(n32125) );
  XOR U32608 ( .A(a[116]), .B(b[27]), .Z(n32321) );
  NANDN U32609 ( .A(n34458), .B(n32321), .Z(n32124) );
  AND U32610 ( .A(n32125), .B(n32124), .Z(n32277) );
  NANDN U32611 ( .A(n38090), .B(n32126), .Z(n32128) );
  XOR U32612 ( .A(b[59]), .B(a[84]), .Z(n32348) );
  NANDN U32613 ( .A(n38130), .B(n32348), .Z(n32127) );
  AND U32614 ( .A(n32128), .B(n32127), .Z(n32276) );
  NANDN U32615 ( .A(n37526), .B(n32129), .Z(n32131) );
  XOR U32616 ( .A(b[51]), .B(a[92]), .Z(n32303) );
  NANDN U32617 ( .A(n37605), .B(n32303), .Z(n32130) );
  NAND U32618 ( .A(n32131), .B(n32130), .Z(n32275) );
  XOR U32619 ( .A(n32276), .B(n32275), .Z(n32278) );
  XOR U32620 ( .A(n32277), .B(n32278), .Z(n32246) );
  NANDN U32621 ( .A(n33866), .B(n32132), .Z(n32134) );
  XOR U32622 ( .A(a[120]), .B(b[23]), .Z(n32381) );
  NANDN U32623 ( .A(n33644), .B(n32381), .Z(n32133) );
  AND U32624 ( .A(n32134), .B(n32133), .Z(n32362) );
  NANDN U32625 ( .A(n32996), .B(n32135), .Z(n32137) );
  XOR U32626 ( .A(a[122]), .B(b[21]), .Z(n32336) );
  NANDN U32627 ( .A(n33271), .B(n32336), .Z(n32136) );
  AND U32628 ( .A(n32137), .B(n32136), .Z(n32361) );
  NANDN U32629 ( .A(n36991), .B(n32138), .Z(n32140) );
  XOR U32630 ( .A(b[45]), .B(a[98]), .Z(n32342) );
  NANDN U32631 ( .A(n37083), .B(n32342), .Z(n32139) );
  NAND U32632 ( .A(n32140), .B(n32139), .Z(n32360) );
  XOR U32633 ( .A(n32361), .B(n32360), .Z(n32363) );
  XNOR U32634 ( .A(n32362), .B(n32363), .Z(n32245) );
  XNOR U32635 ( .A(n32246), .B(n32245), .Z(n32247) );
  XNOR U32636 ( .A(n32248), .B(n32247), .Z(n32236) );
  NANDN U32637 ( .A(n32142), .B(n32141), .Z(n32146) );
  NAND U32638 ( .A(n32144), .B(n32143), .Z(n32145) );
  AND U32639 ( .A(n32146), .B(n32145), .Z(n32233) );
  NANDN U32640 ( .A(n32148), .B(n32147), .Z(n32152) );
  OR U32641 ( .A(n32150), .B(n32149), .Z(n32151) );
  NAND U32642 ( .A(n32152), .B(n32151), .Z(n32234) );
  XNOR U32643 ( .A(n32233), .B(n32234), .Z(n32235) );
  XOR U32644 ( .A(n32236), .B(n32235), .Z(n32264) );
  NANDN U32645 ( .A(n32154), .B(n32153), .Z(n32158) );
  NAND U32646 ( .A(n32156), .B(n32155), .Z(n32157) );
  AND U32647 ( .A(n32158), .B(n32157), .Z(n32263) );
  XNOR U32648 ( .A(n32264), .B(n32263), .Z(n32265) );
  NANDN U32649 ( .A(n32160), .B(n32159), .Z(n32164) );
  NAND U32650 ( .A(n32162), .B(n32161), .Z(n32163) );
  NAND U32651 ( .A(n32164), .B(n32163), .Z(n32266) );
  XNOR U32652 ( .A(n32265), .B(n32266), .Z(n32221) );
  XNOR U32653 ( .A(n32222), .B(n32221), .Z(n32223) );
  XOR U32654 ( .A(n32224), .B(n32223), .Z(n32417) );
  XNOR U32655 ( .A(n32416), .B(n32417), .Z(n32209) );
  XOR U32656 ( .A(n32210), .B(n32209), .Z(n32212) );
  XOR U32657 ( .A(n32211), .B(n32212), .Z(n32205) );
  NANDN U32658 ( .A(n32166), .B(n32165), .Z(n32170) );
  OR U32659 ( .A(n32168), .B(n32167), .Z(n32169) );
  AND U32660 ( .A(n32170), .B(n32169), .Z(n32203) );
  NANDN U32661 ( .A(n32172), .B(n32171), .Z(n32176) );
  NANDN U32662 ( .A(n32174), .B(n32173), .Z(n32175) );
  NAND U32663 ( .A(n32176), .B(n32175), .Z(n32204) );
  XOR U32664 ( .A(n32203), .B(n32204), .Z(n32206) );
  XOR U32665 ( .A(n32205), .B(n32206), .Z(n32198) );
  NANDN U32666 ( .A(n32178), .B(n32177), .Z(n32182) );
  NAND U32667 ( .A(n32180), .B(n32179), .Z(n32181) );
  NAND U32668 ( .A(n32182), .B(n32181), .Z(n32197) );
  XNOR U32669 ( .A(n32198), .B(n32197), .Z(n32200) );
  NANDN U32670 ( .A(n32184), .B(n32183), .Z(n32188) );
  NANDN U32671 ( .A(n32186), .B(n32185), .Z(n32187) );
  AND U32672 ( .A(n32188), .B(n32187), .Z(n32199) );
  XNOR U32673 ( .A(n32200), .B(n32199), .Z(n32191) );
  XOR U32674 ( .A(n32192), .B(n32191), .Z(n32194) );
  XNOR U32675 ( .A(n32193), .B(n32194), .Z(n32189) );
  XOR U32676 ( .A(n32190), .B(n32189), .Z(c[206]) );
  AND U32677 ( .A(n32190), .B(n32189), .Z(n32421) );
  NANDN U32678 ( .A(n32192), .B(n32191), .Z(n32196) );
  OR U32679 ( .A(n32194), .B(n32193), .Z(n32195) );
  AND U32680 ( .A(n32196), .B(n32195), .Z(n32424) );
  NANDN U32681 ( .A(n32198), .B(n32197), .Z(n32202) );
  NAND U32682 ( .A(n32200), .B(n32199), .Z(n32201) );
  AND U32683 ( .A(n32202), .B(n32201), .Z(n32422) );
  NANDN U32684 ( .A(n32204), .B(n32203), .Z(n32208) );
  OR U32685 ( .A(n32206), .B(n32205), .Z(n32207) );
  AND U32686 ( .A(n32208), .B(n32207), .Z(n32431) );
  NANDN U32687 ( .A(n32210), .B(n32209), .Z(n32214) );
  OR U32688 ( .A(n32212), .B(n32211), .Z(n32213) );
  AND U32689 ( .A(n32214), .B(n32213), .Z(n32428) );
  NANDN U32690 ( .A(n32216), .B(n32215), .Z(n32220) );
  OR U32691 ( .A(n32218), .B(n32217), .Z(n32219) );
  AND U32692 ( .A(n32220), .B(n32219), .Z(n32650) );
  NANDN U32693 ( .A(n32222), .B(n32221), .Z(n32226) );
  NANDN U32694 ( .A(n32224), .B(n32223), .Z(n32225) );
  AND U32695 ( .A(n32226), .B(n32225), .Z(n32648) );
  NANDN U32696 ( .A(n32228), .B(n32227), .Z(n32232) );
  NAND U32697 ( .A(n32230), .B(n32229), .Z(n32231) );
  AND U32698 ( .A(n32232), .B(n32231), .Z(n32448) );
  NANDN U32699 ( .A(n32234), .B(n32233), .Z(n32238) );
  NAND U32700 ( .A(n32236), .B(n32235), .Z(n32237) );
  AND U32701 ( .A(n32238), .B(n32237), .Z(n32446) );
  NANDN U32702 ( .A(n32240), .B(n32239), .Z(n32244) );
  NANDN U32703 ( .A(n32242), .B(n32241), .Z(n32243) );
  AND U32704 ( .A(n32244), .B(n32243), .Z(n32602) );
  NANDN U32705 ( .A(n32246), .B(n32245), .Z(n32250) );
  NANDN U32706 ( .A(n32248), .B(n32247), .Z(n32249) );
  AND U32707 ( .A(n32250), .B(n32249), .Z(n32599) );
  NANDN U32708 ( .A(n32252), .B(n32251), .Z(n32256) );
  NANDN U32709 ( .A(n32254), .B(n32253), .Z(n32255) );
  NAND U32710 ( .A(n32256), .B(n32255), .Z(n32600) );
  XNOR U32711 ( .A(n32599), .B(n32600), .Z(n32601) );
  XOR U32712 ( .A(n32602), .B(n32601), .Z(n32447) );
  XOR U32713 ( .A(n32446), .B(n32447), .Z(n32449) );
  XNOR U32714 ( .A(n32448), .B(n32449), .Z(n32647) );
  XNOR U32715 ( .A(n32648), .B(n32647), .Z(n32649) );
  XOR U32716 ( .A(n32650), .B(n32649), .Z(n32644) );
  NANDN U32717 ( .A(n32258), .B(n32257), .Z(n32262) );
  OR U32718 ( .A(n32260), .B(n32259), .Z(n32261) );
  AND U32719 ( .A(n32262), .B(n32261), .Z(n32436) );
  NANDN U32720 ( .A(n32264), .B(n32263), .Z(n32268) );
  NANDN U32721 ( .A(n32266), .B(n32265), .Z(n32267) );
  AND U32722 ( .A(n32268), .B(n32267), .Z(n32435) );
  NANDN U32723 ( .A(n32270), .B(n32269), .Z(n32274) );
  NAND U32724 ( .A(n32272), .B(n32271), .Z(n32273) );
  NAND U32725 ( .A(n32274), .B(n32273), .Z(n32442) );
  NANDN U32726 ( .A(n32276), .B(n32275), .Z(n32280) );
  OR U32727 ( .A(n32278), .B(n32277), .Z(n32279) );
  AND U32728 ( .A(n32280), .B(n32279), .Z(n32618) );
  IV U32729 ( .A(n32299), .Z(n32537) );
  NANDN U32730 ( .A(n32537), .B(n32281), .Z(n32285) );
  NANDN U32731 ( .A(n32283), .B(n32282), .Z(n32284) );
  NAND U32732 ( .A(n32285), .B(n32284), .Z(n32617) );
  XNOR U32733 ( .A(n32618), .B(n32617), .Z(n32620) );
  NANDN U32734 ( .A(n32287), .B(n32286), .Z(n32291) );
  NANDN U32735 ( .A(n32289), .B(n32288), .Z(n32290) );
  AND U32736 ( .A(n32291), .B(n32290), .Z(n32632) );
  XNOR U32737 ( .A(a[127]), .B(b[17]), .Z(n32543) );
  OR U32738 ( .A(n32543), .B(n32292), .Z(n32295) );
  NAND U32739 ( .A(n32544), .B(n32293), .Z(n32294) );
  AND U32740 ( .A(n32295), .B(n32294), .Z(n32558) );
  NANDN U32741 ( .A(n36480), .B(n32296), .Z(n32298) );
  XOR U32742 ( .A(b[41]), .B(a[103]), .Z(n32554) );
  NANDN U32743 ( .A(n36594), .B(n32554), .Z(n32297) );
  NAND U32744 ( .A(n32298), .B(n32297), .Z(n32557) );
  XNOR U32745 ( .A(n32558), .B(n32557), .Z(n32559) );
  AND U32746 ( .A(b[63]), .B(a[79]), .Z(n32534) );
  XOR U32747 ( .A(n32535), .B(n32534), .Z(n32536) );
  XOR U32748 ( .A(n32299), .B(n32536), .Z(n32560) );
  XOR U32749 ( .A(n32559), .B(n32560), .Z(n32629) );
  NANDN U32750 ( .A(n212), .B(n32300), .Z(n32302) );
  XOR U32751 ( .A(b[49]), .B(a[95]), .Z(n32572) );
  NANDN U32752 ( .A(n37432), .B(n32572), .Z(n32301) );
  AND U32753 ( .A(n32302), .B(n32301), .Z(n32590) );
  NANDN U32754 ( .A(n37526), .B(n32303), .Z(n32305) );
  XOR U32755 ( .A(b[51]), .B(a[93]), .Z(n32581) );
  NANDN U32756 ( .A(n37605), .B(n32581), .Z(n32304) );
  AND U32757 ( .A(n32305), .B(n32304), .Z(n32588) );
  NANDN U32758 ( .A(n33875), .B(n32306), .Z(n32308) );
  XOR U32759 ( .A(a[119]), .B(b[25]), .Z(n32464) );
  NANDN U32760 ( .A(n33994), .B(n32464), .Z(n32307) );
  NAND U32761 ( .A(n32308), .B(n32307), .Z(n32587) );
  XNOR U32762 ( .A(n32588), .B(n32587), .Z(n32589) );
  XOR U32763 ( .A(n32590), .B(n32589), .Z(n32630) );
  XNOR U32764 ( .A(n32629), .B(n32630), .Z(n32631) );
  XNOR U32765 ( .A(n32632), .B(n32631), .Z(n32619) );
  XOR U32766 ( .A(n32620), .B(n32619), .Z(n32455) );
  NANDN U32767 ( .A(n32310), .B(n32309), .Z(n32314) );
  NAND U32768 ( .A(n32312), .B(n32311), .Z(n32313) );
  AND U32769 ( .A(n32314), .B(n32313), .Z(n32453) );
  NANDN U32770 ( .A(n35936), .B(n32315), .Z(n32317) );
  XOR U32771 ( .A(a[107]), .B(b[37]), .Z(n32584) );
  NANDN U32772 ( .A(n36047), .B(n32584), .Z(n32316) );
  AND U32773 ( .A(n32317), .B(n32316), .Z(n32565) );
  NANDN U32774 ( .A(n36210), .B(n32318), .Z(n32320) );
  XOR U32775 ( .A(b[39]), .B(a[105]), .Z(n32461) );
  NANDN U32776 ( .A(n36347), .B(n32461), .Z(n32319) );
  AND U32777 ( .A(n32320), .B(n32319), .Z(n32564) );
  NANDN U32778 ( .A(n34223), .B(n32321), .Z(n32323) );
  XOR U32779 ( .A(a[117]), .B(b[27]), .Z(n32473) );
  NANDN U32780 ( .A(n34458), .B(n32473), .Z(n32322) );
  NAND U32781 ( .A(n32323), .B(n32322), .Z(n32563) );
  XOR U32782 ( .A(n32564), .B(n32563), .Z(n32566) );
  XOR U32783 ( .A(n32565), .B(n32566), .Z(n32596) );
  NANDN U32784 ( .A(n34909), .B(n32324), .Z(n32326) );
  XOR U32785 ( .A(a[113]), .B(b[31]), .Z(n32476) );
  NANDN U32786 ( .A(n35145), .B(n32476), .Z(n32325) );
  AND U32787 ( .A(n32326), .B(n32325), .Z(n32530) );
  NANDN U32788 ( .A(n35611), .B(n32327), .Z(n32329) );
  XOR U32789 ( .A(a[109]), .B(b[35]), .Z(n32458) );
  NANDN U32790 ( .A(n35801), .B(n32458), .Z(n32328) );
  AND U32791 ( .A(n32329), .B(n32328), .Z(n32529) );
  NANDN U32792 ( .A(n35260), .B(n32330), .Z(n32332) );
  XOR U32793 ( .A(a[111]), .B(b[33]), .Z(n32467) );
  NANDN U32794 ( .A(n35456), .B(n32467), .Z(n32331) );
  NAND U32795 ( .A(n32332), .B(n32331), .Z(n32528) );
  XOR U32796 ( .A(n32529), .B(n32528), .Z(n32531) );
  XOR U32797 ( .A(n32530), .B(n32531), .Z(n32594) );
  NANDN U32798 ( .A(n32333), .B(n35001), .Z(n32335) );
  XNOR U32799 ( .A(a[115]), .B(b[29]), .Z(n32470) );
  NANDN U32800 ( .A(n32470), .B(n35002), .Z(n32334) );
  AND U32801 ( .A(n32335), .B(n32334), .Z(n32593) );
  XNOR U32802 ( .A(n32594), .B(n32593), .Z(n32595) );
  XNOR U32803 ( .A(n32596), .B(n32595), .Z(n32452) );
  XNOR U32804 ( .A(n32453), .B(n32452), .Z(n32454) );
  XOR U32805 ( .A(n32455), .B(n32454), .Z(n32441) );
  NANDN U32806 ( .A(n32996), .B(n32336), .Z(n32338) );
  XOR U32807 ( .A(a[123]), .B(b[21]), .Z(n32578) );
  NANDN U32808 ( .A(n33271), .B(n32578), .Z(n32337) );
  AND U32809 ( .A(n32338), .B(n32337), .Z(n32506) );
  NANDN U32810 ( .A(n38247), .B(n32339), .Z(n32341) );
  XOR U32811 ( .A(b[61]), .B(a[83]), .Z(n32479) );
  NANDN U32812 ( .A(n38248), .B(n32479), .Z(n32340) );
  AND U32813 ( .A(n32341), .B(n32340), .Z(n32505) );
  NANDN U32814 ( .A(n36991), .B(n32342), .Z(n32344) );
  XOR U32815 ( .A(b[45]), .B(a[99]), .Z(n32495) );
  NANDN U32816 ( .A(n37083), .B(n32495), .Z(n32343) );
  NAND U32817 ( .A(n32344), .B(n32343), .Z(n32504) );
  XOR U32818 ( .A(n32505), .B(n32504), .Z(n32507) );
  XOR U32819 ( .A(n32506), .B(n32507), .Z(n32636) );
  NANDN U32820 ( .A(n37974), .B(n32345), .Z(n32347) );
  XOR U32821 ( .A(b[57]), .B(a[87]), .Z(n32489) );
  NANDN U32822 ( .A(n38031), .B(n32489), .Z(n32346) );
  AND U32823 ( .A(n32347), .B(n32346), .Z(n32518) );
  NANDN U32824 ( .A(n38090), .B(n32348), .Z(n32350) );
  XOR U32825 ( .A(b[59]), .B(a[85]), .Z(n32492) );
  NANDN U32826 ( .A(n38130), .B(n32492), .Z(n32349) );
  AND U32827 ( .A(n32350), .B(n32349), .Z(n32517) );
  NANDN U32828 ( .A(n211), .B(n32351), .Z(n32353) );
  XOR U32829 ( .A(b[47]), .B(a[97]), .Z(n32569) );
  NANDN U32830 ( .A(n37172), .B(n32569), .Z(n32352) );
  NAND U32831 ( .A(n32353), .B(n32352), .Z(n32516) );
  XOR U32832 ( .A(n32517), .B(n32516), .Z(n32519) );
  XNOR U32833 ( .A(n32518), .B(n32519), .Z(n32635) );
  XNOR U32834 ( .A(n32636), .B(n32635), .Z(n32637) );
  NANDN U32835 ( .A(n32355), .B(n32354), .Z(n32359) );
  OR U32836 ( .A(n32357), .B(n32356), .Z(n32358) );
  NAND U32837 ( .A(n32359), .B(n32358), .Z(n32638) );
  XNOR U32838 ( .A(n32637), .B(n32638), .Z(n32611) );
  NANDN U32839 ( .A(n32361), .B(n32360), .Z(n32365) );
  OR U32840 ( .A(n32363), .B(n32362), .Z(n32364) );
  NAND U32841 ( .A(n32365), .B(n32364), .Z(n32612) );
  XNOR U32842 ( .A(n32611), .B(n32612), .Z(n32613) );
  NANDN U32843 ( .A(n32367), .B(n32366), .Z(n32371) );
  OR U32844 ( .A(n32369), .B(n32368), .Z(n32370) );
  NAND U32845 ( .A(n32371), .B(n32370), .Z(n32614) );
  XNOR U32846 ( .A(n32613), .B(n32614), .Z(n32608) );
  NANDN U32847 ( .A(n32483), .B(n32372), .Z(n32374) );
  XOR U32848 ( .A(a[125]), .B(b[19]), .Z(n32482) );
  NANDN U32849 ( .A(n32823), .B(n32482), .Z(n32373) );
  AND U32850 ( .A(n32374), .B(n32373), .Z(n32524) );
  NANDN U32851 ( .A(n38278), .B(n32375), .Z(n32377) );
  XOR U32852 ( .A(b[63]), .B(a[81]), .Z(n32540) );
  NANDN U32853 ( .A(n38279), .B(n32540), .Z(n32376) );
  AND U32854 ( .A(n32377), .B(n32376), .Z(n32523) );
  NANDN U32855 ( .A(n36742), .B(n32378), .Z(n32380) );
  XOR U32856 ( .A(b[43]), .B(a[101]), .Z(n32486) );
  NANDN U32857 ( .A(n36891), .B(n32486), .Z(n32379) );
  NAND U32858 ( .A(n32380), .B(n32379), .Z(n32522) );
  XOR U32859 ( .A(n32523), .B(n32522), .Z(n32525) );
  XOR U32860 ( .A(n32524), .B(n32525), .Z(n32511) );
  NANDN U32861 ( .A(n33866), .B(n32381), .Z(n32383) );
  XOR U32862 ( .A(a[121]), .B(b[23]), .Z(n32575) );
  NANDN U32863 ( .A(n33644), .B(n32575), .Z(n32382) );
  AND U32864 ( .A(n32383), .B(n32382), .Z(n32500) );
  NANDN U32865 ( .A(n37857), .B(n32384), .Z(n32386) );
  XOR U32866 ( .A(b[55]), .B(a[89]), .Z(n32551) );
  NANDN U32867 ( .A(n37911), .B(n32551), .Z(n32385) );
  AND U32868 ( .A(n32386), .B(n32385), .Z(n32499) );
  NANDN U32869 ( .A(n37705), .B(n32387), .Z(n32389) );
  XOR U32870 ( .A(b[53]), .B(a[91]), .Z(n32548) );
  NANDN U32871 ( .A(n37778), .B(n32548), .Z(n32388) );
  NAND U32872 ( .A(n32389), .B(n32388), .Z(n32498) );
  XOR U32873 ( .A(n32499), .B(n32498), .Z(n32501) );
  XNOR U32874 ( .A(n32500), .B(n32501), .Z(n32510) );
  XNOR U32875 ( .A(n32511), .B(n32510), .Z(n32513) );
  NANDN U32876 ( .A(n32391), .B(n32390), .Z(n32395) );
  OR U32877 ( .A(n32393), .B(n32392), .Z(n32394) );
  AND U32878 ( .A(n32395), .B(n32394), .Z(n32512) );
  XOR U32879 ( .A(n32513), .B(n32512), .Z(n32625) );
  NANDN U32880 ( .A(n32397), .B(n32396), .Z(n32401) );
  OR U32881 ( .A(n32399), .B(n32398), .Z(n32400) );
  AND U32882 ( .A(n32401), .B(n32400), .Z(n32624) );
  NANDN U32883 ( .A(n32403), .B(n32402), .Z(n32407) );
  OR U32884 ( .A(n32405), .B(n32404), .Z(n32406) );
  NAND U32885 ( .A(n32407), .B(n32406), .Z(n32623) );
  XOR U32886 ( .A(n32624), .B(n32623), .Z(n32626) );
  XOR U32887 ( .A(n32625), .B(n32626), .Z(n32606) );
  NANDN U32888 ( .A(n32409), .B(n32408), .Z(n32413) );
  NAND U32889 ( .A(n32411), .B(n32410), .Z(n32412) );
  NAND U32890 ( .A(n32413), .B(n32412), .Z(n32605) );
  XNOR U32891 ( .A(n32606), .B(n32605), .Z(n32607) );
  XNOR U32892 ( .A(n32608), .B(n32607), .Z(n32440) );
  XOR U32893 ( .A(n32441), .B(n32440), .Z(n32443) );
  XOR U32894 ( .A(n32442), .B(n32443), .Z(n32434) );
  XOR U32895 ( .A(n32435), .B(n32434), .Z(n32437) );
  XOR U32896 ( .A(n32436), .B(n32437), .Z(n32642) );
  NANDN U32897 ( .A(n32415), .B(n32414), .Z(n32419) );
  NANDN U32898 ( .A(n32417), .B(n32416), .Z(n32418) );
  AND U32899 ( .A(n32419), .B(n32418), .Z(n32641) );
  XNOR U32900 ( .A(n32642), .B(n32641), .Z(n32643) );
  XOR U32901 ( .A(n32644), .B(n32643), .Z(n32429) );
  XNOR U32902 ( .A(n32428), .B(n32429), .Z(n32430) );
  XOR U32903 ( .A(n32431), .B(n32430), .Z(n32423) );
  XOR U32904 ( .A(n32422), .B(n32423), .Z(n32425) );
  XNOR U32905 ( .A(n32424), .B(n32425), .Z(n32420) );
  XOR U32906 ( .A(n32421), .B(n32420), .Z(c[207]) );
  AND U32907 ( .A(n32421), .B(n32420), .Z(n32654) );
  NANDN U32908 ( .A(n32423), .B(n32422), .Z(n32427) );
  OR U32909 ( .A(n32425), .B(n32424), .Z(n32426) );
  AND U32910 ( .A(n32427), .B(n32426), .Z(n32657) );
  NANDN U32911 ( .A(n32429), .B(n32428), .Z(n32433) );
  NANDN U32912 ( .A(n32431), .B(n32430), .Z(n32432) );
  AND U32913 ( .A(n32433), .B(n32432), .Z(n32656) );
  NANDN U32914 ( .A(n32435), .B(n32434), .Z(n32439) );
  OR U32915 ( .A(n32437), .B(n32436), .Z(n32438) );
  AND U32916 ( .A(n32439), .B(n32438), .Z(n32871) );
  NAND U32917 ( .A(n32441), .B(n32440), .Z(n32445) );
  NAND U32918 ( .A(n32443), .B(n32442), .Z(n32444) );
  NAND U32919 ( .A(n32445), .B(n32444), .Z(n32870) );
  XNOR U32920 ( .A(n32871), .B(n32870), .Z(n32873) );
  NANDN U32921 ( .A(n32447), .B(n32446), .Z(n32451) );
  NANDN U32922 ( .A(n32449), .B(n32448), .Z(n32450) );
  AND U32923 ( .A(n32451), .B(n32450), .Z(n32668) );
  NANDN U32924 ( .A(n32453), .B(n32452), .Z(n32457) );
  NANDN U32925 ( .A(n32455), .B(n32454), .Z(n32456) );
  AND U32926 ( .A(n32457), .B(n32456), .Z(n32675) );
  NANDN U32927 ( .A(n35611), .B(n32458), .Z(n32460) );
  XOR U32928 ( .A(a[110]), .B(b[35]), .Z(n32715) );
  NANDN U32929 ( .A(n35801), .B(n32715), .Z(n32459) );
  AND U32930 ( .A(n32460), .B(n32459), .Z(n32819) );
  NANDN U32931 ( .A(n36210), .B(n32461), .Z(n32463) );
  XOR U32932 ( .A(a[106]), .B(b[39]), .Z(n32831) );
  NANDN U32933 ( .A(n36347), .B(n32831), .Z(n32462) );
  AND U32934 ( .A(n32463), .B(n32462), .Z(n32818) );
  NANDN U32935 ( .A(n33875), .B(n32464), .Z(n32466) );
  XOR U32936 ( .A(a[120]), .B(b[25]), .Z(n32769) );
  NANDN U32937 ( .A(n33994), .B(n32769), .Z(n32465) );
  NAND U32938 ( .A(n32466), .B(n32465), .Z(n32817) );
  XOR U32939 ( .A(n32818), .B(n32817), .Z(n32820) );
  XOR U32940 ( .A(n32819), .B(n32820), .Z(n32861) );
  NANDN U32941 ( .A(n35260), .B(n32467), .Z(n32469) );
  XOR U32942 ( .A(a[112]), .B(b[33]), .Z(n32808) );
  NANDN U32943 ( .A(n35456), .B(n32808), .Z(n32468) );
  AND U32944 ( .A(n32469), .B(n32468), .Z(n32789) );
  NANDN U32945 ( .A(n32470), .B(n35001), .Z(n32472) );
  XOR U32946 ( .A(a[116]), .B(b[29]), .Z(n32781) );
  NANDN U32947 ( .A(n34722), .B(n32781), .Z(n32471) );
  AND U32948 ( .A(n32472), .B(n32471), .Z(n32788) );
  NANDN U32949 ( .A(n34223), .B(n32473), .Z(n32475) );
  XOR U32950 ( .A(a[118]), .B(b[27]), .Z(n32718) );
  NANDN U32951 ( .A(n34458), .B(n32718), .Z(n32474) );
  NAND U32952 ( .A(n32475), .B(n32474), .Z(n32787) );
  XOR U32953 ( .A(n32788), .B(n32787), .Z(n32790) );
  XOR U32954 ( .A(n32789), .B(n32790), .Z(n32859) );
  NAND U32955 ( .A(n35309), .B(n32476), .Z(n32478) );
  XNOR U32956 ( .A(a[114]), .B(b[31]), .Z(n32778) );
  NANDN U32957 ( .A(n32778), .B(n35310), .Z(n32477) );
  AND U32958 ( .A(n32478), .B(n32477), .Z(n32858) );
  XNOR U32959 ( .A(n32859), .B(n32858), .Z(n32860) );
  XNOR U32960 ( .A(n32861), .B(n32860), .Z(n32766) );
  NANDN U32961 ( .A(n38247), .B(n32479), .Z(n32481) );
  XOR U32962 ( .A(b[61]), .B(a[84]), .Z(n32721) );
  NANDN U32963 ( .A(n38248), .B(n32721), .Z(n32480) );
  AND U32964 ( .A(n32481), .B(n32480), .Z(n32705) );
  NANDN U32965 ( .A(n32483), .B(n32482), .Z(n32485) );
  XOR U32966 ( .A(a[126]), .B(b[19]), .Z(n32824) );
  NANDN U32967 ( .A(n32823), .B(n32824), .Z(n32484) );
  AND U32968 ( .A(n32485), .B(n32484), .Z(n32704) );
  NANDN U32969 ( .A(n36742), .B(n32486), .Z(n32488) );
  XOR U32970 ( .A(b[43]), .B(a[102]), .Z(n32827) );
  NANDN U32971 ( .A(n36891), .B(n32827), .Z(n32487) );
  NAND U32972 ( .A(n32488), .B(n32487), .Z(n32703) );
  XOR U32973 ( .A(n32704), .B(n32703), .Z(n32706) );
  XOR U32974 ( .A(n32705), .B(n32706), .Z(n32686) );
  NANDN U32975 ( .A(n37974), .B(n32489), .Z(n32491) );
  XOR U32976 ( .A(b[57]), .B(a[88]), .Z(n32784) );
  NANDN U32977 ( .A(n38031), .B(n32784), .Z(n32490) );
  AND U32978 ( .A(n32491), .B(n32490), .Z(n32735) );
  NANDN U32979 ( .A(n38090), .B(n32492), .Z(n32494) );
  XOR U32980 ( .A(b[59]), .B(a[86]), .Z(n32805) );
  NANDN U32981 ( .A(n38130), .B(n32805), .Z(n32493) );
  AND U32982 ( .A(n32494), .B(n32493), .Z(n32734) );
  NANDN U32983 ( .A(n36991), .B(n32495), .Z(n32497) );
  XOR U32984 ( .A(b[45]), .B(a[100]), .Z(n32799) );
  NANDN U32985 ( .A(n37083), .B(n32799), .Z(n32496) );
  NAND U32986 ( .A(n32497), .B(n32496), .Z(n32733) );
  XOR U32987 ( .A(n32734), .B(n32733), .Z(n32736) );
  XNOR U32988 ( .A(n32735), .B(n32736), .Z(n32685) );
  XNOR U32989 ( .A(n32686), .B(n32685), .Z(n32687) );
  NANDN U32990 ( .A(n32499), .B(n32498), .Z(n32503) );
  OR U32991 ( .A(n32501), .B(n32500), .Z(n32502) );
  NAND U32992 ( .A(n32503), .B(n32502), .Z(n32688) );
  XNOR U32993 ( .A(n32687), .B(n32688), .Z(n32764) );
  NANDN U32994 ( .A(n32505), .B(n32504), .Z(n32509) );
  OR U32995 ( .A(n32507), .B(n32506), .Z(n32508) );
  AND U32996 ( .A(n32509), .B(n32508), .Z(n32763) );
  XOR U32997 ( .A(n32764), .B(n32763), .Z(n32765) );
  XOR U32998 ( .A(n32766), .B(n32765), .Z(n32747) );
  NANDN U32999 ( .A(n32511), .B(n32510), .Z(n32515) );
  NAND U33000 ( .A(n32513), .B(n32512), .Z(n32514) );
  AND U33001 ( .A(n32515), .B(n32514), .Z(n32745) );
  NANDN U33002 ( .A(n32517), .B(n32516), .Z(n32521) );
  OR U33003 ( .A(n32519), .B(n32518), .Z(n32520) );
  AND U33004 ( .A(n32521), .B(n32520), .Z(n32698) );
  NANDN U33005 ( .A(n32523), .B(n32522), .Z(n32527) );
  OR U33006 ( .A(n32525), .B(n32524), .Z(n32526) );
  NAND U33007 ( .A(n32527), .B(n32526), .Z(n32697) );
  XNOR U33008 ( .A(n32698), .B(n32697), .Z(n32699) );
  NANDN U33009 ( .A(n32529), .B(n32528), .Z(n32533) );
  OR U33010 ( .A(n32531), .B(n32530), .Z(n32532) );
  AND U33011 ( .A(n32533), .B(n32532), .Z(n32855) );
  NANDN U33012 ( .A(n32535), .B(n32534), .Z(n32539) );
  ANDN U33013 ( .B(n32537), .A(n32536), .Z(n32538) );
  ANDN U33014 ( .B(n32539), .A(n32538), .Z(n32853) );
  NANDN U33015 ( .A(n38278), .B(n32540), .Z(n32542) );
  XOR U33016 ( .A(b[63]), .B(a[82]), .Z(n32796) );
  NANDN U33017 ( .A(n38279), .B(n32796), .Z(n32541) );
  AND U33018 ( .A(n32542), .B(n32541), .Z(n32849) );
  NAND U33019 ( .A(b[63]), .B(a[80]), .Z(n32846) );
  ANDN U33020 ( .B(n32544), .A(n32543), .Z(n32547) );
  NAND U33021 ( .A(b[17]), .B(n32545), .Z(n32546) );
  NANDN U33022 ( .A(n32547), .B(n32546), .Z(n32847) );
  XOR U33023 ( .A(n32846), .B(n32847), .Z(n32848) );
  XNOR U33024 ( .A(n32849), .B(n32848), .Z(n32852) );
  XNOR U33025 ( .A(n32853), .B(n32852), .Z(n32854) );
  XOR U33026 ( .A(n32855), .B(n32854), .Z(n32700) );
  XOR U33027 ( .A(n32699), .B(n32700), .Z(n32746) );
  XOR U33028 ( .A(n32745), .B(n32746), .Z(n32748) );
  XOR U33029 ( .A(n32747), .B(n32748), .Z(n32674) );
  NANDN U33030 ( .A(n37705), .B(n32548), .Z(n32550) );
  XOR U33031 ( .A(b[53]), .B(a[92]), .Z(n32712) );
  NANDN U33032 ( .A(n37778), .B(n32712), .Z(n32549) );
  AND U33033 ( .A(n32550), .B(n32549), .Z(n32842) );
  NANDN U33034 ( .A(n37857), .B(n32551), .Z(n32553) );
  XOR U33035 ( .A(b[55]), .B(a[90]), .Z(n32802) );
  NANDN U33036 ( .A(n37911), .B(n32802), .Z(n32552) );
  AND U33037 ( .A(n32553), .B(n32552), .Z(n32841) );
  NANDN U33038 ( .A(n36480), .B(n32554), .Z(n32556) );
  XOR U33039 ( .A(b[41]), .B(a[104]), .Z(n32834) );
  NANDN U33040 ( .A(n36594), .B(n32834), .Z(n32555) );
  NAND U33041 ( .A(n32556), .B(n32555), .Z(n32840) );
  XOR U33042 ( .A(n32841), .B(n32840), .Z(n32843) );
  XOR U33043 ( .A(n32842), .B(n32843), .Z(n32692) );
  NANDN U33044 ( .A(n32558), .B(n32557), .Z(n32562) );
  NAND U33045 ( .A(n32560), .B(n32559), .Z(n32561) );
  AND U33046 ( .A(n32562), .B(n32561), .Z(n32691) );
  XNOR U33047 ( .A(n32692), .B(n32691), .Z(n32694) );
  NANDN U33048 ( .A(n32564), .B(n32563), .Z(n32568) );
  OR U33049 ( .A(n32566), .B(n32565), .Z(n32567) );
  AND U33050 ( .A(n32568), .B(n32567), .Z(n32693) );
  XOR U33051 ( .A(n32694), .B(n32693), .Z(n32759) );
  NANDN U33052 ( .A(n211), .B(n32569), .Z(n32571) );
  XOR U33053 ( .A(b[47]), .B(a[98]), .Z(n32775) );
  NANDN U33054 ( .A(n37172), .B(n32775), .Z(n32570) );
  AND U33055 ( .A(n32571), .B(n32570), .Z(n32729) );
  NANDN U33056 ( .A(n212), .B(n32572), .Z(n32574) );
  XOR U33057 ( .A(b[49]), .B(a[96]), .Z(n32709) );
  NANDN U33058 ( .A(n37432), .B(n32709), .Z(n32573) );
  AND U33059 ( .A(n32574), .B(n32573), .Z(n32728) );
  NANDN U33060 ( .A(n33866), .B(n32575), .Z(n32577) );
  XOR U33061 ( .A(a[122]), .B(b[23]), .Z(n32772) );
  NANDN U33062 ( .A(n33644), .B(n32772), .Z(n32576) );
  NAND U33063 ( .A(n32577), .B(n32576), .Z(n32727) );
  XOR U33064 ( .A(n32728), .B(n32727), .Z(n32730) );
  XOR U33065 ( .A(n32729), .B(n32730), .Z(n32740) );
  NANDN U33066 ( .A(n32996), .B(n32578), .Z(n32580) );
  XOR U33067 ( .A(a[124]), .B(b[21]), .Z(n32793) );
  NANDN U33068 ( .A(n33271), .B(n32793), .Z(n32579) );
  AND U33069 ( .A(n32580), .B(n32579), .Z(n32813) );
  NANDN U33070 ( .A(n37526), .B(n32581), .Z(n32583) );
  XOR U33071 ( .A(b[51]), .B(a[94]), .Z(n32724) );
  NANDN U33072 ( .A(n37605), .B(n32724), .Z(n32582) );
  AND U33073 ( .A(n32583), .B(n32582), .Z(n32812) );
  NANDN U33074 ( .A(n35936), .B(n32584), .Z(n32586) );
  XOR U33075 ( .A(a[108]), .B(b[37]), .Z(n32837) );
  NANDN U33076 ( .A(n36047), .B(n32837), .Z(n32585) );
  NAND U33077 ( .A(n32586), .B(n32585), .Z(n32811) );
  XOR U33078 ( .A(n32812), .B(n32811), .Z(n32814) );
  XNOR U33079 ( .A(n32813), .B(n32814), .Z(n32739) );
  XNOR U33080 ( .A(n32740), .B(n32739), .Z(n32742) );
  NANDN U33081 ( .A(n32588), .B(n32587), .Z(n32592) );
  NANDN U33082 ( .A(n32590), .B(n32589), .Z(n32591) );
  AND U33083 ( .A(n32592), .B(n32591), .Z(n32741) );
  XOR U33084 ( .A(n32742), .B(n32741), .Z(n32758) );
  NANDN U33085 ( .A(n32594), .B(n32593), .Z(n32598) );
  NANDN U33086 ( .A(n32596), .B(n32595), .Z(n32597) );
  AND U33087 ( .A(n32598), .B(n32597), .Z(n32757) );
  XOR U33088 ( .A(n32758), .B(n32757), .Z(n32760) );
  XNOR U33089 ( .A(n32759), .B(n32760), .Z(n32673) );
  XOR U33090 ( .A(n32674), .B(n32673), .Z(n32676) );
  XNOR U33091 ( .A(n32675), .B(n32676), .Z(n32667) );
  XNOR U33092 ( .A(n32668), .B(n32667), .Z(n32669) );
  NANDN U33093 ( .A(n32600), .B(n32599), .Z(n32604) );
  NANDN U33094 ( .A(n32602), .B(n32601), .Z(n32603) );
  AND U33095 ( .A(n32604), .B(n32603), .Z(n32865) );
  NANDN U33096 ( .A(n32606), .B(n32605), .Z(n32610) );
  NAND U33097 ( .A(n32608), .B(n32607), .Z(n32609) );
  AND U33098 ( .A(n32610), .B(n32609), .Z(n32864) );
  XNOR U33099 ( .A(n32865), .B(n32864), .Z(n32866) );
  NANDN U33100 ( .A(n32612), .B(n32611), .Z(n32616) );
  NANDN U33101 ( .A(n32614), .B(n32613), .Z(n32615) );
  AND U33102 ( .A(n32616), .B(n32615), .Z(n32681) );
  NANDN U33103 ( .A(n32618), .B(n32617), .Z(n32622) );
  NAND U33104 ( .A(n32620), .B(n32619), .Z(n32621) );
  AND U33105 ( .A(n32622), .B(n32621), .Z(n32680) );
  NANDN U33106 ( .A(n32624), .B(n32623), .Z(n32628) );
  OR U33107 ( .A(n32626), .B(n32625), .Z(n32627) );
  AND U33108 ( .A(n32628), .B(n32627), .Z(n32754) );
  NANDN U33109 ( .A(n32630), .B(n32629), .Z(n32634) );
  NANDN U33110 ( .A(n32632), .B(n32631), .Z(n32633) );
  AND U33111 ( .A(n32634), .B(n32633), .Z(n32752) );
  NANDN U33112 ( .A(n32636), .B(n32635), .Z(n32640) );
  NANDN U33113 ( .A(n32638), .B(n32637), .Z(n32639) );
  AND U33114 ( .A(n32640), .B(n32639), .Z(n32751) );
  XNOR U33115 ( .A(n32752), .B(n32751), .Z(n32753) );
  XNOR U33116 ( .A(n32754), .B(n32753), .Z(n32679) );
  XOR U33117 ( .A(n32680), .B(n32679), .Z(n32682) );
  XOR U33118 ( .A(n32681), .B(n32682), .Z(n32867) );
  XOR U33119 ( .A(n32866), .B(n32867), .Z(n32670) );
  XNOR U33120 ( .A(n32669), .B(n32670), .Z(n32872) );
  XOR U33121 ( .A(n32873), .B(n32872), .Z(n32664) );
  NANDN U33122 ( .A(n32642), .B(n32641), .Z(n32646) );
  NANDN U33123 ( .A(n32644), .B(n32643), .Z(n32645) );
  AND U33124 ( .A(n32646), .B(n32645), .Z(n32662) );
  NANDN U33125 ( .A(n32648), .B(n32647), .Z(n32652) );
  NAND U33126 ( .A(n32650), .B(n32649), .Z(n32651) );
  AND U33127 ( .A(n32652), .B(n32651), .Z(n32661) );
  XNOR U33128 ( .A(n32662), .B(n32661), .Z(n32663) );
  XNOR U33129 ( .A(n32664), .B(n32663), .Z(n32655) );
  XOR U33130 ( .A(n32656), .B(n32655), .Z(n32658) );
  XNOR U33131 ( .A(n32657), .B(n32658), .Z(n32653) );
  XOR U33132 ( .A(n32654), .B(n32653), .Z(c[208]) );
  AND U33133 ( .A(n32654), .B(n32653), .Z(n32877) );
  NANDN U33134 ( .A(n32656), .B(n32655), .Z(n32660) );
  OR U33135 ( .A(n32658), .B(n32657), .Z(n32659) );
  AND U33136 ( .A(n32660), .B(n32659), .Z(n32880) );
  NANDN U33137 ( .A(n32662), .B(n32661), .Z(n32666) );
  NANDN U33138 ( .A(n32664), .B(n32663), .Z(n32665) );
  AND U33139 ( .A(n32666), .B(n32665), .Z(n32879) );
  NANDN U33140 ( .A(n32668), .B(n32667), .Z(n32672) );
  NANDN U33141 ( .A(n32670), .B(n32669), .Z(n32671) );
  AND U33142 ( .A(n32672), .B(n32671), .Z(n32884) );
  NANDN U33143 ( .A(n32674), .B(n32673), .Z(n32678) );
  OR U33144 ( .A(n32676), .B(n32675), .Z(n32677) );
  AND U33145 ( .A(n32678), .B(n32677), .Z(n32899) );
  NANDN U33146 ( .A(n32680), .B(n32679), .Z(n32684) );
  NANDN U33147 ( .A(n32682), .B(n32681), .Z(n32683) );
  AND U33148 ( .A(n32684), .B(n32683), .Z(n32897) );
  NANDN U33149 ( .A(n32686), .B(n32685), .Z(n32690) );
  NANDN U33150 ( .A(n32688), .B(n32687), .Z(n32689) );
  AND U33151 ( .A(n32690), .B(n32689), .Z(n32962) );
  NANDN U33152 ( .A(n32692), .B(n32691), .Z(n32696) );
  NAND U33153 ( .A(n32694), .B(n32693), .Z(n32695) );
  NAND U33154 ( .A(n32696), .B(n32695), .Z(n32963) );
  XNOR U33155 ( .A(n32962), .B(n32963), .Z(n32964) );
  NANDN U33156 ( .A(n32698), .B(n32697), .Z(n32702) );
  NANDN U33157 ( .A(n32700), .B(n32699), .Z(n32701) );
  AND U33158 ( .A(n32702), .B(n32701), .Z(n32959) );
  NANDN U33159 ( .A(n32704), .B(n32703), .Z(n32708) );
  OR U33160 ( .A(n32706), .B(n32705), .Z(n32707) );
  AND U33161 ( .A(n32708), .B(n32707), .Z(n32983) );
  NANDN U33162 ( .A(n212), .B(n32709), .Z(n32711) );
  XOR U33163 ( .A(b[49]), .B(a[97]), .Z(n33037) );
  NANDN U33164 ( .A(n37432), .B(n33037), .Z(n32710) );
  AND U33165 ( .A(n32711), .B(n32710), .Z(n33006) );
  NANDN U33166 ( .A(n37705), .B(n32712), .Z(n32714) );
  XOR U33167 ( .A(b[53]), .B(a[93]), .Z(n33025) );
  NANDN U33168 ( .A(n37778), .B(n33025), .Z(n32713) );
  AND U33169 ( .A(n32714), .B(n32713), .Z(n33005) );
  NANDN U33170 ( .A(n35611), .B(n32715), .Z(n32717) );
  XOR U33171 ( .A(a[111]), .B(b[35]), .Z(n33028) );
  NANDN U33172 ( .A(n35801), .B(n33028), .Z(n32716) );
  NAND U33173 ( .A(n32717), .B(n32716), .Z(n33004) );
  XOR U33174 ( .A(n33005), .B(n33004), .Z(n33007) );
  XOR U33175 ( .A(n33006), .B(n33007), .Z(n33077) );
  NANDN U33176 ( .A(n34223), .B(n32718), .Z(n32720) );
  XOR U33177 ( .A(a[119]), .B(b[27]), .Z(n33034) );
  NANDN U33178 ( .A(n34458), .B(n33034), .Z(n32719) );
  AND U33179 ( .A(n32720), .B(n32719), .Z(n32946) );
  NANDN U33180 ( .A(n38247), .B(n32721), .Z(n32723) );
  XOR U33181 ( .A(b[61]), .B(a[85]), .Z(n32929) );
  NANDN U33182 ( .A(n38248), .B(n32929), .Z(n32722) );
  AND U33183 ( .A(n32723), .B(n32722), .Z(n32945) );
  NANDN U33184 ( .A(n37526), .B(n32724), .Z(n32726) );
  XOR U33185 ( .A(b[51]), .B(a[95]), .Z(n33052) );
  NANDN U33186 ( .A(n37605), .B(n33052), .Z(n32725) );
  NAND U33187 ( .A(n32726), .B(n32725), .Z(n32944) );
  XOR U33188 ( .A(n32945), .B(n32944), .Z(n32947) );
  XNOR U33189 ( .A(n32946), .B(n32947), .Z(n33076) );
  XNOR U33190 ( .A(n33077), .B(n33076), .Z(n33078) );
  NANDN U33191 ( .A(n32728), .B(n32727), .Z(n32732) );
  OR U33192 ( .A(n32730), .B(n32729), .Z(n32731) );
  NAND U33193 ( .A(n32732), .B(n32731), .Z(n33079) );
  XNOR U33194 ( .A(n33078), .B(n33079), .Z(n32980) );
  NANDN U33195 ( .A(n32734), .B(n32733), .Z(n32738) );
  OR U33196 ( .A(n32736), .B(n32735), .Z(n32737) );
  NAND U33197 ( .A(n32738), .B(n32737), .Z(n32981) );
  XNOR U33198 ( .A(n32980), .B(n32981), .Z(n32982) );
  XOR U33199 ( .A(n32983), .B(n32982), .Z(n32957) );
  NANDN U33200 ( .A(n32740), .B(n32739), .Z(n32744) );
  NAND U33201 ( .A(n32742), .B(n32741), .Z(n32743) );
  AND U33202 ( .A(n32744), .B(n32743), .Z(n32956) );
  XNOR U33203 ( .A(n32957), .B(n32956), .Z(n32958) );
  XOR U33204 ( .A(n32959), .B(n32958), .Z(n32965) );
  XNOR U33205 ( .A(n32964), .B(n32965), .Z(n32896) );
  XNOR U33206 ( .A(n32897), .B(n32896), .Z(n32898) );
  XOR U33207 ( .A(n32899), .B(n32898), .Z(n32893) );
  NANDN U33208 ( .A(n32746), .B(n32745), .Z(n32750) );
  OR U33209 ( .A(n32748), .B(n32747), .Z(n32749) );
  AND U33210 ( .A(n32750), .B(n32749), .Z(n33087) );
  NANDN U33211 ( .A(n32752), .B(n32751), .Z(n32756) );
  NANDN U33212 ( .A(n32754), .B(n32753), .Z(n32755) );
  NAND U33213 ( .A(n32756), .B(n32755), .Z(n33086) );
  XNOR U33214 ( .A(n33087), .B(n33086), .Z(n33089) );
  NANDN U33215 ( .A(n32758), .B(n32757), .Z(n32762) );
  OR U33216 ( .A(n32760), .B(n32759), .Z(n32761) );
  NAND U33217 ( .A(n32762), .B(n32761), .Z(n33094) );
  NAND U33218 ( .A(n32764), .B(n32763), .Z(n32768) );
  NAND U33219 ( .A(n32766), .B(n32765), .Z(n32767) );
  AND U33220 ( .A(n32768), .B(n32767), .Z(n33093) );
  NANDN U33221 ( .A(n33875), .B(n32769), .Z(n32771) );
  XOR U33222 ( .A(a[121]), .B(b[25]), .Z(n32902) );
  NANDN U33223 ( .A(n33994), .B(n32902), .Z(n32770) );
  AND U33224 ( .A(n32771), .B(n32770), .Z(n33012) );
  NANDN U33225 ( .A(n33866), .B(n32772), .Z(n32774) );
  XOR U33226 ( .A(a[123]), .B(b[23]), .Z(n32905) );
  NANDN U33227 ( .A(n33644), .B(n32905), .Z(n32773) );
  AND U33228 ( .A(n32774), .B(n32773), .Z(n33011) );
  NANDN U33229 ( .A(n211), .B(n32775), .Z(n32777) );
  XOR U33230 ( .A(b[47]), .B(a[99]), .Z(n33022) );
  NANDN U33231 ( .A(n37172), .B(n33022), .Z(n32776) );
  NAND U33232 ( .A(n32777), .B(n32776), .Z(n33010) );
  XOR U33233 ( .A(n33011), .B(n33010), .Z(n33013) );
  XOR U33234 ( .A(n33012), .B(n33013), .Z(n33071) );
  NANDN U33235 ( .A(n32778), .B(n35309), .Z(n32780) );
  XOR U33236 ( .A(a[115]), .B(b[31]), .Z(n33046) );
  NANDN U33237 ( .A(n35145), .B(n33046), .Z(n32779) );
  AND U33238 ( .A(n32780), .B(n32779), .Z(n33066) );
  NANDN U33239 ( .A(n34634), .B(n32781), .Z(n32783) );
  XOR U33240 ( .A(a[117]), .B(b[29]), .Z(n33049) );
  NANDN U33241 ( .A(n34722), .B(n33049), .Z(n32782) );
  AND U33242 ( .A(n32783), .B(n32782), .Z(n33065) );
  NANDN U33243 ( .A(n37974), .B(n32784), .Z(n32786) );
  XOR U33244 ( .A(b[57]), .B(a[89]), .Z(n33058) );
  NANDN U33245 ( .A(n38031), .B(n33058), .Z(n32785) );
  NAND U33246 ( .A(n32786), .B(n32785), .Z(n33064) );
  XOR U33247 ( .A(n33065), .B(n33064), .Z(n33067) );
  XNOR U33248 ( .A(n33066), .B(n33067), .Z(n33070) );
  XNOR U33249 ( .A(n33071), .B(n33070), .Z(n33072) );
  NANDN U33250 ( .A(n32788), .B(n32787), .Z(n32792) );
  OR U33251 ( .A(n32790), .B(n32789), .Z(n32791) );
  NAND U33252 ( .A(n32792), .B(n32791), .Z(n33073) );
  XNOR U33253 ( .A(n33072), .B(n33073), .Z(n33083) );
  NANDN U33254 ( .A(n32996), .B(n32793), .Z(n32795) );
  XOR U33255 ( .A(a[125]), .B(b[21]), .Z(n32995) );
  NANDN U33256 ( .A(n33271), .B(n32995), .Z(n32794) );
  AND U33257 ( .A(n32795), .B(n32794), .Z(n33019) );
  NANDN U33258 ( .A(n38278), .B(n32796), .Z(n32798) );
  XOR U33259 ( .A(b[63]), .B(a[83]), .Z(n32932) );
  NANDN U33260 ( .A(n38279), .B(n32932), .Z(n32797) );
  AND U33261 ( .A(n32798), .B(n32797), .Z(n33017) );
  NANDN U33262 ( .A(n36991), .B(n32799), .Z(n32801) );
  XOR U33263 ( .A(b[45]), .B(a[101]), .Z(n32935) );
  NANDN U33264 ( .A(n37083), .B(n32935), .Z(n32800) );
  NAND U33265 ( .A(n32801), .B(n32800), .Z(n33016) );
  XNOR U33266 ( .A(n33017), .B(n33016), .Z(n33018) );
  XOR U33267 ( .A(n33019), .B(n33018), .Z(n32975) );
  NANDN U33268 ( .A(n37857), .B(n32802), .Z(n32804) );
  XOR U33269 ( .A(b[55]), .B(a[91]), .Z(n33055) );
  NANDN U33270 ( .A(n37911), .B(n33055), .Z(n32803) );
  AND U33271 ( .A(n32804), .B(n32803), .Z(n33042) );
  NANDN U33272 ( .A(n38090), .B(n32805), .Z(n32807) );
  XOR U33273 ( .A(b[59]), .B(a[87]), .Z(n33031) );
  NANDN U33274 ( .A(n38130), .B(n33031), .Z(n32806) );
  AND U33275 ( .A(n32807), .B(n32806), .Z(n33041) );
  NANDN U33276 ( .A(n35260), .B(n32808), .Z(n32810) );
  XOR U33277 ( .A(a[113]), .B(b[33]), .Z(n33061) );
  NANDN U33278 ( .A(n35456), .B(n33061), .Z(n32809) );
  NAND U33279 ( .A(n32810), .B(n32809), .Z(n33040) );
  XOR U33280 ( .A(n33041), .B(n33040), .Z(n33043) );
  XNOR U33281 ( .A(n33042), .B(n33043), .Z(n32974) );
  XOR U33282 ( .A(n32975), .B(n32974), .Z(n32977) );
  NANDN U33283 ( .A(n32812), .B(n32811), .Z(n32816) );
  OR U33284 ( .A(n32814), .B(n32813), .Z(n32815) );
  AND U33285 ( .A(n32816), .B(n32815), .Z(n32976) );
  XOR U33286 ( .A(n32977), .B(n32976), .Z(n33082) );
  XOR U33287 ( .A(n33083), .B(n33082), .Z(n33085) );
  NANDN U33288 ( .A(n32818), .B(n32817), .Z(n32822) );
  OR U33289 ( .A(n32820), .B(n32819), .Z(n32821) );
  AND U33290 ( .A(n32822), .B(n32821), .Z(n32926) );
  XNOR U33291 ( .A(a[127]), .B(b[19]), .Z(n32999) );
  OR U33292 ( .A(n32999), .B(n32823), .Z(n32826) );
  NAND U33293 ( .A(n33000), .B(n32824), .Z(n32825) );
  AND U33294 ( .A(n32826), .B(n32825), .Z(n32939) );
  NANDN U33295 ( .A(n36742), .B(n32827), .Z(n32829) );
  XOR U33296 ( .A(b[43]), .B(a[103]), .Z(n32908) );
  NANDN U33297 ( .A(n36891), .B(n32908), .Z(n32828) );
  NAND U33298 ( .A(n32829), .B(n32828), .Z(n32938) );
  XNOR U33299 ( .A(n32939), .B(n32938), .Z(n32940) );
  AND U33300 ( .A(b[63]), .B(a[81]), .Z(n32911) );
  IV U33301 ( .A(n32830), .Z(n32912) );
  XOR U33302 ( .A(n32911), .B(n32912), .Z(n32913) );
  XOR U33303 ( .A(n32846), .B(n32913), .Z(n32941) );
  XOR U33304 ( .A(n32940), .B(n32941), .Z(n32923) );
  NANDN U33305 ( .A(n36210), .B(n32831), .Z(n32833) );
  XOR U33306 ( .A(a[107]), .B(b[39]), .Z(n32989) );
  NANDN U33307 ( .A(n36347), .B(n32989), .Z(n32832) );
  AND U33308 ( .A(n32833), .B(n32832), .Z(n32920) );
  NANDN U33309 ( .A(n36480), .B(n32834), .Z(n32836) );
  XOR U33310 ( .A(b[41]), .B(a[105]), .Z(n32992) );
  NANDN U33311 ( .A(n36594), .B(n32992), .Z(n32835) );
  AND U33312 ( .A(n32836), .B(n32835), .Z(n32918) );
  NANDN U33313 ( .A(n35936), .B(n32837), .Z(n32839) );
  XOR U33314 ( .A(a[109]), .B(b[37]), .Z(n32986) );
  NANDN U33315 ( .A(n36047), .B(n32986), .Z(n32838) );
  NAND U33316 ( .A(n32839), .B(n32838), .Z(n32917) );
  XNOR U33317 ( .A(n32918), .B(n32917), .Z(n32919) );
  XOR U33318 ( .A(n32920), .B(n32919), .Z(n32924) );
  XNOR U33319 ( .A(n32923), .B(n32924), .Z(n32925) );
  XOR U33320 ( .A(n32926), .B(n32925), .Z(n32968) );
  NANDN U33321 ( .A(n32841), .B(n32840), .Z(n32845) );
  OR U33322 ( .A(n32843), .B(n32842), .Z(n32844) );
  AND U33323 ( .A(n32845), .B(n32844), .Z(n32969) );
  XOR U33324 ( .A(n32968), .B(n32969), .Z(n32971) );
  IV U33325 ( .A(n32846), .Z(n32914) );
  NANDN U33326 ( .A(n32914), .B(n32847), .Z(n32851) );
  NANDN U33327 ( .A(n32849), .B(n32848), .Z(n32850) );
  AND U33328 ( .A(n32851), .B(n32850), .Z(n32970) );
  XOR U33329 ( .A(n32971), .B(n32970), .Z(n33084) );
  XOR U33330 ( .A(n33085), .B(n33084), .Z(n32952) );
  NANDN U33331 ( .A(n32853), .B(n32852), .Z(n32857) );
  NANDN U33332 ( .A(n32855), .B(n32854), .Z(n32856) );
  AND U33333 ( .A(n32857), .B(n32856), .Z(n32951) );
  NANDN U33334 ( .A(n32859), .B(n32858), .Z(n32863) );
  NANDN U33335 ( .A(n32861), .B(n32860), .Z(n32862) );
  AND U33336 ( .A(n32863), .B(n32862), .Z(n32950) );
  XOR U33337 ( .A(n32951), .B(n32950), .Z(n32953) );
  XOR U33338 ( .A(n32952), .B(n32953), .Z(n33092) );
  XOR U33339 ( .A(n33093), .B(n33092), .Z(n33095) );
  XOR U33340 ( .A(n33094), .B(n33095), .Z(n33088) );
  XOR U33341 ( .A(n33089), .B(n33088), .Z(n32891) );
  NANDN U33342 ( .A(n32865), .B(n32864), .Z(n32869) );
  NANDN U33343 ( .A(n32867), .B(n32866), .Z(n32868) );
  AND U33344 ( .A(n32869), .B(n32868), .Z(n32890) );
  XNOR U33345 ( .A(n32891), .B(n32890), .Z(n32892) );
  XOR U33346 ( .A(n32893), .B(n32892), .Z(n32885) );
  XNOR U33347 ( .A(n32884), .B(n32885), .Z(n32886) );
  NANDN U33348 ( .A(n32871), .B(n32870), .Z(n32875) );
  NAND U33349 ( .A(n32873), .B(n32872), .Z(n32874) );
  NAND U33350 ( .A(n32875), .B(n32874), .Z(n32887) );
  XNOR U33351 ( .A(n32886), .B(n32887), .Z(n32878) );
  XOR U33352 ( .A(n32879), .B(n32878), .Z(n32881) );
  XNOR U33353 ( .A(n32880), .B(n32881), .Z(n32876) );
  XOR U33354 ( .A(n32877), .B(n32876), .Z(c[209]) );
  AND U33355 ( .A(n32877), .B(n32876), .Z(n33099) );
  NANDN U33356 ( .A(n32879), .B(n32878), .Z(n32883) );
  OR U33357 ( .A(n32881), .B(n32880), .Z(n32882) );
  AND U33358 ( .A(n32883), .B(n32882), .Z(n33102) );
  NANDN U33359 ( .A(n32885), .B(n32884), .Z(n32889) );
  NANDN U33360 ( .A(n32887), .B(n32886), .Z(n32888) );
  AND U33361 ( .A(n32889), .B(n32888), .Z(n33101) );
  NANDN U33362 ( .A(n32891), .B(n32890), .Z(n32895) );
  NANDN U33363 ( .A(n32893), .B(n32892), .Z(n32894) );
  AND U33364 ( .A(n32895), .B(n32894), .Z(n33109) );
  NANDN U33365 ( .A(n32897), .B(n32896), .Z(n32901) );
  NAND U33366 ( .A(n32899), .B(n32898), .Z(n32900) );
  AND U33367 ( .A(n32901), .B(n32900), .Z(n33106) );
  NANDN U33368 ( .A(n33875), .B(n32902), .Z(n32904) );
  XNOR U33369 ( .A(a[122]), .B(b[25]), .Z(n33154) );
  NANDN U33370 ( .A(n33154), .B(n34298), .Z(n32903) );
  AND U33371 ( .A(n32904), .B(n32903), .Z(n33241) );
  NANDN U33372 ( .A(n33866), .B(n32905), .Z(n32907) );
  XNOR U33373 ( .A(a[124]), .B(b[23]), .Z(n33157) );
  NANDN U33374 ( .A(n33157), .B(n33868), .Z(n32906) );
  AND U33375 ( .A(n32907), .B(n32906), .Z(n33239) );
  NANDN U33376 ( .A(n36742), .B(n32908), .Z(n32910) );
  XOR U33377 ( .A(b[43]), .B(a[104]), .Z(n33232) );
  NANDN U33378 ( .A(n36891), .B(n33232), .Z(n32909) );
  NAND U33379 ( .A(n32910), .B(n32909), .Z(n33238) );
  XNOR U33380 ( .A(n33239), .B(n33238), .Z(n33240) );
  XNOR U33381 ( .A(n33241), .B(n33240), .Z(n33136) );
  NANDN U33382 ( .A(n32912), .B(n32911), .Z(n32916) );
  ANDN U33383 ( .B(n32914), .A(n32913), .Z(n32915) );
  ANDN U33384 ( .B(n32916), .A(n32915), .Z(n33137) );
  XNOR U33385 ( .A(n33136), .B(n33137), .Z(n33139) );
  NANDN U33386 ( .A(n32918), .B(n32917), .Z(n32922) );
  NANDN U33387 ( .A(n32920), .B(n32919), .Z(n32921) );
  NAND U33388 ( .A(n32922), .B(n32921), .Z(n33138) );
  XOR U33389 ( .A(n33139), .B(n33138), .Z(n33149) );
  NANDN U33390 ( .A(n32924), .B(n32923), .Z(n32928) );
  NANDN U33391 ( .A(n32926), .B(n32925), .Z(n32927) );
  AND U33392 ( .A(n32928), .B(n32927), .Z(n33148) );
  XNOR U33393 ( .A(n33149), .B(n33148), .Z(n33150) );
  NANDN U33394 ( .A(n38247), .B(n32929), .Z(n32931) );
  XOR U33395 ( .A(b[61]), .B(a[86]), .Z(n33166) );
  NANDN U33396 ( .A(n38248), .B(n33166), .Z(n32930) );
  AND U33397 ( .A(n32931), .B(n32930), .Z(n33210) );
  NANDN U33398 ( .A(n38278), .B(n32932), .Z(n32934) );
  XOR U33399 ( .A(b[63]), .B(a[84]), .Z(n33229) );
  NANDN U33400 ( .A(n38279), .B(n33229), .Z(n32933) );
  AND U33401 ( .A(n32934), .B(n32933), .Z(n33209) );
  NANDN U33402 ( .A(n36991), .B(n32935), .Z(n32937) );
  XOR U33403 ( .A(b[45]), .B(a[102]), .Z(n33253) );
  NANDN U33404 ( .A(n37083), .B(n33253), .Z(n32936) );
  NAND U33405 ( .A(n32937), .B(n32936), .Z(n33208) );
  XOR U33406 ( .A(n33209), .B(n33208), .Z(n33211) );
  XOR U33407 ( .A(n33210), .B(n33211), .Z(n33197) );
  NANDN U33408 ( .A(n32939), .B(n32938), .Z(n32943) );
  NAND U33409 ( .A(n32941), .B(n32940), .Z(n32942) );
  AND U33410 ( .A(n32943), .B(n32942), .Z(n33196) );
  XNOR U33411 ( .A(n33197), .B(n33196), .Z(n33198) );
  NANDN U33412 ( .A(n32945), .B(n32944), .Z(n32949) );
  OR U33413 ( .A(n32947), .B(n32946), .Z(n32948) );
  NAND U33414 ( .A(n32949), .B(n32948), .Z(n33199) );
  XOR U33415 ( .A(n33198), .B(n33199), .Z(n33151) );
  XNOR U33416 ( .A(n33150), .B(n33151), .Z(n33287) );
  NANDN U33417 ( .A(n32951), .B(n32950), .Z(n32955) );
  OR U33418 ( .A(n32953), .B(n32952), .Z(n32954) );
  NAND U33419 ( .A(n32955), .B(n32954), .Z(n33288) );
  XNOR U33420 ( .A(n33287), .B(n33288), .Z(n33290) );
  NANDN U33421 ( .A(n32957), .B(n32956), .Z(n32961) );
  NANDN U33422 ( .A(n32959), .B(n32958), .Z(n32960) );
  AND U33423 ( .A(n32961), .B(n32960), .Z(n33289) );
  XOR U33424 ( .A(n33290), .B(n33289), .Z(n33301) );
  NANDN U33425 ( .A(n32963), .B(n32962), .Z(n32967) );
  NANDN U33426 ( .A(n32965), .B(n32964), .Z(n32966) );
  AND U33427 ( .A(n32967), .B(n32966), .Z(n33300) );
  NAND U33428 ( .A(n32969), .B(n32968), .Z(n32973) );
  NAND U33429 ( .A(n32971), .B(n32970), .Z(n32972) );
  NAND U33430 ( .A(n32973), .B(n32972), .Z(n33294) );
  NAND U33431 ( .A(n32975), .B(n32974), .Z(n32979) );
  NAND U33432 ( .A(n32977), .B(n32976), .Z(n32978) );
  NAND U33433 ( .A(n32979), .B(n32978), .Z(n33293) );
  XOR U33434 ( .A(n33294), .B(n33293), .Z(n33296) );
  NANDN U33435 ( .A(n32981), .B(n32980), .Z(n32985) );
  NAND U33436 ( .A(n32983), .B(n32982), .Z(n32984) );
  NAND U33437 ( .A(n32985), .B(n32984), .Z(n33295) );
  XOR U33438 ( .A(n33296), .B(n33295), .Z(n33115) );
  NANDN U33439 ( .A(n35936), .B(n32986), .Z(n32988) );
  XOR U33440 ( .A(a[110]), .B(b[37]), .Z(n33250) );
  NANDN U33441 ( .A(n36047), .B(n33250), .Z(n32987) );
  AND U33442 ( .A(n32988), .B(n32987), .Z(n33278) );
  NANDN U33443 ( .A(n36210), .B(n32989), .Z(n32991) );
  XOR U33444 ( .A(a[108]), .B(b[39]), .Z(n33268) );
  NANDN U33445 ( .A(n36347), .B(n33268), .Z(n32990) );
  AND U33446 ( .A(n32991), .B(n32990), .Z(n33276) );
  NANDN U33447 ( .A(n36480), .B(n32992), .Z(n32994) );
  XOR U33448 ( .A(b[41]), .B(a[106]), .Z(n33235) );
  NANDN U33449 ( .A(n36594), .B(n33235), .Z(n32993) );
  NAND U33450 ( .A(n32994), .B(n32993), .Z(n33275) );
  XNOR U33451 ( .A(n33276), .B(n33275), .Z(n33277) );
  XOR U33452 ( .A(n33278), .B(n33277), .Z(n33191) );
  NANDN U33453 ( .A(n32996), .B(n32995), .Z(n32998) );
  XOR U33454 ( .A(a[126]), .B(b[21]), .Z(n33272) );
  NANDN U33455 ( .A(n33271), .B(n33272), .Z(n32997) );
  AND U33456 ( .A(n32998), .B(n32997), .Z(n33284) );
  NAND U33457 ( .A(b[63]), .B(a[82]), .Z(n33281) );
  ANDN U33458 ( .B(n33000), .A(n32999), .Z(n33003) );
  NAND U33459 ( .A(b[19]), .B(n33001), .Z(n33002) );
  NANDN U33460 ( .A(n33003), .B(n33002), .Z(n33282) );
  XOR U33461 ( .A(n33281), .B(n33282), .Z(n33283) );
  XOR U33462 ( .A(n33284), .B(n33283), .Z(n33190) );
  XOR U33463 ( .A(n33191), .B(n33190), .Z(n33193) );
  NANDN U33464 ( .A(n33005), .B(n33004), .Z(n33009) );
  OR U33465 ( .A(n33007), .B(n33006), .Z(n33008) );
  AND U33466 ( .A(n33009), .B(n33008), .Z(n33192) );
  XOR U33467 ( .A(n33193), .B(n33192), .Z(n33204) );
  NANDN U33468 ( .A(n33011), .B(n33010), .Z(n33015) );
  OR U33469 ( .A(n33013), .B(n33012), .Z(n33014) );
  AND U33470 ( .A(n33015), .B(n33014), .Z(n33203) );
  NANDN U33471 ( .A(n33017), .B(n33016), .Z(n33021) );
  NANDN U33472 ( .A(n33019), .B(n33018), .Z(n33020) );
  NAND U33473 ( .A(n33021), .B(n33020), .Z(n33202) );
  XOR U33474 ( .A(n33203), .B(n33202), .Z(n33205) );
  XOR U33475 ( .A(n33204), .B(n33205), .Z(n33144) );
  NANDN U33476 ( .A(n211), .B(n33022), .Z(n33024) );
  XOR U33477 ( .A(b[47]), .B(a[100]), .Z(n33220) );
  NANDN U33478 ( .A(n37172), .B(n33220), .Z(n33023) );
  AND U33479 ( .A(n33024), .B(n33023), .Z(n33174) );
  NANDN U33480 ( .A(n37705), .B(n33025), .Z(n33027) );
  XOR U33481 ( .A(b[53]), .B(a[94]), .Z(n33223) );
  NANDN U33482 ( .A(n37778), .B(n33223), .Z(n33026) );
  AND U33483 ( .A(n33027), .B(n33026), .Z(n33173) );
  NANDN U33484 ( .A(n35611), .B(n33028), .Z(n33030) );
  XNOR U33485 ( .A(a[112]), .B(b[35]), .Z(n33247) );
  NANDN U33486 ( .A(n33247), .B(n35929), .Z(n33029) );
  NAND U33487 ( .A(n33030), .B(n33029), .Z(n33172) );
  XOR U33488 ( .A(n33173), .B(n33172), .Z(n33175) );
  XOR U33489 ( .A(n33174), .B(n33175), .Z(n33131) );
  NANDN U33490 ( .A(n38090), .B(n33031), .Z(n33033) );
  XOR U33491 ( .A(b[59]), .B(a[88]), .Z(n33163) );
  NANDN U33492 ( .A(n38130), .B(n33163), .Z(n33032) );
  AND U33493 ( .A(n33033), .B(n33032), .Z(n33186) );
  NANDN U33494 ( .A(n34223), .B(n33034), .Z(n33036) );
  XOR U33495 ( .A(a[120]), .B(b[27]), .Z(n33262) );
  NANDN U33496 ( .A(n34458), .B(n33262), .Z(n33035) );
  AND U33497 ( .A(n33036), .B(n33035), .Z(n33185) );
  NANDN U33498 ( .A(n212), .B(n33037), .Z(n33039) );
  XOR U33499 ( .A(b[49]), .B(a[98]), .Z(n33160) );
  NANDN U33500 ( .A(n37432), .B(n33160), .Z(n33038) );
  NAND U33501 ( .A(n33039), .B(n33038), .Z(n33184) );
  XOR U33502 ( .A(n33185), .B(n33184), .Z(n33187) );
  XNOR U33503 ( .A(n33186), .B(n33187), .Z(n33130) );
  XNOR U33504 ( .A(n33131), .B(n33130), .Z(n33132) );
  NANDN U33505 ( .A(n33041), .B(n33040), .Z(n33045) );
  OR U33506 ( .A(n33043), .B(n33042), .Z(n33044) );
  NAND U33507 ( .A(n33045), .B(n33044), .Z(n33133) );
  XNOR U33508 ( .A(n33132), .B(n33133), .Z(n33142) );
  NANDN U33509 ( .A(n34909), .B(n33046), .Z(n33048) );
  XOR U33510 ( .A(a[116]), .B(b[31]), .Z(n33256) );
  NANDN U33511 ( .A(n35145), .B(n33256), .Z(n33047) );
  AND U33512 ( .A(n33048), .B(n33047), .Z(n33180) );
  NANDN U33513 ( .A(n34634), .B(n33049), .Z(n33051) );
  XOR U33514 ( .A(a[118]), .B(b[29]), .Z(n33226) );
  NANDN U33515 ( .A(n34722), .B(n33226), .Z(n33050) );
  AND U33516 ( .A(n33051), .B(n33050), .Z(n33179) );
  NANDN U33517 ( .A(n37526), .B(n33052), .Z(n33054) );
  XOR U33518 ( .A(b[51]), .B(a[96]), .Z(n33169) );
  NANDN U33519 ( .A(n37605), .B(n33169), .Z(n33053) );
  NAND U33520 ( .A(n33054), .B(n33053), .Z(n33178) );
  XOR U33521 ( .A(n33179), .B(n33178), .Z(n33181) );
  XOR U33522 ( .A(n33180), .B(n33181), .Z(n33125) );
  NANDN U33523 ( .A(n37857), .B(n33055), .Z(n33057) );
  XOR U33524 ( .A(b[55]), .B(a[92]), .Z(n33259) );
  NANDN U33525 ( .A(n37911), .B(n33259), .Z(n33056) );
  AND U33526 ( .A(n33057), .B(n33056), .Z(n33216) );
  NANDN U33527 ( .A(n37974), .B(n33058), .Z(n33060) );
  XOR U33528 ( .A(b[57]), .B(a[90]), .Z(n33265) );
  NANDN U33529 ( .A(n38031), .B(n33265), .Z(n33059) );
  AND U33530 ( .A(n33060), .B(n33059), .Z(n33215) );
  NANDN U33531 ( .A(n35260), .B(n33061), .Z(n33063) );
  XOR U33532 ( .A(a[114]), .B(b[33]), .Z(n33244) );
  NANDN U33533 ( .A(n35456), .B(n33244), .Z(n33062) );
  NAND U33534 ( .A(n33063), .B(n33062), .Z(n33214) );
  XOR U33535 ( .A(n33215), .B(n33214), .Z(n33217) );
  XNOR U33536 ( .A(n33216), .B(n33217), .Z(n33124) );
  XNOR U33537 ( .A(n33125), .B(n33124), .Z(n33126) );
  NANDN U33538 ( .A(n33065), .B(n33064), .Z(n33069) );
  OR U33539 ( .A(n33067), .B(n33066), .Z(n33068) );
  NAND U33540 ( .A(n33069), .B(n33068), .Z(n33127) );
  XOR U33541 ( .A(n33126), .B(n33127), .Z(n33143) );
  XOR U33542 ( .A(n33142), .B(n33143), .Z(n33145) );
  XOR U33543 ( .A(n33144), .B(n33145), .Z(n33120) );
  NANDN U33544 ( .A(n33071), .B(n33070), .Z(n33075) );
  NANDN U33545 ( .A(n33073), .B(n33072), .Z(n33074) );
  AND U33546 ( .A(n33075), .B(n33074), .Z(n33118) );
  NANDN U33547 ( .A(n33077), .B(n33076), .Z(n33081) );
  NANDN U33548 ( .A(n33079), .B(n33078), .Z(n33080) );
  NAND U33549 ( .A(n33081), .B(n33080), .Z(n33119) );
  XOR U33550 ( .A(n33118), .B(n33119), .Z(n33121) );
  XOR U33551 ( .A(n33120), .B(n33121), .Z(n33113) );
  XNOR U33552 ( .A(n33113), .B(n33112), .Z(n33114) );
  XNOR U33553 ( .A(n33115), .B(n33114), .Z(n33299) );
  XOR U33554 ( .A(n33300), .B(n33299), .Z(n33302) );
  XOR U33555 ( .A(n33301), .B(n33302), .Z(n33308) );
  NANDN U33556 ( .A(n33087), .B(n33086), .Z(n33091) );
  NAND U33557 ( .A(n33089), .B(n33088), .Z(n33090) );
  AND U33558 ( .A(n33091), .B(n33090), .Z(n33305) );
  NAND U33559 ( .A(n33093), .B(n33092), .Z(n33097) );
  NAND U33560 ( .A(n33095), .B(n33094), .Z(n33096) );
  NAND U33561 ( .A(n33097), .B(n33096), .Z(n33306) );
  XNOR U33562 ( .A(n33305), .B(n33306), .Z(n33307) );
  XOR U33563 ( .A(n33308), .B(n33307), .Z(n33107) );
  XNOR U33564 ( .A(n33106), .B(n33107), .Z(n33108) );
  XNOR U33565 ( .A(n33109), .B(n33108), .Z(n33100) );
  XOR U33566 ( .A(n33101), .B(n33100), .Z(n33103) );
  XNOR U33567 ( .A(n33102), .B(n33103), .Z(n33098) );
  XOR U33568 ( .A(n33099), .B(n33098), .Z(c[210]) );
  AND U33569 ( .A(n33099), .B(n33098), .Z(n33312) );
  NANDN U33570 ( .A(n33101), .B(n33100), .Z(n33105) );
  OR U33571 ( .A(n33103), .B(n33102), .Z(n33104) );
  AND U33572 ( .A(n33105), .B(n33104), .Z(n33315) );
  NANDN U33573 ( .A(n33107), .B(n33106), .Z(n33111) );
  NANDN U33574 ( .A(n33109), .B(n33108), .Z(n33110) );
  AND U33575 ( .A(n33111), .B(n33110), .Z(n33314) );
  NANDN U33576 ( .A(n33113), .B(n33112), .Z(n33117) );
  NAND U33577 ( .A(n33115), .B(n33114), .Z(n33116) );
  AND U33578 ( .A(n33117), .B(n33116), .Z(n33334) );
  NANDN U33579 ( .A(n33119), .B(n33118), .Z(n33123) );
  OR U33580 ( .A(n33121), .B(n33120), .Z(n33122) );
  AND U33581 ( .A(n33123), .B(n33122), .Z(n33352) );
  NANDN U33582 ( .A(n33125), .B(n33124), .Z(n33129) );
  NANDN U33583 ( .A(n33127), .B(n33126), .Z(n33128) );
  AND U33584 ( .A(n33129), .B(n33128), .Z(n33338) );
  NANDN U33585 ( .A(n33131), .B(n33130), .Z(n33135) );
  NANDN U33586 ( .A(n33133), .B(n33132), .Z(n33134) );
  NAND U33587 ( .A(n33135), .B(n33134), .Z(n33337) );
  XNOR U33588 ( .A(n33338), .B(n33337), .Z(n33340) );
  NANDN U33589 ( .A(n33137), .B(n33136), .Z(n33141) );
  NAND U33590 ( .A(n33139), .B(n33138), .Z(n33140) );
  AND U33591 ( .A(n33141), .B(n33140), .Z(n33339) );
  XOR U33592 ( .A(n33340), .B(n33339), .Z(n33350) );
  NANDN U33593 ( .A(n33143), .B(n33142), .Z(n33147) );
  OR U33594 ( .A(n33145), .B(n33144), .Z(n33146) );
  AND U33595 ( .A(n33147), .B(n33146), .Z(n33349) );
  XNOR U33596 ( .A(n33350), .B(n33349), .Z(n33351) );
  XNOR U33597 ( .A(n33352), .B(n33351), .Z(n33331) );
  NANDN U33598 ( .A(n33149), .B(n33148), .Z(n33153) );
  NANDN U33599 ( .A(n33151), .B(n33150), .Z(n33152) );
  AND U33600 ( .A(n33153), .B(n33152), .Z(n33357) );
  NANDN U33601 ( .A(n33154), .B(n34297), .Z(n33156) );
  XNOR U33602 ( .A(a[123]), .B(b[25]), .Z(n33370) );
  NANDN U33603 ( .A(n33370), .B(n34298), .Z(n33155) );
  NAND U33604 ( .A(n33156), .B(n33155), .Z(n33393) );
  NANDN U33605 ( .A(n33157), .B(n33492), .Z(n33159) );
  XNOR U33606 ( .A(a[125]), .B(b[23]), .Z(n33493) );
  NANDN U33607 ( .A(n33493), .B(n33868), .Z(n33158) );
  NAND U33608 ( .A(n33159), .B(n33158), .Z(n33392) );
  NAND U33609 ( .A(n37536), .B(n33160), .Z(n33162) );
  XNOR U33610 ( .A(b[49]), .B(a[99]), .Z(n33382) );
  NANDN U33611 ( .A(n33382), .B(n37537), .Z(n33161) );
  NAND U33612 ( .A(n33162), .B(n33161), .Z(n33391) );
  XOR U33613 ( .A(n33392), .B(n33391), .Z(n33394) );
  XNOR U33614 ( .A(n33393), .B(n33394), .Z(n33439) );
  NANDN U33615 ( .A(n38090), .B(n33163), .Z(n33165) );
  XOR U33616 ( .A(b[59]), .B(a[89]), .Z(n33379) );
  NANDN U33617 ( .A(n38130), .B(n33379), .Z(n33164) );
  AND U33618 ( .A(n33165), .B(n33164), .Z(n33504) );
  NANDN U33619 ( .A(n38247), .B(n33166), .Z(n33168) );
  XOR U33620 ( .A(b[61]), .B(a[87]), .Z(n33496) );
  NANDN U33621 ( .A(n38248), .B(n33496), .Z(n33167) );
  AND U33622 ( .A(n33168), .B(n33167), .Z(n33503) );
  NANDN U33623 ( .A(n37526), .B(n33169), .Z(n33171) );
  XOR U33624 ( .A(b[51]), .B(a[97]), .Z(n33426) );
  NANDN U33625 ( .A(n37605), .B(n33426), .Z(n33170) );
  NAND U33626 ( .A(n33171), .B(n33170), .Z(n33502) );
  XOR U33627 ( .A(n33503), .B(n33502), .Z(n33505) );
  XNOR U33628 ( .A(n33504), .B(n33505), .Z(n33438) );
  XOR U33629 ( .A(n33439), .B(n33438), .Z(n33441) );
  NANDN U33630 ( .A(n33173), .B(n33172), .Z(n33177) );
  OR U33631 ( .A(n33175), .B(n33174), .Z(n33176) );
  AND U33632 ( .A(n33177), .B(n33176), .Z(n33440) );
  XOR U33633 ( .A(n33441), .B(n33440), .Z(n33520) );
  NANDN U33634 ( .A(n33179), .B(n33178), .Z(n33183) );
  OR U33635 ( .A(n33181), .B(n33180), .Z(n33182) );
  AND U33636 ( .A(n33183), .B(n33182), .Z(n33519) );
  NANDN U33637 ( .A(n33185), .B(n33184), .Z(n33189) );
  OR U33638 ( .A(n33187), .B(n33186), .Z(n33188) );
  NAND U33639 ( .A(n33189), .B(n33188), .Z(n33518) );
  XOR U33640 ( .A(n33519), .B(n33518), .Z(n33521) );
  XOR U33641 ( .A(n33520), .B(n33521), .Z(n33344) );
  NAND U33642 ( .A(n33191), .B(n33190), .Z(n33195) );
  NAND U33643 ( .A(n33193), .B(n33192), .Z(n33194) );
  NAND U33644 ( .A(n33195), .B(n33194), .Z(n33343) );
  XNOR U33645 ( .A(n33344), .B(n33343), .Z(n33346) );
  NANDN U33646 ( .A(n33197), .B(n33196), .Z(n33201) );
  NANDN U33647 ( .A(n33199), .B(n33198), .Z(n33200) );
  NAND U33648 ( .A(n33201), .B(n33200), .Z(n33345) );
  XOR U33649 ( .A(n33346), .B(n33345), .Z(n33356) );
  NANDN U33650 ( .A(n33203), .B(n33202), .Z(n33207) );
  OR U33651 ( .A(n33205), .B(n33204), .Z(n33206) );
  AND U33652 ( .A(n33207), .B(n33206), .Z(n33474) );
  NANDN U33653 ( .A(n33209), .B(n33208), .Z(n33213) );
  OR U33654 ( .A(n33211), .B(n33210), .Z(n33212) );
  AND U33655 ( .A(n33213), .B(n33212), .Z(n33432) );
  NANDN U33656 ( .A(n33215), .B(n33214), .Z(n33219) );
  OR U33657 ( .A(n33217), .B(n33216), .Z(n33218) );
  NAND U33658 ( .A(n33219), .B(n33218), .Z(n33433) );
  XNOR U33659 ( .A(n33432), .B(n33433), .Z(n33435) );
  NANDN U33660 ( .A(n211), .B(n33220), .Z(n33222) );
  XOR U33661 ( .A(b[47]), .B(a[101]), .Z(n33373) );
  NANDN U33662 ( .A(n37172), .B(n33373), .Z(n33221) );
  AND U33663 ( .A(n33222), .B(n33221), .Z(n33461) );
  NANDN U33664 ( .A(n37705), .B(n33223), .Z(n33225) );
  XOR U33665 ( .A(b[53]), .B(a[95]), .Z(n33444) );
  NANDN U33666 ( .A(n37778), .B(n33444), .Z(n33224) );
  AND U33667 ( .A(n33225), .B(n33224), .Z(n33460) );
  NANDN U33668 ( .A(n34634), .B(n33226), .Z(n33228) );
  XOR U33669 ( .A(a[119]), .B(b[29]), .Z(n33376) );
  NANDN U33670 ( .A(n34722), .B(n33376), .Z(n33227) );
  NAND U33671 ( .A(n33228), .B(n33227), .Z(n33459) );
  XOR U33672 ( .A(n33460), .B(n33459), .Z(n33462) );
  XOR U33673 ( .A(n33461), .B(n33462), .Z(n33466) );
  NANDN U33674 ( .A(n38278), .B(n33229), .Z(n33231) );
  XOR U33675 ( .A(b[63]), .B(a[85]), .Z(n33409) );
  NANDN U33676 ( .A(n38279), .B(n33409), .Z(n33230) );
  AND U33677 ( .A(n33231), .B(n33230), .Z(n33404) );
  NANDN U33678 ( .A(n36742), .B(n33232), .Z(n33234) );
  XOR U33679 ( .A(b[43]), .B(a[105]), .Z(n33499) );
  NANDN U33680 ( .A(n36891), .B(n33499), .Z(n33233) );
  NAND U33681 ( .A(n33234), .B(n33233), .Z(n33403) );
  XNOR U33682 ( .A(n33404), .B(n33403), .Z(n33406) );
  NANDN U33683 ( .A(n36480), .B(n33235), .Z(n33237) );
  XOR U33684 ( .A(b[41]), .B(a[107]), .Z(n33417) );
  NANDN U33685 ( .A(n36594), .B(n33417), .Z(n33236) );
  AND U33686 ( .A(n33237), .B(n33236), .Z(n33454) );
  AND U33687 ( .A(b[63]), .B(a[83]), .Z(n33453) );
  XOR U33688 ( .A(n33454), .B(n33453), .Z(n33456) );
  XOR U33689 ( .A(n33281), .B(n33456), .Z(n33405) );
  XNOR U33690 ( .A(n33406), .B(n33405), .Z(n33465) );
  XNOR U33691 ( .A(n33466), .B(n33465), .Z(n33467) );
  NANDN U33692 ( .A(n33239), .B(n33238), .Z(n33243) );
  NANDN U33693 ( .A(n33241), .B(n33240), .Z(n33242) );
  NAND U33694 ( .A(n33243), .B(n33242), .Z(n33468) );
  XNOR U33695 ( .A(n33467), .B(n33468), .Z(n33434) );
  XOR U33696 ( .A(n33435), .B(n33434), .Z(n33472) );
  NAND U33697 ( .A(n35654), .B(n33244), .Z(n33246) );
  XNOR U33698 ( .A(a[115]), .B(b[33]), .Z(n33483) );
  NANDN U33699 ( .A(n33483), .B(n35655), .Z(n33245) );
  NAND U33700 ( .A(n33246), .B(n33245), .Z(n33363) );
  NANDN U33701 ( .A(n33247), .B(n35928), .Z(n33249) );
  XNOR U33702 ( .A(a[113]), .B(b[35]), .Z(n33450) );
  NANDN U33703 ( .A(n33450), .B(n35929), .Z(n33248) );
  NAND U33704 ( .A(n33249), .B(n33248), .Z(n33361) );
  NANDN U33705 ( .A(n35936), .B(n33250), .Z(n33252) );
  XOR U33706 ( .A(a[111]), .B(b[37]), .Z(n33429) );
  NANDN U33707 ( .A(n36047), .B(n33429), .Z(n33251) );
  AND U33708 ( .A(n33252), .B(n33251), .Z(n33479) );
  NANDN U33709 ( .A(n36991), .B(n33253), .Z(n33255) );
  XOR U33710 ( .A(b[45]), .B(a[103]), .Z(n33423) );
  NANDN U33711 ( .A(n37083), .B(n33423), .Z(n33254) );
  AND U33712 ( .A(n33255), .B(n33254), .Z(n33478) );
  NANDN U33713 ( .A(n34909), .B(n33256), .Z(n33258) );
  XOR U33714 ( .A(a[117]), .B(b[31]), .Z(n33486) );
  NANDN U33715 ( .A(n35145), .B(n33486), .Z(n33257) );
  NAND U33716 ( .A(n33258), .B(n33257), .Z(n33477) );
  XOR U33717 ( .A(n33478), .B(n33477), .Z(n33480) );
  XOR U33718 ( .A(n33479), .B(n33480), .Z(n33362) );
  XOR U33719 ( .A(n33361), .B(n33362), .Z(n33364) );
  XNOR U33720 ( .A(n33363), .B(n33364), .Z(n33399) );
  NANDN U33721 ( .A(n37857), .B(n33259), .Z(n33261) );
  XOR U33722 ( .A(b[55]), .B(a[93]), .Z(n33447) );
  NANDN U33723 ( .A(n37911), .B(n33447), .Z(n33260) );
  AND U33724 ( .A(n33261), .B(n33260), .Z(n33387) );
  NANDN U33725 ( .A(n34223), .B(n33262), .Z(n33264) );
  XOR U33726 ( .A(a[121]), .B(b[27]), .Z(n33367) );
  NANDN U33727 ( .A(n34458), .B(n33367), .Z(n33263) );
  AND U33728 ( .A(n33264), .B(n33263), .Z(n33386) );
  NANDN U33729 ( .A(n37974), .B(n33265), .Z(n33267) );
  XOR U33730 ( .A(b[57]), .B(a[91]), .Z(n33489) );
  NANDN U33731 ( .A(n38031), .B(n33489), .Z(n33266) );
  NAND U33732 ( .A(n33267), .B(n33266), .Z(n33385) );
  XOR U33733 ( .A(n33386), .B(n33385), .Z(n33388) );
  XOR U33734 ( .A(n33387), .B(n33388), .Z(n33398) );
  NANDN U33735 ( .A(n36210), .B(n33268), .Z(n33270) );
  XOR U33736 ( .A(a[109]), .B(b[39]), .Z(n33420) );
  NANDN U33737 ( .A(n36347), .B(n33420), .Z(n33269) );
  AND U33738 ( .A(n33270), .B(n33269), .Z(n33510) );
  XNOR U33739 ( .A(a[127]), .B(b[21]), .Z(n33412) );
  OR U33740 ( .A(n33412), .B(n33271), .Z(n33274) );
  NAND U33741 ( .A(n33413), .B(n33272), .Z(n33273) );
  NAND U33742 ( .A(n33274), .B(n33273), .Z(n33508) );
  XOR U33743 ( .A(n33509), .B(n33508), .Z(n33511) );
  XNOR U33744 ( .A(n33510), .B(n33511), .Z(n33397) );
  XOR U33745 ( .A(n33398), .B(n33397), .Z(n33400) );
  XOR U33746 ( .A(n33399), .B(n33400), .Z(n33516) );
  NANDN U33747 ( .A(n33276), .B(n33275), .Z(n33280) );
  NANDN U33748 ( .A(n33278), .B(n33277), .Z(n33279) );
  AND U33749 ( .A(n33280), .B(n33279), .Z(n33515) );
  IV U33750 ( .A(n33281), .Z(n33455) );
  NANDN U33751 ( .A(n33455), .B(n33282), .Z(n33286) );
  NANDN U33752 ( .A(n33284), .B(n33283), .Z(n33285) );
  NAND U33753 ( .A(n33286), .B(n33285), .Z(n33514) );
  XNOR U33754 ( .A(n33515), .B(n33514), .Z(n33517) );
  XOR U33755 ( .A(n33516), .B(n33517), .Z(n33471) );
  XNOR U33756 ( .A(n33472), .B(n33471), .Z(n33473) );
  XNOR U33757 ( .A(n33474), .B(n33473), .Z(n33355) );
  XOR U33758 ( .A(n33356), .B(n33355), .Z(n33358) );
  XOR U33759 ( .A(n33357), .B(n33358), .Z(n33332) );
  XNOR U33760 ( .A(n33331), .B(n33332), .Z(n33333) );
  XOR U33761 ( .A(n33334), .B(n33333), .Z(n33327) );
  NANDN U33762 ( .A(n33288), .B(n33287), .Z(n33292) );
  NAND U33763 ( .A(n33290), .B(n33289), .Z(n33291) );
  AND U33764 ( .A(n33292), .B(n33291), .Z(n33326) );
  NAND U33765 ( .A(n33294), .B(n33293), .Z(n33298) );
  NAND U33766 ( .A(n33296), .B(n33295), .Z(n33297) );
  NAND U33767 ( .A(n33298), .B(n33297), .Z(n33325) );
  XOR U33768 ( .A(n33326), .B(n33325), .Z(n33328) );
  XOR U33769 ( .A(n33327), .B(n33328), .Z(n33320) );
  NANDN U33770 ( .A(n33300), .B(n33299), .Z(n33304) );
  OR U33771 ( .A(n33302), .B(n33301), .Z(n33303) );
  NAND U33772 ( .A(n33304), .B(n33303), .Z(n33319) );
  XNOR U33773 ( .A(n33320), .B(n33319), .Z(n33322) );
  NANDN U33774 ( .A(n33306), .B(n33305), .Z(n33310) );
  NANDN U33775 ( .A(n33308), .B(n33307), .Z(n33309) );
  AND U33776 ( .A(n33310), .B(n33309), .Z(n33321) );
  XNOR U33777 ( .A(n33322), .B(n33321), .Z(n33313) );
  XOR U33778 ( .A(n33314), .B(n33313), .Z(n33316) );
  XNOR U33779 ( .A(n33315), .B(n33316), .Z(n33311) );
  XOR U33780 ( .A(n33312), .B(n33311), .Z(c[211]) );
  AND U33781 ( .A(n33312), .B(n33311), .Z(n33525) );
  NANDN U33782 ( .A(n33314), .B(n33313), .Z(n33318) );
  OR U33783 ( .A(n33316), .B(n33315), .Z(n33317) );
  AND U33784 ( .A(n33318), .B(n33317), .Z(n33528) );
  NANDN U33785 ( .A(n33320), .B(n33319), .Z(n33324) );
  NAND U33786 ( .A(n33322), .B(n33321), .Z(n33323) );
  AND U33787 ( .A(n33324), .B(n33323), .Z(n33526) );
  NANDN U33788 ( .A(n33326), .B(n33325), .Z(n33330) );
  OR U33789 ( .A(n33328), .B(n33327), .Z(n33329) );
  AND U33790 ( .A(n33330), .B(n33329), .Z(n33535) );
  NANDN U33791 ( .A(n33332), .B(n33331), .Z(n33336) );
  NAND U33792 ( .A(n33334), .B(n33333), .Z(n33335) );
  AND U33793 ( .A(n33336), .B(n33335), .Z(n33532) );
  NANDN U33794 ( .A(n33338), .B(n33337), .Z(n33342) );
  NAND U33795 ( .A(n33340), .B(n33339), .Z(n33341) );
  AND U33796 ( .A(n33342), .B(n33341), .Z(n33722) );
  NANDN U33797 ( .A(n33344), .B(n33343), .Z(n33348) );
  NAND U33798 ( .A(n33346), .B(n33345), .Z(n33347) );
  NAND U33799 ( .A(n33348), .B(n33347), .Z(n33723) );
  XNOR U33800 ( .A(n33722), .B(n33723), .Z(n33725) );
  NANDN U33801 ( .A(n33350), .B(n33349), .Z(n33354) );
  NANDN U33802 ( .A(n33352), .B(n33351), .Z(n33353) );
  NAND U33803 ( .A(n33354), .B(n33353), .Z(n33724) );
  XOR U33804 ( .A(n33725), .B(n33724), .Z(n33719) );
  NANDN U33805 ( .A(n33356), .B(n33355), .Z(n33360) );
  NANDN U33806 ( .A(n33358), .B(n33357), .Z(n33359) );
  AND U33807 ( .A(n33360), .B(n33359), .Z(n33716) );
  NAND U33808 ( .A(n33362), .B(n33361), .Z(n33366) );
  NAND U33809 ( .A(n33364), .B(n33363), .Z(n33365) );
  AND U33810 ( .A(n33366), .B(n33365), .Z(n33677) );
  NANDN U33811 ( .A(n34223), .B(n33367), .Z(n33369) );
  XOR U33812 ( .A(a[122]), .B(b[27]), .Z(n33610) );
  NANDN U33813 ( .A(n34458), .B(n33610), .Z(n33368) );
  AND U33814 ( .A(n33369), .B(n33368), .Z(n33615) );
  NANDN U33815 ( .A(n33370), .B(n34297), .Z(n33372) );
  XOR U33816 ( .A(a[124]), .B(b[25]), .Z(n33656) );
  NANDN U33817 ( .A(n33994), .B(n33656), .Z(n33371) );
  AND U33818 ( .A(n33372), .B(n33371), .Z(n33614) );
  NANDN U33819 ( .A(n211), .B(n33373), .Z(n33375) );
  XOR U33820 ( .A(b[47]), .B(a[102]), .Z(n33659) );
  NANDN U33821 ( .A(n37172), .B(n33659), .Z(n33374) );
  NAND U33822 ( .A(n33375), .B(n33374), .Z(n33613) );
  XOR U33823 ( .A(n33614), .B(n33613), .Z(n33616) );
  XOR U33824 ( .A(n33615), .B(n33616), .Z(n33681) );
  NANDN U33825 ( .A(n34634), .B(n33376), .Z(n33378) );
  XOR U33826 ( .A(a[120]), .B(b[29]), .Z(n33556) );
  NANDN U33827 ( .A(n34722), .B(n33556), .Z(n33377) );
  AND U33828 ( .A(n33378), .B(n33377), .Z(n33621) );
  NANDN U33829 ( .A(n38090), .B(n33379), .Z(n33381) );
  XOR U33830 ( .A(b[59]), .B(a[90]), .Z(n33653) );
  NANDN U33831 ( .A(n38130), .B(n33653), .Z(n33380) );
  AND U33832 ( .A(n33381), .B(n33380), .Z(n33620) );
  NANDN U33833 ( .A(n33382), .B(n37536), .Z(n33384) );
  XOR U33834 ( .A(b[49]), .B(a[100]), .Z(n33550) );
  NANDN U33835 ( .A(n37432), .B(n33550), .Z(n33383) );
  NAND U33836 ( .A(n33384), .B(n33383), .Z(n33619) );
  XOR U33837 ( .A(n33620), .B(n33619), .Z(n33622) );
  XNOR U33838 ( .A(n33621), .B(n33622), .Z(n33680) );
  XNOR U33839 ( .A(n33681), .B(n33680), .Z(n33682) );
  NANDN U33840 ( .A(n33386), .B(n33385), .Z(n33390) );
  OR U33841 ( .A(n33388), .B(n33387), .Z(n33389) );
  NAND U33842 ( .A(n33390), .B(n33389), .Z(n33683) );
  XNOR U33843 ( .A(n33682), .B(n33683), .Z(n33675) );
  NAND U33844 ( .A(n33392), .B(n33391), .Z(n33396) );
  NAND U33845 ( .A(n33394), .B(n33393), .Z(n33395) );
  AND U33846 ( .A(n33396), .B(n33395), .Z(n33674) );
  XOR U33847 ( .A(n33675), .B(n33674), .Z(n33676) );
  XOR U33848 ( .A(n33677), .B(n33676), .Z(n33592) );
  NANDN U33849 ( .A(n33398), .B(n33397), .Z(n33402) );
  NANDN U33850 ( .A(n33400), .B(n33399), .Z(n33401) );
  AND U33851 ( .A(n33402), .B(n33401), .Z(n33589) );
  NANDN U33852 ( .A(n33404), .B(n33403), .Z(n33408) );
  NAND U33853 ( .A(n33406), .B(n33405), .Z(n33407) );
  AND U33854 ( .A(n33408), .B(n33407), .Z(n33632) );
  NANDN U33855 ( .A(n38278), .B(n33409), .Z(n33411) );
  XOR U33856 ( .A(b[63]), .B(a[86]), .Z(n33577) );
  NANDN U33857 ( .A(n38279), .B(n33577), .Z(n33410) );
  AND U33858 ( .A(n33411), .B(n33410), .Z(n33586) );
  NAND U33859 ( .A(b[63]), .B(a[84]), .Z(n33778) );
  ANDN U33860 ( .B(n33413), .A(n33412), .Z(n33416) );
  NAND U33861 ( .A(b[21]), .B(n33414), .Z(n33415) );
  NANDN U33862 ( .A(n33416), .B(n33415), .Z(n33583) );
  XOR U33863 ( .A(n33778), .B(n33583), .Z(n33585) );
  XNOR U33864 ( .A(n33586), .B(n33585), .Z(n33631) );
  XNOR U33865 ( .A(n33632), .B(n33631), .Z(n33633) );
  NANDN U33866 ( .A(n36480), .B(n33417), .Z(n33419) );
  XOR U33867 ( .A(a[108]), .B(b[41]), .Z(n33601) );
  NANDN U33868 ( .A(n36594), .B(n33601), .Z(n33418) );
  AND U33869 ( .A(n33419), .B(n33418), .Z(n33628) );
  NANDN U33870 ( .A(n36210), .B(n33420), .Z(n33422) );
  XOR U33871 ( .A(a[110]), .B(b[39]), .Z(n33559) );
  NANDN U33872 ( .A(n36347), .B(n33559), .Z(n33421) );
  AND U33873 ( .A(n33422), .B(n33421), .Z(n33626) );
  NANDN U33874 ( .A(n36991), .B(n33423), .Z(n33425) );
  XOR U33875 ( .A(b[45]), .B(a[104]), .Z(n33650) );
  NANDN U33876 ( .A(n37083), .B(n33650), .Z(n33424) );
  AND U33877 ( .A(n33425), .B(n33424), .Z(n33574) );
  NANDN U33878 ( .A(n37526), .B(n33426), .Z(n33428) );
  XOR U33879 ( .A(b[51]), .B(a[98]), .Z(n33553) );
  NANDN U33880 ( .A(n37605), .B(n33553), .Z(n33427) );
  AND U33881 ( .A(n33428), .B(n33427), .Z(n33572) );
  NANDN U33882 ( .A(n35936), .B(n33429), .Z(n33431) );
  XOR U33883 ( .A(a[112]), .B(b[37]), .Z(n33568) );
  NANDN U33884 ( .A(n36047), .B(n33568), .Z(n33430) );
  NAND U33885 ( .A(n33431), .B(n33430), .Z(n33571) );
  XNOR U33886 ( .A(n33572), .B(n33571), .Z(n33573) );
  XNOR U33887 ( .A(n33574), .B(n33573), .Z(n33625) );
  XNOR U33888 ( .A(n33626), .B(n33625), .Z(n33627) );
  XOR U33889 ( .A(n33628), .B(n33627), .Z(n33634) );
  XOR U33890 ( .A(n33633), .B(n33634), .Z(n33590) );
  XNOR U33891 ( .A(n33589), .B(n33590), .Z(n33591) );
  XNOR U33892 ( .A(n33592), .B(n33591), .Z(n33710) );
  NANDN U33893 ( .A(n33433), .B(n33432), .Z(n33437) );
  NAND U33894 ( .A(n33435), .B(n33434), .Z(n33436) );
  NAND U33895 ( .A(n33437), .B(n33436), .Z(n33711) );
  XNOR U33896 ( .A(n33710), .B(n33711), .Z(n33713) );
  NAND U33897 ( .A(n33439), .B(n33438), .Z(n33443) );
  NAND U33898 ( .A(n33441), .B(n33440), .Z(n33442) );
  AND U33899 ( .A(n33443), .B(n33442), .Z(n33540) );
  NANDN U33900 ( .A(n37705), .B(n33444), .Z(n33446) );
  XOR U33901 ( .A(b[53]), .B(a[96]), .Z(n33607) );
  NANDN U33902 ( .A(n37778), .B(n33607), .Z(n33445) );
  AND U33903 ( .A(n33446), .B(n33445), .Z(n33639) );
  NANDN U33904 ( .A(n37857), .B(n33447), .Z(n33449) );
  XOR U33905 ( .A(b[55]), .B(a[94]), .Z(n33595) );
  NANDN U33906 ( .A(n37911), .B(n33595), .Z(n33448) );
  AND U33907 ( .A(n33449), .B(n33448), .Z(n33638) );
  NANDN U33908 ( .A(n33450), .B(n35928), .Z(n33452) );
  XOR U33909 ( .A(a[114]), .B(b[35]), .Z(n33604) );
  NANDN U33910 ( .A(n35801), .B(n33604), .Z(n33451) );
  NAND U33911 ( .A(n33452), .B(n33451), .Z(n33637) );
  XOR U33912 ( .A(n33638), .B(n33637), .Z(n33640) );
  XOR U33913 ( .A(n33639), .B(n33640), .Z(n33545) );
  NANDN U33914 ( .A(n33454), .B(n33453), .Z(n33458) );
  NANDN U33915 ( .A(n33456), .B(n33455), .Z(n33457) );
  AND U33916 ( .A(n33458), .B(n33457), .Z(n33544) );
  XNOR U33917 ( .A(n33545), .B(n33544), .Z(n33547) );
  NANDN U33918 ( .A(n33460), .B(n33459), .Z(n33464) );
  OR U33919 ( .A(n33462), .B(n33461), .Z(n33463) );
  AND U33920 ( .A(n33464), .B(n33463), .Z(n33546) );
  XOR U33921 ( .A(n33547), .B(n33546), .Z(n33539) );
  NANDN U33922 ( .A(n33466), .B(n33465), .Z(n33470) );
  NANDN U33923 ( .A(n33468), .B(n33467), .Z(n33469) );
  AND U33924 ( .A(n33470), .B(n33469), .Z(n33538) );
  XOR U33925 ( .A(n33539), .B(n33538), .Z(n33541) );
  XNOR U33926 ( .A(n33540), .B(n33541), .Z(n33712) );
  XOR U33927 ( .A(n33713), .B(n33712), .Z(n33707) );
  NANDN U33928 ( .A(n33472), .B(n33471), .Z(n33476) );
  NANDN U33929 ( .A(n33474), .B(n33473), .Z(n33475) );
  AND U33930 ( .A(n33476), .B(n33475), .Z(n33704) );
  NANDN U33931 ( .A(n33478), .B(n33477), .Z(n33482) );
  OR U33932 ( .A(n33480), .B(n33479), .Z(n33481) );
  AND U33933 ( .A(n33482), .B(n33481), .Z(n33689) );
  NANDN U33934 ( .A(n33483), .B(n35654), .Z(n33485) );
  XOR U33935 ( .A(a[116]), .B(b[33]), .Z(n33562) );
  NANDN U33936 ( .A(n35456), .B(n33562), .Z(n33484) );
  AND U33937 ( .A(n33485), .B(n33484), .Z(n33664) );
  NANDN U33938 ( .A(n34909), .B(n33486), .Z(n33488) );
  XOR U33939 ( .A(a[118]), .B(b[31]), .Z(n33565) );
  NANDN U33940 ( .A(n35145), .B(n33565), .Z(n33487) );
  AND U33941 ( .A(n33488), .B(n33487), .Z(n33663) );
  NANDN U33942 ( .A(n37974), .B(n33489), .Z(n33491) );
  XOR U33943 ( .A(b[57]), .B(a[92]), .Z(n33598) );
  NANDN U33944 ( .A(n38031), .B(n33598), .Z(n33490) );
  NAND U33945 ( .A(n33491), .B(n33490), .Z(n33662) );
  XOR U33946 ( .A(n33663), .B(n33662), .Z(n33665) );
  XOR U33947 ( .A(n33664), .B(n33665), .Z(n33687) );
  NANDN U33948 ( .A(n33493), .B(n33492), .Z(n33495) );
  XOR U33949 ( .A(a[126]), .B(b[23]), .Z(n33643) );
  NANDN U33950 ( .A(n33644), .B(n33643), .Z(n33494) );
  AND U33951 ( .A(n33495), .B(n33494), .Z(n33670) );
  NANDN U33952 ( .A(n38247), .B(n33496), .Z(n33498) );
  XOR U33953 ( .A(b[61]), .B(a[88]), .Z(n33647) );
  NANDN U33954 ( .A(n38248), .B(n33647), .Z(n33497) );
  AND U33955 ( .A(n33498), .B(n33497), .Z(n33669) );
  NANDN U33956 ( .A(n36742), .B(n33499), .Z(n33501) );
  XOR U33957 ( .A(b[43]), .B(a[106]), .Z(n33580) );
  NANDN U33958 ( .A(n36891), .B(n33580), .Z(n33500) );
  NAND U33959 ( .A(n33501), .B(n33500), .Z(n33668) );
  XOR U33960 ( .A(n33669), .B(n33668), .Z(n33671) );
  XNOR U33961 ( .A(n33670), .B(n33671), .Z(n33686) );
  XNOR U33962 ( .A(n33687), .B(n33686), .Z(n33688) );
  XOR U33963 ( .A(n33689), .B(n33688), .Z(n33694) );
  NANDN U33964 ( .A(n33503), .B(n33502), .Z(n33507) );
  OR U33965 ( .A(n33505), .B(n33504), .Z(n33506) );
  AND U33966 ( .A(n33507), .B(n33506), .Z(n33693) );
  NANDN U33967 ( .A(n33509), .B(n33508), .Z(n33513) );
  OR U33968 ( .A(n33511), .B(n33510), .Z(n33512) );
  NAND U33969 ( .A(n33513), .B(n33512), .Z(n33692) );
  XOR U33970 ( .A(n33693), .B(n33692), .Z(n33695) );
  XOR U33971 ( .A(n33694), .B(n33695), .Z(n33699) );
  XNOR U33972 ( .A(n33699), .B(n33698), .Z(n33700) );
  NANDN U33973 ( .A(n33519), .B(n33518), .Z(n33523) );
  OR U33974 ( .A(n33521), .B(n33520), .Z(n33522) );
  NAND U33975 ( .A(n33523), .B(n33522), .Z(n33701) );
  XOR U33976 ( .A(n33700), .B(n33701), .Z(n33705) );
  XNOR U33977 ( .A(n33704), .B(n33705), .Z(n33706) );
  XOR U33978 ( .A(n33707), .B(n33706), .Z(n33717) );
  XNOR U33979 ( .A(n33716), .B(n33717), .Z(n33718) );
  XOR U33980 ( .A(n33719), .B(n33718), .Z(n33533) );
  XNOR U33981 ( .A(n33532), .B(n33533), .Z(n33534) );
  XOR U33982 ( .A(n33535), .B(n33534), .Z(n33527) );
  XOR U33983 ( .A(n33526), .B(n33527), .Z(n33529) );
  XNOR U33984 ( .A(n33528), .B(n33529), .Z(n33524) );
  XOR U33985 ( .A(n33525), .B(n33524), .Z(c[212]) );
  AND U33986 ( .A(n33525), .B(n33524), .Z(n33729) );
  NANDN U33987 ( .A(n33527), .B(n33526), .Z(n33531) );
  OR U33988 ( .A(n33529), .B(n33528), .Z(n33530) );
  AND U33989 ( .A(n33531), .B(n33530), .Z(n33732) );
  NANDN U33990 ( .A(n33533), .B(n33532), .Z(n33537) );
  NANDN U33991 ( .A(n33535), .B(n33534), .Z(n33536) );
  AND U33992 ( .A(n33537), .B(n33536), .Z(n33731) );
  NANDN U33993 ( .A(n33539), .B(n33538), .Z(n33543) );
  NANDN U33994 ( .A(n33541), .B(n33540), .Z(n33542) );
  AND U33995 ( .A(n33543), .B(n33542), .Z(n33914) );
  NANDN U33996 ( .A(n33545), .B(n33544), .Z(n33549) );
  NAND U33997 ( .A(n33547), .B(n33546), .Z(n33548) );
  AND U33998 ( .A(n33549), .B(n33548), .Z(n33798) );
  NANDN U33999 ( .A(n212), .B(n33550), .Z(n33552) );
  XOR U34000 ( .A(b[49]), .B(a[101]), .Z(n33827) );
  NANDN U34001 ( .A(n37432), .B(n33827), .Z(n33551) );
  AND U34002 ( .A(n33552), .B(n33551), .Z(n33781) );
  NANDN U34003 ( .A(n37526), .B(n33553), .Z(n33555) );
  XOR U34004 ( .A(b[51]), .B(a[99]), .Z(n33887) );
  NANDN U34005 ( .A(n37605), .B(n33887), .Z(n33554) );
  AND U34006 ( .A(n33555), .B(n33554), .Z(n33780) );
  NANDN U34007 ( .A(n34634), .B(n33556), .Z(n33558) );
  XOR U34008 ( .A(a[121]), .B(b[29]), .Z(n33766) );
  NANDN U34009 ( .A(n34722), .B(n33766), .Z(n33557) );
  NAND U34010 ( .A(n33558), .B(n33557), .Z(n33779) );
  XOR U34011 ( .A(n33780), .B(n33779), .Z(n33782) );
  XOR U34012 ( .A(n33781), .B(n33782), .Z(n33788) );
  NANDN U34013 ( .A(n36210), .B(n33559), .Z(n33561) );
  XOR U34014 ( .A(a[111]), .B(b[39]), .Z(n33860) );
  NANDN U34015 ( .A(n36347), .B(n33860), .Z(n33560) );
  AND U34016 ( .A(n33561), .B(n33560), .Z(n33892) );
  NANDN U34017 ( .A(n35260), .B(n33562), .Z(n33564) );
  XOR U34018 ( .A(a[117]), .B(b[33]), .Z(n33833) );
  NANDN U34019 ( .A(n35456), .B(n33833), .Z(n33563) );
  AND U34020 ( .A(n33564), .B(n33563), .Z(n33891) );
  NANDN U34021 ( .A(n34909), .B(n33565), .Z(n33567) );
  XOR U34022 ( .A(a[119]), .B(b[31]), .Z(n33857) );
  NANDN U34023 ( .A(n35145), .B(n33857), .Z(n33566) );
  NAND U34024 ( .A(n33567), .B(n33566), .Z(n33890) );
  XOR U34025 ( .A(n33891), .B(n33890), .Z(n33893) );
  XOR U34026 ( .A(n33892), .B(n33893), .Z(n33786) );
  NAND U34027 ( .A(n36238), .B(n33568), .Z(n33570) );
  XNOR U34028 ( .A(a[113]), .B(b[37]), .Z(n33836) );
  NANDN U34029 ( .A(n33836), .B(n36239), .Z(n33569) );
  AND U34030 ( .A(n33570), .B(n33569), .Z(n33785) );
  XNOR U34031 ( .A(n33786), .B(n33785), .Z(n33787) );
  XNOR U34032 ( .A(n33788), .B(n33787), .Z(n33797) );
  XNOR U34033 ( .A(n33798), .B(n33797), .Z(n33799) );
  NANDN U34034 ( .A(n33572), .B(n33571), .Z(n33576) );
  NANDN U34035 ( .A(n33574), .B(n33573), .Z(n33575) );
  AND U34036 ( .A(n33576), .B(n33575), .Z(n33898) );
  NANDN U34037 ( .A(n38278), .B(n33577), .Z(n33579) );
  XOR U34038 ( .A(b[63]), .B(a[87]), .Z(n33863) );
  NANDN U34039 ( .A(n38279), .B(n33863), .Z(n33578) );
  AND U34040 ( .A(n33579), .B(n33578), .Z(n33816) );
  NANDN U34041 ( .A(n36742), .B(n33580), .Z(n33582) );
  XOR U34042 ( .A(b[43]), .B(a[107]), .Z(n33839) );
  NANDN U34043 ( .A(n36891), .B(n33839), .Z(n33581) );
  NAND U34044 ( .A(n33582), .B(n33581), .Z(n33815) );
  XNOR U34045 ( .A(n33816), .B(n33815), .Z(n33818) );
  IV U34046 ( .A(n33778), .Z(n33584) );
  AND U34047 ( .A(b[63]), .B(a[85]), .Z(n33776) );
  XOR U34048 ( .A(n33775), .B(n33776), .Z(n33777) );
  XOR U34049 ( .A(n33584), .B(n33777), .Z(n33817) );
  XOR U34050 ( .A(n33818), .B(n33817), .Z(n33897) );
  NANDN U34051 ( .A(n33584), .B(n33583), .Z(n33588) );
  NANDN U34052 ( .A(n33586), .B(n33585), .Z(n33587) );
  AND U34053 ( .A(n33588), .B(n33587), .Z(n33896) );
  XOR U34054 ( .A(n33897), .B(n33896), .Z(n33899) );
  XOR U34055 ( .A(n33898), .B(n33899), .Z(n33800) );
  XOR U34056 ( .A(n33799), .B(n33800), .Z(n33915) );
  XNOR U34057 ( .A(n33914), .B(n33915), .Z(n33917) );
  NANDN U34058 ( .A(n33590), .B(n33589), .Z(n33594) );
  NANDN U34059 ( .A(n33592), .B(n33591), .Z(n33593) );
  AND U34060 ( .A(n33594), .B(n33593), .Z(n33916) );
  XOR U34061 ( .A(n33917), .B(n33916), .Z(n33928) );
  NANDN U34062 ( .A(n37857), .B(n33595), .Z(n33597) );
  XOR U34063 ( .A(b[55]), .B(a[95]), .Z(n33854) );
  NANDN U34064 ( .A(n37911), .B(n33854), .Z(n33596) );
  AND U34065 ( .A(n33597), .B(n33596), .Z(n33823) );
  NANDN U34066 ( .A(n37974), .B(n33598), .Z(n33600) );
  XOR U34067 ( .A(b[57]), .B(a[93]), .Z(n33881) );
  NANDN U34068 ( .A(n38031), .B(n33881), .Z(n33599) );
  AND U34069 ( .A(n33600), .B(n33599), .Z(n33822) );
  NANDN U34070 ( .A(n36480), .B(n33601), .Z(n33603) );
  XOR U34071 ( .A(a[109]), .B(b[41]), .Z(n33845) );
  NANDN U34072 ( .A(n36594), .B(n33845), .Z(n33602) );
  NAND U34073 ( .A(n33603), .B(n33602), .Z(n33821) );
  XOR U34074 ( .A(n33822), .B(n33821), .Z(n33824) );
  XOR U34075 ( .A(n33823), .B(n33824), .Z(n33903) );
  NANDN U34076 ( .A(n35611), .B(n33604), .Z(n33606) );
  XOR U34077 ( .A(a[115]), .B(b[35]), .Z(n33842) );
  NANDN U34078 ( .A(n35801), .B(n33842), .Z(n33605) );
  AND U34079 ( .A(n33606), .B(n33605), .Z(n33850) );
  NANDN U34080 ( .A(n37705), .B(n33607), .Z(n33609) );
  XOR U34081 ( .A(b[53]), .B(a[97]), .Z(n33830) );
  NANDN U34082 ( .A(n37778), .B(n33830), .Z(n33608) );
  AND U34083 ( .A(n33609), .B(n33608), .Z(n33849) );
  NANDN U34084 ( .A(n34223), .B(n33610), .Z(n33612) );
  XOR U34085 ( .A(a[123]), .B(b[27]), .Z(n33769) );
  NANDN U34086 ( .A(n34458), .B(n33769), .Z(n33611) );
  NAND U34087 ( .A(n33612), .B(n33611), .Z(n33848) );
  XOR U34088 ( .A(n33849), .B(n33848), .Z(n33851) );
  XNOR U34089 ( .A(n33850), .B(n33851), .Z(n33902) );
  XNOR U34090 ( .A(n33903), .B(n33902), .Z(n33904) );
  NANDN U34091 ( .A(n33614), .B(n33613), .Z(n33618) );
  OR U34092 ( .A(n33616), .B(n33615), .Z(n33617) );
  NAND U34093 ( .A(n33618), .B(n33617), .Z(n33905) );
  XNOR U34094 ( .A(n33904), .B(n33905), .Z(n33809) );
  NANDN U34095 ( .A(n33620), .B(n33619), .Z(n33624) );
  OR U34096 ( .A(n33622), .B(n33621), .Z(n33623) );
  NAND U34097 ( .A(n33624), .B(n33623), .Z(n33810) );
  XNOR U34098 ( .A(n33809), .B(n33810), .Z(n33812) );
  NANDN U34099 ( .A(n33626), .B(n33625), .Z(n33630) );
  NANDN U34100 ( .A(n33628), .B(n33627), .Z(n33629) );
  AND U34101 ( .A(n33630), .B(n33629), .Z(n33811) );
  XOR U34102 ( .A(n33812), .B(n33811), .Z(n33805) );
  NANDN U34103 ( .A(n33632), .B(n33631), .Z(n33636) );
  NANDN U34104 ( .A(n33634), .B(n33633), .Z(n33635) );
  AND U34105 ( .A(n33636), .B(n33635), .Z(n33804) );
  NANDN U34106 ( .A(n33638), .B(n33637), .Z(n33642) );
  OR U34107 ( .A(n33640), .B(n33639), .Z(n33641) );
  AND U34108 ( .A(n33642), .B(n33641), .Z(n33911) );
  NANDN U34109 ( .A(n33866), .B(n33643), .Z(n33646) );
  XOR U34110 ( .A(a[127]), .B(b[23]), .Z(n33867) );
  NANDN U34111 ( .A(n33644), .B(n33867), .Z(n33645) );
  AND U34112 ( .A(n33646), .B(n33645), .Z(n33763) );
  NANDN U34113 ( .A(n38247), .B(n33647), .Z(n33649) );
  XOR U34114 ( .A(b[61]), .B(a[89]), .Z(n33871) );
  NANDN U34115 ( .A(n38248), .B(n33871), .Z(n33648) );
  AND U34116 ( .A(n33649), .B(n33648), .Z(n33761) );
  NANDN U34117 ( .A(n36991), .B(n33650), .Z(n33652) );
  XOR U34118 ( .A(b[45]), .B(a[105]), .Z(n33878) );
  NANDN U34119 ( .A(n37083), .B(n33878), .Z(n33651) );
  NAND U34120 ( .A(n33652), .B(n33651), .Z(n33760) );
  XNOR U34121 ( .A(n33761), .B(n33760), .Z(n33762) );
  XOR U34122 ( .A(n33763), .B(n33762), .Z(n33909) );
  NANDN U34123 ( .A(n38090), .B(n33653), .Z(n33655) );
  XOR U34124 ( .A(b[59]), .B(a[91]), .Z(n33884) );
  NANDN U34125 ( .A(n38130), .B(n33884), .Z(n33654) );
  AND U34126 ( .A(n33655), .B(n33654), .Z(n33756) );
  NANDN U34127 ( .A(n33875), .B(n33656), .Z(n33658) );
  XOR U34128 ( .A(a[125]), .B(b[25]), .Z(n33874) );
  NANDN U34129 ( .A(n33994), .B(n33874), .Z(n33657) );
  AND U34130 ( .A(n33658), .B(n33657), .Z(n33755) );
  NANDN U34131 ( .A(n211), .B(n33659), .Z(n33661) );
  XOR U34132 ( .A(b[47]), .B(a[103]), .Z(n33772) );
  NANDN U34133 ( .A(n37172), .B(n33772), .Z(n33660) );
  NAND U34134 ( .A(n33661), .B(n33660), .Z(n33754) );
  XOR U34135 ( .A(n33755), .B(n33754), .Z(n33757) );
  XNOR U34136 ( .A(n33756), .B(n33757), .Z(n33908) );
  XOR U34137 ( .A(n33909), .B(n33908), .Z(n33910) );
  XOR U34138 ( .A(n33911), .B(n33910), .Z(n33794) );
  NANDN U34139 ( .A(n33663), .B(n33662), .Z(n33667) );
  OR U34140 ( .A(n33665), .B(n33664), .Z(n33666) );
  AND U34141 ( .A(n33667), .B(n33666), .Z(n33792) );
  NANDN U34142 ( .A(n33669), .B(n33668), .Z(n33673) );
  OR U34143 ( .A(n33671), .B(n33670), .Z(n33672) );
  NAND U34144 ( .A(n33673), .B(n33672), .Z(n33791) );
  XNOR U34145 ( .A(n33792), .B(n33791), .Z(n33793) );
  XNOR U34146 ( .A(n33794), .B(n33793), .Z(n33803) );
  XOR U34147 ( .A(n33804), .B(n33803), .Z(n33806) );
  XOR U34148 ( .A(n33805), .B(n33806), .Z(n33922) );
  NAND U34149 ( .A(n33675), .B(n33674), .Z(n33679) );
  NAND U34150 ( .A(n33677), .B(n33676), .Z(n33678) );
  AND U34151 ( .A(n33679), .B(n33678), .Z(n33921) );
  NANDN U34152 ( .A(n33681), .B(n33680), .Z(n33685) );
  NANDN U34153 ( .A(n33683), .B(n33682), .Z(n33684) );
  AND U34154 ( .A(n33685), .B(n33684), .Z(n33749) );
  NANDN U34155 ( .A(n33687), .B(n33686), .Z(n33691) );
  NAND U34156 ( .A(n33689), .B(n33688), .Z(n33690) );
  NAND U34157 ( .A(n33691), .B(n33690), .Z(n33748) );
  XNOR U34158 ( .A(n33749), .B(n33748), .Z(n33750) );
  NANDN U34159 ( .A(n33693), .B(n33692), .Z(n33697) );
  OR U34160 ( .A(n33695), .B(n33694), .Z(n33696) );
  NAND U34161 ( .A(n33697), .B(n33696), .Z(n33751) );
  XNOR U34162 ( .A(n33750), .B(n33751), .Z(n33920) );
  XOR U34163 ( .A(n33921), .B(n33920), .Z(n33923) );
  XOR U34164 ( .A(n33922), .B(n33923), .Z(n33927) );
  NANDN U34165 ( .A(n33699), .B(n33698), .Z(n33703) );
  NANDN U34166 ( .A(n33701), .B(n33700), .Z(n33702) );
  AND U34167 ( .A(n33703), .B(n33702), .Z(n33926) );
  XOR U34168 ( .A(n33927), .B(n33926), .Z(n33929) );
  XOR U34169 ( .A(n33928), .B(n33929), .Z(n33745) );
  NANDN U34170 ( .A(n33705), .B(n33704), .Z(n33709) );
  NANDN U34171 ( .A(n33707), .B(n33706), .Z(n33708) );
  AND U34172 ( .A(n33709), .B(n33708), .Z(n33743) );
  NANDN U34173 ( .A(n33711), .B(n33710), .Z(n33715) );
  NAND U34174 ( .A(n33713), .B(n33712), .Z(n33714) );
  AND U34175 ( .A(n33715), .B(n33714), .Z(n33742) );
  XNOR U34176 ( .A(n33743), .B(n33742), .Z(n33744) );
  XNOR U34177 ( .A(n33745), .B(n33744), .Z(n33738) );
  NANDN U34178 ( .A(n33717), .B(n33716), .Z(n33721) );
  NANDN U34179 ( .A(n33719), .B(n33718), .Z(n33720) );
  AND U34180 ( .A(n33721), .B(n33720), .Z(n33737) );
  NANDN U34181 ( .A(n33723), .B(n33722), .Z(n33727) );
  NAND U34182 ( .A(n33725), .B(n33724), .Z(n33726) );
  AND U34183 ( .A(n33727), .B(n33726), .Z(n33736) );
  XOR U34184 ( .A(n33737), .B(n33736), .Z(n33739) );
  XNOR U34185 ( .A(n33738), .B(n33739), .Z(n33730) );
  XOR U34186 ( .A(n33731), .B(n33730), .Z(n33733) );
  XNOR U34187 ( .A(n33732), .B(n33733), .Z(n33728) );
  XOR U34188 ( .A(n33729), .B(n33728), .Z(c[213]) );
  AND U34189 ( .A(n33729), .B(n33728), .Z(n33933) );
  NANDN U34190 ( .A(n33731), .B(n33730), .Z(n33735) );
  OR U34191 ( .A(n33733), .B(n33732), .Z(n33734) );
  AND U34192 ( .A(n33735), .B(n33734), .Z(n33936) );
  NANDN U34193 ( .A(n33737), .B(n33736), .Z(n33741) );
  NANDN U34194 ( .A(n33739), .B(n33738), .Z(n33740) );
  AND U34195 ( .A(n33741), .B(n33740), .Z(n33935) );
  NANDN U34196 ( .A(n33743), .B(n33742), .Z(n33747) );
  NANDN U34197 ( .A(n33745), .B(n33744), .Z(n33746) );
  AND U34198 ( .A(n33747), .B(n33746), .Z(n34121) );
  NANDN U34199 ( .A(n33749), .B(n33748), .Z(n33753) );
  NANDN U34200 ( .A(n33751), .B(n33750), .Z(n33752) );
  AND U34201 ( .A(n33753), .B(n33752), .Z(n33955) );
  NANDN U34202 ( .A(n33755), .B(n33754), .Z(n33759) );
  OR U34203 ( .A(n33757), .B(n33756), .Z(n33758) );
  AND U34204 ( .A(n33759), .B(n33758), .Z(n34017) );
  NANDN U34205 ( .A(n33761), .B(n33760), .Z(n33765) );
  NANDN U34206 ( .A(n33763), .B(n33762), .Z(n33764) );
  NAND U34207 ( .A(n33765), .B(n33764), .Z(n34016) );
  XNOR U34208 ( .A(n34017), .B(n34016), .Z(n34019) );
  NANDN U34209 ( .A(n34634), .B(n33766), .Z(n33768) );
  XOR U34210 ( .A(a[122]), .B(b[29]), .Z(n34043) );
  NANDN U34211 ( .A(n34722), .B(n34043), .Z(n33767) );
  AND U34212 ( .A(n33768), .B(n33767), .Z(n33979) );
  NANDN U34213 ( .A(n34223), .B(n33769), .Z(n33771) );
  XOR U34214 ( .A(a[124]), .B(b[27]), .Z(n34064) );
  NANDN U34215 ( .A(n34458), .B(n34064), .Z(n33770) );
  AND U34216 ( .A(n33771), .B(n33770), .Z(n33977) );
  NANDN U34217 ( .A(n211), .B(n33772), .Z(n33774) );
  XOR U34218 ( .A(b[47]), .B(a[104]), .Z(n34046) );
  NANDN U34219 ( .A(n37172), .B(n34046), .Z(n33773) );
  NAND U34220 ( .A(n33774), .B(n33773), .Z(n33976) );
  XNOR U34221 ( .A(n33977), .B(n33976), .Z(n33978) );
  XNOR U34222 ( .A(n33979), .B(n33978), .Z(n34095) );
  XOR U34223 ( .A(n34095), .B(n34094), .Z(n34097) );
  NANDN U34224 ( .A(n33780), .B(n33779), .Z(n33784) );
  OR U34225 ( .A(n33782), .B(n33781), .Z(n33783) );
  NAND U34226 ( .A(n33784), .B(n33783), .Z(n34096) );
  XOR U34227 ( .A(n34097), .B(n34096), .Z(n34018) );
  XOR U34228 ( .A(n34019), .B(n34018), .Z(n33965) );
  NANDN U34229 ( .A(n33786), .B(n33785), .Z(n33790) );
  NANDN U34230 ( .A(n33788), .B(n33787), .Z(n33789) );
  NAND U34231 ( .A(n33790), .B(n33789), .Z(n33964) );
  XNOR U34232 ( .A(n33965), .B(n33964), .Z(n33967) );
  NANDN U34233 ( .A(n33792), .B(n33791), .Z(n33796) );
  NANDN U34234 ( .A(n33794), .B(n33793), .Z(n33795) );
  AND U34235 ( .A(n33796), .B(n33795), .Z(n33966) );
  XOR U34236 ( .A(n33967), .B(n33966), .Z(n33953) );
  NANDN U34237 ( .A(n33798), .B(n33797), .Z(n33802) );
  NANDN U34238 ( .A(n33800), .B(n33799), .Z(n33801) );
  AND U34239 ( .A(n33802), .B(n33801), .Z(n33952) );
  XNOR U34240 ( .A(n33953), .B(n33952), .Z(n33954) );
  XOR U34241 ( .A(n33955), .B(n33954), .Z(n33948) );
  NANDN U34242 ( .A(n33804), .B(n33803), .Z(n33808) );
  OR U34243 ( .A(n33806), .B(n33805), .Z(n33807) );
  AND U34244 ( .A(n33808), .B(n33807), .Z(n33946) );
  NANDN U34245 ( .A(n33810), .B(n33809), .Z(n33814) );
  NAND U34246 ( .A(n33812), .B(n33811), .Z(n33813) );
  AND U34247 ( .A(n33814), .B(n33813), .Z(n33961) );
  NANDN U34248 ( .A(n33816), .B(n33815), .Z(n33820) );
  NAND U34249 ( .A(n33818), .B(n33817), .Z(n33819) );
  AND U34250 ( .A(n33820), .B(n33819), .Z(n34101) );
  NANDN U34251 ( .A(n33822), .B(n33821), .Z(n33826) );
  OR U34252 ( .A(n33824), .B(n33823), .Z(n33825) );
  NAND U34253 ( .A(n33826), .B(n33825), .Z(n34100) );
  XNOR U34254 ( .A(n34101), .B(n34100), .Z(n34103) );
  NANDN U34255 ( .A(n212), .B(n33827), .Z(n33829) );
  XOR U34256 ( .A(b[49]), .B(a[102]), .Z(n34070) );
  NANDN U34257 ( .A(n37432), .B(n34070), .Z(n33828) );
  AND U34258 ( .A(n33829), .B(n33828), .Z(n34084) );
  NANDN U34259 ( .A(n37705), .B(n33830), .Z(n33832) );
  XOR U34260 ( .A(b[53]), .B(a[98]), .Z(n34055) );
  NANDN U34261 ( .A(n37778), .B(n34055), .Z(n33831) );
  AND U34262 ( .A(n33832), .B(n33831), .Z(n34083) );
  NANDN U34263 ( .A(n35260), .B(n33833), .Z(n33835) );
  XOR U34264 ( .A(a[118]), .B(b[33]), .Z(n34052) );
  NANDN U34265 ( .A(n35456), .B(n34052), .Z(n33834) );
  NAND U34266 ( .A(n33835), .B(n33834), .Z(n34082) );
  XOR U34267 ( .A(n34083), .B(n34082), .Z(n34085) );
  XOR U34268 ( .A(n34084), .B(n34085), .Z(n34012) );
  NANDN U34269 ( .A(n33836), .B(n36238), .Z(n33838) );
  XOR U34270 ( .A(a[114]), .B(b[37]), .Z(n34028) );
  NANDN U34271 ( .A(n36047), .B(n34028), .Z(n33837) );
  AND U34272 ( .A(n33838), .B(n33837), .Z(n34036) );
  NANDN U34273 ( .A(n36742), .B(n33839), .Z(n33841) );
  XOR U34274 ( .A(b[43]), .B(a[108]), .Z(n34007) );
  NANDN U34275 ( .A(n36891), .B(n34007), .Z(n33840) );
  AND U34276 ( .A(n33841), .B(n33840), .Z(n34035) );
  NANDN U34277 ( .A(n35611), .B(n33842), .Z(n33844) );
  XOR U34278 ( .A(a[116]), .B(b[35]), .Z(n34049) );
  NANDN U34279 ( .A(n35801), .B(n34049), .Z(n33843) );
  NAND U34280 ( .A(n33844), .B(n33843), .Z(n34034) );
  XOR U34281 ( .A(n34035), .B(n34034), .Z(n34037) );
  XOR U34282 ( .A(n34036), .B(n34037), .Z(n34011) );
  NAND U34283 ( .A(n36735), .B(n33845), .Z(n33847) );
  XNOR U34284 ( .A(a[110]), .B(b[41]), .Z(n34001) );
  NANDN U34285 ( .A(n34001), .B(n36733), .Z(n33846) );
  AND U34286 ( .A(n33847), .B(n33846), .Z(n34010) );
  XOR U34287 ( .A(n34011), .B(n34010), .Z(n34013) );
  XNOR U34288 ( .A(n34012), .B(n34013), .Z(n34102) );
  XOR U34289 ( .A(n34103), .B(n34102), .Z(n33973) );
  NANDN U34290 ( .A(n33849), .B(n33848), .Z(n33853) );
  OR U34291 ( .A(n33851), .B(n33850), .Z(n33852) );
  AND U34292 ( .A(n33853), .B(n33852), .Z(n34108) );
  NANDN U34293 ( .A(n37857), .B(n33854), .Z(n33856) );
  XOR U34294 ( .A(b[55]), .B(a[96]), .Z(n34022) );
  NANDN U34295 ( .A(n37911), .B(n34022), .Z(n33855) );
  AND U34296 ( .A(n33856), .B(n33855), .Z(n33990) );
  NANDN U34297 ( .A(n34909), .B(n33857), .Z(n33859) );
  XOR U34298 ( .A(a[120]), .B(b[31]), .Z(n34040) );
  NANDN U34299 ( .A(n35145), .B(n34040), .Z(n33858) );
  AND U34300 ( .A(n33859), .B(n33858), .Z(n33989) );
  NANDN U34301 ( .A(n36210), .B(n33860), .Z(n33862) );
  XOR U34302 ( .A(a[112]), .B(b[39]), .Z(n34004) );
  NANDN U34303 ( .A(n36347), .B(n34004), .Z(n33861) );
  NAND U34304 ( .A(n33862), .B(n33861), .Z(n33988) );
  XOR U34305 ( .A(n33989), .B(n33988), .Z(n33991) );
  XOR U34306 ( .A(n33990), .B(n33991), .Z(n34107) );
  NANDN U34307 ( .A(n38278), .B(n33863), .Z(n33865) );
  XOR U34308 ( .A(b[63]), .B(a[88]), .Z(n34067) );
  NANDN U34309 ( .A(n38279), .B(n34067), .Z(n33864) );
  AND U34310 ( .A(n33865), .B(n33864), .Z(n34033) );
  NAND U34311 ( .A(b[63]), .B(a[86]), .Z(n34266) );
  ANDN U34312 ( .B(n33867), .A(n33866), .Z(n33870) );
  NAND U34313 ( .A(b[23]), .B(n33868), .Z(n33869) );
  NANDN U34314 ( .A(n33870), .B(n33869), .Z(n34031) );
  XOR U34315 ( .A(n34266), .B(n34031), .Z(n34032) );
  XOR U34316 ( .A(n34033), .B(n34032), .Z(n34106) );
  XOR U34317 ( .A(n34107), .B(n34106), .Z(n34109) );
  XNOR U34318 ( .A(n34108), .B(n34109), .Z(n33970) );
  NANDN U34319 ( .A(n38247), .B(n33871), .Z(n33873) );
  XOR U34320 ( .A(b[61]), .B(a[90]), .Z(n34076) );
  NANDN U34321 ( .A(n38248), .B(n34076), .Z(n33872) );
  AND U34322 ( .A(n33873), .B(n33872), .Z(n33984) );
  NANDN U34323 ( .A(n33875), .B(n33874), .Z(n33877) );
  XOR U34324 ( .A(a[126]), .B(b[25]), .Z(n33995) );
  NANDN U34325 ( .A(n33994), .B(n33995), .Z(n33876) );
  AND U34326 ( .A(n33877), .B(n33876), .Z(n33983) );
  NANDN U34327 ( .A(n36991), .B(n33878), .Z(n33880) );
  XOR U34328 ( .A(b[45]), .B(a[106]), .Z(n33998) );
  NANDN U34329 ( .A(n37083), .B(n33998), .Z(n33879) );
  NAND U34330 ( .A(n33880), .B(n33879), .Z(n33982) );
  XOR U34331 ( .A(n33983), .B(n33982), .Z(n33985) );
  XOR U34332 ( .A(n33984), .B(n33985), .Z(n34089) );
  NANDN U34333 ( .A(n37974), .B(n33881), .Z(n33883) );
  XOR U34334 ( .A(b[57]), .B(a[94]), .Z(n34025) );
  NANDN U34335 ( .A(n38031), .B(n34025), .Z(n33882) );
  AND U34336 ( .A(n33883), .B(n33882), .Z(n34060) );
  NANDN U34337 ( .A(n38090), .B(n33884), .Z(n33886) );
  XOR U34338 ( .A(b[59]), .B(a[92]), .Z(n34073) );
  NANDN U34339 ( .A(n38130), .B(n34073), .Z(n33885) );
  AND U34340 ( .A(n33886), .B(n33885), .Z(n34059) );
  NANDN U34341 ( .A(n37526), .B(n33887), .Z(n33889) );
  XOR U34342 ( .A(b[51]), .B(a[100]), .Z(n34079) );
  NANDN U34343 ( .A(n37605), .B(n34079), .Z(n33888) );
  NAND U34344 ( .A(n33889), .B(n33888), .Z(n34058) );
  XOR U34345 ( .A(n34059), .B(n34058), .Z(n34061) );
  XNOR U34346 ( .A(n34060), .B(n34061), .Z(n34088) );
  XNOR U34347 ( .A(n34089), .B(n34088), .Z(n34090) );
  NANDN U34348 ( .A(n33891), .B(n33890), .Z(n33895) );
  OR U34349 ( .A(n33893), .B(n33892), .Z(n33894) );
  NAND U34350 ( .A(n33895), .B(n33894), .Z(n34091) );
  XOR U34351 ( .A(n34090), .B(n34091), .Z(n33971) );
  XNOR U34352 ( .A(n33970), .B(n33971), .Z(n33972) );
  XNOR U34353 ( .A(n33973), .B(n33972), .Z(n33958) );
  NANDN U34354 ( .A(n33897), .B(n33896), .Z(n33901) );
  NANDN U34355 ( .A(n33899), .B(n33898), .Z(n33900) );
  AND U34356 ( .A(n33901), .B(n33900), .Z(n34115) );
  NANDN U34357 ( .A(n33903), .B(n33902), .Z(n33907) );
  NANDN U34358 ( .A(n33905), .B(n33904), .Z(n33906) );
  AND U34359 ( .A(n33907), .B(n33906), .Z(n34113) );
  NAND U34360 ( .A(n33909), .B(n33908), .Z(n33913) );
  NAND U34361 ( .A(n33911), .B(n33910), .Z(n33912) );
  NAND U34362 ( .A(n33913), .B(n33912), .Z(n34112) );
  XNOR U34363 ( .A(n34113), .B(n34112), .Z(n34114) );
  XOR U34364 ( .A(n34115), .B(n34114), .Z(n33959) );
  XNOR U34365 ( .A(n33958), .B(n33959), .Z(n33960) );
  XOR U34366 ( .A(n33961), .B(n33960), .Z(n33947) );
  XOR U34367 ( .A(n33946), .B(n33947), .Z(n33949) );
  XOR U34368 ( .A(n33948), .B(n33949), .Z(n33942) );
  NANDN U34369 ( .A(n33915), .B(n33914), .Z(n33919) );
  NAND U34370 ( .A(n33917), .B(n33916), .Z(n33918) );
  AND U34371 ( .A(n33919), .B(n33918), .Z(n33940) );
  NANDN U34372 ( .A(n33921), .B(n33920), .Z(n33925) );
  OR U34373 ( .A(n33923), .B(n33922), .Z(n33924) );
  NAND U34374 ( .A(n33925), .B(n33924), .Z(n33941) );
  XOR U34375 ( .A(n33940), .B(n33941), .Z(n33943) );
  XOR U34376 ( .A(n33942), .B(n33943), .Z(n34119) );
  NANDN U34377 ( .A(n33927), .B(n33926), .Z(n33931) );
  OR U34378 ( .A(n33929), .B(n33928), .Z(n33930) );
  AND U34379 ( .A(n33931), .B(n33930), .Z(n34118) );
  XNOR U34380 ( .A(n34119), .B(n34118), .Z(n34120) );
  XNOR U34381 ( .A(n34121), .B(n34120), .Z(n33934) );
  XOR U34382 ( .A(n33935), .B(n33934), .Z(n33937) );
  XNOR U34383 ( .A(n33936), .B(n33937), .Z(n33932) );
  XOR U34384 ( .A(n33933), .B(n33932), .Z(c[214]) );
  AND U34385 ( .A(n33933), .B(n33932), .Z(n34125) );
  NANDN U34386 ( .A(n33935), .B(n33934), .Z(n33939) );
  OR U34387 ( .A(n33937), .B(n33936), .Z(n33938) );
  AND U34388 ( .A(n33939), .B(n33938), .Z(n34128) );
  NANDN U34389 ( .A(n33941), .B(n33940), .Z(n33945) );
  OR U34390 ( .A(n33943), .B(n33942), .Z(n33944) );
  AND U34391 ( .A(n33945), .B(n33944), .Z(n34134) );
  NANDN U34392 ( .A(n33947), .B(n33946), .Z(n33951) );
  OR U34393 ( .A(n33949), .B(n33948), .Z(n33950) );
  AND U34394 ( .A(n33951), .B(n33950), .Z(n34132) );
  NANDN U34395 ( .A(n33953), .B(n33952), .Z(n33957) );
  NAND U34396 ( .A(n33955), .B(n33954), .Z(n33956) );
  AND U34397 ( .A(n33957), .B(n33956), .Z(n34141) );
  NANDN U34398 ( .A(n33959), .B(n33958), .Z(n33963) );
  NANDN U34399 ( .A(n33961), .B(n33960), .Z(n33962) );
  AND U34400 ( .A(n33963), .B(n33962), .Z(n34138) );
  NANDN U34401 ( .A(n33965), .B(n33964), .Z(n33969) );
  NAND U34402 ( .A(n33967), .B(n33966), .Z(n33968) );
  AND U34403 ( .A(n33969), .B(n33968), .Z(n34309) );
  NANDN U34404 ( .A(n33971), .B(n33970), .Z(n33975) );
  NANDN U34405 ( .A(n33973), .B(n33972), .Z(n33974) );
  AND U34406 ( .A(n33975), .B(n33974), .Z(n34308) );
  NANDN U34407 ( .A(n33977), .B(n33976), .Z(n33981) );
  NANDN U34408 ( .A(n33979), .B(n33978), .Z(n33980) );
  AND U34409 ( .A(n33981), .B(n33980), .Z(n34157) );
  NANDN U34410 ( .A(n33983), .B(n33982), .Z(n33987) );
  OR U34411 ( .A(n33985), .B(n33984), .Z(n33986) );
  NAND U34412 ( .A(n33987), .B(n33986), .Z(n34156) );
  XNOR U34413 ( .A(n34157), .B(n34156), .Z(n34159) );
  NANDN U34414 ( .A(n33989), .B(n33988), .Z(n33993) );
  OR U34415 ( .A(n33991), .B(n33990), .Z(n33992) );
  AND U34416 ( .A(n33993), .B(n33992), .Z(n34304) );
  XNOR U34417 ( .A(a[127]), .B(b[25]), .Z(n34296) );
  OR U34418 ( .A(n34296), .B(n33994), .Z(n33997) );
  NAND U34419 ( .A(n34297), .B(n33995), .Z(n33996) );
  AND U34420 ( .A(n33997), .B(n33996), .Z(n34254) );
  NANDN U34421 ( .A(n36991), .B(n33998), .Z(n34000) );
  XOR U34422 ( .A(b[45]), .B(a[107]), .Z(n34195) );
  NANDN U34423 ( .A(n37083), .B(n34195), .Z(n33999) );
  NAND U34424 ( .A(n34000), .B(n33999), .Z(n34253) );
  XNOR U34425 ( .A(n34254), .B(n34253), .Z(n34256) );
  XOR U34426 ( .A(n34266), .B(n34267), .Z(n34269) );
  AND U34427 ( .A(b[63]), .B(a[87]), .Z(n34268) );
  XOR U34428 ( .A(n34269), .B(n34268), .Z(n34255) );
  XOR U34429 ( .A(n34256), .B(n34255), .Z(n34301) );
  NANDN U34430 ( .A(n34001), .B(n36735), .Z(n34003) );
  XOR U34431 ( .A(a[111]), .B(b[41]), .Z(n34260) );
  NANDN U34432 ( .A(n36594), .B(n34260), .Z(n34002) );
  AND U34433 ( .A(n34003), .B(n34002), .Z(n34275) );
  NANDN U34434 ( .A(n36210), .B(n34004), .Z(n34006) );
  XOR U34435 ( .A(a[113]), .B(b[39]), .Z(n34263) );
  NANDN U34436 ( .A(n36347), .B(n34263), .Z(n34005) );
  AND U34437 ( .A(n34006), .B(n34005), .Z(n34273) );
  NANDN U34438 ( .A(n36742), .B(n34007), .Z(n34009) );
  XOR U34439 ( .A(b[43]), .B(a[109]), .Z(n34257) );
  NANDN U34440 ( .A(n36891), .B(n34257), .Z(n34008) );
  NAND U34441 ( .A(n34009), .B(n34008), .Z(n34272) );
  XNOR U34442 ( .A(n34273), .B(n34272), .Z(n34274) );
  XOR U34443 ( .A(n34275), .B(n34274), .Z(n34302) );
  XNOR U34444 ( .A(n34301), .B(n34302), .Z(n34303) );
  XNOR U34445 ( .A(n34304), .B(n34303), .Z(n34158) );
  XOR U34446 ( .A(n34159), .B(n34158), .Z(n34175) );
  NANDN U34447 ( .A(n34011), .B(n34010), .Z(n34015) );
  OR U34448 ( .A(n34013), .B(n34012), .Z(n34014) );
  NAND U34449 ( .A(n34015), .B(n34014), .Z(n34174) );
  XNOR U34450 ( .A(n34175), .B(n34174), .Z(n34176) );
  NANDN U34451 ( .A(n34017), .B(n34016), .Z(n34021) );
  NAND U34452 ( .A(n34019), .B(n34018), .Z(n34020) );
  NAND U34453 ( .A(n34021), .B(n34020), .Z(n34177) );
  XNOR U34454 ( .A(n34176), .B(n34177), .Z(n34307) );
  XOR U34455 ( .A(n34308), .B(n34307), .Z(n34310) );
  XOR U34456 ( .A(n34309), .B(n34310), .Z(n34147) );
  NANDN U34457 ( .A(n37857), .B(n34022), .Z(n34024) );
  XOR U34458 ( .A(b[55]), .B(a[97]), .Z(n34213) );
  NANDN U34459 ( .A(n37911), .B(n34213), .Z(n34023) );
  AND U34460 ( .A(n34024), .B(n34023), .Z(n34231) );
  NANDN U34461 ( .A(n37974), .B(n34025), .Z(n34027) );
  XOR U34462 ( .A(b[57]), .B(a[95]), .Z(n34189) );
  NANDN U34463 ( .A(n38031), .B(n34189), .Z(n34026) );
  AND U34464 ( .A(n34027), .B(n34026), .Z(n34230) );
  NANDN U34465 ( .A(n35936), .B(n34028), .Z(n34030) );
  XOR U34466 ( .A(a[115]), .B(b[37]), .Z(n34216) );
  NANDN U34467 ( .A(n36047), .B(n34216), .Z(n34029) );
  NAND U34468 ( .A(n34030), .B(n34029), .Z(n34229) );
  XOR U34469 ( .A(n34230), .B(n34229), .Z(n34232) );
  XOR U34470 ( .A(n34231), .B(n34232), .Z(n34163) );
  XNOR U34471 ( .A(n34163), .B(n34162), .Z(n34165) );
  NANDN U34472 ( .A(n34035), .B(n34034), .Z(n34039) );
  OR U34473 ( .A(n34037), .B(n34036), .Z(n34038) );
  AND U34474 ( .A(n34039), .B(n34038), .Z(n34164) );
  XOR U34475 ( .A(n34165), .B(n34164), .Z(n34152) );
  NANDN U34476 ( .A(n34909), .B(n34040), .Z(n34042) );
  XOR U34477 ( .A(a[121]), .B(b[31]), .Z(n34284) );
  NANDN U34478 ( .A(n35145), .B(n34284), .Z(n34041) );
  AND U34479 ( .A(n34042), .B(n34041), .Z(n34249) );
  NANDN U34480 ( .A(n34634), .B(n34043), .Z(n34045) );
  XOR U34481 ( .A(a[123]), .B(b[29]), .Z(n34287) );
  NANDN U34482 ( .A(n34722), .B(n34287), .Z(n34044) );
  AND U34483 ( .A(n34045), .B(n34044), .Z(n34248) );
  NANDN U34484 ( .A(n211), .B(n34046), .Z(n34048) );
  XOR U34485 ( .A(b[47]), .B(a[105]), .Z(n34226) );
  NANDN U34486 ( .A(n37172), .B(n34226), .Z(n34047) );
  NAND U34487 ( .A(n34048), .B(n34047), .Z(n34247) );
  XOR U34488 ( .A(n34248), .B(n34247), .Z(n34250) );
  XOR U34489 ( .A(n34249), .B(n34250), .Z(n34236) );
  NANDN U34490 ( .A(n35611), .B(n34049), .Z(n34051) );
  XOR U34491 ( .A(a[117]), .B(b[35]), .Z(n34180) );
  NANDN U34492 ( .A(n35801), .B(n34180), .Z(n34050) );
  AND U34493 ( .A(n34051), .B(n34050), .Z(n34200) );
  NANDN U34494 ( .A(n35260), .B(n34052), .Z(n34054) );
  XOR U34495 ( .A(a[119]), .B(b[33]), .Z(n34183) );
  NANDN U34496 ( .A(n35456), .B(n34183), .Z(n34053) );
  AND U34497 ( .A(n34054), .B(n34053), .Z(n34199) );
  NANDN U34498 ( .A(n37705), .B(n34055), .Z(n34057) );
  XOR U34499 ( .A(b[53]), .B(a[99]), .Z(n34210) );
  NANDN U34500 ( .A(n37778), .B(n34210), .Z(n34056) );
  NAND U34501 ( .A(n34057), .B(n34056), .Z(n34198) );
  XOR U34502 ( .A(n34199), .B(n34198), .Z(n34201) );
  XNOR U34503 ( .A(n34200), .B(n34201), .Z(n34235) );
  XNOR U34504 ( .A(n34236), .B(n34235), .Z(n34238) );
  NANDN U34505 ( .A(n34059), .B(n34058), .Z(n34063) );
  OR U34506 ( .A(n34061), .B(n34060), .Z(n34062) );
  AND U34507 ( .A(n34063), .B(n34062), .Z(n34237) );
  XOR U34508 ( .A(n34238), .B(n34237), .Z(n34151) );
  NANDN U34509 ( .A(n34223), .B(n34064), .Z(n34066) );
  XOR U34510 ( .A(a[125]), .B(b[27]), .Z(n34222) );
  NANDN U34511 ( .A(n34458), .B(n34222), .Z(n34065) );
  AND U34512 ( .A(n34066), .B(n34065), .Z(n34206) );
  NANDN U34513 ( .A(n38278), .B(n34067), .Z(n34069) );
  XOR U34514 ( .A(b[63]), .B(a[89]), .Z(n34293) );
  NANDN U34515 ( .A(n38279), .B(n34293), .Z(n34068) );
  AND U34516 ( .A(n34069), .B(n34068), .Z(n34205) );
  NANDN U34517 ( .A(n212), .B(n34070), .Z(n34072) );
  XOR U34518 ( .A(b[49]), .B(a[103]), .Z(n34290) );
  NANDN U34519 ( .A(n37432), .B(n34290), .Z(n34071) );
  NAND U34520 ( .A(n34072), .B(n34071), .Z(n34204) );
  XOR U34521 ( .A(n34205), .B(n34204), .Z(n34207) );
  XOR U34522 ( .A(n34206), .B(n34207), .Z(n34242) );
  NANDN U34523 ( .A(n38090), .B(n34073), .Z(n34075) );
  XOR U34524 ( .A(b[59]), .B(a[93]), .Z(n34192) );
  NANDN U34525 ( .A(n38130), .B(n34192), .Z(n34074) );
  AND U34526 ( .A(n34075), .B(n34074), .Z(n34280) );
  NANDN U34527 ( .A(n38247), .B(n34076), .Z(n34078) );
  XOR U34528 ( .A(b[61]), .B(a[91]), .Z(n34219) );
  NANDN U34529 ( .A(n38248), .B(n34219), .Z(n34077) );
  AND U34530 ( .A(n34078), .B(n34077), .Z(n34279) );
  NANDN U34531 ( .A(n37526), .B(n34079), .Z(n34081) );
  XOR U34532 ( .A(b[51]), .B(a[101]), .Z(n34186) );
  NANDN U34533 ( .A(n37605), .B(n34186), .Z(n34080) );
  NAND U34534 ( .A(n34081), .B(n34080), .Z(n34278) );
  XOR U34535 ( .A(n34279), .B(n34278), .Z(n34281) );
  XNOR U34536 ( .A(n34280), .B(n34281), .Z(n34241) );
  XNOR U34537 ( .A(n34242), .B(n34241), .Z(n34244) );
  NANDN U34538 ( .A(n34083), .B(n34082), .Z(n34087) );
  OR U34539 ( .A(n34085), .B(n34084), .Z(n34086) );
  AND U34540 ( .A(n34087), .B(n34086), .Z(n34243) );
  XNOR U34541 ( .A(n34244), .B(n34243), .Z(n34150) );
  XOR U34542 ( .A(n34151), .B(n34150), .Z(n34153) );
  XOR U34543 ( .A(n34152), .B(n34153), .Z(n34170) );
  NANDN U34544 ( .A(n34089), .B(n34088), .Z(n34093) );
  NANDN U34545 ( .A(n34091), .B(n34090), .Z(n34092) );
  AND U34546 ( .A(n34093), .B(n34092), .Z(n34169) );
  NAND U34547 ( .A(n34095), .B(n34094), .Z(n34099) );
  NAND U34548 ( .A(n34097), .B(n34096), .Z(n34098) );
  AND U34549 ( .A(n34099), .B(n34098), .Z(n34168) );
  XOR U34550 ( .A(n34169), .B(n34168), .Z(n34171) );
  XOR U34551 ( .A(n34170), .B(n34171), .Z(n34316) );
  NANDN U34552 ( .A(n34101), .B(n34100), .Z(n34105) );
  NAND U34553 ( .A(n34103), .B(n34102), .Z(n34104) );
  AND U34554 ( .A(n34105), .B(n34104), .Z(n34314) );
  NANDN U34555 ( .A(n34107), .B(n34106), .Z(n34111) );
  NANDN U34556 ( .A(n34109), .B(n34108), .Z(n34110) );
  AND U34557 ( .A(n34111), .B(n34110), .Z(n34313) );
  XNOR U34558 ( .A(n34314), .B(n34313), .Z(n34315) );
  XNOR U34559 ( .A(n34316), .B(n34315), .Z(n34144) );
  NANDN U34560 ( .A(n34113), .B(n34112), .Z(n34117) );
  NANDN U34561 ( .A(n34115), .B(n34114), .Z(n34116) );
  NAND U34562 ( .A(n34117), .B(n34116), .Z(n34145) );
  XNOR U34563 ( .A(n34144), .B(n34145), .Z(n34146) );
  XOR U34564 ( .A(n34147), .B(n34146), .Z(n34139) );
  XNOR U34565 ( .A(n34138), .B(n34139), .Z(n34140) );
  XOR U34566 ( .A(n34141), .B(n34140), .Z(n34133) );
  XOR U34567 ( .A(n34132), .B(n34133), .Z(n34135) );
  XOR U34568 ( .A(n34134), .B(n34135), .Z(n34127) );
  NANDN U34569 ( .A(n34119), .B(n34118), .Z(n34123) );
  NANDN U34570 ( .A(n34121), .B(n34120), .Z(n34122) );
  NAND U34571 ( .A(n34123), .B(n34122), .Z(n34126) );
  XOR U34572 ( .A(n34127), .B(n34126), .Z(n34129) );
  XNOR U34573 ( .A(n34128), .B(n34129), .Z(n34124) );
  XOR U34574 ( .A(n34125), .B(n34124), .Z(c[215]) );
  AND U34575 ( .A(n34125), .B(n34124), .Z(n34320) );
  NANDN U34576 ( .A(n34127), .B(n34126), .Z(n34131) );
  OR U34577 ( .A(n34129), .B(n34128), .Z(n34130) );
  AND U34578 ( .A(n34131), .B(n34130), .Z(n34323) );
  NANDN U34579 ( .A(n34133), .B(n34132), .Z(n34137) );
  OR U34580 ( .A(n34135), .B(n34134), .Z(n34136) );
  AND U34581 ( .A(n34137), .B(n34136), .Z(n34321) );
  NANDN U34582 ( .A(n34139), .B(n34138), .Z(n34143) );
  NANDN U34583 ( .A(n34141), .B(n34140), .Z(n34142) );
  AND U34584 ( .A(n34143), .B(n34142), .Z(n34329) );
  NANDN U34585 ( .A(n34145), .B(n34144), .Z(n34149) );
  NANDN U34586 ( .A(n34147), .B(n34146), .Z(n34148) );
  AND U34587 ( .A(n34149), .B(n34148), .Z(n34327) );
  NANDN U34588 ( .A(n34151), .B(n34150), .Z(n34155) );
  OR U34589 ( .A(n34153), .B(n34152), .Z(n34154) );
  AND U34590 ( .A(n34155), .B(n34154), .Z(n34501) );
  NANDN U34591 ( .A(n34157), .B(n34156), .Z(n34161) );
  NAND U34592 ( .A(n34159), .B(n34158), .Z(n34160) );
  AND U34593 ( .A(n34161), .B(n34160), .Z(n34500) );
  NANDN U34594 ( .A(n34163), .B(n34162), .Z(n34167) );
  NAND U34595 ( .A(n34165), .B(n34164), .Z(n34166) );
  AND U34596 ( .A(n34167), .B(n34166), .Z(n34499) );
  XOR U34597 ( .A(n34500), .B(n34499), .Z(n34502) );
  XOR U34598 ( .A(n34501), .B(n34502), .Z(n34340) );
  NANDN U34599 ( .A(n34169), .B(n34168), .Z(n34173) );
  OR U34600 ( .A(n34171), .B(n34170), .Z(n34172) );
  NAND U34601 ( .A(n34173), .B(n34172), .Z(n34339) );
  XNOR U34602 ( .A(n34340), .B(n34339), .Z(n34341) );
  NANDN U34603 ( .A(n34175), .B(n34174), .Z(n34179) );
  NANDN U34604 ( .A(n34177), .B(n34176), .Z(n34178) );
  AND U34605 ( .A(n34179), .B(n34178), .Z(n34496) );
  NANDN U34606 ( .A(n35611), .B(n34180), .Z(n34182) );
  XOR U34607 ( .A(a[118]), .B(b[35]), .Z(n34472) );
  NANDN U34608 ( .A(n35801), .B(n34472), .Z(n34181) );
  AND U34609 ( .A(n34182), .B(n34181), .Z(n34454) );
  NANDN U34610 ( .A(n35260), .B(n34183), .Z(n34185) );
  XOR U34611 ( .A(a[120]), .B(b[33]), .Z(n34366) );
  NANDN U34612 ( .A(n35456), .B(n34366), .Z(n34184) );
  AND U34613 ( .A(n34185), .B(n34184), .Z(n34453) );
  NANDN U34614 ( .A(n37526), .B(n34186), .Z(n34188) );
  XOR U34615 ( .A(b[51]), .B(a[102]), .Z(n34363) );
  NANDN U34616 ( .A(n37605), .B(n34363), .Z(n34187) );
  NAND U34617 ( .A(n34188), .B(n34187), .Z(n34452) );
  XOR U34618 ( .A(n34453), .B(n34452), .Z(n34455) );
  XOR U34619 ( .A(n34454), .B(n34455), .Z(n34352) );
  NANDN U34620 ( .A(n37974), .B(n34189), .Z(n34191) );
  XOR U34621 ( .A(b[57]), .B(a[96]), .Z(n34469) );
  NANDN U34622 ( .A(n38031), .B(n34469), .Z(n34190) );
  AND U34623 ( .A(n34191), .B(n34190), .Z(n34383) );
  NANDN U34624 ( .A(n38090), .B(n34192), .Z(n34194) );
  XOR U34625 ( .A(b[59]), .B(a[94]), .Z(n34369) );
  NANDN U34626 ( .A(n38130), .B(n34369), .Z(n34193) );
  AND U34627 ( .A(n34194), .B(n34193), .Z(n34382) );
  NANDN U34628 ( .A(n36991), .B(n34195), .Z(n34197) );
  XOR U34629 ( .A(b[45]), .B(a[108]), .Z(n34372) );
  NANDN U34630 ( .A(n37083), .B(n34372), .Z(n34196) );
  NAND U34631 ( .A(n34197), .B(n34196), .Z(n34381) );
  XOR U34632 ( .A(n34382), .B(n34381), .Z(n34384) );
  XNOR U34633 ( .A(n34383), .B(n34384), .Z(n34351) );
  XNOR U34634 ( .A(n34352), .B(n34351), .Z(n34353) );
  NANDN U34635 ( .A(n34199), .B(n34198), .Z(n34203) );
  OR U34636 ( .A(n34201), .B(n34200), .Z(n34202) );
  NAND U34637 ( .A(n34203), .B(n34202), .Z(n34354) );
  XNOR U34638 ( .A(n34353), .B(n34354), .Z(n34487) );
  NANDN U34639 ( .A(n34205), .B(n34204), .Z(n34209) );
  OR U34640 ( .A(n34207), .B(n34206), .Z(n34208) );
  NAND U34641 ( .A(n34209), .B(n34208), .Z(n34488) );
  XNOR U34642 ( .A(n34487), .B(n34488), .Z(n34489) );
  NANDN U34643 ( .A(n37705), .B(n34210), .Z(n34212) );
  XOR U34644 ( .A(b[53]), .B(a[100]), .Z(n34399) );
  NANDN U34645 ( .A(n37778), .B(n34399), .Z(n34211) );
  AND U34646 ( .A(n34212), .B(n34211), .Z(n34377) );
  NANDN U34647 ( .A(n37857), .B(n34213), .Z(n34215) );
  XOR U34648 ( .A(b[55]), .B(a[98]), .Z(n34466) );
  NANDN U34649 ( .A(n37911), .B(n34466), .Z(n34214) );
  AND U34650 ( .A(n34215), .B(n34214), .Z(n34376) );
  NANDN U34651 ( .A(n35936), .B(n34216), .Z(n34218) );
  XOR U34652 ( .A(a[116]), .B(b[37]), .Z(n34405) );
  NANDN U34653 ( .A(n36047), .B(n34405), .Z(n34217) );
  NAND U34654 ( .A(n34218), .B(n34217), .Z(n34375) );
  XOR U34655 ( .A(n34376), .B(n34375), .Z(n34378) );
  XOR U34656 ( .A(n34377), .B(n34378), .Z(n34476) );
  NANDN U34657 ( .A(n38247), .B(n34219), .Z(n34221) );
  XOR U34658 ( .A(b[61]), .B(a[92]), .Z(n34357) );
  NANDN U34659 ( .A(n38248), .B(n34357), .Z(n34220) );
  AND U34660 ( .A(n34221), .B(n34220), .Z(n34448) );
  NANDN U34661 ( .A(n34223), .B(n34222), .Z(n34225) );
  XOR U34662 ( .A(a[126]), .B(b[27]), .Z(n34459) );
  NANDN U34663 ( .A(n34458), .B(n34459), .Z(n34224) );
  AND U34664 ( .A(n34225), .B(n34224), .Z(n34447) );
  NANDN U34665 ( .A(n211), .B(n34226), .Z(n34228) );
  XOR U34666 ( .A(b[47]), .B(a[106]), .Z(n34462) );
  NANDN U34667 ( .A(n37172), .B(n34462), .Z(n34227) );
  NAND U34668 ( .A(n34228), .B(n34227), .Z(n34446) );
  XOR U34669 ( .A(n34447), .B(n34446), .Z(n34449) );
  XNOR U34670 ( .A(n34448), .B(n34449), .Z(n34475) );
  XNOR U34671 ( .A(n34476), .B(n34475), .Z(n34477) );
  NANDN U34672 ( .A(n34230), .B(n34229), .Z(n34234) );
  OR U34673 ( .A(n34232), .B(n34231), .Z(n34233) );
  NAND U34674 ( .A(n34234), .B(n34233), .Z(n34478) );
  XOR U34675 ( .A(n34477), .B(n34478), .Z(n34490) );
  XNOR U34676 ( .A(n34489), .B(n34490), .Z(n34430) );
  NANDN U34677 ( .A(n34236), .B(n34235), .Z(n34240) );
  NAND U34678 ( .A(n34238), .B(n34237), .Z(n34239) );
  AND U34679 ( .A(n34240), .B(n34239), .Z(n34429) );
  NANDN U34680 ( .A(n34242), .B(n34241), .Z(n34246) );
  NAND U34681 ( .A(n34244), .B(n34243), .Z(n34245) );
  NAND U34682 ( .A(n34246), .B(n34245), .Z(n34428) );
  XOR U34683 ( .A(n34429), .B(n34428), .Z(n34431) );
  XNOR U34684 ( .A(n34430), .B(n34431), .Z(n34493) );
  NANDN U34685 ( .A(n34248), .B(n34247), .Z(n34252) );
  OR U34686 ( .A(n34250), .B(n34249), .Z(n34251) );
  AND U34687 ( .A(n34252), .B(n34251), .Z(n34482) );
  XNOR U34688 ( .A(n34482), .B(n34481), .Z(n34484) );
  NANDN U34689 ( .A(n36742), .B(n34257), .Z(n34259) );
  XOR U34690 ( .A(a[110]), .B(b[43]), .Z(n34393) );
  NANDN U34691 ( .A(n36891), .B(n34393), .Z(n34258) );
  AND U34692 ( .A(n34259), .B(n34258), .Z(n34443) );
  NANDN U34693 ( .A(n36480), .B(n34260), .Z(n34262) );
  XOR U34694 ( .A(a[112]), .B(b[41]), .Z(n34396) );
  NANDN U34695 ( .A(n36594), .B(n34396), .Z(n34261) );
  AND U34696 ( .A(n34262), .B(n34261), .Z(n34441) );
  NANDN U34697 ( .A(n36210), .B(n34263), .Z(n34265) );
  XOR U34698 ( .A(a[114]), .B(b[39]), .Z(n34402) );
  NANDN U34699 ( .A(n36347), .B(n34402), .Z(n34264) );
  NAND U34700 ( .A(n34265), .B(n34264), .Z(n34440) );
  XNOR U34701 ( .A(n34441), .B(n34440), .Z(n34442) );
  XNOR U34702 ( .A(n34443), .B(n34442), .Z(n34423) );
  OR U34703 ( .A(n34267), .B(n34266), .Z(n34271) );
  NAND U34704 ( .A(n34269), .B(n34268), .Z(n34270) );
  NAND U34705 ( .A(n34271), .B(n34270), .Z(n34422) );
  XOR U34706 ( .A(n34423), .B(n34422), .Z(n34425) );
  NANDN U34707 ( .A(n34273), .B(n34272), .Z(n34277) );
  NANDN U34708 ( .A(n34275), .B(n34274), .Z(n34276) );
  NAND U34709 ( .A(n34277), .B(n34276), .Z(n34424) );
  XOR U34710 ( .A(n34425), .B(n34424), .Z(n34483) );
  XOR U34711 ( .A(n34484), .B(n34483), .Z(n34437) );
  NANDN U34712 ( .A(n34279), .B(n34278), .Z(n34283) );
  OR U34713 ( .A(n34281), .B(n34280), .Z(n34282) );
  AND U34714 ( .A(n34283), .B(n34282), .Z(n34347) );
  NANDN U34715 ( .A(n34909), .B(n34284), .Z(n34286) );
  XOR U34716 ( .A(a[122]), .B(b[31]), .Z(n34360) );
  NANDN U34717 ( .A(n35145), .B(n34360), .Z(n34285) );
  AND U34718 ( .A(n34286), .B(n34285), .Z(n34389) );
  NANDN U34719 ( .A(n34634), .B(n34287), .Z(n34289) );
  XOR U34720 ( .A(a[124]), .B(b[29]), .Z(n34408) );
  NANDN U34721 ( .A(n34722), .B(n34408), .Z(n34288) );
  AND U34722 ( .A(n34289), .B(n34288), .Z(n34388) );
  NANDN U34723 ( .A(n212), .B(n34290), .Z(n34292) );
  XOR U34724 ( .A(b[49]), .B(a[104]), .Z(n34414) );
  NANDN U34725 ( .A(n37432), .B(n34414), .Z(n34291) );
  NAND U34726 ( .A(n34292), .B(n34291), .Z(n34387) );
  XOR U34727 ( .A(n34388), .B(n34387), .Z(n34390) );
  XOR U34728 ( .A(n34389), .B(n34390), .Z(n34346) );
  NANDN U34729 ( .A(n38278), .B(n34293), .Z(n34295) );
  XOR U34730 ( .A(b[63]), .B(a[90]), .Z(n34411) );
  NANDN U34731 ( .A(n38279), .B(n34411), .Z(n34294) );
  AND U34732 ( .A(n34295), .B(n34294), .Z(n34419) );
  NAND U34733 ( .A(b[63]), .B(a[88]), .Z(n34465) );
  ANDN U34734 ( .B(n34297), .A(n34296), .Z(n34300) );
  NAND U34735 ( .A(b[25]), .B(n34298), .Z(n34299) );
  NANDN U34736 ( .A(n34300), .B(n34299), .Z(n34417) );
  XOR U34737 ( .A(n34465), .B(n34417), .Z(n34418) );
  XOR U34738 ( .A(n34419), .B(n34418), .Z(n34345) );
  XOR U34739 ( .A(n34346), .B(n34345), .Z(n34348) );
  XNOR U34740 ( .A(n34347), .B(n34348), .Z(n34434) );
  NANDN U34741 ( .A(n34302), .B(n34301), .Z(n34306) );
  NANDN U34742 ( .A(n34304), .B(n34303), .Z(n34305) );
  NAND U34743 ( .A(n34306), .B(n34305), .Z(n34435) );
  XNOR U34744 ( .A(n34434), .B(n34435), .Z(n34436) );
  XOR U34745 ( .A(n34437), .B(n34436), .Z(n34494) );
  XNOR U34746 ( .A(n34493), .B(n34494), .Z(n34495) );
  XOR U34747 ( .A(n34496), .B(n34495), .Z(n34342) );
  XNOR U34748 ( .A(n34341), .B(n34342), .Z(n34335) );
  NANDN U34749 ( .A(n34308), .B(n34307), .Z(n34312) );
  OR U34750 ( .A(n34310), .B(n34309), .Z(n34311) );
  AND U34751 ( .A(n34312), .B(n34311), .Z(n34334) );
  NANDN U34752 ( .A(n34314), .B(n34313), .Z(n34318) );
  NANDN U34753 ( .A(n34316), .B(n34315), .Z(n34317) );
  AND U34754 ( .A(n34318), .B(n34317), .Z(n34333) );
  XOR U34755 ( .A(n34334), .B(n34333), .Z(n34336) );
  XOR U34756 ( .A(n34335), .B(n34336), .Z(n34328) );
  XOR U34757 ( .A(n34327), .B(n34328), .Z(n34330) );
  XOR U34758 ( .A(n34329), .B(n34330), .Z(n34322) );
  XOR U34759 ( .A(n34321), .B(n34322), .Z(n34324) );
  XNOR U34760 ( .A(n34323), .B(n34324), .Z(n34319) );
  XOR U34761 ( .A(n34320), .B(n34319), .Z(c[216]) );
  AND U34762 ( .A(n34320), .B(n34319), .Z(n34506) );
  NANDN U34763 ( .A(n34322), .B(n34321), .Z(n34326) );
  OR U34764 ( .A(n34324), .B(n34323), .Z(n34325) );
  AND U34765 ( .A(n34326), .B(n34325), .Z(n34509) );
  NANDN U34766 ( .A(n34328), .B(n34327), .Z(n34332) );
  NANDN U34767 ( .A(n34330), .B(n34329), .Z(n34331) );
  AND U34768 ( .A(n34332), .B(n34331), .Z(n34508) );
  NANDN U34769 ( .A(n34334), .B(n34333), .Z(n34338) );
  NANDN U34770 ( .A(n34336), .B(n34335), .Z(n34337) );
  AND U34771 ( .A(n34338), .B(n34337), .Z(n34516) );
  NANDN U34772 ( .A(n34340), .B(n34339), .Z(n34344) );
  NANDN U34773 ( .A(n34342), .B(n34341), .Z(n34343) );
  AND U34774 ( .A(n34344), .B(n34343), .Z(n34514) );
  NANDN U34775 ( .A(n34346), .B(n34345), .Z(n34350) );
  NANDN U34776 ( .A(n34348), .B(n34347), .Z(n34349) );
  AND U34777 ( .A(n34350), .B(n34349), .Z(n34533) );
  NANDN U34778 ( .A(n34352), .B(n34351), .Z(n34356) );
  NANDN U34779 ( .A(n34354), .B(n34353), .Z(n34355) );
  AND U34780 ( .A(n34356), .B(n34355), .Z(n34678) );
  NANDN U34781 ( .A(n38247), .B(n34357), .Z(n34359) );
  XOR U34782 ( .A(b[61]), .B(a[93]), .Z(n34637) );
  NANDN U34783 ( .A(n38248), .B(n34637), .Z(n34358) );
  AND U34784 ( .A(n34359), .B(n34358), .Z(n34602) );
  NANDN U34785 ( .A(n34909), .B(n34360), .Z(n34362) );
  XOR U34786 ( .A(a[123]), .B(b[31]), .Z(n34573) );
  NANDN U34787 ( .A(n35145), .B(n34573), .Z(n34361) );
  AND U34788 ( .A(n34362), .B(n34361), .Z(n34601) );
  NANDN U34789 ( .A(n37526), .B(n34363), .Z(n34365) );
  XOR U34790 ( .A(b[51]), .B(a[103]), .Z(n34570) );
  NANDN U34791 ( .A(n37605), .B(n34570), .Z(n34364) );
  NAND U34792 ( .A(n34365), .B(n34364), .Z(n34600) );
  XOR U34793 ( .A(n34601), .B(n34600), .Z(n34603) );
  XOR U34794 ( .A(n34602), .B(n34603), .Z(n34664) );
  NANDN U34795 ( .A(n35260), .B(n34366), .Z(n34368) );
  XOR U34796 ( .A(a[121]), .B(b[33]), .Z(n34567) );
  NANDN U34797 ( .A(n35456), .B(n34567), .Z(n34367) );
  AND U34798 ( .A(n34368), .B(n34367), .Z(n34584) );
  NANDN U34799 ( .A(n38090), .B(n34369), .Z(n34371) );
  XOR U34800 ( .A(b[59]), .B(a[95]), .Z(n34576) );
  NANDN U34801 ( .A(n38130), .B(n34576), .Z(n34370) );
  AND U34802 ( .A(n34371), .B(n34370), .Z(n34583) );
  NANDN U34803 ( .A(n36991), .B(n34372), .Z(n34374) );
  XOR U34804 ( .A(b[45]), .B(a[109]), .Z(n34624) );
  NANDN U34805 ( .A(n37083), .B(n34624), .Z(n34373) );
  NAND U34806 ( .A(n34374), .B(n34373), .Z(n34582) );
  XOR U34807 ( .A(n34583), .B(n34582), .Z(n34585) );
  XNOR U34808 ( .A(n34584), .B(n34585), .Z(n34663) );
  XNOR U34809 ( .A(n34664), .B(n34663), .Z(n34666) );
  NANDN U34810 ( .A(n34376), .B(n34375), .Z(n34380) );
  OR U34811 ( .A(n34378), .B(n34377), .Z(n34379) );
  AND U34812 ( .A(n34380), .B(n34379), .Z(n34665) );
  XOR U34813 ( .A(n34666), .B(n34665), .Z(n34545) );
  NANDN U34814 ( .A(n34382), .B(n34381), .Z(n34386) );
  OR U34815 ( .A(n34384), .B(n34383), .Z(n34385) );
  AND U34816 ( .A(n34386), .B(n34385), .Z(n34544) );
  NANDN U34817 ( .A(n34388), .B(n34387), .Z(n34392) );
  OR U34818 ( .A(n34390), .B(n34389), .Z(n34391) );
  NAND U34819 ( .A(n34392), .B(n34391), .Z(n34543) );
  XOR U34820 ( .A(n34544), .B(n34543), .Z(n34546) );
  XOR U34821 ( .A(n34545), .B(n34546), .Z(n34676) );
  NANDN U34822 ( .A(n36742), .B(n34393), .Z(n34395) );
  XOR U34823 ( .A(a[111]), .B(b[43]), .Z(n34555) );
  NANDN U34824 ( .A(n36891), .B(n34555), .Z(n34394) );
  AND U34825 ( .A(n34395), .B(n34394), .Z(n34596) );
  NANDN U34826 ( .A(n36480), .B(n34396), .Z(n34398) );
  XOR U34827 ( .A(a[113]), .B(b[41]), .Z(n34552) );
  NANDN U34828 ( .A(n36594), .B(n34552), .Z(n34397) );
  AND U34829 ( .A(n34398), .B(n34397), .Z(n34595) );
  NAND U34830 ( .A(n37849), .B(n34399), .Z(n34401) );
  XNOR U34831 ( .A(b[53]), .B(a[101]), .Z(n34558) );
  NANDN U34832 ( .A(n34558), .B(n37850), .Z(n34400) );
  NAND U34833 ( .A(n34401), .B(n34400), .Z(n34652) );
  NANDN U34834 ( .A(n36210), .B(n34402), .Z(n34404) );
  XOR U34835 ( .A(a[115]), .B(b[39]), .Z(n34549) );
  NANDN U34836 ( .A(n36347), .B(n34549), .Z(n34403) );
  NAND U34837 ( .A(n34404), .B(n34403), .Z(n34651) );
  XOR U34838 ( .A(n34652), .B(n34651), .Z(n34654) );
  NAND U34839 ( .A(n36238), .B(n34405), .Z(n34407) );
  XNOR U34840 ( .A(a[117]), .B(b[37]), .Z(n34561) );
  NANDN U34841 ( .A(n34561), .B(n36239), .Z(n34406) );
  NAND U34842 ( .A(n34407), .B(n34406), .Z(n34653) );
  XOR U34843 ( .A(n34654), .B(n34653), .Z(n34594) );
  XOR U34844 ( .A(n34595), .B(n34594), .Z(n34597) );
  XOR U34845 ( .A(n34596), .B(n34597), .Z(n34540) );
  NANDN U34846 ( .A(n34634), .B(n34408), .Z(n34410) );
  XOR U34847 ( .A(a[125]), .B(b[29]), .Z(n34633) );
  NANDN U34848 ( .A(n34722), .B(n34633), .Z(n34409) );
  AND U34849 ( .A(n34410), .B(n34409), .Z(n34608) );
  NANDN U34850 ( .A(n38278), .B(n34411), .Z(n34413) );
  XOR U34851 ( .A(b[63]), .B(a[91]), .Z(n34643) );
  NANDN U34852 ( .A(n38279), .B(n34643), .Z(n34412) );
  AND U34853 ( .A(n34413), .B(n34412), .Z(n34607) );
  NANDN U34854 ( .A(n212), .B(n34414), .Z(n34416) );
  XOR U34855 ( .A(b[49]), .B(a[105]), .Z(n34579) );
  NANDN U34856 ( .A(n37432), .B(n34579), .Z(n34415) );
  NAND U34857 ( .A(n34416), .B(n34415), .Z(n34606) );
  XOR U34858 ( .A(n34607), .B(n34606), .Z(n34609) );
  XOR U34859 ( .A(n34608), .B(n34609), .Z(n34538) );
  IV U34860 ( .A(n34465), .Z(n34621) );
  NANDN U34861 ( .A(n34621), .B(n34417), .Z(n34421) );
  NANDN U34862 ( .A(n34419), .B(n34418), .Z(n34420) );
  AND U34863 ( .A(n34421), .B(n34420), .Z(n34537) );
  XNOR U34864 ( .A(n34538), .B(n34537), .Z(n34539) );
  XNOR U34865 ( .A(n34540), .B(n34539), .Z(n34675) );
  XNOR U34866 ( .A(n34676), .B(n34675), .Z(n34677) );
  XNOR U34867 ( .A(n34678), .B(n34677), .Z(n34531) );
  NAND U34868 ( .A(n34423), .B(n34422), .Z(n34427) );
  NAND U34869 ( .A(n34425), .B(n34424), .Z(n34426) );
  NAND U34870 ( .A(n34427), .B(n34426), .Z(n34532) );
  XOR U34871 ( .A(n34531), .B(n34532), .Z(n34534) );
  XOR U34872 ( .A(n34533), .B(n34534), .Z(n34688) );
  NANDN U34873 ( .A(n34429), .B(n34428), .Z(n34433) );
  NANDN U34874 ( .A(n34431), .B(n34430), .Z(n34432) );
  AND U34875 ( .A(n34433), .B(n34432), .Z(n34687) );
  XNOR U34876 ( .A(n34688), .B(n34687), .Z(n34690) );
  NANDN U34877 ( .A(n34435), .B(n34434), .Z(n34439) );
  NANDN U34878 ( .A(n34437), .B(n34436), .Z(n34438) );
  AND U34879 ( .A(n34439), .B(n34438), .Z(n34527) );
  NANDN U34880 ( .A(n34441), .B(n34440), .Z(n34445) );
  NANDN U34881 ( .A(n34443), .B(n34442), .Z(n34444) );
  AND U34882 ( .A(n34445), .B(n34444), .Z(n34670) );
  NANDN U34883 ( .A(n34447), .B(n34446), .Z(n34451) );
  OR U34884 ( .A(n34449), .B(n34448), .Z(n34450) );
  NAND U34885 ( .A(n34451), .B(n34450), .Z(n34669) );
  XNOR U34886 ( .A(n34670), .B(n34669), .Z(n34672) );
  NANDN U34887 ( .A(n34453), .B(n34452), .Z(n34457) );
  OR U34888 ( .A(n34455), .B(n34454), .Z(n34456) );
  AND U34889 ( .A(n34457), .B(n34456), .Z(n34660) );
  XNOR U34890 ( .A(a[127]), .B(b[27]), .Z(n34646) );
  OR U34891 ( .A(n34646), .B(n34458), .Z(n34461) );
  NAND U34892 ( .A(n34647), .B(n34459), .Z(n34460) );
  AND U34893 ( .A(n34461), .B(n34460), .Z(n34589) );
  NANDN U34894 ( .A(n211), .B(n34462), .Z(n34464) );
  XOR U34895 ( .A(b[47]), .B(a[107]), .Z(n34640) );
  NANDN U34896 ( .A(n37172), .B(n34640), .Z(n34463) );
  NAND U34897 ( .A(n34464), .B(n34463), .Z(n34588) );
  XNOR U34898 ( .A(n34589), .B(n34588), .Z(n34590) );
  AND U34899 ( .A(b[63]), .B(a[89]), .Z(n34618) );
  XOR U34900 ( .A(n34619), .B(n34618), .Z(n34620) );
  XOR U34901 ( .A(n34465), .B(n34620), .Z(n34591) );
  XOR U34902 ( .A(n34590), .B(n34591), .Z(n34657) );
  NANDN U34903 ( .A(n37857), .B(n34466), .Z(n34468) );
  XOR U34904 ( .A(b[55]), .B(a[99]), .Z(n34627) );
  NANDN U34905 ( .A(n37911), .B(n34627), .Z(n34467) );
  AND U34906 ( .A(n34468), .B(n34467), .Z(n34615) );
  NANDN U34907 ( .A(n37974), .B(n34469), .Z(n34471) );
  XOR U34908 ( .A(b[57]), .B(a[97]), .Z(n34630) );
  NANDN U34909 ( .A(n38031), .B(n34630), .Z(n34470) );
  AND U34910 ( .A(n34471), .B(n34470), .Z(n34613) );
  NANDN U34911 ( .A(n35611), .B(n34472), .Z(n34474) );
  XOR U34912 ( .A(a[119]), .B(b[35]), .Z(n34564) );
  NANDN U34913 ( .A(n35801), .B(n34564), .Z(n34473) );
  NAND U34914 ( .A(n34474), .B(n34473), .Z(n34612) );
  XNOR U34915 ( .A(n34613), .B(n34612), .Z(n34614) );
  XOR U34916 ( .A(n34615), .B(n34614), .Z(n34658) );
  XNOR U34917 ( .A(n34657), .B(n34658), .Z(n34659) );
  XNOR U34918 ( .A(n34660), .B(n34659), .Z(n34671) );
  XOR U34919 ( .A(n34672), .B(n34671), .Z(n34682) );
  NANDN U34920 ( .A(n34476), .B(n34475), .Z(n34480) );
  NANDN U34921 ( .A(n34478), .B(n34477), .Z(n34479) );
  NAND U34922 ( .A(n34480), .B(n34479), .Z(n34681) );
  XNOR U34923 ( .A(n34682), .B(n34681), .Z(n34684) );
  NANDN U34924 ( .A(n34482), .B(n34481), .Z(n34486) );
  NAND U34925 ( .A(n34484), .B(n34483), .Z(n34485) );
  AND U34926 ( .A(n34486), .B(n34485), .Z(n34683) );
  XOR U34927 ( .A(n34684), .B(n34683), .Z(n34526) );
  NANDN U34928 ( .A(n34488), .B(n34487), .Z(n34492) );
  NANDN U34929 ( .A(n34490), .B(n34489), .Z(n34491) );
  AND U34930 ( .A(n34492), .B(n34491), .Z(n34525) );
  XOR U34931 ( .A(n34526), .B(n34525), .Z(n34528) );
  XNOR U34932 ( .A(n34527), .B(n34528), .Z(n34689) );
  XOR U34933 ( .A(n34690), .B(n34689), .Z(n34522) );
  NANDN U34934 ( .A(n34494), .B(n34493), .Z(n34498) );
  NANDN U34935 ( .A(n34496), .B(n34495), .Z(n34497) );
  AND U34936 ( .A(n34498), .B(n34497), .Z(n34520) );
  NANDN U34937 ( .A(n34500), .B(n34499), .Z(n34504) );
  OR U34938 ( .A(n34502), .B(n34501), .Z(n34503) );
  AND U34939 ( .A(n34504), .B(n34503), .Z(n34519) );
  XNOR U34940 ( .A(n34520), .B(n34519), .Z(n34521) );
  XNOR U34941 ( .A(n34522), .B(n34521), .Z(n34513) );
  XNOR U34942 ( .A(n34514), .B(n34513), .Z(n34515) );
  XNOR U34943 ( .A(n34516), .B(n34515), .Z(n34507) );
  XOR U34944 ( .A(n34508), .B(n34507), .Z(n34510) );
  XNOR U34945 ( .A(n34509), .B(n34510), .Z(n34505) );
  XOR U34946 ( .A(n34506), .B(n34505), .Z(c[217]) );
  AND U34947 ( .A(n34506), .B(n34505), .Z(n34694) );
  NANDN U34948 ( .A(n34508), .B(n34507), .Z(n34512) );
  OR U34949 ( .A(n34510), .B(n34509), .Z(n34511) );
  AND U34950 ( .A(n34512), .B(n34511), .Z(n34697) );
  NANDN U34951 ( .A(n34514), .B(n34513), .Z(n34518) );
  NANDN U34952 ( .A(n34516), .B(n34515), .Z(n34517) );
  AND U34953 ( .A(n34518), .B(n34517), .Z(n34696) );
  NANDN U34954 ( .A(n34520), .B(n34519), .Z(n34524) );
  NANDN U34955 ( .A(n34522), .B(n34521), .Z(n34523) );
  AND U34956 ( .A(n34524), .B(n34523), .Z(n34704) );
  NANDN U34957 ( .A(n34526), .B(n34525), .Z(n34530) );
  NANDN U34958 ( .A(n34528), .B(n34527), .Z(n34529) );
  AND U34959 ( .A(n34530), .B(n34529), .Z(n34708) );
  NANDN U34960 ( .A(n34532), .B(n34531), .Z(n34536) );
  OR U34961 ( .A(n34534), .B(n34533), .Z(n34535) );
  AND U34962 ( .A(n34536), .B(n34535), .Z(n34707) );
  XNOR U34963 ( .A(n34708), .B(n34707), .Z(n34710) );
  NANDN U34964 ( .A(n34538), .B(n34537), .Z(n34542) );
  NANDN U34965 ( .A(n34540), .B(n34539), .Z(n34541) );
  AND U34966 ( .A(n34542), .B(n34541), .Z(n34810) );
  NANDN U34967 ( .A(n34544), .B(n34543), .Z(n34548) );
  OR U34968 ( .A(n34546), .B(n34545), .Z(n34547) );
  AND U34969 ( .A(n34548), .B(n34547), .Z(n34808) );
  NANDN U34970 ( .A(n36210), .B(n34549), .Z(n34551) );
  XOR U34971 ( .A(a[116]), .B(b[39]), .Z(n34762) );
  NANDN U34972 ( .A(n36347), .B(n34762), .Z(n34550) );
  AND U34973 ( .A(n34551), .B(n34550), .Z(n34767) );
  NANDN U34974 ( .A(n36480), .B(n34552), .Z(n34554) );
  XOR U34975 ( .A(a[114]), .B(b[41]), .Z(n34753) );
  NANDN U34976 ( .A(n36594), .B(n34753), .Z(n34553) );
  AND U34977 ( .A(n34554), .B(n34553), .Z(n34766) );
  NANDN U34978 ( .A(n36742), .B(n34555), .Z(n34557) );
  XOR U34979 ( .A(a[112]), .B(b[43]), .Z(n34756) );
  NANDN U34980 ( .A(n36891), .B(n34756), .Z(n34556) );
  AND U34981 ( .A(n34557), .B(n34556), .Z(n34861) );
  NANDN U34982 ( .A(n34558), .B(n37849), .Z(n34560) );
  XOR U34983 ( .A(b[53]), .B(a[102]), .Z(n34750) );
  NANDN U34984 ( .A(n37778), .B(n34750), .Z(n34559) );
  AND U34985 ( .A(n34560), .B(n34559), .Z(n34859) );
  NANDN U34986 ( .A(n34561), .B(n36238), .Z(n34563) );
  XOR U34987 ( .A(a[118]), .B(b[37]), .Z(n34759) );
  NANDN U34988 ( .A(n36047), .B(n34759), .Z(n34562) );
  NAND U34989 ( .A(n34563), .B(n34562), .Z(n34858) );
  XNOR U34990 ( .A(n34859), .B(n34858), .Z(n34860) );
  XNOR U34991 ( .A(n34861), .B(n34860), .Z(n34765) );
  XOR U34992 ( .A(n34766), .B(n34765), .Z(n34768) );
  XOR U34993 ( .A(n34767), .B(n34768), .Z(n34797) );
  NANDN U34994 ( .A(n35611), .B(n34564), .Z(n34566) );
  XOR U34995 ( .A(a[120]), .B(b[35]), .Z(n34744) );
  NANDN U34996 ( .A(n35801), .B(n34744), .Z(n34565) );
  AND U34997 ( .A(n34566), .B(n34565), .Z(n34833) );
  NANDN U34998 ( .A(n35260), .B(n34567), .Z(n34569) );
  XOR U34999 ( .A(a[122]), .B(b[33]), .Z(n34845) );
  NANDN U35000 ( .A(n35456), .B(n34845), .Z(n34568) );
  AND U35001 ( .A(n34569), .B(n34568), .Z(n34832) );
  NANDN U35002 ( .A(n37526), .B(n34570), .Z(n34572) );
  XOR U35003 ( .A(b[51]), .B(a[104]), .Z(n34735) );
  NANDN U35004 ( .A(n37605), .B(n34735), .Z(n34571) );
  NAND U35005 ( .A(n34572), .B(n34571), .Z(n34831) );
  XOR U35006 ( .A(n34832), .B(n34831), .Z(n34834) );
  XOR U35007 ( .A(n34833), .B(n34834), .Z(n34796) );
  NANDN U35008 ( .A(n34909), .B(n34573), .Z(n34575) );
  XOR U35009 ( .A(a[124]), .B(b[31]), .Z(n34719) );
  NANDN U35010 ( .A(n35145), .B(n34719), .Z(n34574) );
  AND U35011 ( .A(n34575), .B(n34574), .Z(n34773) );
  NANDN U35012 ( .A(n38090), .B(n34576), .Z(n34578) );
  XOR U35013 ( .A(b[59]), .B(a[96]), .Z(n34729) );
  NANDN U35014 ( .A(n38130), .B(n34729), .Z(n34577) );
  AND U35015 ( .A(n34578), .B(n34577), .Z(n34772) );
  NANDN U35016 ( .A(n212), .B(n34579), .Z(n34581) );
  XOR U35017 ( .A(b[49]), .B(a[106]), .Z(n34747) );
  NANDN U35018 ( .A(n37432), .B(n34747), .Z(n34580) );
  NAND U35019 ( .A(n34581), .B(n34580), .Z(n34771) );
  XOR U35020 ( .A(n34772), .B(n34771), .Z(n34774) );
  XNOR U35021 ( .A(n34773), .B(n34774), .Z(n34795) );
  XOR U35022 ( .A(n34796), .B(n34795), .Z(n34798) );
  XOR U35023 ( .A(n34797), .B(n34798), .Z(n34786) );
  NANDN U35024 ( .A(n34583), .B(n34582), .Z(n34587) );
  OR U35025 ( .A(n34585), .B(n34584), .Z(n34586) );
  AND U35026 ( .A(n34587), .B(n34586), .Z(n34784) );
  NANDN U35027 ( .A(n34589), .B(n34588), .Z(n34593) );
  NAND U35028 ( .A(n34591), .B(n34590), .Z(n34592) );
  NAND U35029 ( .A(n34593), .B(n34592), .Z(n34783) );
  XNOR U35030 ( .A(n34784), .B(n34783), .Z(n34785) );
  XNOR U35031 ( .A(n34786), .B(n34785), .Z(n34807) );
  XNOR U35032 ( .A(n34808), .B(n34807), .Z(n34809) );
  XOR U35033 ( .A(n34810), .B(n34809), .Z(n34803) );
  NANDN U35034 ( .A(n34595), .B(n34594), .Z(n34599) );
  OR U35035 ( .A(n34597), .B(n34596), .Z(n34598) );
  AND U35036 ( .A(n34599), .B(n34598), .Z(n34821) );
  NANDN U35037 ( .A(n34601), .B(n34600), .Z(n34605) );
  OR U35038 ( .A(n34603), .B(n34602), .Z(n34604) );
  AND U35039 ( .A(n34605), .B(n34604), .Z(n34820) );
  NANDN U35040 ( .A(n34607), .B(n34606), .Z(n34611) );
  OR U35041 ( .A(n34609), .B(n34608), .Z(n34610) );
  NAND U35042 ( .A(n34611), .B(n34610), .Z(n34819) );
  XOR U35043 ( .A(n34820), .B(n34819), .Z(n34822) );
  XOR U35044 ( .A(n34821), .B(n34822), .Z(n34715) );
  NANDN U35045 ( .A(n34613), .B(n34612), .Z(n34617) );
  NANDN U35046 ( .A(n34615), .B(n34614), .Z(n34616) );
  AND U35047 ( .A(n34617), .B(n34616), .Z(n34827) );
  NANDN U35048 ( .A(n34619), .B(n34618), .Z(n34623) );
  ANDN U35049 ( .B(n34621), .A(n34620), .Z(n34622) );
  ANDN U35050 ( .B(n34623), .A(n34622), .Z(n34826) );
  NANDN U35051 ( .A(n36991), .B(n34624), .Z(n34626) );
  XOR U35052 ( .A(b[45]), .B(a[110]), .Z(n34726) );
  NANDN U35053 ( .A(n37083), .B(n34726), .Z(n34625) );
  AND U35054 ( .A(n34626), .B(n34625), .Z(n34741) );
  NANDN U35055 ( .A(n37857), .B(n34627), .Z(n34629) );
  XOR U35056 ( .A(b[55]), .B(a[100]), .Z(n34848) );
  NANDN U35057 ( .A(n37911), .B(n34848), .Z(n34628) );
  AND U35058 ( .A(n34629), .B(n34628), .Z(n34739) );
  NANDN U35059 ( .A(n37974), .B(n34630), .Z(n34632) );
  XOR U35060 ( .A(b[57]), .B(a[98]), .Z(n34842) );
  NANDN U35061 ( .A(n38031), .B(n34842), .Z(n34631) );
  NAND U35062 ( .A(n34632), .B(n34631), .Z(n34738) );
  XNOR U35063 ( .A(n34739), .B(n34738), .Z(n34740) );
  XNOR U35064 ( .A(n34741), .B(n34740), .Z(n34825) );
  XOR U35065 ( .A(n34826), .B(n34825), .Z(n34828) );
  XOR U35066 ( .A(n34827), .B(n34828), .Z(n34714) );
  NANDN U35067 ( .A(n34634), .B(n34633), .Z(n34636) );
  XOR U35068 ( .A(a[126]), .B(b[29]), .Z(n34723) );
  NANDN U35069 ( .A(n34722), .B(n34723), .Z(n34635) );
  AND U35070 ( .A(n34636), .B(n34635), .Z(n34779) );
  NANDN U35071 ( .A(n38247), .B(n34637), .Z(n34639) );
  XOR U35072 ( .A(b[61]), .B(a[94]), .Z(n34732) );
  NANDN U35073 ( .A(n38248), .B(n34732), .Z(n34638) );
  AND U35074 ( .A(n34639), .B(n34638), .Z(n34778) );
  NANDN U35075 ( .A(n211), .B(n34640), .Z(n34642) );
  XOR U35076 ( .A(b[47]), .B(a[108]), .Z(n34854) );
  NANDN U35077 ( .A(n37172), .B(n34854), .Z(n34641) );
  NAND U35078 ( .A(n34642), .B(n34641), .Z(n34777) );
  XOR U35079 ( .A(n34778), .B(n34777), .Z(n34780) );
  XOR U35080 ( .A(n34779), .B(n34780), .Z(n34790) );
  NANDN U35081 ( .A(n38278), .B(n34643), .Z(n34645) );
  XOR U35082 ( .A(b[63]), .B(a[92]), .Z(n34851) );
  NANDN U35083 ( .A(n38279), .B(n34851), .Z(n34644) );
  AND U35084 ( .A(n34645), .B(n34644), .Z(n34839) );
  NAND U35085 ( .A(b[63]), .B(a[90]), .Z(n34857) );
  ANDN U35086 ( .B(n34647), .A(n34646), .Z(n34650) );
  NAND U35087 ( .A(b[27]), .B(n34648), .Z(n34649) );
  NANDN U35088 ( .A(n34650), .B(n34649), .Z(n34837) );
  XOR U35089 ( .A(n34857), .B(n34837), .Z(n34838) );
  XOR U35090 ( .A(n34839), .B(n34838), .Z(n34789) );
  XNOR U35091 ( .A(n34790), .B(n34789), .Z(n34791) );
  NAND U35092 ( .A(n34652), .B(n34651), .Z(n34656) );
  NAND U35093 ( .A(n34654), .B(n34653), .Z(n34655) );
  NAND U35094 ( .A(n34656), .B(n34655), .Z(n34792) );
  XNOR U35095 ( .A(n34791), .B(n34792), .Z(n34713) );
  XOR U35096 ( .A(n34714), .B(n34713), .Z(n34716) );
  XOR U35097 ( .A(n34715), .B(n34716), .Z(n34815) );
  NANDN U35098 ( .A(n34658), .B(n34657), .Z(n34662) );
  NANDN U35099 ( .A(n34660), .B(n34659), .Z(n34661) );
  AND U35100 ( .A(n34662), .B(n34661), .Z(n34814) );
  NANDN U35101 ( .A(n34664), .B(n34663), .Z(n34668) );
  NAND U35102 ( .A(n34666), .B(n34665), .Z(n34667) );
  AND U35103 ( .A(n34668), .B(n34667), .Z(n34813) );
  XOR U35104 ( .A(n34814), .B(n34813), .Z(n34816) );
  XOR U35105 ( .A(n34815), .B(n34816), .Z(n34802) );
  NANDN U35106 ( .A(n34670), .B(n34669), .Z(n34674) );
  NAND U35107 ( .A(n34672), .B(n34671), .Z(n34673) );
  AND U35108 ( .A(n34674), .B(n34673), .Z(n34801) );
  XOR U35109 ( .A(n34802), .B(n34801), .Z(n34804) );
  XOR U35110 ( .A(n34803), .B(n34804), .Z(n34867) );
  NANDN U35111 ( .A(n34676), .B(n34675), .Z(n34680) );
  NANDN U35112 ( .A(n34678), .B(n34677), .Z(n34679) );
  AND U35113 ( .A(n34680), .B(n34679), .Z(n34864) );
  NANDN U35114 ( .A(n34682), .B(n34681), .Z(n34686) );
  NAND U35115 ( .A(n34684), .B(n34683), .Z(n34685) );
  NAND U35116 ( .A(n34686), .B(n34685), .Z(n34865) );
  XNOR U35117 ( .A(n34864), .B(n34865), .Z(n34866) );
  XNOR U35118 ( .A(n34867), .B(n34866), .Z(n34709) );
  XOR U35119 ( .A(n34710), .B(n34709), .Z(n34702) );
  NANDN U35120 ( .A(n34688), .B(n34687), .Z(n34692) );
  NAND U35121 ( .A(n34690), .B(n34689), .Z(n34691) );
  AND U35122 ( .A(n34692), .B(n34691), .Z(n34701) );
  XNOR U35123 ( .A(n34702), .B(n34701), .Z(n34703) );
  XNOR U35124 ( .A(n34704), .B(n34703), .Z(n34695) );
  XOR U35125 ( .A(n34696), .B(n34695), .Z(n34698) );
  XNOR U35126 ( .A(n34697), .B(n34698), .Z(n34693) );
  XOR U35127 ( .A(n34694), .B(n34693), .Z(c[218]) );
  AND U35128 ( .A(n34694), .B(n34693), .Z(n34871) );
  NANDN U35129 ( .A(n34696), .B(n34695), .Z(n34700) );
  OR U35130 ( .A(n34698), .B(n34697), .Z(n34699) );
  AND U35131 ( .A(n34700), .B(n34699), .Z(n34874) );
  NANDN U35132 ( .A(n34702), .B(n34701), .Z(n34706) );
  NANDN U35133 ( .A(n34704), .B(n34703), .Z(n34705) );
  AND U35134 ( .A(n34706), .B(n34705), .Z(n34873) );
  NANDN U35135 ( .A(n34708), .B(n34707), .Z(n34712) );
  NAND U35136 ( .A(n34710), .B(n34709), .Z(n34711) );
  AND U35137 ( .A(n34712), .B(n34711), .Z(n34880) );
  NANDN U35138 ( .A(n34714), .B(n34713), .Z(n34718) );
  OR U35139 ( .A(n34716), .B(n34715), .Z(n34717) );
  AND U35140 ( .A(n34718), .B(n34717), .Z(n34942) );
  NANDN U35141 ( .A(n34909), .B(n34719), .Z(n34721) );
  XOR U35142 ( .A(a[125]), .B(b[31]), .Z(n34908) );
  NANDN U35143 ( .A(n35145), .B(n34908), .Z(n34720) );
  AND U35144 ( .A(n34721), .B(n34720), .Z(n34981) );
  XNOR U35145 ( .A(a[127]), .B(b[29]), .Z(n35000) );
  OR U35146 ( .A(n35000), .B(n34722), .Z(n34725) );
  NAND U35147 ( .A(n35001), .B(n34723), .Z(n34724) );
  AND U35148 ( .A(n34725), .B(n34724), .Z(n34980) );
  NANDN U35149 ( .A(n36991), .B(n34726), .Z(n34728) );
  XOR U35150 ( .A(b[45]), .B(a[111]), .Z(n35011) );
  NANDN U35151 ( .A(n37083), .B(n35011), .Z(n34727) );
  NAND U35152 ( .A(n34728), .B(n34727), .Z(n34979) );
  XOR U35153 ( .A(n34980), .B(n34979), .Z(n34982) );
  XOR U35154 ( .A(n34981), .B(n34982), .Z(n35042) );
  NANDN U35155 ( .A(n38090), .B(n34729), .Z(n34731) );
  XOR U35156 ( .A(b[59]), .B(a[97]), .Z(n35014) );
  NANDN U35157 ( .A(n38130), .B(n35014), .Z(n34730) );
  AND U35158 ( .A(n34731), .B(n34730), .Z(n34975) );
  NANDN U35159 ( .A(n38247), .B(n34732), .Z(n34734) );
  XOR U35160 ( .A(b[61]), .B(a[95]), .Z(n35017) );
  NANDN U35161 ( .A(n38248), .B(n35017), .Z(n34733) );
  AND U35162 ( .A(n34734), .B(n34733), .Z(n34974) );
  NANDN U35163 ( .A(n37526), .B(n34735), .Z(n34737) );
  XOR U35164 ( .A(b[51]), .B(a[105]), .Z(n34958) );
  NANDN U35165 ( .A(n37605), .B(n34958), .Z(n34736) );
  NAND U35166 ( .A(n34737), .B(n34736), .Z(n34973) );
  XOR U35167 ( .A(n34974), .B(n34973), .Z(n34976) );
  XNOR U35168 ( .A(n34975), .B(n34976), .Z(n35041) );
  XNOR U35169 ( .A(n35042), .B(n35041), .Z(n35044) );
  NANDN U35170 ( .A(n34739), .B(n34738), .Z(n34743) );
  NANDN U35171 ( .A(n34741), .B(n34740), .Z(n34742) );
  AND U35172 ( .A(n34743), .B(n34742), .Z(n35043) );
  XOR U35173 ( .A(n35044), .B(n35043), .Z(n34947) );
  NANDN U35174 ( .A(n35611), .B(n34744), .Z(n34746) );
  XOR U35175 ( .A(a[121]), .B(b[35]), .Z(n34967) );
  NANDN U35176 ( .A(n35801), .B(n34967), .Z(n34745) );
  AND U35177 ( .A(n34746), .B(n34745), .Z(n34987) );
  NANDN U35178 ( .A(n212), .B(n34747), .Z(n34749) );
  XOR U35179 ( .A(b[49]), .B(a[107]), .Z(n35020) );
  NANDN U35180 ( .A(n37432), .B(n35020), .Z(n34748) );
  AND U35181 ( .A(n34749), .B(n34748), .Z(n34986) );
  NANDN U35182 ( .A(n37705), .B(n34750), .Z(n34752) );
  XOR U35183 ( .A(b[53]), .B(a[103]), .Z(n35005) );
  NANDN U35184 ( .A(n37778), .B(n35005), .Z(n34751) );
  NAND U35185 ( .A(n34752), .B(n34751), .Z(n34985) );
  XOR U35186 ( .A(n34986), .B(n34985), .Z(n34988) );
  XOR U35187 ( .A(n34987), .B(n34988), .Z(n34904) );
  NANDN U35188 ( .A(n36480), .B(n34753), .Z(n34755) );
  XOR U35189 ( .A(a[115]), .B(b[41]), .Z(n34964) );
  NANDN U35190 ( .A(n36594), .B(n34964), .Z(n34754) );
  AND U35191 ( .A(n34755), .B(n34754), .Z(n34926) );
  NANDN U35192 ( .A(n36742), .B(n34756), .Z(n34758) );
  XOR U35193 ( .A(a[113]), .B(b[43]), .Z(n34955) );
  NANDN U35194 ( .A(n36891), .B(n34955), .Z(n34757) );
  AND U35195 ( .A(n34758), .B(n34757), .Z(n34925) );
  NANDN U35196 ( .A(n35936), .B(n34759), .Z(n34761) );
  XOR U35197 ( .A(a[119]), .B(b[37]), .Z(n34970) );
  NANDN U35198 ( .A(n36047), .B(n34970), .Z(n34760) );
  NAND U35199 ( .A(n34761), .B(n34760), .Z(n34924) );
  XOR U35200 ( .A(n34925), .B(n34924), .Z(n34927) );
  XOR U35201 ( .A(n34926), .B(n34927), .Z(n34903) );
  NAND U35202 ( .A(n36490), .B(n34762), .Z(n34764) );
  XNOR U35203 ( .A(a[117]), .B(b[39]), .Z(n34961) );
  NANDN U35204 ( .A(n34961), .B(n36491), .Z(n34763) );
  AND U35205 ( .A(n34764), .B(n34763), .Z(n34902) );
  XOR U35206 ( .A(n34903), .B(n34902), .Z(n34905) );
  XNOR U35207 ( .A(n34904), .B(n34905), .Z(n34946) );
  XNOR U35208 ( .A(n34947), .B(n34946), .Z(n34949) );
  NANDN U35209 ( .A(n34766), .B(n34765), .Z(n34770) );
  OR U35210 ( .A(n34768), .B(n34767), .Z(n34769) );
  AND U35211 ( .A(n34770), .B(n34769), .Z(n35032) );
  NANDN U35212 ( .A(n34772), .B(n34771), .Z(n34776) );
  OR U35213 ( .A(n34774), .B(n34773), .Z(n34775) );
  AND U35214 ( .A(n34776), .B(n34775), .Z(n35030) );
  NANDN U35215 ( .A(n34778), .B(n34777), .Z(n34782) );
  OR U35216 ( .A(n34780), .B(n34779), .Z(n34781) );
  NAND U35217 ( .A(n34782), .B(n34781), .Z(n35029) );
  XNOR U35218 ( .A(n35030), .B(n35029), .Z(n35031) );
  XNOR U35219 ( .A(n35032), .B(n35031), .Z(n34948) );
  XOR U35220 ( .A(n34949), .B(n34948), .Z(n34941) );
  NANDN U35221 ( .A(n34784), .B(n34783), .Z(n34788) );
  NANDN U35222 ( .A(n34786), .B(n34785), .Z(n34787) );
  AND U35223 ( .A(n34788), .B(n34787), .Z(n34898) );
  NANDN U35224 ( .A(n34790), .B(n34789), .Z(n34794) );
  NANDN U35225 ( .A(n34792), .B(n34791), .Z(n34793) );
  AND U35226 ( .A(n34794), .B(n34793), .Z(n34897) );
  NANDN U35227 ( .A(n34796), .B(n34795), .Z(n34800) );
  OR U35228 ( .A(n34798), .B(n34797), .Z(n34799) );
  NAND U35229 ( .A(n34800), .B(n34799), .Z(n34896) );
  XOR U35230 ( .A(n34897), .B(n34896), .Z(n34899) );
  XNOR U35231 ( .A(n34898), .B(n34899), .Z(n34940) );
  XOR U35232 ( .A(n34941), .B(n34940), .Z(n34943) );
  XOR U35233 ( .A(n34942), .B(n34943), .Z(n34885) );
  NANDN U35234 ( .A(n34802), .B(n34801), .Z(n34806) );
  OR U35235 ( .A(n34804), .B(n34803), .Z(n34805) );
  AND U35236 ( .A(n34806), .B(n34805), .Z(n34884) );
  XNOR U35237 ( .A(n34885), .B(n34884), .Z(n34887) );
  NANDN U35238 ( .A(n34808), .B(n34807), .Z(n34812) );
  NAND U35239 ( .A(n34810), .B(n34809), .Z(n34811) );
  AND U35240 ( .A(n34812), .B(n34811), .Z(n34893) );
  NANDN U35241 ( .A(n34814), .B(n34813), .Z(n34818) );
  OR U35242 ( .A(n34816), .B(n34815), .Z(n34817) );
  AND U35243 ( .A(n34818), .B(n34817), .Z(n34891) );
  NANDN U35244 ( .A(n34820), .B(n34819), .Z(n34824) );
  OR U35245 ( .A(n34822), .B(n34821), .Z(n34823) );
  AND U35246 ( .A(n34824), .B(n34823), .Z(n34937) );
  NANDN U35247 ( .A(n34826), .B(n34825), .Z(n34830) );
  OR U35248 ( .A(n34828), .B(n34827), .Z(n34829) );
  AND U35249 ( .A(n34830), .B(n34829), .Z(n34935) );
  NANDN U35250 ( .A(n34832), .B(n34831), .Z(n34836) );
  OR U35251 ( .A(n34834), .B(n34833), .Z(n34835) );
  AND U35252 ( .A(n34836), .B(n34835), .Z(n34931) );
  IV U35253 ( .A(n34857), .Z(n34994) );
  NANDN U35254 ( .A(n34994), .B(n34837), .Z(n34841) );
  NANDN U35255 ( .A(n34839), .B(n34838), .Z(n34840) );
  NAND U35256 ( .A(n34841), .B(n34840), .Z(n34930) );
  XNOR U35257 ( .A(n34931), .B(n34930), .Z(n34933) );
  NANDN U35258 ( .A(n37974), .B(n34842), .Z(n34844) );
  XOR U35259 ( .A(b[57]), .B(a[99]), .Z(n34912) );
  NANDN U35260 ( .A(n38031), .B(n34912), .Z(n34843) );
  AND U35261 ( .A(n34844), .B(n34843), .Z(n35026) );
  NANDN U35262 ( .A(n35260), .B(n34845), .Z(n34847) );
  XOR U35263 ( .A(a[123]), .B(b[33]), .Z(n34952) );
  NANDN U35264 ( .A(n35456), .B(n34952), .Z(n34846) );
  AND U35265 ( .A(n34847), .B(n34846), .Z(n35024) );
  NANDN U35266 ( .A(n37857), .B(n34848), .Z(n34850) );
  XOR U35267 ( .A(b[55]), .B(a[101]), .Z(n35008) );
  NANDN U35268 ( .A(n37911), .B(n35008), .Z(n34849) );
  NAND U35269 ( .A(n34850), .B(n34849), .Z(n35023) );
  XNOR U35270 ( .A(n35024), .B(n35023), .Z(n35025) );
  XNOR U35271 ( .A(n35026), .B(n35025), .Z(n35036) );
  NANDN U35272 ( .A(n38278), .B(n34851), .Z(n34853) );
  XOR U35273 ( .A(b[63]), .B(a[93]), .Z(n34997) );
  NANDN U35274 ( .A(n38279), .B(n34997), .Z(n34852) );
  AND U35275 ( .A(n34853), .B(n34852), .Z(n34919) );
  NANDN U35276 ( .A(n211), .B(n34854), .Z(n34856) );
  XOR U35277 ( .A(b[47]), .B(a[109]), .Z(n34915) );
  NANDN U35278 ( .A(n37172), .B(n34915), .Z(n34855) );
  NAND U35279 ( .A(n34856), .B(n34855), .Z(n34918) );
  XNOR U35280 ( .A(n34919), .B(n34918), .Z(n34921) );
  AND U35281 ( .A(b[63]), .B(a[91]), .Z(n34991) );
  XOR U35282 ( .A(n34991), .B(n34992), .Z(n34993) );
  XOR U35283 ( .A(n34857), .B(n34993), .Z(n34920) );
  XOR U35284 ( .A(n34921), .B(n34920), .Z(n35035) );
  XOR U35285 ( .A(n35036), .B(n35035), .Z(n35038) );
  NANDN U35286 ( .A(n34859), .B(n34858), .Z(n34863) );
  NANDN U35287 ( .A(n34861), .B(n34860), .Z(n34862) );
  NAND U35288 ( .A(n34863), .B(n34862), .Z(n35037) );
  XOR U35289 ( .A(n35038), .B(n35037), .Z(n34932) );
  XOR U35290 ( .A(n34933), .B(n34932), .Z(n34934) );
  XNOR U35291 ( .A(n34935), .B(n34934), .Z(n34936) );
  XNOR U35292 ( .A(n34937), .B(n34936), .Z(n34890) );
  XNOR U35293 ( .A(n34891), .B(n34890), .Z(n34892) );
  XNOR U35294 ( .A(n34893), .B(n34892), .Z(n34886) );
  XOR U35295 ( .A(n34887), .B(n34886), .Z(n34879) );
  NANDN U35296 ( .A(n34865), .B(n34864), .Z(n34869) );
  NANDN U35297 ( .A(n34867), .B(n34866), .Z(n34868) );
  AND U35298 ( .A(n34869), .B(n34868), .Z(n34878) );
  XOR U35299 ( .A(n34879), .B(n34878), .Z(n34881) );
  XNOR U35300 ( .A(n34880), .B(n34881), .Z(n34872) );
  XOR U35301 ( .A(n34873), .B(n34872), .Z(n34875) );
  XNOR U35302 ( .A(n34874), .B(n34875), .Z(n34870) );
  XOR U35303 ( .A(n34871), .B(n34870), .Z(c[219]) );
  AND U35304 ( .A(n34871), .B(n34870), .Z(n35048) );
  NANDN U35305 ( .A(n34873), .B(n34872), .Z(n34877) );
  OR U35306 ( .A(n34875), .B(n34874), .Z(n34876) );
  AND U35307 ( .A(n34877), .B(n34876), .Z(n35051) );
  NANDN U35308 ( .A(n34879), .B(n34878), .Z(n34883) );
  NANDN U35309 ( .A(n34881), .B(n34880), .Z(n34882) );
  AND U35310 ( .A(n34883), .B(n34882), .Z(n35050) );
  NANDN U35311 ( .A(n34885), .B(n34884), .Z(n34889) );
  NAND U35312 ( .A(n34887), .B(n34886), .Z(n34888) );
  AND U35313 ( .A(n34889), .B(n34888), .Z(n35057) );
  NANDN U35314 ( .A(n34891), .B(n34890), .Z(n34895) );
  NANDN U35315 ( .A(n34893), .B(n34892), .Z(n34894) );
  AND U35316 ( .A(n34895), .B(n34894), .Z(n35056) );
  NANDN U35317 ( .A(n34897), .B(n34896), .Z(n34901) );
  NANDN U35318 ( .A(n34899), .B(n34898), .Z(n34900) );
  AND U35319 ( .A(n34901), .B(n34900), .Z(n35069) );
  NANDN U35320 ( .A(n34903), .B(n34902), .Z(n34907) );
  OR U35321 ( .A(n34905), .B(n34904), .Z(n34906) );
  AND U35322 ( .A(n34907), .B(n34906), .Z(n35080) );
  NANDN U35323 ( .A(n34909), .B(n34908), .Z(n34911) );
  XOR U35324 ( .A(a[126]), .B(b[31]), .Z(n35146) );
  NANDN U35325 ( .A(n35145), .B(n35146), .Z(n34910) );
  AND U35326 ( .A(n34911), .B(n34910), .Z(n35169) );
  NANDN U35327 ( .A(n37974), .B(n34912), .Z(n34914) );
  XOR U35328 ( .A(b[57]), .B(a[100]), .Z(n35182) );
  NANDN U35329 ( .A(n38031), .B(n35182), .Z(n34913) );
  AND U35330 ( .A(n34914), .B(n34913), .Z(n35168) );
  NANDN U35331 ( .A(n211), .B(n34915), .Z(n34917) );
  XOR U35332 ( .A(b[47]), .B(a[110]), .Z(n35149) );
  NANDN U35333 ( .A(n37172), .B(n35149), .Z(n34916) );
  NAND U35334 ( .A(n34917), .B(n34916), .Z(n35167) );
  XOR U35335 ( .A(n35168), .B(n35167), .Z(n35170) );
  XOR U35336 ( .A(n35169), .B(n35170), .Z(n35086) );
  NANDN U35337 ( .A(n34919), .B(n34918), .Z(n34923) );
  NAND U35338 ( .A(n34921), .B(n34920), .Z(n34922) );
  AND U35339 ( .A(n34923), .B(n34922), .Z(n35085) );
  XNOR U35340 ( .A(n35086), .B(n35085), .Z(n35087) );
  NANDN U35341 ( .A(n34925), .B(n34924), .Z(n34929) );
  OR U35342 ( .A(n34927), .B(n34926), .Z(n34928) );
  NAND U35343 ( .A(n34929), .B(n34928), .Z(n35088) );
  XNOR U35344 ( .A(n35087), .B(n35088), .Z(n35079) );
  XNOR U35345 ( .A(n35080), .B(n35079), .Z(n35081) );
  XNOR U35346 ( .A(n35081), .B(n35082), .Z(n35067) );
  NANDN U35347 ( .A(n34935), .B(n34934), .Z(n34939) );
  NANDN U35348 ( .A(n34937), .B(n34936), .Z(n34938) );
  NAND U35349 ( .A(n34939), .B(n34938), .Z(n35068) );
  XOR U35350 ( .A(n35067), .B(n35068), .Z(n35070) );
  XOR U35351 ( .A(n35069), .B(n35070), .Z(n35064) );
  NANDN U35352 ( .A(n34941), .B(n34940), .Z(n34945) );
  OR U35353 ( .A(n34943), .B(n34942), .Z(n34944) );
  AND U35354 ( .A(n34945), .B(n34944), .Z(n35061) );
  NANDN U35355 ( .A(n34947), .B(n34946), .Z(n34951) );
  NAND U35356 ( .A(n34949), .B(n34948), .Z(n34950) );
  AND U35357 ( .A(n34951), .B(n34950), .Z(n35133) );
  NANDN U35358 ( .A(n35260), .B(n34952), .Z(n34954) );
  XOR U35359 ( .A(a[124]), .B(b[33]), .Z(n35155) );
  NANDN U35360 ( .A(n35456), .B(n35155), .Z(n34953) );
  AND U35361 ( .A(n34954), .B(n34953), .Z(n35193) );
  NANDN U35362 ( .A(n36742), .B(n34955), .Z(n34957) );
  XOR U35363 ( .A(a[114]), .B(b[43]), .Z(n35124) );
  NANDN U35364 ( .A(n36891), .B(n35124), .Z(n34956) );
  AND U35365 ( .A(n34957), .B(n34956), .Z(n35192) );
  NANDN U35366 ( .A(n37526), .B(n34958), .Z(n34960) );
  XOR U35367 ( .A(b[51]), .B(a[106]), .Z(n35127) );
  NANDN U35368 ( .A(n37605), .B(n35127), .Z(n34959) );
  NAND U35369 ( .A(n34960), .B(n34959), .Z(n35191) );
  XOR U35370 ( .A(n35192), .B(n35191), .Z(n35194) );
  XOR U35371 ( .A(n35193), .B(n35194), .Z(n35093) );
  NANDN U35372 ( .A(n34961), .B(n36490), .Z(n34963) );
  XOR U35373 ( .A(a[118]), .B(b[39]), .Z(n35179) );
  NANDN U35374 ( .A(n36347), .B(n35179), .Z(n34962) );
  AND U35375 ( .A(n34963), .B(n34962), .Z(n35163) );
  NANDN U35376 ( .A(n36480), .B(n34964), .Z(n34966) );
  XOR U35377 ( .A(a[116]), .B(b[41]), .Z(n35121) );
  NANDN U35378 ( .A(n36594), .B(n35121), .Z(n34965) );
  AND U35379 ( .A(n34966), .B(n34965), .Z(n35162) );
  NANDN U35380 ( .A(n35611), .B(n34967), .Z(n34969) );
  XOR U35381 ( .A(a[122]), .B(b[35]), .Z(n35152) );
  NANDN U35382 ( .A(n35801), .B(n35152), .Z(n34968) );
  NAND U35383 ( .A(n34969), .B(n34968), .Z(n35161) );
  XOR U35384 ( .A(n35162), .B(n35161), .Z(n35164) );
  XOR U35385 ( .A(n35163), .B(n35164), .Z(n35092) );
  NAND U35386 ( .A(n36238), .B(n34970), .Z(n34972) );
  XNOR U35387 ( .A(a[120]), .B(b[37]), .Z(n35185) );
  NANDN U35388 ( .A(n35185), .B(n36239), .Z(n34971) );
  AND U35389 ( .A(n34972), .B(n34971), .Z(n35091) );
  XOR U35390 ( .A(n35092), .B(n35091), .Z(n35094) );
  XOR U35391 ( .A(n35093), .B(n35094), .Z(n35199) );
  NANDN U35392 ( .A(n34974), .B(n34973), .Z(n34978) );
  OR U35393 ( .A(n34976), .B(n34975), .Z(n34977) );
  AND U35394 ( .A(n34978), .B(n34977), .Z(n35198) );
  NANDN U35395 ( .A(n34980), .B(n34979), .Z(n34984) );
  OR U35396 ( .A(n34982), .B(n34981), .Z(n34983) );
  NAND U35397 ( .A(n34984), .B(n34983), .Z(n35197) );
  XOR U35398 ( .A(n35198), .B(n35197), .Z(n35200) );
  XOR U35399 ( .A(n35199), .B(n35200), .Z(n35138) );
  NANDN U35400 ( .A(n34986), .B(n34985), .Z(n34990) );
  OR U35401 ( .A(n34988), .B(n34987), .Z(n34989) );
  AND U35402 ( .A(n34990), .B(n34989), .Z(n35211) );
  NANDN U35403 ( .A(n34992), .B(n34991), .Z(n34996) );
  ANDN U35404 ( .B(n34994), .A(n34993), .Z(n34995) );
  ANDN U35405 ( .B(n34996), .A(n34995), .Z(n35210) );
  NANDN U35406 ( .A(n38278), .B(n34997), .Z(n34999) );
  XOR U35407 ( .A(b[63]), .B(a[94]), .Z(n35114) );
  NANDN U35408 ( .A(n38279), .B(n35114), .Z(n34998) );
  AND U35409 ( .A(n34999), .B(n34998), .Z(n35105) );
  NAND U35410 ( .A(b[63]), .B(a[92]), .Z(n35120) );
  ANDN U35411 ( .B(n35001), .A(n35000), .Z(n35004) );
  NAND U35412 ( .A(b[29]), .B(n35002), .Z(n35003) );
  NANDN U35413 ( .A(n35004), .B(n35003), .Z(n35103) );
  XOR U35414 ( .A(n35120), .B(n35103), .Z(n35104) );
  XNOR U35415 ( .A(n35105), .B(n35104), .Z(n35209) );
  XOR U35416 ( .A(n35210), .B(n35209), .Z(n35212) );
  XOR U35417 ( .A(n35211), .B(n35212), .Z(n35137) );
  NANDN U35418 ( .A(n37705), .B(n35005), .Z(n35007) );
  XOR U35419 ( .A(b[53]), .B(a[104]), .Z(n35173) );
  NANDN U35420 ( .A(n37778), .B(n35173), .Z(n35006) );
  AND U35421 ( .A(n35007), .B(n35006), .Z(n35099) );
  NANDN U35422 ( .A(n37857), .B(n35008), .Z(n35010) );
  XOR U35423 ( .A(b[55]), .B(a[102]), .Z(n35176) );
  NANDN U35424 ( .A(n37911), .B(n35176), .Z(n35009) );
  AND U35425 ( .A(n35010), .B(n35009), .Z(n35098) );
  NANDN U35426 ( .A(n36991), .B(n35011), .Z(n35013) );
  XOR U35427 ( .A(a[112]), .B(b[45]), .Z(n35158) );
  NANDN U35428 ( .A(n37083), .B(n35158), .Z(n35012) );
  NAND U35429 ( .A(n35013), .B(n35012), .Z(n35097) );
  XOR U35430 ( .A(n35098), .B(n35097), .Z(n35100) );
  XOR U35431 ( .A(n35099), .B(n35100), .Z(n35204) );
  NANDN U35432 ( .A(n38090), .B(n35014), .Z(n35016) );
  XOR U35433 ( .A(b[59]), .B(a[98]), .Z(n35188) );
  NANDN U35434 ( .A(n38130), .B(n35188), .Z(n35015) );
  AND U35435 ( .A(n35016), .B(n35015), .Z(n35110) );
  NANDN U35436 ( .A(n38247), .B(n35017), .Z(n35019) );
  XOR U35437 ( .A(b[61]), .B(a[96]), .Z(n35142) );
  NANDN U35438 ( .A(n38248), .B(n35142), .Z(n35018) );
  AND U35439 ( .A(n35019), .B(n35018), .Z(n35109) );
  NANDN U35440 ( .A(n212), .B(n35020), .Z(n35022) );
  XOR U35441 ( .A(b[49]), .B(a[108]), .Z(n35117) );
  NANDN U35442 ( .A(n37432), .B(n35117), .Z(n35021) );
  NAND U35443 ( .A(n35022), .B(n35021), .Z(n35108) );
  XOR U35444 ( .A(n35109), .B(n35108), .Z(n35111) );
  XNOR U35445 ( .A(n35110), .B(n35111), .Z(n35203) );
  XNOR U35446 ( .A(n35204), .B(n35203), .Z(n35205) );
  NANDN U35447 ( .A(n35024), .B(n35023), .Z(n35028) );
  NANDN U35448 ( .A(n35026), .B(n35025), .Z(n35027) );
  NAND U35449 ( .A(n35028), .B(n35027), .Z(n35206) );
  XNOR U35450 ( .A(n35205), .B(n35206), .Z(n35136) );
  XOR U35451 ( .A(n35137), .B(n35136), .Z(n35139) );
  XOR U35452 ( .A(n35138), .B(n35139), .Z(n35131) );
  NANDN U35453 ( .A(n35030), .B(n35029), .Z(n35034) );
  NANDN U35454 ( .A(n35032), .B(n35031), .Z(n35033) );
  AND U35455 ( .A(n35034), .B(n35033), .Z(n35076) );
  NAND U35456 ( .A(n35036), .B(n35035), .Z(n35040) );
  NAND U35457 ( .A(n35038), .B(n35037), .Z(n35039) );
  AND U35458 ( .A(n35040), .B(n35039), .Z(n35074) );
  NANDN U35459 ( .A(n35042), .B(n35041), .Z(n35046) );
  NAND U35460 ( .A(n35044), .B(n35043), .Z(n35045) );
  AND U35461 ( .A(n35046), .B(n35045), .Z(n35073) );
  XNOR U35462 ( .A(n35074), .B(n35073), .Z(n35075) );
  XNOR U35463 ( .A(n35076), .B(n35075), .Z(n35130) );
  XNOR U35464 ( .A(n35131), .B(n35130), .Z(n35132) );
  XOR U35465 ( .A(n35133), .B(n35132), .Z(n35062) );
  XNOR U35466 ( .A(n35061), .B(n35062), .Z(n35063) );
  XNOR U35467 ( .A(n35064), .B(n35063), .Z(n35055) );
  XOR U35468 ( .A(n35056), .B(n35055), .Z(n35058) );
  XNOR U35469 ( .A(n35057), .B(n35058), .Z(n35049) );
  XOR U35470 ( .A(n35050), .B(n35049), .Z(n35052) );
  XNOR U35471 ( .A(n35051), .B(n35052), .Z(n35047) );
  XOR U35472 ( .A(n35048), .B(n35047), .Z(c[220]) );
  AND U35473 ( .A(n35048), .B(n35047), .Z(n35216) );
  NANDN U35474 ( .A(n35050), .B(n35049), .Z(n35054) );
  OR U35475 ( .A(n35052), .B(n35051), .Z(n35053) );
  AND U35476 ( .A(n35054), .B(n35053), .Z(n35219) );
  NANDN U35477 ( .A(n35056), .B(n35055), .Z(n35060) );
  OR U35478 ( .A(n35058), .B(n35057), .Z(n35059) );
  AND U35479 ( .A(n35060), .B(n35059), .Z(n35217) );
  NANDN U35480 ( .A(n35062), .B(n35061), .Z(n35066) );
  NANDN U35481 ( .A(n35064), .B(n35063), .Z(n35065) );
  AND U35482 ( .A(n35066), .B(n35065), .Z(n35225) );
  NANDN U35483 ( .A(n35068), .B(n35067), .Z(n35072) );
  OR U35484 ( .A(n35070), .B(n35069), .Z(n35071) );
  AND U35485 ( .A(n35072), .B(n35071), .Z(n35224) );
  NANDN U35486 ( .A(n35074), .B(n35073), .Z(n35078) );
  NANDN U35487 ( .A(n35076), .B(n35075), .Z(n35077) );
  AND U35488 ( .A(n35078), .B(n35077), .Z(n35380) );
  NANDN U35489 ( .A(n35080), .B(n35079), .Z(n35084) );
  NANDN U35490 ( .A(n35082), .B(n35081), .Z(n35083) );
  AND U35491 ( .A(n35084), .B(n35083), .Z(n35377) );
  NANDN U35492 ( .A(n35086), .B(n35085), .Z(n35090) );
  NANDN U35493 ( .A(n35088), .B(n35087), .Z(n35089) );
  AND U35494 ( .A(n35090), .B(n35089), .Z(n35243) );
  NANDN U35495 ( .A(n35092), .B(n35091), .Z(n35096) );
  OR U35496 ( .A(n35094), .B(n35093), .Z(n35095) );
  AND U35497 ( .A(n35096), .B(n35095), .Z(n35241) );
  NANDN U35498 ( .A(n35098), .B(n35097), .Z(n35102) );
  OR U35499 ( .A(n35100), .B(n35099), .Z(n35101) );
  AND U35500 ( .A(n35102), .B(n35101), .Z(n35354) );
  IV U35501 ( .A(n35120), .Z(n35343) );
  NANDN U35502 ( .A(n35343), .B(n35103), .Z(n35107) );
  NANDN U35503 ( .A(n35105), .B(n35104), .Z(n35106) );
  NAND U35504 ( .A(n35107), .B(n35106), .Z(n35353) );
  XNOR U35505 ( .A(n35354), .B(n35353), .Z(n35355) );
  NANDN U35506 ( .A(n35109), .B(n35108), .Z(n35113) );
  OR U35507 ( .A(n35111), .B(n35110), .Z(n35112) );
  AND U35508 ( .A(n35113), .B(n35112), .Z(n35275) );
  NANDN U35509 ( .A(n38278), .B(n35114), .Z(n35116) );
  XOR U35510 ( .A(b[63]), .B(a[95]), .Z(n35305) );
  NANDN U35511 ( .A(n38279), .B(n35305), .Z(n35115) );
  AND U35512 ( .A(n35116), .B(n35115), .Z(n35288) );
  NANDN U35513 ( .A(n212), .B(n35117), .Z(n35119) );
  XOR U35514 ( .A(b[49]), .B(a[109]), .Z(n35263) );
  NANDN U35515 ( .A(n37432), .B(n35263), .Z(n35118) );
  NAND U35516 ( .A(n35119), .B(n35118), .Z(n35287) );
  XNOR U35517 ( .A(n35288), .B(n35287), .Z(n35289) );
  AND U35518 ( .A(b[63]), .B(a[93]), .Z(n35341) );
  XNOR U35519 ( .A(n35340), .B(n35341), .Z(n35342) );
  XOR U35520 ( .A(n35120), .B(n35342), .Z(n35290) );
  XOR U35521 ( .A(n35289), .B(n35290), .Z(n35272) );
  NANDN U35522 ( .A(n36480), .B(n35121), .Z(n35123) );
  XOR U35523 ( .A(a[117]), .B(b[41]), .Z(n35253) );
  NANDN U35524 ( .A(n36594), .B(n35253), .Z(n35122) );
  AND U35525 ( .A(n35123), .B(n35122), .Z(n35337) );
  NANDN U35526 ( .A(n36742), .B(n35124), .Z(n35126) );
  XOR U35527 ( .A(a[115]), .B(b[43]), .Z(n35319) );
  NANDN U35528 ( .A(n36891), .B(n35319), .Z(n35125) );
  AND U35529 ( .A(n35126), .B(n35125), .Z(n35335) );
  NANDN U35530 ( .A(n37526), .B(n35127), .Z(n35129) );
  XOR U35531 ( .A(b[51]), .B(a[107]), .Z(n35284) );
  NANDN U35532 ( .A(n37605), .B(n35284), .Z(n35128) );
  NAND U35533 ( .A(n35129), .B(n35128), .Z(n35334) );
  XNOR U35534 ( .A(n35335), .B(n35334), .Z(n35336) );
  XOR U35535 ( .A(n35337), .B(n35336), .Z(n35273) );
  XNOR U35536 ( .A(n35272), .B(n35273), .Z(n35274) );
  XOR U35537 ( .A(n35275), .B(n35274), .Z(n35356) );
  XOR U35538 ( .A(n35355), .B(n35356), .Z(n35242) );
  XOR U35539 ( .A(n35241), .B(n35242), .Z(n35244) );
  XOR U35540 ( .A(n35243), .B(n35244), .Z(n35378) );
  XNOR U35541 ( .A(n35377), .B(n35378), .Z(n35379) );
  XNOR U35542 ( .A(n35380), .B(n35379), .Z(n35232) );
  NANDN U35543 ( .A(n35131), .B(n35130), .Z(n35135) );
  NANDN U35544 ( .A(n35133), .B(n35132), .Z(n35134) );
  AND U35545 ( .A(n35135), .B(n35134), .Z(n35230) );
  NANDN U35546 ( .A(n35137), .B(n35136), .Z(n35141) );
  OR U35547 ( .A(n35139), .B(n35138), .Z(n35140) );
  AND U35548 ( .A(n35141), .B(n35140), .Z(n35373) );
  NANDN U35549 ( .A(n38247), .B(n35142), .Z(n35144) );
  XOR U35550 ( .A(b[61]), .B(a[97]), .Z(n35256) );
  NANDN U35551 ( .A(n38248), .B(n35256), .Z(n35143) );
  AND U35552 ( .A(n35144), .B(n35143), .Z(n35330) );
  XNOR U35553 ( .A(a[127]), .B(b[31]), .Z(n35308) );
  OR U35554 ( .A(n35308), .B(n35145), .Z(n35148) );
  NAND U35555 ( .A(n35309), .B(n35146), .Z(n35147) );
  AND U35556 ( .A(n35148), .B(n35147), .Z(n35329) );
  NANDN U35557 ( .A(n211), .B(n35149), .Z(n35151) );
  XOR U35558 ( .A(b[47]), .B(a[111]), .Z(n35316) );
  NANDN U35559 ( .A(n37172), .B(n35316), .Z(n35150) );
  NAND U35560 ( .A(n35151), .B(n35150), .Z(n35328) );
  XOR U35561 ( .A(n35329), .B(n35328), .Z(n35331) );
  XOR U35562 ( .A(n35330), .B(n35331), .Z(n35366) );
  NANDN U35563 ( .A(n35611), .B(n35152), .Z(n35154) );
  XOR U35564 ( .A(a[123]), .B(b[35]), .Z(n35281) );
  NANDN U35565 ( .A(n35801), .B(n35281), .Z(n35153) );
  AND U35566 ( .A(n35154), .B(n35153), .Z(n35295) );
  NANDN U35567 ( .A(n35260), .B(n35155), .Z(n35157) );
  XOR U35568 ( .A(a[125]), .B(b[33]), .Z(n35259) );
  NANDN U35569 ( .A(n35456), .B(n35259), .Z(n35156) );
  AND U35570 ( .A(n35157), .B(n35156), .Z(n35294) );
  NANDN U35571 ( .A(n36991), .B(n35158), .Z(n35160) );
  XOR U35572 ( .A(a[113]), .B(b[45]), .Z(n35313) );
  NANDN U35573 ( .A(n37083), .B(n35313), .Z(n35159) );
  NAND U35574 ( .A(n35160), .B(n35159), .Z(n35293) );
  XOR U35575 ( .A(n35294), .B(n35293), .Z(n35296) );
  XNOR U35576 ( .A(n35295), .B(n35296), .Z(n35365) );
  XNOR U35577 ( .A(n35366), .B(n35365), .Z(n35367) );
  NANDN U35578 ( .A(n35162), .B(n35161), .Z(n35166) );
  OR U35579 ( .A(n35164), .B(n35163), .Z(n35165) );
  NAND U35580 ( .A(n35166), .B(n35165), .Z(n35368) );
  XNOR U35581 ( .A(n35367), .B(n35368), .Z(n35299) );
  NANDN U35582 ( .A(n35168), .B(n35167), .Z(n35172) );
  OR U35583 ( .A(n35170), .B(n35169), .Z(n35171) );
  NAND U35584 ( .A(n35172), .B(n35171), .Z(n35300) );
  XNOR U35585 ( .A(n35299), .B(n35300), .Z(n35301) );
  NANDN U35586 ( .A(n37705), .B(n35173), .Z(n35175) );
  XOR U35587 ( .A(b[53]), .B(a[105]), .Z(n35247) );
  NANDN U35588 ( .A(n37778), .B(n35247), .Z(n35174) );
  AND U35589 ( .A(n35175), .B(n35174), .Z(n35324) );
  NANDN U35590 ( .A(n37857), .B(n35176), .Z(n35178) );
  XOR U35591 ( .A(b[55]), .B(a[103]), .Z(n35350) );
  NANDN U35592 ( .A(n37911), .B(n35350), .Z(n35177) );
  AND U35593 ( .A(n35178), .B(n35177), .Z(n35323) );
  NANDN U35594 ( .A(n36210), .B(n35179), .Z(n35181) );
  XOR U35595 ( .A(a[119]), .B(b[39]), .Z(n35347) );
  NANDN U35596 ( .A(n36347), .B(n35347), .Z(n35180) );
  NAND U35597 ( .A(n35181), .B(n35180), .Z(n35322) );
  XOR U35598 ( .A(n35323), .B(n35322), .Z(n35325) );
  XOR U35599 ( .A(n35324), .B(n35325), .Z(n35360) );
  NANDN U35600 ( .A(n37974), .B(n35182), .Z(n35184) );
  XOR U35601 ( .A(b[57]), .B(a[101]), .Z(n35250) );
  NANDN U35602 ( .A(n38031), .B(n35250), .Z(n35183) );
  AND U35603 ( .A(n35184), .B(n35183), .Z(n35268) );
  NANDN U35604 ( .A(n35185), .B(n36238), .Z(n35187) );
  XOR U35605 ( .A(a[121]), .B(b[37]), .Z(n35278) );
  NANDN U35606 ( .A(n36047), .B(n35278), .Z(n35186) );
  AND U35607 ( .A(n35187), .B(n35186), .Z(n35267) );
  NANDN U35608 ( .A(n38090), .B(n35188), .Z(n35190) );
  XOR U35609 ( .A(b[59]), .B(a[99]), .Z(n35344) );
  NANDN U35610 ( .A(n38130), .B(n35344), .Z(n35189) );
  NAND U35611 ( .A(n35190), .B(n35189), .Z(n35266) );
  XOR U35612 ( .A(n35267), .B(n35266), .Z(n35269) );
  XNOR U35613 ( .A(n35268), .B(n35269), .Z(n35359) );
  XNOR U35614 ( .A(n35360), .B(n35359), .Z(n35361) );
  NANDN U35615 ( .A(n35192), .B(n35191), .Z(n35196) );
  OR U35616 ( .A(n35194), .B(n35193), .Z(n35195) );
  NAND U35617 ( .A(n35196), .B(n35195), .Z(n35362) );
  XOR U35618 ( .A(n35361), .B(n35362), .Z(n35302) );
  XNOR U35619 ( .A(n35301), .B(n35302), .Z(n35371) );
  NANDN U35620 ( .A(n35198), .B(n35197), .Z(n35202) );
  OR U35621 ( .A(n35200), .B(n35199), .Z(n35201) );
  AND U35622 ( .A(n35202), .B(n35201), .Z(n35237) );
  NANDN U35623 ( .A(n35204), .B(n35203), .Z(n35208) );
  NANDN U35624 ( .A(n35206), .B(n35205), .Z(n35207) );
  AND U35625 ( .A(n35208), .B(n35207), .Z(n35236) );
  NANDN U35626 ( .A(n35210), .B(n35209), .Z(n35214) );
  OR U35627 ( .A(n35212), .B(n35211), .Z(n35213) );
  AND U35628 ( .A(n35214), .B(n35213), .Z(n35235) );
  XOR U35629 ( .A(n35236), .B(n35235), .Z(n35238) );
  XOR U35630 ( .A(n35237), .B(n35238), .Z(n35372) );
  XOR U35631 ( .A(n35371), .B(n35372), .Z(n35374) );
  XNOR U35632 ( .A(n35373), .B(n35374), .Z(n35229) );
  XNOR U35633 ( .A(n35230), .B(n35229), .Z(n35231) );
  XNOR U35634 ( .A(n35232), .B(n35231), .Z(n35223) );
  XOR U35635 ( .A(n35224), .B(n35223), .Z(n35226) );
  XOR U35636 ( .A(n35225), .B(n35226), .Z(n35218) );
  XOR U35637 ( .A(n35217), .B(n35218), .Z(n35220) );
  XNOR U35638 ( .A(n35219), .B(n35220), .Z(n35215) );
  XOR U35639 ( .A(n35216), .B(n35215), .Z(c[221]) );
  AND U35640 ( .A(n35216), .B(n35215), .Z(n35384) );
  NANDN U35641 ( .A(n35218), .B(n35217), .Z(n35222) );
  OR U35642 ( .A(n35220), .B(n35219), .Z(n35221) );
  AND U35643 ( .A(n35222), .B(n35221), .Z(n35387) );
  NANDN U35644 ( .A(n35224), .B(n35223), .Z(n35228) );
  NANDN U35645 ( .A(n35226), .B(n35225), .Z(n35227) );
  AND U35646 ( .A(n35228), .B(n35227), .Z(n35386) );
  NANDN U35647 ( .A(n35230), .B(n35229), .Z(n35234) );
  NAND U35648 ( .A(n35232), .B(n35231), .Z(n35233) );
  AND U35649 ( .A(n35234), .B(n35233), .Z(n35394) );
  NANDN U35650 ( .A(n35236), .B(n35235), .Z(n35240) );
  NANDN U35651 ( .A(n35238), .B(n35237), .Z(n35239) );
  AND U35652 ( .A(n35240), .B(n35239), .Z(n35532) );
  NANDN U35653 ( .A(n35242), .B(n35241), .Z(n35246) );
  NANDN U35654 ( .A(n35244), .B(n35243), .Z(n35245) );
  AND U35655 ( .A(n35246), .B(n35245), .Z(n35530) );
  NANDN U35656 ( .A(n37705), .B(n35247), .Z(n35249) );
  XOR U35657 ( .A(b[53]), .B(a[106]), .Z(n35496) );
  NANDN U35658 ( .A(n37778), .B(n35496), .Z(n35248) );
  AND U35659 ( .A(n35249), .B(n35248), .Z(n35443) );
  NANDN U35660 ( .A(n37974), .B(n35250), .Z(n35252) );
  XOR U35661 ( .A(b[57]), .B(a[102]), .Z(n35478) );
  NANDN U35662 ( .A(n38031), .B(n35478), .Z(n35251) );
  AND U35663 ( .A(n35252), .B(n35251), .Z(n35442) );
  NANDN U35664 ( .A(n36480), .B(n35253), .Z(n35255) );
  XOR U35665 ( .A(a[118]), .B(b[41]), .Z(n35447) );
  NANDN U35666 ( .A(n36594), .B(n35447), .Z(n35254) );
  NAND U35667 ( .A(n35255), .B(n35254), .Z(n35441) );
  XOR U35668 ( .A(n35442), .B(n35441), .Z(n35444) );
  XOR U35669 ( .A(n35443), .B(n35444), .Z(n35436) );
  NANDN U35670 ( .A(n38247), .B(n35256), .Z(n35258) );
  XOR U35671 ( .A(b[61]), .B(a[98]), .Z(n35490) );
  NANDN U35672 ( .A(n38248), .B(n35490), .Z(n35257) );
  AND U35673 ( .A(n35258), .B(n35257), .Z(n35486) );
  NANDN U35674 ( .A(n35260), .B(n35259), .Z(n35262) );
  XOR U35675 ( .A(a[126]), .B(b[33]), .Z(n35457) );
  NANDN U35676 ( .A(n35456), .B(n35457), .Z(n35261) );
  AND U35677 ( .A(n35262), .B(n35261), .Z(n35485) );
  NANDN U35678 ( .A(n212), .B(n35263), .Z(n35265) );
  XOR U35679 ( .A(b[49]), .B(a[110]), .Z(n35460) );
  NANDN U35680 ( .A(n37432), .B(n35460), .Z(n35264) );
  NAND U35681 ( .A(n35265), .B(n35264), .Z(n35484) );
  XOR U35682 ( .A(n35485), .B(n35484), .Z(n35487) );
  XNOR U35683 ( .A(n35486), .B(n35487), .Z(n35435) );
  XNOR U35684 ( .A(n35436), .B(n35435), .Z(n35437) );
  NANDN U35685 ( .A(n35267), .B(n35266), .Z(n35271) );
  OR U35686 ( .A(n35269), .B(n35268), .Z(n35270) );
  NAND U35687 ( .A(n35271), .B(n35270), .Z(n35438) );
  XNOR U35688 ( .A(n35437), .B(n35438), .Z(n35405) );
  NANDN U35689 ( .A(n35273), .B(n35272), .Z(n35277) );
  NANDN U35690 ( .A(n35275), .B(n35274), .Z(n35276) );
  NAND U35691 ( .A(n35277), .B(n35276), .Z(n35406) );
  XNOR U35692 ( .A(n35405), .B(n35406), .Z(n35407) );
  NANDN U35693 ( .A(n35936), .B(n35278), .Z(n35280) );
  XOR U35694 ( .A(a[122]), .B(b[37]), .Z(n35493) );
  NANDN U35695 ( .A(n36047), .B(n35493), .Z(n35279) );
  AND U35696 ( .A(n35280), .B(n35279), .Z(n35465) );
  NANDN U35697 ( .A(n35611), .B(n35281), .Z(n35283) );
  XOR U35698 ( .A(a[124]), .B(b[35]), .Z(n35499) );
  NANDN U35699 ( .A(n35801), .B(n35499), .Z(n35282) );
  AND U35700 ( .A(n35283), .B(n35282), .Z(n35464) );
  NANDN U35701 ( .A(n37526), .B(n35284), .Z(n35286) );
  XOR U35702 ( .A(b[51]), .B(a[108]), .Z(n35505) );
  NANDN U35703 ( .A(n37605), .B(n35505), .Z(n35285) );
  NAND U35704 ( .A(n35286), .B(n35285), .Z(n35463) );
  XOR U35705 ( .A(n35464), .B(n35463), .Z(n35466) );
  XOR U35706 ( .A(n35465), .B(n35466), .Z(n35420) );
  NANDN U35707 ( .A(n35288), .B(n35287), .Z(n35292) );
  NAND U35708 ( .A(n35290), .B(n35289), .Z(n35291) );
  AND U35709 ( .A(n35292), .B(n35291), .Z(n35417) );
  NANDN U35710 ( .A(n35294), .B(n35293), .Z(n35298) );
  OR U35711 ( .A(n35296), .B(n35295), .Z(n35297) );
  NAND U35712 ( .A(n35298), .B(n35297), .Z(n35418) );
  XNOR U35713 ( .A(n35417), .B(n35418), .Z(n35419) );
  XOR U35714 ( .A(n35420), .B(n35419), .Z(n35408) );
  XOR U35715 ( .A(n35407), .B(n35408), .Z(n35531) );
  XOR U35716 ( .A(n35530), .B(n35531), .Z(n35533) );
  XOR U35717 ( .A(n35532), .B(n35533), .Z(n35398) );
  NANDN U35718 ( .A(n35300), .B(n35299), .Z(n35304) );
  NANDN U35719 ( .A(n35302), .B(n35301), .Z(n35303) );
  AND U35720 ( .A(n35304), .B(n35303), .Z(n35529) );
  NANDN U35721 ( .A(n38278), .B(n35305), .Z(n35307) );
  XOR U35722 ( .A(b[63]), .B(a[96]), .Z(n35502) );
  NANDN U35723 ( .A(n38279), .B(n35502), .Z(n35306) );
  AND U35724 ( .A(n35307), .B(n35306), .Z(n35511) );
  NAND U35725 ( .A(b[63]), .B(a[94]), .Z(n35508) );
  ANDN U35726 ( .B(n35309), .A(n35308), .Z(n35312) );
  NAND U35727 ( .A(b[31]), .B(n35310), .Z(n35311) );
  NANDN U35728 ( .A(n35312), .B(n35311), .Z(n35509) );
  XOR U35729 ( .A(n35508), .B(n35509), .Z(n35510) );
  XOR U35730 ( .A(n35511), .B(n35510), .Z(n35425) );
  NANDN U35731 ( .A(n36991), .B(n35313), .Z(n35315) );
  XOR U35732 ( .A(a[114]), .B(b[45]), .Z(n35472) );
  NANDN U35733 ( .A(n37083), .B(n35472), .Z(n35314) );
  AND U35734 ( .A(n35315), .B(n35314), .Z(n35516) );
  NANDN U35735 ( .A(n211), .B(n35316), .Z(n35318) );
  XOR U35736 ( .A(b[47]), .B(a[112]), .Z(n35469) );
  NANDN U35737 ( .A(n37172), .B(n35469), .Z(n35317) );
  AND U35738 ( .A(n35318), .B(n35317), .Z(n35515) );
  NANDN U35739 ( .A(n36742), .B(n35319), .Z(n35321) );
  XOR U35740 ( .A(a[116]), .B(b[43]), .Z(n35481) );
  NANDN U35741 ( .A(n36891), .B(n35481), .Z(n35320) );
  NAND U35742 ( .A(n35321), .B(n35320), .Z(n35514) );
  XOR U35743 ( .A(n35515), .B(n35514), .Z(n35517) );
  XOR U35744 ( .A(n35516), .B(n35517), .Z(n35424) );
  NANDN U35745 ( .A(n35323), .B(n35322), .Z(n35327) );
  OR U35746 ( .A(n35325), .B(n35324), .Z(n35326) );
  AND U35747 ( .A(n35327), .B(n35326), .Z(n35423) );
  XOR U35748 ( .A(n35424), .B(n35423), .Z(n35426) );
  XOR U35749 ( .A(n35425), .B(n35426), .Z(n35413) );
  NANDN U35750 ( .A(n35329), .B(n35328), .Z(n35333) );
  OR U35751 ( .A(n35331), .B(n35330), .Z(n35332) );
  AND U35752 ( .A(n35333), .B(n35332), .Z(n35412) );
  NANDN U35753 ( .A(n35335), .B(n35334), .Z(n35339) );
  NANDN U35754 ( .A(n35337), .B(n35336), .Z(n35338) );
  AND U35755 ( .A(n35339), .B(n35338), .Z(n35432) );
  NANDN U35756 ( .A(n38090), .B(n35344), .Z(n35346) );
  XOR U35757 ( .A(b[59]), .B(a[100]), .Z(n35453) );
  NANDN U35758 ( .A(n38130), .B(n35453), .Z(n35345) );
  AND U35759 ( .A(n35346), .B(n35345), .Z(n35523) );
  NANDN U35760 ( .A(n36210), .B(n35347), .Z(n35349) );
  XOR U35761 ( .A(a[120]), .B(b[39]), .Z(n35450) );
  NANDN U35762 ( .A(n36347), .B(n35450), .Z(n35348) );
  AND U35763 ( .A(n35349), .B(n35348), .Z(n35521) );
  NANDN U35764 ( .A(n37857), .B(n35350), .Z(n35352) );
  XOR U35765 ( .A(b[55]), .B(a[104]), .Z(n35475) );
  NANDN U35766 ( .A(n37911), .B(n35475), .Z(n35351) );
  NAND U35767 ( .A(n35352), .B(n35351), .Z(n35520) );
  XNOR U35768 ( .A(n35521), .B(n35520), .Z(n35522) );
  XNOR U35769 ( .A(n35523), .B(n35522), .Z(n35429) );
  XNOR U35770 ( .A(n35430), .B(n35429), .Z(n35431) );
  XNOR U35771 ( .A(n35432), .B(n35431), .Z(n35411) );
  XOR U35772 ( .A(n35412), .B(n35411), .Z(n35414) );
  XOR U35773 ( .A(n35413), .B(n35414), .Z(n35526) );
  NANDN U35774 ( .A(n35354), .B(n35353), .Z(n35358) );
  NANDN U35775 ( .A(n35356), .B(n35355), .Z(n35357) );
  AND U35776 ( .A(n35358), .B(n35357), .Z(n35401) );
  NANDN U35777 ( .A(n35360), .B(n35359), .Z(n35364) );
  NANDN U35778 ( .A(n35362), .B(n35361), .Z(n35363) );
  AND U35779 ( .A(n35364), .B(n35363), .Z(n35400) );
  NANDN U35780 ( .A(n35366), .B(n35365), .Z(n35370) );
  NANDN U35781 ( .A(n35368), .B(n35367), .Z(n35369) );
  NAND U35782 ( .A(n35370), .B(n35369), .Z(n35399) );
  XOR U35783 ( .A(n35400), .B(n35399), .Z(n35402) );
  XNOR U35784 ( .A(n35401), .B(n35402), .Z(n35527) );
  XOR U35785 ( .A(n35526), .B(n35527), .Z(n35528) );
  XOR U35786 ( .A(n35529), .B(n35528), .Z(n35395) );
  NANDN U35787 ( .A(n35372), .B(n35371), .Z(n35376) );
  OR U35788 ( .A(n35374), .B(n35373), .Z(n35375) );
  AND U35789 ( .A(n35376), .B(n35375), .Z(n35396) );
  XOR U35790 ( .A(n35395), .B(n35396), .Z(n35397) );
  XOR U35791 ( .A(n35398), .B(n35397), .Z(n35391) );
  NANDN U35792 ( .A(n35378), .B(n35377), .Z(n35382) );
  NANDN U35793 ( .A(n35380), .B(n35379), .Z(n35381) );
  AND U35794 ( .A(n35382), .B(n35381), .Z(n35392) );
  XOR U35795 ( .A(n35391), .B(n35392), .Z(n35393) );
  XOR U35796 ( .A(n35394), .B(n35393), .Z(n35385) );
  XOR U35797 ( .A(n35386), .B(n35385), .Z(n35388) );
  XNOR U35798 ( .A(n35387), .B(n35388), .Z(n35383) );
  XOR U35799 ( .A(n35384), .B(n35383), .Z(c[222]) );
  AND U35800 ( .A(n35384), .B(n35383), .Z(n35537) );
  NANDN U35801 ( .A(n35386), .B(n35385), .Z(n35390) );
  OR U35802 ( .A(n35388), .B(n35387), .Z(n35389) );
  AND U35803 ( .A(n35390), .B(n35389), .Z(n35540) );
  NANDN U35804 ( .A(n35400), .B(n35399), .Z(n35404) );
  NANDN U35805 ( .A(n35402), .B(n35401), .Z(n35403) );
  AND U35806 ( .A(n35404), .B(n35403), .Z(n35687) );
  NANDN U35807 ( .A(n35406), .B(n35405), .Z(n35410) );
  NANDN U35808 ( .A(n35408), .B(n35407), .Z(n35409) );
  AND U35809 ( .A(n35410), .B(n35409), .Z(n35686) );
  NANDN U35810 ( .A(n35412), .B(n35411), .Z(n35416) );
  NANDN U35811 ( .A(n35414), .B(n35413), .Z(n35415) );
  AND U35812 ( .A(n35416), .B(n35415), .Z(n35685) );
  XOR U35813 ( .A(n35686), .B(n35685), .Z(n35688) );
  XOR U35814 ( .A(n35687), .B(n35688), .Z(n35546) );
  NANDN U35815 ( .A(n35418), .B(n35417), .Z(n35422) );
  NANDN U35816 ( .A(n35420), .B(n35419), .Z(n35421) );
  NAND U35817 ( .A(n35422), .B(n35421), .Z(n35675) );
  NANDN U35818 ( .A(n35424), .B(n35423), .Z(n35428) );
  NANDN U35819 ( .A(n35426), .B(n35425), .Z(n35427) );
  NAND U35820 ( .A(n35428), .B(n35427), .Z(n35673) );
  NANDN U35821 ( .A(n35430), .B(n35429), .Z(n35434) );
  NANDN U35822 ( .A(n35432), .B(n35431), .Z(n35433) );
  AND U35823 ( .A(n35434), .B(n35433), .Z(n35674) );
  XOR U35824 ( .A(n35673), .B(n35674), .Z(n35676) );
  XNOR U35825 ( .A(n35675), .B(n35676), .Z(n35680) );
  NANDN U35826 ( .A(n35436), .B(n35435), .Z(n35440) );
  NANDN U35827 ( .A(n35438), .B(n35437), .Z(n35439) );
  AND U35828 ( .A(n35440), .B(n35439), .Z(n35679) );
  XOR U35829 ( .A(n35680), .B(n35679), .Z(n35681) );
  NANDN U35830 ( .A(n35442), .B(n35441), .Z(n35446) );
  OR U35831 ( .A(n35444), .B(n35443), .Z(n35445) );
  AND U35832 ( .A(n35446), .B(n35445), .Z(n35551) );
  NANDN U35833 ( .A(n36480), .B(n35447), .Z(n35449) );
  XOR U35834 ( .A(a[119]), .B(b[41]), .Z(n35664) );
  NANDN U35835 ( .A(n36594), .B(n35664), .Z(n35448) );
  AND U35836 ( .A(n35449), .B(n35448), .Z(n35577) );
  NANDN U35837 ( .A(n36210), .B(n35450), .Z(n35452) );
  XOR U35838 ( .A(a[121]), .B(b[39]), .Z(n35670) );
  NANDN U35839 ( .A(n36347), .B(n35670), .Z(n35451) );
  AND U35840 ( .A(n35452), .B(n35451), .Z(n35575) );
  NANDN U35841 ( .A(n38090), .B(n35453), .Z(n35455) );
  XOR U35842 ( .A(b[59]), .B(a[101]), .Z(n35604) );
  NANDN U35843 ( .A(n38130), .B(n35604), .Z(n35454) );
  NAND U35844 ( .A(n35455), .B(n35454), .Z(n35574) );
  XNOR U35845 ( .A(n35575), .B(n35574), .Z(n35576) );
  XNOR U35846 ( .A(n35577), .B(n35576), .Z(n35621) );
  XNOR U35847 ( .A(a[127]), .B(b[33]), .Z(n35653) );
  OR U35848 ( .A(n35653), .B(n35456), .Z(n35459) );
  NAND U35849 ( .A(n35654), .B(n35457), .Z(n35458) );
  AND U35850 ( .A(n35459), .B(n35458), .Z(n35645) );
  NANDN U35851 ( .A(n212), .B(n35460), .Z(n35462) );
  XOR U35852 ( .A(b[49]), .B(a[111]), .Z(n35607) );
  NANDN U35853 ( .A(n37432), .B(n35607), .Z(n35461) );
  NAND U35854 ( .A(n35462), .B(n35461), .Z(n35644) );
  XNOR U35855 ( .A(n35645), .B(n35644), .Z(n35647) );
  AND U35856 ( .A(b[63]), .B(a[95]), .Z(n35580) );
  XOR U35857 ( .A(n35581), .B(n35580), .Z(n35582) );
  XOR U35858 ( .A(n35508), .B(n35582), .Z(n35646) );
  XOR U35859 ( .A(n35647), .B(n35646), .Z(n35620) );
  XOR U35860 ( .A(n35621), .B(n35620), .Z(n35623) );
  NANDN U35861 ( .A(n35464), .B(n35463), .Z(n35468) );
  OR U35862 ( .A(n35466), .B(n35465), .Z(n35467) );
  NAND U35863 ( .A(n35468), .B(n35467), .Z(n35622) );
  XOR U35864 ( .A(n35623), .B(n35622), .Z(n35640) );
  NANDN U35865 ( .A(n211), .B(n35469), .Z(n35471) );
  XOR U35866 ( .A(b[47]), .B(a[113]), .Z(n35667) );
  NANDN U35867 ( .A(n37172), .B(n35667), .Z(n35470) );
  AND U35868 ( .A(n35471), .B(n35470), .Z(n35558) );
  NANDN U35869 ( .A(n36991), .B(n35472), .Z(n35474) );
  XOR U35870 ( .A(a[115]), .B(b[45]), .Z(n35658) );
  NANDN U35871 ( .A(n37083), .B(n35658), .Z(n35473) );
  AND U35872 ( .A(n35474), .B(n35473), .Z(n35557) );
  NANDN U35873 ( .A(n37857), .B(n35475), .Z(n35477) );
  XOR U35874 ( .A(b[55]), .B(a[105]), .Z(n35592) );
  NANDN U35875 ( .A(n37911), .B(n35592), .Z(n35476) );
  AND U35876 ( .A(n35477), .B(n35476), .Z(n35598) );
  NANDN U35877 ( .A(n37974), .B(n35478), .Z(n35480) );
  XOR U35878 ( .A(b[57]), .B(a[103]), .Z(n35601) );
  NANDN U35879 ( .A(n38031), .B(n35601), .Z(n35479) );
  AND U35880 ( .A(n35480), .B(n35479), .Z(n35596) );
  NANDN U35881 ( .A(n36742), .B(n35481), .Z(n35483) );
  XOR U35882 ( .A(a[117]), .B(b[43]), .Z(n35661) );
  NANDN U35883 ( .A(n36891), .B(n35661), .Z(n35482) );
  NAND U35884 ( .A(n35483), .B(n35482), .Z(n35595) );
  XNOR U35885 ( .A(n35596), .B(n35595), .Z(n35597) );
  XNOR U35886 ( .A(n35598), .B(n35597), .Z(n35556) );
  XOR U35887 ( .A(n35557), .B(n35556), .Z(n35559) );
  XOR U35888 ( .A(n35558), .B(n35559), .Z(n35639) );
  NANDN U35889 ( .A(n35485), .B(n35484), .Z(n35489) );
  OR U35890 ( .A(n35487), .B(n35486), .Z(n35488) );
  AND U35891 ( .A(n35489), .B(n35488), .Z(n35638) );
  XOR U35892 ( .A(n35639), .B(n35638), .Z(n35641) );
  XNOR U35893 ( .A(n35640), .B(n35641), .Z(n35550) );
  XNOR U35894 ( .A(n35551), .B(n35550), .Z(n35552) );
  NANDN U35895 ( .A(n38247), .B(n35490), .Z(n35492) );
  XOR U35896 ( .A(b[61]), .B(a[99]), .Z(n35614) );
  NANDN U35897 ( .A(n38248), .B(n35614), .Z(n35491) );
  AND U35898 ( .A(n35492), .B(n35491), .Z(n35565) );
  NANDN U35899 ( .A(n35936), .B(n35493), .Z(n35495) );
  XOR U35900 ( .A(a[123]), .B(b[37]), .Z(n35589) );
  NANDN U35901 ( .A(n36047), .B(n35589), .Z(n35494) );
  AND U35902 ( .A(n35495), .B(n35494), .Z(n35563) );
  NANDN U35903 ( .A(n37705), .B(n35496), .Z(n35498) );
  XOR U35904 ( .A(b[53]), .B(a[107]), .Z(n35586) );
  NANDN U35905 ( .A(n37778), .B(n35586), .Z(n35497) );
  NAND U35906 ( .A(n35498), .B(n35497), .Z(n35562) );
  XNOR U35907 ( .A(n35563), .B(n35562), .Z(n35564) );
  XOR U35908 ( .A(n35565), .B(n35564), .Z(n35627) );
  NANDN U35909 ( .A(n35611), .B(n35499), .Z(n35501) );
  XOR U35910 ( .A(a[125]), .B(b[35]), .Z(n35610) );
  NANDN U35911 ( .A(n35801), .B(n35610), .Z(n35500) );
  AND U35912 ( .A(n35501), .B(n35500), .Z(n35570) );
  NANDN U35913 ( .A(n38278), .B(n35502), .Z(n35504) );
  XOR U35914 ( .A(b[63]), .B(a[97]), .Z(n35650) );
  NANDN U35915 ( .A(n38279), .B(n35650), .Z(n35503) );
  AND U35916 ( .A(n35504), .B(n35503), .Z(n35569) );
  NANDN U35917 ( .A(n37526), .B(n35505), .Z(n35507) );
  XOR U35918 ( .A(b[51]), .B(a[109]), .Z(n35617) );
  NANDN U35919 ( .A(n37605), .B(n35617), .Z(n35506) );
  NAND U35920 ( .A(n35507), .B(n35506), .Z(n35568) );
  XOR U35921 ( .A(n35569), .B(n35568), .Z(n35571) );
  XNOR U35922 ( .A(n35570), .B(n35571), .Z(n35626) );
  XOR U35923 ( .A(n35627), .B(n35626), .Z(n35629) );
  IV U35924 ( .A(n35508), .Z(n35583) );
  NANDN U35925 ( .A(n35583), .B(n35509), .Z(n35513) );
  NANDN U35926 ( .A(n35511), .B(n35510), .Z(n35512) );
  AND U35927 ( .A(n35513), .B(n35512), .Z(n35628) );
  XOR U35928 ( .A(n35629), .B(n35628), .Z(n35635) );
  NANDN U35929 ( .A(n35515), .B(n35514), .Z(n35519) );
  OR U35930 ( .A(n35517), .B(n35516), .Z(n35518) );
  AND U35931 ( .A(n35519), .B(n35518), .Z(n35633) );
  NANDN U35932 ( .A(n35521), .B(n35520), .Z(n35525) );
  NANDN U35933 ( .A(n35523), .B(n35522), .Z(n35524) );
  NAND U35934 ( .A(n35525), .B(n35524), .Z(n35632) );
  XNOR U35935 ( .A(n35633), .B(n35632), .Z(n35634) );
  XOR U35936 ( .A(n35635), .B(n35634), .Z(n35553) );
  XOR U35937 ( .A(n35552), .B(n35553), .Z(n35682) );
  XNOR U35938 ( .A(n35681), .B(n35682), .Z(n35544) );
  XOR U35939 ( .A(n35544), .B(n35545), .Z(n35547) );
  XOR U35940 ( .A(n35546), .B(n35547), .Z(n35692) );
  NANDN U35941 ( .A(n35531), .B(n35530), .Z(n35535) );
  OR U35942 ( .A(n35533), .B(n35532), .Z(n35534) );
  NAND U35943 ( .A(n35535), .B(n35534), .Z(n35691) );
  XOR U35944 ( .A(n35692), .B(n35691), .Z(n35694) );
  XNOR U35945 ( .A(n35693), .B(n35694), .Z(n35538) );
  XOR U35946 ( .A(n35539), .B(n35538), .Z(n35541) );
  XNOR U35947 ( .A(n35540), .B(n35541), .Z(n35536) );
  XOR U35948 ( .A(n35537), .B(n35536), .Z(c[223]) );
  AND U35949 ( .A(n35537), .B(n35536), .Z(n35698) );
  NANDN U35950 ( .A(n35539), .B(n35538), .Z(n35543) );
  OR U35951 ( .A(n35541), .B(n35540), .Z(n35542) );
  AND U35952 ( .A(n35543), .B(n35542), .Z(n35701) );
  NANDN U35953 ( .A(n35545), .B(n35544), .Z(n35549) );
  OR U35954 ( .A(n35547), .B(n35546), .Z(n35548) );
  AND U35955 ( .A(n35549), .B(n35548), .Z(n35843) );
  NANDN U35956 ( .A(n35551), .B(n35550), .Z(n35555) );
  NANDN U35957 ( .A(n35553), .B(n35552), .Z(n35554) );
  AND U35958 ( .A(n35555), .B(n35554), .Z(n35706) );
  NANDN U35959 ( .A(n35557), .B(n35556), .Z(n35561) );
  OR U35960 ( .A(n35559), .B(n35558), .Z(n35560) );
  AND U35961 ( .A(n35561), .B(n35560), .Z(n35725) );
  NANDN U35962 ( .A(n35563), .B(n35562), .Z(n35567) );
  NANDN U35963 ( .A(n35565), .B(n35564), .Z(n35566) );
  AND U35964 ( .A(n35567), .B(n35566), .Z(n35724) );
  NANDN U35965 ( .A(n35569), .B(n35568), .Z(n35573) );
  OR U35966 ( .A(n35571), .B(n35570), .Z(n35572) );
  NAND U35967 ( .A(n35573), .B(n35572), .Z(n35723) );
  XOR U35968 ( .A(n35724), .B(n35723), .Z(n35726) );
  XOR U35969 ( .A(n35725), .B(n35726), .Z(n35755) );
  NANDN U35970 ( .A(n35575), .B(n35574), .Z(n35579) );
  NANDN U35971 ( .A(n35577), .B(n35576), .Z(n35578) );
  AND U35972 ( .A(n35579), .B(n35578), .Z(n35825) );
  NANDN U35973 ( .A(n35581), .B(n35580), .Z(n35585) );
  ANDN U35974 ( .B(n35583), .A(n35582), .Z(n35584) );
  ANDN U35975 ( .B(n35585), .A(n35584), .Z(n35824) );
  NANDN U35976 ( .A(n37705), .B(n35586), .Z(n35588) );
  XOR U35977 ( .A(b[53]), .B(a[108]), .Z(n35789) );
  NANDN U35978 ( .A(n37778), .B(n35789), .Z(n35587) );
  AND U35979 ( .A(n35588), .B(n35587), .Z(n35768) );
  NANDN U35980 ( .A(n35936), .B(n35589), .Z(n35591) );
  XOR U35981 ( .A(a[124]), .B(b[37]), .Z(n35808) );
  NANDN U35982 ( .A(n36047), .B(n35808), .Z(n35590) );
  AND U35983 ( .A(n35591), .B(n35590), .Z(n35766) );
  NANDN U35984 ( .A(n37857), .B(n35592), .Z(n35594) );
  XOR U35985 ( .A(b[55]), .B(a[106]), .Z(n35777) );
  NANDN U35986 ( .A(n37911), .B(n35777), .Z(n35593) );
  NAND U35987 ( .A(n35594), .B(n35593), .Z(n35765) );
  XNOR U35988 ( .A(n35766), .B(n35765), .Z(n35767) );
  XNOR U35989 ( .A(n35768), .B(n35767), .Z(n35823) );
  XOR U35990 ( .A(n35824), .B(n35823), .Z(n35826) );
  XOR U35991 ( .A(n35825), .B(n35826), .Z(n35754) );
  NANDN U35992 ( .A(n35596), .B(n35595), .Z(n35600) );
  NANDN U35993 ( .A(n35598), .B(n35597), .Z(n35599) );
  AND U35994 ( .A(n35600), .B(n35599), .Z(n35831) );
  NANDN U35995 ( .A(n37974), .B(n35601), .Z(n35603) );
  XOR U35996 ( .A(b[57]), .B(a[104]), .Z(n35780) );
  NANDN U35997 ( .A(n38031), .B(n35780), .Z(n35602) );
  AND U35998 ( .A(n35603), .B(n35602), .Z(n35773) );
  NANDN U35999 ( .A(n38090), .B(n35604), .Z(n35606) );
  XOR U36000 ( .A(b[59]), .B(a[102]), .Z(n35811) );
  NANDN U36001 ( .A(n38130), .B(n35811), .Z(n35605) );
  AND U36002 ( .A(n35606), .B(n35605), .Z(n35772) );
  NANDN U36003 ( .A(n212), .B(n35607), .Z(n35609) );
  XOR U36004 ( .A(b[49]), .B(a[112]), .Z(n35805) );
  NANDN U36005 ( .A(n37432), .B(n35805), .Z(n35608) );
  NAND U36006 ( .A(n35609), .B(n35608), .Z(n35771) );
  XOR U36007 ( .A(n35772), .B(n35771), .Z(n35774) );
  XOR U36008 ( .A(n35773), .B(n35774), .Z(n35830) );
  NANDN U36009 ( .A(n35611), .B(n35610), .Z(n35613) );
  XOR U36010 ( .A(a[126]), .B(b[35]), .Z(n35802) );
  NANDN U36011 ( .A(n35801), .B(n35802), .Z(n35612) );
  AND U36012 ( .A(n35613), .B(n35612), .Z(n35749) );
  NANDN U36013 ( .A(n38247), .B(n35614), .Z(n35616) );
  XOR U36014 ( .A(b[61]), .B(a[100]), .Z(n35798) );
  NANDN U36015 ( .A(n38248), .B(n35798), .Z(n35615) );
  AND U36016 ( .A(n35616), .B(n35615), .Z(n35748) );
  NANDN U36017 ( .A(n37526), .B(n35617), .Z(n35619) );
  XOR U36018 ( .A(b[51]), .B(a[110]), .Z(n35744) );
  NANDN U36019 ( .A(n37605), .B(n35744), .Z(n35618) );
  NAND U36020 ( .A(n35619), .B(n35618), .Z(n35747) );
  XOR U36021 ( .A(n35748), .B(n35747), .Z(n35750) );
  XNOR U36022 ( .A(n35749), .B(n35750), .Z(n35829) );
  XOR U36023 ( .A(n35830), .B(n35829), .Z(n35832) );
  XNOR U36024 ( .A(n35831), .B(n35832), .Z(n35753) );
  XOR U36025 ( .A(n35754), .B(n35753), .Z(n35756) );
  XOR U36026 ( .A(n35755), .B(n35756), .Z(n35720) );
  NAND U36027 ( .A(n35621), .B(n35620), .Z(n35625) );
  NAND U36028 ( .A(n35623), .B(n35622), .Z(n35624) );
  AND U36029 ( .A(n35625), .B(n35624), .Z(n35718) );
  NAND U36030 ( .A(n35627), .B(n35626), .Z(n35631) );
  NAND U36031 ( .A(n35629), .B(n35628), .Z(n35630) );
  AND U36032 ( .A(n35631), .B(n35630), .Z(n35717) );
  XNOR U36033 ( .A(n35718), .B(n35717), .Z(n35719) );
  XNOR U36034 ( .A(n35720), .B(n35719), .Z(n35705) );
  XNOR U36035 ( .A(n35706), .B(n35705), .Z(n35708) );
  NANDN U36036 ( .A(n35633), .B(n35632), .Z(n35637) );
  NANDN U36037 ( .A(n35635), .B(n35634), .Z(n35636) );
  AND U36038 ( .A(n35637), .B(n35636), .Z(n35714) );
  NANDN U36039 ( .A(n35639), .B(n35638), .Z(n35643) );
  OR U36040 ( .A(n35641), .B(n35640), .Z(n35642) );
  AND U36041 ( .A(n35643), .B(n35642), .Z(n35711) );
  NANDN U36042 ( .A(n35645), .B(n35644), .Z(n35649) );
  NAND U36043 ( .A(n35647), .B(n35646), .Z(n35648) );
  AND U36044 ( .A(n35649), .B(n35648), .Z(n35730) );
  NANDN U36045 ( .A(n38278), .B(n35650), .Z(n35652) );
  XOR U36046 ( .A(b[63]), .B(a[98]), .Z(n35741) );
  NANDN U36047 ( .A(n38279), .B(n35741), .Z(n35651) );
  AND U36048 ( .A(n35652), .B(n35651), .Z(n35820) );
  NAND U36049 ( .A(b[63]), .B(a[96]), .Z(n35817) );
  ANDN U36050 ( .B(n35654), .A(n35653), .Z(n35657) );
  NAND U36051 ( .A(b[33]), .B(n35655), .Z(n35656) );
  NANDN U36052 ( .A(n35657), .B(n35656), .Z(n35818) );
  XOR U36053 ( .A(n35817), .B(n35818), .Z(n35819) );
  XNOR U36054 ( .A(n35820), .B(n35819), .Z(n35729) );
  XNOR U36055 ( .A(n35730), .B(n35729), .Z(n35731) );
  NANDN U36056 ( .A(n36991), .B(n35658), .Z(n35660) );
  XOR U36057 ( .A(a[116]), .B(b[45]), .Z(n35783) );
  NANDN U36058 ( .A(n37083), .B(n35783), .Z(n35659) );
  AND U36059 ( .A(n35660), .B(n35659), .Z(n35762) );
  NANDN U36060 ( .A(n36742), .B(n35661), .Z(n35663) );
  XOR U36061 ( .A(a[118]), .B(b[43]), .Z(n35786) );
  NANDN U36062 ( .A(n36891), .B(n35786), .Z(n35662) );
  AND U36063 ( .A(n35663), .B(n35662), .Z(n35760) );
  NANDN U36064 ( .A(n36480), .B(n35664), .Z(n35666) );
  XOR U36065 ( .A(a[120]), .B(b[41]), .Z(n35795) );
  NANDN U36066 ( .A(n36594), .B(n35795), .Z(n35665) );
  AND U36067 ( .A(n35666), .B(n35665), .Z(n35738) );
  NANDN U36068 ( .A(n211), .B(n35667), .Z(n35669) );
  XOR U36069 ( .A(a[114]), .B(b[47]), .Z(n35814) );
  NANDN U36070 ( .A(n37172), .B(n35814), .Z(n35668) );
  AND U36071 ( .A(n35669), .B(n35668), .Z(n35736) );
  NANDN U36072 ( .A(n36210), .B(n35670), .Z(n35672) );
  XOR U36073 ( .A(a[122]), .B(b[39]), .Z(n35792) );
  NANDN U36074 ( .A(n36347), .B(n35792), .Z(n35671) );
  NAND U36075 ( .A(n35672), .B(n35671), .Z(n35735) );
  XNOR U36076 ( .A(n35736), .B(n35735), .Z(n35737) );
  XNOR U36077 ( .A(n35738), .B(n35737), .Z(n35759) );
  XNOR U36078 ( .A(n35760), .B(n35759), .Z(n35761) );
  XOR U36079 ( .A(n35762), .B(n35761), .Z(n35732) );
  XOR U36080 ( .A(n35731), .B(n35732), .Z(n35712) );
  XNOR U36081 ( .A(n35711), .B(n35712), .Z(n35713) );
  XNOR U36082 ( .A(n35714), .B(n35713), .Z(n35707) );
  XOR U36083 ( .A(n35708), .B(n35707), .Z(n35837) );
  NAND U36084 ( .A(n35674), .B(n35673), .Z(n35678) );
  NAND U36085 ( .A(n35676), .B(n35675), .Z(n35677) );
  AND U36086 ( .A(n35678), .B(n35677), .Z(n35836) );
  NAND U36087 ( .A(n35680), .B(n35679), .Z(n35684) );
  NANDN U36088 ( .A(n35682), .B(n35681), .Z(n35683) );
  AND U36089 ( .A(n35684), .B(n35683), .Z(n35835) );
  XOR U36090 ( .A(n35836), .B(n35835), .Z(n35838) );
  XOR U36091 ( .A(n35837), .B(n35838), .Z(n35842) );
  NANDN U36092 ( .A(n35686), .B(n35685), .Z(n35690) );
  OR U36093 ( .A(n35688), .B(n35687), .Z(n35689) );
  AND U36094 ( .A(n35690), .B(n35689), .Z(n35841) );
  XOR U36095 ( .A(n35842), .B(n35841), .Z(n35844) );
  XOR U36096 ( .A(n35843), .B(n35844), .Z(n35700) );
  NANDN U36097 ( .A(n35692), .B(n35691), .Z(n35696) );
  NANDN U36098 ( .A(n35694), .B(n35693), .Z(n35695) );
  NAND U36099 ( .A(n35696), .B(n35695), .Z(n35699) );
  XOR U36100 ( .A(n35700), .B(n35699), .Z(n35702) );
  XNOR U36101 ( .A(n35701), .B(n35702), .Z(n35697) );
  XOR U36102 ( .A(n35698), .B(n35697), .Z(c[224]) );
  AND U36103 ( .A(n35698), .B(n35697), .Z(n35848) );
  NANDN U36104 ( .A(n35700), .B(n35699), .Z(n35704) );
  OR U36105 ( .A(n35702), .B(n35701), .Z(n35703) );
  AND U36106 ( .A(n35704), .B(n35703), .Z(n35851) );
  NANDN U36107 ( .A(n35706), .B(n35705), .Z(n35710) );
  NAND U36108 ( .A(n35708), .B(n35707), .Z(n35709) );
  AND U36109 ( .A(n35710), .B(n35709), .Z(n35856) );
  NANDN U36110 ( .A(n35712), .B(n35711), .Z(n35716) );
  NANDN U36111 ( .A(n35714), .B(n35713), .Z(n35715) );
  AND U36112 ( .A(n35716), .B(n35715), .Z(n35862) );
  NANDN U36113 ( .A(n35718), .B(n35717), .Z(n35722) );
  NANDN U36114 ( .A(n35720), .B(n35719), .Z(n35721) );
  NAND U36115 ( .A(n35722), .B(n35721), .Z(n35861) );
  XNOR U36116 ( .A(n35862), .B(n35861), .Z(n35863) );
  NANDN U36117 ( .A(n35724), .B(n35723), .Z(n35728) );
  OR U36118 ( .A(n35726), .B(n35725), .Z(n35727) );
  AND U36119 ( .A(n35728), .B(n35727), .Z(n35990) );
  NANDN U36120 ( .A(n35730), .B(n35729), .Z(n35734) );
  NANDN U36121 ( .A(n35732), .B(n35731), .Z(n35733) );
  AND U36122 ( .A(n35734), .B(n35733), .Z(n35988) );
  NANDN U36123 ( .A(n35736), .B(n35735), .Z(n35740) );
  NANDN U36124 ( .A(n35738), .B(n35737), .Z(n35739) );
  AND U36125 ( .A(n35740), .B(n35739), .Z(n35909) );
  NANDN U36126 ( .A(n38278), .B(n35741), .Z(n35743) );
  XOR U36127 ( .A(b[63]), .B(a[99]), .Z(n35924) );
  NANDN U36128 ( .A(n38279), .B(n35924), .Z(n35742) );
  AND U36129 ( .A(n35743), .B(n35742), .Z(n35874) );
  NANDN U36130 ( .A(n37526), .B(n35744), .Z(n35746) );
  XOR U36131 ( .A(b[51]), .B(a[111]), .Z(n35939) );
  NANDN U36132 ( .A(n37605), .B(n35939), .Z(n35745) );
  NAND U36133 ( .A(n35746), .B(n35745), .Z(n35873) );
  XNOR U36134 ( .A(n35874), .B(n35873), .Z(n35876) );
  AND U36135 ( .A(b[63]), .B(a[97]), .Z(n35960) );
  XOR U36136 ( .A(n35961), .B(n35960), .Z(n35962) );
  XOR U36137 ( .A(n35817), .B(n35962), .Z(n35875) );
  XOR U36138 ( .A(n35876), .B(n35875), .Z(n35907) );
  NANDN U36139 ( .A(n35748), .B(n35747), .Z(n35752) );
  OR U36140 ( .A(n35750), .B(n35749), .Z(n35751) );
  AND U36141 ( .A(n35752), .B(n35751), .Z(n35906) );
  XNOR U36142 ( .A(n35907), .B(n35906), .Z(n35908) );
  XNOR U36143 ( .A(n35909), .B(n35908), .Z(n35987) );
  XNOR U36144 ( .A(n35988), .B(n35987), .Z(n35989) );
  XNOR U36145 ( .A(n35990), .B(n35989), .Z(n35995) );
  NANDN U36146 ( .A(n35754), .B(n35753), .Z(n35758) );
  OR U36147 ( .A(n35756), .B(n35755), .Z(n35757) );
  AND U36148 ( .A(n35758), .B(n35757), .Z(n35993) );
  NANDN U36149 ( .A(n35760), .B(n35759), .Z(n35764) );
  NANDN U36150 ( .A(n35762), .B(n35761), .Z(n35763) );
  AND U36151 ( .A(n35764), .B(n35763), .Z(n35869) );
  NANDN U36152 ( .A(n35766), .B(n35765), .Z(n35770) );
  NANDN U36153 ( .A(n35768), .B(n35767), .Z(n35769) );
  AND U36154 ( .A(n35770), .B(n35769), .Z(n35868) );
  NANDN U36155 ( .A(n35772), .B(n35771), .Z(n35776) );
  OR U36156 ( .A(n35774), .B(n35773), .Z(n35775) );
  NAND U36157 ( .A(n35776), .B(n35775), .Z(n35867) );
  XOR U36158 ( .A(n35868), .B(n35867), .Z(n35870) );
  XOR U36159 ( .A(n35869), .B(n35870), .Z(n35977) );
  NANDN U36160 ( .A(n37857), .B(n35777), .Z(n35779) );
  XOR U36161 ( .A(b[55]), .B(a[107]), .Z(n35972) );
  NANDN U36162 ( .A(n37911), .B(n35972), .Z(n35778) );
  AND U36163 ( .A(n35779), .B(n35778), .Z(n35956) );
  NANDN U36164 ( .A(n37974), .B(n35780), .Z(n35782) );
  XOR U36165 ( .A(b[57]), .B(a[105]), .Z(n35882) );
  NANDN U36166 ( .A(n38031), .B(n35882), .Z(n35781) );
  AND U36167 ( .A(n35782), .B(n35781), .Z(n35955) );
  NANDN U36168 ( .A(n36991), .B(n35783), .Z(n35785) );
  XOR U36169 ( .A(a[117]), .B(b[45]), .Z(n35888) );
  NANDN U36170 ( .A(n37083), .B(n35888), .Z(n35784) );
  NAND U36171 ( .A(n35785), .B(n35784), .Z(n35954) );
  XOR U36172 ( .A(n35955), .B(n35954), .Z(n35957) );
  XOR U36173 ( .A(n35956), .B(n35957), .Z(n35915) );
  NANDN U36174 ( .A(n36742), .B(n35786), .Z(n35788) );
  XNOR U36175 ( .A(a[119]), .B(b[43]), .Z(n35897) );
  NANDN U36176 ( .A(n35897), .B(n36963), .Z(n35787) );
  AND U36177 ( .A(n35788), .B(n35787), .Z(n35944) );
  NANDN U36178 ( .A(n37705), .B(n35789), .Z(n35791) );
  XOR U36179 ( .A(b[53]), .B(a[109]), .Z(n35879) );
  NANDN U36180 ( .A(n37778), .B(n35879), .Z(n35790) );
  AND U36181 ( .A(n35791), .B(n35790), .Z(n35943) );
  NANDN U36182 ( .A(n36210), .B(n35792), .Z(n35794) );
  XOR U36183 ( .A(a[123]), .B(b[39]), .Z(n35932) );
  NANDN U36184 ( .A(n36347), .B(n35932), .Z(n35793) );
  NAND U36185 ( .A(n35794), .B(n35793), .Z(n35942) );
  XOR U36186 ( .A(n35943), .B(n35942), .Z(n35945) );
  XOR U36187 ( .A(n35944), .B(n35945), .Z(n35913) );
  NAND U36188 ( .A(n36735), .B(n35795), .Z(n35797) );
  XNOR U36189 ( .A(a[121]), .B(b[41]), .Z(n35894) );
  NANDN U36190 ( .A(n35894), .B(n36733), .Z(n35796) );
  AND U36191 ( .A(n35797), .B(n35796), .Z(n35912) );
  XNOR U36192 ( .A(n35913), .B(n35912), .Z(n35914) );
  XNOR U36193 ( .A(n35915), .B(n35914), .Z(n35975) );
  NAND U36194 ( .A(n37921), .B(n35798), .Z(n35800) );
  XNOR U36195 ( .A(b[61]), .B(a[101]), .Z(n35969) );
  NANDN U36196 ( .A(n35969), .B(n37864), .Z(n35799) );
  NAND U36197 ( .A(n35800), .B(n35799), .Z(n35949) );
  XNOR U36198 ( .A(a[127]), .B(b[35]), .Z(n35927) );
  OR U36199 ( .A(n35927), .B(n35801), .Z(n35804) );
  NAND U36200 ( .A(n35928), .B(n35802), .Z(n35803) );
  NAND U36201 ( .A(n35804), .B(n35803), .Z(n35948) );
  XOR U36202 ( .A(n35949), .B(n35948), .Z(n35951) );
  NANDN U36203 ( .A(n212), .B(n35805), .Z(n35807) );
  XOR U36204 ( .A(b[49]), .B(a[113]), .Z(n35891) );
  NANDN U36205 ( .A(n37432), .B(n35891), .Z(n35806) );
  NAND U36206 ( .A(n35807), .B(n35806), .Z(n35950) );
  XOR U36207 ( .A(n35951), .B(n35950), .Z(n35919) );
  NANDN U36208 ( .A(n35936), .B(n35808), .Z(n35810) );
  XOR U36209 ( .A(a[125]), .B(b[37]), .Z(n35935) );
  NANDN U36210 ( .A(n36047), .B(n35935), .Z(n35809) );
  AND U36211 ( .A(n35810), .B(n35809), .Z(n35902) );
  NANDN U36212 ( .A(n38090), .B(n35811), .Z(n35813) );
  XOR U36213 ( .A(b[59]), .B(a[103]), .Z(n35966) );
  NANDN U36214 ( .A(n38130), .B(n35966), .Z(n35812) );
  AND U36215 ( .A(n35813), .B(n35812), .Z(n35901) );
  NANDN U36216 ( .A(n211), .B(n35814), .Z(n35816) );
  XOR U36217 ( .A(a[115]), .B(b[47]), .Z(n35885) );
  NANDN U36218 ( .A(n37172), .B(n35885), .Z(n35815) );
  NAND U36219 ( .A(n35816), .B(n35815), .Z(n35900) );
  XOR U36220 ( .A(n35901), .B(n35900), .Z(n35903) );
  XNOR U36221 ( .A(n35902), .B(n35903), .Z(n35918) );
  XNOR U36222 ( .A(n35919), .B(n35918), .Z(n35920) );
  IV U36223 ( .A(n35817), .Z(n35963) );
  NANDN U36224 ( .A(n35963), .B(n35818), .Z(n35822) );
  NANDN U36225 ( .A(n35820), .B(n35819), .Z(n35821) );
  NAND U36226 ( .A(n35822), .B(n35821), .Z(n35921) );
  XOR U36227 ( .A(n35920), .B(n35921), .Z(n35976) );
  XOR U36228 ( .A(n35975), .B(n35976), .Z(n35978) );
  XOR U36229 ( .A(n35977), .B(n35978), .Z(n35984) );
  NANDN U36230 ( .A(n35824), .B(n35823), .Z(n35828) );
  OR U36231 ( .A(n35826), .B(n35825), .Z(n35827) );
  AND U36232 ( .A(n35828), .B(n35827), .Z(n35982) );
  NANDN U36233 ( .A(n35830), .B(n35829), .Z(n35834) );
  NANDN U36234 ( .A(n35832), .B(n35831), .Z(n35833) );
  AND U36235 ( .A(n35834), .B(n35833), .Z(n35981) );
  XNOR U36236 ( .A(n35982), .B(n35981), .Z(n35983) );
  XOR U36237 ( .A(n35984), .B(n35983), .Z(n35994) );
  XOR U36238 ( .A(n35993), .B(n35994), .Z(n35996) );
  XOR U36239 ( .A(n35995), .B(n35996), .Z(n35864) );
  XNOR U36240 ( .A(n35863), .B(n35864), .Z(n35855) );
  XNOR U36241 ( .A(n35856), .B(n35855), .Z(n35858) );
  NANDN U36242 ( .A(n35836), .B(n35835), .Z(n35840) );
  OR U36243 ( .A(n35838), .B(n35837), .Z(n35839) );
  AND U36244 ( .A(n35840), .B(n35839), .Z(n35857) );
  XOR U36245 ( .A(n35858), .B(n35857), .Z(n35850) );
  NANDN U36246 ( .A(n35842), .B(n35841), .Z(n35846) );
  OR U36247 ( .A(n35844), .B(n35843), .Z(n35845) );
  AND U36248 ( .A(n35846), .B(n35845), .Z(n35849) );
  XOR U36249 ( .A(n35850), .B(n35849), .Z(n35852) );
  XNOR U36250 ( .A(n35851), .B(n35852), .Z(n35847) );
  XOR U36251 ( .A(n35848), .B(n35847), .Z(c[225]) );
  AND U36252 ( .A(n35848), .B(n35847), .Z(n36000) );
  NANDN U36253 ( .A(n35850), .B(n35849), .Z(n35854) );
  OR U36254 ( .A(n35852), .B(n35851), .Z(n35853) );
  AND U36255 ( .A(n35854), .B(n35853), .Z(n36003) );
  NANDN U36256 ( .A(n35856), .B(n35855), .Z(n35860) );
  NAND U36257 ( .A(n35858), .B(n35857), .Z(n35859) );
  AND U36258 ( .A(n35860), .B(n35859), .Z(n36001) );
  NANDN U36259 ( .A(n35862), .B(n35861), .Z(n35866) );
  NANDN U36260 ( .A(n35864), .B(n35863), .Z(n35865) );
  AND U36261 ( .A(n35866), .B(n35865), .Z(n36009) );
  NANDN U36262 ( .A(n35868), .B(n35867), .Z(n35872) );
  OR U36263 ( .A(n35870), .B(n35869), .Z(n35871) );
  AND U36264 ( .A(n35872), .B(n35871), .Z(n36131) );
  NANDN U36265 ( .A(n35874), .B(n35873), .Z(n35878) );
  NAND U36266 ( .A(n35876), .B(n35875), .Z(n35877) );
  AND U36267 ( .A(n35878), .B(n35877), .Z(n36096) );
  NANDN U36268 ( .A(n37705), .B(n35879), .Z(n35881) );
  XOR U36269 ( .A(b[53]), .B(a[110]), .Z(n36069) );
  NANDN U36270 ( .A(n37778), .B(n36069), .Z(n35880) );
  AND U36271 ( .A(n35881), .B(n35880), .Z(n36089) );
  NANDN U36272 ( .A(n37974), .B(n35882), .Z(n35884) );
  XOR U36273 ( .A(b[57]), .B(a[106]), .Z(n36072) );
  NANDN U36274 ( .A(n38031), .B(n36072), .Z(n35883) );
  AND U36275 ( .A(n35884), .B(n35883), .Z(n36088) );
  NANDN U36276 ( .A(n211), .B(n35885), .Z(n35887) );
  XOR U36277 ( .A(a[116]), .B(b[47]), .Z(n36111) );
  NANDN U36278 ( .A(n37172), .B(n36111), .Z(n35886) );
  NAND U36279 ( .A(n35887), .B(n35886), .Z(n36087) );
  XOR U36280 ( .A(n36088), .B(n36087), .Z(n36090) );
  XOR U36281 ( .A(n36089), .B(n36090), .Z(n36102) );
  NANDN U36282 ( .A(n36991), .B(n35888), .Z(n35890) );
  XOR U36283 ( .A(a[118]), .B(b[45]), .Z(n36075) );
  NANDN U36284 ( .A(n37083), .B(n36075), .Z(n35889) );
  AND U36285 ( .A(n35890), .B(n35889), .Z(n36119) );
  NANDN U36286 ( .A(n212), .B(n35891), .Z(n35893) );
  XOR U36287 ( .A(b[49]), .B(a[114]), .Z(n36060) );
  NANDN U36288 ( .A(n37432), .B(n36060), .Z(n35892) );
  AND U36289 ( .A(n35893), .B(n35892), .Z(n36118) );
  NANDN U36290 ( .A(n35894), .B(n36735), .Z(n35896) );
  XOR U36291 ( .A(a[122]), .B(b[41]), .Z(n36063) );
  NANDN U36292 ( .A(n36594), .B(n36063), .Z(n35895) );
  NAND U36293 ( .A(n35896), .B(n35895), .Z(n36117) );
  XOR U36294 ( .A(n36118), .B(n36117), .Z(n36120) );
  XOR U36295 ( .A(n36119), .B(n36120), .Z(n36100) );
  NANDN U36296 ( .A(n35897), .B(n36962), .Z(n35899) );
  XNOR U36297 ( .A(a[120]), .B(b[43]), .Z(n36078) );
  NANDN U36298 ( .A(n36078), .B(n36963), .Z(n35898) );
  AND U36299 ( .A(n35899), .B(n35898), .Z(n36099) );
  XNOR U36300 ( .A(n36100), .B(n36099), .Z(n36101) );
  XNOR U36301 ( .A(n36102), .B(n36101), .Z(n36093) );
  NANDN U36302 ( .A(n35901), .B(n35900), .Z(n35905) );
  OR U36303 ( .A(n35903), .B(n35902), .Z(n35904) );
  NAND U36304 ( .A(n35905), .B(n35904), .Z(n36094) );
  XNOR U36305 ( .A(n36093), .B(n36094), .Z(n36095) );
  XOR U36306 ( .A(n36096), .B(n36095), .Z(n36130) );
  NANDN U36307 ( .A(n35907), .B(n35906), .Z(n35911) );
  NAND U36308 ( .A(n35909), .B(n35908), .Z(n35910) );
  AND U36309 ( .A(n35911), .B(n35910), .Z(n36129) );
  XOR U36310 ( .A(n36130), .B(n36129), .Z(n36132) );
  XOR U36311 ( .A(n36131), .B(n36132), .Z(n36021) );
  NANDN U36312 ( .A(n35913), .B(n35912), .Z(n35917) );
  NANDN U36313 ( .A(n35915), .B(n35914), .Z(n35916) );
  AND U36314 ( .A(n35917), .B(n35916), .Z(n36025) );
  NANDN U36315 ( .A(n35919), .B(n35918), .Z(n35923) );
  NANDN U36316 ( .A(n35921), .B(n35920), .Z(n35922) );
  NAND U36317 ( .A(n35923), .B(n35922), .Z(n36026) );
  XNOR U36318 ( .A(n36025), .B(n36026), .Z(n36028) );
  NANDN U36319 ( .A(n38278), .B(n35924), .Z(n35926) );
  XOR U36320 ( .A(b[63]), .B(a[100]), .Z(n36108) );
  NANDN U36321 ( .A(n38279), .B(n36108), .Z(n35925) );
  AND U36322 ( .A(n35926), .B(n35925), .Z(n36116) );
  NAND U36323 ( .A(b[63]), .B(a[98]), .Z(n36185) );
  ANDN U36324 ( .B(n35928), .A(n35927), .Z(n35931) );
  NAND U36325 ( .A(b[35]), .B(n35929), .Z(n35930) );
  NANDN U36326 ( .A(n35931), .B(n35930), .Z(n36114) );
  XOR U36327 ( .A(n36185), .B(n36114), .Z(n36115) );
  XOR U36328 ( .A(n36116), .B(n36115), .Z(n36031) );
  NANDN U36329 ( .A(n36210), .B(n35932), .Z(n35934) );
  XOR U36330 ( .A(a[124]), .B(b[39]), .Z(n36066) );
  NANDN U36331 ( .A(n36347), .B(n36066), .Z(n35933) );
  AND U36332 ( .A(n35934), .B(n35933), .Z(n36043) );
  NANDN U36333 ( .A(n35936), .B(n35935), .Z(n35938) );
  XOR U36334 ( .A(a[126]), .B(b[37]), .Z(n36048) );
  NANDN U36335 ( .A(n36047), .B(n36048), .Z(n35937) );
  AND U36336 ( .A(n35938), .B(n35937), .Z(n36042) );
  NANDN U36337 ( .A(n37526), .B(n35939), .Z(n35941) );
  XOR U36338 ( .A(b[51]), .B(a[112]), .Z(n36051) );
  NANDN U36339 ( .A(n37605), .B(n36051), .Z(n35940) );
  NAND U36340 ( .A(n35941), .B(n35940), .Z(n36041) );
  XOR U36341 ( .A(n36042), .B(n36041), .Z(n36044) );
  XNOR U36342 ( .A(n36043), .B(n36044), .Z(n36032) );
  XOR U36343 ( .A(n36031), .B(n36032), .Z(n36033) );
  NANDN U36344 ( .A(n35943), .B(n35942), .Z(n35947) );
  OR U36345 ( .A(n35945), .B(n35944), .Z(n35946) );
  NAND U36346 ( .A(n35947), .B(n35946), .Z(n36034) );
  XOR U36347 ( .A(n36033), .B(n36034), .Z(n36124) );
  NAND U36348 ( .A(n35949), .B(n35948), .Z(n35953) );
  NAND U36349 ( .A(n35951), .B(n35950), .Z(n35952) );
  NAND U36350 ( .A(n35953), .B(n35952), .Z(n36123) );
  XOR U36351 ( .A(n36124), .B(n36123), .Z(n36126) );
  NANDN U36352 ( .A(n35955), .B(n35954), .Z(n35959) );
  OR U36353 ( .A(n35957), .B(n35956), .Z(n35958) );
  AND U36354 ( .A(n35959), .B(n35958), .Z(n36037) );
  NANDN U36355 ( .A(n35961), .B(n35960), .Z(n35965) );
  ANDN U36356 ( .B(n35963), .A(n35962), .Z(n35964) );
  ANDN U36357 ( .B(n35965), .A(n35964), .Z(n36036) );
  NANDN U36358 ( .A(n38090), .B(n35966), .Z(n35968) );
  XOR U36359 ( .A(b[59]), .B(a[104]), .Z(n36057) );
  NANDN U36360 ( .A(n38130), .B(n36057), .Z(n35967) );
  AND U36361 ( .A(n35968), .B(n35967), .Z(n36084) );
  NANDN U36362 ( .A(n35969), .B(n37921), .Z(n35971) );
  XOR U36363 ( .A(b[61]), .B(a[102]), .Z(n36105) );
  NANDN U36364 ( .A(n38248), .B(n36105), .Z(n35970) );
  AND U36365 ( .A(n35971), .B(n35970), .Z(n36082) );
  NANDN U36366 ( .A(n37857), .B(n35972), .Z(n35974) );
  XOR U36367 ( .A(b[55]), .B(a[108]), .Z(n36054) );
  NANDN U36368 ( .A(n37911), .B(n36054), .Z(n35973) );
  NAND U36369 ( .A(n35974), .B(n35973), .Z(n36081) );
  XNOR U36370 ( .A(n36082), .B(n36081), .Z(n36083) );
  XNOR U36371 ( .A(n36084), .B(n36083), .Z(n36035) );
  XOR U36372 ( .A(n36036), .B(n36035), .Z(n36038) );
  XOR U36373 ( .A(n36037), .B(n36038), .Z(n36125) );
  XOR U36374 ( .A(n36126), .B(n36125), .Z(n36027) );
  XOR U36375 ( .A(n36028), .B(n36027), .Z(n36020) );
  NANDN U36376 ( .A(n35976), .B(n35975), .Z(n35980) );
  OR U36377 ( .A(n35978), .B(n35977), .Z(n35979) );
  NAND U36378 ( .A(n35980), .B(n35979), .Z(n36019) );
  XOR U36379 ( .A(n36020), .B(n36019), .Z(n36022) );
  XOR U36380 ( .A(n36021), .B(n36022), .Z(n36015) );
  NANDN U36381 ( .A(n35982), .B(n35981), .Z(n35986) );
  NANDN U36382 ( .A(n35984), .B(n35983), .Z(n35985) );
  AND U36383 ( .A(n35986), .B(n35985), .Z(n36014) );
  NANDN U36384 ( .A(n35988), .B(n35987), .Z(n35992) );
  NANDN U36385 ( .A(n35990), .B(n35989), .Z(n35991) );
  NAND U36386 ( .A(n35992), .B(n35991), .Z(n36013) );
  XOR U36387 ( .A(n36014), .B(n36013), .Z(n36016) );
  XOR U36388 ( .A(n36015), .B(n36016), .Z(n36008) );
  NANDN U36389 ( .A(n35994), .B(n35993), .Z(n35998) );
  NANDN U36390 ( .A(n35996), .B(n35995), .Z(n35997) );
  AND U36391 ( .A(n35998), .B(n35997), .Z(n36007) );
  XOR U36392 ( .A(n36008), .B(n36007), .Z(n36010) );
  XOR U36393 ( .A(n36009), .B(n36010), .Z(n36002) );
  XOR U36394 ( .A(n36001), .B(n36002), .Z(n36004) );
  XNOR U36395 ( .A(n36003), .B(n36004), .Z(n35999) );
  XOR U36396 ( .A(n36000), .B(n35999), .Z(c[226]) );
  AND U36397 ( .A(n36000), .B(n35999), .Z(n36136) );
  NANDN U36398 ( .A(n36002), .B(n36001), .Z(n36006) );
  OR U36399 ( .A(n36004), .B(n36003), .Z(n36005) );
  AND U36400 ( .A(n36006), .B(n36005), .Z(n36139) );
  NANDN U36401 ( .A(n36008), .B(n36007), .Z(n36012) );
  NANDN U36402 ( .A(n36010), .B(n36009), .Z(n36011) );
  AND U36403 ( .A(n36012), .B(n36011), .Z(n36138) );
  NANDN U36404 ( .A(n36014), .B(n36013), .Z(n36018) );
  OR U36405 ( .A(n36016), .B(n36015), .Z(n36017) );
  AND U36406 ( .A(n36018), .B(n36017), .Z(n36145) );
  NANDN U36407 ( .A(n36020), .B(n36019), .Z(n36024) );
  OR U36408 ( .A(n36022), .B(n36021), .Z(n36023) );
  AND U36409 ( .A(n36024), .B(n36023), .Z(n36144) );
  NANDN U36410 ( .A(n36026), .B(n36025), .Z(n36030) );
  NAND U36411 ( .A(n36028), .B(n36027), .Z(n36029) );
  AND U36412 ( .A(n36030), .B(n36029), .Z(n36151) );
  NANDN U36413 ( .A(n36036), .B(n36035), .Z(n36040) );
  OR U36414 ( .A(n36038), .B(n36037), .Z(n36039) );
  AND U36415 ( .A(n36040), .B(n36039), .Z(n36260) );
  XNOR U36416 ( .A(n36261), .B(n36260), .Z(n36263) );
  NANDN U36417 ( .A(n36042), .B(n36041), .Z(n36046) );
  OR U36418 ( .A(n36044), .B(n36043), .Z(n36045) );
  AND U36419 ( .A(n36046), .B(n36045), .Z(n36250) );
  XNOR U36420 ( .A(a[127]), .B(b[37]), .Z(n36237) );
  OR U36421 ( .A(n36237), .B(n36047), .Z(n36050) );
  NAND U36422 ( .A(n36238), .B(n36048), .Z(n36049) );
  AND U36423 ( .A(n36050), .B(n36049), .Z(n36168) );
  NANDN U36424 ( .A(n37526), .B(n36051), .Z(n36053) );
  XOR U36425 ( .A(b[51]), .B(a[113]), .Z(n36216) );
  NANDN U36426 ( .A(n37605), .B(n36216), .Z(n36052) );
  NAND U36427 ( .A(n36053), .B(n36052), .Z(n36167) );
  XNOR U36428 ( .A(n36168), .B(n36167), .Z(n36169) );
  AND U36429 ( .A(b[63]), .B(a[99]), .Z(n36183) );
  XNOR U36430 ( .A(n36183), .B(n36182), .Z(n36184) );
  XNOR U36431 ( .A(n36185), .B(n36184), .Z(n36170) );
  XOR U36432 ( .A(n36169), .B(n36170), .Z(n36248) );
  NANDN U36433 ( .A(n37857), .B(n36054), .Z(n36056) );
  XOR U36434 ( .A(b[55]), .B(a[109]), .Z(n36200) );
  NANDN U36435 ( .A(n37911), .B(n36200), .Z(n36055) );
  AND U36436 ( .A(n36056), .B(n36055), .Z(n36191) );
  NANDN U36437 ( .A(n38090), .B(n36057), .Z(n36059) );
  XOR U36438 ( .A(b[59]), .B(a[105]), .Z(n36225) );
  NANDN U36439 ( .A(n38130), .B(n36225), .Z(n36058) );
  AND U36440 ( .A(n36059), .B(n36058), .Z(n36189) );
  NANDN U36441 ( .A(n212), .B(n36060), .Z(n36062) );
  XOR U36442 ( .A(b[49]), .B(a[115]), .Z(n36176) );
  NANDN U36443 ( .A(n37432), .B(n36176), .Z(n36061) );
  NAND U36444 ( .A(n36062), .B(n36061), .Z(n36188) );
  XNOR U36445 ( .A(n36189), .B(n36188), .Z(n36190) );
  XOR U36446 ( .A(n36191), .B(n36190), .Z(n36249) );
  XOR U36447 ( .A(n36248), .B(n36249), .Z(n36251) );
  XOR U36448 ( .A(n36250), .B(n36251), .Z(n36257) );
  NANDN U36449 ( .A(n36480), .B(n36063), .Z(n36065) );
  XOR U36450 ( .A(a[123]), .B(b[41]), .Z(n36228) );
  NANDN U36451 ( .A(n36594), .B(n36228), .Z(n36064) );
  AND U36452 ( .A(n36065), .B(n36064), .Z(n36163) );
  NANDN U36453 ( .A(n36210), .B(n36066), .Z(n36068) );
  XOR U36454 ( .A(a[125]), .B(b[39]), .Z(n36209) );
  NANDN U36455 ( .A(n36347), .B(n36209), .Z(n36067) );
  AND U36456 ( .A(n36068), .B(n36067), .Z(n36162) );
  NANDN U36457 ( .A(n37705), .B(n36069), .Z(n36071) );
  XOR U36458 ( .A(b[53]), .B(a[111]), .Z(n36231) );
  NANDN U36459 ( .A(n37778), .B(n36231), .Z(n36070) );
  NAND U36460 ( .A(n36071), .B(n36070), .Z(n36161) );
  XOR U36461 ( .A(n36162), .B(n36161), .Z(n36164) );
  XOR U36462 ( .A(n36163), .B(n36164), .Z(n36195) );
  NANDN U36463 ( .A(n37974), .B(n36072), .Z(n36074) );
  XOR U36464 ( .A(b[57]), .B(a[107]), .Z(n36203) );
  NANDN U36465 ( .A(n38031), .B(n36203), .Z(n36073) );
  AND U36466 ( .A(n36074), .B(n36073), .Z(n36244) );
  NANDN U36467 ( .A(n36991), .B(n36075), .Z(n36077) );
  XOR U36468 ( .A(a[119]), .B(b[45]), .Z(n36179) );
  NANDN U36469 ( .A(n37083), .B(n36179), .Z(n36076) );
  AND U36470 ( .A(n36077), .B(n36076), .Z(n36243) );
  NANDN U36471 ( .A(n36078), .B(n36962), .Z(n36080) );
  XOR U36472 ( .A(a[121]), .B(b[43]), .Z(n36206) );
  NANDN U36473 ( .A(n36891), .B(n36206), .Z(n36079) );
  NAND U36474 ( .A(n36080), .B(n36079), .Z(n36242) );
  XOR U36475 ( .A(n36243), .B(n36242), .Z(n36245) );
  XNOR U36476 ( .A(n36244), .B(n36245), .Z(n36194) );
  XNOR U36477 ( .A(n36195), .B(n36194), .Z(n36196) );
  NANDN U36478 ( .A(n36082), .B(n36081), .Z(n36086) );
  NANDN U36479 ( .A(n36084), .B(n36083), .Z(n36085) );
  NAND U36480 ( .A(n36086), .B(n36085), .Z(n36197) );
  XNOR U36481 ( .A(n36196), .B(n36197), .Z(n36254) );
  NANDN U36482 ( .A(n36088), .B(n36087), .Z(n36092) );
  OR U36483 ( .A(n36090), .B(n36089), .Z(n36091) );
  NAND U36484 ( .A(n36092), .B(n36091), .Z(n36255) );
  XNOR U36485 ( .A(n36254), .B(n36255), .Z(n36256) );
  XNOR U36486 ( .A(n36257), .B(n36256), .Z(n36262) );
  XOR U36487 ( .A(n36263), .B(n36262), .Z(n36150) );
  NANDN U36488 ( .A(n36094), .B(n36093), .Z(n36098) );
  NAND U36489 ( .A(n36096), .B(n36095), .Z(n36097) );
  AND U36490 ( .A(n36098), .B(n36097), .Z(n36268) );
  NANDN U36491 ( .A(n36100), .B(n36099), .Z(n36104) );
  NANDN U36492 ( .A(n36102), .B(n36101), .Z(n36103) );
  AND U36493 ( .A(n36104), .B(n36103), .Z(n36267) );
  NANDN U36494 ( .A(n38247), .B(n36105), .Z(n36107) );
  XOR U36495 ( .A(b[61]), .B(a[103]), .Z(n36213) );
  NANDN U36496 ( .A(n38248), .B(n36213), .Z(n36106) );
  AND U36497 ( .A(n36107), .B(n36106), .Z(n36221) );
  NANDN U36498 ( .A(n38278), .B(n36108), .Z(n36110) );
  XOR U36499 ( .A(b[63]), .B(a[101]), .Z(n36234) );
  NANDN U36500 ( .A(n38279), .B(n36234), .Z(n36109) );
  AND U36501 ( .A(n36110), .B(n36109), .Z(n36220) );
  NANDN U36502 ( .A(n211), .B(n36111), .Z(n36113) );
  XOR U36503 ( .A(a[117]), .B(b[47]), .Z(n36173) );
  NANDN U36504 ( .A(n37172), .B(n36173), .Z(n36112) );
  NAND U36505 ( .A(n36113), .B(n36112), .Z(n36219) );
  XOR U36506 ( .A(n36220), .B(n36219), .Z(n36222) );
  XOR U36507 ( .A(n36221), .B(n36222), .Z(n36156) );
  XNOR U36508 ( .A(n36156), .B(n36155), .Z(n36157) );
  NANDN U36509 ( .A(n36118), .B(n36117), .Z(n36122) );
  OR U36510 ( .A(n36120), .B(n36119), .Z(n36121) );
  NAND U36511 ( .A(n36122), .B(n36121), .Z(n36158) );
  XNOR U36512 ( .A(n36157), .B(n36158), .Z(n36266) );
  XOR U36513 ( .A(n36267), .B(n36266), .Z(n36269) );
  XNOR U36514 ( .A(n36268), .B(n36269), .Z(n36149) );
  XOR U36515 ( .A(n36150), .B(n36149), .Z(n36152) );
  XOR U36516 ( .A(n36151), .B(n36152), .Z(n36275) );
  NAND U36517 ( .A(n36124), .B(n36123), .Z(n36128) );
  NAND U36518 ( .A(n36126), .B(n36125), .Z(n36127) );
  AND U36519 ( .A(n36128), .B(n36127), .Z(n36272) );
  NANDN U36520 ( .A(n36130), .B(n36129), .Z(n36134) );
  OR U36521 ( .A(n36132), .B(n36131), .Z(n36133) );
  NAND U36522 ( .A(n36134), .B(n36133), .Z(n36273) );
  XNOR U36523 ( .A(n36272), .B(n36273), .Z(n36274) );
  XNOR U36524 ( .A(n36275), .B(n36274), .Z(n36143) );
  XOR U36525 ( .A(n36144), .B(n36143), .Z(n36146) );
  XNOR U36526 ( .A(n36145), .B(n36146), .Z(n36137) );
  XOR U36527 ( .A(n36138), .B(n36137), .Z(n36140) );
  XNOR U36528 ( .A(n36139), .B(n36140), .Z(n36135) );
  XOR U36529 ( .A(n36136), .B(n36135), .Z(c[227]) );
  AND U36530 ( .A(n36136), .B(n36135), .Z(n36279) );
  NANDN U36531 ( .A(n36138), .B(n36137), .Z(n36142) );
  OR U36532 ( .A(n36140), .B(n36139), .Z(n36141) );
  AND U36533 ( .A(n36142), .B(n36141), .Z(n36282) );
  NANDN U36534 ( .A(n36144), .B(n36143), .Z(n36148) );
  NANDN U36535 ( .A(n36146), .B(n36145), .Z(n36147) );
  AND U36536 ( .A(n36148), .B(n36147), .Z(n36281) );
  NANDN U36537 ( .A(n36150), .B(n36149), .Z(n36154) );
  OR U36538 ( .A(n36152), .B(n36151), .Z(n36153) );
  AND U36539 ( .A(n36154), .B(n36153), .Z(n36406) );
  NANDN U36540 ( .A(n36156), .B(n36155), .Z(n36160) );
  NANDN U36541 ( .A(n36158), .B(n36157), .Z(n36159) );
  AND U36542 ( .A(n36160), .B(n36159), .Z(n36383) );
  NANDN U36543 ( .A(n36162), .B(n36161), .Z(n36166) );
  OR U36544 ( .A(n36164), .B(n36163), .Z(n36165) );
  AND U36545 ( .A(n36166), .B(n36165), .Z(n36388) );
  NANDN U36546 ( .A(n36168), .B(n36167), .Z(n36172) );
  NAND U36547 ( .A(n36170), .B(n36169), .Z(n36171) );
  NAND U36548 ( .A(n36172), .B(n36171), .Z(n36387) );
  XNOR U36549 ( .A(n36388), .B(n36387), .Z(n36390) );
  NANDN U36550 ( .A(n211), .B(n36173), .Z(n36175) );
  XOR U36551 ( .A(a[118]), .B(b[47]), .Z(n36354) );
  NANDN U36552 ( .A(n37172), .B(n36354), .Z(n36174) );
  AND U36553 ( .A(n36175), .B(n36174), .Z(n36307) );
  NANDN U36554 ( .A(n212), .B(n36176), .Z(n36178) );
  XOR U36555 ( .A(a[116]), .B(b[49]), .Z(n36360) );
  NANDN U36556 ( .A(n37432), .B(n36360), .Z(n36177) );
  AND U36557 ( .A(n36178), .B(n36177), .Z(n36305) );
  NANDN U36558 ( .A(n36991), .B(n36179), .Z(n36181) );
  XOR U36559 ( .A(a[120]), .B(b[45]), .Z(n36357) );
  NANDN U36560 ( .A(n37083), .B(n36357), .Z(n36180) );
  NAND U36561 ( .A(n36181), .B(n36180), .Z(n36304) );
  XNOR U36562 ( .A(n36305), .B(n36304), .Z(n36306) );
  XNOR U36563 ( .A(n36307), .B(n36306), .Z(n36376) );
  ANDN U36564 ( .B(n36183), .A(n36182), .Z(n36187) );
  NANDN U36565 ( .A(n36185), .B(n36184), .Z(n36186) );
  NANDN U36566 ( .A(n36187), .B(n36186), .Z(n36375) );
  XOR U36567 ( .A(n36376), .B(n36375), .Z(n36378) );
  NANDN U36568 ( .A(n36189), .B(n36188), .Z(n36193) );
  NANDN U36569 ( .A(n36191), .B(n36190), .Z(n36192) );
  NAND U36570 ( .A(n36193), .B(n36192), .Z(n36377) );
  XOR U36571 ( .A(n36378), .B(n36377), .Z(n36389) );
  XOR U36572 ( .A(n36390), .B(n36389), .Z(n36382) );
  NANDN U36573 ( .A(n36195), .B(n36194), .Z(n36199) );
  NANDN U36574 ( .A(n36197), .B(n36196), .Z(n36198) );
  NAND U36575 ( .A(n36199), .B(n36198), .Z(n36381) );
  XOR U36576 ( .A(n36382), .B(n36381), .Z(n36384) );
  XOR U36577 ( .A(n36383), .B(n36384), .Z(n36294) );
  NANDN U36578 ( .A(n37857), .B(n36200), .Z(n36202) );
  XOR U36579 ( .A(b[55]), .B(a[110]), .Z(n36329) );
  NANDN U36580 ( .A(n37911), .B(n36329), .Z(n36201) );
  AND U36581 ( .A(n36202), .B(n36201), .Z(n36371) );
  NANDN U36582 ( .A(n37974), .B(n36203), .Z(n36205) );
  XOR U36583 ( .A(b[57]), .B(a[108]), .Z(n36363) );
  NANDN U36584 ( .A(n38031), .B(n36363), .Z(n36204) );
  AND U36585 ( .A(n36205), .B(n36204), .Z(n36370) );
  NANDN U36586 ( .A(n36742), .B(n36206), .Z(n36208) );
  XOR U36587 ( .A(a[122]), .B(b[43]), .Z(n36366) );
  NANDN U36588 ( .A(n36891), .B(n36366), .Z(n36207) );
  NAND U36589 ( .A(n36208), .B(n36207), .Z(n36369) );
  XOR U36590 ( .A(n36370), .B(n36369), .Z(n36372) );
  XOR U36591 ( .A(n36371), .B(n36372), .Z(n36400) );
  NANDN U36592 ( .A(n36210), .B(n36209), .Z(n36212) );
  XOR U36593 ( .A(a[126]), .B(b[39]), .Z(n36348) );
  NANDN U36594 ( .A(n36347), .B(n36348), .Z(n36211) );
  AND U36595 ( .A(n36212), .B(n36211), .Z(n36340) );
  NANDN U36596 ( .A(n38247), .B(n36213), .Z(n36215) );
  XOR U36597 ( .A(b[61]), .B(a[104]), .Z(n36344) );
  NANDN U36598 ( .A(n38248), .B(n36344), .Z(n36214) );
  AND U36599 ( .A(n36215), .B(n36214), .Z(n36339) );
  NANDN U36600 ( .A(n37526), .B(n36216), .Z(n36218) );
  XOR U36601 ( .A(b[51]), .B(a[114]), .Z(n36324) );
  NANDN U36602 ( .A(n37605), .B(n36324), .Z(n36217) );
  NAND U36603 ( .A(n36218), .B(n36217), .Z(n36338) );
  XOR U36604 ( .A(n36339), .B(n36338), .Z(n36341) );
  XNOR U36605 ( .A(n36340), .B(n36341), .Z(n36399) );
  XNOR U36606 ( .A(n36400), .B(n36399), .Z(n36401) );
  NANDN U36607 ( .A(n36220), .B(n36219), .Z(n36224) );
  OR U36608 ( .A(n36222), .B(n36221), .Z(n36223) );
  NAND U36609 ( .A(n36224), .B(n36223), .Z(n36402) );
  XNOR U36610 ( .A(n36401), .B(n36402), .Z(n36298) );
  NANDN U36611 ( .A(n38090), .B(n36225), .Z(n36227) );
  XOR U36612 ( .A(b[59]), .B(a[106]), .Z(n36335) );
  NANDN U36613 ( .A(n38130), .B(n36335), .Z(n36226) );
  AND U36614 ( .A(n36227), .B(n36226), .Z(n36312) );
  NANDN U36615 ( .A(n36480), .B(n36228), .Z(n36230) );
  XOR U36616 ( .A(a[124]), .B(b[41]), .Z(n36332) );
  NANDN U36617 ( .A(n36594), .B(n36332), .Z(n36229) );
  AND U36618 ( .A(n36230), .B(n36229), .Z(n36311) );
  NANDN U36619 ( .A(n37705), .B(n36231), .Z(n36233) );
  XOR U36620 ( .A(b[53]), .B(a[112]), .Z(n36351) );
  NANDN U36621 ( .A(n37778), .B(n36351), .Z(n36232) );
  NAND U36622 ( .A(n36233), .B(n36232), .Z(n36310) );
  XOR U36623 ( .A(n36311), .B(n36310), .Z(n36313) );
  XOR U36624 ( .A(n36312), .B(n36313), .Z(n36394) );
  NANDN U36625 ( .A(n38278), .B(n36234), .Z(n36236) );
  XOR U36626 ( .A(b[63]), .B(a[102]), .Z(n36321) );
  NANDN U36627 ( .A(n38279), .B(n36321), .Z(n36235) );
  AND U36628 ( .A(n36236), .B(n36235), .Z(n36318) );
  NAND U36629 ( .A(b[63]), .B(a[100]), .Z(n36328) );
  ANDN U36630 ( .B(n36238), .A(n36237), .Z(n36241) );
  NAND U36631 ( .A(b[37]), .B(n36239), .Z(n36240) );
  NANDN U36632 ( .A(n36241), .B(n36240), .Z(n36316) );
  XOR U36633 ( .A(n36328), .B(n36316), .Z(n36317) );
  XOR U36634 ( .A(n36318), .B(n36317), .Z(n36393) );
  XNOR U36635 ( .A(n36394), .B(n36393), .Z(n36395) );
  NANDN U36636 ( .A(n36243), .B(n36242), .Z(n36247) );
  OR U36637 ( .A(n36245), .B(n36244), .Z(n36246) );
  NAND U36638 ( .A(n36247), .B(n36246), .Z(n36396) );
  XOR U36639 ( .A(n36395), .B(n36396), .Z(n36299) );
  XNOR U36640 ( .A(n36298), .B(n36299), .Z(n36301) );
  NANDN U36641 ( .A(n36249), .B(n36248), .Z(n36253) );
  OR U36642 ( .A(n36251), .B(n36250), .Z(n36252) );
  AND U36643 ( .A(n36253), .B(n36252), .Z(n36300) );
  XOR U36644 ( .A(n36301), .B(n36300), .Z(n36293) );
  NANDN U36645 ( .A(n36255), .B(n36254), .Z(n36259) );
  NANDN U36646 ( .A(n36257), .B(n36256), .Z(n36258) );
  AND U36647 ( .A(n36259), .B(n36258), .Z(n36292) );
  XOR U36648 ( .A(n36293), .B(n36292), .Z(n36295) );
  XOR U36649 ( .A(n36294), .B(n36295), .Z(n36288) );
  NANDN U36650 ( .A(n36261), .B(n36260), .Z(n36265) );
  NAND U36651 ( .A(n36263), .B(n36262), .Z(n36264) );
  AND U36652 ( .A(n36265), .B(n36264), .Z(n36287) );
  NANDN U36653 ( .A(n36267), .B(n36266), .Z(n36271) );
  OR U36654 ( .A(n36269), .B(n36268), .Z(n36270) );
  NAND U36655 ( .A(n36271), .B(n36270), .Z(n36286) );
  XOR U36656 ( .A(n36287), .B(n36286), .Z(n36289) );
  XNOR U36657 ( .A(n36288), .B(n36289), .Z(n36405) );
  XNOR U36658 ( .A(n36406), .B(n36405), .Z(n36408) );
  NANDN U36659 ( .A(n36273), .B(n36272), .Z(n36277) );
  NANDN U36660 ( .A(n36275), .B(n36274), .Z(n36276) );
  AND U36661 ( .A(n36277), .B(n36276), .Z(n36407) );
  XNOR U36662 ( .A(n36408), .B(n36407), .Z(n36280) );
  XOR U36663 ( .A(n36281), .B(n36280), .Z(n36283) );
  XNOR U36664 ( .A(n36282), .B(n36283), .Z(n36278) );
  XOR U36665 ( .A(n36279), .B(n36278), .Z(c[228]) );
  AND U36666 ( .A(n36279), .B(n36278), .Z(n36412) );
  NANDN U36667 ( .A(n36281), .B(n36280), .Z(n36285) );
  OR U36668 ( .A(n36283), .B(n36282), .Z(n36284) );
  AND U36669 ( .A(n36285), .B(n36284), .Z(n36415) );
  NANDN U36670 ( .A(n36287), .B(n36286), .Z(n36291) );
  OR U36671 ( .A(n36289), .B(n36288), .Z(n36290) );
  AND U36672 ( .A(n36291), .B(n36290), .Z(n36422) );
  NANDN U36673 ( .A(n36293), .B(n36292), .Z(n36297) );
  OR U36674 ( .A(n36295), .B(n36294), .Z(n36296) );
  AND U36675 ( .A(n36297), .B(n36296), .Z(n36419) );
  NANDN U36676 ( .A(n36299), .B(n36298), .Z(n36303) );
  NAND U36677 ( .A(n36301), .B(n36300), .Z(n36302) );
  AND U36678 ( .A(n36303), .B(n36302), .Z(n36434) );
  NANDN U36679 ( .A(n36305), .B(n36304), .Z(n36309) );
  NANDN U36680 ( .A(n36307), .B(n36306), .Z(n36308) );
  AND U36681 ( .A(n36309), .B(n36308), .Z(n36507) );
  NANDN U36682 ( .A(n36311), .B(n36310), .Z(n36315) );
  OR U36683 ( .A(n36313), .B(n36312), .Z(n36314) );
  NAND U36684 ( .A(n36315), .B(n36314), .Z(n36506) );
  XNOR U36685 ( .A(n36507), .B(n36506), .Z(n36509) );
  IV U36686 ( .A(n36328), .Z(n36527) );
  NANDN U36687 ( .A(n36527), .B(n36316), .Z(n36320) );
  NANDN U36688 ( .A(n36318), .B(n36317), .Z(n36319) );
  AND U36689 ( .A(n36320), .B(n36319), .Z(n36458) );
  NANDN U36690 ( .A(n38278), .B(n36321), .Z(n36323) );
  XOR U36691 ( .A(b[63]), .B(a[103]), .Z(n36486) );
  NANDN U36692 ( .A(n38279), .B(n36486), .Z(n36322) );
  AND U36693 ( .A(n36323), .B(n36322), .Z(n36495) );
  NANDN U36694 ( .A(n37526), .B(n36324), .Z(n36326) );
  XOR U36695 ( .A(b[51]), .B(a[115]), .Z(n36464) );
  NANDN U36696 ( .A(n37605), .B(n36464), .Z(n36325) );
  NAND U36697 ( .A(n36326), .B(n36325), .Z(n36494) );
  XNOR U36698 ( .A(n36495), .B(n36494), .Z(n36496) );
  IV U36699 ( .A(n36327), .Z(n36525) );
  AND U36700 ( .A(b[63]), .B(a[101]), .Z(n36524) );
  XOR U36701 ( .A(n36525), .B(n36524), .Z(n36526) );
  XOR U36702 ( .A(n36328), .B(n36526), .Z(n36497) );
  XOR U36703 ( .A(n36496), .B(n36497), .Z(n36455) );
  NANDN U36704 ( .A(n37857), .B(n36329), .Z(n36331) );
  XOR U36705 ( .A(b[55]), .B(a[111]), .Z(n36461) );
  NANDN U36706 ( .A(n37911), .B(n36461), .Z(n36330) );
  AND U36707 ( .A(n36331), .B(n36330), .Z(n36521) );
  NANDN U36708 ( .A(n36480), .B(n36332), .Z(n36334) );
  XOR U36709 ( .A(a[125]), .B(b[41]), .Z(n36479) );
  NANDN U36710 ( .A(n36594), .B(n36479), .Z(n36333) );
  AND U36711 ( .A(n36334), .B(n36333), .Z(n36519) );
  NANDN U36712 ( .A(n38090), .B(n36335), .Z(n36337) );
  XOR U36713 ( .A(b[59]), .B(a[107]), .Z(n36467) );
  NANDN U36714 ( .A(n38130), .B(n36467), .Z(n36336) );
  NAND U36715 ( .A(n36337), .B(n36336), .Z(n36518) );
  XNOR U36716 ( .A(n36519), .B(n36518), .Z(n36520) );
  XOR U36717 ( .A(n36521), .B(n36520), .Z(n36456) );
  XNOR U36718 ( .A(n36455), .B(n36456), .Z(n36457) );
  XNOR U36719 ( .A(n36458), .B(n36457), .Z(n36508) );
  XOR U36720 ( .A(n36509), .B(n36508), .Z(n36446) );
  NANDN U36721 ( .A(n36339), .B(n36338), .Z(n36343) );
  OR U36722 ( .A(n36341), .B(n36340), .Z(n36342) );
  AND U36723 ( .A(n36343), .B(n36342), .Z(n36450) );
  NANDN U36724 ( .A(n38247), .B(n36344), .Z(n36346) );
  XOR U36725 ( .A(b[61]), .B(a[105]), .Z(n36470) );
  NANDN U36726 ( .A(n38248), .B(n36470), .Z(n36345) );
  AND U36727 ( .A(n36346), .B(n36345), .Z(n36542) );
  XNOR U36728 ( .A(a[127]), .B(b[39]), .Z(n36489) );
  OR U36729 ( .A(n36489), .B(n36347), .Z(n36350) );
  NAND U36730 ( .A(n36490), .B(n36348), .Z(n36349) );
  AND U36731 ( .A(n36350), .B(n36349), .Z(n36540) );
  NANDN U36732 ( .A(n37705), .B(n36351), .Z(n36353) );
  XOR U36733 ( .A(b[53]), .B(a[113]), .Z(n36483) );
  NANDN U36734 ( .A(n37778), .B(n36483), .Z(n36352) );
  NAND U36735 ( .A(n36353), .B(n36352), .Z(n36539) );
  XNOR U36736 ( .A(n36540), .B(n36539), .Z(n36541) );
  XNOR U36737 ( .A(n36542), .B(n36541), .Z(n36449) );
  XNOR U36738 ( .A(n36450), .B(n36449), .Z(n36452) );
  NANDN U36739 ( .A(n211), .B(n36354), .Z(n36356) );
  XOR U36740 ( .A(a[119]), .B(b[47]), .Z(n36530) );
  NANDN U36741 ( .A(n37172), .B(n36530), .Z(n36355) );
  AND U36742 ( .A(n36356), .B(n36355), .Z(n36515) );
  NANDN U36743 ( .A(n36991), .B(n36357), .Z(n36359) );
  XOR U36744 ( .A(a[121]), .B(b[45]), .Z(n36533) );
  NANDN U36745 ( .A(n37083), .B(n36533), .Z(n36358) );
  AND U36746 ( .A(n36359), .B(n36358), .Z(n36513) );
  NANDN U36747 ( .A(n212), .B(n36360), .Z(n36362) );
  XOR U36748 ( .A(a[117]), .B(b[49]), .Z(n36473) );
  NANDN U36749 ( .A(n37432), .B(n36473), .Z(n36361) );
  AND U36750 ( .A(n36362), .B(n36361), .Z(n36503) );
  NANDN U36751 ( .A(n37974), .B(n36363), .Z(n36365) );
  XOR U36752 ( .A(b[57]), .B(a[109]), .Z(n36536) );
  NANDN U36753 ( .A(n38031), .B(n36536), .Z(n36364) );
  AND U36754 ( .A(n36365), .B(n36364), .Z(n36501) );
  NANDN U36755 ( .A(n36742), .B(n36366), .Z(n36368) );
  XOR U36756 ( .A(a[123]), .B(b[43]), .Z(n36476) );
  NANDN U36757 ( .A(n36891), .B(n36476), .Z(n36367) );
  NAND U36758 ( .A(n36368), .B(n36367), .Z(n36500) );
  XNOR U36759 ( .A(n36501), .B(n36500), .Z(n36502) );
  XNOR U36760 ( .A(n36503), .B(n36502), .Z(n36512) );
  XNOR U36761 ( .A(n36513), .B(n36512), .Z(n36514) );
  XNOR U36762 ( .A(n36515), .B(n36514), .Z(n36451) );
  XOR U36763 ( .A(n36452), .B(n36451), .Z(n36444) );
  NANDN U36764 ( .A(n36370), .B(n36369), .Z(n36374) );
  OR U36765 ( .A(n36372), .B(n36371), .Z(n36373) );
  AND U36766 ( .A(n36374), .B(n36373), .Z(n36443) );
  XNOR U36767 ( .A(n36444), .B(n36443), .Z(n36445) );
  XNOR U36768 ( .A(n36446), .B(n36445), .Z(n36431) );
  NAND U36769 ( .A(n36376), .B(n36375), .Z(n36380) );
  NAND U36770 ( .A(n36378), .B(n36377), .Z(n36379) );
  NAND U36771 ( .A(n36380), .B(n36379), .Z(n36432) );
  XNOR U36772 ( .A(n36431), .B(n36432), .Z(n36433) );
  XNOR U36773 ( .A(n36434), .B(n36433), .Z(n36427) );
  NANDN U36774 ( .A(n36382), .B(n36381), .Z(n36386) );
  OR U36775 ( .A(n36384), .B(n36383), .Z(n36385) );
  AND U36776 ( .A(n36386), .B(n36385), .Z(n36426) );
  NANDN U36777 ( .A(n36388), .B(n36387), .Z(n36392) );
  NAND U36778 ( .A(n36390), .B(n36389), .Z(n36391) );
  AND U36779 ( .A(n36392), .B(n36391), .Z(n36439) );
  NANDN U36780 ( .A(n36394), .B(n36393), .Z(n36398) );
  NANDN U36781 ( .A(n36396), .B(n36395), .Z(n36397) );
  AND U36782 ( .A(n36398), .B(n36397), .Z(n36438) );
  NANDN U36783 ( .A(n36400), .B(n36399), .Z(n36404) );
  NANDN U36784 ( .A(n36402), .B(n36401), .Z(n36403) );
  NAND U36785 ( .A(n36404), .B(n36403), .Z(n36437) );
  XOR U36786 ( .A(n36438), .B(n36437), .Z(n36440) );
  XNOR U36787 ( .A(n36439), .B(n36440), .Z(n36425) );
  XOR U36788 ( .A(n36426), .B(n36425), .Z(n36428) );
  XOR U36789 ( .A(n36427), .B(n36428), .Z(n36420) );
  XNOR U36790 ( .A(n36419), .B(n36420), .Z(n36421) );
  XNOR U36791 ( .A(n36422), .B(n36421), .Z(n36413) );
  NANDN U36792 ( .A(n36406), .B(n36405), .Z(n36410) );
  NAND U36793 ( .A(n36408), .B(n36407), .Z(n36409) );
  NAND U36794 ( .A(n36410), .B(n36409), .Z(n36414) );
  XOR U36795 ( .A(n36413), .B(n36414), .Z(n36416) );
  XNOR U36796 ( .A(n36415), .B(n36416), .Z(n36411) );
  XOR U36797 ( .A(n36412), .B(n36411), .Z(c[229]) );
  AND U36798 ( .A(n36412), .B(n36411), .Z(n36546) );
  NANDN U36799 ( .A(n36414), .B(n36413), .Z(n36418) );
  OR U36800 ( .A(n36416), .B(n36415), .Z(n36417) );
  AND U36801 ( .A(n36418), .B(n36417), .Z(n36549) );
  NANDN U36802 ( .A(n36420), .B(n36419), .Z(n36424) );
  NANDN U36803 ( .A(n36422), .B(n36421), .Z(n36423) );
  AND U36804 ( .A(n36424), .B(n36423), .Z(n36548) );
  NANDN U36805 ( .A(n36426), .B(n36425), .Z(n36430) );
  NANDN U36806 ( .A(n36428), .B(n36427), .Z(n36429) );
  AND U36807 ( .A(n36430), .B(n36429), .Z(n36556) );
  NANDN U36808 ( .A(n36432), .B(n36431), .Z(n36436) );
  NANDN U36809 ( .A(n36434), .B(n36433), .Z(n36435) );
  AND U36810 ( .A(n36436), .B(n36435), .Z(n36554) );
  NANDN U36811 ( .A(n36438), .B(n36437), .Z(n36442) );
  NANDN U36812 ( .A(n36440), .B(n36439), .Z(n36441) );
  AND U36813 ( .A(n36442), .B(n36441), .Z(n36562) );
  NANDN U36814 ( .A(n36444), .B(n36443), .Z(n36448) );
  NANDN U36815 ( .A(n36446), .B(n36445), .Z(n36447) );
  AND U36816 ( .A(n36448), .B(n36447), .Z(n36560) );
  NANDN U36817 ( .A(n36450), .B(n36449), .Z(n36454) );
  NAND U36818 ( .A(n36452), .B(n36451), .Z(n36453) );
  AND U36819 ( .A(n36454), .B(n36453), .Z(n36664) );
  NANDN U36820 ( .A(n36456), .B(n36455), .Z(n36460) );
  NANDN U36821 ( .A(n36458), .B(n36457), .Z(n36459) );
  AND U36822 ( .A(n36460), .B(n36459), .Z(n36663) );
  NANDN U36823 ( .A(n37857), .B(n36461), .Z(n36463) );
  XOR U36824 ( .A(b[55]), .B(a[112]), .Z(n36608) );
  NANDN U36825 ( .A(n37911), .B(n36608), .Z(n36462) );
  AND U36826 ( .A(n36463), .B(n36462), .Z(n36640) );
  NANDN U36827 ( .A(n37526), .B(n36464), .Z(n36466) );
  XOR U36828 ( .A(b[51]), .B(a[116]), .Z(n36629) );
  NANDN U36829 ( .A(n37605), .B(n36629), .Z(n36465) );
  AND U36830 ( .A(n36466), .B(n36465), .Z(n36639) );
  NANDN U36831 ( .A(n38090), .B(n36467), .Z(n36469) );
  XOR U36832 ( .A(b[59]), .B(a[108]), .Z(n36617) );
  NANDN U36833 ( .A(n38130), .B(n36617), .Z(n36468) );
  AND U36834 ( .A(n36469), .B(n36468), .Z(n36586) );
  NANDN U36835 ( .A(n38247), .B(n36470), .Z(n36472) );
  XOR U36836 ( .A(b[61]), .B(a[106]), .Z(n36602) );
  NANDN U36837 ( .A(n38248), .B(n36602), .Z(n36471) );
  AND U36838 ( .A(n36472), .B(n36471), .Z(n36584) );
  NANDN U36839 ( .A(n212), .B(n36473), .Z(n36475) );
  XOR U36840 ( .A(a[118]), .B(b[49]), .Z(n36626) );
  NANDN U36841 ( .A(n37432), .B(n36626), .Z(n36474) );
  NAND U36842 ( .A(n36475), .B(n36474), .Z(n36583) );
  XNOR U36843 ( .A(n36584), .B(n36583), .Z(n36585) );
  XNOR U36844 ( .A(n36586), .B(n36585), .Z(n36638) );
  XOR U36845 ( .A(n36639), .B(n36638), .Z(n36641) );
  XOR U36846 ( .A(n36640), .B(n36641), .Z(n36658) );
  NANDN U36847 ( .A(n36742), .B(n36476), .Z(n36478) );
  XOR U36848 ( .A(a[124]), .B(b[43]), .Z(n36620) );
  NANDN U36849 ( .A(n36891), .B(n36620), .Z(n36477) );
  AND U36850 ( .A(n36478), .B(n36477), .Z(n36579) );
  NANDN U36851 ( .A(n36480), .B(n36479), .Z(n36482) );
  XOR U36852 ( .A(a[126]), .B(b[41]), .Z(n36595) );
  NANDN U36853 ( .A(n36594), .B(n36595), .Z(n36481) );
  AND U36854 ( .A(n36482), .B(n36481), .Z(n36578) );
  NANDN U36855 ( .A(n37705), .B(n36483), .Z(n36485) );
  XOR U36856 ( .A(b[53]), .B(a[114]), .Z(n36598) );
  NANDN U36857 ( .A(n37778), .B(n36598), .Z(n36484) );
  NAND U36858 ( .A(n36485), .B(n36484), .Z(n36577) );
  XOR U36859 ( .A(n36578), .B(n36577), .Z(n36580) );
  XOR U36860 ( .A(n36579), .B(n36580), .Z(n36657) );
  NANDN U36861 ( .A(n38278), .B(n36486), .Z(n36488) );
  XOR U36862 ( .A(b[63]), .B(a[104]), .Z(n36605) );
  NANDN U36863 ( .A(n38279), .B(n36605), .Z(n36487) );
  AND U36864 ( .A(n36488), .B(n36487), .Z(n36591) );
  NAND U36865 ( .A(b[63]), .B(a[102]), .Z(n36601) );
  ANDN U36866 ( .B(n36490), .A(n36489), .Z(n36493) );
  NAND U36867 ( .A(b[39]), .B(n36491), .Z(n36492) );
  NANDN U36868 ( .A(n36493), .B(n36492), .Z(n36589) );
  XOR U36869 ( .A(n36601), .B(n36589), .Z(n36590) );
  XOR U36870 ( .A(n36591), .B(n36590), .Z(n36656) );
  XOR U36871 ( .A(n36657), .B(n36656), .Z(n36659) );
  XOR U36872 ( .A(n36658), .B(n36659), .Z(n36647) );
  NANDN U36873 ( .A(n36495), .B(n36494), .Z(n36499) );
  NAND U36874 ( .A(n36497), .B(n36496), .Z(n36498) );
  AND U36875 ( .A(n36499), .B(n36498), .Z(n36645) );
  NANDN U36876 ( .A(n36501), .B(n36500), .Z(n36505) );
  NANDN U36877 ( .A(n36503), .B(n36502), .Z(n36504) );
  NAND U36878 ( .A(n36505), .B(n36504), .Z(n36644) );
  XNOR U36879 ( .A(n36645), .B(n36644), .Z(n36646) );
  XNOR U36880 ( .A(n36647), .B(n36646), .Z(n36662) );
  XOR U36881 ( .A(n36663), .B(n36662), .Z(n36665) );
  XOR U36882 ( .A(n36664), .B(n36665), .Z(n36568) );
  NANDN U36883 ( .A(n36507), .B(n36506), .Z(n36511) );
  NAND U36884 ( .A(n36509), .B(n36508), .Z(n36510) );
  AND U36885 ( .A(n36511), .B(n36510), .Z(n36565) );
  NANDN U36886 ( .A(n36513), .B(n36512), .Z(n36517) );
  NANDN U36887 ( .A(n36515), .B(n36514), .Z(n36516) );
  AND U36888 ( .A(n36517), .B(n36516), .Z(n36573) );
  NANDN U36889 ( .A(n36519), .B(n36518), .Z(n36523) );
  NANDN U36890 ( .A(n36521), .B(n36520), .Z(n36522) );
  AND U36891 ( .A(n36523), .B(n36522), .Z(n36652) );
  NANDN U36892 ( .A(n36525), .B(n36524), .Z(n36529) );
  ANDN U36893 ( .B(n36527), .A(n36526), .Z(n36528) );
  ANDN U36894 ( .B(n36529), .A(n36528), .Z(n36651) );
  NANDN U36895 ( .A(n211), .B(n36530), .Z(n36532) );
  XOR U36896 ( .A(a[120]), .B(b[47]), .Z(n36635) );
  NANDN U36897 ( .A(n37172), .B(n36635), .Z(n36531) );
  AND U36898 ( .A(n36532), .B(n36531), .Z(n36614) );
  NANDN U36899 ( .A(n36991), .B(n36533), .Z(n36535) );
  XOR U36900 ( .A(a[122]), .B(b[45]), .Z(n36632) );
  NANDN U36901 ( .A(n37083), .B(n36632), .Z(n36534) );
  AND U36902 ( .A(n36535), .B(n36534), .Z(n36612) );
  NANDN U36903 ( .A(n37974), .B(n36536), .Z(n36538) );
  XOR U36904 ( .A(b[57]), .B(a[110]), .Z(n36623) );
  NANDN U36905 ( .A(n38031), .B(n36623), .Z(n36537) );
  NAND U36906 ( .A(n36538), .B(n36537), .Z(n36611) );
  XNOR U36907 ( .A(n36612), .B(n36611), .Z(n36613) );
  XNOR U36908 ( .A(n36614), .B(n36613), .Z(n36650) );
  XOR U36909 ( .A(n36651), .B(n36650), .Z(n36653) );
  XOR U36910 ( .A(n36652), .B(n36653), .Z(n36572) );
  NANDN U36911 ( .A(n36540), .B(n36539), .Z(n36544) );
  NANDN U36912 ( .A(n36542), .B(n36541), .Z(n36543) );
  AND U36913 ( .A(n36544), .B(n36543), .Z(n36571) );
  XOR U36914 ( .A(n36572), .B(n36571), .Z(n36574) );
  XOR U36915 ( .A(n36573), .B(n36574), .Z(n36566) );
  XNOR U36916 ( .A(n36565), .B(n36566), .Z(n36567) );
  XNOR U36917 ( .A(n36568), .B(n36567), .Z(n36559) );
  XNOR U36918 ( .A(n36560), .B(n36559), .Z(n36561) );
  XNOR U36919 ( .A(n36562), .B(n36561), .Z(n36553) );
  XNOR U36920 ( .A(n36554), .B(n36553), .Z(n36555) );
  XNOR U36921 ( .A(n36556), .B(n36555), .Z(n36547) );
  XOR U36922 ( .A(n36548), .B(n36547), .Z(n36550) );
  XNOR U36923 ( .A(n36549), .B(n36550), .Z(n36545) );
  XOR U36924 ( .A(n36546), .B(n36545), .Z(c[230]) );
  AND U36925 ( .A(n36546), .B(n36545), .Z(n36669) );
  NANDN U36926 ( .A(n36548), .B(n36547), .Z(n36552) );
  OR U36927 ( .A(n36550), .B(n36549), .Z(n36551) );
  AND U36928 ( .A(n36552), .B(n36551), .Z(n36672) );
  NANDN U36929 ( .A(n36554), .B(n36553), .Z(n36558) );
  NANDN U36930 ( .A(n36556), .B(n36555), .Z(n36557) );
  AND U36931 ( .A(n36558), .B(n36557), .Z(n36671) );
  NANDN U36932 ( .A(n36560), .B(n36559), .Z(n36564) );
  NANDN U36933 ( .A(n36562), .B(n36561), .Z(n36563) );
  AND U36934 ( .A(n36564), .B(n36563), .Z(n36679) );
  NANDN U36935 ( .A(n36566), .B(n36565), .Z(n36570) );
  NANDN U36936 ( .A(n36568), .B(n36567), .Z(n36569) );
  AND U36937 ( .A(n36570), .B(n36569), .Z(n36677) );
  NANDN U36938 ( .A(n36572), .B(n36571), .Z(n36576) );
  NANDN U36939 ( .A(n36574), .B(n36573), .Z(n36575) );
  AND U36940 ( .A(n36576), .B(n36575), .Z(n36790) );
  NANDN U36941 ( .A(n36578), .B(n36577), .Z(n36582) );
  OR U36942 ( .A(n36580), .B(n36579), .Z(n36581) );
  AND U36943 ( .A(n36582), .B(n36581), .Z(n36764) );
  NANDN U36944 ( .A(n36584), .B(n36583), .Z(n36588) );
  NANDN U36945 ( .A(n36586), .B(n36585), .Z(n36587) );
  NAND U36946 ( .A(n36588), .B(n36587), .Z(n36763) );
  XNOR U36947 ( .A(n36764), .B(n36763), .Z(n36766) );
  IV U36948 ( .A(n36601), .Z(n36730) );
  NANDN U36949 ( .A(n36730), .B(n36589), .Z(n36593) );
  NANDN U36950 ( .A(n36591), .B(n36590), .Z(n36592) );
  AND U36951 ( .A(n36593), .B(n36592), .Z(n36778) );
  XNOR U36952 ( .A(a[127]), .B(b[41]), .Z(n36734) );
  OR U36953 ( .A(n36734), .B(n36594), .Z(n36597) );
  NAND U36954 ( .A(n36735), .B(n36595), .Z(n36596) );
  AND U36955 ( .A(n36597), .B(n36596), .Z(n36752) );
  NANDN U36956 ( .A(n37705), .B(n36598), .Z(n36600) );
  XOR U36957 ( .A(b[53]), .B(a[115]), .Z(n36748) );
  NANDN U36958 ( .A(n37778), .B(n36748), .Z(n36599) );
  NAND U36959 ( .A(n36600), .B(n36599), .Z(n36751) );
  XNOR U36960 ( .A(n36752), .B(n36751), .Z(n36753) );
  AND U36961 ( .A(b[63]), .B(a[103]), .Z(n36727) );
  XOR U36962 ( .A(n36728), .B(n36727), .Z(n36729) );
  XOR U36963 ( .A(n36601), .B(n36729), .Z(n36754) );
  XOR U36964 ( .A(n36753), .B(n36754), .Z(n36775) );
  NANDN U36965 ( .A(n38247), .B(n36602), .Z(n36604) );
  XOR U36966 ( .A(b[61]), .B(a[107]), .Z(n36745) );
  NANDN U36967 ( .A(n38248), .B(n36745), .Z(n36603) );
  AND U36968 ( .A(n36604), .B(n36603), .Z(n36718) );
  NANDN U36969 ( .A(n38278), .B(n36605), .Z(n36607) );
  XOR U36970 ( .A(b[63]), .B(a[105]), .Z(n36738) );
  NANDN U36971 ( .A(n38279), .B(n36738), .Z(n36606) );
  AND U36972 ( .A(n36607), .B(n36606), .Z(n36716) );
  NANDN U36973 ( .A(n37857), .B(n36608), .Z(n36610) );
  XOR U36974 ( .A(b[55]), .B(a[113]), .Z(n36700) );
  NANDN U36975 ( .A(n37911), .B(n36700), .Z(n36609) );
  NAND U36976 ( .A(n36610), .B(n36609), .Z(n36715) );
  XNOR U36977 ( .A(n36716), .B(n36715), .Z(n36717) );
  XOR U36978 ( .A(n36718), .B(n36717), .Z(n36776) );
  XNOR U36979 ( .A(n36775), .B(n36776), .Z(n36777) );
  XNOR U36980 ( .A(n36778), .B(n36777), .Z(n36765) );
  XOR U36981 ( .A(n36766), .B(n36765), .Z(n36788) );
  NANDN U36982 ( .A(n36612), .B(n36611), .Z(n36616) );
  NANDN U36983 ( .A(n36614), .B(n36613), .Z(n36615) );
  AND U36984 ( .A(n36616), .B(n36615), .Z(n36688) );
  NANDN U36985 ( .A(n38090), .B(n36617), .Z(n36619) );
  XOR U36986 ( .A(b[59]), .B(a[109]), .Z(n36697) );
  NANDN U36987 ( .A(n38130), .B(n36697), .Z(n36618) );
  AND U36988 ( .A(n36619), .B(n36618), .Z(n36723) );
  NANDN U36989 ( .A(n36742), .B(n36620), .Z(n36622) );
  XOR U36990 ( .A(a[125]), .B(b[43]), .Z(n36741) );
  NANDN U36991 ( .A(n36891), .B(n36741), .Z(n36621) );
  AND U36992 ( .A(n36622), .B(n36621), .Z(n36722) );
  NANDN U36993 ( .A(n37974), .B(n36623), .Z(n36625) );
  XOR U36994 ( .A(b[57]), .B(a[111]), .Z(n36694) );
  NANDN U36995 ( .A(n38031), .B(n36694), .Z(n36624) );
  NAND U36996 ( .A(n36625), .B(n36624), .Z(n36721) );
  XOR U36997 ( .A(n36722), .B(n36721), .Z(n36724) );
  XOR U36998 ( .A(n36723), .B(n36724), .Z(n36772) );
  NANDN U36999 ( .A(n212), .B(n36626), .Z(n36628) );
  XNOR U37000 ( .A(a[119]), .B(b[49]), .Z(n36712) );
  NANDN U37001 ( .A(n36712), .B(n37537), .Z(n36627) );
  AND U37002 ( .A(n36628), .B(n36627), .Z(n36759) );
  NANDN U37003 ( .A(n37526), .B(n36629), .Z(n36631) );
  XOR U37004 ( .A(b[51]), .B(a[117]), .Z(n36706) );
  NANDN U37005 ( .A(n37605), .B(n36706), .Z(n36630) );
  AND U37006 ( .A(n36631), .B(n36630), .Z(n36758) );
  NANDN U37007 ( .A(n36991), .B(n36632), .Z(n36634) );
  XOR U37008 ( .A(a[123]), .B(b[45]), .Z(n36709) );
  NANDN U37009 ( .A(n37083), .B(n36709), .Z(n36633) );
  NAND U37010 ( .A(n36634), .B(n36633), .Z(n36757) );
  XOR U37011 ( .A(n36758), .B(n36757), .Z(n36760) );
  XOR U37012 ( .A(n36759), .B(n36760), .Z(n36770) );
  NAND U37013 ( .A(n37294), .B(n36635), .Z(n36637) );
  XNOR U37014 ( .A(a[121]), .B(b[47]), .Z(n36703) );
  NANDN U37015 ( .A(n36703), .B(n37341), .Z(n36636) );
  AND U37016 ( .A(n36637), .B(n36636), .Z(n36769) );
  XNOR U37017 ( .A(n36770), .B(n36769), .Z(n36771) );
  XOR U37018 ( .A(n36772), .B(n36771), .Z(n36689) );
  XNOR U37019 ( .A(n36688), .B(n36689), .Z(n36690) );
  NANDN U37020 ( .A(n36639), .B(n36638), .Z(n36643) );
  OR U37021 ( .A(n36641), .B(n36640), .Z(n36642) );
  NAND U37022 ( .A(n36643), .B(n36642), .Z(n36691) );
  XNOR U37023 ( .A(n36690), .B(n36691), .Z(n36787) );
  XNOR U37024 ( .A(n36788), .B(n36787), .Z(n36789) );
  XNOR U37025 ( .A(n36790), .B(n36789), .Z(n36684) );
  NANDN U37026 ( .A(n36645), .B(n36644), .Z(n36649) );
  NANDN U37027 ( .A(n36647), .B(n36646), .Z(n36648) );
  AND U37028 ( .A(n36649), .B(n36648), .Z(n36783) );
  NANDN U37029 ( .A(n36651), .B(n36650), .Z(n36655) );
  OR U37030 ( .A(n36653), .B(n36652), .Z(n36654) );
  AND U37031 ( .A(n36655), .B(n36654), .Z(n36782) );
  NANDN U37032 ( .A(n36657), .B(n36656), .Z(n36661) );
  OR U37033 ( .A(n36659), .B(n36658), .Z(n36660) );
  AND U37034 ( .A(n36661), .B(n36660), .Z(n36781) );
  XOR U37035 ( .A(n36782), .B(n36781), .Z(n36784) );
  XOR U37036 ( .A(n36783), .B(n36784), .Z(n36683) );
  NANDN U37037 ( .A(n36663), .B(n36662), .Z(n36667) );
  OR U37038 ( .A(n36665), .B(n36664), .Z(n36666) );
  AND U37039 ( .A(n36667), .B(n36666), .Z(n36682) );
  XOR U37040 ( .A(n36683), .B(n36682), .Z(n36685) );
  XNOR U37041 ( .A(n36684), .B(n36685), .Z(n36676) );
  XNOR U37042 ( .A(n36677), .B(n36676), .Z(n36678) );
  XNOR U37043 ( .A(n36679), .B(n36678), .Z(n36670) );
  XOR U37044 ( .A(n36671), .B(n36670), .Z(n36673) );
  XNOR U37045 ( .A(n36672), .B(n36673), .Z(n36668) );
  XOR U37046 ( .A(n36669), .B(n36668), .Z(c[231]) );
  AND U37047 ( .A(n36669), .B(n36668), .Z(n36794) );
  NANDN U37048 ( .A(n36671), .B(n36670), .Z(n36675) );
  OR U37049 ( .A(n36673), .B(n36672), .Z(n36674) );
  AND U37050 ( .A(n36675), .B(n36674), .Z(n36797) );
  NANDN U37051 ( .A(n36677), .B(n36676), .Z(n36681) );
  NANDN U37052 ( .A(n36679), .B(n36678), .Z(n36680) );
  AND U37053 ( .A(n36681), .B(n36680), .Z(n36796) );
  NANDN U37054 ( .A(n36683), .B(n36682), .Z(n36687) );
  NANDN U37055 ( .A(n36685), .B(n36684), .Z(n36686) );
  AND U37056 ( .A(n36687), .B(n36686), .Z(n36804) );
  NANDN U37057 ( .A(n36689), .B(n36688), .Z(n36693) );
  NANDN U37058 ( .A(n36691), .B(n36690), .Z(n36692) );
  AND U37059 ( .A(n36693), .B(n36692), .Z(n36815) );
  NANDN U37060 ( .A(n37974), .B(n36694), .Z(n36696) );
  XOR U37061 ( .A(b[57]), .B(a[112]), .Z(n36870) );
  NANDN U37062 ( .A(n38031), .B(n36870), .Z(n36695) );
  AND U37063 ( .A(n36696), .B(n36695), .Z(n36851) );
  NANDN U37064 ( .A(n38090), .B(n36697), .Z(n36699) );
  XOR U37065 ( .A(b[59]), .B(a[110]), .Z(n36873) );
  NANDN U37066 ( .A(n38130), .B(n36873), .Z(n36698) );
  AND U37067 ( .A(n36699), .B(n36698), .Z(n36850) );
  NANDN U37068 ( .A(n37857), .B(n36700), .Z(n36702) );
  XOR U37069 ( .A(b[55]), .B(a[114]), .Z(n36895) );
  NANDN U37070 ( .A(n37911), .B(n36895), .Z(n36701) );
  NAND U37071 ( .A(n36702), .B(n36701), .Z(n36849) );
  XOR U37072 ( .A(n36850), .B(n36849), .Z(n36852) );
  XOR U37073 ( .A(n36851), .B(n36852), .Z(n36833) );
  NANDN U37074 ( .A(n36703), .B(n37294), .Z(n36705) );
  XOR U37075 ( .A(a[122]), .B(b[47]), .Z(n36885) );
  NANDN U37076 ( .A(n37172), .B(n36885), .Z(n36704) );
  AND U37077 ( .A(n36705), .B(n36704), .Z(n36900) );
  NANDN U37078 ( .A(n37526), .B(n36706), .Z(n36708) );
  XOR U37079 ( .A(a[118]), .B(b[51]), .Z(n36876) );
  NANDN U37080 ( .A(n37605), .B(n36876), .Z(n36707) );
  AND U37081 ( .A(n36708), .B(n36707), .Z(n36899) );
  NANDN U37082 ( .A(n36991), .B(n36709), .Z(n36711) );
  XOR U37083 ( .A(a[124]), .B(b[45]), .Z(n36888) );
  NANDN U37084 ( .A(n37083), .B(n36888), .Z(n36710) );
  NAND U37085 ( .A(n36711), .B(n36710), .Z(n36898) );
  XOR U37086 ( .A(n36899), .B(n36898), .Z(n36901) );
  XOR U37087 ( .A(n36900), .B(n36901), .Z(n36832) );
  NANDN U37088 ( .A(n36712), .B(n37536), .Z(n36714) );
  XNOR U37089 ( .A(a[120]), .B(b[49]), .Z(n36882) );
  NANDN U37090 ( .A(n36882), .B(n37537), .Z(n36713) );
  AND U37091 ( .A(n36714), .B(n36713), .Z(n36831) );
  XOR U37092 ( .A(n36832), .B(n36831), .Z(n36834) );
  XOR U37093 ( .A(n36833), .B(n36834), .Z(n36821) );
  NANDN U37094 ( .A(n36716), .B(n36715), .Z(n36720) );
  NANDN U37095 ( .A(n36718), .B(n36717), .Z(n36719) );
  AND U37096 ( .A(n36720), .B(n36719), .Z(n36820) );
  NANDN U37097 ( .A(n36722), .B(n36721), .Z(n36726) );
  OR U37098 ( .A(n36724), .B(n36723), .Z(n36725) );
  AND U37099 ( .A(n36726), .B(n36725), .Z(n36846) );
  NANDN U37100 ( .A(n36728), .B(n36727), .Z(n36732) );
  ANDN U37101 ( .B(n36730), .A(n36729), .Z(n36731) );
  ANDN U37102 ( .B(n36732), .A(n36731), .Z(n36844) );
  NAND U37103 ( .A(b[41]), .B(n36733), .Z(n36737) );
  ANDN U37104 ( .B(n36735), .A(n36734), .Z(n36736) );
  ANDN U37105 ( .B(n36737), .A(n36736), .Z(n36857) );
  NAND U37106 ( .A(b[63]), .B(a[104]), .Z(n36942) );
  NANDN U37107 ( .A(n38278), .B(n36738), .Z(n36740) );
  XOR U37108 ( .A(b[63]), .B(a[106]), .Z(n36864) );
  NANDN U37109 ( .A(n38279), .B(n36864), .Z(n36739) );
  NAND U37110 ( .A(n36740), .B(n36739), .Z(n36855) );
  XOR U37111 ( .A(n36942), .B(n36855), .Z(n36856) );
  XNOR U37112 ( .A(n36857), .B(n36856), .Z(n36843) );
  XNOR U37113 ( .A(n36844), .B(n36843), .Z(n36845) );
  XNOR U37114 ( .A(n36846), .B(n36845), .Z(n36819) );
  XOR U37115 ( .A(n36820), .B(n36819), .Z(n36822) );
  XOR U37116 ( .A(n36821), .B(n36822), .Z(n36814) );
  NANDN U37117 ( .A(n36742), .B(n36741), .Z(n36744) );
  XOR U37118 ( .A(a[126]), .B(b[43]), .Z(n36892) );
  NANDN U37119 ( .A(n36891), .B(n36892), .Z(n36743) );
  AND U37120 ( .A(n36744), .B(n36743), .Z(n36860) );
  NANDN U37121 ( .A(n38247), .B(n36745), .Z(n36747) );
  XOR U37122 ( .A(b[61]), .B(a[108]), .Z(n36879) );
  NANDN U37123 ( .A(n38248), .B(n36879), .Z(n36746) );
  AND U37124 ( .A(n36747), .B(n36746), .Z(n36859) );
  NANDN U37125 ( .A(n37705), .B(n36748), .Z(n36750) );
  XOR U37126 ( .A(b[53]), .B(a[116]), .Z(n36867) );
  NANDN U37127 ( .A(n37778), .B(n36867), .Z(n36749) );
  NAND U37128 ( .A(n36750), .B(n36749), .Z(n36858) );
  XOR U37129 ( .A(n36859), .B(n36858), .Z(n36861) );
  XOR U37130 ( .A(n36860), .B(n36861), .Z(n36826) );
  NANDN U37131 ( .A(n36752), .B(n36751), .Z(n36756) );
  NAND U37132 ( .A(n36754), .B(n36753), .Z(n36755) );
  AND U37133 ( .A(n36756), .B(n36755), .Z(n36825) );
  XNOR U37134 ( .A(n36826), .B(n36825), .Z(n36827) );
  NANDN U37135 ( .A(n36758), .B(n36757), .Z(n36762) );
  OR U37136 ( .A(n36760), .B(n36759), .Z(n36761) );
  NAND U37137 ( .A(n36762), .B(n36761), .Z(n36828) );
  XNOR U37138 ( .A(n36827), .B(n36828), .Z(n36813) );
  XOR U37139 ( .A(n36814), .B(n36813), .Z(n36816) );
  XOR U37140 ( .A(n36815), .B(n36816), .Z(n36809) );
  NANDN U37141 ( .A(n36764), .B(n36763), .Z(n36768) );
  NAND U37142 ( .A(n36766), .B(n36765), .Z(n36767) );
  AND U37143 ( .A(n36768), .B(n36767), .Z(n36840) );
  NANDN U37144 ( .A(n36770), .B(n36769), .Z(n36774) );
  NANDN U37145 ( .A(n36772), .B(n36771), .Z(n36773) );
  AND U37146 ( .A(n36774), .B(n36773), .Z(n36838) );
  NANDN U37147 ( .A(n36776), .B(n36775), .Z(n36780) );
  NANDN U37148 ( .A(n36778), .B(n36777), .Z(n36779) );
  AND U37149 ( .A(n36780), .B(n36779), .Z(n36837) );
  XNOR U37150 ( .A(n36838), .B(n36837), .Z(n36839) );
  XOR U37151 ( .A(n36840), .B(n36839), .Z(n36808) );
  NANDN U37152 ( .A(n36782), .B(n36781), .Z(n36786) );
  OR U37153 ( .A(n36784), .B(n36783), .Z(n36785) );
  NAND U37154 ( .A(n36786), .B(n36785), .Z(n36807) );
  XOR U37155 ( .A(n36808), .B(n36807), .Z(n36810) );
  XOR U37156 ( .A(n36809), .B(n36810), .Z(n36802) );
  NANDN U37157 ( .A(n36788), .B(n36787), .Z(n36792) );
  NANDN U37158 ( .A(n36790), .B(n36789), .Z(n36791) );
  NAND U37159 ( .A(n36792), .B(n36791), .Z(n36801) );
  XNOR U37160 ( .A(n36802), .B(n36801), .Z(n36803) );
  XNOR U37161 ( .A(n36804), .B(n36803), .Z(n36795) );
  XOR U37162 ( .A(n36796), .B(n36795), .Z(n36798) );
  XNOR U37163 ( .A(n36797), .B(n36798), .Z(n36793) );
  XOR U37164 ( .A(n36794), .B(n36793), .Z(c[232]) );
  AND U37165 ( .A(n36794), .B(n36793), .Z(n36905) );
  NANDN U37166 ( .A(n36796), .B(n36795), .Z(n36800) );
  OR U37167 ( .A(n36798), .B(n36797), .Z(n36799) );
  AND U37168 ( .A(n36800), .B(n36799), .Z(n36908) );
  NANDN U37169 ( .A(n36802), .B(n36801), .Z(n36806) );
  NANDN U37170 ( .A(n36804), .B(n36803), .Z(n36805) );
  AND U37171 ( .A(n36806), .B(n36805), .Z(n36907) );
  NANDN U37172 ( .A(n36808), .B(n36807), .Z(n36812) );
  OR U37173 ( .A(n36810), .B(n36809), .Z(n36811) );
  AND U37174 ( .A(n36812), .B(n36811), .Z(n36914) );
  NANDN U37175 ( .A(n36814), .B(n36813), .Z(n36818) );
  OR U37176 ( .A(n36816), .B(n36815), .Z(n36817) );
  AND U37177 ( .A(n36818), .B(n36817), .Z(n36913) );
  NANDN U37178 ( .A(n36820), .B(n36819), .Z(n36824) );
  OR U37179 ( .A(n36822), .B(n36821), .Z(n36823) );
  AND U37180 ( .A(n36824), .B(n36823), .Z(n37014) );
  NANDN U37181 ( .A(n36826), .B(n36825), .Z(n36830) );
  NANDN U37182 ( .A(n36828), .B(n36827), .Z(n36829) );
  AND U37183 ( .A(n36830), .B(n36829), .Z(n37013) );
  NANDN U37184 ( .A(n36832), .B(n36831), .Z(n36836) );
  OR U37185 ( .A(n36834), .B(n36833), .Z(n36835) );
  NAND U37186 ( .A(n36836), .B(n36835), .Z(n37012) );
  XOR U37187 ( .A(n37013), .B(n37012), .Z(n37015) );
  XNOR U37188 ( .A(n37014), .B(n37015), .Z(n36920) );
  NANDN U37189 ( .A(n36838), .B(n36837), .Z(n36842) );
  NAND U37190 ( .A(n36840), .B(n36839), .Z(n36841) );
  AND U37191 ( .A(n36842), .B(n36841), .Z(n36919) );
  NANDN U37192 ( .A(n36844), .B(n36843), .Z(n36848) );
  NANDN U37193 ( .A(n36846), .B(n36845), .Z(n36847) );
  AND U37194 ( .A(n36848), .B(n36847), .Z(n36926) );
  NANDN U37195 ( .A(n36850), .B(n36849), .Z(n36854) );
  OR U37196 ( .A(n36852), .B(n36851), .Z(n36853) );
  AND U37197 ( .A(n36854), .B(n36853), .Z(n37007) );
  XNOR U37198 ( .A(n37007), .B(n37006), .Z(n37009) );
  NANDN U37199 ( .A(n36859), .B(n36858), .Z(n36863) );
  OR U37200 ( .A(n36861), .B(n36860), .Z(n36862) );
  AND U37201 ( .A(n36863), .B(n36862), .Z(n37003) );
  NANDN U37202 ( .A(n38278), .B(n36864), .Z(n36866) );
  XOR U37203 ( .A(b[63]), .B(a[107]), .Z(n36958) );
  NANDN U37204 ( .A(n38279), .B(n36958), .Z(n36865) );
  AND U37205 ( .A(n36866), .B(n36865), .Z(n36955) );
  NANDN U37206 ( .A(n37705), .B(n36867), .Z(n36869) );
  XOR U37207 ( .A(b[53]), .B(a[117]), .Z(n36969) );
  NANDN U37208 ( .A(n37778), .B(n36969), .Z(n36868) );
  NAND U37209 ( .A(n36869), .B(n36868), .Z(n36954) );
  XNOR U37210 ( .A(n36955), .B(n36954), .Z(n36957) );
  XOR U37211 ( .A(n36942), .B(n36943), .Z(n36945) );
  AND U37212 ( .A(b[63]), .B(a[105]), .Z(n36944) );
  XOR U37213 ( .A(n36945), .B(n36944), .Z(n36956) );
  XOR U37214 ( .A(n36957), .B(n36956), .Z(n37000) );
  NANDN U37215 ( .A(n37974), .B(n36870), .Z(n36872) );
  XOR U37216 ( .A(b[57]), .B(a[113]), .Z(n36966) );
  NANDN U37217 ( .A(n38031), .B(n36966), .Z(n36871) );
  AND U37218 ( .A(n36872), .B(n36871), .Z(n36997) );
  NANDN U37219 ( .A(n38090), .B(n36873), .Z(n36875) );
  XOR U37220 ( .A(b[59]), .B(a[111]), .Z(n36981) );
  NANDN U37221 ( .A(n38130), .B(n36981), .Z(n36874) );
  AND U37222 ( .A(n36875), .B(n36874), .Z(n36995) );
  NANDN U37223 ( .A(n37526), .B(n36876), .Z(n36878) );
  XOR U37224 ( .A(a[119]), .B(b[51]), .Z(n36972) );
  NANDN U37225 ( .A(n37605), .B(n36972), .Z(n36877) );
  NAND U37226 ( .A(n36878), .B(n36877), .Z(n36994) );
  XNOR U37227 ( .A(n36995), .B(n36994), .Z(n36996) );
  XOR U37228 ( .A(n36997), .B(n36996), .Z(n37001) );
  XNOR U37229 ( .A(n37000), .B(n37001), .Z(n37002) );
  XNOR U37230 ( .A(n37003), .B(n37002), .Z(n37008) );
  XOR U37231 ( .A(n37009), .B(n37008), .Z(n36925) );
  NANDN U37232 ( .A(n38247), .B(n36879), .Z(n36881) );
  XOR U37233 ( .A(b[61]), .B(a[109]), .Z(n36975) );
  NANDN U37234 ( .A(n38248), .B(n36975), .Z(n36880) );
  AND U37235 ( .A(n36881), .B(n36880), .Z(n36938) );
  NANDN U37236 ( .A(n36882), .B(n37536), .Z(n36884) );
  XOR U37237 ( .A(a[121]), .B(b[49]), .Z(n36978) );
  NANDN U37238 ( .A(n37432), .B(n36978), .Z(n36883) );
  AND U37239 ( .A(n36884), .B(n36883), .Z(n36937) );
  NANDN U37240 ( .A(n211), .B(n36885), .Z(n36887) );
  XOR U37241 ( .A(a[123]), .B(b[47]), .Z(n36987) );
  NANDN U37242 ( .A(n37172), .B(n36987), .Z(n36886) );
  NAND U37243 ( .A(n36887), .B(n36886), .Z(n36936) );
  XOR U37244 ( .A(n36937), .B(n36936), .Z(n36939) );
  XOR U37245 ( .A(n36938), .B(n36939), .Z(n36931) );
  NANDN U37246 ( .A(n36991), .B(n36888), .Z(n36890) );
  XOR U37247 ( .A(a[125]), .B(b[45]), .Z(n36990) );
  NANDN U37248 ( .A(n37083), .B(n36990), .Z(n36889) );
  AND U37249 ( .A(n36890), .B(n36889), .Z(n36950) );
  XNOR U37250 ( .A(a[127]), .B(b[43]), .Z(n36961) );
  OR U37251 ( .A(n36961), .B(n36891), .Z(n36894) );
  NAND U37252 ( .A(n36962), .B(n36892), .Z(n36893) );
  AND U37253 ( .A(n36894), .B(n36893), .Z(n36949) );
  NANDN U37254 ( .A(n37857), .B(n36895), .Z(n36897) );
  XOR U37255 ( .A(b[55]), .B(a[115]), .Z(n36984) );
  NANDN U37256 ( .A(n37911), .B(n36984), .Z(n36896) );
  NAND U37257 ( .A(n36897), .B(n36896), .Z(n36948) );
  XOR U37258 ( .A(n36949), .B(n36948), .Z(n36951) );
  XNOR U37259 ( .A(n36950), .B(n36951), .Z(n36930) );
  XNOR U37260 ( .A(n36931), .B(n36930), .Z(n36932) );
  NANDN U37261 ( .A(n36899), .B(n36898), .Z(n36903) );
  OR U37262 ( .A(n36901), .B(n36900), .Z(n36902) );
  NAND U37263 ( .A(n36903), .B(n36902), .Z(n36933) );
  XNOR U37264 ( .A(n36932), .B(n36933), .Z(n36924) );
  XOR U37265 ( .A(n36925), .B(n36924), .Z(n36927) );
  XNOR U37266 ( .A(n36926), .B(n36927), .Z(n36918) );
  XOR U37267 ( .A(n36919), .B(n36918), .Z(n36921) );
  XNOR U37268 ( .A(n36920), .B(n36921), .Z(n36912) );
  XOR U37269 ( .A(n36913), .B(n36912), .Z(n36915) );
  XNOR U37270 ( .A(n36914), .B(n36915), .Z(n36906) );
  XOR U37271 ( .A(n36907), .B(n36906), .Z(n36909) );
  XNOR U37272 ( .A(n36908), .B(n36909), .Z(n36904) );
  XOR U37273 ( .A(n36905), .B(n36904), .Z(c[233]) );
  AND U37274 ( .A(n36905), .B(n36904), .Z(n37019) );
  NANDN U37275 ( .A(n36907), .B(n36906), .Z(n36911) );
  OR U37276 ( .A(n36909), .B(n36908), .Z(n36910) );
  AND U37277 ( .A(n36911), .B(n36910), .Z(n37022) );
  NANDN U37278 ( .A(n36913), .B(n36912), .Z(n36917) );
  NANDN U37279 ( .A(n36915), .B(n36914), .Z(n36916) );
  AND U37280 ( .A(n36917), .B(n36916), .Z(n37021) );
  NANDN U37281 ( .A(n36919), .B(n36918), .Z(n36923) );
  NANDN U37282 ( .A(n36921), .B(n36920), .Z(n36922) );
  AND U37283 ( .A(n36923), .B(n36922), .Z(n37118) );
  NANDN U37284 ( .A(n36925), .B(n36924), .Z(n36929) );
  NANDN U37285 ( .A(n36927), .B(n36926), .Z(n36928) );
  AND U37286 ( .A(n36929), .B(n36928), .Z(n37111) );
  NANDN U37287 ( .A(n36931), .B(n36930), .Z(n36935) );
  NANDN U37288 ( .A(n36933), .B(n36932), .Z(n36934) );
  AND U37289 ( .A(n36935), .B(n36934), .Z(n37027) );
  NANDN U37290 ( .A(n36937), .B(n36936), .Z(n36941) );
  OR U37291 ( .A(n36939), .B(n36938), .Z(n36940) );
  AND U37292 ( .A(n36941), .B(n36940), .Z(n37105) );
  OR U37293 ( .A(n36943), .B(n36942), .Z(n36947) );
  NAND U37294 ( .A(n36945), .B(n36944), .Z(n36946) );
  AND U37295 ( .A(n36947), .B(n36946), .Z(n37103) );
  NANDN U37296 ( .A(n36949), .B(n36948), .Z(n36953) );
  OR U37297 ( .A(n36951), .B(n36950), .Z(n36952) );
  NAND U37298 ( .A(n36953), .B(n36952), .Z(n37104) );
  XOR U37299 ( .A(n37103), .B(n37104), .Z(n37106) );
  XNOR U37300 ( .A(n37105), .B(n37106), .Z(n37026) );
  XNOR U37301 ( .A(n37027), .B(n37026), .Z(n37028) );
  NANDN U37302 ( .A(n38278), .B(n36958), .Z(n36960) );
  XOR U37303 ( .A(b[63]), .B(a[108]), .Z(n37091) );
  NANDN U37304 ( .A(n38279), .B(n37091), .Z(n36959) );
  AND U37305 ( .A(n36960), .B(n36959), .Z(n37079) );
  NAND U37306 ( .A(b[63]), .B(a[106]), .Z(n37179) );
  ANDN U37307 ( .B(n36962), .A(n36961), .Z(n36965) );
  NAND U37308 ( .A(b[43]), .B(n36963), .Z(n36964) );
  NANDN U37309 ( .A(n36965), .B(n36964), .Z(n37077) );
  XOR U37310 ( .A(n37179), .B(n37077), .Z(n37078) );
  XNOR U37311 ( .A(n37079), .B(n37078), .Z(n37038) );
  NANDN U37312 ( .A(n37974), .B(n36966), .Z(n36968) );
  XOR U37313 ( .A(b[57]), .B(a[114]), .Z(n37068) );
  NANDN U37314 ( .A(n38031), .B(n37068), .Z(n36967) );
  AND U37315 ( .A(n36968), .B(n36967), .Z(n37053) );
  NANDN U37316 ( .A(n37705), .B(n36969), .Z(n36971) );
  XOR U37317 ( .A(b[53]), .B(a[118]), .Z(n37087) );
  NANDN U37318 ( .A(n37778), .B(n37087), .Z(n36970) );
  AND U37319 ( .A(n36971), .B(n36970), .Z(n37051) );
  NANDN U37320 ( .A(n37526), .B(n36972), .Z(n36974) );
  XOR U37321 ( .A(a[120]), .B(b[51]), .Z(n37074) );
  NANDN U37322 ( .A(n37605), .B(n37074), .Z(n36973) );
  NAND U37323 ( .A(n36974), .B(n36973), .Z(n37050) );
  XNOR U37324 ( .A(n37051), .B(n37050), .Z(n37052) );
  XOR U37325 ( .A(n37053), .B(n37052), .Z(n37039) );
  XOR U37326 ( .A(n37038), .B(n37039), .Z(n37041) );
  XOR U37327 ( .A(n37040), .B(n37041), .Z(n37098) );
  NANDN U37328 ( .A(n38247), .B(n36975), .Z(n36977) );
  XOR U37329 ( .A(b[61]), .B(a[110]), .Z(n37080) );
  NANDN U37330 ( .A(n38248), .B(n37080), .Z(n36976) );
  AND U37331 ( .A(n36977), .B(n36976), .Z(n37046) );
  NANDN U37332 ( .A(n212), .B(n36978), .Z(n36980) );
  XOR U37333 ( .A(a[122]), .B(b[49]), .Z(n37062) );
  NANDN U37334 ( .A(n37432), .B(n37062), .Z(n36979) );
  AND U37335 ( .A(n36980), .B(n36979), .Z(n37045) );
  NANDN U37336 ( .A(n38090), .B(n36981), .Z(n36983) );
  XOR U37337 ( .A(b[59]), .B(a[112]), .Z(n37071) );
  NANDN U37338 ( .A(n38130), .B(n37071), .Z(n36982) );
  NAND U37339 ( .A(n36983), .B(n36982), .Z(n37044) );
  XOR U37340 ( .A(n37045), .B(n37044), .Z(n37047) );
  XOR U37341 ( .A(n37046), .B(n37047), .Z(n37033) );
  NANDN U37342 ( .A(n37857), .B(n36984), .Z(n36986) );
  XOR U37343 ( .A(b[55]), .B(a[116]), .Z(n37094) );
  NANDN U37344 ( .A(n37911), .B(n37094), .Z(n36985) );
  AND U37345 ( .A(n36986), .B(n36985), .Z(n37058) );
  NANDN U37346 ( .A(n211), .B(n36987), .Z(n36989) );
  XOR U37347 ( .A(a[124]), .B(b[47]), .Z(n37065) );
  NANDN U37348 ( .A(n37172), .B(n37065), .Z(n36988) );
  AND U37349 ( .A(n36989), .B(n36988), .Z(n37057) );
  NANDN U37350 ( .A(n36991), .B(n36990), .Z(n36993) );
  XOR U37351 ( .A(a[126]), .B(b[45]), .Z(n37084) );
  NANDN U37352 ( .A(n37083), .B(n37084), .Z(n36992) );
  NAND U37353 ( .A(n36993), .B(n36992), .Z(n37056) );
  XOR U37354 ( .A(n37057), .B(n37056), .Z(n37059) );
  XNOR U37355 ( .A(n37058), .B(n37059), .Z(n37032) );
  XNOR U37356 ( .A(n37033), .B(n37032), .Z(n37034) );
  NANDN U37357 ( .A(n36995), .B(n36994), .Z(n36999) );
  NANDN U37358 ( .A(n36997), .B(n36996), .Z(n36998) );
  NAND U37359 ( .A(n36999), .B(n36998), .Z(n37035) );
  XNOR U37360 ( .A(n37034), .B(n37035), .Z(n37097) );
  XNOR U37361 ( .A(n37098), .B(n37097), .Z(n37099) );
  NANDN U37362 ( .A(n37001), .B(n37000), .Z(n37005) );
  NANDN U37363 ( .A(n37003), .B(n37002), .Z(n37004) );
  NAND U37364 ( .A(n37005), .B(n37004), .Z(n37100) );
  XOR U37365 ( .A(n37099), .B(n37100), .Z(n37029) );
  XNOR U37366 ( .A(n37028), .B(n37029), .Z(n37109) );
  NANDN U37367 ( .A(n37007), .B(n37006), .Z(n37011) );
  NAND U37368 ( .A(n37009), .B(n37008), .Z(n37010) );
  NAND U37369 ( .A(n37011), .B(n37010), .Z(n37110) );
  XOR U37370 ( .A(n37109), .B(n37110), .Z(n37112) );
  XOR U37371 ( .A(n37111), .B(n37112), .Z(n37116) );
  NANDN U37372 ( .A(n37013), .B(n37012), .Z(n37017) );
  NANDN U37373 ( .A(n37015), .B(n37014), .Z(n37016) );
  AND U37374 ( .A(n37017), .B(n37016), .Z(n37115) );
  XNOR U37375 ( .A(n37116), .B(n37115), .Z(n37117) );
  XNOR U37376 ( .A(n37118), .B(n37117), .Z(n37020) );
  XOR U37377 ( .A(n37021), .B(n37020), .Z(n37023) );
  XNOR U37378 ( .A(n37022), .B(n37023), .Z(n37018) );
  XOR U37379 ( .A(n37019), .B(n37018), .Z(c[234]) );
  AND U37380 ( .A(n37019), .B(n37018), .Z(n37122) );
  NANDN U37381 ( .A(n37021), .B(n37020), .Z(n37025) );
  OR U37382 ( .A(n37023), .B(n37022), .Z(n37024) );
  AND U37383 ( .A(n37025), .B(n37024), .Z(n37125) );
  NANDN U37384 ( .A(n37027), .B(n37026), .Z(n37031) );
  NANDN U37385 ( .A(n37029), .B(n37028), .Z(n37030) );
  AND U37386 ( .A(n37031), .B(n37030), .Z(n37129) );
  NANDN U37387 ( .A(n37033), .B(n37032), .Z(n37037) );
  NANDN U37388 ( .A(n37035), .B(n37034), .Z(n37036) );
  AND U37389 ( .A(n37037), .B(n37036), .Z(n37142) );
  NANDN U37390 ( .A(n37039), .B(n37038), .Z(n37043) );
  OR U37391 ( .A(n37041), .B(n37040), .Z(n37042) );
  AND U37392 ( .A(n37043), .B(n37042), .Z(n37141) );
  XNOR U37393 ( .A(n37142), .B(n37141), .Z(n37144) );
  NANDN U37394 ( .A(n37045), .B(n37044), .Z(n37049) );
  OR U37395 ( .A(n37047), .B(n37046), .Z(n37048) );
  AND U37396 ( .A(n37049), .B(n37048), .Z(n37217) );
  NANDN U37397 ( .A(n37051), .B(n37050), .Z(n37055) );
  NANDN U37398 ( .A(n37053), .B(n37052), .Z(n37054) );
  AND U37399 ( .A(n37055), .B(n37054), .Z(n37215) );
  NANDN U37400 ( .A(n37057), .B(n37056), .Z(n37061) );
  OR U37401 ( .A(n37059), .B(n37058), .Z(n37060) );
  AND U37402 ( .A(n37061), .B(n37060), .Z(n37219) );
  NANDN U37403 ( .A(n212), .B(n37062), .Z(n37064) );
  XOR U37404 ( .A(a[123]), .B(b[49]), .Z(n37168) );
  NANDN U37405 ( .A(n37432), .B(n37168), .Z(n37063) );
  AND U37406 ( .A(n37064), .B(n37063), .Z(n37150) );
  NANDN U37407 ( .A(n211), .B(n37065), .Z(n37067) );
  XOR U37408 ( .A(a[125]), .B(b[47]), .Z(n37171) );
  NANDN U37409 ( .A(n37172), .B(n37171), .Z(n37066) );
  AND U37410 ( .A(n37067), .B(n37066), .Z(n37148) );
  NAND U37411 ( .A(n38076), .B(n37068), .Z(n37070) );
  XNOR U37412 ( .A(b[57]), .B(a[115]), .Z(n37175) );
  NANDN U37413 ( .A(n37175), .B(n38077), .Z(n37069) );
  NAND U37414 ( .A(n37070), .B(n37069), .Z(n37210) );
  NAND U37415 ( .A(n38174), .B(n37071), .Z(n37073) );
  XNOR U37416 ( .A(b[59]), .B(a[113]), .Z(n37159) );
  NANDN U37417 ( .A(n37159), .B(n38175), .Z(n37072) );
  NAND U37418 ( .A(n37073), .B(n37072), .Z(n37209) );
  NANDN U37419 ( .A(n37526), .B(n37074), .Z(n37076) );
  XOR U37420 ( .A(a[121]), .B(b[51]), .Z(n37153) );
  NANDN U37421 ( .A(n37605), .B(n37153), .Z(n37075) );
  NAND U37422 ( .A(n37076), .B(n37075), .Z(n37208) );
  XOR U37423 ( .A(n37209), .B(n37208), .Z(n37211) );
  XOR U37424 ( .A(n37210), .B(n37211), .Z(n37147) );
  XNOR U37425 ( .A(n37148), .B(n37147), .Z(n37149) );
  XOR U37426 ( .A(n37150), .B(n37149), .Z(n37218) );
  XOR U37427 ( .A(n37219), .B(n37218), .Z(n37221) );
  NANDN U37428 ( .A(n38247), .B(n37080), .Z(n37082) );
  XOR U37429 ( .A(b[61]), .B(a[111]), .Z(n37162) );
  NANDN U37430 ( .A(n38248), .B(n37162), .Z(n37081) );
  AND U37431 ( .A(n37082), .B(n37081), .Z(n37186) );
  XNOR U37432 ( .A(a[127]), .B(b[45]), .Z(n37201) );
  OR U37433 ( .A(n37201), .B(n37083), .Z(n37086) );
  NAND U37434 ( .A(n37202), .B(n37084), .Z(n37085) );
  AND U37435 ( .A(n37086), .B(n37085), .Z(n37185) );
  NANDN U37436 ( .A(n37705), .B(n37087), .Z(n37089) );
  XOR U37437 ( .A(b[53]), .B(a[119]), .Z(n37156) );
  NANDN U37438 ( .A(n37778), .B(n37156), .Z(n37088) );
  NAND U37439 ( .A(n37089), .B(n37088), .Z(n37184) );
  XOR U37440 ( .A(n37185), .B(n37184), .Z(n37187) );
  XOR U37441 ( .A(n37186), .B(n37187), .Z(n37191) );
  AND U37442 ( .A(b[63]), .B(a[107]), .Z(n37181) );
  XOR U37443 ( .A(n37090), .B(n37181), .Z(n37178) );
  XOR U37444 ( .A(n37179), .B(n37178), .Z(n37196) );
  NAND U37445 ( .A(n38262), .B(n37091), .Z(n37093) );
  XNOR U37446 ( .A(b[63]), .B(a[109]), .Z(n37205) );
  NANDN U37447 ( .A(n37205), .B(n38264), .Z(n37092) );
  AND U37448 ( .A(n37093), .B(n37092), .Z(n37197) );
  XOR U37449 ( .A(n37196), .B(n37197), .Z(n37198) );
  NAND U37450 ( .A(n37984), .B(n37094), .Z(n37096) );
  XNOR U37451 ( .A(b[55]), .B(a[117]), .Z(n37165) );
  NANDN U37452 ( .A(n37165), .B(n37985), .Z(n37095) );
  NAND U37453 ( .A(n37096), .B(n37095), .Z(n37199) );
  XNOR U37454 ( .A(n37198), .B(n37199), .Z(n37190) );
  XNOR U37455 ( .A(n37191), .B(n37190), .Z(n37192) );
  XOR U37456 ( .A(n37193), .B(n37192), .Z(n37220) );
  XOR U37457 ( .A(n37221), .B(n37220), .Z(n37214) );
  XOR U37458 ( .A(n37215), .B(n37214), .Z(n37216) );
  XOR U37459 ( .A(n37217), .B(n37216), .Z(n37143) );
  XOR U37460 ( .A(n37144), .B(n37143), .Z(n37138) );
  NANDN U37461 ( .A(n37098), .B(n37097), .Z(n37102) );
  NANDN U37462 ( .A(n37100), .B(n37099), .Z(n37101) );
  AND U37463 ( .A(n37102), .B(n37101), .Z(n37135) );
  NANDN U37464 ( .A(n37104), .B(n37103), .Z(n37108) );
  NANDN U37465 ( .A(n37106), .B(n37105), .Z(n37107) );
  NAND U37466 ( .A(n37108), .B(n37107), .Z(n37136) );
  XNOR U37467 ( .A(n37135), .B(n37136), .Z(n37137) );
  XOR U37468 ( .A(n37138), .B(n37137), .Z(n37130) );
  XNOR U37469 ( .A(n37129), .B(n37130), .Z(n37132) );
  NANDN U37470 ( .A(n37110), .B(n37109), .Z(n37114) );
  OR U37471 ( .A(n37112), .B(n37111), .Z(n37113) );
  AND U37472 ( .A(n37114), .B(n37113), .Z(n37131) );
  XOR U37473 ( .A(n37132), .B(n37131), .Z(n37124) );
  NANDN U37474 ( .A(n37116), .B(n37115), .Z(n37120) );
  NAND U37475 ( .A(n37118), .B(n37117), .Z(n37119) );
  AND U37476 ( .A(n37120), .B(n37119), .Z(n37123) );
  XOR U37477 ( .A(n37124), .B(n37123), .Z(n37126) );
  XNOR U37478 ( .A(n37125), .B(n37126), .Z(n37121) );
  XOR U37479 ( .A(n37122), .B(n37121), .Z(c[235]) );
  AND U37480 ( .A(n37122), .B(n37121), .Z(n37225) );
  NANDN U37481 ( .A(n37124), .B(n37123), .Z(n37128) );
  OR U37482 ( .A(n37126), .B(n37125), .Z(n37127) );
  AND U37483 ( .A(n37128), .B(n37127), .Z(n37228) );
  NANDN U37484 ( .A(n37130), .B(n37129), .Z(n37134) );
  NAND U37485 ( .A(n37132), .B(n37131), .Z(n37133) );
  AND U37486 ( .A(n37134), .B(n37133), .Z(n37226) );
  NANDN U37487 ( .A(n37136), .B(n37135), .Z(n37140) );
  NANDN U37488 ( .A(n37138), .B(n37137), .Z(n37139) );
  AND U37489 ( .A(n37140), .B(n37139), .Z(n37234) );
  NANDN U37490 ( .A(n37142), .B(n37141), .Z(n37146) );
  NAND U37491 ( .A(n37144), .B(n37143), .Z(n37145) );
  AND U37492 ( .A(n37146), .B(n37145), .Z(n37233) );
  NANDN U37493 ( .A(n37148), .B(n37147), .Z(n37152) );
  NANDN U37494 ( .A(n37150), .B(n37149), .Z(n37151) );
  AND U37495 ( .A(n37152), .B(n37151), .Z(n37246) );
  NANDN U37496 ( .A(n37526), .B(n37153), .Z(n37155) );
  XOR U37497 ( .A(a[122]), .B(b[51]), .Z(n37269) );
  NANDN U37498 ( .A(n37605), .B(n37269), .Z(n37154) );
  AND U37499 ( .A(n37155), .B(n37154), .Z(n37283) );
  NANDN U37500 ( .A(n37705), .B(n37156), .Z(n37158) );
  XOR U37501 ( .A(a[120]), .B(b[53]), .Z(n37272) );
  NANDN U37502 ( .A(n37778), .B(n37272), .Z(n37157) );
  AND U37503 ( .A(n37158), .B(n37157), .Z(n37282) );
  NANDN U37504 ( .A(n37159), .B(n38174), .Z(n37161) );
  XOR U37505 ( .A(b[59]), .B(a[114]), .Z(n37263) );
  NANDN U37506 ( .A(n38130), .B(n37263), .Z(n37160) );
  AND U37507 ( .A(n37161), .B(n37160), .Z(n37290) );
  NANDN U37508 ( .A(n38247), .B(n37162), .Z(n37164) );
  XOR U37509 ( .A(b[61]), .B(a[112]), .Z(n37266) );
  NANDN U37510 ( .A(n38248), .B(n37266), .Z(n37163) );
  AND U37511 ( .A(n37164), .B(n37163), .Z(n37288) );
  NANDN U37512 ( .A(n37165), .B(n37984), .Z(n37167) );
  XOR U37513 ( .A(b[55]), .B(a[118]), .Z(n37260) );
  NANDN U37514 ( .A(n37911), .B(n37260), .Z(n37166) );
  NAND U37515 ( .A(n37167), .B(n37166), .Z(n37287) );
  XNOR U37516 ( .A(n37288), .B(n37287), .Z(n37289) );
  XNOR U37517 ( .A(n37290), .B(n37289), .Z(n37281) );
  XOR U37518 ( .A(n37282), .B(n37281), .Z(n37284) );
  XOR U37519 ( .A(n37283), .B(n37284), .Z(n37306) );
  NANDN U37520 ( .A(n212), .B(n37168), .Z(n37170) );
  XOR U37521 ( .A(a[124]), .B(b[49]), .Z(n37254) );
  NANDN U37522 ( .A(n37432), .B(n37254), .Z(n37169) );
  AND U37523 ( .A(n37170), .B(n37169), .Z(n37277) );
  NANDN U37524 ( .A(n211), .B(n37171), .Z(n37174) );
  XOR U37525 ( .A(a[126]), .B(b[47]), .Z(n37293) );
  NANDN U37526 ( .A(n37172), .B(n37293), .Z(n37173) );
  AND U37527 ( .A(n37174), .B(n37173), .Z(n37276) );
  NANDN U37528 ( .A(n37175), .B(n38076), .Z(n37177) );
  XOR U37529 ( .A(b[57]), .B(a[116]), .Z(n37297) );
  NANDN U37530 ( .A(n38031), .B(n37297), .Z(n37176) );
  NAND U37531 ( .A(n37177), .B(n37176), .Z(n37275) );
  XOR U37532 ( .A(n37276), .B(n37275), .Z(n37278) );
  XOR U37533 ( .A(n37277), .B(n37278), .Z(n37304) );
  NANDN U37534 ( .A(n37179), .B(n37178), .Z(n37183) );
  ANDN U37535 ( .B(n37181), .A(n37180), .Z(n37182) );
  ANDN U37536 ( .B(n37183), .A(n37182), .Z(n37303) );
  XNOR U37537 ( .A(n37304), .B(n37303), .Z(n37305) );
  XNOR U37538 ( .A(n37306), .B(n37305), .Z(n37244) );
  NANDN U37539 ( .A(n37185), .B(n37184), .Z(n37189) );
  OR U37540 ( .A(n37187), .B(n37186), .Z(n37188) );
  NAND U37541 ( .A(n37189), .B(n37188), .Z(n37245) );
  XOR U37542 ( .A(n37244), .B(n37245), .Z(n37247) );
  XNOR U37543 ( .A(n37246), .B(n37247), .Z(n37240) );
  NANDN U37544 ( .A(n37191), .B(n37190), .Z(n37195) );
  NAND U37545 ( .A(n37193), .B(n37192), .Z(n37194) );
  AND U37546 ( .A(n37195), .B(n37194), .Z(n37239) );
  NAND U37547 ( .A(b[45]), .B(n37200), .Z(n37204) );
  ANDN U37548 ( .B(n37202), .A(n37201), .Z(n37203) );
  ANDN U37549 ( .B(n37204), .A(n37203), .Z(n37302) );
  NAND U37550 ( .A(b[63]), .B(a[108]), .Z(n37337) );
  NANDN U37551 ( .A(n37205), .B(n38262), .Z(n37207) );
  XOR U37552 ( .A(b[63]), .B(a[110]), .Z(n37257) );
  NANDN U37553 ( .A(n38279), .B(n37257), .Z(n37206) );
  NAND U37554 ( .A(n37207), .B(n37206), .Z(n37300) );
  XOR U37555 ( .A(n37337), .B(n37300), .Z(n37301) );
  XOR U37556 ( .A(n37302), .B(n37301), .Z(n37250) );
  NAND U37557 ( .A(n37209), .B(n37208), .Z(n37213) );
  NAND U37558 ( .A(n37211), .B(n37210), .Z(n37212) );
  AND U37559 ( .A(n37213), .B(n37212), .Z(n37251) );
  XOR U37560 ( .A(n37250), .B(n37251), .Z(n37252) );
  XNOR U37561 ( .A(n37253), .B(n37252), .Z(n37238) );
  XOR U37562 ( .A(n37239), .B(n37238), .Z(n37241) );
  XNOR U37563 ( .A(n37240), .B(n37241), .Z(n37311) );
  NAND U37564 ( .A(n37219), .B(n37218), .Z(n37223) );
  NAND U37565 ( .A(n37221), .B(n37220), .Z(n37222) );
  NAND U37566 ( .A(n37223), .B(n37222), .Z(n37309) );
  XOR U37567 ( .A(n37310), .B(n37309), .Z(n37312) );
  XNOR U37568 ( .A(n37311), .B(n37312), .Z(n37232) );
  XOR U37569 ( .A(n37233), .B(n37232), .Z(n37235) );
  XOR U37570 ( .A(n37234), .B(n37235), .Z(n37227) );
  XOR U37571 ( .A(n37226), .B(n37227), .Z(n37229) );
  XNOR U37572 ( .A(n37228), .B(n37229), .Z(n37224) );
  XOR U37573 ( .A(n37225), .B(n37224), .Z(c[236]) );
  AND U37574 ( .A(n37225), .B(n37224), .Z(n37316) );
  NANDN U37575 ( .A(n37227), .B(n37226), .Z(n37231) );
  OR U37576 ( .A(n37229), .B(n37228), .Z(n37230) );
  AND U37577 ( .A(n37231), .B(n37230), .Z(n37319) );
  NANDN U37578 ( .A(n37233), .B(n37232), .Z(n37237) );
  NANDN U37579 ( .A(n37235), .B(n37234), .Z(n37236) );
  AND U37580 ( .A(n37237), .B(n37236), .Z(n37318) );
  NANDN U37581 ( .A(n37239), .B(n37238), .Z(n37243) );
  NANDN U37582 ( .A(n37241), .B(n37240), .Z(n37242) );
  AND U37583 ( .A(n37243), .B(n37242), .Z(n37403) );
  NANDN U37584 ( .A(n37245), .B(n37244), .Z(n37249) );
  NANDN U37585 ( .A(n37247), .B(n37246), .Z(n37248) );
  AND U37586 ( .A(n37249), .B(n37248), .Z(n37323) );
  XNOR U37587 ( .A(n37323), .B(n37324), .Z(n37325) );
  NANDN U37588 ( .A(n212), .B(n37254), .Z(n37256) );
  XOR U37589 ( .A(a[125]), .B(b[49]), .Z(n37367) );
  NANDN U37590 ( .A(n37432), .B(n37367), .Z(n37255) );
  AND U37591 ( .A(n37256), .B(n37255), .Z(n37381) );
  NANDN U37592 ( .A(n38278), .B(n37257), .Z(n37259) );
  XOR U37593 ( .A(b[63]), .B(a[111]), .Z(n37345) );
  NANDN U37594 ( .A(n38279), .B(n37345), .Z(n37258) );
  AND U37595 ( .A(n37259), .B(n37258), .Z(n37380) );
  NANDN U37596 ( .A(n37857), .B(n37260), .Z(n37262) );
  XOR U37597 ( .A(b[55]), .B(a[119]), .Z(n37364) );
  NANDN U37598 ( .A(n37911), .B(n37364), .Z(n37261) );
  NAND U37599 ( .A(n37262), .B(n37261), .Z(n37379) );
  XOR U37600 ( .A(n37380), .B(n37379), .Z(n37382) );
  XOR U37601 ( .A(n37381), .B(n37382), .Z(n37332) );
  NANDN U37602 ( .A(n38090), .B(n37263), .Z(n37265) );
  XOR U37603 ( .A(b[59]), .B(a[115]), .Z(n37352) );
  NANDN U37604 ( .A(n38130), .B(n37352), .Z(n37264) );
  AND U37605 ( .A(n37265), .B(n37264), .Z(n37375) );
  NANDN U37606 ( .A(n38247), .B(n37266), .Z(n37268) );
  XOR U37607 ( .A(b[61]), .B(a[113]), .Z(n37355) );
  NANDN U37608 ( .A(n38248), .B(n37355), .Z(n37267) );
  AND U37609 ( .A(n37268), .B(n37267), .Z(n37374) );
  NANDN U37610 ( .A(n37526), .B(n37269), .Z(n37271) );
  XOR U37611 ( .A(a[123]), .B(b[51]), .Z(n37370) );
  NANDN U37612 ( .A(n37605), .B(n37370), .Z(n37270) );
  NAND U37613 ( .A(n37271), .B(n37270), .Z(n37373) );
  XOR U37614 ( .A(n37374), .B(n37373), .Z(n37376) );
  XOR U37615 ( .A(n37375), .B(n37376), .Z(n37330) );
  NAND U37616 ( .A(n37849), .B(n37272), .Z(n37274) );
  XNOR U37617 ( .A(a[121]), .B(b[53]), .Z(n37361) );
  NANDN U37618 ( .A(n37361), .B(n37850), .Z(n37273) );
  AND U37619 ( .A(n37274), .B(n37273), .Z(n37329) );
  XNOR U37620 ( .A(n37330), .B(n37329), .Z(n37331) );
  XNOR U37621 ( .A(n37332), .B(n37331), .Z(n37391) );
  NANDN U37622 ( .A(n37276), .B(n37275), .Z(n37280) );
  OR U37623 ( .A(n37278), .B(n37277), .Z(n37279) );
  NAND U37624 ( .A(n37280), .B(n37279), .Z(n37392) );
  XNOR U37625 ( .A(n37391), .B(n37392), .Z(n37394) );
  NANDN U37626 ( .A(n37282), .B(n37281), .Z(n37286) );
  OR U37627 ( .A(n37284), .B(n37283), .Z(n37285) );
  AND U37628 ( .A(n37286), .B(n37285), .Z(n37393) );
  XOR U37629 ( .A(n37394), .B(n37393), .Z(n37400) );
  NANDN U37630 ( .A(n37288), .B(n37287), .Z(n37292) );
  NANDN U37631 ( .A(n37290), .B(n37289), .Z(n37291) );
  AND U37632 ( .A(n37292), .B(n37291), .Z(n37385) );
  AND U37633 ( .A(b[63]), .B(a[109]), .Z(n37335) );
  XNOR U37634 ( .A(n37336), .B(n37335), .Z(n37338) );
  XOR U37635 ( .A(n37337), .B(n37338), .Z(n37348) );
  NAND U37636 ( .A(n37294), .B(n37293), .Z(n37296) );
  XOR U37637 ( .A(a[127]), .B(b[47]), .Z(n37342) );
  NAND U37638 ( .A(n37341), .B(n37342), .Z(n37295) );
  AND U37639 ( .A(n37296), .B(n37295), .Z(n37349) );
  XOR U37640 ( .A(n37348), .B(n37349), .Z(n37350) );
  NAND U37641 ( .A(n38076), .B(n37297), .Z(n37299) );
  XNOR U37642 ( .A(b[57]), .B(a[117]), .Z(n37358) );
  NANDN U37643 ( .A(n37358), .B(n38077), .Z(n37298) );
  NAND U37644 ( .A(n37299), .B(n37298), .Z(n37351) );
  XOR U37645 ( .A(n37350), .B(n37351), .Z(n37386) );
  XNOR U37646 ( .A(n37385), .B(n37386), .Z(n37388) );
  XOR U37647 ( .A(n37388), .B(n37387), .Z(n37398) );
  NANDN U37648 ( .A(n37304), .B(n37303), .Z(n37308) );
  NANDN U37649 ( .A(n37306), .B(n37305), .Z(n37307) );
  AND U37650 ( .A(n37308), .B(n37307), .Z(n37397) );
  XNOR U37651 ( .A(n37398), .B(n37397), .Z(n37399) );
  XOR U37652 ( .A(n37400), .B(n37399), .Z(n37326) );
  XOR U37653 ( .A(n37325), .B(n37326), .Z(n37404) );
  XNOR U37654 ( .A(n37403), .B(n37404), .Z(n37406) );
  NANDN U37655 ( .A(n37310), .B(n37309), .Z(n37314) );
  NANDN U37656 ( .A(n37312), .B(n37311), .Z(n37313) );
  AND U37657 ( .A(n37314), .B(n37313), .Z(n37405) );
  XNOR U37658 ( .A(n37406), .B(n37405), .Z(n37317) );
  XOR U37659 ( .A(n37318), .B(n37317), .Z(n37320) );
  XNOR U37660 ( .A(n37319), .B(n37320), .Z(n37315) );
  XOR U37661 ( .A(n37316), .B(n37315), .Z(c[237]) );
  AND U37662 ( .A(n37316), .B(n37315), .Z(n37410) );
  NANDN U37663 ( .A(n37318), .B(n37317), .Z(n37322) );
  OR U37664 ( .A(n37320), .B(n37319), .Z(n37321) );
  AND U37665 ( .A(n37322), .B(n37321), .Z(n37413) );
  NANDN U37666 ( .A(n37324), .B(n37323), .Z(n37328) );
  NANDN U37667 ( .A(n37326), .B(n37325), .Z(n37327) );
  AND U37668 ( .A(n37328), .B(n37327), .Z(n37419) );
  NANDN U37669 ( .A(n37330), .B(n37329), .Z(n37334) );
  NANDN U37670 ( .A(n37332), .B(n37331), .Z(n37333) );
  AND U37671 ( .A(n37334), .B(n37333), .Z(n37490) );
  NANDN U37672 ( .A(n37336), .B(n37335), .Z(n37340) );
  ANDN U37673 ( .B(n37338), .A(n37337), .Z(n37339) );
  ANDN U37674 ( .B(n37340), .A(n37339), .Z(n37479) );
  NAND U37675 ( .A(b[47]), .B(n37341), .Z(n37344) );
  ANDN U37676 ( .B(n37342), .A(n211), .Z(n37343) );
  ANDN U37677 ( .B(n37344), .A(n37343), .Z(n37459) );
  NAND U37678 ( .A(b[63]), .B(a[110]), .Z(n37468) );
  NANDN U37679 ( .A(n38278), .B(n37345), .Z(n37347) );
  XOR U37680 ( .A(b[63]), .B(a[112]), .Z(n37462) );
  NANDN U37681 ( .A(n38279), .B(n37462), .Z(n37346) );
  NAND U37682 ( .A(n37347), .B(n37346), .Z(n37457) );
  XOR U37683 ( .A(n37468), .B(n37457), .Z(n37458) );
  XNOR U37684 ( .A(n37459), .B(n37458), .Z(n37478) );
  XNOR U37685 ( .A(n37479), .B(n37478), .Z(n37480) );
  XOR U37686 ( .A(n37480), .B(n37481), .Z(n37491) );
  XNOR U37687 ( .A(n37490), .B(n37491), .Z(n37493) );
  NANDN U37688 ( .A(n38090), .B(n37352), .Z(n37354) );
  XOR U37689 ( .A(b[59]), .B(a[116]), .Z(n37469) );
  NANDN U37690 ( .A(n38130), .B(n37469), .Z(n37353) );
  AND U37691 ( .A(n37354), .B(n37353), .Z(n37441) );
  NANDN U37692 ( .A(n38247), .B(n37355), .Z(n37357) );
  XOR U37693 ( .A(b[61]), .B(a[114]), .Z(n37472) );
  NANDN U37694 ( .A(n38248), .B(n37472), .Z(n37356) );
  AND U37695 ( .A(n37357), .B(n37356), .Z(n37440) );
  NANDN U37696 ( .A(n37358), .B(n38076), .Z(n37360) );
  XOR U37697 ( .A(b[57]), .B(a[118]), .Z(n37465) );
  NANDN U37698 ( .A(n38031), .B(n37465), .Z(n37359) );
  NAND U37699 ( .A(n37360), .B(n37359), .Z(n37439) );
  XOR U37700 ( .A(n37440), .B(n37439), .Z(n37442) );
  XOR U37701 ( .A(n37441), .B(n37442), .Z(n37453) );
  NANDN U37702 ( .A(n37361), .B(n37849), .Z(n37363) );
  XOR U37703 ( .A(a[122]), .B(b[53]), .Z(n37475) );
  NANDN U37704 ( .A(n37778), .B(n37475), .Z(n37362) );
  AND U37705 ( .A(n37363), .B(n37362), .Z(n37447) );
  NANDN U37706 ( .A(n37857), .B(n37364), .Z(n37366) );
  XOR U37707 ( .A(b[55]), .B(a[120]), .Z(n37436) );
  NANDN U37708 ( .A(n37911), .B(n37436), .Z(n37365) );
  AND U37709 ( .A(n37366), .B(n37365), .Z(n37446) );
  NANDN U37710 ( .A(n212), .B(n37367), .Z(n37369) );
  XOR U37711 ( .A(a[126]), .B(b[49]), .Z(n37433) );
  NANDN U37712 ( .A(n37432), .B(n37433), .Z(n37368) );
  NAND U37713 ( .A(n37369), .B(n37368), .Z(n37445) );
  XOR U37714 ( .A(n37446), .B(n37445), .Z(n37448) );
  XOR U37715 ( .A(n37447), .B(n37448), .Z(n37452) );
  NAND U37716 ( .A(n37733), .B(n37370), .Z(n37372) );
  XNOR U37717 ( .A(a[124]), .B(b[51]), .Z(n37429) );
  NANDN U37718 ( .A(n37429), .B(n37734), .Z(n37371) );
  AND U37719 ( .A(n37372), .B(n37371), .Z(n37451) );
  XOR U37720 ( .A(n37452), .B(n37451), .Z(n37454) );
  XOR U37721 ( .A(n37453), .B(n37454), .Z(n37487) );
  NANDN U37722 ( .A(n37374), .B(n37373), .Z(n37378) );
  OR U37723 ( .A(n37376), .B(n37375), .Z(n37377) );
  AND U37724 ( .A(n37378), .B(n37377), .Z(n37485) );
  NANDN U37725 ( .A(n37380), .B(n37379), .Z(n37384) );
  OR U37726 ( .A(n37382), .B(n37381), .Z(n37383) );
  NAND U37727 ( .A(n37384), .B(n37383), .Z(n37484) );
  XNOR U37728 ( .A(n37485), .B(n37484), .Z(n37486) );
  XNOR U37729 ( .A(n37487), .B(n37486), .Z(n37492) );
  XOR U37730 ( .A(n37493), .B(n37492), .Z(n37425) );
  NANDN U37731 ( .A(n37386), .B(n37385), .Z(n37390) );
  NAND U37732 ( .A(n37388), .B(n37387), .Z(n37389) );
  AND U37733 ( .A(n37390), .B(n37389), .Z(n37424) );
  NANDN U37734 ( .A(n37392), .B(n37391), .Z(n37396) );
  NAND U37735 ( .A(n37394), .B(n37393), .Z(n37395) );
  NAND U37736 ( .A(n37396), .B(n37395), .Z(n37423) );
  XOR U37737 ( .A(n37424), .B(n37423), .Z(n37426) );
  XOR U37738 ( .A(n37425), .B(n37426), .Z(n37418) );
  NANDN U37739 ( .A(n37398), .B(n37397), .Z(n37402) );
  NANDN U37740 ( .A(n37400), .B(n37399), .Z(n37401) );
  NAND U37741 ( .A(n37402), .B(n37401), .Z(n37417) );
  XOR U37742 ( .A(n37418), .B(n37417), .Z(n37420) );
  XOR U37743 ( .A(n37419), .B(n37420), .Z(n37412) );
  NANDN U37744 ( .A(n37404), .B(n37403), .Z(n37408) );
  NAND U37745 ( .A(n37406), .B(n37405), .Z(n37407) );
  AND U37746 ( .A(n37408), .B(n37407), .Z(n37411) );
  XOR U37747 ( .A(n37412), .B(n37411), .Z(n37414) );
  XNOR U37748 ( .A(n37413), .B(n37414), .Z(n37409) );
  XOR U37749 ( .A(n37410), .B(n37409), .Z(c[238]) );
  AND U37750 ( .A(n37410), .B(n37409), .Z(n37497) );
  NANDN U37751 ( .A(n37412), .B(n37411), .Z(n37416) );
  OR U37752 ( .A(n37414), .B(n37413), .Z(n37415) );
  AND U37753 ( .A(n37416), .B(n37415), .Z(n37500) );
  NANDN U37754 ( .A(n37418), .B(n37417), .Z(n37422) );
  OR U37755 ( .A(n37420), .B(n37419), .Z(n37421) );
  AND U37756 ( .A(n37422), .B(n37421), .Z(n37498) );
  NANDN U37757 ( .A(n37424), .B(n37423), .Z(n37428) );
  OR U37758 ( .A(n37426), .B(n37425), .Z(n37427) );
  AND U37759 ( .A(n37428), .B(n37427), .Z(n37507) );
  NANDN U37760 ( .A(n37429), .B(n37733), .Z(n37431) );
  XOR U37761 ( .A(a[125]), .B(b[51]), .Z(n37525) );
  NANDN U37762 ( .A(n37605), .B(n37525), .Z(n37430) );
  AND U37763 ( .A(n37431), .B(n37430), .Z(n37542) );
  XNOR U37764 ( .A(a[127]), .B(b[49]), .Z(n37535) );
  OR U37765 ( .A(n37535), .B(n37432), .Z(n37435) );
  NAND U37766 ( .A(n37536), .B(n37433), .Z(n37434) );
  AND U37767 ( .A(n37435), .B(n37434), .Z(n37541) );
  NANDN U37768 ( .A(n37857), .B(n37436), .Z(n37438) );
  XOR U37769 ( .A(b[55]), .B(a[121]), .Z(n37564) );
  NANDN U37770 ( .A(n37911), .B(n37564), .Z(n37437) );
  NAND U37771 ( .A(n37438), .B(n37437), .Z(n37540) );
  XOR U37772 ( .A(n37541), .B(n37540), .Z(n37543) );
  XOR U37773 ( .A(n37542), .B(n37543), .Z(n37568) );
  NANDN U37774 ( .A(n37440), .B(n37439), .Z(n37444) );
  OR U37775 ( .A(n37442), .B(n37441), .Z(n37443) );
  AND U37776 ( .A(n37444), .B(n37443), .Z(n37567) );
  XNOR U37777 ( .A(n37568), .B(n37567), .Z(n37570) );
  NANDN U37778 ( .A(n37446), .B(n37445), .Z(n37450) );
  OR U37779 ( .A(n37448), .B(n37447), .Z(n37449) );
  AND U37780 ( .A(n37450), .B(n37449), .Z(n37569) );
  XOR U37781 ( .A(n37570), .B(n37569), .Z(n37581) );
  NANDN U37782 ( .A(n37452), .B(n37451), .Z(n37456) );
  OR U37783 ( .A(n37454), .B(n37453), .Z(n37455) );
  AND U37784 ( .A(n37456), .B(n37455), .Z(n37579) );
  IV U37785 ( .A(n37468), .Z(n37555) );
  NANDN U37786 ( .A(n37555), .B(n37457), .Z(n37461) );
  NANDN U37787 ( .A(n37459), .B(n37458), .Z(n37460) );
  AND U37788 ( .A(n37461), .B(n37460), .Z(n37576) );
  NANDN U37789 ( .A(n38278), .B(n37462), .Z(n37464) );
  XOR U37790 ( .A(b[63]), .B(a[113]), .Z(n37532) );
  NANDN U37791 ( .A(n38279), .B(n37532), .Z(n37463) );
  AND U37792 ( .A(n37464), .B(n37463), .Z(n37517) );
  NANDN U37793 ( .A(n37974), .B(n37465), .Z(n37467) );
  XOR U37794 ( .A(b[57]), .B(a[119]), .Z(n37558) );
  NANDN U37795 ( .A(n38031), .B(n37558), .Z(n37466) );
  NAND U37796 ( .A(n37467), .B(n37466), .Z(n37516) );
  XNOR U37797 ( .A(n37517), .B(n37516), .Z(n37518) );
  AND U37798 ( .A(b[63]), .B(a[111]), .Z(n37552) );
  XOR U37799 ( .A(n37553), .B(n37552), .Z(n37554) );
  XOR U37800 ( .A(n37468), .B(n37554), .Z(n37519) );
  XOR U37801 ( .A(n37518), .B(n37519), .Z(n37573) );
  NANDN U37802 ( .A(n38090), .B(n37469), .Z(n37471) );
  XOR U37803 ( .A(b[59]), .B(a[117]), .Z(n37529) );
  NANDN U37804 ( .A(n38130), .B(n37529), .Z(n37470) );
  AND U37805 ( .A(n37471), .B(n37470), .Z(n37549) );
  NANDN U37806 ( .A(n38247), .B(n37472), .Z(n37474) );
  XOR U37807 ( .A(b[61]), .B(a[115]), .Z(n37561) );
  NANDN U37808 ( .A(n38248), .B(n37561), .Z(n37473) );
  AND U37809 ( .A(n37474), .B(n37473), .Z(n37547) );
  NANDN U37810 ( .A(n37705), .B(n37475), .Z(n37477) );
  XOR U37811 ( .A(a[123]), .B(b[53]), .Z(n37522) );
  NANDN U37812 ( .A(n37778), .B(n37522), .Z(n37476) );
  NAND U37813 ( .A(n37477), .B(n37476), .Z(n37546) );
  XNOR U37814 ( .A(n37547), .B(n37546), .Z(n37548) );
  XOR U37815 ( .A(n37549), .B(n37548), .Z(n37574) );
  XNOR U37816 ( .A(n37573), .B(n37574), .Z(n37575) );
  XOR U37817 ( .A(n37576), .B(n37575), .Z(n37580) );
  XOR U37818 ( .A(n37579), .B(n37580), .Z(n37582) );
  XOR U37819 ( .A(n37581), .B(n37582), .Z(n37513) );
  NANDN U37820 ( .A(n37479), .B(n37478), .Z(n37483) );
  NANDN U37821 ( .A(n37481), .B(n37480), .Z(n37482) );
  AND U37822 ( .A(n37483), .B(n37482), .Z(n37510) );
  NANDN U37823 ( .A(n37485), .B(n37484), .Z(n37489) );
  NANDN U37824 ( .A(n37487), .B(n37486), .Z(n37488) );
  NAND U37825 ( .A(n37489), .B(n37488), .Z(n37511) );
  XNOR U37826 ( .A(n37510), .B(n37511), .Z(n37512) );
  XNOR U37827 ( .A(n37513), .B(n37512), .Z(n37504) );
  NANDN U37828 ( .A(n37491), .B(n37490), .Z(n37495) );
  NAND U37829 ( .A(n37493), .B(n37492), .Z(n37494) );
  NAND U37830 ( .A(n37495), .B(n37494), .Z(n37505) );
  XNOR U37831 ( .A(n37504), .B(n37505), .Z(n37506) );
  XOR U37832 ( .A(n37507), .B(n37506), .Z(n37499) );
  XOR U37833 ( .A(n37498), .B(n37499), .Z(n37501) );
  XNOR U37834 ( .A(n37500), .B(n37501), .Z(n37496) );
  XOR U37835 ( .A(n37497), .B(n37496), .Z(c[239]) );
  AND U37836 ( .A(n37497), .B(n37496), .Z(n37586) );
  NANDN U37837 ( .A(n37499), .B(n37498), .Z(n37503) );
  OR U37838 ( .A(n37501), .B(n37500), .Z(n37502) );
  AND U37839 ( .A(n37503), .B(n37502), .Z(n37589) );
  NANDN U37840 ( .A(n37505), .B(n37504), .Z(n37509) );
  NANDN U37841 ( .A(n37507), .B(n37506), .Z(n37508) );
  AND U37842 ( .A(n37509), .B(n37508), .Z(n37588) );
  NANDN U37843 ( .A(n37511), .B(n37510), .Z(n37515) );
  NANDN U37844 ( .A(n37513), .B(n37512), .Z(n37514) );
  AND U37845 ( .A(n37515), .B(n37514), .Z(n37596) );
  NANDN U37846 ( .A(n37517), .B(n37516), .Z(n37521) );
  NAND U37847 ( .A(n37519), .B(n37518), .Z(n37520) );
  AND U37848 ( .A(n37521), .B(n37520), .Z(n37658) );
  NANDN U37849 ( .A(n37705), .B(n37522), .Z(n37524) );
  XOR U37850 ( .A(a[124]), .B(b[53]), .Z(n37618) );
  NANDN U37851 ( .A(n37778), .B(n37618), .Z(n37523) );
  AND U37852 ( .A(n37524), .B(n37523), .Z(n37647) );
  NANDN U37853 ( .A(n37526), .B(n37525), .Z(n37528) );
  XOR U37854 ( .A(a[126]), .B(b[51]), .Z(n37606) );
  NANDN U37855 ( .A(n37605), .B(n37606), .Z(n37527) );
  AND U37856 ( .A(n37528), .B(n37527), .Z(n37646) );
  NANDN U37857 ( .A(n38090), .B(n37529), .Z(n37531) );
  XOR U37858 ( .A(b[59]), .B(a[118]), .Z(n37609) );
  NANDN U37859 ( .A(n38130), .B(n37609), .Z(n37530) );
  NAND U37860 ( .A(n37531), .B(n37530), .Z(n37645) );
  XOR U37861 ( .A(n37646), .B(n37645), .Z(n37648) );
  XOR U37862 ( .A(n37647), .B(n37648), .Z(n37634) );
  NANDN U37863 ( .A(n38278), .B(n37532), .Z(n37534) );
  XOR U37864 ( .A(b[63]), .B(a[114]), .Z(n37621) );
  NANDN U37865 ( .A(n38279), .B(n37621), .Z(n37533) );
  AND U37866 ( .A(n37534), .B(n37533), .Z(n37654) );
  NAND U37867 ( .A(b[63]), .B(a[112]), .Z(n37651) );
  ANDN U37868 ( .B(n37536), .A(n37535), .Z(n37539) );
  NAND U37869 ( .A(b[49]), .B(n37537), .Z(n37538) );
  NANDN U37870 ( .A(n37539), .B(n37538), .Z(n37652) );
  XOR U37871 ( .A(n37651), .B(n37652), .Z(n37653) );
  XOR U37872 ( .A(n37654), .B(n37653), .Z(n37633) );
  XNOR U37873 ( .A(n37634), .B(n37633), .Z(n37636) );
  NANDN U37874 ( .A(n37541), .B(n37540), .Z(n37545) );
  OR U37875 ( .A(n37543), .B(n37542), .Z(n37544) );
  AND U37876 ( .A(n37545), .B(n37544), .Z(n37635) );
  XNOR U37877 ( .A(n37636), .B(n37635), .Z(n37657) );
  XNOR U37878 ( .A(n37658), .B(n37657), .Z(n37660) );
  NANDN U37879 ( .A(n37547), .B(n37546), .Z(n37551) );
  NANDN U37880 ( .A(n37549), .B(n37548), .Z(n37550) );
  AND U37881 ( .A(n37551), .B(n37550), .Z(n37642) );
  NANDN U37882 ( .A(n37553), .B(n37552), .Z(n37557) );
  ANDN U37883 ( .B(n37555), .A(n37554), .Z(n37556) );
  ANDN U37884 ( .B(n37557), .A(n37556), .Z(n37640) );
  NANDN U37885 ( .A(n37974), .B(n37558), .Z(n37560) );
  XOR U37886 ( .A(b[57]), .B(a[120]), .Z(n37624) );
  NANDN U37887 ( .A(n38031), .B(n37624), .Z(n37559) );
  AND U37888 ( .A(n37560), .B(n37559), .Z(n37630) );
  NANDN U37889 ( .A(n38247), .B(n37561), .Z(n37563) );
  XOR U37890 ( .A(b[61]), .B(a[116]), .Z(n37612) );
  NANDN U37891 ( .A(n38248), .B(n37612), .Z(n37562) );
  AND U37892 ( .A(n37563), .B(n37562), .Z(n37628) );
  NANDN U37893 ( .A(n37857), .B(n37564), .Z(n37566) );
  XOR U37894 ( .A(a[122]), .B(b[55]), .Z(n37615) );
  NANDN U37895 ( .A(n37911), .B(n37615), .Z(n37565) );
  NAND U37896 ( .A(n37566), .B(n37565), .Z(n37627) );
  XNOR U37897 ( .A(n37628), .B(n37627), .Z(n37629) );
  XNOR U37898 ( .A(n37630), .B(n37629), .Z(n37639) );
  XNOR U37899 ( .A(n37640), .B(n37639), .Z(n37641) );
  XNOR U37900 ( .A(n37642), .B(n37641), .Z(n37659) );
  XOR U37901 ( .A(n37660), .B(n37659), .Z(n37602) );
  NANDN U37902 ( .A(n37568), .B(n37567), .Z(n37572) );
  NAND U37903 ( .A(n37570), .B(n37569), .Z(n37571) );
  AND U37904 ( .A(n37572), .B(n37571), .Z(n37600) );
  NANDN U37905 ( .A(n37574), .B(n37573), .Z(n37578) );
  NANDN U37906 ( .A(n37576), .B(n37575), .Z(n37577) );
  AND U37907 ( .A(n37578), .B(n37577), .Z(n37599) );
  XNOR U37908 ( .A(n37600), .B(n37599), .Z(n37601) );
  XNOR U37909 ( .A(n37602), .B(n37601), .Z(n37593) );
  NANDN U37910 ( .A(n37580), .B(n37579), .Z(n37584) );
  OR U37911 ( .A(n37582), .B(n37581), .Z(n37583) );
  NAND U37912 ( .A(n37584), .B(n37583), .Z(n37594) );
  XNOR U37913 ( .A(n37593), .B(n37594), .Z(n37595) );
  XNOR U37914 ( .A(n37596), .B(n37595), .Z(n37587) );
  XOR U37915 ( .A(n37588), .B(n37587), .Z(n37590) );
  XNOR U37916 ( .A(n37589), .B(n37590), .Z(n37585) );
  XOR U37917 ( .A(n37586), .B(n37585), .Z(c[240]) );
  AND U37918 ( .A(n37586), .B(n37585), .Z(n37664) );
  NANDN U37919 ( .A(n37588), .B(n37587), .Z(n37592) );
  OR U37920 ( .A(n37590), .B(n37589), .Z(n37591) );
  AND U37921 ( .A(n37592), .B(n37591), .Z(n37667) );
  NANDN U37922 ( .A(n37594), .B(n37593), .Z(n37598) );
  NANDN U37923 ( .A(n37596), .B(n37595), .Z(n37597) );
  AND U37924 ( .A(n37598), .B(n37597), .Z(n37666) );
  NANDN U37925 ( .A(n37600), .B(n37599), .Z(n37604) );
  NANDN U37926 ( .A(n37602), .B(n37601), .Z(n37603) );
  AND U37927 ( .A(n37604), .B(n37603), .Z(n37674) );
  XNOR U37928 ( .A(a[127]), .B(b[51]), .Z(n37732) );
  OR U37929 ( .A(n37732), .B(n37605), .Z(n37608) );
  NAND U37930 ( .A(n37733), .B(n37606), .Z(n37607) );
  AND U37931 ( .A(n37608), .B(n37607), .Z(n37718) );
  NANDN U37932 ( .A(n38090), .B(n37609), .Z(n37611) );
  XOR U37933 ( .A(b[59]), .B(a[119]), .Z(n37714) );
  NANDN U37934 ( .A(n38130), .B(n37714), .Z(n37610) );
  NAND U37935 ( .A(n37611), .B(n37610), .Z(n37717) );
  XNOR U37936 ( .A(n37718), .B(n37717), .Z(n37720) );
  AND U37937 ( .A(b[63]), .B(a[113]), .Z(n37723) );
  XOR U37938 ( .A(n37724), .B(n37723), .Z(n37725) );
  XOR U37939 ( .A(n37651), .B(n37725), .Z(n37719) );
  XOR U37940 ( .A(n37720), .B(n37719), .Z(n37690) );
  NANDN U37941 ( .A(n38247), .B(n37612), .Z(n37614) );
  XOR U37942 ( .A(b[61]), .B(a[117]), .Z(n37711) );
  NANDN U37943 ( .A(n38248), .B(n37711), .Z(n37613) );
  AND U37944 ( .A(n37614), .B(n37613), .Z(n37739) );
  NANDN U37945 ( .A(n37857), .B(n37615), .Z(n37617) );
  XOR U37946 ( .A(a[123]), .B(b[55]), .Z(n37701) );
  NANDN U37947 ( .A(n37911), .B(n37701), .Z(n37616) );
  AND U37948 ( .A(n37617), .B(n37616), .Z(n37738) );
  NANDN U37949 ( .A(n37705), .B(n37618), .Z(n37620) );
  XOR U37950 ( .A(a[125]), .B(b[53]), .Z(n37704) );
  NANDN U37951 ( .A(n37778), .B(n37704), .Z(n37619) );
  AND U37952 ( .A(n37620), .B(n37619), .Z(n37698) );
  NANDN U37953 ( .A(n38278), .B(n37621), .Z(n37623) );
  XOR U37954 ( .A(b[63]), .B(a[115]), .Z(n37729) );
  NANDN U37955 ( .A(n38279), .B(n37729), .Z(n37622) );
  AND U37956 ( .A(n37623), .B(n37622), .Z(n37696) );
  NANDN U37957 ( .A(n37974), .B(n37624), .Z(n37626) );
  XOR U37958 ( .A(b[57]), .B(a[121]), .Z(n37708) );
  NANDN U37959 ( .A(n38031), .B(n37708), .Z(n37625) );
  NAND U37960 ( .A(n37626), .B(n37625), .Z(n37695) );
  XNOR U37961 ( .A(n37696), .B(n37695), .Z(n37697) );
  XNOR U37962 ( .A(n37698), .B(n37697), .Z(n37737) );
  XOR U37963 ( .A(n37738), .B(n37737), .Z(n37740) );
  XNOR U37964 ( .A(n37739), .B(n37740), .Z(n37689) );
  XNOR U37965 ( .A(n37690), .B(n37689), .Z(n37692) );
  NANDN U37966 ( .A(n37628), .B(n37627), .Z(n37632) );
  NANDN U37967 ( .A(n37630), .B(n37629), .Z(n37631) );
  AND U37968 ( .A(n37632), .B(n37631), .Z(n37691) );
  XOR U37969 ( .A(n37692), .B(n37691), .Z(n37678) );
  NANDN U37970 ( .A(n37634), .B(n37633), .Z(n37638) );
  NAND U37971 ( .A(n37636), .B(n37635), .Z(n37637) );
  AND U37972 ( .A(n37638), .B(n37637), .Z(n37677) );
  XNOR U37973 ( .A(n37678), .B(n37677), .Z(n37680) );
  NANDN U37974 ( .A(n37640), .B(n37639), .Z(n37644) );
  NANDN U37975 ( .A(n37642), .B(n37641), .Z(n37643) );
  AND U37976 ( .A(n37644), .B(n37643), .Z(n37686) );
  NANDN U37977 ( .A(n37646), .B(n37645), .Z(n37650) );
  OR U37978 ( .A(n37648), .B(n37647), .Z(n37649) );
  AND U37979 ( .A(n37650), .B(n37649), .Z(n37684) );
  IV U37980 ( .A(n37651), .Z(n37726) );
  NANDN U37981 ( .A(n37726), .B(n37652), .Z(n37656) );
  NANDN U37982 ( .A(n37654), .B(n37653), .Z(n37655) );
  NAND U37983 ( .A(n37656), .B(n37655), .Z(n37683) );
  XNOR U37984 ( .A(n37684), .B(n37683), .Z(n37685) );
  XNOR U37985 ( .A(n37686), .B(n37685), .Z(n37679) );
  XOR U37986 ( .A(n37680), .B(n37679), .Z(n37672) );
  NANDN U37987 ( .A(n37658), .B(n37657), .Z(n37662) );
  NAND U37988 ( .A(n37660), .B(n37659), .Z(n37661) );
  AND U37989 ( .A(n37662), .B(n37661), .Z(n37671) );
  XNOR U37990 ( .A(n37672), .B(n37671), .Z(n37673) );
  XNOR U37991 ( .A(n37674), .B(n37673), .Z(n37665) );
  XOR U37992 ( .A(n37666), .B(n37665), .Z(n37668) );
  XNOR U37993 ( .A(n37667), .B(n37668), .Z(n37663) );
  XOR U37994 ( .A(n37664), .B(n37663), .Z(c[241]) );
  AND U37995 ( .A(n37664), .B(n37663), .Z(n37744) );
  NANDN U37996 ( .A(n37666), .B(n37665), .Z(n37670) );
  OR U37997 ( .A(n37668), .B(n37667), .Z(n37669) );
  AND U37998 ( .A(n37670), .B(n37669), .Z(n37747) );
  NANDN U37999 ( .A(n37672), .B(n37671), .Z(n37676) );
  NANDN U38000 ( .A(n37674), .B(n37673), .Z(n37675) );
  AND U38001 ( .A(n37676), .B(n37675), .Z(n37746) );
  NANDN U38002 ( .A(n37678), .B(n37677), .Z(n37682) );
  NAND U38003 ( .A(n37680), .B(n37679), .Z(n37681) );
  AND U38004 ( .A(n37682), .B(n37681), .Z(n37753) );
  NANDN U38005 ( .A(n37684), .B(n37683), .Z(n37688) );
  NANDN U38006 ( .A(n37686), .B(n37685), .Z(n37687) );
  AND U38007 ( .A(n37688), .B(n37687), .Z(n37751) );
  NANDN U38008 ( .A(n37690), .B(n37689), .Z(n37694) );
  NAND U38009 ( .A(n37692), .B(n37691), .Z(n37693) );
  AND U38010 ( .A(n37694), .B(n37693), .Z(n37806) );
  NANDN U38011 ( .A(n37696), .B(n37695), .Z(n37700) );
  NANDN U38012 ( .A(n37698), .B(n37697), .Z(n37699) );
  AND U38013 ( .A(n37700), .B(n37699), .Z(n37798) );
  NANDN U38014 ( .A(n37857), .B(n37701), .Z(n37703) );
  XOR U38015 ( .A(a[124]), .B(b[55]), .Z(n37772) );
  NANDN U38016 ( .A(n37911), .B(n37772), .Z(n37702) );
  AND U38017 ( .A(n37703), .B(n37702), .Z(n37788) );
  NANDN U38018 ( .A(n37705), .B(n37704), .Z(n37707) );
  XOR U38019 ( .A(a[126]), .B(b[53]), .Z(n37779) );
  NANDN U38020 ( .A(n37778), .B(n37779), .Z(n37706) );
  AND U38021 ( .A(n37707), .B(n37706), .Z(n37786) );
  NANDN U38022 ( .A(n37974), .B(n37708), .Z(n37710) );
  XOR U38023 ( .A(b[57]), .B(a[122]), .Z(n37769) );
  NANDN U38024 ( .A(n38031), .B(n37769), .Z(n37709) );
  AND U38025 ( .A(n37710), .B(n37709), .Z(n37760) );
  NANDN U38026 ( .A(n38247), .B(n37711), .Z(n37713) );
  XOR U38027 ( .A(b[61]), .B(a[118]), .Z(n37766) );
  NANDN U38028 ( .A(n38248), .B(n37766), .Z(n37712) );
  AND U38029 ( .A(n37713), .B(n37712), .Z(n37758) );
  NANDN U38030 ( .A(n38090), .B(n37714), .Z(n37716) );
  XOR U38031 ( .A(b[59]), .B(a[120]), .Z(n37782) );
  NANDN U38032 ( .A(n38130), .B(n37782), .Z(n37715) );
  NAND U38033 ( .A(n37716), .B(n37715), .Z(n37757) );
  XNOR U38034 ( .A(n37758), .B(n37757), .Z(n37759) );
  XNOR U38035 ( .A(n37760), .B(n37759), .Z(n37785) );
  XNOR U38036 ( .A(n37786), .B(n37785), .Z(n37787) );
  XNOR U38037 ( .A(n37788), .B(n37787), .Z(n37797) );
  XNOR U38038 ( .A(n37798), .B(n37797), .Z(n37800) );
  NANDN U38039 ( .A(n37718), .B(n37717), .Z(n37722) );
  NAND U38040 ( .A(n37720), .B(n37719), .Z(n37721) );
  AND U38041 ( .A(n37722), .B(n37721), .Z(n37794) );
  NANDN U38042 ( .A(n37724), .B(n37723), .Z(n37728) );
  ANDN U38043 ( .B(n37726), .A(n37725), .Z(n37727) );
  ANDN U38044 ( .B(n37728), .A(n37727), .Z(n37792) );
  NANDN U38045 ( .A(n38278), .B(n37729), .Z(n37731) );
  XOR U38046 ( .A(b[63]), .B(a[116]), .Z(n37775) );
  NANDN U38047 ( .A(n38279), .B(n37775), .Z(n37730) );
  AND U38048 ( .A(n37731), .B(n37730), .Z(n37765) );
  NAND U38049 ( .A(b[63]), .B(a[114]), .Z(n37830) );
  ANDN U38050 ( .B(n37733), .A(n37732), .Z(n37736) );
  NAND U38051 ( .A(b[51]), .B(n37734), .Z(n37735) );
  NANDN U38052 ( .A(n37736), .B(n37735), .Z(n37763) );
  XOR U38053 ( .A(n37830), .B(n37763), .Z(n37764) );
  XNOR U38054 ( .A(n37765), .B(n37764), .Z(n37791) );
  XNOR U38055 ( .A(n37792), .B(n37791), .Z(n37793) );
  XNOR U38056 ( .A(n37794), .B(n37793), .Z(n37799) );
  XOR U38057 ( .A(n37800), .B(n37799), .Z(n37804) );
  NANDN U38058 ( .A(n37738), .B(n37737), .Z(n37742) );
  OR U38059 ( .A(n37740), .B(n37739), .Z(n37741) );
  AND U38060 ( .A(n37742), .B(n37741), .Z(n37803) );
  XNOR U38061 ( .A(n37804), .B(n37803), .Z(n37805) );
  XOR U38062 ( .A(n37806), .B(n37805), .Z(n37752) );
  XOR U38063 ( .A(n37751), .B(n37752), .Z(n37754) );
  XNOR U38064 ( .A(n37753), .B(n37754), .Z(n37745) );
  XOR U38065 ( .A(n37746), .B(n37745), .Z(n37748) );
  XNOR U38066 ( .A(n37747), .B(n37748), .Z(n37743) );
  XOR U38067 ( .A(n37744), .B(n37743), .Z(c[242]) );
  AND U38068 ( .A(n37744), .B(n37743), .Z(n37810) );
  NANDN U38069 ( .A(n37746), .B(n37745), .Z(n37750) );
  OR U38070 ( .A(n37748), .B(n37747), .Z(n37749) );
  AND U38071 ( .A(n37750), .B(n37749), .Z(n37813) );
  NANDN U38072 ( .A(n37752), .B(n37751), .Z(n37756) );
  NANDN U38073 ( .A(n37754), .B(n37753), .Z(n37755) );
  AND U38074 ( .A(n37756), .B(n37755), .Z(n37812) );
  NANDN U38075 ( .A(n37758), .B(n37757), .Z(n37762) );
  NANDN U38076 ( .A(n37760), .B(n37759), .Z(n37761) );
  AND U38077 ( .A(n37762), .B(n37761), .Z(n37872) );
  XNOR U38078 ( .A(n37872), .B(n37871), .Z(n37874) );
  NANDN U38079 ( .A(n38247), .B(n37766), .Z(n37768) );
  XOR U38080 ( .A(b[61]), .B(a[119]), .Z(n37863) );
  NANDN U38081 ( .A(n38248), .B(n37863), .Z(n37767) );
  AND U38082 ( .A(n37768), .B(n37767), .Z(n37868) );
  NANDN U38083 ( .A(n37974), .B(n37769), .Z(n37771) );
  XOR U38084 ( .A(b[57]), .B(a[123]), .Z(n37853) );
  NANDN U38085 ( .A(n38031), .B(n37853), .Z(n37770) );
  AND U38086 ( .A(n37771), .B(n37770), .Z(n37842) );
  NANDN U38087 ( .A(n37857), .B(n37772), .Z(n37774) );
  XOR U38088 ( .A(a[125]), .B(b[55]), .Z(n37856) );
  NANDN U38089 ( .A(n37911), .B(n37856), .Z(n37773) );
  AND U38090 ( .A(n37774), .B(n37773), .Z(n37840) );
  NANDN U38091 ( .A(n38278), .B(n37775), .Z(n37777) );
  XOR U38092 ( .A(b[63]), .B(a[117]), .Z(n37845) );
  NANDN U38093 ( .A(n38279), .B(n37845), .Z(n37776) );
  NAND U38094 ( .A(n37777), .B(n37776), .Z(n37839) );
  XNOR U38095 ( .A(n37840), .B(n37839), .Z(n37841) );
  XNOR U38096 ( .A(n37842), .B(n37841), .Z(n37867) );
  XNOR U38097 ( .A(n37868), .B(n37867), .Z(n37870) );
  XNOR U38098 ( .A(a[127]), .B(b[53]), .Z(n37848) );
  OR U38099 ( .A(n37848), .B(n37778), .Z(n37781) );
  NAND U38100 ( .A(n37849), .B(n37779), .Z(n37780) );
  AND U38101 ( .A(n37781), .B(n37780), .Z(n37834) );
  NANDN U38102 ( .A(n38090), .B(n37782), .Z(n37784) );
  XOR U38103 ( .A(b[59]), .B(a[121]), .Z(n37860) );
  NANDN U38104 ( .A(n38130), .B(n37860), .Z(n37783) );
  NAND U38105 ( .A(n37784), .B(n37783), .Z(n37833) );
  XNOR U38106 ( .A(n37834), .B(n37833), .Z(n37835) );
  AND U38107 ( .A(b[63]), .B(a[115]), .Z(n37832) );
  XOR U38108 ( .A(n37831), .B(n37832), .Z(n37829) );
  XNOR U38109 ( .A(n37830), .B(n37829), .Z(n37836) );
  XOR U38110 ( .A(n37835), .B(n37836), .Z(n37869) );
  XOR U38111 ( .A(n37870), .B(n37869), .Z(n37873) );
  XOR U38112 ( .A(n37874), .B(n37873), .Z(n37825) );
  NANDN U38113 ( .A(n37786), .B(n37785), .Z(n37790) );
  NANDN U38114 ( .A(n37788), .B(n37787), .Z(n37789) );
  AND U38115 ( .A(n37790), .B(n37789), .Z(n37823) );
  NANDN U38116 ( .A(n37792), .B(n37791), .Z(n37796) );
  NANDN U38117 ( .A(n37794), .B(n37793), .Z(n37795) );
  NAND U38118 ( .A(n37796), .B(n37795), .Z(n37824) );
  XOR U38119 ( .A(n37823), .B(n37824), .Z(n37826) );
  XOR U38120 ( .A(n37825), .B(n37826), .Z(n37818) );
  NANDN U38121 ( .A(n37798), .B(n37797), .Z(n37802) );
  NAND U38122 ( .A(n37800), .B(n37799), .Z(n37801) );
  NAND U38123 ( .A(n37802), .B(n37801), .Z(n37817) );
  XNOR U38124 ( .A(n37818), .B(n37817), .Z(n37820) );
  NANDN U38125 ( .A(n37804), .B(n37803), .Z(n37808) );
  NANDN U38126 ( .A(n37806), .B(n37805), .Z(n37807) );
  AND U38127 ( .A(n37808), .B(n37807), .Z(n37819) );
  XNOR U38128 ( .A(n37820), .B(n37819), .Z(n37811) );
  XOR U38129 ( .A(n37812), .B(n37811), .Z(n37814) );
  XNOR U38130 ( .A(n37813), .B(n37814), .Z(n37809) );
  XOR U38131 ( .A(n37810), .B(n37809), .Z(c[243]) );
  AND U38132 ( .A(n37810), .B(n37809), .Z(n37878) );
  NANDN U38133 ( .A(n37812), .B(n37811), .Z(n37816) );
  OR U38134 ( .A(n37814), .B(n37813), .Z(n37815) );
  AND U38135 ( .A(n37816), .B(n37815), .Z(n37881) );
  NANDN U38136 ( .A(n37818), .B(n37817), .Z(n37822) );
  NAND U38137 ( .A(n37820), .B(n37819), .Z(n37821) );
  AND U38138 ( .A(n37822), .B(n37821), .Z(n37879) );
  NANDN U38139 ( .A(n37824), .B(n37823), .Z(n37828) );
  OR U38140 ( .A(n37826), .B(n37825), .Z(n37827) );
  AND U38141 ( .A(n37828), .B(n37827), .Z(n37888) );
  NANDN U38142 ( .A(n37834), .B(n37833), .Z(n37838) );
  NAND U38143 ( .A(n37836), .B(n37835), .Z(n37837) );
  NAND U38144 ( .A(n37838), .B(n37837), .Z(n37894) );
  XNOR U38145 ( .A(n37893), .B(n37894), .Z(n37896) );
  NANDN U38146 ( .A(n37840), .B(n37839), .Z(n37844) );
  NANDN U38147 ( .A(n37842), .B(n37841), .Z(n37843) );
  AND U38148 ( .A(n37844), .B(n37843), .Z(n37895) );
  XOR U38149 ( .A(n37896), .B(n37895), .Z(n37892) );
  NANDN U38150 ( .A(n38278), .B(n37845), .Z(n37847) );
  XOR U38151 ( .A(b[63]), .B(a[118]), .Z(n37925) );
  NANDN U38152 ( .A(n38279), .B(n37925), .Z(n37846) );
  AND U38153 ( .A(n37847), .B(n37846), .Z(n37931) );
  NAND U38154 ( .A(b[63]), .B(a[116]), .Z(n37965) );
  ANDN U38155 ( .B(n37849), .A(n37848), .Z(n37852) );
  NAND U38156 ( .A(b[53]), .B(n37850), .Z(n37851) );
  NANDN U38157 ( .A(n37852), .B(n37851), .Z(n37928) );
  XOR U38158 ( .A(n37965), .B(n37928), .Z(n37930) );
  XOR U38159 ( .A(n37931), .B(n37930), .Z(n37901) );
  NANDN U38160 ( .A(n37974), .B(n37853), .Z(n37855) );
  XOR U38161 ( .A(a[124]), .B(b[57]), .Z(n37918) );
  NANDN U38162 ( .A(n38031), .B(n37918), .Z(n37854) );
  AND U38163 ( .A(n37855), .B(n37854), .Z(n37907) );
  NANDN U38164 ( .A(n37857), .B(n37856), .Z(n37859) );
  XOR U38165 ( .A(a[126]), .B(b[55]), .Z(n37912) );
  NANDN U38166 ( .A(n37911), .B(n37912), .Z(n37858) );
  AND U38167 ( .A(n37859), .B(n37858), .Z(n37906) );
  NANDN U38168 ( .A(n38090), .B(n37860), .Z(n37862) );
  XOR U38169 ( .A(b[59]), .B(a[122]), .Z(n37915) );
  NANDN U38170 ( .A(n38130), .B(n37915), .Z(n37861) );
  NAND U38171 ( .A(n37862), .B(n37861), .Z(n37905) );
  XOR U38172 ( .A(n37906), .B(n37905), .Z(n37908) );
  XOR U38173 ( .A(n37907), .B(n37908), .Z(n37900) );
  NAND U38174 ( .A(n37921), .B(n37863), .Z(n37866) );
  XNOR U38175 ( .A(b[61]), .B(a[120]), .Z(n37922) );
  NANDN U38176 ( .A(n37922), .B(n37864), .Z(n37865) );
  AND U38177 ( .A(n37866), .B(n37865), .Z(n37899) );
  XOR U38178 ( .A(n37900), .B(n37899), .Z(n37902) );
  XOR U38179 ( .A(n37901), .B(n37902), .Z(n37889) );
  XOR U38180 ( .A(n37889), .B(n37890), .Z(n37891) );
  XOR U38181 ( .A(n37892), .B(n37891), .Z(n37885) );
  NANDN U38182 ( .A(n37872), .B(n37871), .Z(n37876) );
  NAND U38183 ( .A(n37874), .B(n37873), .Z(n37875) );
  AND U38184 ( .A(n37876), .B(n37875), .Z(n37886) );
  XOR U38185 ( .A(n37885), .B(n37886), .Z(n37887) );
  XOR U38186 ( .A(n37888), .B(n37887), .Z(n37880) );
  XOR U38187 ( .A(n37879), .B(n37880), .Z(n37882) );
  XNOR U38188 ( .A(n37881), .B(n37882), .Z(n37877) );
  XOR U38189 ( .A(n37878), .B(n37877), .Z(c[244]) );
  AND U38190 ( .A(n37878), .B(n37877), .Z(n37935) );
  NANDN U38191 ( .A(n37880), .B(n37879), .Z(n37884) );
  OR U38192 ( .A(n37882), .B(n37881), .Z(n37883) );
  AND U38193 ( .A(n37884), .B(n37883), .Z(n37938) );
  NANDN U38194 ( .A(n37894), .B(n37893), .Z(n37898) );
  NAND U38195 ( .A(n37896), .B(n37895), .Z(n37897) );
  AND U38196 ( .A(n37898), .B(n37897), .Z(n37943) );
  NANDN U38197 ( .A(n37900), .B(n37899), .Z(n37904) );
  NANDN U38198 ( .A(n37902), .B(n37901), .Z(n37903) );
  AND U38199 ( .A(n37904), .B(n37903), .Z(n37951) );
  NANDN U38200 ( .A(n37906), .B(n37905), .Z(n37910) );
  OR U38201 ( .A(n37908), .B(n37907), .Z(n37909) );
  AND U38202 ( .A(n37910), .B(n37909), .Z(n37956) );
  XNOR U38203 ( .A(a[127]), .B(b[55]), .Z(n37983) );
  OR U38204 ( .A(n37983), .B(n37911), .Z(n37914) );
  NAND U38205 ( .A(n37984), .B(n37912), .Z(n37913) );
  AND U38206 ( .A(n37914), .B(n37913), .Z(n37961) );
  NANDN U38207 ( .A(n38090), .B(n37915), .Z(n37917) );
  XOR U38208 ( .A(b[59]), .B(a[123]), .Z(n37970) );
  NANDN U38209 ( .A(n38130), .B(n37970), .Z(n37916) );
  NAND U38210 ( .A(n37917), .B(n37916), .Z(n37960) );
  XNOR U38211 ( .A(n37961), .B(n37960), .Z(n37963) );
  IV U38212 ( .A(n37965), .Z(n37929) );
  XOR U38213 ( .A(n37964), .B(n37929), .Z(n37967) );
  AND U38214 ( .A(b[63]), .B(a[117]), .Z(n37966) );
  XOR U38215 ( .A(n37967), .B(n37966), .Z(n37962) );
  XOR U38216 ( .A(n37963), .B(n37962), .Z(n37954) );
  NANDN U38217 ( .A(n37974), .B(n37918), .Z(n37920) );
  XOR U38218 ( .A(a[125]), .B(b[57]), .Z(n37973) );
  NANDN U38219 ( .A(n38031), .B(n37973), .Z(n37919) );
  AND U38220 ( .A(n37920), .B(n37919), .Z(n37991) );
  NANDN U38221 ( .A(n37922), .B(n37921), .Z(n37924) );
  XOR U38222 ( .A(b[61]), .B(a[121]), .Z(n37977) );
  NANDN U38223 ( .A(n38248), .B(n37977), .Z(n37923) );
  AND U38224 ( .A(n37924), .B(n37923), .Z(n37989) );
  NANDN U38225 ( .A(n38278), .B(n37925), .Z(n37927) );
  XOR U38226 ( .A(b[63]), .B(a[119]), .Z(n37980) );
  NANDN U38227 ( .A(n38279), .B(n37980), .Z(n37926) );
  NAND U38228 ( .A(n37927), .B(n37926), .Z(n37988) );
  XNOR U38229 ( .A(n37989), .B(n37988), .Z(n37990) );
  XOR U38230 ( .A(n37991), .B(n37990), .Z(n37955) );
  XOR U38231 ( .A(n37954), .B(n37955), .Z(n37957) );
  XOR U38232 ( .A(n37956), .B(n37957), .Z(n37949) );
  NANDN U38233 ( .A(n37929), .B(n37928), .Z(n37933) );
  NANDN U38234 ( .A(n37931), .B(n37930), .Z(n37932) );
  AND U38235 ( .A(n37933), .B(n37932), .Z(n37948) );
  XNOR U38236 ( .A(n37949), .B(n37948), .Z(n37950) );
  XNOR U38237 ( .A(n37951), .B(n37950), .Z(n37942) );
  XOR U38238 ( .A(n37943), .B(n37942), .Z(n37945) );
  XNOR U38239 ( .A(n37944), .B(n37945), .Z(n37936) );
  XOR U38240 ( .A(n37937), .B(n37936), .Z(n37939) );
  XNOR U38241 ( .A(n37938), .B(n37939), .Z(n37934) );
  XOR U38242 ( .A(n37935), .B(n37934), .Z(c[245]) );
  AND U38243 ( .A(n37935), .B(n37934), .Z(n37995) );
  NANDN U38244 ( .A(n37937), .B(n37936), .Z(n37941) );
  OR U38245 ( .A(n37939), .B(n37938), .Z(n37940) );
  AND U38246 ( .A(n37941), .B(n37940), .Z(n37998) );
  NANDN U38247 ( .A(n37943), .B(n37942), .Z(n37947) );
  NANDN U38248 ( .A(n37945), .B(n37944), .Z(n37946) );
  AND U38249 ( .A(n37947), .B(n37946), .Z(n37997) );
  NANDN U38250 ( .A(n37949), .B(n37948), .Z(n37953) );
  NANDN U38251 ( .A(n37951), .B(n37950), .Z(n37952) );
  AND U38252 ( .A(n37953), .B(n37952), .Z(n38005) );
  NANDN U38253 ( .A(n37955), .B(n37954), .Z(n37959) );
  OR U38254 ( .A(n37957), .B(n37956), .Z(n37958) );
  AND U38255 ( .A(n37959), .B(n37958), .Z(n38002) );
  NANDN U38256 ( .A(n37965), .B(n37964), .Z(n37969) );
  NAND U38257 ( .A(n37967), .B(n37966), .Z(n37968) );
  NAND U38258 ( .A(n37969), .B(n37968), .Z(n38009) );
  XNOR U38259 ( .A(n38008), .B(n38009), .Z(n38010) );
  NANDN U38260 ( .A(n38090), .B(n37970), .Z(n37972) );
  XOR U38261 ( .A(b[59]), .B(a[124]), .Z(n38028) );
  NANDN U38262 ( .A(n38130), .B(n38028), .Z(n37971) );
  AND U38263 ( .A(n37972), .B(n37971), .Z(n38016) );
  NANDN U38264 ( .A(n37974), .B(n37973), .Z(n37976) );
  XOR U38265 ( .A(a[126]), .B(b[57]), .Z(n38032) );
  NANDN U38266 ( .A(n38031), .B(n38032), .Z(n37975) );
  AND U38267 ( .A(n37976), .B(n37975), .Z(n38015) );
  NANDN U38268 ( .A(n38247), .B(n37977), .Z(n37979) );
  XOR U38269 ( .A(b[61]), .B(a[122]), .Z(n38035) );
  NANDN U38270 ( .A(n38248), .B(n38035), .Z(n37978) );
  NAND U38271 ( .A(n37979), .B(n37978), .Z(n38014) );
  XOR U38272 ( .A(n38015), .B(n38014), .Z(n38017) );
  XOR U38273 ( .A(n38016), .B(n38017), .Z(n38041) );
  NANDN U38274 ( .A(n38278), .B(n37980), .Z(n37982) );
  XOR U38275 ( .A(b[63]), .B(a[120]), .Z(n38025) );
  NANDN U38276 ( .A(n38279), .B(n38025), .Z(n37981) );
  AND U38277 ( .A(n37982), .B(n37981), .Z(n38022) );
  NAND U38278 ( .A(b[63]), .B(a[118]), .Z(n38039) );
  ANDN U38279 ( .B(n37984), .A(n37983), .Z(n37987) );
  NAND U38280 ( .A(b[55]), .B(n37985), .Z(n37986) );
  NANDN U38281 ( .A(n37987), .B(n37986), .Z(n38020) );
  XOR U38282 ( .A(n38039), .B(n38020), .Z(n38021) );
  XOR U38283 ( .A(n38022), .B(n38021), .Z(n38040) );
  XNOR U38284 ( .A(n38041), .B(n38040), .Z(n38042) );
  NANDN U38285 ( .A(n37989), .B(n37988), .Z(n37993) );
  NANDN U38286 ( .A(n37991), .B(n37990), .Z(n37992) );
  NAND U38287 ( .A(n37993), .B(n37992), .Z(n38043) );
  XOR U38288 ( .A(n38042), .B(n38043), .Z(n38011) );
  XOR U38289 ( .A(n38010), .B(n38011), .Z(n38003) );
  XNOR U38290 ( .A(n38002), .B(n38003), .Z(n38004) );
  XNOR U38291 ( .A(n38005), .B(n38004), .Z(n37996) );
  XOR U38292 ( .A(n37997), .B(n37996), .Z(n37999) );
  XNOR U38293 ( .A(n37998), .B(n37999), .Z(n37994) );
  XOR U38294 ( .A(n37995), .B(n37994), .Z(c[246]) );
  AND U38295 ( .A(n37995), .B(n37994), .Z(n38047) );
  NANDN U38296 ( .A(n37997), .B(n37996), .Z(n38001) );
  OR U38297 ( .A(n37999), .B(n37998), .Z(n38000) );
  AND U38298 ( .A(n38001), .B(n38000), .Z(n38050) );
  NANDN U38299 ( .A(n38003), .B(n38002), .Z(n38007) );
  NANDN U38300 ( .A(n38005), .B(n38004), .Z(n38006) );
  AND U38301 ( .A(n38007), .B(n38006), .Z(n38049) );
  NANDN U38302 ( .A(n38009), .B(n38008), .Z(n38013) );
  NANDN U38303 ( .A(n38011), .B(n38010), .Z(n38012) );
  AND U38304 ( .A(n38013), .B(n38012), .Z(n38057) );
  NANDN U38305 ( .A(n38015), .B(n38014), .Z(n38019) );
  OR U38306 ( .A(n38017), .B(n38016), .Z(n38018) );
  AND U38307 ( .A(n38019), .B(n38018), .Z(n38062) );
  IV U38308 ( .A(n38039), .Z(n38083) );
  NANDN U38309 ( .A(n38083), .B(n38020), .Z(n38024) );
  NANDN U38310 ( .A(n38022), .B(n38021), .Z(n38023) );
  AND U38311 ( .A(n38024), .B(n38023), .Z(n38061) );
  NANDN U38312 ( .A(n38278), .B(n38025), .Z(n38027) );
  XOR U38313 ( .A(b[63]), .B(a[121]), .Z(n38072) );
  NANDN U38314 ( .A(n38279), .B(n38072), .Z(n38026) );
  AND U38315 ( .A(n38027), .B(n38026), .Z(n38096) );
  NANDN U38316 ( .A(n38090), .B(n38028), .Z(n38030) );
  XOR U38317 ( .A(b[59]), .B(a[125]), .Z(n38089) );
  NANDN U38318 ( .A(n38130), .B(n38089), .Z(n38029) );
  AND U38319 ( .A(n38030), .B(n38029), .Z(n38094) );
  XNOR U38320 ( .A(a[127]), .B(b[57]), .Z(n38075) );
  OR U38321 ( .A(n38075), .B(n38031), .Z(n38034) );
  NAND U38322 ( .A(n38076), .B(n38032), .Z(n38033) );
  AND U38323 ( .A(n38034), .B(n38033), .Z(n38067) );
  NANDN U38324 ( .A(n38247), .B(n38035), .Z(n38037) );
  XOR U38325 ( .A(b[61]), .B(a[123]), .Z(n38086) );
  NANDN U38326 ( .A(n38248), .B(n38086), .Z(n38036) );
  NAND U38327 ( .A(n38037), .B(n38036), .Z(n38066) );
  XNOR U38328 ( .A(n38067), .B(n38066), .Z(n38068) );
  IV U38329 ( .A(n38038), .Z(n38081) );
  AND U38330 ( .A(b[63]), .B(a[119]), .Z(n38080) );
  XOR U38331 ( .A(n38081), .B(n38080), .Z(n38082) );
  XOR U38332 ( .A(n38039), .B(n38082), .Z(n38069) );
  XOR U38333 ( .A(n38068), .B(n38069), .Z(n38093) );
  XNOR U38334 ( .A(n38094), .B(n38093), .Z(n38095) );
  XNOR U38335 ( .A(n38096), .B(n38095), .Z(n38060) );
  XOR U38336 ( .A(n38061), .B(n38060), .Z(n38063) );
  XOR U38337 ( .A(n38062), .B(n38063), .Z(n38055) );
  NANDN U38338 ( .A(n38041), .B(n38040), .Z(n38045) );
  NANDN U38339 ( .A(n38043), .B(n38042), .Z(n38044) );
  NAND U38340 ( .A(n38045), .B(n38044), .Z(n38054) );
  XNOR U38341 ( .A(n38055), .B(n38054), .Z(n38056) );
  XNOR U38342 ( .A(n38057), .B(n38056), .Z(n38048) );
  XOR U38343 ( .A(n38049), .B(n38048), .Z(n38051) );
  XNOR U38344 ( .A(n38050), .B(n38051), .Z(n38046) );
  XOR U38345 ( .A(n38047), .B(n38046), .Z(c[247]) );
  AND U38346 ( .A(n38047), .B(n38046), .Z(n38100) );
  NANDN U38347 ( .A(n38049), .B(n38048), .Z(n38053) );
  OR U38348 ( .A(n38051), .B(n38050), .Z(n38052) );
  AND U38349 ( .A(n38053), .B(n38052), .Z(n38103) );
  NANDN U38350 ( .A(n38055), .B(n38054), .Z(n38059) );
  NANDN U38351 ( .A(n38057), .B(n38056), .Z(n38058) );
  AND U38352 ( .A(n38059), .B(n38058), .Z(n38102) );
  NANDN U38353 ( .A(n38061), .B(n38060), .Z(n38065) );
  OR U38354 ( .A(n38063), .B(n38062), .Z(n38064) );
  AND U38355 ( .A(n38065), .B(n38064), .Z(n38109) );
  NANDN U38356 ( .A(n38067), .B(n38066), .Z(n38071) );
  NAND U38357 ( .A(n38069), .B(n38068), .Z(n38070) );
  AND U38358 ( .A(n38071), .B(n38070), .Z(n38114) );
  NANDN U38359 ( .A(n38278), .B(n38072), .Z(n38074) );
  XOR U38360 ( .A(b[63]), .B(a[122]), .Z(n38137) );
  NANDN U38361 ( .A(n38279), .B(n38137), .Z(n38073) );
  AND U38362 ( .A(n38074), .B(n38073), .Z(n38127) );
  NAND U38363 ( .A(b[63]), .B(a[120]), .Z(n38140) );
  ANDN U38364 ( .B(n38076), .A(n38075), .Z(n38079) );
  NAND U38365 ( .A(b[57]), .B(n38077), .Z(n38078) );
  NANDN U38366 ( .A(n38079), .B(n38078), .Z(n38125) );
  XOR U38367 ( .A(n38140), .B(n38125), .Z(n38126) );
  XNOR U38368 ( .A(n38127), .B(n38126), .Z(n38113) );
  XNOR U38369 ( .A(n38114), .B(n38113), .Z(n38116) );
  NANDN U38370 ( .A(n38081), .B(n38080), .Z(n38085) );
  ANDN U38371 ( .B(n38083), .A(n38082), .Z(n38084) );
  ANDN U38372 ( .B(n38085), .A(n38084), .Z(n38122) );
  NANDN U38373 ( .A(n38247), .B(n38086), .Z(n38088) );
  XOR U38374 ( .A(b[61]), .B(a[124]), .Z(n38134) );
  NANDN U38375 ( .A(n38248), .B(n38134), .Z(n38087) );
  AND U38376 ( .A(n38088), .B(n38087), .Z(n38120) );
  NANDN U38377 ( .A(n38090), .B(n38089), .Z(n38092) );
  XOR U38378 ( .A(a[126]), .B(b[59]), .Z(n38131) );
  NANDN U38379 ( .A(n38130), .B(n38131), .Z(n38091) );
  NAND U38380 ( .A(n38092), .B(n38091), .Z(n38119) );
  XNOR U38381 ( .A(n38120), .B(n38119), .Z(n38121) );
  XNOR U38382 ( .A(n38122), .B(n38121), .Z(n38115) );
  XOR U38383 ( .A(n38116), .B(n38115), .Z(n38108) );
  NANDN U38384 ( .A(n38094), .B(n38093), .Z(n38098) );
  NANDN U38385 ( .A(n38096), .B(n38095), .Z(n38097) );
  AND U38386 ( .A(n38098), .B(n38097), .Z(n38107) );
  XOR U38387 ( .A(n38108), .B(n38107), .Z(n38110) );
  XNOR U38388 ( .A(n38109), .B(n38110), .Z(n38101) );
  XOR U38389 ( .A(n38102), .B(n38101), .Z(n38104) );
  XNOR U38390 ( .A(n38103), .B(n38104), .Z(n38099) );
  XOR U38391 ( .A(n38100), .B(n38099), .Z(c[248]) );
  AND U38392 ( .A(n38100), .B(n38099), .Z(n38142) );
  NANDN U38393 ( .A(n38102), .B(n38101), .Z(n38106) );
  OR U38394 ( .A(n38104), .B(n38103), .Z(n38105) );
  AND U38395 ( .A(n38106), .B(n38105), .Z(n38145) );
  NANDN U38396 ( .A(n38108), .B(n38107), .Z(n38112) );
  NANDN U38397 ( .A(n38110), .B(n38109), .Z(n38111) );
  AND U38398 ( .A(n38112), .B(n38111), .Z(n38144) );
  NANDN U38399 ( .A(n38114), .B(n38113), .Z(n38118) );
  NAND U38400 ( .A(n38116), .B(n38115), .Z(n38117) );
  AND U38401 ( .A(n38118), .B(n38117), .Z(n38180) );
  NANDN U38402 ( .A(n38120), .B(n38119), .Z(n38124) );
  NANDN U38403 ( .A(n38122), .B(n38121), .Z(n38123) );
  AND U38404 ( .A(n38124), .B(n38123), .Z(n38179) );
  IV U38405 ( .A(n38140), .Z(n38165) );
  NANDN U38406 ( .A(n38165), .B(n38125), .Z(n38129) );
  NANDN U38407 ( .A(n38127), .B(n38126), .Z(n38128) );
  AND U38408 ( .A(n38129), .B(n38128), .Z(n38152) );
  XNOR U38409 ( .A(a[127]), .B(b[59]), .Z(n38173) );
  OR U38410 ( .A(n38173), .B(n38130), .Z(n38133) );
  NAND U38411 ( .A(n38174), .B(n38131), .Z(n38132) );
  AND U38412 ( .A(n38133), .B(n38132), .Z(n38150) );
  NANDN U38413 ( .A(n38247), .B(n38134), .Z(n38136) );
  XOR U38414 ( .A(b[61]), .B(a[125]), .Z(n38161) );
  NANDN U38415 ( .A(n38248), .B(n38161), .Z(n38135) );
  AND U38416 ( .A(n38136), .B(n38135), .Z(n38156) );
  NANDN U38417 ( .A(n38278), .B(n38137), .Z(n38139) );
  XOR U38418 ( .A(b[63]), .B(a[123]), .Z(n38170) );
  NANDN U38419 ( .A(n38279), .B(n38170), .Z(n38138) );
  NAND U38420 ( .A(n38139), .B(n38138), .Z(n38155) );
  XNOR U38421 ( .A(n38156), .B(n38155), .Z(n38157) );
  AND U38422 ( .A(b[63]), .B(a[121]), .Z(n38166) );
  XOR U38423 ( .A(n38167), .B(n38166), .Z(n38164) );
  XOR U38424 ( .A(n38140), .B(n38164), .Z(n38158) );
  XOR U38425 ( .A(n38157), .B(n38158), .Z(n38149) );
  XNOR U38426 ( .A(n38150), .B(n38149), .Z(n38151) );
  XNOR U38427 ( .A(n38152), .B(n38151), .Z(n38178) );
  XOR U38428 ( .A(n38179), .B(n38178), .Z(n38181) );
  XNOR U38429 ( .A(n38180), .B(n38181), .Z(n38143) );
  XOR U38430 ( .A(n38144), .B(n38143), .Z(n38146) );
  XNOR U38431 ( .A(n38145), .B(n38146), .Z(n38141) );
  XOR U38432 ( .A(n38142), .B(n38141), .Z(c[249]) );
  AND U38433 ( .A(n38142), .B(n38141), .Z(n38185) );
  NANDN U38434 ( .A(n38144), .B(n38143), .Z(n38148) );
  OR U38435 ( .A(n38146), .B(n38145), .Z(n38147) );
  AND U38436 ( .A(n38148), .B(n38147), .Z(n38188) );
  NANDN U38437 ( .A(n38150), .B(n38149), .Z(n38154) );
  NANDN U38438 ( .A(n38152), .B(n38151), .Z(n38153) );
  AND U38439 ( .A(n38154), .B(n38153), .Z(n38194) );
  NANDN U38440 ( .A(n38156), .B(n38155), .Z(n38160) );
  NAND U38441 ( .A(n38158), .B(n38157), .Z(n38159) );
  AND U38442 ( .A(n38160), .B(n38159), .Z(n38193) );
  NANDN U38443 ( .A(n38247), .B(n38161), .Z(n38163) );
  XOR U38444 ( .A(b[61]), .B(a[126]), .Z(n38207) );
  NANDN U38445 ( .A(n38248), .B(n38207), .Z(n38162) );
  AND U38446 ( .A(n38163), .B(n38162), .Z(n38199) );
  ANDN U38447 ( .B(n38165), .A(n38164), .Z(n38169) );
  NANDN U38448 ( .A(n38167), .B(n38166), .Z(n38168) );
  NANDN U38449 ( .A(n38169), .B(n38168), .Z(n38198) );
  XNOR U38450 ( .A(n38199), .B(n38198), .Z(n38200) );
  NANDN U38451 ( .A(n38278), .B(n38170), .Z(n38172) );
  XOR U38452 ( .A(b[63]), .B(a[124]), .Z(n38204) );
  NANDN U38453 ( .A(n38279), .B(n38204), .Z(n38171) );
  AND U38454 ( .A(n38172), .B(n38171), .Z(n38214) );
  NAND U38455 ( .A(b[63]), .B(a[122]), .Z(n38211) );
  ANDN U38456 ( .B(n38174), .A(n38173), .Z(n38177) );
  NAND U38457 ( .A(b[59]), .B(n38175), .Z(n38176) );
  NANDN U38458 ( .A(n38177), .B(n38176), .Z(n38212) );
  XOR U38459 ( .A(n38211), .B(n38212), .Z(n38213) );
  XOR U38460 ( .A(n38214), .B(n38213), .Z(n38201) );
  XNOR U38461 ( .A(n38200), .B(n38201), .Z(n38192) );
  XOR U38462 ( .A(n38193), .B(n38192), .Z(n38195) );
  XOR U38463 ( .A(n38194), .B(n38195), .Z(n38187) );
  NANDN U38464 ( .A(n38179), .B(n38178), .Z(n38183) );
  OR U38465 ( .A(n38181), .B(n38180), .Z(n38182) );
  AND U38466 ( .A(n38183), .B(n38182), .Z(n38186) );
  XOR U38467 ( .A(n38187), .B(n38186), .Z(n38189) );
  XNOR U38468 ( .A(n38188), .B(n38189), .Z(n38184) );
  XOR U38469 ( .A(n38185), .B(n38184), .Z(c[250]) );
  AND U38470 ( .A(n38185), .B(n38184), .Z(n38218) );
  NANDN U38471 ( .A(n38187), .B(n38186), .Z(n38191) );
  OR U38472 ( .A(n38189), .B(n38188), .Z(n38190) );
  AND U38473 ( .A(n38191), .B(n38190), .Z(n38221) );
  NANDN U38474 ( .A(n38193), .B(n38192), .Z(n38197) );
  OR U38475 ( .A(n38195), .B(n38194), .Z(n38196) );
  AND U38476 ( .A(n38197), .B(n38196), .Z(n38219) );
  NANDN U38477 ( .A(n38199), .B(n38198), .Z(n38203) );
  NANDN U38478 ( .A(n38201), .B(n38200), .Z(n38202) );
  AND U38479 ( .A(n38203), .B(n38202), .Z(n38227) );
  NANDN U38480 ( .A(n38278), .B(n38204), .Z(n38206) );
  XOR U38481 ( .A(b[63]), .B(a[125]), .Z(n38243) );
  NANDN U38482 ( .A(n38279), .B(n38243), .Z(n38205) );
  AND U38483 ( .A(n38206), .B(n38205), .Z(n38232) );
  NANDN U38484 ( .A(n38247), .B(n38207), .Z(n38209) );
  XOR U38485 ( .A(a[127]), .B(b[61]), .Z(n38246) );
  NANDN U38486 ( .A(n38248), .B(n38246), .Z(n38208) );
  NAND U38487 ( .A(n38209), .B(n38208), .Z(n38231) );
  XNOR U38488 ( .A(n38232), .B(n38231), .Z(n38234) );
  IV U38489 ( .A(n38210), .Z(n38238) );
  AND U38490 ( .A(b[63]), .B(a[123]), .Z(n38237) );
  XOR U38491 ( .A(n38238), .B(n38237), .Z(n38239) );
  XOR U38492 ( .A(n38211), .B(n38239), .Z(n38233) );
  XOR U38493 ( .A(n38234), .B(n38233), .Z(n38226) );
  IV U38494 ( .A(n38211), .Z(n38240) );
  NANDN U38495 ( .A(n38240), .B(n38212), .Z(n38216) );
  NANDN U38496 ( .A(n38214), .B(n38213), .Z(n38215) );
  AND U38497 ( .A(n38216), .B(n38215), .Z(n38225) );
  XOR U38498 ( .A(n38226), .B(n38225), .Z(n38228) );
  XOR U38499 ( .A(n38227), .B(n38228), .Z(n38220) );
  XOR U38500 ( .A(n38219), .B(n38220), .Z(n38222) );
  XNOR U38501 ( .A(n38221), .B(n38222), .Z(n38217) );
  XOR U38502 ( .A(n38218), .B(n38217), .Z(c[251]) );
  AND U38503 ( .A(n38218), .B(n38217), .Z(n38252) );
  NANDN U38504 ( .A(n38220), .B(n38219), .Z(n38224) );
  OR U38505 ( .A(n38222), .B(n38221), .Z(n38223) );
  AND U38506 ( .A(n38224), .B(n38223), .Z(n38255) );
  NANDN U38507 ( .A(n38226), .B(n38225), .Z(n38230) );
  NANDN U38508 ( .A(n38228), .B(n38227), .Z(n38229) );
  AND U38509 ( .A(n38230), .B(n38229), .Z(n38254) );
  NANDN U38510 ( .A(n38232), .B(n38231), .Z(n38236) );
  NAND U38511 ( .A(n38234), .B(n38233), .Z(n38235) );
  AND U38512 ( .A(n38236), .B(n38235), .Z(n38269) );
  NANDN U38513 ( .A(n38238), .B(n38237), .Z(n38242) );
  ANDN U38514 ( .B(n38240), .A(n38239), .Z(n38241) );
  ANDN U38515 ( .B(n38242), .A(n38241), .Z(n38268) );
  NAND U38516 ( .A(n38262), .B(n38243), .Z(n38245) );
  XNOR U38517 ( .A(b[63]), .B(a[126]), .Z(n38263) );
  NANDN U38518 ( .A(n38263), .B(n38264), .Z(n38244) );
  NAND U38519 ( .A(n38245), .B(n38244), .Z(n38260) );
  NAND U38520 ( .A(b[63]), .B(a[124]), .Z(n38275) );
  NANDN U38521 ( .A(n38247), .B(n38246), .Z(n38250) );
  NANDN U38522 ( .A(n38248), .B(b[61]), .Z(n38249) );
  NAND U38523 ( .A(n38250), .B(n38249), .Z(n38259) );
  XOR U38524 ( .A(n38275), .B(n38259), .Z(n38261) );
  XOR U38525 ( .A(n38260), .B(n38261), .Z(n38267) );
  XOR U38526 ( .A(n38268), .B(n38267), .Z(n38270) );
  XNOR U38527 ( .A(n38269), .B(n38270), .Z(n38253) );
  XOR U38528 ( .A(n38254), .B(n38253), .Z(n38256) );
  XNOR U38529 ( .A(n38255), .B(n38256), .Z(n38251) );
  XOR U38530 ( .A(n38252), .B(n38251), .Z(c[252]) );
  AND U38531 ( .A(n38252), .B(n38251), .Z(n38283) );
  NANDN U38532 ( .A(n38254), .B(n38253), .Z(n38258) );
  OR U38533 ( .A(n38256), .B(n38255), .Z(n38257) );
  AND U38534 ( .A(n38258), .B(n38257), .Z(n38293) );
  NANDN U38535 ( .A(n38263), .B(n38262), .Z(n38266) );
  XOR U38536 ( .A(a[127]), .B(b[63]), .Z(n38277) );
  NAND U38537 ( .A(n38264), .B(n38277), .Z(n38265) );
  NAND U38538 ( .A(n38266), .B(n38265), .Z(n38284) );
  AND U38539 ( .A(b[63]), .B(a[125]), .Z(n38274) );
  XOR U38540 ( .A(n38273), .B(n38274), .Z(n38276) );
  XOR U38541 ( .A(n38276), .B(n38275), .Z(n38285) );
  XOR U38542 ( .A(n38284), .B(n38285), .Z(n38287) );
  XOR U38543 ( .A(n38286), .B(n38287), .Z(n38290) );
  NANDN U38544 ( .A(n38268), .B(n38267), .Z(n38272) );
  OR U38545 ( .A(n38270), .B(n38269), .Z(n38271) );
  AND U38546 ( .A(n38272), .B(n38271), .Z(n38291) );
  XOR U38547 ( .A(n38290), .B(n38291), .Z(n38292) );
  XOR U38548 ( .A(n38293), .B(n38292), .Z(n38282) );
  XOR U38549 ( .A(n38283), .B(n38282), .Z(c[253]) );
  AND U38550 ( .A(b[63]), .B(a[126]), .Z(n38297) );
  NANDN U38551 ( .A(n38278), .B(n38277), .Z(n38281) );
  NANDN U38552 ( .A(n38279), .B(b[63]), .Z(n38280) );
  NAND U38553 ( .A(n38281), .B(n38280), .Z(n38298) );
  XNOR U38554 ( .A(n38297), .B(n38298), .Z(n38300) );
  XOR U38555 ( .A(n38299), .B(n38300), .Z(n38303) );
  AND U38556 ( .A(n38283), .B(n38282), .Z(n38302) );
  XNOR U38557 ( .A(n38303), .B(n38302), .Z(n38295) );
  NANDN U38558 ( .A(n38285), .B(n38284), .Z(n38289) );
  NANDN U38559 ( .A(n38287), .B(n38286), .Z(n38288) );
  AND U38560 ( .A(n38289), .B(n38288), .Z(n38304) );
  IV U38561 ( .A(n38305), .Z(n38301) );
  XOR U38562 ( .A(n38304), .B(n38301), .Z(n38294) );
  XNOR U38563 ( .A(n38295), .B(n38294), .Z(c[254]) );
endmodule

