
module Data_Mem ( clk, rst, data_mem_in_wire, data_mem_out_wire, mem_source, 
        addr, data_in, data_out );
  input [2047:0] data_mem_in_wire;
  output [2047:0] data_mem_out_wire;
  input [3:0] mem_source;
  input [31:0] addr;
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst;
  wire   N37, N38, N39, N40, N41, N42, N714, N715, N716, N717, N718, N719,
         N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730,
         N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741,
         N742, N743, N744, N745, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272;
  assign N37 = addr[2];
  assign N38 = addr[3];
  assign N39 = addr[4];
  assign N40 = addr[5];
  assign N41 = addr[6];
  assign N42 = addr[7];

  DFF \memory_reg[0][31]  ( .D(n7761), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[31]), .Q(data_mem_out_wire[31]) );
  DFF \memory_reg[0][30]  ( .D(n7760), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[30]), .Q(data_mem_out_wire[30]) );
  DFF \memory_reg[0][29]  ( .D(n7759), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[29]), .Q(data_mem_out_wire[29]) );
  DFF \memory_reg[0][28]  ( .D(n7758), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[28]), .Q(data_mem_out_wire[28]) );
  DFF \memory_reg[0][27]  ( .D(n7757), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[27]), .Q(data_mem_out_wire[27]) );
  DFF \memory_reg[0][26]  ( .D(n7756), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[26]), .Q(data_mem_out_wire[26]) );
  DFF \memory_reg[0][25]  ( .D(n7755), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[25]), .Q(data_mem_out_wire[25]) );
  DFF \memory_reg[0][24]  ( .D(n7754), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[24]), .Q(data_mem_out_wire[24]) );
  DFF \memory_reg[0][23]  ( .D(n7753), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[23]), .Q(data_mem_out_wire[23]) );
  DFF \memory_reg[0][22]  ( .D(n7752), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[22]), .Q(data_mem_out_wire[22]) );
  DFF \memory_reg[0][21]  ( .D(n7751), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[21]), .Q(data_mem_out_wire[21]) );
  DFF \memory_reg[0][20]  ( .D(n7750), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[20]), .Q(data_mem_out_wire[20]) );
  DFF \memory_reg[0][19]  ( .D(n7749), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[19]), .Q(data_mem_out_wire[19]) );
  DFF \memory_reg[0][18]  ( .D(n7748), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[18]), .Q(data_mem_out_wire[18]) );
  DFF \memory_reg[0][17]  ( .D(n7747), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[17]), .Q(data_mem_out_wire[17]) );
  DFF \memory_reg[0][16]  ( .D(n7746), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[16]), .Q(data_mem_out_wire[16]) );
  DFF \memory_reg[0][15]  ( .D(n7745), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[15]), .Q(data_mem_out_wire[15]) );
  DFF \memory_reg[0][14]  ( .D(n7744), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[14]), .Q(data_mem_out_wire[14]) );
  DFF \memory_reg[0][13]  ( .D(n7743), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[13]), .Q(data_mem_out_wire[13]) );
  DFF \memory_reg[0][12]  ( .D(n7742), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[12]), .Q(data_mem_out_wire[12]) );
  DFF \memory_reg[0][11]  ( .D(n7741), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[11]), .Q(data_mem_out_wire[11]) );
  DFF \memory_reg[0][10]  ( .D(n7740), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[10]), .Q(data_mem_out_wire[10]) );
  DFF \memory_reg[0][9]  ( .D(n7739), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[9]), .Q(data_mem_out_wire[9]) );
  DFF \memory_reg[0][8]  ( .D(n7738), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[8]), .Q(data_mem_out_wire[8]) );
  DFF \memory_reg[0][7]  ( .D(n7737), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[7]), .Q(data_mem_out_wire[7]) );
  DFF \memory_reg[0][6]  ( .D(n7736), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[6]), .Q(data_mem_out_wire[6]) );
  DFF \memory_reg[0][5]  ( .D(n7735), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[5]), .Q(data_mem_out_wire[5]) );
  DFF \memory_reg[0][4]  ( .D(n7734), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[4]), .Q(data_mem_out_wire[4]) );
  DFF \memory_reg[0][3]  ( .D(n7733), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[3]), .Q(data_mem_out_wire[3]) );
  DFF \memory_reg[0][2]  ( .D(n7732), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2]), .Q(data_mem_out_wire[2]) );
  DFF \memory_reg[0][1]  ( .D(n7731), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1]), .Q(data_mem_out_wire[1]) );
  DFF \memory_reg[0][0]  ( .D(n7730), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[0]), .Q(data_mem_out_wire[0]) );
  DFF \memory_reg[1][31]  ( .D(n7729), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[63]), .Q(data_mem_out_wire[63]) );
  DFF \memory_reg[1][30]  ( .D(n7728), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[62]), .Q(data_mem_out_wire[62]) );
  DFF \memory_reg[1][29]  ( .D(n7727), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[61]), .Q(data_mem_out_wire[61]) );
  DFF \memory_reg[1][28]  ( .D(n7726), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[60]), .Q(data_mem_out_wire[60]) );
  DFF \memory_reg[1][27]  ( .D(n7725), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[59]), .Q(data_mem_out_wire[59]) );
  DFF \memory_reg[1][26]  ( .D(n7724), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[58]), .Q(data_mem_out_wire[58]) );
  DFF \memory_reg[1][25]  ( .D(n7723), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[57]), .Q(data_mem_out_wire[57]) );
  DFF \memory_reg[1][24]  ( .D(n7722), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[56]), .Q(data_mem_out_wire[56]) );
  DFF \memory_reg[1][23]  ( .D(n7721), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[55]), .Q(data_mem_out_wire[55]) );
  DFF \memory_reg[1][22]  ( .D(n7720), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[54]), .Q(data_mem_out_wire[54]) );
  DFF \memory_reg[1][21]  ( .D(n7719), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[53]), .Q(data_mem_out_wire[53]) );
  DFF \memory_reg[1][20]  ( .D(n7718), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[52]), .Q(data_mem_out_wire[52]) );
  DFF \memory_reg[1][19]  ( .D(n7717), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[51]), .Q(data_mem_out_wire[51]) );
  DFF \memory_reg[1][18]  ( .D(n7716), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[50]), .Q(data_mem_out_wire[50]) );
  DFF \memory_reg[1][17]  ( .D(n7715), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[49]), .Q(data_mem_out_wire[49]) );
  DFF \memory_reg[1][16]  ( .D(n7714), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[48]), .Q(data_mem_out_wire[48]) );
  DFF \memory_reg[1][15]  ( .D(n7713), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[47]), .Q(data_mem_out_wire[47]) );
  DFF \memory_reg[1][14]  ( .D(n7712), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[46]), .Q(data_mem_out_wire[46]) );
  DFF \memory_reg[1][13]  ( .D(n7711), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[45]), .Q(data_mem_out_wire[45]) );
  DFF \memory_reg[1][12]  ( .D(n7710), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[44]), .Q(data_mem_out_wire[44]) );
  DFF \memory_reg[1][11]  ( .D(n7709), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[43]), .Q(data_mem_out_wire[43]) );
  DFF \memory_reg[1][10]  ( .D(n7708), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[42]), .Q(data_mem_out_wire[42]) );
  DFF \memory_reg[1][9]  ( .D(n7707), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[41]), .Q(data_mem_out_wire[41]) );
  DFF \memory_reg[1][8]  ( .D(n7706), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[40]), .Q(data_mem_out_wire[40]) );
  DFF \memory_reg[1][7]  ( .D(n7705), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[39]), .Q(data_mem_out_wire[39]) );
  DFF \memory_reg[1][6]  ( .D(n7704), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[38]), .Q(data_mem_out_wire[38]) );
  DFF \memory_reg[1][5]  ( .D(n7703), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[37]), .Q(data_mem_out_wire[37]) );
  DFF \memory_reg[1][4]  ( .D(n7702), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[36]), .Q(data_mem_out_wire[36]) );
  DFF \memory_reg[1][3]  ( .D(n7701), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[35]), .Q(data_mem_out_wire[35]) );
  DFF \memory_reg[1][2]  ( .D(n7700), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[34]), .Q(data_mem_out_wire[34]) );
  DFF \memory_reg[1][1]  ( .D(n7699), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[33]), .Q(data_mem_out_wire[33]) );
  DFF \memory_reg[1][0]  ( .D(n7698), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[32]), .Q(data_mem_out_wire[32]) );
  DFF \memory_reg[2][31]  ( .D(n7697), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[95]), .Q(data_mem_out_wire[95]) );
  DFF \memory_reg[2][30]  ( .D(n7696), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[94]), .Q(data_mem_out_wire[94]) );
  DFF \memory_reg[2][29]  ( .D(n7695), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[93]), .Q(data_mem_out_wire[93]) );
  DFF \memory_reg[2][28]  ( .D(n7694), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[92]), .Q(data_mem_out_wire[92]) );
  DFF \memory_reg[2][27]  ( .D(n7693), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[91]), .Q(data_mem_out_wire[91]) );
  DFF \memory_reg[2][26]  ( .D(n7692), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[90]), .Q(data_mem_out_wire[90]) );
  DFF \memory_reg[2][25]  ( .D(n7691), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[89]), .Q(data_mem_out_wire[89]) );
  DFF \memory_reg[2][24]  ( .D(n7690), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[88]), .Q(data_mem_out_wire[88]) );
  DFF \memory_reg[2][23]  ( .D(n7689), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[87]), .Q(data_mem_out_wire[87]) );
  DFF \memory_reg[2][22]  ( .D(n7688), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[86]), .Q(data_mem_out_wire[86]) );
  DFF \memory_reg[2][21]  ( .D(n7687), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[85]), .Q(data_mem_out_wire[85]) );
  DFF \memory_reg[2][20]  ( .D(n7686), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[84]), .Q(data_mem_out_wire[84]) );
  DFF \memory_reg[2][19]  ( .D(n7685), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[83]), .Q(data_mem_out_wire[83]) );
  DFF \memory_reg[2][18]  ( .D(n7684), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[82]), .Q(data_mem_out_wire[82]) );
  DFF \memory_reg[2][17]  ( .D(n7683), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[81]), .Q(data_mem_out_wire[81]) );
  DFF \memory_reg[2][16]  ( .D(n7682), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[80]), .Q(data_mem_out_wire[80]) );
  DFF \memory_reg[2][15]  ( .D(n7681), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[79]), .Q(data_mem_out_wire[79]) );
  DFF \memory_reg[2][14]  ( .D(n7680), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[78]), .Q(data_mem_out_wire[78]) );
  DFF \memory_reg[2][13]  ( .D(n7679), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[77]), .Q(data_mem_out_wire[77]) );
  DFF \memory_reg[2][12]  ( .D(n7678), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[76]), .Q(data_mem_out_wire[76]) );
  DFF \memory_reg[2][11]  ( .D(n7677), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[75]), .Q(data_mem_out_wire[75]) );
  DFF \memory_reg[2][10]  ( .D(n7676), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[74]), .Q(data_mem_out_wire[74]) );
  DFF \memory_reg[2][9]  ( .D(n7675), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[73]), .Q(data_mem_out_wire[73]) );
  DFF \memory_reg[2][8]  ( .D(n7674), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[72]), .Q(data_mem_out_wire[72]) );
  DFF \memory_reg[2][7]  ( .D(n7673), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[71]), .Q(data_mem_out_wire[71]) );
  DFF \memory_reg[2][6]  ( .D(n7672), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[70]), .Q(data_mem_out_wire[70]) );
  DFF \memory_reg[2][5]  ( .D(n7671), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[69]), .Q(data_mem_out_wire[69]) );
  DFF \memory_reg[2][4]  ( .D(n7670), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[68]), .Q(data_mem_out_wire[68]) );
  DFF \memory_reg[2][3]  ( .D(n7669), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[67]), .Q(data_mem_out_wire[67]) );
  DFF \memory_reg[2][2]  ( .D(n7668), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[66]), .Q(data_mem_out_wire[66]) );
  DFF \memory_reg[2][1]  ( .D(n7667), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[65]), .Q(data_mem_out_wire[65]) );
  DFF \memory_reg[2][0]  ( .D(n7666), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[64]), .Q(data_mem_out_wire[64]) );
  DFF \memory_reg[3][31]  ( .D(n7665), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[127]), .Q(data_mem_out_wire[127]) );
  DFF \memory_reg[3][30]  ( .D(n7664), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[126]), .Q(data_mem_out_wire[126]) );
  DFF \memory_reg[3][29]  ( .D(n7663), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[125]), .Q(data_mem_out_wire[125]) );
  DFF \memory_reg[3][28]  ( .D(n7662), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[124]), .Q(data_mem_out_wire[124]) );
  DFF \memory_reg[3][27]  ( .D(n7661), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[123]), .Q(data_mem_out_wire[123]) );
  DFF \memory_reg[3][26]  ( .D(n7660), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[122]), .Q(data_mem_out_wire[122]) );
  DFF \memory_reg[3][25]  ( .D(n7659), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[121]), .Q(data_mem_out_wire[121]) );
  DFF \memory_reg[3][24]  ( .D(n7658), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[120]), .Q(data_mem_out_wire[120]) );
  DFF \memory_reg[3][23]  ( .D(n7657), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[119]), .Q(data_mem_out_wire[119]) );
  DFF \memory_reg[3][22]  ( .D(n7656), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[118]), .Q(data_mem_out_wire[118]) );
  DFF \memory_reg[3][21]  ( .D(n7655), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[117]), .Q(data_mem_out_wire[117]) );
  DFF \memory_reg[3][20]  ( .D(n7654), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[116]), .Q(data_mem_out_wire[116]) );
  DFF \memory_reg[3][19]  ( .D(n7653), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[115]), .Q(data_mem_out_wire[115]) );
  DFF \memory_reg[3][18]  ( .D(n7652), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[114]), .Q(data_mem_out_wire[114]) );
  DFF \memory_reg[3][17]  ( .D(n7651), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[113]), .Q(data_mem_out_wire[113]) );
  DFF \memory_reg[3][16]  ( .D(n7650), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[112]), .Q(data_mem_out_wire[112]) );
  DFF \memory_reg[3][15]  ( .D(n7649), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[111]), .Q(data_mem_out_wire[111]) );
  DFF \memory_reg[3][14]  ( .D(n7648), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[110]), .Q(data_mem_out_wire[110]) );
  DFF \memory_reg[3][13]  ( .D(n7647), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[109]), .Q(data_mem_out_wire[109]) );
  DFF \memory_reg[3][12]  ( .D(n7646), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[108]), .Q(data_mem_out_wire[108]) );
  DFF \memory_reg[3][11]  ( .D(n7645), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[107]), .Q(data_mem_out_wire[107]) );
  DFF \memory_reg[3][10]  ( .D(n7644), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[106]), .Q(data_mem_out_wire[106]) );
  DFF \memory_reg[3][9]  ( .D(n7643), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[105]), .Q(data_mem_out_wire[105]) );
  DFF \memory_reg[3][8]  ( .D(n7642), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[104]), .Q(data_mem_out_wire[104]) );
  DFF \memory_reg[3][7]  ( .D(n7641), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[103]), .Q(data_mem_out_wire[103]) );
  DFF \memory_reg[3][6]  ( .D(n7640), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[102]), .Q(data_mem_out_wire[102]) );
  DFF \memory_reg[3][5]  ( .D(n7639), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[101]), .Q(data_mem_out_wire[101]) );
  DFF \memory_reg[3][4]  ( .D(n7638), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[100]), .Q(data_mem_out_wire[100]) );
  DFF \memory_reg[3][3]  ( .D(n7637), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[99]), .Q(data_mem_out_wire[99]) );
  DFF \memory_reg[3][2]  ( .D(n7636), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[98]), .Q(data_mem_out_wire[98]) );
  DFF \memory_reg[3][1]  ( .D(n7635), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[97]), .Q(data_mem_out_wire[97]) );
  DFF \memory_reg[3][0]  ( .D(n7634), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[96]), .Q(data_mem_out_wire[96]) );
  DFF \memory_reg[4][31]  ( .D(n7633), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[159]), .Q(data_mem_out_wire[159]) );
  DFF \memory_reg[4][30]  ( .D(n7632), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[158]), .Q(data_mem_out_wire[158]) );
  DFF \memory_reg[4][29]  ( .D(n7631), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[157]), .Q(data_mem_out_wire[157]) );
  DFF \memory_reg[4][28]  ( .D(n7630), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[156]), .Q(data_mem_out_wire[156]) );
  DFF \memory_reg[4][27]  ( .D(n7629), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[155]), .Q(data_mem_out_wire[155]) );
  DFF \memory_reg[4][26]  ( .D(n7628), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[154]), .Q(data_mem_out_wire[154]) );
  DFF \memory_reg[4][25]  ( .D(n7627), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[153]), .Q(data_mem_out_wire[153]) );
  DFF \memory_reg[4][24]  ( .D(n7626), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[152]), .Q(data_mem_out_wire[152]) );
  DFF \memory_reg[4][23]  ( .D(n7625), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[151]), .Q(data_mem_out_wire[151]) );
  DFF \memory_reg[4][22]  ( .D(n7624), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[150]), .Q(data_mem_out_wire[150]) );
  DFF \memory_reg[4][21]  ( .D(n7623), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[149]), .Q(data_mem_out_wire[149]) );
  DFF \memory_reg[4][20]  ( .D(n7622), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[148]), .Q(data_mem_out_wire[148]) );
  DFF \memory_reg[4][19]  ( .D(n7621), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[147]), .Q(data_mem_out_wire[147]) );
  DFF \memory_reg[4][18]  ( .D(n7620), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[146]), .Q(data_mem_out_wire[146]) );
  DFF \memory_reg[4][17]  ( .D(n7619), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[145]), .Q(data_mem_out_wire[145]) );
  DFF \memory_reg[4][16]  ( .D(n7618), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[144]), .Q(data_mem_out_wire[144]) );
  DFF \memory_reg[4][15]  ( .D(n7617), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[143]), .Q(data_mem_out_wire[143]) );
  DFF \memory_reg[4][14]  ( .D(n7616), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[142]), .Q(data_mem_out_wire[142]) );
  DFF \memory_reg[4][13]  ( .D(n7615), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[141]), .Q(data_mem_out_wire[141]) );
  DFF \memory_reg[4][12]  ( .D(n7614), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[140]), .Q(data_mem_out_wire[140]) );
  DFF \memory_reg[4][11]  ( .D(n7613), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[139]), .Q(data_mem_out_wire[139]) );
  DFF \memory_reg[4][10]  ( .D(n7612), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[138]), .Q(data_mem_out_wire[138]) );
  DFF \memory_reg[4][9]  ( .D(n7611), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[137]), .Q(data_mem_out_wire[137]) );
  DFF \memory_reg[4][8]  ( .D(n7610), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[136]), .Q(data_mem_out_wire[136]) );
  DFF \memory_reg[4][7]  ( .D(n7609), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[135]), .Q(data_mem_out_wire[135]) );
  DFF \memory_reg[4][6]  ( .D(n7608), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[134]), .Q(data_mem_out_wire[134]) );
  DFF \memory_reg[4][5]  ( .D(n7607), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[133]), .Q(data_mem_out_wire[133]) );
  DFF \memory_reg[4][4]  ( .D(n7606), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[132]), .Q(data_mem_out_wire[132]) );
  DFF \memory_reg[4][3]  ( .D(n7605), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[131]), .Q(data_mem_out_wire[131]) );
  DFF \memory_reg[4][2]  ( .D(n7604), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[130]), .Q(data_mem_out_wire[130]) );
  DFF \memory_reg[4][1]  ( .D(n7603), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[129]), .Q(data_mem_out_wire[129]) );
  DFF \memory_reg[4][0]  ( .D(n7602), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[128]), .Q(data_mem_out_wire[128]) );
  DFF \memory_reg[5][31]  ( .D(n7601), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[191]), .Q(data_mem_out_wire[191]) );
  DFF \memory_reg[5][30]  ( .D(n7600), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[190]), .Q(data_mem_out_wire[190]) );
  DFF \memory_reg[5][29]  ( .D(n7599), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[189]), .Q(data_mem_out_wire[189]) );
  DFF \memory_reg[5][28]  ( .D(n7598), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[188]), .Q(data_mem_out_wire[188]) );
  DFF \memory_reg[5][27]  ( .D(n7597), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[187]), .Q(data_mem_out_wire[187]) );
  DFF \memory_reg[5][26]  ( .D(n7596), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[186]), .Q(data_mem_out_wire[186]) );
  DFF \memory_reg[5][25]  ( .D(n7595), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[185]), .Q(data_mem_out_wire[185]) );
  DFF \memory_reg[5][24]  ( .D(n7594), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[184]), .Q(data_mem_out_wire[184]) );
  DFF \memory_reg[5][23]  ( .D(n7593), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[183]), .Q(data_mem_out_wire[183]) );
  DFF \memory_reg[5][22]  ( .D(n7592), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[182]), .Q(data_mem_out_wire[182]) );
  DFF \memory_reg[5][21]  ( .D(n7591), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[181]), .Q(data_mem_out_wire[181]) );
  DFF \memory_reg[5][20]  ( .D(n7590), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[180]), .Q(data_mem_out_wire[180]) );
  DFF \memory_reg[5][19]  ( .D(n7589), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[179]), .Q(data_mem_out_wire[179]) );
  DFF \memory_reg[5][18]  ( .D(n7588), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[178]), .Q(data_mem_out_wire[178]) );
  DFF \memory_reg[5][17]  ( .D(n7587), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[177]), .Q(data_mem_out_wire[177]) );
  DFF \memory_reg[5][16]  ( .D(n7586), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[176]), .Q(data_mem_out_wire[176]) );
  DFF \memory_reg[5][15]  ( .D(n7585), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[175]), .Q(data_mem_out_wire[175]) );
  DFF \memory_reg[5][14]  ( .D(n7584), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[174]), .Q(data_mem_out_wire[174]) );
  DFF \memory_reg[5][13]  ( .D(n7583), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[173]), .Q(data_mem_out_wire[173]) );
  DFF \memory_reg[5][12]  ( .D(n7582), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[172]), .Q(data_mem_out_wire[172]) );
  DFF \memory_reg[5][11]  ( .D(n7581), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[171]), .Q(data_mem_out_wire[171]) );
  DFF \memory_reg[5][10]  ( .D(n7580), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[170]), .Q(data_mem_out_wire[170]) );
  DFF \memory_reg[5][9]  ( .D(n7579), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[169]), .Q(data_mem_out_wire[169]) );
  DFF \memory_reg[5][8]  ( .D(n7578), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[168]), .Q(data_mem_out_wire[168]) );
  DFF \memory_reg[5][7]  ( .D(n7577), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[167]), .Q(data_mem_out_wire[167]) );
  DFF \memory_reg[5][6]  ( .D(n7576), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[166]), .Q(data_mem_out_wire[166]) );
  DFF \memory_reg[5][5]  ( .D(n7575), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[165]), .Q(data_mem_out_wire[165]) );
  DFF \memory_reg[5][4]  ( .D(n7574), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[164]), .Q(data_mem_out_wire[164]) );
  DFF \memory_reg[5][3]  ( .D(n7573), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[163]), .Q(data_mem_out_wire[163]) );
  DFF \memory_reg[5][2]  ( .D(n7572), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[162]), .Q(data_mem_out_wire[162]) );
  DFF \memory_reg[5][1]  ( .D(n7571), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[161]), .Q(data_mem_out_wire[161]) );
  DFF \memory_reg[5][0]  ( .D(n7570), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[160]), .Q(data_mem_out_wire[160]) );
  DFF \memory_reg[6][31]  ( .D(n7569), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[223]), .Q(data_mem_out_wire[223]) );
  DFF \memory_reg[6][30]  ( .D(n7568), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[222]), .Q(data_mem_out_wire[222]) );
  DFF \memory_reg[6][29]  ( .D(n7567), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[221]), .Q(data_mem_out_wire[221]) );
  DFF \memory_reg[6][28]  ( .D(n7566), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[220]), .Q(data_mem_out_wire[220]) );
  DFF \memory_reg[6][27]  ( .D(n7565), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[219]), .Q(data_mem_out_wire[219]) );
  DFF \memory_reg[6][26]  ( .D(n7564), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[218]), .Q(data_mem_out_wire[218]) );
  DFF \memory_reg[6][25]  ( .D(n7563), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[217]), .Q(data_mem_out_wire[217]) );
  DFF \memory_reg[6][24]  ( .D(n7562), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[216]), .Q(data_mem_out_wire[216]) );
  DFF \memory_reg[6][23]  ( .D(n7561), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[215]), .Q(data_mem_out_wire[215]) );
  DFF \memory_reg[6][22]  ( .D(n7560), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[214]), .Q(data_mem_out_wire[214]) );
  DFF \memory_reg[6][21]  ( .D(n7559), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[213]), .Q(data_mem_out_wire[213]) );
  DFF \memory_reg[6][20]  ( .D(n7558), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[212]), .Q(data_mem_out_wire[212]) );
  DFF \memory_reg[6][19]  ( .D(n7557), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[211]), .Q(data_mem_out_wire[211]) );
  DFF \memory_reg[6][18]  ( .D(n7556), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[210]), .Q(data_mem_out_wire[210]) );
  DFF \memory_reg[6][17]  ( .D(n7555), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[209]), .Q(data_mem_out_wire[209]) );
  DFF \memory_reg[6][16]  ( .D(n7554), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[208]), .Q(data_mem_out_wire[208]) );
  DFF \memory_reg[6][15]  ( .D(n7553), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[207]), .Q(data_mem_out_wire[207]) );
  DFF \memory_reg[6][14]  ( .D(n7552), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[206]), .Q(data_mem_out_wire[206]) );
  DFF \memory_reg[6][13]  ( .D(n7551), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[205]), .Q(data_mem_out_wire[205]) );
  DFF \memory_reg[6][12]  ( .D(n7550), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[204]), .Q(data_mem_out_wire[204]) );
  DFF \memory_reg[6][11]  ( .D(n7549), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[203]), .Q(data_mem_out_wire[203]) );
  DFF \memory_reg[6][10]  ( .D(n7548), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[202]), .Q(data_mem_out_wire[202]) );
  DFF \memory_reg[6][9]  ( .D(n7547), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[201]), .Q(data_mem_out_wire[201]) );
  DFF \memory_reg[6][8]  ( .D(n7546), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[200]), .Q(data_mem_out_wire[200]) );
  DFF \memory_reg[6][7]  ( .D(n7545), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[199]), .Q(data_mem_out_wire[199]) );
  DFF \memory_reg[6][6]  ( .D(n7544), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[198]), .Q(data_mem_out_wire[198]) );
  DFF \memory_reg[6][5]  ( .D(n7543), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[197]), .Q(data_mem_out_wire[197]) );
  DFF \memory_reg[6][4]  ( .D(n7542), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[196]), .Q(data_mem_out_wire[196]) );
  DFF \memory_reg[6][3]  ( .D(n7541), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[195]), .Q(data_mem_out_wire[195]) );
  DFF \memory_reg[6][2]  ( .D(n7540), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[194]), .Q(data_mem_out_wire[194]) );
  DFF \memory_reg[6][1]  ( .D(n7539), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[193]), .Q(data_mem_out_wire[193]) );
  DFF \memory_reg[6][0]  ( .D(n7538), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[192]), .Q(data_mem_out_wire[192]) );
  DFF \memory_reg[7][31]  ( .D(n7537), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[255]), .Q(data_mem_out_wire[255]) );
  DFF \memory_reg[7][30]  ( .D(n7536), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[254]), .Q(data_mem_out_wire[254]) );
  DFF \memory_reg[7][29]  ( .D(n7535), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[253]), .Q(data_mem_out_wire[253]) );
  DFF \memory_reg[7][28]  ( .D(n7534), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[252]), .Q(data_mem_out_wire[252]) );
  DFF \memory_reg[7][27]  ( .D(n7533), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[251]), .Q(data_mem_out_wire[251]) );
  DFF \memory_reg[7][26]  ( .D(n7532), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[250]), .Q(data_mem_out_wire[250]) );
  DFF \memory_reg[7][25]  ( .D(n7531), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[249]), .Q(data_mem_out_wire[249]) );
  DFF \memory_reg[7][24]  ( .D(n7530), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[248]), .Q(data_mem_out_wire[248]) );
  DFF \memory_reg[7][23]  ( .D(n7529), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[247]), .Q(data_mem_out_wire[247]) );
  DFF \memory_reg[7][22]  ( .D(n7528), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[246]), .Q(data_mem_out_wire[246]) );
  DFF \memory_reg[7][21]  ( .D(n7527), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[245]), .Q(data_mem_out_wire[245]) );
  DFF \memory_reg[7][20]  ( .D(n7526), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[244]), .Q(data_mem_out_wire[244]) );
  DFF \memory_reg[7][19]  ( .D(n7525), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[243]), .Q(data_mem_out_wire[243]) );
  DFF \memory_reg[7][18]  ( .D(n7524), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[242]), .Q(data_mem_out_wire[242]) );
  DFF \memory_reg[7][17]  ( .D(n7523), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[241]), .Q(data_mem_out_wire[241]) );
  DFF \memory_reg[7][16]  ( .D(n7522), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[240]), .Q(data_mem_out_wire[240]) );
  DFF \memory_reg[7][15]  ( .D(n7521), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[239]), .Q(data_mem_out_wire[239]) );
  DFF \memory_reg[7][14]  ( .D(n7520), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[238]), .Q(data_mem_out_wire[238]) );
  DFF \memory_reg[7][13]  ( .D(n7519), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[237]), .Q(data_mem_out_wire[237]) );
  DFF \memory_reg[7][12]  ( .D(n7518), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[236]), .Q(data_mem_out_wire[236]) );
  DFF \memory_reg[7][11]  ( .D(n7517), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[235]), .Q(data_mem_out_wire[235]) );
  DFF \memory_reg[7][10]  ( .D(n7516), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[234]), .Q(data_mem_out_wire[234]) );
  DFF \memory_reg[7][9]  ( .D(n7515), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[233]), .Q(data_mem_out_wire[233]) );
  DFF \memory_reg[7][8]  ( .D(n7514), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[232]), .Q(data_mem_out_wire[232]) );
  DFF \memory_reg[7][7]  ( .D(n7513), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[231]), .Q(data_mem_out_wire[231]) );
  DFF \memory_reg[7][6]  ( .D(n7512), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[230]), .Q(data_mem_out_wire[230]) );
  DFF \memory_reg[7][5]  ( .D(n7511), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[229]), .Q(data_mem_out_wire[229]) );
  DFF \memory_reg[7][4]  ( .D(n7510), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[228]), .Q(data_mem_out_wire[228]) );
  DFF \memory_reg[7][3]  ( .D(n7509), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[227]), .Q(data_mem_out_wire[227]) );
  DFF \memory_reg[7][2]  ( .D(n7508), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[226]), .Q(data_mem_out_wire[226]) );
  DFF \memory_reg[7][1]  ( .D(n7507), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[225]), .Q(data_mem_out_wire[225]) );
  DFF \memory_reg[7][0]  ( .D(n7506), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[224]), .Q(data_mem_out_wire[224]) );
  DFF \memory_reg[8][31]  ( .D(n7505), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[287]), .Q(data_mem_out_wire[287]) );
  DFF \memory_reg[8][30]  ( .D(n7504), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[286]), .Q(data_mem_out_wire[286]) );
  DFF \memory_reg[8][29]  ( .D(n7503), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[285]), .Q(data_mem_out_wire[285]) );
  DFF \memory_reg[8][28]  ( .D(n7502), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[284]), .Q(data_mem_out_wire[284]) );
  DFF \memory_reg[8][27]  ( .D(n7501), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[283]), .Q(data_mem_out_wire[283]) );
  DFF \memory_reg[8][26]  ( .D(n7500), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[282]), .Q(data_mem_out_wire[282]) );
  DFF \memory_reg[8][25]  ( .D(n7499), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[281]), .Q(data_mem_out_wire[281]) );
  DFF \memory_reg[8][24]  ( .D(n7498), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[280]), .Q(data_mem_out_wire[280]) );
  DFF \memory_reg[8][23]  ( .D(n7497), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[279]), .Q(data_mem_out_wire[279]) );
  DFF \memory_reg[8][22]  ( .D(n7496), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[278]), .Q(data_mem_out_wire[278]) );
  DFF \memory_reg[8][21]  ( .D(n7495), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[277]), .Q(data_mem_out_wire[277]) );
  DFF \memory_reg[8][20]  ( .D(n7494), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[276]), .Q(data_mem_out_wire[276]) );
  DFF \memory_reg[8][19]  ( .D(n7493), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[275]), .Q(data_mem_out_wire[275]) );
  DFF \memory_reg[8][18]  ( .D(n7492), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[274]), .Q(data_mem_out_wire[274]) );
  DFF \memory_reg[8][17]  ( .D(n7491), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[273]), .Q(data_mem_out_wire[273]) );
  DFF \memory_reg[8][16]  ( .D(n7490), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[272]), .Q(data_mem_out_wire[272]) );
  DFF \memory_reg[8][15]  ( .D(n7489), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[271]), .Q(data_mem_out_wire[271]) );
  DFF \memory_reg[8][14]  ( .D(n7488), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[270]), .Q(data_mem_out_wire[270]) );
  DFF \memory_reg[8][13]  ( .D(n7487), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[269]), .Q(data_mem_out_wire[269]) );
  DFF \memory_reg[8][12]  ( .D(n7486), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[268]), .Q(data_mem_out_wire[268]) );
  DFF \memory_reg[8][11]  ( .D(n7485), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[267]), .Q(data_mem_out_wire[267]) );
  DFF \memory_reg[8][10]  ( .D(n7484), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[266]), .Q(data_mem_out_wire[266]) );
  DFF \memory_reg[8][9]  ( .D(n7483), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[265]), .Q(data_mem_out_wire[265]) );
  DFF \memory_reg[8][8]  ( .D(n7482), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[264]), .Q(data_mem_out_wire[264]) );
  DFF \memory_reg[8][7]  ( .D(n7481), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[263]), .Q(data_mem_out_wire[263]) );
  DFF \memory_reg[8][6]  ( .D(n7480), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[262]), .Q(data_mem_out_wire[262]) );
  DFF \memory_reg[8][5]  ( .D(n7479), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[261]), .Q(data_mem_out_wire[261]) );
  DFF \memory_reg[8][4]  ( .D(n7478), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[260]), .Q(data_mem_out_wire[260]) );
  DFF \memory_reg[8][3]  ( .D(n7477), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[259]), .Q(data_mem_out_wire[259]) );
  DFF \memory_reg[8][2]  ( .D(n7476), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[258]), .Q(data_mem_out_wire[258]) );
  DFF \memory_reg[8][1]  ( .D(n7475), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[257]), .Q(data_mem_out_wire[257]) );
  DFF \memory_reg[8][0]  ( .D(n7474), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[256]), .Q(data_mem_out_wire[256]) );
  DFF \memory_reg[9][31]  ( .D(n7473), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[319]), .Q(data_mem_out_wire[319]) );
  DFF \memory_reg[9][30]  ( .D(n7472), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[318]), .Q(data_mem_out_wire[318]) );
  DFF \memory_reg[9][29]  ( .D(n7471), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[317]), .Q(data_mem_out_wire[317]) );
  DFF \memory_reg[9][28]  ( .D(n7470), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[316]), .Q(data_mem_out_wire[316]) );
  DFF \memory_reg[9][27]  ( .D(n7469), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[315]), .Q(data_mem_out_wire[315]) );
  DFF \memory_reg[9][26]  ( .D(n7468), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[314]), .Q(data_mem_out_wire[314]) );
  DFF \memory_reg[9][25]  ( .D(n7467), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[313]), .Q(data_mem_out_wire[313]) );
  DFF \memory_reg[9][24]  ( .D(n7466), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[312]), .Q(data_mem_out_wire[312]) );
  DFF \memory_reg[9][23]  ( .D(n7465), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[311]), .Q(data_mem_out_wire[311]) );
  DFF \memory_reg[9][22]  ( .D(n7464), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[310]), .Q(data_mem_out_wire[310]) );
  DFF \memory_reg[9][21]  ( .D(n7463), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[309]), .Q(data_mem_out_wire[309]) );
  DFF \memory_reg[9][20]  ( .D(n7462), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[308]), .Q(data_mem_out_wire[308]) );
  DFF \memory_reg[9][19]  ( .D(n7461), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[307]), .Q(data_mem_out_wire[307]) );
  DFF \memory_reg[9][18]  ( .D(n7460), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[306]), .Q(data_mem_out_wire[306]) );
  DFF \memory_reg[9][17]  ( .D(n7459), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[305]), .Q(data_mem_out_wire[305]) );
  DFF \memory_reg[9][16]  ( .D(n7458), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[304]), .Q(data_mem_out_wire[304]) );
  DFF \memory_reg[9][15]  ( .D(n7457), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[303]), .Q(data_mem_out_wire[303]) );
  DFF \memory_reg[9][14]  ( .D(n7456), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[302]), .Q(data_mem_out_wire[302]) );
  DFF \memory_reg[9][13]  ( .D(n7455), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[301]), .Q(data_mem_out_wire[301]) );
  DFF \memory_reg[9][12]  ( .D(n7454), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[300]), .Q(data_mem_out_wire[300]) );
  DFF \memory_reg[9][11]  ( .D(n7453), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[299]), .Q(data_mem_out_wire[299]) );
  DFF \memory_reg[9][10]  ( .D(n7452), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[298]), .Q(data_mem_out_wire[298]) );
  DFF \memory_reg[9][9]  ( .D(n7451), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[297]), .Q(data_mem_out_wire[297]) );
  DFF \memory_reg[9][8]  ( .D(n7450), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[296]), .Q(data_mem_out_wire[296]) );
  DFF \memory_reg[9][7]  ( .D(n7449), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[295]), .Q(data_mem_out_wire[295]) );
  DFF \memory_reg[9][6]  ( .D(n7448), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[294]), .Q(data_mem_out_wire[294]) );
  DFF \memory_reg[9][5]  ( .D(n7447), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[293]), .Q(data_mem_out_wire[293]) );
  DFF \memory_reg[9][4]  ( .D(n7446), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[292]), .Q(data_mem_out_wire[292]) );
  DFF \memory_reg[9][3]  ( .D(n7445), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[291]), .Q(data_mem_out_wire[291]) );
  DFF \memory_reg[9][2]  ( .D(n7444), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[290]), .Q(data_mem_out_wire[290]) );
  DFF \memory_reg[9][1]  ( .D(n7443), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[289]), .Q(data_mem_out_wire[289]) );
  DFF \memory_reg[9][0]  ( .D(n7442), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[288]), .Q(data_mem_out_wire[288]) );
  DFF \memory_reg[10][31]  ( .D(n7441), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[351]), .Q(data_mem_out_wire[351]) );
  DFF \memory_reg[10][30]  ( .D(n7440), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[350]), .Q(data_mem_out_wire[350]) );
  DFF \memory_reg[10][29]  ( .D(n7439), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[349]), .Q(data_mem_out_wire[349]) );
  DFF \memory_reg[10][28]  ( .D(n7438), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[348]), .Q(data_mem_out_wire[348]) );
  DFF \memory_reg[10][27]  ( .D(n7437), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[347]), .Q(data_mem_out_wire[347]) );
  DFF \memory_reg[10][26]  ( .D(n7436), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[346]), .Q(data_mem_out_wire[346]) );
  DFF \memory_reg[10][25]  ( .D(n7435), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[345]), .Q(data_mem_out_wire[345]) );
  DFF \memory_reg[10][24]  ( .D(n7434), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[344]), .Q(data_mem_out_wire[344]) );
  DFF \memory_reg[10][23]  ( .D(n7433), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[343]), .Q(data_mem_out_wire[343]) );
  DFF \memory_reg[10][22]  ( .D(n7432), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[342]), .Q(data_mem_out_wire[342]) );
  DFF \memory_reg[10][21]  ( .D(n7431), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[341]), .Q(data_mem_out_wire[341]) );
  DFF \memory_reg[10][20]  ( .D(n7430), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[340]), .Q(data_mem_out_wire[340]) );
  DFF \memory_reg[10][19]  ( .D(n7429), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[339]), .Q(data_mem_out_wire[339]) );
  DFF \memory_reg[10][18]  ( .D(n7428), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[338]), .Q(data_mem_out_wire[338]) );
  DFF \memory_reg[10][17]  ( .D(n7427), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[337]), .Q(data_mem_out_wire[337]) );
  DFF \memory_reg[10][16]  ( .D(n7426), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[336]), .Q(data_mem_out_wire[336]) );
  DFF \memory_reg[10][15]  ( .D(n7425), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[335]), .Q(data_mem_out_wire[335]) );
  DFF \memory_reg[10][14]  ( .D(n7424), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[334]), .Q(data_mem_out_wire[334]) );
  DFF \memory_reg[10][13]  ( .D(n7423), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[333]), .Q(data_mem_out_wire[333]) );
  DFF \memory_reg[10][12]  ( .D(n7422), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[332]), .Q(data_mem_out_wire[332]) );
  DFF \memory_reg[10][11]  ( .D(n7421), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[331]), .Q(data_mem_out_wire[331]) );
  DFF \memory_reg[10][10]  ( .D(n7420), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[330]), .Q(data_mem_out_wire[330]) );
  DFF \memory_reg[10][9]  ( .D(n7419), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[329]), .Q(data_mem_out_wire[329]) );
  DFF \memory_reg[10][8]  ( .D(n7418), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[328]), .Q(data_mem_out_wire[328]) );
  DFF \memory_reg[10][7]  ( .D(n7417), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[327]), .Q(data_mem_out_wire[327]) );
  DFF \memory_reg[10][6]  ( .D(n7416), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[326]), .Q(data_mem_out_wire[326]) );
  DFF \memory_reg[10][5]  ( .D(n7415), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[325]), .Q(data_mem_out_wire[325]) );
  DFF \memory_reg[10][4]  ( .D(n7414), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[324]), .Q(data_mem_out_wire[324]) );
  DFF \memory_reg[10][3]  ( .D(n7413), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[323]), .Q(data_mem_out_wire[323]) );
  DFF \memory_reg[10][2]  ( .D(n7412), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[322]), .Q(data_mem_out_wire[322]) );
  DFF \memory_reg[10][1]  ( .D(n7411), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[321]), .Q(data_mem_out_wire[321]) );
  DFF \memory_reg[10][0]  ( .D(n7410), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[320]), .Q(data_mem_out_wire[320]) );
  DFF \memory_reg[11][31]  ( .D(n7409), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[383]), .Q(data_mem_out_wire[383]) );
  DFF \memory_reg[11][30]  ( .D(n7408), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[382]), .Q(data_mem_out_wire[382]) );
  DFF \memory_reg[11][29]  ( .D(n7407), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[381]), .Q(data_mem_out_wire[381]) );
  DFF \memory_reg[11][28]  ( .D(n7406), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[380]), .Q(data_mem_out_wire[380]) );
  DFF \memory_reg[11][27]  ( .D(n7405), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[379]), .Q(data_mem_out_wire[379]) );
  DFF \memory_reg[11][26]  ( .D(n7404), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[378]), .Q(data_mem_out_wire[378]) );
  DFF \memory_reg[11][25]  ( .D(n7403), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[377]), .Q(data_mem_out_wire[377]) );
  DFF \memory_reg[11][24]  ( .D(n7402), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[376]), .Q(data_mem_out_wire[376]) );
  DFF \memory_reg[11][23]  ( .D(n7401), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[375]), .Q(data_mem_out_wire[375]) );
  DFF \memory_reg[11][22]  ( .D(n7400), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[374]), .Q(data_mem_out_wire[374]) );
  DFF \memory_reg[11][21]  ( .D(n7399), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[373]), .Q(data_mem_out_wire[373]) );
  DFF \memory_reg[11][20]  ( .D(n7398), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[372]), .Q(data_mem_out_wire[372]) );
  DFF \memory_reg[11][19]  ( .D(n7397), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[371]), .Q(data_mem_out_wire[371]) );
  DFF \memory_reg[11][18]  ( .D(n7396), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[370]), .Q(data_mem_out_wire[370]) );
  DFF \memory_reg[11][17]  ( .D(n7395), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[369]), .Q(data_mem_out_wire[369]) );
  DFF \memory_reg[11][16]  ( .D(n7394), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[368]), .Q(data_mem_out_wire[368]) );
  DFF \memory_reg[11][15]  ( .D(n7393), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[367]), .Q(data_mem_out_wire[367]) );
  DFF \memory_reg[11][14]  ( .D(n7392), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[366]), .Q(data_mem_out_wire[366]) );
  DFF \memory_reg[11][13]  ( .D(n7391), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[365]), .Q(data_mem_out_wire[365]) );
  DFF \memory_reg[11][12]  ( .D(n7390), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[364]), .Q(data_mem_out_wire[364]) );
  DFF \memory_reg[11][11]  ( .D(n7389), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[363]), .Q(data_mem_out_wire[363]) );
  DFF \memory_reg[11][10]  ( .D(n7388), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[362]), .Q(data_mem_out_wire[362]) );
  DFF \memory_reg[11][9]  ( .D(n7387), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[361]), .Q(data_mem_out_wire[361]) );
  DFF \memory_reg[11][8]  ( .D(n7386), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[360]), .Q(data_mem_out_wire[360]) );
  DFF \memory_reg[11][7]  ( .D(n7385), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[359]), .Q(data_mem_out_wire[359]) );
  DFF \memory_reg[11][6]  ( .D(n7384), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[358]), .Q(data_mem_out_wire[358]) );
  DFF \memory_reg[11][5]  ( .D(n7383), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[357]), .Q(data_mem_out_wire[357]) );
  DFF \memory_reg[11][4]  ( .D(n7382), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[356]), .Q(data_mem_out_wire[356]) );
  DFF \memory_reg[11][3]  ( .D(n7381), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[355]), .Q(data_mem_out_wire[355]) );
  DFF \memory_reg[11][2]  ( .D(n7380), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[354]), .Q(data_mem_out_wire[354]) );
  DFF \memory_reg[11][1]  ( .D(n7379), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[353]), .Q(data_mem_out_wire[353]) );
  DFF \memory_reg[11][0]  ( .D(n7378), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[352]), .Q(data_mem_out_wire[352]) );
  DFF \memory_reg[12][31]  ( .D(n7377), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[415]), .Q(data_mem_out_wire[415]) );
  DFF \memory_reg[12][30]  ( .D(n7376), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[414]), .Q(data_mem_out_wire[414]) );
  DFF \memory_reg[12][29]  ( .D(n7375), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[413]), .Q(data_mem_out_wire[413]) );
  DFF \memory_reg[12][28]  ( .D(n7374), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[412]), .Q(data_mem_out_wire[412]) );
  DFF \memory_reg[12][27]  ( .D(n7373), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[411]), .Q(data_mem_out_wire[411]) );
  DFF \memory_reg[12][26]  ( .D(n7372), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[410]), .Q(data_mem_out_wire[410]) );
  DFF \memory_reg[12][25]  ( .D(n7371), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[409]), .Q(data_mem_out_wire[409]) );
  DFF \memory_reg[12][24]  ( .D(n7370), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[408]), .Q(data_mem_out_wire[408]) );
  DFF \memory_reg[12][23]  ( .D(n7369), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[407]), .Q(data_mem_out_wire[407]) );
  DFF \memory_reg[12][22]  ( .D(n7368), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[406]), .Q(data_mem_out_wire[406]) );
  DFF \memory_reg[12][21]  ( .D(n7367), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[405]), .Q(data_mem_out_wire[405]) );
  DFF \memory_reg[12][20]  ( .D(n7366), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[404]), .Q(data_mem_out_wire[404]) );
  DFF \memory_reg[12][19]  ( .D(n7365), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[403]), .Q(data_mem_out_wire[403]) );
  DFF \memory_reg[12][18]  ( .D(n7364), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[402]), .Q(data_mem_out_wire[402]) );
  DFF \memory_reg[12][17]  ( .D(n7363), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[401]), .Q(data_mem_out_wire[401]) );
  DFF \memory_reg[12][16]  ( .D(n7362), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[400]), .Q(data_mem_out_wire[400]) );
  DFF \memory_reg[12][15]  ( .D(n7361), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[399]), .Q(data_mem_out_wire[399]) );
  DFF \memory_reg[12][14]  ( .D(n7360), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[398]), .Q(data_mem_out_wire[398]) );
  DFF \memory_reg[12][13]  ( .D(n7359), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[397]), .Q(data_mem_out_wire[397]) );
  DFF \memory_reg[12][12]  ( .D(n7358), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[396]), .Q(data_mem_out_wire[396]) );
  DFF \memory_reg[12][11]  ( .D(n7357), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[395]), .Q(data_mem_out_wire[395]) );
  DFF \memory_reg[12][10]  ( .D(n7356), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[394]), .Q(data_mem_out_wire[394]) );
  DFF \memory_reg[12][9]  ( .D(n7355), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[393]), .Q(data_mem_out_wire[393]) );
  DFF \memory_reg[12][8]  ( .D(n7354), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[392]), .Q(data_mem_out_wire[392]) );
  DFF \memory_reg[12][7]  ( .D(n7353), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[391]), .Q(data_mem_out_wire[391]) );
  DFF \memory_reg[12][6]  ( .D(n7352), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[390]), .Q(data_mem_out_wire[390]) );
  DFF \memory_reg[12][5]  ( .D(n7351), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[389]), .Q(data_mem_out_wire[389]) );
  DFF \memory_reg[12][4]  ( .D(n7350), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[388]), .Q(data_mem_out_wire[388]) );
  DFF \memory_reg[12][3]  ( .D(n7349), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[387]), .Q(data_mem_out_wire[387]) );
  DFF \memory_reg[12][2]  ( .D(n7348), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[386]), .Q(data_mem_out_wire[386]) );
  DFF \memory_reg[12][1]  ( .D(n7347), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[385]), .Q(data_mem_out_wire[385]) );
  DFF \memory_reg[12][0]  ( .D(n7346), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[384]), .Q(data_mem_out_wire[384]) );
  DFF \memory_reg[13][31]  ( .D(n7345), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[447]), .Q(data_mem_out_wire[447]) );
  DFF \memory_reg[13][30]  ( .D(n7344), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[446]), .Q(data_mem_out_wire[446]) );
  DFF \memory_reg[13][29]  ( .D(n7343), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[445]), .Q(data_mem_out_wire[445]) );
  DFF \memory_reg[13][28]  ( .D(n7342), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[444]), .Q(data_mem_out_wire[444]) );
  DFF \memory_reg[13][27]  ( .D(n7341), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[443]), .Q(data_mem_out_wire[443]) );
  DFF \memory_reg[13][26]  ( .D(n7340), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[442]), .Q(data_mem_out_wire[442]) );
  DFF \memory_reg[13][25]  ( .D(n7339), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[441]), .Q(data_mem_out_wire[441]) );
  DFF \memory_reg[13][24]  ( .D(n7338), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[440]), .Q(data_mem_out_wire[440]) );
  DFF \memory_reg[13][23]  ( .D(n7337), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[439]), .Q(data_mem_out_wire[439]) );
  DFF \memory_reg[13][22]  ( .D(n7336), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[438]), .Q(data_mem_out_wire[438]) );
  DFF \memory_reg[13][21]  ( .D(n7335), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[437]), .Q(data_mem_out_wire[437]) );
  DFF \memory_reg[13][20]  ( .D(n7334), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[436]), .Q(data_mem_out_wire[436]) );
  DFF \memory_reg[13][19]  ( .D(n7333), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[435]), .Q(data_mem_out_wire[435]) );
  DFF \memory_reg[13][18]  ( .D(n7332), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[434]), .Q(data_mem_out_wire[434]) );
  DFF \memory_reg[13][17]  ( .D(n7331), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[433]), .Q(data_mem_out_wire[433]) );
  DFF \memory_reg[13][16]  ( .D(n7330), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[432]), .Q(data_mem_out_wire[432]) );
  DFF \memory_reg[13][15]  ( .D(n7329), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[431]), .Q(data_mem_out_wire[431]) );
  DFF \memory_reg[13][14]  ( .D(n7328), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[430]), .Q(data_mem_out_wire[430]) );
  DFF \memory_reg[13][13]  ( .D(n7327), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[429]), .Q(data_mem_out_wire[429]) );
  DFF \memory_reg[13][12]  ( .D(n7326), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[428]), .Q(data_mem_out_wire[428]) );
  DFF \memory_reg[13][11]  ( .D(n7325), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[427]), .Q(data_mem_out_wire[427]) );
  DFF \memory_reg[13][10]  ( .D(n7324), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[426]), .Q(data_mem_out_wire[426]) );
  DFF \memory_reg[13][9]  ( .D(n7323), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[425]), .Q(data_mem_out_wire[425]) );
  DFF \memory_reg[13][8]  ( .D(n7322), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[424]), .Q(data_mem_out_wire[424]) );
  DFF \memory_reg[13][7]  ( .D(n7321), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[423]), .Q(data_mem_out_wire[423]) );
  DFF \memory_reg[13][6]  ( .D(n7320), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[422]), .Q(data_mem_out_wire[422]) );
  DFF \memory_reg[13][5]  ( .D(n7319), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[421]), .Q(data_mem_out_wire[421]) );
  DFF \memory_reg[13][4]  ( .D(n7318), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[420]), .Q(data_mem_out_wire[420]) );
  DFF \memory_reg[13][3]  ( .D(n7317), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[419]), .Q(data_mem_out_wire[419]) );
  DFF \memory_reg[13][2]  ( .D(n7316), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[418]), .Q(data_mem_out_wire[418]) );
  DFF \memory_reg[13][1]  ( .D(n7315), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[417]), .Q(data_mem_out_wire[417]) );
  DFF \memory_reg[13][0]  ( .D(n7314), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[416]), .Q(data_mem_out_wire[416]) );
  DFF \memory_reg[14][31]  ( .D(n7313), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[479]), .Q(data_mem_out_wire[479]) );
  DFF \memory_reg[14][30]  ( .D(n7312), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[478]), .Q(data_mem_out_wire[478]) );
  DFF \memory_reg[14][29]  ( .D(n7311), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[477]), .Q(data_mem_out_wire[477]) );
  DFF \memory_reg[14][28]  ( .D(n7310), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[476]), .Q(data_mem_out_wire[476]) );
  DFF \memory_reg[14][27]  ( .D(n7309), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[475]), .Q(data_mem_out_wire[475]) );
  DFF \memory_reg[14][26]  ( .D(n7308), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[474]), .Q(data_mem_out_wire[474]) );
  DFF \memory_reg[14][25]  ( .D(n7307), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[473]), .Q(data_mem_out_wire[473]) );
  DFF \memory_reg[14][24]  ( .D(n7306), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[472]), .Q(data_mem_out_wire[472]) );
  DFF \memory_reg[14][23]  ( .D(n7305), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[471]), .Q(data_mem_out_wire[471]) );
  DFF \memory_reg[14][22]  ( .D(n7304), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[470]), .Q(data_mem_out_wire[470]) );
  DFF \memory_reg[14][21]  ( .D(n7303), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[469]), .Q(data_mem_out_wire[469]) );
  DFF \memory_reg[14][20]  ( .D(n7302), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[468]), .Q(data_mem_out_wire[468]) );
  DFF \memory_reg[14][19]  ( .D(n7301), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[467]), .Q(data_mem_out_wire[467]) );
  DFF \memory_reg[14][18]  ( .D(n7300), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[466]), .Q(data_mem_out_wire[466]) );
  DFF \memory_reg[14][17]  ( .D(n7299), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[465]), .Q(data_mem_out_wire[465]) );
  DFF \memory_reg[14][16]  ( .D(n7298), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[464]), .Q(data_mem_out_wire[464]) );
  DFF \memory_reg[14][15]  ( .D(n7297), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[463]), .Q(data_mem_out_wire[463]) );
  DFF \memory_reg[14][14]  ( .D(n7296), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[462]), .Q(data_mem_out_wire[462]) );
  DFF \memory_reg[14][13]  ( .D(n7295), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[461]), .Q(data_mem_out_wire[461]) );
  DFF \memory_reg[14][12]  ( .D(n7294), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[460]), .Q(data_mem_out_wire[460]) );
  DFF \memory_reg[14][11]  ( .D(n7293), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[459]), .Q(data_mem_out_wire[459]) );
  DFF \memory_reg[14][10]  ( .D(n7292), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[458]), .Q(data_mem_out_wire[458]) );
  DFF \memory_reg[14][9]  ( .D(n7291), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[457]), .Q(data_mem_out_wire[457]) );
  DFF \memory_reg[14][8]  ( .D(n7290), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[456]), .Q(data_mem_out_wire[456]) );
  DFF \memory_reg[14][7]  ( .D(n7289), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[455]), .Q(data_mem_out_wire[455]) );
  DFF \memory_reg[14][6]  ( .D(n7288), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[454]), .Q(data_mem_out_wire[454]) );
  DFF \memory_reg[14][5]  ( .D(n7287), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[453]), .Q(data_mem_out_wire[453]) );
  DFF \memory_reg[14][4]  ( .D(n7286), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[452]), .Q(data_mem_out_wire[452]) );
  DFF \memory_reg[14][3]  ( .D(n7285), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[451]), .Q(data_mem_out_wire[451]) );
  DFF \memory_reg[14][2]  ( .D(n7284), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[450]), .Q(data_mem_out_wire[450]) );
  DFF \memory_reg[14][1]  ( .D(n7283), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[449]), .Q(data_mem_out_wire[449]) );
  DFF \memory_reg[14][0]  ( .D(n7282), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[448]), .Q(data_mem_out_wire[448]) );
  DFF \memory_reg[15][31]  ( .D(n7281), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[511]), .Q(data_mem_out_wire[511]) );
  DFF \memory_reg[15][30]  ( .D(n7280), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[510]), .Q(data_mem_out_wire[510]) );
  DFF \memory_reg[15][29]  ( .D(n7279), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[509]), .Q(data_mem_out_wire[509]) );
  DFF \memory_reg[15][28]  ( .D(n7278), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[508]), .Q(data_mem_out_wire[508]) );
  DFF \memory_reg[15][27]  ( .D(n7277), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[507]), .Q(data_mem_out_wire[507]) );
  DFF \memory_reg[15][26]  ( .D(n7276), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[506]), .Q(data_mem_out_wire[506]) );
  DFF \memory_reg[15][25]  ( .D(n7275), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[505]), .Q(data_mem_out_wire[505]) );
  DFF \memory_reg[15][24]  ( .D(n7274), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[504]), .Q(data_mem_out_wire[504]) );
  DFF \memory_reg[15][23]  ( .D(n7273), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[503]), .Q(data_mem_out_wire[503]) );
  DFF \memory_reg[15][22]  ( .D(n7272), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[502]), .Q(data_mem_out_wire[502]) );
  DFF \memory_reg[15][21]  ( .D(n7271), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[501]), .Q(data_mem_out_wire[501]) );
  DFF \memory_reg[15][20]  ( .D(n7270), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[500]), .Q(data_mem_out_wire[500]) );
  DFF \memory_reg[15][19]  ( .D(n7269), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[499]), .Q(data_mem_out_wire[499]) );
  DFF \memory_reg[15][18]  ( .D(n7268), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[498]), .Q(data_mem_out_wire[498]) );
  DFF \memory_reg[15][17]  ( .D(n7267), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[497]), .Q(data_mem_out_wire[497]) );
  DFF \memory_reg[15][16]  ( .D(n7266), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[496]), .Q(data_mem_out_wire[496]) );
  DFF \memory_reg[15][15]  ( .D(n7265), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[495]), .Q(data_mem_out_wire[495]) );
  DFF \memory_reg[15][14]  ( .D(n7264), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[494]), .Q(data_mem_out_wire[494]) );
  DFF \memory_reg[15][13]  ( .D(n7263), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[493]), .Q(data_mem_out_wire[493]) );
  DFF \memory_reg[15][12]  ( .D(n7262), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[492]), .Q(data_mem_out_wire[492]) );
  DFF \memory_reg[15][11]  ( .D(n7261), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[491]), .Q(data_mem_out_wire[491]) );
  DFF \memory_reg[15][10]  ( .D(n7260), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[490]), .Q(data_mem_out_wire[490]) );
  DFF \memory_reg[15][9]  ( .D(n7259), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[489]), .Q(data_mem_out_wire[489]) );
  DFF \memory_reg[15][8]  ( .D(n7258), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[488]), .Q(data_mem_out_wire[488]) );
  DFF \memory_reg[15][7]  ( .D(n7257), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[487]), .Q(data_mem_out_wire[487]) );
  DFF \memory_reg[15][6]  ( .D(n7256), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[486]), .Q(data_mem_out_wire[486]) );
  DFF \memory_reg[15][5]  ( .D(n7255), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[485]), .Q(data_mem_out_wire[485]) );
  DFF \memory_reg[15][4]  ( .D(n7254), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[484]), .Q(data_mem_out_wire[484]) );
  DFF \memory_reg[15][3]  ( .D(n7253), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[483]), .Q(data_mem_out_wire[483]) );
  DFF \memory_reg[15][2]  ( .D(n7252), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[482]), .Q(data_mem_out_wire[482]) );
  DFF \memory_reg[15][1]  ( .D(n7251), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[481]), .Q(data_mem_out_wire[481]) );
  DFF \memory_reg[15][0]  ( .D(n7250), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[480]), .Q(data_mem_out_wire[480]) );
  DFF \memory_reg[16][31]  ( .D(n7249), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[543]), .Q(data_mem_out_wire[543]) );
  DFF \memory_reg[16][30]  ( .D(n7248), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[542]), .Q(data_mem_out_wire[542]) );
  DFF \memory_reg[16][29]  ( .D(n7247), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[541]), .Q(data_mem_out_wire[541]) );
  DFF \memory_reg[16][28]  ( .D(n7246), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[540]), .Q(data_mem_out_wire[540]) );
  DFF \memory_reg[16][27]  ( .D(n7245), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[539]), .Q(data_mem_out_wire[539]) );
  DFF \memory_reg[16][26]  ( .D(n7244), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[538]), .Q(data_mem_out_wire[538]) );
  DFF \memory_reg[16][25]  ( .D(n7243), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[537]), .Q(data_mem_out_wire[537]) );
  DFF \memory_reg[16][24]  ( .D(n7242), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[536]), .Q(data_mem_out_wire[536]) );
  DFF \memory_reg[16][23]  ( .D(n7241), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[535]), .Q(data_mem_out_wire[535]) );
  DFF \memory_reg[16][22]  ( .D(n7240), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[534]), .Q(data_mem_out_wire[534]) );
  DFF \memory_reg[16][21]  ( .D(n7239), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[533]), .Q(data_mem_out_wire[533]) );
  DFF \memory_reg[16][20]  ( .D(n7238), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[532]), .Q(data_mem_out_wire[532]) );
  DFF \memory_reg[16][19]  ( .D(n7237), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[531]), .Q(data_mem_out_wire[531]) );
  DFF \memory_reg[16][18]  ( .D(n7236), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[530]), .Q(data_mem_out_wire[530]) );
  DFF \memory_reg[16][17]  ( .D(n7235), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[529]), .Q(data_mem_out_wire[529]) );
  DFF \memory_reg[16][16]  ( .D(n7234), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[528]), .Q(data_mem_out_wire[528]) );
  DFF \memory_reg[16][15]  ( .D(n7233), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[527]), .Q(data_mem_out_wire[527]) );
  DFF \memory_reg[16][14]  ( .D(n7232), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[526]), .Q(data_mem_out_wire[526]) );
  DFF \memory_reg[16][13]  ( .D(n7231), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[525]), .Q(data_mem_out_wire[525]) );
  DFF \memory_reg[16][12]  ( .D(n7230), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[524]), .Q(data_mem_out_wire[524]) );
  DFF \memory_reg[16][11]  ( .D(n7229), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[523]), .Q(data_mem_out_wire[523]) );
  DFF \memory_reg[16][10]  ( .D(n7228), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[522]), .Q(data_mem_out_wire[522]) );
  DFF \memory_reg[16][9]  ( .D(n7227), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[521]), .Q(data_mem_out_wire[521]) );
  DFF \memory_reg[16][8]  ( .D(n7226), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[520]), .Q(data_mem_out_wire[520]) );
  DFF \memory_reg[16][7]  ( .D(n7225), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[519]), .Q(data_mem_out_wire[519]) );
  DFF \memory_reg[16][6]  ( .D(n7224), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[518]), .Q(data_mem_out_wire[518]) );
  DFF \memory_reg[16][5]  ( .D(n7223), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[517]), .Q(data_mem_out_wire[517]) );
  DFF \memory_reg[16][4]  ( .D(n7222), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[516]), .Q(data_mem_out_wire[516]) );
  DFF \memory_reg[16][3]  ( .D(n7221), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[515]), .Q(data_mem_out_wire[515]) );
  DFF \memory_reg[16][2]  ( .D(n7220), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[514]), .Q(data_mem_out_wire[514]) );
  DFF \memory_reg[16][1]  ( .D(n7219), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[513]), .Q(data_mem_out_wire[513]) );
  DFF \memory_reg[16][0]  ( .D(n7218), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[512]), .Q(data_mem_out_wire[512]) );
  DFF \memory_reg[17][31]  ( .D(n7217), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[575]), .Q(data_mem_out_wire[575]) );
  DFF \memory_reg[17][30]  ( .D(n7216), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[574]), .Q(data_mem_out_wire[574]) );
  DFF \memory_reg[17][29]  ( .D(n7215), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[573]), .Q(data_mem_out_wire[573]) );
  DFF \memory_reg[17][28]  ( .D(n7214), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[572]), .Q(data_mem_out_wire[572]) );
  DFF \memory_reg[17][27]  ( .D(n7213), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[571]), .Q(data_mem_out_wire[571]) );
  DFF \memory_reg[17][26]  ( .D(n7212), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[570]), .Q(data_mem_out_wire[570]) );
  DFF \memory_reg[17][25]  ( .D(n7211), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[569]), .Q(data_mem_out_wire[569]) );
  DFF \memory_reg[17][24]  ( .D(n7210), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[568]), .Q(data_mem_out_wire[568]) );
  DFF \memory_reg[17][23]  ( .D(n7209), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[567]), .Q(data_mem_out_wire[567]) );
  DFF \memory_reg[17][22]  ( .D(n7208), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[566]), .Q(data_mem_out_wire[566]) );
  DFF \memory_reg[17][21]  ( .D(n7207), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[565]), .Q(data_mem_out_wire[565]) );
  DFF \memory_reg[17][20]  ( .D(n7206), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[564]), .Q(data_mem_out_wire[564]) );
  DFF \memory_reg[17][19]  ( .D(n7205), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[563]), .Q(data_mem_out_wire[563]) );
  DFF \memory_reg[17][18]  ( .D(n7204), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[562]), .Q(data_mem_out_wire[562]) );
  DFF \memory_reg[17][17]  ( .D(n7203), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[561]), .Q(data_mem_out_wire[561]) );
  DFF \memory_reg[17][16]  ( .D(n7202), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[560]), .Q(data_mem_out_wire[560]) );
  DFF \memory_reg[17][15]  ( .D(n7201), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[559]), .Q(data_mem_out_wire[559]) );
  DFF \memory_reg[17][14]  ( .D(n7200), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[558]), .Q(data_mem_out_wire[558]) );
  DFF \memory_reg[17][13]  ( .D(n7199), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[557]), .Q(data_mem_out_wire[557]) );
  DFF \memory_reg[17][12]  ( .D(n7198), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[556]), .Q(data_mem_out_wire[556]) );
  DFF \memory_reg[17][11]  ( .D(n7197), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[555]), .Q(data_mem_out_wire[555]) );
  DFF \memory_reg[17][10]  ( .D(n7196), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[554]), .Q(data_mem_out_wire[554]) );
  DFF \memory_reg[17][9]  ( .D(n7195), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[553]), .Q(data_mem_out_wire[553]) );
  DFF \memory_reg[17][8]  ( .D(n7194), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[552]), .Q(data_mem_out_wire[552]) );
  DFF \memory_reg[17][7]  ( .D(n7193), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[551]), .Q(data_mem_out_wire[551]) );
  DFF \memory_reg[17][6]  ( .D(n7192), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[550]), .Q(data_mem_out_wire[550]) );
  DFF \memory_reg[17][5]  ( .D(n7191), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[549]), .Q(data_mem_out_wire[549]) );
  DFF \memory_reg[17][4]  ( .D(n7190), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[548]), .Q(data_mem_out_wire[548]) );
  DFF \memory_reg[17][3]  ( .D(n7189), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[547]), .Q(data_mem_out_wire[547]) );
  DFF \memory_reg[17][2]  ( .D(n7188), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[546]), .Q(data_mem_out_wire[546]) );
  DFF \memory_reg[17][1]  ( .D(n7187), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[545]), .Q(data_mem_out_wire[545]) );
  DFF \memory_reg[17][0]  ( .D(n7186), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[544]), .Q(data_mem_out_wire[544]) );
  DFF \memory_reg[18][31]  ( .D(n7185), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[607]), .Q(data_mem_out_wire[607]) );
  DFF \memory_reg[18][30]  ( .D(n7184), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[606]), .Q(data_mem_out_wire[606]) );
  DFF \memory_reg[18][29]  ( .D(n7183), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[605]), .Q(data_mem_out_wire[605]) );
  DFF \memory_reg[18][28]  ( .D(n7182), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[604]), .Q(data_mem_out_wire[604]) );
  DFF \memory_reg[18][27]  ( .D(n7181), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[603]), .Q(data_mem_out_wire[603]) );
  DFF \memory_reg[18][26]  ( .D(n7180), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[602]), .Q(data_mem_out_wire[602]) );
  DFF \memory_reg[18][25]  ( .D(n7179), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[601]), .Q(data_mem_out_wire[601]) );
  DFF \memory_reg[18][24]  ( .D(n7178), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[600]), .Q(data_mem_out_wire[600]) );
  DFF \memory_reg[18][23]  ( .D(n7177), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[599]), .Q(data_mem_out_wire[599]) );
  DFF \memory_reg[18][22]  ( .D(n7176), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[598]), .Q(data_mem_out_wire[598]) );
  DFF \memory_reg[18][21]  ( .D(n7175), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[597]), .Q(data_mem_out_wire[597]) );
  DFF \memory_reg[18][20]  ( .D(n7174), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[596]), .Q(data_mem_out_wire[596]) );
  DFF \memory_reg[18][19]  ( .D(n7173), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[595]), .Q(data_mem_out_wire[595]) );
  DFF \memory_reg[18][18]  ( .D(n7172), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[594]), .Q(data_mem_out_wire[594]) );
  DFF \memory_reg[18][17]  ( .D(n7171), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[593]), .Q(data_mem_out_wire[593]) );
  DFF \memory_reg[18][16]  ( .D(n7170), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[592]), .Q(data_mem_out_wire[592]) );
  DFF \memory_reg[18][15]  ( .D(n7169), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[591]), .Q(data_mem_out_wire[591]) );
  DFF \memory_reg[18][14]  ( .D(n7168), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[590]), .Q(data_mem_out_wire[590]) );
  DFF \memory_reg[18][13]  ( .D(n7167), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[589]), .Q(data_mem_out_wire[589]) );
  DFF \memory_reg[18][12]  ( .D(n7166), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[588]), .Q(data_mem_out_wire[588]) );
  DFF \memory_reg[18][11]  ( .D(n7165), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[587]), .Q(data_mem_out_wire[587]) );
  DFF \memory_reg[18][10]  ( .D(n7164), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[586]), .Q(data_mem_out_wire[586]) );
  DFF \memory_reg[18][9]  ( .D(n7163), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[585]), .Q(data_mem_out_wire[585]) );
  DFF \memory_reg[18][8]  ( .D(n7162), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[584]), .Q(data_mem_out_wire[584]) );
  DFF \memory_reg[18][7]  ( .D(n7161), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[583]), .Q(data_mem_out_wire[583]) );
  DFF \memory_reg[18][6]  ( .D(n7160), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[582]), .Q(data_mem_out_wire[582]) );
  DFF \memory_reg[18][5]  ( .D(n7159), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[581]), .Q(data_mem_out_wire[581]) );
  DFF \memory_reg[18][4]  ( .D(n7158), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[580]), .Q(data_mem_out_wire[580]) );
  DFF \memory_reg[18][3]  ( .D(n7157), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[579]), .Q(data_mem_out_wire[579]) );
  DFF \memory_reg[18][2]  ( .D(n7156), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[578]), .Q(data_mem_out_wire[578]) );
  DFF \memory_reg[18][1]  ( .D(n7155), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[577]), .Q(data_mem_out_wire[577]) );
  DFF \memory_reg[18][0]  ( .D(n7154), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[576]), .Q(data_mem_out_wire[576]) );
  DFF \memory_reg[19][31]  ( .D(n7153), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[639]), .Q(data_mem_out_wire[639]) );
  DFF \memory_reg[19][30]  ( .D(n7152), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[638]), .Q(data_mem_out_wire[638]) );
  DFF \memory_reg[19][29]  ( .D(n7151), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[637]), .Q(data_mem_out_wire[637]) );
  DFF \memory_reg[19][28]  ( .D(n7150), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[636]), .Q(data_mem_out_wire[636]) );
  DFF \memory_reg[19][27]  ( .D(n7149), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[635]), .Q(data_mem_out_wire[635]) );
  DFF \memory_reg[19][26]  ( .D(n7148), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[634]), .Q(data_mem_out_wire[634]) );
  DFF \memory_reg[19][25]  ( .D(n7147), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[633]), .Q(data_mem_out_wire[633]) );
  DFF \memory_reg[19][24]  ( .D(n7146), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[632]), .Q(data_mem_out_wire[632]) );
  DFF \memory_reg[19][23]  ( .D(n7145), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[631]), .Q(data_mem_out_wire[631]) );
  DFF \memory_reg[19][22]  ( .D(n7144), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[630]), .Q(data_mem_out_wire[630]) );
  DFF \memory_reg[19][21]  ( .D(n7143), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[629]), .Q(data_mem_out_wire[629]) );
  DFF \memory_reg[19][20]  ( .D(n7142), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[628]), .Q(data_mem_out_wire[628]) );
  DFF \memory_reg[19][19]  ( .D(n7141), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[627]), .Q(data_mem_out_wire[627]) );
  DFF \memory_reg[19][18]  ( .D(n7140), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[626]), .Q(data_mem_out_wire[626]) );
  DFF \memory_reg[19][17]  ( .D(n7139), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[625]), .Q(data_mem_out_wire[625]) );
  DFF \memory_reg[19][16]  ( .D(n7138), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[624]), .Q(data_mem_out_wire[624]) );
  DFF \memory_reg[19][15]  ( .D(n7137), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[623]), .Q(data_mem_out_wire[623]) );
  DFF \memory_reg[19][14]  ( .D(n7136), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[622]), .Q(data_mem_out_wire[622]) );
  DFF \memory_reg[19][13]  ( .D(n7135), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[621]), .Q(data_mem_out_wire[621]) );
  DFF \memory_reg[19][12]  ( .D(n7134), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[620]), .Q(data_mem_out_wire[620]) );
  DFF \memory_reg[19][11]  ( .D(n7133), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[619]), .Q(data_mem_out_wire[619]) );
  DFF \memory_reg[19][10]  ( .D(n7132), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[618]), .Q(data_mem_out_wire[618]) );
  DFF \memory_reg[19][9]  ( .D(n7131), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[617]), .Q(data_mem_out_wire[617]) );
  DFF \memory_reg[19][8]  ( .D(n7130), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[616]), .Q(data_mem_out_wire[616]) );
  DFF \memory_reg[19][7]  ( .D(n7129), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[615]), .Q(data_mem_out_wire[615]) );
  DFF \memory_reg[19][6]  ( .D(n7128), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[614]), .Q(data_mem_out_wire[614]) );
  DFF \memory_reg[19][5]  ( .D(n7127), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[613]), .Q(data_mem_out_wire[613]) );
  DFF \memory_reg[19][4]  ( .D(n7126), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[612]), .Q(data_mem_out_wire[612]) );
  DFF \memory_reg[19][3]  ( .D(n7125), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[611]), .Q(data_mem_out_wire[611]) );
  DFF \memory_reg[19][2]  ( .D(n7124), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[610]), .Q(data_mem_out_wire[610]) );
  DFF \memory_reg[19][1]  ( .D(n7123), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[609]), .Q(data_mem_out_wire[609]) );
  DFF \memory_reg[19][0]  ( .D(n7122), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[608]), .Q(data_mem_out_wire[608]) );
  DFF \memory_reg[20][31]  ( .D(n7121), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[671]), .Q(data_mem_out_wire[671]) );
  DFF \memory_reg[20][30]  ( .D(n7120), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[670]), .Q(data_mem_out_wire[670]) );
  DFF \memory_reg[20][29]  ( .D(n7119), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[669]), .Q(data_mem_out_wire[669]) );
  DFF \memory_reg[20][28]  ( .D(n7118), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[668]), .Q(data_mem_out_wire[668]) );
  DFF \memory_reg[20][27]  ( .D(n7117), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[667]), .Q(data_mem_out_wire[667]) );
  DFF \memory_reg[20][26]  ( .D(n7116), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[666]), .Q(data_mem_out_wire[666]) );
  DFF \memory_reg[20][25]  ( .D(n7115), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[665]), .Q(data_mem_out_wire[665]) );
  DFF \memory_reg[20][24]  ( .D(n7114), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[664]), .Q(data_mem_out_wire[664]) );
  DFF \memory_reg[20][23]  ( .D(n7113), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[663]), .Q(data_mem_out_wire[663]) );
  DFF \memory_reg[20][22]  ( .D(n7112), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[662]), .Q(data_mem_out_wire[662]) );
  DFF \memory_reg[20][21]  ( .D(n7111), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[661]), .Q(data_mem_out_wire[661]) );
  DFF \memory_reg[20][20]  ( .D(n7110), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[660]), .Q(data_mem_out_wire[660]) );
  DFF \memory_reg[20][19]  ( .D(n7109), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[659]), .Q(data_mem_out_wire[659]) );
  DFF \memory_reg[20][18]  ( .D(n7108), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[658]), .Q(data_mem_out_wire[658]) );
  DFF \memory_reg[20][17]  ( .D(n7107), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[657]), .Q(data_mem_out_wire[657]) );
  DFF \memory_reg[20][16]  ( .D(n7106), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[656]), .Q(data_mem_out_wire[656]) );
  DFF \memory_reg[20][15]  ( .D(n7105), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[655]), .Q(data_mem_out_wire[655]) );
  DFF \memory_reg[20][14]  ( .D(n7104), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[654]), .Q(data_mem_out_wire[654]) );
  DFF \memory_reg[20][13]  ( .D(n7103), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[653]), .Q(data_mem_out_wire[653]) );
  DFF \memory_reg[20][12]  ( .D(n7102), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[652]), .Q(data_mem_out_wire[652]) );
  DFF \memory_reg[20][11]  ( .D(n7101), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[651]), .Q(data_mem_out_wire[651]) );
  DFF \memory_reg[20][10]  ( .D(n7100), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[650]), .Q(data_mem_out_wire[650]) );
  DFF \memory_reg[20][9]  ( .D(n7099), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[649]), .Q(data_mem_out_wire[649]) );
  DFF \memory_reg[20][8]  ( .D(n7098), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[648]), .Q(data_mem_out_wire[648]) );
  DFF \memory_reg[20][7]  ( .D(n7097), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[647]), .Q(data_mem_out_wire[647]) );
  DFF \memory_reg[20][6]  ( .D(n7096), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[646]), .Q(data_mem_out_wire[646]) );
  DFF \memory_reg[20][5]  ( .D(n7095), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[645]), .Q(data_mem_out_wire[645]) );
  DFF \memory_reg[20][4]  ( .D(n7094), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[644]), .Q(data_mem_out_wire[644]) );
  DFF \memory_reg[20][3]  ( .D(n7093), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[643]), .Q(data_mem_out_wire[643]) );
  DFF \memory_reg[20][2]  ( .D(n7092), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[642]), .Q(data_mem_out_wire[642]) );
  DFF \memory_reg[20][1]  ( .D(n7091), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[641]), .Q(data_mem_out_wire[641]) );
  DFF \memory_reg[20][0]  ( .D(n7090), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[640]), .Q(data_mem_out_wire[640]) );
  DFF \memory_reg[21][31]  ( .D(n7089), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[703]), .Q(data_mem_out_wire[703]) );
  DFF \memory_reg[21][30]  ( .D(n7088), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[702]), .Q(data_mem_out_wire[702]) );
  DFF \memory_reg[21][29]  ( .D(n7087), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[701]), .Q(data_mem_out_wire[701]) );
  DFF \memory_reg[21][28]  ( .D(n7086), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[700]), .Q(data_mem_out_wire[700]) );
  DFF \memory_reg[21][27]  ( .D(n7085), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[699]), .Q(data_mem_out_wire[699]) );
  DFF \memory_reg[21][26]  ( .D(n7084), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[698]), .Q(data_mem_out_wire[698]) );
  DFF \memory_reg[21][25]  ( .D(n7083), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[697]), .Q(data_mem_out_wire[697]) );
  DFF \memory_reg[21][24]  ( .D(n7082), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[696]), .Q(data_mem_out_wire[696]) );
  DFF \memory_reg[21][23]  ( .D(n7081), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[695]), .Q(data_mem_out_wire[695]) );
  DFF \memory_reg[21][22]  ( .D(n7080), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[694]), .Q(data_mem_out_wire[694]) );
  DFF \memory_reg[21][21]  ( .D(n7079), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[693]), .Q(data_mem_out_wire[693]) );
  DFF \memory_reg[21][20]  ( .D(n7078), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[692]), .Q(data_mem_out_wire[692]) );
  DFF \memory_reg[21][19]  ( .D(n7077), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[691]), .Q(data_mem_out_wire[691]) );
  DFF \memory_reg[21][18]  ( .D(n7076), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[690]), .Q(data_mem_out_wire[690]) );
  DFF \memory_reg[21][17]  ( .D(n7075), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[689]), .Q(data_mem_out_wire[689]) );
  DFF \memory_reg[21][16]  ( .D(n7074), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[688]), .Q(data_mem_out_wire[688]) );
  DFF \memory_reg[21][15]  ( .D(n7073), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[687]), .Q(data_mem_out_wire[687]) );
  DFF \memory_reg[21][14]  ( .D(n7072), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[686]), .Q(data_mem_out_wire[686]) );
  DFF \memory_reg[21][13]  ( .D(n7071), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[685]), .Q(data_mem_out_wire[685]) );
  DFF \memory_reg[21][12]  ( .D(n7070), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[684]), .Q(data_mem_out_wire[684]) );
  DFF \memory_reg[21][11]  ( .D(n7069), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[683]), .Q(data_mem_out_wire[683]) );
  DFF \memory_reg[21][10]  ( .D(n7068), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[682]), .Q(data_mem_out_wire[682]) );
  DFF \memory_reg[21][9]  ( .D(n7067), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[681]), .Q(data_mem_out_wire[681]) );
  DFF \memory_reg[21][8]  ( .D(n7066), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[680]), .Q(data_mem_out_wire[680]) );
  DFF \memory_reg[21][7]  ( .D(n7065), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[679]), .Q(data_mem_out_wire[679]) );
  DFF \memory_reg[21][6]  ( .D(n7064), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[678]), .Q(data_mem_out_wire[678]) );
  DFF \memory_reg[21][5]  ( .D(n7063), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[677]), .Q(data_mem_out_wire[677]) );
  DFF \memory_reg[21][4]  ( .D(n7062), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[676]), .Q(data_mem_out_wire[676]) );
  DFF \memory_reg[21][3]  ( .D(n7061), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[675]), .Q(data_mem_out_wire[675]) );
  DFF \memory_reg[21][2]  ( .D(n7060), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[674]), .Q(data_mem_out_wire[674]) );
  DFF \memory_reg[21][1]  ( .D(n7059), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[673]), .Q(data_mem_out_wire[673]) );
  DFF \memory_reg[21][0]  ( .D(n7058), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[672]), .Q(data_mem_out_wire[672]) );
  DFF \memory_reg[22][31]  ( .D(n7057), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[735]), .Q(data_mem_out_wire[735]) );
  DFF \memory_reg[22][30]  ( .D(n7056), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[734]), .Q(data_mem_out_wire[734]) );
  DFF \memory_reg[22][29]  ( .D(n7055), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[733]), .Q(data_mem_out_wire[733]) );
  DFF \memory_reg[22][28]  ( .D(n7054), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[732]), .Q(data_mem_out_wire[732]) );
  DFF \memory_reg[22][27]  ( .D(n7053), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[731]), .Q(data_mem_out_wire[731]) );
  DFF \memory_reg[22][26]  ( .D(n7052), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[730]), .Q(data_mem_out_wire[730]) );
  DFF \memory_reg[22][25]  ( .D(n7051), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[729]), .Q(data_mem_out_wire[729]) );
  DFF \memory_reg[22][24]  ( .D(n7050), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[728]), .Q(data_mem_out_wire[728]) );
  DFF \memory_reg[22][23]  ( .D(n7049), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[727]), .Q(data_mem_out_wire[727]) );
  DFF \memory_reg[22][22]  ( .D(n7048), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[726]), .Q(data_mem_out_wire[726]) );
  DFF \memory_reg[22][21]  ( .D(n7047), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[725]), .Q(data_mem_out_wire[725]) );
  DFF \memory_reg[22][20]  ( .D(n7046), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[724]), .Q(data_mem_out_wire[724]) );
  DFF \memory_reg[22][19]  ( .D(n7045), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[723]), .Q(data_mem_out_wire[723]) );
  DFF \memory_reg[22][18]  ( .D(n7044), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[722]), .Q(data_mem_out_wire[722]) );
  DFF \memory_reg[22][17]  ( .D(n7043), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[721]), .Q(data_mem_out_wire[721]) );
  DFF \memory_reg[22][16]  ( .D(n7042), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[720]), .Q(data_mem_out_wire[720]) );
  DFF \memory_reg[22][15]  ( .D(n7041), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[719]), .Q(data_mem_out_wire[719]) );
  DFF \memory_reg[22][14]  ( .D(n7040), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[718]), .Q(data_mem_out_wire[718]) );
  DFF \memory_reg[22][13]  ( .D(n7039), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[717]), .Q(data_mem_out_wire[717]) );
  DFF \memory_reg[22][12]  ( .D(n7038), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[716]), .Q(data_mem_out_wire[716]) );
  DFF \memory_reg[22][11]  ( .D(n7037), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[715]), .Q(data_mem_out_wire[715]) );
  DFF \memory_reg[22][10]  ( .D(n7036), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[714]), .Q(data_mem_out_wire[714]) );
  DFF \memory_reg[22][9]  ( .D(n7035), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[713]), .Q(data_mem_out_wire[713]) );
  DFF \memory_reg[22][8]  ( .D(n7034), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[712]), .Q(data_mem_out_wire[712]) );
  DFF \memory_reg[22][7]  ( .D(n7033), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[711]), .Q(data_mem_out_wire[711]) );
  DFF \memory_reg[22][6]  ( .D(n7032), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[710]), .Q(data_mem_out_wire[710]) );
  DFF \memory_reg[22][5]  ( .D(n7031), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[709]), .Q(data_mem_out_wire[709]) );
  DFF \memory_reg[22][4]  ( .D(n7030), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[708]), .Q(data_mem_out_wire[708]) );
  DFF \memory_reg[22][3]  ( .D(n7029), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[707]), .Q(data_mem_out_wire[707]) );
  DFF \memory_reg[22][2]  ( .D(n7028), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[706]), .Q(data_mem_out_wire[706]) );
  DFF \memory_reg[22][1]  ( .D(n7027), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[705]), .Q(data_mem_out_wire[705]) );
  DFF \memory_reg[22][0]  ( .D(n7026), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[704]), .Q(data_mem_out_wire[704]) );
  DFF \memory_reg[23][31]  ( .D(n7025), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[767]), .Q(data_mem_out_wire[767]) );
  DFF \memory_reg[23][30]  ( .D(n7024), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[766]), .Q(data_mem_out_wire[766]) );
  DFF \memory_reg[23][29]  ( .D(n7023), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[765]), .Q(data_mem_out_wire[765]) );
  DFF \memory_reg[23][28]  ( .D(n7022), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[764]), .Q(data_mem_out_wire[764]) );
  DFF \memory_reg[23][27]  ( .D(n7021), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[763]), .Q(data_mem_out_wire[763]) );
  DFF \memory_reg[23][26]  ( .D(n7020), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[762]), .Q(data_mem_out_wire[762]) );
  DFF \memory_reg[23][25]  ( .D(n7019), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[761]), .Q(data_mem_out_wire[761]) );
  DFF \memory_reg[23][24]  ( .D(n7018), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[760]), .Q(data_mem_out_wire[760]) );
  DFF \memory_reg[23][23]  ( .D(n7017), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[759]), .Q(data_mem_out_wire[759]) );
  DFF \memory_reg[23][22]  ( .D(n7016), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[758]), .Q(data_mem_out_wire[758]) );
  DFF \memory_reg[23][21]  ( .D(n7015), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[757]), .Q(data_mem_out_wire[757]) );
  DFF \memory_reg[23][20]  ( .D(n7014), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[756]), .Q(data_mem_out_wire[756]) );
  DFF \memory_reg[23][19]  ( .D(n7013), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[755]), .Q(data_mem_out_wire[755]) );
  DFF \memory_reg[23][18]  ( .D(n7012), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[754]), .Q(data_mem_out_wire[754]) );
  DFF \memory_reg[23][17]  ( .D(n7011), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[753]), .Q(data_mem_out_wire[753]) );
  DFF \memory_reg[23][16]  ( .D(n7010), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[752]), .Q(data_mem_out_wire[752]) );
  DFF \memory_reg[23][15]  ( .D(n7009), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[751]), .Q(data_mem_out_wire[751]) );
  DFF \memory_reg[23][14]  ( .D(n7008), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[750]), .Q(data_mem_out_wire[750]) );
  DFF \memory_reg[23][13]  ( .D(n7007), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[749]), .Q(data_mem_out_wire[749]) );
  DFF \memory_reg[23][12]  ( .D(n7006), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[748]), .Q(data_mem_out_wire[748]) );
  DFF \memory_reg[23][11]  ( .D(n7005), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[747]), .Q(data_mem_out_wire[747]) );
  DFF \memory_reg[23][10]  ( .D(n7004), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[746]), .Q(data_mem_out_wire[746]) );
  DFF \memory_reg[23][9]  ( .D(n7003), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[745]), .Q(data_mem_out_wire[745]) );
  DFF \memory_reg[23][8]  ( .D(n7002), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[744]), .Q(data_mem_out_wire[744]) );
  DFF \memory_reg[23][7]  ( .D(n7001), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[743]), .Q(data_mem_out_wire[743]) );
  DFF \memory_reg[23][6]  ( .D(n7000), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[742]), .Q(data_mem_out_wire[742]) );
  DFF \memory_reg[23][5]  ( .D(n6999), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[741]), .Q(data_mem_out_wire[741]) );
  DFF \memory_reg[23][4]  ( .D(n6998), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[740]), .Q(data_mem_out_wire[740]) );
  DFF \memory_reg[23][3]  ( .D(n6997), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[739]), .Q(data_mem_out_wire[739]) );
  DFF \memory_reg[23][2]  ( .D(n6996), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[738]), .Q(data_mem_out_wire[738]) );
  DFF \memory_reg[23][1]  ( .D(n6995), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[737]), .Q(data_mem_out_wire[737]) );
  DFF \memory_reg[23][0]  ( .D(n6994), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[736]), .Q(data_mem_out_wire[736]) );
  DFF \memory_reg[24][31]  ( .D(n6993), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[799]), .Q(data_mem_out_wire[799]) );
  DFF \memory_reg[24][30]  ( .D(n6992), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[798]), .Q(data_mem_out_wire[798]) );
  DFF \memory_reg[24][29]  ( .D(n6991), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[797]), .Q(data_mem_out_wire[797]) );
  DFF \memory_reg[24][28]  ( .D(n6990), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[796]), .Q(data_mem_out_wire[796]) );
  DFF \memory_reg[24][27]  ( .D(n6989), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[795]), .Q(data_mem_out_wire[795]) );
  DFF \memory_reg[24][26]  ( .D(n6988), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[794]), .Q(data_mem_out_wire[794]) );
  DFF \memory_reg[24][25]  ( .D(n6987), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[793]), .Q(data_mem_out_wire[793]) );
  DFF \memory_reg[24][24]  ( .D(n6986), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[792]), .Q(data_mem_out_wire[792]) );
  DFF \memory_reg[24][23]  ( .D(n6985), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[791]), .Q(data_mem_out_wire[791]) );
  DFF \memory_reg[24][22]  ( .D(n6984), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[790]), .Q(data_mem_out_wire[790]) );
  DFF \memory_reg[24][21]  ( .D(n6983), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[789]), .Q(data_mem_out_wire[789]) );
  DFF \memory_reg[24][20]  ( .D(n6982), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[788]), .Q(data_mem_out_wire[788]) );
  DFF \memory_reg[24][19]  ( .D(n6981), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[787]), .Q(data_mem_out_wire[787]) );
  DFF \memory_reg[24][18]  ( .D(n6980), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[786]), .Q(data_mem_out_wire[786]) );
  DFF \memory_reg[24][17]  ( .D(n6979), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[785]), .Q(data_mem_out_wire[785]) );
  DFF \memory_reg[24][16]  ( .D(n6978), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[784]), .Q(data_mem_out_wire[784]) );
  DFF \memory_reg[24][15]  ( .D(n6977), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[783]), .Q(data_mem_out_wire[783]) );
  DFF \memory_reg[24][14]  ( .D(n6976), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[782]), .Q(data_mem_out_wire[782]) );
  DFF \memory_reg[24][13]  ( .D(n6975), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[781]), .Q(data_mem_out_wire[781]) );
  DFF \memory_reg[24][12]  ( .D(n6974), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[780]), .Q(data_mem_out_wire[780]) );
  DFF \memory_reg[24][11]  ( .D(n6973), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[779]), .Q(data_mem_out_wire[779]) );
  DFF \memory_reg[24][10]  ( .D(n6972), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[778]), .Q(data_mem_out_wire[778]) );
  DFF \memory_reg[24][9]  ( .D(n6971), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[777]), .Q(data_mem_out_wire[777]) );
  DFF \memory_reg[24][8]  ( .D(n6970), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[776]), .Q(data_mem_out_wire[776]) );
  DFF \memory_reg[24][7]  ( .D(n6969), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[775]), .Q(data_mem_out_wire[775]) );
  DFF \memory_reg[24][6]  ( .D(n6968), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[774]), .Q(data_mem_out_wire[774]) );
  DFF \memory_reg[24][5]  ( .D(n6967), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[773]), .Q(data_mem_out_wire[773]) );
  DFF \memory_reg[24][4]  ( .D(n6966), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[772]), .Q(data_mem_out_wire[772]) );
  DFF \memory_reg[24][3]  ( .D(n6965), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[771]), .Q(data_mem_out_wire[771]) );
  DFF \memory_reg[24][2]  ( .D(n6964), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[770]), .Q(data_mem_out_wire[770]) );
  DFF \memory_reg[24][1]  ( .D(n6963), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[769]), .Q(data_mem_out_wire[769]) );
  DFF \memory_reg[24][0]  ( .D(n6962), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[768]), .Q(data_mem_out_wire[768]) );
  DFF \memory_reg[25][31]  ( .D(n6961), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[831]), .Q(data_mem_out_wire[831]) );
  DFF \memory_reg[25][30]  ( .D(n6960), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[830]), .Q(data_mem_out_wire[830]) );
  DFF \memory_reg[25][29]  ( .D(n6959), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[829]), .Q(data_mem_out_wire[829]) );
  DFF \memory_reg[25][28]  ( .D(n6958), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[828]), .Q(data_mem_out_wire[828]) );
  DFF \memory_reg[25][27]  ( .D(n6957), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[827]), .Q(data_mem_out_wire[827]) );
  DFF \memory_reg[25][26]  ( .D(n6956), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[826]), .Q(data_mem_out_wire[826]) );
  DFF \memory_reg[25][25]  ( .D(n6955), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[825]), .Q(data_mem_out_wire[825]) );
  DFF \memory_reg[25][24]  ( .D(n6954), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[824]), .Q(data_mem_out_wire[824]) );
  DFF \memory_reg[25][23]  ( .D(n6953), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[823]), .Q(data_mem_out_wire[823]) );
  DFF \memory_reg[25][22]  ( .D(n6952), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[822]), .Q(data_mem_out_wire[822]) );
  DFF \memory_reg[25][21]  ( .D(n6951), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[821]), .Q(data_mem_out_wire[821]) );
  DFF \memory_reg[25][20]  ( .D(n6950), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[820]), .Q(data_mem_out_wire[820]) );
  DFF \memory_reg[25][19]  ( .D(n6949), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[819]), .Q(data_mem_out_wire[819]) );
  DFF \memory_reg[25][18]  ( .D(n6948), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[818]), .Q(data_mem_out_wire[818]) );
  DFF \memory_reg[25][17]  ( .D(n6947), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[817]), .Q(data_mem_out_wire[817]) );
  DFF \memory_reg[25][16]  ( .D(n6946), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[816]), .Q(data_mem_out_wire[816]) );
  DFF \memory_reg[25][15]  ( .D(n6945), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[815]), .Q(data_mem_out_wire[815]) );
  DFF \memory_reg[25][14]  ( .D(n6944), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[814]), .Q(data_mem_out_wire[814]) );
  DFF \memory_reg[25][13]  ( .D(n6943), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[813]), .Q(data_mem_out_wire[813]) );
  DFF \memory_reg[25][12]  ( .D(n6942), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[812]), .Q(data_mem_out_wire[812]) );
  DFF \memory_reg[25][11]  ( .D(n6941), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[811]), .Q(data_mem_out_wire[811]) );
  DFF \memory_reg[25][10]  ( .D(n6940), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[810]), .Q(data_mem_out_wire[810]) );
  DFF \memory_reg[25][9]  ( .D(n6939), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[809]), .Q(data_mem_out_wire[809]) );
  DFF \memory_reg[25][8]  ( .D(n6938), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[808]), .Q(data_mem_out_wire[808]) );
  DFF \memory_reg[25][7]  ( .D(n6937), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[807]), .Q(data_mem_out_wire[807]) );
  DFF \memory_reg[25][6]  ( .D(n6936), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[806]), .Q(data_mem_out_wire[806]) );
  DFF \memory_reg[25][5]  ( .D(n6935), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[805]), .Q(data_mem_out_wire[805]) );
  DFF \memory_reg[25][4]  ( .D(n6934), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[804]), .Q(data_mem_out_wire[804]) );
  DFF \memory_reg[25][3]  ( .D(n6933), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[803]), .Q(data_mem_out_wire[803]) );
  DFF \memory_reg[25][2]  ( .D(n6932), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[802]), .Q(data_mem_out_wire[802]) );
  DFF \memory_reg[25][1]  ( .D(n6931), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[801]), .Q(data_mem_out_wire[801]) );
  DFF \memory_reg[25][0]  ( .D(n6930), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[800]), .Q(data_mem_out_wire[800]) );
  DFF \memory_reg[26][31]  ( .D(n6929), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[863]), .Q(data_mem_out_wire[863]) );
  DFF \memory_reg[26][30]  ( .D(n6928), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[862]), .Q(data_mem_out_wire[862]) );
  DFF \memory_reg[26][29]  ( .D(n6927), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[861]), .Q(data_mem_out_wire[861]) );
  DFF \memory_reg[26][28]  ( .D(n6926), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[860]), .Q(data_mem_out_wire[860]) );
  DFF \memory_reg[26][27]  ( .D(n6925), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[859]), .Q(data_mem_out_wire[859]) );
  DFF \memory_reg[26][26]  ( .D(n6924), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[858]), .Q(data_mem_out_wire[858]) );
  DFF \memory_reg[26][25]  ( .D(n6923), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[857]), .Q(data_mem_out_wire[857]) );
  DFF \memory_reg[26][24]  ( .D(n6922), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[856]), .Q(data_mem_out_wire[856]) );
  DFF \memory_reg[26][23]  ( .D(n6921), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[855]), .Q(data_mem_out_wire[855]) );
  DFF \memory_reg[26][22]  ( .D(n6920), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[854]), .Q(data_mem_out_wire[854]) );
  DFF \memory_reg[26][21]  ( .D(n6919), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[853]), .Q(data_mem_out_wire[853]) );
  DFF \memory_reg[26][20]  ( .D(n6918), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[852]), .Q(data_mem_out_wire[852]) );
  DFF \memory_reg[26][19]  ( .D(n6917), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[851]), .Q(data_mem_out_wire[851]) );
  DFF \memory_reg[26][18]  ( .D(n6916), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[850]), .Q(data_mem_out_wire[850]) );
  DFF \memory_reg[26][17]  ( .D(n6915), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[849]), .Q(data_mem_out_wire[849]) );
  DFF \memory_reg[26][16]  ( .D(n6914), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[848]), .Q(data_mem_out_wire[848]) );
  DFF \memory_reg[26][15]  ( .D(n6913), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[847]), .Q(data_mem_out_wire[847]) );
  DFF \memory_reg[26][14]  ( .D(n6912), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[846]), .Q(data_mem_out_wire[846]) );
  DFF \memory_reg[26][13]  ( .D(n6911), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[845]), .Q(data_mem_out_wire[845]) );
  DFF \memory_reg[26][12]  ( .D(n6910), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[844]), .Q(data_mem_out_wire[844]) );
  DFF \memory_reg[26][11]  ( .D(n6909), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[843]), .Q(data_mem_out_wire[843]) );
  DFF \memory_reg[26][10]  ( .D(n6908), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[842]), .Q(data_mem_out_wire[842]) );
  DFF \memory_reg[26][9]  ( .D(n6907), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[841]), .Q(data_mem_out_wire[841]) );
  DFF \memory_reg[26][8]  ( .D(n6906), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[840]), .Q(data_mem_out_wire[840]) );
  DFF \memory_reg[26][7]  ( .D(n6905), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[839]), .Q(data_mem_out_wire[839]) );
  DFF \memory_reg[26][6]  ( .D(n6904), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[838]), .Q(data_mem_out_wire[838]) );
  DFF \memory_reg[26][5]  ( .D(n6903), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[837]), .Q(data_mem_out_wire[837]) );
  DFF \memory_reg[26][4]  ( .D(n6902), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[836]), .Q(data_mem_out_wire[836]) );
  DFF \memory_reg[26][3]  ( .D(n6901), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[835]), .Q(data_mem_out_wire[835]) );
  DFF \memory_reg[26][2]  ( .D(n6900), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[834]), .Q(data_mem_out_wire[834]) );
  DFF \memory_reg[26][1]  ( .D(n6899), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[833]), .Q(data_mem_out_wire[833]) );
  DFF \memory_reg[26][0]  ( .D(n6898), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[832]), .Q(data_mem_out_wire[832]) );
  DFF \memory_reg[27][31]  ( .D(n6897), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[895]), .Q(data_mem_out_wire[895]) );
  DFF \memory_reg[27][30]  ( .D(n6896), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[894]), .Q(data_mem_out_wire[894]) );
  DFF \memory_reg[27][29]  ( .D(n6895), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[893]), .Q(data_mem_out_wire[893]) );
  DFF \memory_reg[27][28]  ( .D(n6894), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[892]), .Q(data_mem_out_wire[892]) );
  DFF \memory_reg[27][27]  ( .D(n6893), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[891]), .Q(data_mem_out_wire[891]) );
  DFF \memory_reg[27][26]  ( .D(n6892), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[890]), .Q(data_mem_out_wire[890]) );
  DFF \memory_reg[27][25]  ( .D(n6891), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[889]), .Q(data_mem_out_wire[889]) );
  DFF \memory_reg[27][24]  ( .D(n6890), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[888]), .Q(data_mem_out_wire[888]) );
  DFF \memory_reg[27][23]  ( .D(n6889), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[887]), .Q(data_mem_out_wire[887]) );
  DFF \memory_reg[27][22]  ( .D(n6888), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[886]), .Q(data_mem_out_wire[886]) );
  DFF \memory_reg[27][21]  ( .D(n6887), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[885]), .Q(data_mem_out_wire[885]) );
  DFF \memory_reg[27][20]  ( .D(n6886), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[884]), .Q(data_mem_out_wire[884]) );
  DFF \memory_reg[27][19]  ( .D(n6885), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[883]), .Q(data_mem_out_wire[883]) );
  DFF \memory_reg[27][18]  ( .D(n6884), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[882]), .Q(data_mem_out_wire[882]) );
  DFF \memory_reg[27][17]  ( .D(n6883), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[881]), .Q(data_mem_out_wire[881]) );
  DFF \memory_reg[27][16]  ( .D(n6882), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[880]), .Q(data_mem_out_wire[880]) );
  DFF \memory_reg[27][15]  ( .D(n6881), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[879]), .Q(data_mem_out_wire[879]) );
  DFF \memory_reg[27][14]  ( .D(n6880), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[878]), .Q(data_mem_out_wire[878]) );
  DFF \memory_reg[27][13]  ( .D(n6879), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[877]), .Q(data_mem_out_wire[877]) );
  DFF \memory_reg[27][12]  ( .D(n6878), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[876]), .Q(data_mem_out_wire[876]) );
  DFF \memory_reg[27][11]  ( .D(n6877), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[875]), .Q(data_mem_out_wire[875]) );
  DFF \memory_reg[27][10]  ( .D(n6876), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[874]), .Q(data_mem_out_wire[874]) );
  DFF \memory_reg[27][9]  ( .D(n6875), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[873]), .Q(data_mem_out_wire[873]) );
  DFF \memory_reg[27][8]  ( .D(n6874), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[872]), .Q(data_mem_out_wire[872]) );
  DFF \memory_reg[27][7]  ( .D(n6873), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[871]), .Q(data_mem_out_wire[871]) );
  DFF \memory_reg[27][6]  ( .D(n6872), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[870]), .Q(data_mem_out_wire[870]) );
  DFF \memory_reg[27][5]  ( .D(n6871), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[869]), .Q(data_mem_out_wire[869]) );
  DFF \memory_reg[27][4]  ( .D(n6870), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[868]), .Q(data_mem_out_wire[868]) );
  DFF \memory_reg[27][3]  ( .D(n6869), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[867]), .Q(data_mem_out_wire[867]) );
  DFF \memory_reg[27][2]  ( .D(n6868), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[866]), .Q(data_mem_out_wire[866]) );
  DFF \memory_reg[27][1]  ( .D(n6867), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[865]), .Q(data_mem_out_wire[865]) );
  DFF \memory_reg[27][0]  ( .D(n6866), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[864]), .Q(data_mem_out_wire[864]) );
  DFF \memory_reg[28][31]  ( .D(n6865), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[927]), .Q(data_mem_out_wire[927]) );
  DFF \memory_reg[28][30]  ( .D(n6864), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[926]), .Q(data_mem_out_wire[926]) );
  DFF \memory_reg[28][29]  ( .D(n6863), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[925]), .Q(data_mem_out_wire[925]) );
  DFF \memory_reg[28][28]  ( .D(n6862), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[924]), .Q(data_mem_out_wire[924]) );
  DFF \memory_reg[28][27]  ( .D(n6861), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[923]), .Q(data_mem_out_wire[923]) );
  DFF \memory_reg[28][26]  ( .D(n6860), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[922]), .Q(data_mem_out_wire[922]) );
  DFF \memory_reg[28][25]  ( .D(n6859), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[921]), .Q(data_mem_out_wire[921]) );
  DFF \memory_reg[28][24]  ( .D(n6858), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[920]), .Q(data_mem_out_wire[920]) );
  DFF \memory_reg[28][23]  ( .D(n6857), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[919]), .Q(data_mem_out_wire[919]) );
  DFF \memory_reg[28][22]  ( .D(n6856), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[918]), .Q(data_mem_out_wire[918]) );
  DFF \memory_reg[28][21]  ( .D(n6855), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[917]), .Q(data_mem_out_wire[917]) );
  DFF \memory_reg[28][20]  ( .D(n6854), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[916]), .Q(data_mem_out_wire[916]) );
  DFF \memory_reg[28][19]  ( .D(n6853), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[915]), .Q(data_mem_out_wire[915]) );
  DFF \memory_reg[28][18]  ( .D(n6852), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[914]), .Q(data_mem_out_wire[914]) );
  DFF \memory_reg[28][17]  ( .D(n6851), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[913]), .Q(data_mem_out_wire[913]) );
  DFF \memory_reg[28][16]  ( .D(n6850), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[912]), .Q(data_mem_out_wire[912]) );
  DFF \memory_reg[28][15]  ( .D(n6849), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[911]), .Q(data_mem_out_wire[911]) );
  DFF \memory_reg[28][14]  ( .D(n6848), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[910]), .Q(data_mem_out_wire[910]) );
  DFF \memory_reg[28][13]  ( .D(n6847), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[909]), .Q(data_mem_out_wire[909]) );
  DFF \memory_reg[28][12]  ( .D(n6846), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[908]), .Q(data_mem_out_wire[908]) );
  DFF \memory_reg[28][11]  ( .D(n6845), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[907]), .Q(data_mem_out_wire[907]) );
  DFF \memory_reg[28][10]  ( .D(n6844), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[906]), .Q(data_mem_out_wire[906]) );
  DFF \memory_reg[28][9]  ( .D(n6843), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[905]), .Q(data_mem_out_wire[905]) );
  DFF \memory_reg[28][8]  ( .D(n6842), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[904]), .Q(data_mem_out_wire[904]) );
  DFF \memory_reg[28][7]  ( .D(n6841), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[903]), .Q(data_mem_out_wire[903]) );
  DFF \memory_reg[28][6]  ( .D(n6840), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[902]), .Q(data_mem_out_wire[902]) );
  DFF \memory_reg[28][5]  ( .D(n6839), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[901]), .Q(data_mem_out_wire[901]) );
  DFF \memory_reg[28][4]  ( .D(n6838), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[900]), .Q(data_mem_out_wire[900]) );
  DFF \memory_reg[28][3]  ( .D(n6837), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[899]), .Q(data_mem_out_wire[899]) );
  DFF \memory_reg[28][2]  ( .D(n6836), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[898]), .Q(data_mem_out_wire[898]) );
  DFF \memory_reg[28][1]  ( .D(n6835), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[897]), .Q(data_mem_out_wire[897]) );
  DFF \memory_reg[28][0]  ( .D(n6834), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[896]), .Q(data_mem_out_wire[896]) );
  DFF \memory_reg[29][31]  ( .D(n6833), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[959]), .Q(data_mem_out_wire[959]) );
  DFF \memory_reg[29][30]  ( .D(n6832), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[958]), .Q(data_mem_out_wire[958]) );
  DFF \memory_reg[29][29]  ( .D(n6831), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[957]), .Q(data_mem_out_wire[957]) );
  DFF \memory_reg[29][28]  ( .D(n6830), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[956]), .Q(data_mem_out_wire[956]) );
  DFF \memory_reg[29][27]  ( .D(n6829), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[955]), .Q(data_mem_out_wire[955]) );
  DFF \memory_reg[29][26]  ( .D(n6828), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[954]), .Q(data_mem_out_wire[954]) );
  DFF \memory_reg[29][25]  ( .D(n6827), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[953]), .Q(data_mem_out_wire[953]) );
  DFF \memory_reg[29][24]  ( .D(n6826), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[952]), .Q(data_mem_out_wire[952]) );
  DFF \memory_reg[29][23]  ( .D(n6825), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[951]), .Q(data_mem_out_wire[951]) );
  DFF \memory_reg[29][22]  ( .D(n6824), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[950]), .Q(data_mem_out_wire[950]) );
  DFF \memory_reg[29][21]  ( .D(n6823), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[949]), .Q(data_mem_out_wire[949]) );
  DFF \memory_reg[29][20]  ( .D(n6822), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[948]), .Q(data_mem_out_wire[948]) );
  DFF \memory_reg[29][19]  ( .D(n6821), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[947]), .Q(data_mem_out_wire[947]) );
  DFF \memory_reg[29][18]  ( .D(n6820), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[946]), .Q(data_mem_out_wire[946]) );
  DFF \memory_reg[29][17]  ( .D(n6819), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[945]), .Q(data_mem_out_wire[945]) );
  DFF \memory_reg[29][16]  ( .D(n6818), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[944]), .Q(data_mem_out_wire[944]) );
  DFF \memory_reg[29][15]  ( .D(n6817), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[943]), .Q(data_mem_out_wire[943]) );
  DFF \memory_reg[29][14]  ( .D(n6816), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[942]), .Q(data_mem_out_wire[942]) );
  DFF \memory_reg[29][13]  ( .D(n6815), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[941]), .Q(data_mem_out_wire[941]) );
  DFF \memory_reg[29][12]  ( .D(n6814), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[940]), .Q(data_mem_out_wire[940]) );
  DFF \memory_reg[29][11]  ( .D(n6813), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[939]), .Q(data_mem_out_wire[939]) );
  DFF \memory_reg[29][10]  ( .D(n6812), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[938]), .Q(data_mem_out_wire[938]) );
  DFF \memory_reg[29][9]  ( .D(n6811), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[937]), .Q(data_mem_out_wire[937]) );
  DFF \memory_reg[29][8]  ( .D(n6810), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[936]), .Q(data_mem_out_wire[936]) );
  DFF \memory_reg[29][7]  ( .D(n6809), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[935]), .Q(data_mem_out_wire[935]) );
  DFF \memory_reg[29][6]  ( .D(n6808), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[934]), .Q(data_mem_out_wire[934]) );
  DFF \memory_reg[29][5]  ( .D(n6807), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[933]), .Q(data_mem_out_wire[933]) );
  DFF \memory_reg[29][4]  ( .D(n6806), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[932]), .Q(data_mem_out_wire[932]) );
  DFF \memory_reg[29][3]  ( .D(n6805), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[931]), .Q(data_mem_out_wire[931]) );
  DFF \memory_reg[29][2]  ( .D(n6804), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[930]), .Q(data_mem_out_wire[930]) );
  DFF \memory_reg[29][1]  ( .D(n6803), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[929]), .Q(data_mem_out_wire[929]) );
  DFF \memory_reg[29][0]  ( .D(n6802), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[928]), .Q(data_mem_out_wire[928]) );
  DFF \memory_reg[30][31]  ( .D(n6801), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[991]), .Q(data_mem_out_wire[991]) );
  DFF \memory_reg[30][30]  ( .D(n6800), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[990]), .Q(data_mem_out_wire[990]) );
  DFF \memory_reg[30][29]  ( .D(n6799), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[989]), .Q(data_mem_out_wire[989]) );
  DFF \memory_reg[30][28]  ( .D(n6798), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[988]), .Q(data_mem_out_wire[988]) );
  DFF \memory_reg[30][27]  ( .D(n6797), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[987]), .Q(data_mem_out_wire[987]) );
  DFF \memory_reg[30][26]  ( .D(n6796), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[986]), .Q(data_mem_out_wire[986]) );
  DFF \memory_reg[30][25]  ( .D(n6795), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[985]), .Q(data_mem_out_wire[985]) );
  DFF \memory_reg[30][24]  ( .D(n6794), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[984]), .Q(data_mem_out_wire[984]) );
  DFF \memory_reg[30][23]  ( .D(n6793), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[983]), .Q(data_mem_out_wire[983]) );
  DFF \memory_reg[30][22]  ( .D(n6792), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[982]), .Q(data_mem_out_wire[982]) );
  DFF \memory_reg[30][21]  ( .D(n6791), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[981]), .Q(data_mem_out_wire[981]) );
  DFF \memory_reg[30][20]  ( .D(n6790), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[980]), .Q(data_mem_out_wire[980]) );
  DFF \memory_reg[30][19]  ( .D(n6789), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[979]), .Q(data_mem_out_wire[979]) );
  DFF \memory_reg[30][18]  ( .D(n6788), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[978]), .Q(data_mem_out_wire[978]) );
  DFF \memory_reg[30][17]  ( .D(n6787), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[977]), .Q(data_mem_out_wire[977]) );
  DFF \memory_reg[30][16]  ( .D(n6786), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[976]), .Q(data_mem_out_wire[976]) );
  DFF \memory_reg[30][15]  ( .D(n6785), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[975]), .Q(data_mem_out_wire[975]) );
  DFF \memory_reg[30][14]  ( .D(n6784), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[974]), .Q(data_mem_out_wire[974]) );
  DFF \memory_reg[30][13]  ( .D(n6783), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[973]), .Q(data_mem_out_wire[973]) );
  DFF \memory_reg[30][12]  ( .D(n6782), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[972]), .Q(data_mem_out_wire[972]) );
  DFF \memory_reg[30][11]  ( .D(n6781), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[971]), .Q(data_mem_out_wire[971]) );
  DFF \memory_reg[30][10]  ( .D(n6780), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[970]), .Q(data_mem_out_wire[970]) );
  DFF \memory_reg[30][9]  ( .D(n6779), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[969]), .Q(data_mem_out_wire[969]) );
  DFF \memory_reg[30][8]  ( .D(n6778), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[968]), .Q(data_mem_out_wire[968]) );
  DFF \memory_reg[30][7]  ( .D(n6777), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[967]), .Q(data_mem_out_wire[967]) );
  DFF \memory_reg[30][6]  ( .D(n6776), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[966]), .Q(data_mem_out_wire[966]) );
  DFF \memory_reg[30][5]  ( .D(n6775), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[965]), .Q(data_mem_out_wire[965]) );
  DFF \memory_reg[30][4]  ( .D(n6774), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[964]), .Q(data_mem_out_wire[964]) );
  DFF \memory_reg[30][3]  ( .D(n6773), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[963]), .Q(data_mem_out_wire[963]) );
  DFF \memory_reg[30][2]  ( .D(n6772), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[962]), .Q(data_mem_out_wire[962]) );
  DFF \memory_reg[30][1]  ( .D(n6771), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[961]), .Q(data_mem_out_wire[961]) );
  DFF \memory_reg[30][0]  ( .D(n6770), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[960]), .Q(data_mem_out_wire[960]) );
  DFF \memory_reg[31][31]  ( .D(n6769), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1023]), .Q(data_mem_out_wire[1023]) );
  DFF \memory_reg[31][30]  ( .D(n6768), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1022]), .Q(data_mem_out_wire[1022]) );
  DFF \memory_reg[31][29]  ( .D(n6767), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1021]), .Q(data_mem_out_wire[1021]) );
  DFF \memory_reg[31][28]  ( .D(n6766), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1020]), .Q(data_mem_out_wire[1020]) );
  DFF \memory_reg[31][27]  ( .D(n6765), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1019]), .Q(data_mem_out_wire[1019]) );
  DFF \memory_reg[31][26]  ( .D(n6764), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1018]), .Q(data_mem_out_wire[1018]) );
  DFF \memory_reg[31][25]  ( .D(n6763), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1017]), .Q(data_mem_out_wire[1017]) );
  DFF \memory_reg[31][24]  ( .D(n6762), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1016]), .Q(data_mem_out_wire[1016]) );
  DFF \memory_reg[31][23]  ( .D(n6761), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1015]), .Q(data_mem_out_wire[1015]) );
  DFF \memory_reg[31][22]  ( .D(n6760), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1014]), .Q(data_mem_out_wire[1014]) );
  DFF \memory_reg[31][21]  ( .D(n6759), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1013]), .Q(data_mem_out_wire[1013]) );
  DFF \memory_reg[31][20]  ( .D(n6758), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1012]), .Q(data_mem_out_wire[1012]) );
  DFF \memory_reg[31][19]  ( .D(n6757), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1011]), .Q(data_mem_out_wire[1011]) );
  DFF \memory_reg[31][18]  ( .D(n6756), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1010]), .Q(data_mem_out_wire[1010]) );
  DFF \memory_reg[31][17]  ( .D(n6755), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1009]), .Q(data_mem_out_wire[1009]) );
  DFF \memory_reg[31][16]  ( .D(n6754), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1008]), .Q(data_mem_out_wire[1008]) );
  DFF \memory_reg[31][15]  ( .D(n6753), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1007]), .Q(data_mem_out_wire[1007]) );
  DFF \memory_reg[31][14]  ( .D(n6752), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1006]), .Q(data_mem_out_wire[1006]) );
  DFF \memory_reg[31][13]  ( .D(n6751), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1005]), .Q(data_mem_out_wire[1005]) );
  DFF \memory_reg[31][12]  ( .D(n6750), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1004]), .Q(data_mem_out_wire[1004]) );
  DFF \memory_reg[31][11]  ( .D(n6749), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1003]), .Q(data_mem_out_wire[1003]) );
  DFF \memory_reg[31][10]  ( .D(n6748), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1002]), .Q(data_mem_out_wire[1002]) );
  DFF \memory_reg[31][9]  ( .D(n6747), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1001]), .Q(data_mem_out_wire[1001]) );
  DFF \memory_reg[31][8]  ( .D(n6746), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1000]), .Q(data_mem_out_wire[1000]) );
  DFF \memory_reg[31][7]  ( .D(n6745), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[999]), .Q(data_mem_out_wire[999]) );
  DFF \memory_reg[31][6]  ( .D(n6744), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[998]), .Q(data_mem_out_wire[998]) );
  DFF \memory_reg[31][5]  ( .D(n6743), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[997]), .Q(data_mem_out_wire[997]) );
  DFF \memory_reg[31][4]  ( .D(n6742), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[996]), .Q(data_mem_out_wire[996]) );
  DFF \memory_reg[31][3]  ( .D(n6741), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[995]), .Q(data_mem_out_wire[995]) );
  DFF \memory_reg[31][2]  ( .D(n6740), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[994]), .Q(data_mem_out_wire[994]) );
  DFF \memory_reg[31][1]  ( .D(n6739), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[993]), .Q(data_mem_out_wire[993]) );
  DFF \memory_reg[31][0]  ( .D(n6738), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[992]), .Q(data_mem_out_wire[992]) );
  DFF \memory_reg[32][31]  ( .D(n6737), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1055]), .Q(data_mem_out_wire[1055]) );
  DFF \memory_reg[32][30]  ( .D(n6736), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1054]), .Q(data_mem_out_wire[1054]) );
  DFF \memory_reg[32][29]  ( .D(n6735), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1053]), .Q(data_mem_out_wire[1053]) );
  DFF \memory_reg[32][28]  ( .D(n6734), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1052]), .Q(data_mem_out_wire[1052]) );
  DFF \memory_reg[32][27]  ( .D(n6733), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1051]), .Q(data_mem_out_wire[1051]) );
  DFF \memory_reg[32][26]  ( .D(n6732), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1050]), .Q(data_mem_out_wire[1050]) );
  DFF \memory_reg[32][25]  ( .D(n6731), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1049]), .Q(data_mem_out_wire[1049]) );
  DFF \memory_reg[32][24]  ( .D(n6730), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1048]), .Q(data_mem_out_wire[1048]) );
  DFF \memory_reg[32][23]  ( .D(n6729), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1047]), .Q(data_mem_out_wire[1047]) );
  DFF \memory_reg[32][22]  ( .D(n6728), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1046]), .Q(data_mem_out_wire[1046]) );
  DFF \memory_reg[32][21]  ( .D(n6727), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1045]), .Q(data_mem_out_wire[1045]) );
  DFF \memory_reg[32][20]  ( .D(n6726), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1044]), .Q(data_mem_out_wire[1044]) );
  DFF \memory_reg[32][19]  ( .D(n6725), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1043]), .Q(data_mem_out_wire[1043]) );
  DFF \memory_reg[32][18]  ( .D(n6724), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1042]), .Q(data_mem_out_wire[1042]) );
  DFF \memory_reg[32][17]  ( .D(n6723), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1041]), .Q(data_mem_out_wire[1041]) );
  DFF \memory_reg[32][16]  ( .D(n6722), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1040]), .Q(data_mem_out_wire[1040]) );
  DFF \memory_reg[32][15]  ( .D(n6721), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1039]), .Q(data_mem_out_wire[1039]) );
  DFF \memory_reg[32][14]  ( .D(n6720), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1038]), .Q(data_mem_out_wire[1038]) );
  DFF \memory_reg[32][13]  ( .D(n6719), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1037]), .Q(data_mem_out_wire[1037]) );
  DFF \memory_reg[32][12]  ( .D(n6718), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1036]), .Q(data_mem_out_wire[1036]) );
  DFF \memory_reg[32][11]  ( .D(n6717), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1035]), .Q(data_mem_out_wire[1035]) );
  DFF \memory_reg[32][10]  ( .D(n6716), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1034]), .Q(data_mem_out_wire[1034]) );
  DFF \memory_reg[32][9]  ( .D(n6715), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1033]), .Q(data_mem_out_wire[1033]) );
  DFF \memory_reg[32][8]  ( .D(n6714), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1032]), .Q(data_mem_out_wire[1032]) );
  DFF \memory_reg[32][7]  ( .D(n6713), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1031]), .Q(data_mem_out_wire[1031]) );
  DFF \memory_reg[32][6]  ( .D(n6712), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1030]), .Q(data_mem_out_wire[1030]) );
  DFF \memory_reg[32][5]  ( .D(n6711), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1029]), .Q(data_mem_out_wire[1029]) );
  DFF \memory_reg[32][4]  ( .D(n6710), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1028]), .Q(data_mem_out_wire[1028]) );
  DFF \memory_reg[32][3]  ( .D(n6709), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1027]), .Q(data_mem_out_wire[1027]) );
  DFF \memory_reg[32][2]  ( .D(n6708), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1026]), .Q(data_mem_out_wire[1026]) );
  DFF \memory_reg[32][1]  ( .D(n6707), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1025]), .Q(data_mem_out_wire[1025]) );
  DFF \memory_reg[32][0]  ( .D(n6706), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1024]), .Q(data_mem_out_wire[1024]) );
  DFF \memory_reg[33][31]  ( .D(n6705), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1087]), .Q(data_mem_out_wire[1087]) );
  DFF \memory_reg[33][30]  ( .D(n6704), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1086]), .Q(data_mem_out_wire[1086]) );
  DFF \memory_reg[33][29]  ( .D(n6703), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1085]), .Q(data_mem_out_wire[1085]) );
  DFF \memory_reg[33][28]  ( .D(n6702), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1084]), .Q(data_mem_out_wire[1084]) );
  DFF \memory_reg[33][27]  ( .D(n6701), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1083]), .Q(data_mem_out_wire[1083]) );
  DFF \memory_reg[33][26]  ( .D(n6700), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1082]), .Q(data_mem_out_wire[1082]) );
  DFF \memory_reg[33][25]  ( .D(n6699), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1081]), .Q(data_mem_out_wire[1081]) );
  DFF \memory_reg[33][24]  ( .D(n6698), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1080]), .Q(data_mem_out_wire[1080]) );
  DFF \memory_reg[33][23]  ( .D(n6697), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1079]), .Q(data_mem_out_wire[1079]) );
  DFF \memory_reg[33][22]  ( .D(n6696), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1078]), .Q(data_mem_out_wire[1078]) );
  DFF \memory_reg[33][21]  ( .D(n6695), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1077]), .Q(data_mem_out_wire[1077]) );
  DFF \memory_reg[33][20]  ( .D(n6694), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1076]), .Q(data_mem_out_wire[1076]) );
  DFF \memory_reg[33][19]  ( .D(n6693), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1075]), .Q(data_mem_out_wire[1075]) );
  DFF \memory_reg[33][18]  ( .D(n6692), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1074]), .Q(data_mem_out_wire[1074]) );
  DFF \memory_reg[33][17]  ( .D(n6691), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1073]), .Q(data_mem_out_wire[1073]) );
  DFF \memory_reg[33][16]  ( .D(n6690), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1072]), .Q(data_mem_out_wire[1072]) );
  DFF \memory_reg[33][15]  ( .D(n6689), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1071]), .Q(data_mem_out_wire[1071]) );
  DFF \memory_reg[33][14]  ( .D(n6688), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1070]), .Q(data_mem_out_wire[1070]) );
  DFF \memory_reg[33][13]  ( .D(n6687), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1069]), .Q(data_mem_out_wire[1069]) );
  DFF \memory_reg[33][12]  ( .D(n6686), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1068]), .Q(data_mem_out_wire[1068]) );
  DFF \memory_reg[33][11]  ( .D(n6685), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1067]), .Q(data_mem_out_wire[1067]) );
  DFF \memory_reg[33][10]  ( .D(n6684), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1066]), .Q(data_mem_out_wire[1066]) );
  DFF \memory_reg[33][9]  ( .D(n6683), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1065]), .Q(data_mem_out_wire[1065]) );
  DFF \memory_reg[33][8]  ( .D(n6682), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1064]), .Q(data_mem_out_wire[1064]) );
  DFF \memory_reg[33][7]  ( .D(n6681), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1063]), .Q(data_mem_out_wire[1063]) );
  DFF \memory_reg[33][6]  ( .D(n6680), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1062]), .Q(data_mem_out_wire[1062]) );
  DFF \memory_reg[33][5]  ( .D(n6679), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1061]), .Q(data_mem_out_wire[1061]) );
  DFF \memory_reg[33][4]  ( .D(n6678), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1060]), .Q(data_mem_out_wire[1060]) );
  DFF \memory_reg[33][3]  ( .D(n6677), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1059]), .Q(data_mem_out_wire[1059]) );
  DFF \memory_reg[33][2]  ( .D(n6676), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1058]), .Q(data_mem_out_wire[1058]) );
  DFF \memory_reg[33][1]  ( .D(n6675), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1057]), .Q(data_mem_out_wire[1057]) );
  DFF \memory_reg[33][0]  ( .D(n6674), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1056]), .Q(data_mem_out_wire[1056]) );
  DFF \memory_reg[34][31]  ( .D(n6673), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1119]), .Q(data_mem_out_wire[1119]) );
  DFF \memory_reg[34][30]  ( .D(n6672), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1118]), .Q(data_mem_out_wire[1118]) );
  DFF \memory_reg[34][29]  ( .D(n6671), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1117]), .Q(data_mem_out_wire[1117]) );
  DFF \memory_reg[34][28]  ( .D(n6670), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1116]), .Q(data_mem_out_wire[1116]) );
  DFF \memory_reg[34][27]  ( .D(n6669), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1115]), .Q(data_mem_out_wire[1115]) );
  DFF \memory_reg[34][26]  ( .D(n6668), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1114]), .Q(data_mem_out_wire[1114]) );
  DFF \memory_reg[34][25]  ( .D(n6667), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1113]), .Q(data_mem_out_wire[1113]) );
  DFF \memory_reg[34][24]  ( .D(n6666), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1112]), .Q(data_mem_out_wire[1112]) );
  DFF \memory_reg[34][23]  ( .D(n6665), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1111]), .Q(data_mem_out_wire[1111]) );
  DFF \memory_reg[34][22]  ( .D(n6664), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1110]), .Q(data_mem_out_wire[1110]) );
  DFF \memory_reg[34][21]  ( .D(n6663), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1109]), .Q(data_mem_out_wire[1109]) );
  DFF \memory_reg[34][20]  ( .D(n6662), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1108]), .Q(data_mem_out_wire[1108]) );
  DFF \memory_reg[34][19]  ( .D(n6661), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1107]), .Q(data_mem_out_wire[1107]) );
  DFF \memory_reg[34][18]  ( .D(n6660), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1106]), .Q(data_mem_out_wire[1106]) );
  DFF \memory_reg[34][17]  ( .D(n6659), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1105]), .Q(data_mem_out_wire[1105]) );
  DFF \memory_reg[34][16]  ( .D(n6658), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1104]), .Q(data_mem_out_wire[1104]) );
  DFF \memory_reg[34][15]  ( .D(n6657), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1103]), .Q(data_mem_out_wire[1103]) );
  DFF \memory_reg[34][14]  ( .D(n6656), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1102]), .Q(data_mem_out_wire[1102]) );
  DFF \memory_reg[34][13]  ( .D(n6655), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1101]), .Q(data_mem_out_wire[1101]) );
  DFF \memory_reg[34][12]  ( .D(n6654), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1100]), .Q(data_mem_out_wire[1100]) );
  DFF \memory_reg[34][11]  ( .D(n6653), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1099]), .Q(data_mem_out_wire[1099]) );
  DFF \memory_reg[34][10]  ( .D(n6652), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1098]), .Q(data_mem_out_wire[1098]) );
  DFF \memory_reg[34][9]  ( .D(n6651), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1097]), .Q(data_mem_out_wire[1097]) );
  DFF \memory_reg[34][8]  ( .D(n6650), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1096]), .Q(data_mem_out_wire[1096]) );
  DFF \memory_reg[34][7]  ( .D(n6649), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1095]), .Q(data_mem_out_wire[1095]) );
  DFF \memory_reg[34][6]  ( .D(n6648), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1094]), .Q(data_mem_out_wire[1094]) );
  DFF \memory_reg[34][5]  ( .D(n6647), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1093]), .Q(data_mem_out_wire[1093]) );
  DFF \memory_reg[34][4]  ( .D(n6646), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1092]), .Q(data_mem_out_wire[1092]) );
  DFF \memory_reg[34][3]  ( .D(n6645), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1091]), .Q(data_mem_out_wire[1091]) );
  DFF \memory_reg[34][2]  ( .D(n6644), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1090]), .Q(data_mem_out_wire[1090]) );
  DFF \memory_reg[34][1]  ( .D(n6643), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1089]), .Q(data_mem_out_wire[1089]) );
  DFF \memory_reg[34][0]  ( .D(n6642), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1088]), .Q(data_mem_out_wire[1088]) );
  DFF \memory_reg[35][31]  ( .D(n6641), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1151]), .Q(data_mem_out_wire[1151]) );
  DFF \memory_reg[35][30]  ( .D(n6640), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1150]), .Q(data_mem_out_wire[1150]) );
  DFF \memory_reg[35][29]  ( .D(n6639), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1149]), .Q(data_mem_out_wire[1149]) );
  DFF \memory_reg[35][28]  ( .D(n6638), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1148]), .Q(data_mem_out_wire[1148]) );
  DFF \memory_reg[35][27]  ( .D(n6637), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1147]), .Q(data_mem_out_wire[1147]) );
  DFF \memory_reg[35][26]  ( .D(n6636), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1146]), .Q(data_mem_out_wire[1146]) );
  DFF \memory_reg[35][25]  ( .D(n6635), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1145]), .Q(data_mem_out_wire[1145]) );
  DFF \memory_reg[35][24]  ( .D(n6634), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1144]), .Q(data_mem_out_wire[1144]) );
  DFF \memory_reg[35][23]  ( .D(n6633), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1143]), .Q(data_mem_out_wire[1143]) );
  DFF \memory_reg[35][22]  ( .D(n6632), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1142]), .Q(data_mem_out_wire[1142]) );
  DFF \memory_reg[35][21]  ( .D(n6631), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1141]), .Q(data_mem_out_wire[1141]) );
  DFF \memory_reg[35][20]  ( .D(n6630), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1140]), .Q(data_mem_out_wire[1140]) );
  DFF \memory_reg[35][19]  ( .D(n6629), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1139]), .Q(data_mem_out_wire[1139]) );
  DFF \memory_reg[35][18]  ( .D(n6628), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1138]), .Q(data_mem_out_wire[1138]) );
  DFF \memory_reg[35][17]  ( .D(n6627), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1137]), .Q(data_mem_out_wire[1137]) );
  DFF \memory_reg[35][16]  ( .D(n6626), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1136]), .Q(data_mem_out_wire[1136]) );
  DFF \memory_reg[35][15]  ( .D(n6625), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1135]), .Q(data_mem_out_wire[1135]) );
  DFF \memory_reg[35][14]  ( .D(n6624), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1134]), .Q(data_mem_out_wire[1134]) );
  DFF \memory_reg[35][13]  ( .D(n6623), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1133]), .Q(data_mem_out_wire[1133]) );
  DFF \memory_reg[35][12]  ( .D(n6622), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1132]), .Q(data_mem_out_wire[1132]) );
  DFF \memory_reg[35][11]  ( .D(n6621), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1131]), .Q(data_mem_out_wire[1131]) );
  DFF \memory_reg[35][10]  ( .D(n6620), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1130]), .Q(data_mem_out_wire[1130]) );
  DFF \memory_reg[35][9]  ( .D(n6619), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1129]), .Q(data_mem_out_wire[1129]) );
  DFF \memory_reg[35][8]  ( .D(n6618), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1128]), .Q(data_mem_out_wire[1128]) );
  DFF \memory_reg[35][7]  ( .D(n6617), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1127]), .Q(data_mem_out_wire[1127]) );
  DFF \memory_reg[35][6]  ( .D(n6616), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1126]), .Q(data_mem_out_wire[1126]) );
  DFF \memory_reg[35][5]  ( .D(n6615), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1125]), .Q(data_mem_out_wire[1125]) );
  DFF \memory_reg[35][4]  ( .D(n6614), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1124]), .Q(data_mem_out_wire[1124]) );
  DFF \memory_reg[35][3]  ( .D(n6613), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1123]), .Q(data_mem_out_wire[1123]) );
  DFF \memory_reg[35][2]  ( .D(n6612), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1122]), .Q(data_mem_out_wire[1122]) );
  DFF \memory_reg[35][1]  ( .D(n6611), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1121]), .Q(data_mem_out_wire[1121]) );
  DFF \memory_reg[35][0]  ( .D(n6610), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1120]), .Q(data_mem_out_wire[1120]) );
  DFF \memory_reg[36][31]  ( .D(n6609), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1183]), .Q(data_mem_out_wire[1183]) );
  DFF \memory_reg[36][30]  ( .D(n6608), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1182]), .Q(data_mem_out_wire[1182]) );
  DFF \memory_reg[36][29]  ( .D(n6607), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1181]), .Q(data_mem_out_wire[1181]) );
  DFF \memory_reg[36][28]  ( .D(n6606), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1180]), .Q(data_mem_out_wire[1180]) );
  DFF \memory_reg[36][27]  ( .D(n6605), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1179]), .Q(data_mem_out_wire[1179]) );
  DFF \memory_reg[36][26]  ( .D(n6604), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1178]), .Q(data_mem_out_wire[1178]) );
  DFF \memory_reg[36][25]  ( .D(n6603), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1177]), .Q(data_mem_out_wire[1177]) );
  DFF \memory_reg[36][24]  ( .D(n6602), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1176]), .Q(data_mem_out_wire[1176]) );
  DFF \memory_reg[36][23]  ( .D(n6601), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1175]), .Q(data_mem_out_wire[1175]) );
  DFF \memory_reg[36][22]  ( .D(n6600), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1174]), .Q(data_mem_out_wire[1174]) );
  DFF \memory_reg[36][21]  ( .D(n6599), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1173]), .Q(data_mem_out_wire[1173]) );
  DFF \memory_reg[36][20]  ( .D(n6598), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1172]), .Q(data_mem_out_wire[1172]) );
  DFF \memory_reg[36][19]  ( .D(n6597), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1171]), .Q(data_mem_out_wire[1171]) );
  DFF \memory_reg[36][18]  ( .D(n6596), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1170]), .Q(data_mem_out_wire[1170]) );
  DFF \memory_reg[36][17]  ( .D(n6595), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1169]), .Q(data_mem_out_wire[1169]) );
  DFF \memory_reg[36][16]  ( .D(n6594), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1168]), .Q(data_mem_out_wire[1168]) );
  DFF \memory_reg[36][15]  ( .D(n6593), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1167]), .Q(data_mem_out_wire[1167]) );
  DFF \memory_reg[36][14]  ( .D(n6592), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1166]), .Q(data_mem_out_wire[1166]) );
  DFF \memory_reg[36][13]  ( .D(n6591), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1165]), .Q(data_mem_out_wire[1165]) );
  DFF \memory_reg[36][12]  ( .D(n6590), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1164]), .Q(data_mem_out_wire[1164]) );
  DFF \memory_reg[36][11]  ( .D(n6589), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1163]), .Q(data_mem_out_wire[1163]) );
  DFF \memory_reg[36][10]  ( .D(n6588), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1162]), .Q(data_mem_out_wire[1162]) );
  DFF \memory_reg[36][9]  ( .D(n6587), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1161]), .Q(data_mem_out_wire[1161]) );
  DFF \memory_reg[36][8]  ( .D(n6586), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1160]), .Q(data_mem_out_wire[1160]) );
  DFF \memory_reg[36][7]  ( .D(n6585), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1159]), .Q(data_mem_out_wire[1159]) );
  DFF \memory_reg[36][6]  ( .D(n6584), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1158]), .Q(data_mem_out_wire[1158]) );
  DFF \memory_reg[36][5]  ( .D(n6583), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1157]), .Q(data_mem_out_wire[1157]) );
  DFF \memory_reg[36][4]  ( .D(n6582), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1156]), .Q(data_mem_out_wire[1156]) );
  DFF \memory_reg[36][3]  ( .D(n6581), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1155]), .Q(data_mem_out_wire[1155]) );
  DFF \memory_reg[36][2]  ( .D(n6580), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1154]), .Q(data_mem_out_wire[1154]) );
  DFF \memory_reg[36][1]  ( .D(n6579), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1153]), .Q(data_mem_out_wire[1153]) );
  DFF \memory_reg[36][0]  ( .D(n6578), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1152]), .Q(data_mem_out_wire[1152]) );
  DFF \memory_reg[37][31]  ( .D(n6577), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1215]), .Q(data_mem_out_wire[1215]) );
  DFF \memory_reg[37][30]  ( .D(n6576), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1214]), .Q(data_mem_out_wire[1214]) );
  DFF \memory_reg[37][29]  ( .D(n6575), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1213]), .Q(data_mem_out_wire[1213]) );
  DFF \memory_reg[37][28]  ( .D(n6574), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1212]), .Q(data_mem_out_wire[1212]) );
  DFF \memory_reg[37][27]  ( .D(n6573), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1211]), .Q(data_mem_out_wire[1211]) );
  DFF \memory_reg[37][26]  ( .D(n6572), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1210]), .Q(data_mem_out_wire[1210]) );
  DFF \memory_reg[37][25]  ( .D(n6571), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1209]), .Q(data_mem_out_wire[1209]) );
  DFF \memory_reg[37][24]  ( .D(n6570), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1208]), .Q(data_mem_out_wire[1208]) );
  DFF \memory_reg[37][23]  ( .D(n6569), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1207]), .Q(data_mem_out_wire[1207]) );
  DFF \memory_reg[37][22]  ( .D(n6568), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1206]), .Q(data_mem_out_wire[1206]) );
  DFF \memory_reg[37][21]  ( .D(n6567), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1205]), .Q(data_mem_out_wire[1205]) );
  DFF \memory_reg[37][20]  ( .D(n6566), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1204]), .Q(data_mem_out_wire[1204]) );
  DFF \memory_reg[37][19]  ( .D(n6565), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1203]), .Q(data_mem_out_wire[1203]) );
  DFF \memory_reg[37][18]  ( .D(n6564), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1202]), .Q(data_mem_out_wire[1202]) );
  DFF \memory_reg[37][17]  ( .D(n6563), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1201]), .Q(data_mem_out_wire[1201]) );
  DFF \memory_reg[37][16]  ( .D(n6562), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1200]), .Q(data_mem_out_wire[1200]) );
  DFF \memory_reg[37][15]  ( .D(n6561), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1199]), .Q(data_mem_out_wire[1199]) );
  DFF \memory_reg[37][14]  ( .D(n6560), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1198]), .Q(data_mem_out_wire[1198]) );
  DFF \memory_reg[37][13]  ( .D(n6559), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1197]), .Q(data_mem_out_wire[1197]) );
  DFF \memory_reg[37][12]  ( .D(n6558), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1196]), .Q(data_mem_out_wire[1196]) );
  DFF \memory_reg[37][11]  ( .D(n6557), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1195]), .Q(data_mem_out_wire[1195]) );
  DFF \memory_reg[37][10]  ( .D(n6556), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1194]), .Q(data_mem_out_wire[1194]) );
  DFF \memory_reg[37][9]  ( .D(n6555), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1193]), .Q(data_mem_out_wire[1193]) );
  DFF \memory_reg[37][8]  ( .D(n6554), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1192]), .Q(data_mem_out_wire[1192]) );
  DFF \memory_reg[37][7]  ( .D(n6553), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1191]), .Q(data_mem_out_wire[1191]) );
  DFF \memory_reg[37][6]  ( .D(n6552), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1190]), .Q(data_mem_out_wire[1190]) );
  DFF \memory_reg[37][5]  ( .D(n6551), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1189]), .Q(data_mem_out_wire[1189]) );
  DFF \memory_reg[37][4]  ( .D(n6550), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1188]), .Q(data_mem_out_wire[1188]) );
  DFF \memory_reg[37][3]  ( .D(n6549), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1187]), .Q(data_mem_out_wire[1187]) );
  DFF \memory_reg[37][2]  ( .D(n6548), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1186]), .Q(data_mem_out_wire[1186]) );
  DFF \memory_reg[37][1]  ( .D(n6547), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1185]), .Q(data_mem_out_wire[1185]) );
  DFF \memory_reg[37][0]  ( .D(n6546), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1184]), .Q(data_mem_out_wire[1184]) );
  DFF \memory_reg[38][31]  ( .D(n6545), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1247]), .Q(data_mem_out_wire[1247]) );
  DFF \memory_reg[38][30]  ( .D(n6544), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1246]), .Q(data_mem_out_wire[1246]) );
  DFF \memory_reg[38][29]  ( .D(n6543), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1245]), .Q(data_mem_out_wire[1245]) );
  DFF \memory_reg[38][28]  ( .D(n6542), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1244]), .Q(data_mem_out_wire[1244]) );
  DFF \memory_reg[38][27]  ( .D(n6541), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1243]), .Q(data_mem_out_wire[1243]) );
  DFF \memory_reg[38][26]  ( .D(n6540), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1242]), .Q(data_mem_out_wire[1242]) );
  DFF \memory_reg[38][25]  ( .D(n6539), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1241]), .Q(data_mem_out_wire[1241]) );
  DFF \memory_reg[38][24]  ( .D(n6538), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1240]), .Q(data_mem_out_wire[1240]) );
  DFF \memory_reg[38][23]  ( .D(n6537), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1239]), .Q(data_mem_out_wire[1239]) );
  DFF \memory_reg[38][22]  ( .D(n6536), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1238]), .Q(data_mem_out_wire[1238]) );
  DFF \memory_reg[38][21]  ( .D(n6535), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1237]), .Q(data_mem_out_wire[1237]) );
  DFF \memory_reg[38][20]  ( .D(n6534), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1236]), .Q(data_mem_out_wire[1236]) );
  DFF \memory_reg[38][19]  ( .D(n6533), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1235]), .Q(data_mem_out_wire[1235]) );
  DFF \memory_reg[38][18]  ( .D(n6532), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1234]), .Q(data_mem_out_wire[1234]) );
  DFF \memory_reg[38][17]  ( .D(n6531), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1233]), .Q(data_mem_out_wire[1233]) );
  DFF \memory_reg[38][16]  ( .D(n6530), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1232]), .Q(data_mem_out_wire[1232]) );
  DFF \memory_reg[38][15]  ( .D(n6529), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1231]), .Q(data_mem_out_wire[1231]) );
  DFF \memory_reg[38][14]  ( .D(n6528), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1230]), .Q(data_mem_out_wire[1230]) );
  DFF \memory_reg[38][13]  ( .D(n6527), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1229]), .Q(data_mem_out_wire[1229]) );
  DFF \memory_reg[38][12]  ( .D(n6526), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1228]), .Q(data_mem_out_wire[1228]) );
  DFF \memory_reg[38][11]  ( .D(n6525), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1227]), .Q(data_mem_out_wire[1227]) );
  DFF \memory_reg[38][10]  ( .D(n6524), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1226]), .Q(data_mem_out_wire[1226]) );
  DFF \memory_reg[38][9]  ( .D(n6523), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1225]), .Q(data_mem_out_wire[1225]) );
  DFF \memory_reg[38][8]  ( .D(n6522), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1224]), .Q(data_mem_out_wire[1224]) );
  DFF \memory_reg[38][7]  ( .D(n6521), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1223]), .Q(data_mem_out_wire[1223]) );
  DFF \memory_reg[38][6]  ( .D(n6520), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1222]), .Q(data_mem_out_wire[1222]) );
  DFF \memory_reg[38][5]  ( .D(n6519), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1221]), .Q(data_mem_out_wire[1221]) );
  DFF \memory_reg[38][4]  ( .D(n6518), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1220]), .Q(data_mem_out_wire[1220]) );
  DFF \memory_reg[38][3]  ( .D(n6517), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1219]), .Q(data_mem_out_wire[1219]) );
  DFF \memory_reg[38][2]  ( .D(n6516), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1218]), .Q(data_mem_out_wire[1218]) );
  DFF \memory_reg[38][1]  ( .D(n6515), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1217]), .Q(data_mem_out_wire[1217]) );
  DFF \memory_reg[38][0]  ( .D(n6514), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1216]), .Q(data_mem_out_wire[1216]) );
  DFF \memory_reg[39][31]  ( .D(n6513), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1279]), .Q(data_mem_out_wire[1279]) );
  DFF \memory_reg[39][30]  ( .D(n6512), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1278]), .Q(data_mem_out_wire[1278]) );
  DFF \memory_reg[39][29]  ( .D(n6511), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1277]), .Q(data_mem_out_wire[1277]) );
  DFF \memory_reg[39][28]  ( .D(n6510), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1276]), .Q(data_mem_out_wire[1276]) );
  DFF \memory_reg[39][27]  ( .D(n6509), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1275]), .Q(data_mem_out_wire[1275]) );
  DFF \memory_reg[39][26]  ( .D(n6508), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1274]), .Q(data_mem_out_wire[1274]) );
  DFF \memory_reg[39][25]  ( .D(n6507), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1273]), .Q(data_mem_out_wire[1273]) );
  DFF \memory_reg[39][24]  ( .D(n6506), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1272]), .Q(data_mem_out_wire[1272]) );
  DFF \memory_reg[39][23]  ( .D(n6505), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1271]), .Q(data_mem_out_wire[1271]) );
  DFF \memory_reg[39][22]  ( .D(n6504), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1270]), .Q(data_mem_out_wire[1270]) );
  DFF \memory_reg[39][21]  ( .D(n6503), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1269]), .Q(data_mem_out_wire[1269]) );
  DFF \memory_reg[39][20]  ( .D(n6502), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1268]), .Q(data_mem_out_wire[1268]) );
  DFF \memory_reg[39][19]  ( .D(n6501), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1267]), .Q(data_mem_out_wire[1267]) );
  DFF \memory_reg[39][18]  ( .D(n6500), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1266]), .Q(data_mem_out_wire[1266]) );
  DFF \memory_reg[39][17]  ( .D(n6499), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1265]), .Q(data_mem_out_wire[1265]) );
  DFF \memory_reg[39][16]  ( .D(n6498), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1264]), .Q(data_mem_out_wire[1264]) );
  DFF \memory_reg[39][15]  ( .D(n6497), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1263]), .Q(data_mem_out_wire[1263]) );
  DFF \memory_reg[39][14]  ( .D(n6496), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1262]), .Q(data_mem_out_wire[1262]) );
  DFF \memory_reg[39][13]  ( .D(n6495), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1261]), .Q(data_mem_out_wire[1261]) );
  DFF \memory_reg[39][12]  ( .D(n6494), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1260]), .Q(data_mem_out_wire[1260]) );
  DFF \memory_reg[39][11]  ( .D(n6493), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1259]), .Q(data_mem_out_wire[1259]) );
  DFF \memory_reg[39][10]  ( .D(n6492), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1258]), .Q(data_mem_out_wire[1258]) );
  DFF \memory_reg[39][9]  ( .D(n6491), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1257]), .Q(data_mem_out_wire[1257]) );
  DFF \memory_reg[39][8]  ( .D(n6490), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1256]), .Q(data_mem_out_wire[1256]) );
  DFF \memory_reg[39][7]  ( .D(n6489), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1255]), .Q(data_mem_out_wire[1255]) );
  DFF \memory_reg[39][6]  ( .D(n6488), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1254]), .Q(data_mem_out_wire[1254]) );
  DFF \memory_reg[39][5]  ( .D(n6487), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1253]), .Q(data_mem_out_wire[1253]) );
  DFF \memory_reg[39][4]  ( .D(n6486), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1252]), .Q(data_mem_out_wire[1252]) );
  DFF \memory_reg[39][3]  ( .D(n6485), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1251]), .Q(data_mem_out_wire[1251]) );
  DFF \memory_reg[39][2]  ( .D(n6484), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1250]), .Q(data_mem_out_wire[1250]) );
  DFF \memory_reg[39][1]  ( .D(n6483), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1249]), .Q(data_mem_out_wire[1249]) );
  DFF \memory_reg[39][0]  ( .D(n6482), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1248]), .Q(data_mem_out_wire[1248]) );
  DFF \memory_reg[40][31]  ( .D(n6481), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1311]), .Q(data_mem_out_wire[1311]) );
  DFF \memory_reg[40][30]  ( .D(n6480), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1310]), .Q(data_mem_out_wire[1310]) );
  DFF \memory_reg[40][29]  ( .D(n6479), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1309]), .Q(data_mem_out_wire[1309]) );
  DFF \memory_reg[40][28]  ( .D(n6478), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1308]), .Q(data_mem_out_wire[1308]) );
  DFF \memory_reg[40][27]  ( .D(n6477), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1307]), .Q(data_mem_out_wire[1307]) );
  DFF \memory_reg[40][26]  ( .D(n6476), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1306]), .Q(data_mem_out_wire[1306]) );
  DFF \memory_reg[40][25]  ( .D(n6475), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1305]), .Q(data_mem_out_wire[1305]) );
  DFF \memory_reg[40][24]  ( .D(n6474), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1304]), .Q(data_mem_out_wire[1304]) );
  DFF \memory_reg[40][23]  ( .D(n6473), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1303]), .Q(data_mem_out_wire[1303]) );
  DFF \memory_reg[40][22]  ( .D(n6472), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1302]), .Q(data_mem_out_wire[1302]) );
  DFF \memory_reg[40][21]  ( .D(n6471), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1301]), .Q(data_mem_out_wire[1301]) );
  DFF \memory_reg[40][20]  ( .D(n6470), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1300]), .Q(data_mem_out_wire[1300]) );
  DFF \memory_reg[40][19]  ( .D(n6469), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1299]), .Q(data_mem_out_wire[1299]) );
  DFF \memory_reg[40][18]  ( .D(n6468), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1298]), .Q(data_mem_out_wire[1298]) );
  DFF \memory_reg[40][17]  ( .D(n6467), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1297]), .Q(data_mem_out_wire[1297]) );
  DFF \memory_reg[40][16]  ( .D(n6466), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1296]), .Q(data_mem_out_wire[1296]) );
  DFF \memory_reg[40][15]  ( .D(n6465), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1295]), .Q(data_mem_out_wire[1295]) );
  DFF \memory_reg[40][14]  ( .D(n6464), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1294]), .Q(data_mem_out_wire[1294]) );
  DFF \memory_reg[40][13]  ( .D(n6463), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1293]), .Q(data_mem_out_wire[1293]) );
  DFF \memory_reg[40][12]  ( .D(n6462), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1292]), .Q(data_mem_out_wire[1292]) );
  DFF \memory_reg[40][11]  ( .D(n6461), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1291]), .Q(data_mem_out_wire[1291]) );
  DFF \memory_reg[40][10]  ( .D(n6460), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1290]), .Q(data_mem_out_wire[1290]) );
  DFF \memory_reg[40][9]  ( .D(n6459), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1289]), .Q(data_mem_out_wire[1289]) );
  DFF \memory_reg[40][8]  ( .D(n6458), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1288]), .Q(data_mem_out_wire[1288]) );
  DFF \memory_reg[40][7]  ( .D(n6457), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1287]), .Q(data_mem_out_wire[1287]) );
  DFF \memory_reg[40][6]  ( .D(n6456), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1286]), .Q(data_mem_out_wire[1286]) );
  DFF \memory_reg[40][5]  ( .D(n6455), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1285]), .Q(data_mem_out_wire[1285]) );
  DFF \memory_reg[40][4]  ( .D(n6454), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1284]), .Q(data_mem_out_wire[1284]) );
  DFF \memory_reg[40][3]  ( .D(n6453), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1283]), .Q(data_mem_out_wire[1283]) );
  DFF \memory_reg[40][2]  ( .D(n6452), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1282]), .Q(data_mem_out_wire[1282]) );
  DFF \memory_reg[40][1]  ( .D(n6451), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1281]), .Q(data_mem_out_wire[1281]) );
  DFF \memory_reg[40][0]  ( .D(n6450), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1280]), .Q(data_mem_out_wire[1280]) );
  DFF \memory_reg[41][31]  ( .D(n6449), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1343]), .Q(data_mem_out_wire[1343]) );
  DFF \memory_reg[41][30]  ( .D(n6448), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1342]), .Q(data_mem_out_wire[1342]) );
  DFF \memory_reg[41][29]  ( .D(n6447), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1341]), .Q(data_mem_out_wire[1341]) );
  DFF \memory_reg[41][28]  ( .D(n6446), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1340]), .Q(data_mem_out_wire[1340]) );
  DFF \memory_reg[41][27]  ( .D(n6445), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1339]), .Q(data_mem_out_wire[1339]) );
  DFF \memory_reg[41][26]  ( .D(n6444), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1338]), .Q(data_mem_out_wire[1338]) );
  DFF \memory_reg[41][25]  ( .D(n6443), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1337]), .Q(data_mem_out_wire[1337]) );
  DFF \memory_reg[41][24]  ( .D(n6442), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1336]), .Q(data_mem_out_wire[1336]) );
  DFF \memory_reg[41][23]  ( .D(n6441), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1335]), .Q(data_mem_out_wire[1335]) );
  DFF \memory_reg[41][22]  ( .D(n6440), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1334]), .Q(data_mem_out_wire[1334]) );
  DFF \memory_reg[41][21]  ( .D(n6439), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1333]), .Q(data_mem_out_wire[1333]) );
  DFF \memory_reg[41][20]  ( .D(n6438), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1332]), .Q(data_mem_out_wire[1332]) );
  DFF \memory_reg[41][19]  ( .D(n6437), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1331]), .Q(data_mem_out_wire[1331]) );
  DFF \memory_reg[41][18]  ( .D(n6436), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1330]), .Q(data_mem_out_wire[1330]) );
  DFF \memory_reg[41][17]  ( .D(n6435), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1329]), .Q(data_mem_out_wire[1329]) );
  DFF \memory_reg[41][16]  ( .D(n6434), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1328]), .Q(data_mem_out_wire[1328]) );
  DFF \memory_reg[41][15]  ( .D(n6433), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1327]), .Q(data_mem_out_wire[1327]) );
  DFF \memory_reg[41][14]  ( .D(n6432), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1326]), .Q(data_mem_out_wire[1326]) );
  DFF \memory_reg[41][13]  ( .D(n6431), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1325]), .Q(data_mem_out_wire[1325]) );
  DFF \memory_reg[41][12]  ( .D(n6430), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1324]), .Q(data_mem_out_wire[1324]) );
  DFF \memory_reg[41][11]  ( .D(n6429), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1323]), .Q(data_mem_out_wire[1323]) );
  DFF \memory_reg[41][10]  ( .D(n6428), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1322]), .Q(data_mem_out_wire[1322]) );
  DFF \memory_reg[41][9]  ( .D(n6427), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1321]), .Q(data_mem_out_wire[1321]) );
  DFF \memory_reg[41][8]  ( .D(n6426), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1320]), .Q(data_mem_out_wire[1320]) );
  DFF \memory_reg[41][7]  ( .D(n6425), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1319]), .Q(data_mem_out_wire[1319]) );
  DFF \memory_reg[41][6]  ( .D(n6424), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1318]), .Q(data_mem_out_wire[1318]) );
  DFF \memory_reg[41][5]  ( .D(n6423), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1317]), .Q(data_mem_out_wire[1317]) );
  DFF \memory_reg[41][4]  ( .D(n6422), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1316]), .Q(data_mem_out_wire[1316]) );
  DFF \memory_reg[41][3]  ( .D(n6421), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1315]), .Q(data_mem_out_wire[1315]) );
  DFF \memory_reg[41][2]  ( .D(n6420), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1314]), .Q(data_mem_out_wire[1314]) );
  DFF \memory_reg[41][1]  ( .D(n6419), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1313]), .Q(data_mem_out_wire[1313]) );
  DFF \memory_reg[41][0]  ( .D(n6418), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1312]), .Q(data_mem_out_wire[1312]) );
  DFF \memory_reg[42][31]  ( .D(n6417), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1375]), .Q(data_mem_out_wire[1375]) );
  DFF \memory_reg[42][30]  ( .D(n6416), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1374]), .Q(data_mem_out_wire[1374]) );
  DFF \memory_reg[42][29]  ( .D(n6415), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1373]), .Q(data_mem_out_wire[1373]) );
  DFF \memory_reg[42][28]  ( .D(n6414), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1372]), .Q(data_mem_out_wire[1372]) );
  DFF \memory_reg[42][27]  ( .D(n6413), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1371]), .Q(data_mem_out_wire[1371]) );
  DFF \memory_reg[42][26]  ( .D(n6412), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1370]), .Q(data_mem_out_wire[1370]) );
  DFF \memory_reg[42][25]  ( .D(n6411), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1369]), .Q(data_mem_out_wire[1369]) );
  DFF \memory_reg[42][24]  ( .D(n6410), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1368]), .Q(data_mem_out_wire[1368]) );
  DFF \memory_reg[42][23]  ( .D(n6409), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1367]), .Q(data_mem_out_wire[1367]) );
  DFF \memory_reg[42][22]  ( .D(n6408), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1366]), .Q(data_mem_out_wire[1366]) );
  DFF \memory_reg[42][21]  ( .D(n6407), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1365]), .Q(data_mem_out_wire[1365]) );
  DFF \memory_reg[42][20]  ( .D(n6406), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1364]), .Q(data_mem_out_wire[1364]) );
  DFF \memory_reg[42][19]  ( .D(n6405), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1363]), .Q(data_mem_out_wire[1363]) );
  DFF \memory_reg[42][18]  ( .D(n6404), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1362]), .Q(data_mem_out_wire[1362]) );
  DFF \memory_reg[42][17]  ( .D(n6403), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1361]), .Q(data_mem_out_wire[1361]) );
  DFF \memory_reg[42][16]  ( .D(n6402), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1360]), .Q(data_mem_out_wire[1360]) );
  DFF \memory_reg[42][15]  ( .D(n6401), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1359]), .Q(data_mem_out_wire[1359]) );
  DFF \memory_reg[42][14]  ( .D(n6400), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1358]), .Q(data_mem_out_wire[1358]) );
  DFF \memory_reg[42][13]  ( .D(n6399), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1357]), .Q(data_mem_out_wire[1357]) );
  DFF \memory_reg[42][12]  ( .D(n6398), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1356]), .Q(data_mem_out_wire[1356]) );
  DFF \memory_reg[42][11]  ( .D(n6397), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1355]), .Q(data_mem_out_wire[1355]) );
  DFF \memory_reg[42][10]  ( .D(n6396), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1354]), .Q(data_mem_out_wire[1354]) );
  DFF \memory_reg[42][9]  ( .D(n6395), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1353]), .Q(data_mem_out_wire[1353]) );
  DFF \memory_reg[42][8]  ( .D(n6394), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1352]), .Q(data_mem_out_wire[1352]) );
  DFF \memory_reg[42][7]  ( .D(n6393), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1351]), .Q(data_mem_out_wire[1351]) );
  DFF \memory_reg[42][6]  ( .D(n6392), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1350]), .Q(data_mem_out_wire[1350]) );
  DFF \memory_reg[42][5]  ( .D(n6391), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1349]), .Q(data_mem_out_wire[1349]) );
  DFF \memory_reg[42][4]  ( .D(n6390), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1348]), .Q(data_mem_out_wire[1348]) );
  DFF \memory_reg[42][3]  ( .D(n6389), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1347]), .Q(data_mem_out_wire[1347]) );
  DFF \memory_reg[42][2]  ( .D(n6388), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1346]), .Q(data_mem_out_wire[1346]) );
  DFF \memory_reg[42][1]  ( .D(n6387), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1345]), .Q(data_mem_out_wire[1345]) );
  DFF \memory_reg[42][0]  ( .D(n6386), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1344]), .Q(data_mem_out_wire[1344]) );
  DFF \memory_reg[43][31]  ( .D(n6385), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1407]), .Q(data_mem_out_wire[1407]) );
  DFF \memory_reg[43][30]  ( .D(n6384), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1406]), .Q(data_mem_out_wire[1406]) );
  DFF \memory_reg[43][29]  ( .D(n6383), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1405]), .Q(data_mem_out_wire[1405]) );
  DFF \memory_reg[43][28]  ( .D(n6382), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1404]), .Q(data_mem_out_wire[1404]) );
  DFF \memory_reg[43][27]  ( .D(n6381), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1403]), .Q(data_mem_out_wire[1403]) );
  DFF \memory_reg[43][26]  ( .D(n6380), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1402]), .Q(data_mem_out_wire[1402]) );
  DFF \memory_reg[43][25]  ( .D(n6379), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1401]), .Q(data_mem_out_wire[1401]) );
  DFF \memory_reg[43][24]  ( .D(n6378), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1400]), .Q(data_mem_out_wire[1400]) );
  DFF \memory_reg[43][23]  ( .D(n6377), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1399]), .Q(data_mem_out_wire[1399]) );
  DFF \memory_reg[43][22]  ( .D(n6376), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1398]), .Q(data_mem_out_wire[1398]) );
  DFF \memory_reg[43][21]  ( .D(n6375), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1397]), .Q(data_mem_out_wire[1397]) );
  DFF \memory_reg[43][20]  ( .D(n6374), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1396]), .Q(data_mem_out_wire[1396]) );
  DFF \memory_reg[43][19]  ( .D(n6373), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1395]), .Q(data_mem_out_wire[1395]) );
  DFF \memory_reg[43][18]  ( .D(n6372), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1394]), .Q(data_mem_out_wire[1394]) );
  DFF \memory_reg[43][17]  ( .D(n6371), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1393]), .Q(data_mem_out_wire[1393]) );
  DFF \memory_reg[43][16]  ( .D(n6370), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1392]), .Q(data_mem_out_wire[1392]) );
  DFF \memory_reg[43][15]  ( .D(n6369), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1391]), .Q(data_mem_out_wire[1391]) );
  DFF \memory_reg[43][14]  ( .D(n6368), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1390]), .Q(data_mem_out_wire[1390]) );
  DFF \memory_reg[43][13]  ( .D(n6367), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1389]), .Q(data_mem_out_wire[1389]) );
  DFF \memory_reg[43][12]  ( .D(n6366), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1388]), .Q(data_mem_out_wire[1388]) );
  DFF \memory_reg[43][11]  ( .D(n6365), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1387]), .Q(data_mem_out_wire[1387]) );
  DFF \memory_reg[43][10]  ( .D(n6364), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1386]), .Q(data_mem_out_wire[1386]) );
  DFF \memory_reg[43][9]  ( .D(n6363), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1385]), .Q(data_mem_out_wire[1385]) );
  DFF \memory_reg[43][8]  ( .D(n6362), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1384]), .Q(data_mem_out_wire[1384]) );
  DFF \memory_reg[43][7]  ( .D(n6361), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1383]), .Q(data_mem_out_wire[1383]) );
  DFF \memory_reg[43][6]  ( .D(n6360), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1382]), .Q(data_mem_out_wire[1382]) );
  DFF \memory_reg[43][5]  ( .D(n6359), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1381]), .Q(data_mem_out_wire[1381]) );
  DFF \memory_reg[43][4]  ( .D(n6358), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1380]), .Q(data_mem_out_wire[1380]) );
  DFF \memory_reg[43][3]  ( .D(n6357), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1379]), .Q(data_mem_out_wire[1379]) );
  DFF \memory_reg[43][2]  ( .D(n6356), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1378]), .Q(data_mem_out_wire[1378]) );
  DFF \memory_reg[43][1]  ( .D(n6355), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1377]), .Q(data_mem_out_wire[1377]) );
  DFF \memory_reg[43][0]  ( .D(n6354), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1376]), .Q(data_mem_out_wire[1376]) );
  DFF \memory_reg[44][31]  ( .D(n6353), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1439]), .Q(data_mem_out_wire[1439]) );
  DFF \memory_reg[44][30]  ( .D(n6352), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1438]), .Q(data_mem_out_wire[1438]) );
  DFF \memory_reg[44][29]  ( .D(n6351), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1437]), .Q(data_mem_out_wire[1437]) );
  DFF \memory_reg[44][28]  ( .D(n6350), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1436]), .Q(data_mem_out_wire[1436]) );
  DFF \memory_reg[44][27]  ( .D(n6349), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1435]), .Q(data_mem_out_wire[1435]) );
  DFF \memory_reg[44][26]  ( .D(n6348), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1434]), .Q(data_mem_out_wire[1434]) );
  DFF \memory_reg[44][25]  ( .D(n6347), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1433]), .Q(data_mem_out_wire[1433]) );
  DFF \memory_reg[44][24]  ( .D(n6346), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1432]), .Q(data_mem_out_wire[1432]) );
  DFF \memory_reg[44][23]  ( .D(n6345), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1431]), .Q(data_mem_out_wire[1431]) );
  DFF \memory_reg[44][22]  ( .D(n6344), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1430]), .Q(data_mem_out_wire[1430]) );
  DFF \memory_reg[44][21]  ( .D(n6343), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1429]), .Q(data_mem_out_wire[1429]) );
  DFF \memory_reg[44][20]  ( .D(n6342), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1428]), .Q(data_mem_out_wire[1428]) );
  DFF \memory_reg[44][19]  ( .D(n6341), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1427]), .Q(data_mem_out_wire[1427]) );
  DFF \memory_reg[44][18]  ( .D(n6340), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1426]), .Q(data_mem_out_wire[1426]) );
  DFF \memory_reg[44][17]  ( .D(n6339), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1425]), .Q(data_mem_out_wire[1425]) );
  DFF \memory_reg[44][16]  ( .D(n6338), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1424]), .Q(data_mem_out_wire[1424]) );
  DFF \memory_reg[44][15]  ( .D(n6337), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1423]), .Q(data_mem_out_wire[1423]) );
  DFF \memory_reg[44][14]  ( .D(n6336), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1422]), .Q(data_mem_out_wire[1422]) );
  DFF \memory_reg[44][13]  ( .D(n6335), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1421]), .Q(data_mem_out_wire[1421]) );
  DFF \memory_reg[44][12]  ( .D(n6334), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1420]), .Q(data_mem_out_wire[1420]) );
  DFF \memory_reg[44][11]  ( .D(n6333), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1419]), .Q(data_mem_out_wire[1419]) );
  DFF \memory_reg[44][10]  ( .D(n6332), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1418]), .Q(data_mem_out_wire[1418]) );
  DFF \memory_reg[44][9]  ( .D(n6331), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1417]), .Q(data_mem_out_wire[1417]) );
  DFF \memory_reg[44][8]  ( .D(n6330), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1416]), .Q(data_mem_out_wire[1416]) );
  DFF \memory_reg[44][7]  ( .D(n6329), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1415]), .Q(data_mem_out_wire[1415]) );
  DFF \memory_reg[44][6]  ( .D(n6328), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1414]), .Q(data_mem_out_wire[1414]) );
  DFF \memory_reg[44][5]  ( .D(n6327), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1413]), .Q(data_mem_out_wire[1413]) );
  DFF \memory_reg[44][4]  ( .D(n6326), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1412]), .Q(data_mem_out_wire[1412]) );
  DFF \memory_reg[44][3]  ( .D(n6325), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1411]), .Q(data_mem_out_wire[1411]) );
  DFF \memory_reg[44][2]  ( .D(n6324), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1410]), .Q(data_mem_out_wire[1410]) );
  DFF \memory_reg[44][1]  ( .D(n6323), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1409]), .Q(data_mem_out_wire[1409]) );
  DFF \memory_reg[44][0]  ( .D(n6322), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1408]), .Q(data_mem_out_wire[1408]) );
  DFF \memory_reg[45][31]  ( .D(n6321), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1471]), .Q(data_mem_out_wire[1471]) );
  DFF \memory_reg[45][30]  ( .D(n6320), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1470]), .Q(data_mem_out_wire[1470]) );
  DFF \memory_reg[45][29]  ( .D(n6319), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1469]), .Q(data_mem_out_wire[1469]) );
  DFF \memory_reg[45][28]  ( .D(n6318), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1468]), .Q(data_mem_out_wire[1468]) );
  DFF \memory_reg[45][27]  ( .D(n6317), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1467]), .Q(data_mem_out_wire[1467]) );
  DFF \memory_reg[45][26]  ( .D(n6316), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1466]), .Q(data_mem_out_wire[1466]) );
  DFF \memory_reg[45][25]  ( .D(n6315), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1465]), .Q(data_mem_out_wire[1465]) );
  DFF \memory_reg[45][24]  ( .D(n6314), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1464]), .Q(data_mem_out_wire[1464]) );
  DFF \memory_reg[45][23]  ( .D(n6313), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1463]), .Q(data_mem_out_wire[1463]) );
  DFF \memory_reg[45][22]  ( .D(n6312), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1462]), .Q(data_mem_out_wire[1462]) );
  DFF \memory_reg[45][21]  ( .D(n6311), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1461]), .Q(data_mem_out_wire[1461]) );
  DFF \memory_reg[45][20]  ( .D(n6310), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1460]), .Q(data_mem_out_wire[1460]) );
  DFF \memory_reg[45][19]  ( .D(n6309), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1459]), .Q(data_mem_out_wire[1459]) );
  DFF \memory_reg[45][18]  ( .D(n6308), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1458]), .Q(data_mem_out_wire[1458]) );
  DFF \memory_reg[45][17]  ( .D(n6307), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1457]), .Q(data_mem_out_wire[1457]) );
  DFF \memory_reg[45][16]  ( .D(n6306), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1456]), .Q(data_mem_out_wire[1456]) );
  DFF \memory_reg[45][15]  ( .D(n6305), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1455]), .Q(data_mem_out_wire[1455]) );
  DFF \memory_reg[45][14]  ( .D(n6304), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1454]), .Q(data_mem_out_wire[1454]) );
  DFF \memory_reg[45][13]  ( .D(n6303), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1453]), .Q(data_mem_out_wire[1453]) );
  DFF \memory_reg[45][12]  ( .D(n6302), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1452]), .Q(data_mem_out_wire[1452]) );
  DFF \memory_reg[45][11]  ( .D(n6301), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1451]), .Q(data_mem_out_wire[1451]) );
  DFF \memory_reg[45][10]  ( .D(n6300), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1450]), .Q(data_mem_out_wire[1450]) );
  DFF \memory_reg[45][9]  ( .D(n6299), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1449]), .Q(data_mem_out_wire[1449]) );
  DFF \memory_reg[45][8]  ( .D(n6298), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1448]), .Q(data_mem_out_wire[1448]) );
  DFF \memory_reg[45][7]  ( .D(n6297), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1447]), .Q(data_mem_out_wire[1447]) );
  DFF \memory_reg[45][6]  ( .D(n6296), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1446]), .Q(data_mem_out_wire[1446]) );
  DFF \memory_reg[45][5]  ( .D(n6295), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1445]), .Q(data_mem_out_wire[1445]) );
  DFF \memory_reg[45][4]  ( .D(n6294), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1444]), .Q(data_mem_out_wire[1444]) );
  DFF \memory_reg[45][3]  ( .D(n6293), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1443]), .Q(data_mem_out_wire[1443]) );
  DFF \memory_reg[45][2]  ( .D(n6292), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1442]), .Q(data_mem_out_wire[1442]) );
  DFF \memory_reg[45][1]  ( .D(n6291), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1441]), .Q(data_mem_out_wire[1441]) );
  DFF \memory_reg[45][0]  ( .D(n6290), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1440]), .Q(data_mem_out_wire[1440]) );
  DFF \memory_reg[46][31]  ( .D(n6289), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1503]), .Q(data_mem_out_wire[1503]) );
  DFF \memory_reg[46][30]  ( .D(n6288), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1502]), .Q(data_mem_out_wire[1502]) );
  DFF \memory_reg[46][29]  ( .D(n6287), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1501]), .Q(data_mem_out_wire[1501]) );
  DFF \memory_reg[46][28]  ( .D(n6286), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1500]), .Q(data_mem_out_wire[1500]) );
  DFF \memory_reg[46][27]  ( .D(n6285), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1499]), .Q(data_mem_out_wire[1499]) );
  DFF \memory_reg[46][26]  ( .D(n6284), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1498]), .Q(data_mem_out_wire[1498]) );
  DFF \memory_reg[46][25]  ( .D(n6283), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1497]), .Q(data_mem_out_wire[1497]) );
  DFF \memory_reg[46][24]  ( .D(n6282), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1496]), .Q(data_mem_out_wire[1496]) );
  DFF \memory_reg[46][23]  ( .D(n6281), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1495]), .Q(data_mem_out_wire[1495]) );
  DFF \memory_reg[46][22]  ( .D(n6280), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1494]), .Q(data_mem_out_wire[1494]) );
  DFF \memory_reg[46][21]  ( .D(n6279), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1493]), .Q(data_mem_out_wire[1493]) );
  DFF \memory_reg[46][20]  ( .D(n6278), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1492]), .Q(data_mem_out_wire[1492]) );
  DFF \memory_reg[46][19]  ( .D(n6277), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1491]), .Q(data_mem_out_wire[1491]) );
  DFF \memory_reg[46][18]  ( .D(n6276), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1490]), .Q(data_mem_out_wire[1490]) );
  DFF \memory_reg[46][17]  ( .D(n6275), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1489]), .Q(data_mem_out_wire[1489]) );
  DFF \memory_reg[46][16]  ( .D(n6274), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1488]), .Q(data_mem_out_wire[1488]) );
  DFF \memory_reg[46][15]  ( .D(n6273), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1487]), .Q(data_mem_out_wire[1487]) );
  DFF \memory_reg[46][14]  ( .D(n6272), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1486]), .Q(data_mem_out_wire[1486]) );
  DFF \memory_reg[46][13]  ( .D(n6271), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1485]), .Q(data_mem_out_wire[1485]) );
  DFF \memory_reg[46][12]  ( .D(n6270), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1484]), .Q(data_mem_out_wire[1484]) );
  DFF \memory_reg[46][11]  ( .D(n6269), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1483]), .Q(data_mem_out_wire[1483]) );
  DFF \memory_reg[46][10]  ( .D(n6268), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1482]), .Q(data_mem_out_wire[1482]) );
  DFF \memory_reg[46][9]  ( .D(n6267), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1481]), .Q(data_mem_out_wire[1481]) );
  DFF \memory_reg[46][8]  ( .D(n6266), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1480]), .Q(data_mem_out_wire[1480]) );
  DFF \memory_reg[46][7]  ( .D(n6265), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1479]), .Q(data_mem_out_wire[1479]) );
  DFF \memory_reg[46][6]  ( .D(n6264), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1478]), .Q(data_mem_out_wire[1478]) );
  DFF \memory_reg[46][5]  ( .D(n6263), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1477]), .Q(data_mem_out_wire[1477]) );
  DFF \memory_reg[46][4]  ( .D(n6262), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1476]), .Q(data_mem_out_wire[1476]) );
  DFF \memory_reg[46][3]  ( .D(n6261), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1475]), .Q(data_mem_out_wire[1475]) );
  DFF \memory_reg[46][2]  ( .D(n6260), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1474]), .Q(data_mem_out_wire[1474]) );
  DFF \memory_reg[46][1]  ( .D(n6259), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1473]), .Q(data_mem_out_wire[1473]) );
  DFF \memory_reg[46][0]  ( .D(n6258), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1472]), .Q(data_mem_out_wire[1472]) );
  DFF \memory_reg[47][31]  ( .D(n6257), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1535]), .Q(data_mem_out_wire[1535]) );
  DFF \memory_reg[47][30]  ( .D(n6256), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1534]), .Q(data_mem_out_wire[1534]) );
  DFF \memory_reg[47][29]  ( .D(n6255), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1533]), .Q(data_mem_out_wire[1533]) );
  DFF \memory_reg[47][28]  ( .D(n6254), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1532]), .Q(data_mem_out_wire[1532]) );
  DFF \memory_reg[47][27]  ( .D(n6253), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1531]), .Q(data_mem_out_wire[1531]) );
  DFF \memory_reg[47][26]  ( .D(n6252), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1530]), .Q(data_mem_out_wire[1530]) );
  DFF \memory_reg[47][25]  ( .D(n6251), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1529]), .Q(data_mem_out_wire[1529]) );
  DFF \memory_reg[47][24]  ( .D(n6250), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1528]), .Q(data_mem_out_wire[1528]) );
  DFF \memory_reg[47][23]  ( .D(n6249), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1527]), .Q(data_mem_out_wire[1527]) );
  DFF \memory_reg[47][22]  ( .D(n6248), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1526]), .Q(data_mem_out_wire[1526]) );
  DFF \memory_reg[47][21]  ( .D(n6247), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1525]), .Q(data_mem_out_wire[1525]) );
  DFF \memory_reg[47][20]  ( .D(n6246), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1524]), .Q(data_mem_out_wire[1524]) );
  DFF \memory_reg[47][19]  ( .D(n6245), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1523]), .Q(data_mem_out_wire[1523]) );
  DFF \memory_reg[47][18]  ( .D(n6244), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1522]), .Q(data_mem_out_wire[1522]) );
  DFF \memory_reg[47][17]  ( .D(n6243), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1521]), .Q(data_mem_out_wire[1521]) );
  DFF \memory_reg[47][16]  ( .D(n6242), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1520]), .Q(data_mem_out_wire[1520]) );
  DFF \memory_reg[47][15]  ( .D(n6241), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1519]), .Q(data_mem_out_wire[1519]) );
  DFF \memory_reg[47][14]  ( .D(n6240), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1518]), .Q(data_mem_out_wire[1518]) );
  DFF \memory_reg[47][13]  ( .D(n6239), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1517]), .Q(data_mem_out_wire[1517]) );
  DFF \memory_reg[47][12]  ( .D(n6238), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1516]), .Q(data_mem_out_wire[1516]) );
  DFF \memory_reg[47][11]  ( .D(n6237), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1515]), .Q(data_mem_out_wire[1515]) );
  DFF \memory_reg[47][10]  ( .D(n6236), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1514]), .Q(data_mem_out_wire[1514]) );
  DFF \memory_reg[47][9]  ( .D(n6235), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1513]), .Q(data_mem_out_wire[1513]) );
  DFF \memory_reg[47][8]  ( .D(n6234), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1512]), .Q(data_mem_out_wire[1512]) );
  DFF \memory_reg[47][7]  ( .D(n6233), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1511]), .Q(data_mem_out_wire[1511]) );
  DFF \memory_reg[47][6]  ( .D(n6232), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1510]), .Q(data_mem_out_wire[1510]) );
  DFF \memory_reg[47][5]  ( .D(n6231), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1509]), .Q(data_mem_out_wire[1509]) );
  DFF \memory_reg[47][4]  ( .D(n6230), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1508]), .Q(data_mem_out_wire[1508]) );
  DFF \memory_reg[47][3]  ( .D(n6229), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1507]), .Q(data_mem_out_wire[1507]) );
  DFF \memory_reg[47][2]  ( .D(n6228), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1506]), .Q(data_mem_out_wire[1506]) );
  DFF \memory_reg[47][1]  ( .D(n6227), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1505]), .Q(data_mem_out_wire[1505]) );
  DFF \memory_reg[47][0]  ( .D(n6226), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1504]), .Q(data_mem_out_wire[1504]) );
  DFF \memory_reg[48][31]  ( .D(n6225), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1567]), .Q(data_mem_out_wire[1567]) );
  DFF \memory_reg[48][30]  ( .D(n6224), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1566]), .Q(data_mem_out_wire[1566]) );
  DFF \memory_reg[48][29]  ( .D(n6223), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1565]), .Q(data_mem_out_wire[1565]) );
  DFF \memory_reg[48][28]  ( .D(n6222), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1564]), .Q(data_mem_out_wire[1564]) );
  DFF \memory_reg[48][27]  ( .D(n6221), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1563]), .Q(data_mem_out_wire[1563]) );
  DFF \memory_reg[48][26]  ( .D(n6220), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1562]), .Q(data_mem_out_wire[1562]) );
  DFF \memory_reg[48][25]  ( .D(n6219), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1561]), .Q(data_mem_out_wire[1561]) );
  DFF \memory_reg[48][24]  ( .D(n6218), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1560]), .Q(data_mem_out_wire[1560]) );
  DFF \memory_reg[48][23]  ( .D(n6217), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1559]), .Q(data_mem_out_wire[1559]) );
  DFF \memory_reg[48][22]  ( .D(n6216), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1558]), .Q(data_mem_out_wire[1558]) );
  DFF \memory_reg[48][21]  ( .D(n6215), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1557]), .Q(data_mem_out_wire[1557]) );
  DFF \memory_reg[48][20]  ( .D(n6214), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1556]), .Q(data_mem_out_wire[1556]) );
  DFF \memory_reg[48][19]  ( .D(n6213), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1555]), .Q(data_mem_out_wire[1555]) );
  DFF \memory_reg[48][18]  ( .D(n6212), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1554]), .Q(data_mem_out_wire[1554]) );
  DFF \memory_reg[48][17]  ( .D(n6211), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1553]), .Q(data_mem_out_wire[1553]) );
  DFF \memory_reg[48][16]  ( .D(n6210), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1552]), .Q(data_mem_out_wire[1552]) );
  DFF \memory_reg[48][15]  ( .D(n6209), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1551]), .Q(data_mem_out_wire[1551]) );
  DFF \memory_reg[48][14]  ( .D(n6208), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1550]), .Q(data_mem_out_wire[1550]) );
  DFF \memory_reg[48][13]  ( .D(n6207), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1549]), .Q(data_mem_out_wire[1549]) );
  DFF \memory_reg[48][12]  ( .D(n6206), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1548]), .Q(data_mem_out_wire[1548]) );
  DFF \memory_reg[48][11]  ( .D(n6205), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1547]), .Q(data_mem_out_wire[1547]) );
  DFF \memory_reg[48][10]  ( .D(n6204), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1546]), .Q(data_mem_out_wire[1546]) );
  DFF \memory_reg[48][9]  ( .D(n6203), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1545]), .Q(data_mem_out_wire[1545]) );
  DFF \memory_reg[48][8]  ( .D(n6202), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1544]), .Q(data_mem_out_wire[1544]) );
  DFF \memory_reg[48][7]  ( .D(n6201), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1543]), .Q(data_mem_out_wire[1543]) );
  DFF \memory_reg[48][6]  ( .D(n6200), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1542]), .Q(data_mem_out_wire[1542]) );
  DFF \memory_reg[48][5]  ( .D(n6199), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1541]), .Q(data_mem_out_wire[1541]) );
  DFF \memory_reg[48][4]  ( .D(n6198), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1540]), .Q(data_mem_out_wire[1540]) );
  DFF \memory_reg[48][3]  ( .D(n6197), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1539]), .Q(data_mem_out_wire[1539]) );
  DFF \memory_reg[48][2]  ( .D(n6196), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1538]), .Q(data_mem_out_wire[1538]) );
  DFF \memory_reg[48][1]  ( .D(n6195), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1537]), .Q(data_mem_out_wire[1537]) );
  DFF \memory_reg[48][0]  ( .D(n6194), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1536]), .Q(data_mem_out_wire[1536]) );
  DFF \memory_reg[49][31]  ( .D(n6193), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1599]), .Q(data_mem_out_wire[1599]) );
  DFF \memory_reg[49][30]  ( .D(n6192), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1598]), .Q(data_mem_out_wire[1598]) );
  DFF \memory_reg[49][29]  ( .D(n6191), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1597]), .Q(data_mem_out_wire[1597]) );
  DFF \memory_reg[49][28]  ( .D(n6190), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1596]), .Q(data_mem_out_wire[1596]) );
  DFF \memory_reg[49][27]  ( .D(n6189), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1595]), .Q(data_mem_out_wire[1595]) );
  DFF \memory_reg[49][26]  ( .D(n6188), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1594]), .Q(data_mem_out_wire[1594]) );
  DFF \memory_reg[49][25]  ( .D(n6187), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1593]), .Q(data_mem_out_wire[1593]) );
  DFF \memory_reg[49][24]  ( .D(n6186), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1592]), .Q(data_mem_out_wire[1592]) );
  DFF \memory_reg[49][23]  ( .D(n6185), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1591]), .Q(data_mem_out_wire[1591]) );
  DFF \memory_reg[49][22]  ( .D(n6184), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1590]), .Q(data_mem_out_wire[1590]) );
  DFF \memory_reg[49][21]  ( .D(n6183), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1589]), .Q(data_mem_out_wire[1589]) );
  DFF \memory_reg[49][20]  ( .D(n6182), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1588]), .Q(data_mem_out_wire[1588]) );
  DFF \memory_reg[49][19]  ( .D(n6181), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1587]), .Q(data_mem_out_wire[1587]) );
  DFF \memory_reg[49][18]  ( .D(n6180), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1586]), .Q(data_mem_out_wire[1586]) );
  DFF \memory_reg[49][17]  ( .D(n6179), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1585]), .Q(data_mem_out_wire[1585]) );
  DFF \memory_reg[49][16]  ( .D(n6178), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1584]), .Q(data_mem_out_wire[1584]) );
  DFF \memory_reg[49][15]  ( .D(n6177), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1583]), .Q(data_mem_out_wire[1583]) );
  DFF \memory_reg[49][14]  ( .D(n6176), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1582]), .Q(data_mem_out_wire[1582]) );
  DFF \memory_reg[49][13]  ( .D(n6175), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1581]), .Q(data_mem_out_wire[1581]) );
  DFF \memory_reg[49][12]  ( .D(n6174), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1580]), .Q(data_mem_out_wire[1580]) );
  DFF \memory_reg[49][11]  ( .D(n6173), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1579]), .Q(data_mem_out_wire[1579]) );
  DFF \memory_reg[49][10]  ( .D(n6172), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1578]), .Q(data_mem_out_wire[1578]) );
  DFF \memory_reg[49][9]  ( .D(n6171), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1577]), .Q(data_mem_out_wire[1577]) );
  DFF \memory_reg[49][8]  ( .D(n6170), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1576]), .Q(data_mem_out_wire[1576]) );
  DFF \memory_reg[49][7]  ( .D(n6169), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1575]), .Q(data_mem_out_wire[1575]) );
  DFF \memory_reg[49][6]  ( .D(n6168), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1574]), .Q(data_mem_out_wire[1574]) );
  DFF \memory_reg[49][5]  ( .D(n6167), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1573]), .Q(data_mem_out_wire[1573]) );
  DFF \memory_reg[49][4]  ( .D(n6166), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1572]), .Q(data_mem_out_wire[1572]) );
  DFF \memory_reg[49][3]  ( .D(n6165), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1571]), .Q(data_mem_out_wire[1571]) );
  DFF \memory_reg[49][2]  ( .D(n6164), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1570]), .Q(data_mem_out_wire[1570]) );
  DFF \memory_reg[49][1]  ( .D(n6163), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1569]), .Q(data_mem_out_wire[1569]) );
  DFF \memory_reg[49][0]  ( .D(n6162), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1568]), .Q(data_mem_out_wire[1568]) );
  DFF \memory_reg[50][31]  ( .D(n6161), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1631]), .Q(data_mem_out_wire[1631]) );
  DFF \memory_reg[50][30]  ( .D(n6160), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1630]), .Q(data_mem_out_wire[1630]) );
  DFF \memory_reg[50][29]  ( .D(n6159), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1629]), .Q(data_mem_out_wire[1629]) );
  DFF \memory_reg[50][28]  ( .D(n6158), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1628]), .Q(data_mem_out_wire[1628]) );
  DFF \memory_reg[50][27]  ( .D(n6157), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1627]), .Q(data_mem_out_wire[1627]) );
  DFF \memory_reg[50][26]  ( .D(n6156), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1626]), .Q(data_mem_out_wire[1626]) );
  DFF \memory_reg[50][25]  ( .D(n6155), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1625]), .Q(data_mem_out_wire[1625]) );
  DFF \memory_reg[50][24]  ( .D(n6154), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1624]), .Q(data_mem_out_wire[1624]) );
  DFF \memory_reg[50][23]  ( .D(n6153), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1623]), .Q(data_mem_out_wire[1623]) );
  DFF \memory_reg[50][22]  ( .D(n6152), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1622]), .Q(data_mem_out_wire[1622]) );
  DFF \memory_reg[50][21]  ( .D(n6151), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1621]), .Q(data_mem_out_wire[1621]) );
  DFF \memory_reg[50][20]  ( .D(n6150), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1620]), .Q(data_mem_out_wire[1620]) );
  DFF \memory_reg[50][19]  ( .D(n6149), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1619]), .Q(data_mem_out_wire[1619]) );
  DFF \memory_reg[50][18]  ( .D(n6148), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1618]), .Q(data_mem_out_wire[1618]) );
  DFF \memory_reg[50][17]  ( .D(n6147), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1617]), .Q(data_mem_out_wire[1617]) );
  DFF \memory_reg[50][16]  ( .D(n6146), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1616]), .Q(data_mem_out_wire[1616]) );
  DFF \memory_reg[50][15]  ( .D(n6145), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1615]), .Q(data_mem_out_wire[1615]) );
  DFF \memory_reg[50][14]  ( .D(n6144), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1614]), .Q(data_mem_out_wire[1614]) );
  DFF \memory_reg[50][13]  ( .D(n6143), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1613]), .Q(data_mem_out_wire[1613]) );
  DFF \memory_reg[50][12]  ( .D(n6142), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1612]), .Q(data_mem_out_wire[1612]) );
  DFF \memory_reg[50][11]  ( .D(n6141), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1611]), .Q(data_mem_out_wire[1611]) );
  DFF \memory_reg[50][10]  ( .D(n6140), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1610]), .Q(data_mem_out_wire[1610]) );
  DFF \memory_reg[50][9]  ( .D(n6139), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1609]), .Q(data_mem_out_wire[1609]) );
  DFF \memory_reg[50][8]  ( .D(n6138), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1608]), .Q(data_mem_out_wire[1608]) );
  DFF \memory_reg[50][7]  ( .D(n6137), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1607]), .Q(data_mem_out_wire[1607]) );
  DFF \memory_reg[50][6]  ( .D(n6136), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1606]), .Q(data_mem_out_wire[1606]) );
  DFF \memory_reg[50][5]  ( .D(n6135), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1605]), .Q(data_mem_out_wire[1605]) );
  DFF \memory_reg[50][4]  ( .D(n6134), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1604]), .Q(data_mem_out_wire[1604]) );
  DFF \memory_reg[50][3]  ( .D(n6133), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1603]), .Q(data_mem_out_wire[1603]) );
  DFF \memory_reg[50][2]  ( .D(n6132), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1602]), .Q(data_mem_out_wire[1602]) );
  DFF \memory_reg[50][1]  ( .D(n6131), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1601]), .Q(data_mem_out_wire[1601]) );
  DFF \memory_reg[50][0]  ( .D(n6130), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1600]), .Q(data_mem_out_wire[1600]) );
  DFF \memory_reg[51][31]  ( .D(n6129), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1663]), .Q(data_mem_out_wire[1663]) );
  DFF \memory_reg[51][30]  ( .D(n6128), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1662]), .Q(data_mem_out_wire[1662]) );
  DFF \memory_reg[51][29]  ( .D(n6127), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1661]), .Q(data_mem_out_wire[1661]) );
  DFF \memory_reg[51][28]  ( .D(n6126), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1660]), .Q(data_mem_out_wire[1660]) );
  DFF \memory_reg[51][27]  ( .D(n6125), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1659]), .Q(data_mem_out_wire[1659]) );
  DFF \memory_reg[51][26]  ( .D(n6124), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1658]), .Q(data_mem_out_wire[1658]) );
  DFF \memory_reg[51][25]  ( .D(n6123), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1657]), .Q(data_mem_out_wire[1657]) );
  DFF \memory_reg[51][24]  ( .D(n6122), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1656]), .Q(data_mem_out_wire[1656]) );
  DFF \memory_reg[51][23]  ( .D(n6121), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1655]), .Q(data_mem_out_wire[1655]) );
  DFF \memory_reg[51][22]  ( .D(n6120), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1654]), .Q(data_mem_out_wire[1654]) );
  DFF \memory_reg[51][21]  ( .D(n6119), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1653]), .Q(data_mem_out_wire[1653]) );
  DFF \memory_reg[51][20]  ( .D(n6118), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1652]), .Q(data_mem_out_wire[1652]) );
  DFF \memory_reg[51][19]  ( .D(n6117), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1651]), .Q(data_mem_out_wire[1651]) );
  DFF \memory_reg[51][18]  ( .D(n6116), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1650]), .Q(data_mem_out_wire[1650]) );
  DFF \memory_reg[51][17]  ( .D(n6115), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1649]), .Q(data_mem_out_wire[1649]) );
  DFF \memory_reg[51][16]  ( .D(n6114), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1648]), .Q(data_mem_out_wire[1648]) );
  DFF \memory_reg[51][15]  ( .D(n6113), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1647]), .Q(data_mem_out_wire[1647]) );
  DFF \memory_reg[51][14]  ( .D(n6112), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1646]), .Q(data_mem_out_wire[1646]) );
  DFF \memory_reg[51][13]  ( .D(n6111), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1645]), .Q(data_mem_out_wire[1645]) );
  DFF \memory_reg[51][12]  ( .D(n6110), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1644]), .Q(data_mem_out_wire[1644]) );
  DFF \memory_reg[51][11]  ( .D(n6109), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1643]), .Q(data_mem_out_wire[1643]) );
  DFF \memory_reg[51][10]  ( .D(n6108), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1642]), .Q(data_mem_out_wire[1642]) );
  DFF \memory_reg[51][9]  ( .D(n6107), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1641]), .Q(data_mem_out_wire[1641]) );
  DFF \memory_reg[51][8]  ( .D(n6106), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1640]), .Q(data_mem_out_wire[1640]) );
  DFF \memory_reg[51][7]  ( .D(n6105), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1639]), .Q(data_mem_out_wire[1639]) );
  DFF \memory_reg[51][6]  ( .D(n6104), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1638]), .Q(data_mem_out_wire[1638]) );
  DFF \memory_reg[51][5]  ( .D(n6103), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1637]), .Q(data_mem_out_wire[1637]) );
  DFF \memory_reg[51][4]  ( .D(n6102), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1636]), .Q(data_mem_out_wire[1636]) );
  DFF \memory_reg[51][3]  ( .D(n6101), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1635]), .Q(data_mem_out_wire[1635]) );
  DFF \memory_reg[51][2]  ( .D(n6100), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1634]), .Q(data_mem_out_wire[1634]) );
  DFF \memory_reg[51][1]  ( .D(n6099), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1633]), .Q(data_mem_out_wire[1633]) );
  DFF \memory_reg[51][0]  ( .D(n6098), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1632]), .Q(data_mem_out_wire[1632]) );
  DFF \memory_reg[52][31]  ( .D(n6097), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1695]), .Q(data_mem_out_wire[1695]) );
  DFF \memory_reg[52][30]  ( .D(n6096), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1694]), .Q(data_mem_out_wire[1694]) );
  DFF \memory_reg[52][29]  ( .D(n6095), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1693]), .Q(data_mem_out_wire[1693]) );
  DFF \memory_reg[52][28]  ( .D(n6094), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1692]), .Q(data_mem_out_wire[1692]) );
  DFF \memory_reg[52][27]  ( .D(n6093), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1691]), .Q(data_mem_out_wire[1691]) );
  DFF \memory_reg[52][26]  ( .D(n6092), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1690]), .Q(data_mem_out_wire[1690]) );
  DFF \memory_reg[52][25]  ( .D(n6091), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1689]), .Q(data_mem_out_wire[1689]) );
  DFF \memory_reg[52][24]  ( .D(n6090), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1688]), .Q(data_mem_out_wire[1688]) );
  DFF \memory_reg[52][23]  ( .D(n6089), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1687]), .Q(data_mem_out_wire[1687]) );
  DFF \memory_reg[52][22]  ( .D(n6088), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1686]), .Q(data_mem_out_wire[1686]) );
  DFF \memory_reg[52][21]  ( .D(n6087), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1685]), .Q(data_mem_out_wire[1685]) );
  DFF \memory_reg[52][20]  ( .D(n6086), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1684]), .Q(data_mem_out_wire[1684]) );
  DFF \memory_reg[52][19]  ( .D(n6085), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1683]), .Q(data_mem_out_wire[1683]) );
  DFF \memory_reg[52][18]  ( .D(n6084), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1682]), .Q(data_mem_out_wire[1682]) );
  DFF \memory_reg[52][17]  ( .D(n6083), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1681]), .Q(data_mem_out_wire[1681]) );
  DFF \memory_reg[52][16]  ( .D(n6082), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1680]), .Q(data_mem_out_wire[1680]) );
  DFF \memory_reg[52][15]  ( .D(n6081), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1679]), .Q(data_mem_out_wire[1679]) );
  DFF \memory_reg[52][14]  ( .D(n6080), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1678]), .Q(data_mem_out_wire[1678]) );
  DFF \memory_reg[52][13]  ( .D(n6079), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1677]), .Q(data_mem_out_wire[1677]) );
  DFF \memory_reg[52][12]  ( .D(n6078), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1676]), .Q(data_mem_out_wire[1676]) );
  DFF \memory_reg[52][11]  ( .D(n6077), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1675]), .Q(data_mem_out_wire[1675]) );
  DFF \memory_reg[52][10]  ( .D(n6076), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1674]), .Q(data_mem_out_wire[1674]) );
  DFF \memory_reg[52][9]  ( .D(n6075), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1673]), .Q(data_mem_out_wire[1673]) );
  DFF \memory_reg[52][8]  ( .D(n6074), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1672]), .Q(data_mem_out_wire[1672]) );
  DFF \memory_reg[52][7]  ( .D(n6073), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1671]), .Q(data_mem_out_wire[1671]) );
  DFF \memory_reg[52][6]  ( .D(n6072), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1670]), .Q(data_mem_out_wire[1670]) );
  DFF \memory_reg[52][5]  ( .D(n6071), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1669]), .Q(data_mem_out_wire[1669]) );
  DFF \memory_reg[52][4]  ( .D(n6070), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1668]), .Q(data_mem_out_wire[1668]) );
  DFF \memory_reg[52][3]  ( .D(n6069), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1667]), .Q(data_mem_out_wire[1667]) );
  DFF \memory_reg[52][2]  ( .D(n6068), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1666]), .Q(data_mem_out_wire[1666]) );
  DFF \memory_reg[52][1]  ( .D(n6067), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1665]), .Q(data_mem_out_wire[1665]) );
  DFF \memory_reg[52][0]  ( .D(n6066), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1664]), .Q(data_mem_out_wire[1664]) );
  DFF \memory_reg[53][31]  ( .D(n6065), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1727]), .Q(data_mem_out_wire[1727]) );
  DFF \memory_reg[53][30]  ( .D(n6064), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1726]), .Q(data_mem_out_wire[1726]) );
  DFF \memory_reg[53][29]  ( .D(n6063), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1725]), .Q(data_mem_out_wire[1725]) );
  DFF \memory_reg[53][28]  ( .D(n6062), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1724]), .Q(data_mem_out_wire[1724]) );
  DFF \memory_reg[53][27]  ( .D(n6061), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1723]), .Q(data_mem_out_wire[1723]) );
  DFF \memory_reg[53][26]  ( .D(n6060), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1722]), .Q(data_mem_out_wire[1722]) );
  DFF \memory_reg[53][25]  ( .D(n6059), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1721]), .Q(data_mem_out_wire[1721]) );
  DFF \memory_reg[53][24]  ( .D(n6058), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1720]), .Q(data_mem_out_wire[1720]) );
  DFF \memory_reg[53][23]  ( .D(n6057), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1719]), .Q(data_mem_out_wire[1719]) );
  DFF \memory_reg[53][22]  ( .D(n6056), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1718]), .Q(data_mem_out_wire[1718]) );
  DFF \memory_reg[53][21]  ( .D(n6055), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1717]), .Q(data_mem_out_wire[1717]) );
  DFF \memory_reg[53][20]  ( .D(n6054), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1716]), .Q(data_mem_out_wire[1716]) );
  DFF \memory_reg[53][19]  ( .D(n6053), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1715]), .Q(data_mem_out_wire[1715]) );
  DFF \memory_reg[53][18]  ( .D(n6052), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1714]), .Q(data_mem_out_wire[1714]) );
  DFF \memory_reg[53][17]  ( .D(n6051), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1713]), .Q(data_mem_out_wire[1713]) );
  DFF \memory_reg[53][16]  ( .D(n6050), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1712]), .Q(data_mem_out_wire[1712]) );
  DFF \memory_reg[53][15]  ( .D(n6049), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1711]), .Q(data_mem_out_wire[1711]) );
  DFF \memory_reg[53][14]  ( .D(n6048), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1710]), .Q(data_mem_out_wire[1710]) );
  DFF \memory_reg[53][13]  ( .D(n6047), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1709]), .Q(data_mem_out_wire[1709]) );
  DFF \memory_reg[53][12]  ( .D(n6046), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1708]), .Q(data_mem_out_wire[1708]) );
  DFF \memory_reg[53][11]  ( .D(n6045), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1707]), .Q(data_mem_out_wire[1707]) );
  DFF \memory_reg[53][10]  ( .D(n6044), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1706]), .Q(data_mem_out_wire[1706]) );
  DFF \memory_reg[53][9]  ( .D(n6043), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1705]), .Q(data_mem_out_wire[1705]) );
  DFF \memory_reg[53][8]  ( .D(n6042), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1704]), .Q(data_mem_out_wire[1704]) );
  DFF \memory_reg[53][7]  ( .D(n6041), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1703]), .Q(data_mem_out_wire[1703]) );
  DFF \memory_reg[53][6]  ( .D(n6040), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1702]), .Q(data_mem_out_wire[1702]) );
  DFF \memory_reg[53][5]  ( .D(n6039), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1701]), .Q(data_mem_out_wire[1701]) );
  DFF \memory_reg[53][4]  ( .D(n6038), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1700]), .Q(data_mem_out_wire[1700]) );
  DFF \memory_reg[53][3]  ( .D(n6037), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1699]), .Q(data_mem_out_wire[1699]) );
  DFF \memory_reg[53][2]  ( .D(n6036), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1698]), .Q(data_mem_out_wire[1698]) );
  DFF \memory_reg[53][1]  ( .D(n6035), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1697]), .Q(data_mem_out_wire[1697]) );
  DFF \memory_reg[53][0]  ( .D(n6034), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1696]), .Q(data_mem_out_wire[1696]) );
  DFF \memory_reg[54][31]  ( .D(n6033), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1759]), .Q(data_mem_out_wire[1759]) );
  DFF \memory_reg[54][30]  ( .D(n6032), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1758]), .Q(data_mem_out_wire[1758]) );
  DFF \memory_reg[54][29]  ( .D(n6031), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1757]), .Q(data_mem_out_wire[1757]) );
  DFF \memory_reg[54][28]  ( .D(n6030), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1756]), .Q(data_mem_out_wire[1756]) );
  DFF \memory_reg[54][27]  ( .D(n6029), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1755]), .Q(data_mem_out_wire[1755]) );
  DFF \memory_reg[54][26]  ( .D(n6028), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1754]), .Q(data_mem_out_wire[1754]) );
  DFF \memory_reg[54][25]  ( .D(n6027), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1753]), .Q(data_mem_out_wire[1753]) );
  DFF \memory_reg[54][24]  ( .D(n6026), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1752]), .Q(data_mem_out_wire[1752]) );
  DFF \memory_reg[54][23]  ( .D(n6025), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1751]), .Q(data_mem_out_wire[1751]) );
  DFF \memory_reg[54][22]  ( .D(n6024), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1750]), .Q(data_mem_out_wire[1750]) );
  DFF \memory_reg[54][21]  ( .D(n6023), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1749]), .Q(data_mem_out_wire[1749]) );
  DFF \memory_reg[54][20]  ( .D(n6022), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1748]), .Q(data_mem_out_wire[1748]) );
  DFF \memory_reg[54][19]  ( .D(n6021), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1747]), .Q(data_mem_out_wire[1747]) );
  DFF \memory_reg[54][18]  ( .D(n6020), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1746]), .Q(data_mem_out_wire[1746]) );
  DFF \memory_reg[54][17]  ( .D(n6019), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1745]), .Q(data_mem_out_wire[1745]) );
  DFF \memory_reg[54][16]  ( .D(n6018), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1744]), .Q(data_mem_out_wire[1744]) );
  DFF \memory_reg[54][15]  ( .D(n6017), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1743]), .Q(data_mem_out_wire[1743]) );
  DFF \memory_reg[54][14]  ( .D(n6016), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1742]), .Q(data_mem_out_wire[1742]) );
  DFF \memory_reg[54][13]  ( .D(n6015), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1741]), .Q(data_mem_out_wire[1741]) );
  DFF \memory_reg[54][12]  ( .D(n6014), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1740]), .Q(data_mem_out_wire[1740]) );
  DFF \memory_reg[54][11]  ( .D(n6013), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1739]), .Q(data_mem_out_wire[1739]) );
  DFF \memory_reg[54][10]  ( .D(n6012), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1738]), .Q(data_mem_out_wire[1738]) );
  DFF \memory_reg[54][9]  ( .D(n6011), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1737]), .Q(data_mem_out_wire[1737]) );
  DFF \memory_reg[54][8]  ( .D(n6010), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1736]), .Q(data_mem_out_wire[1736]) );
  DFF \memory_reg[54][7]  ( .D(n6009), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1735]), .Q(data_mem_out_wire[1735]) );
  DFF \memory_reg[54][6]  ( .D(n6008), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1734]), .Q(data_mem_out_wire[1734]) );
  DFF \memory_reg[54][5]  ( .D(n6007), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1733]), .Q(data_mem_out_wire[1733]) );
  DFF \memory_reg[54][4]  ( .D(n6006), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1732]), .Q(data_mem_out_wire[1732]) );
  DFF \memory_reg[54][3]  ( .D(n6005), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1731]), .Q(data_mem_out_wire[1731]) );
  DFF \memory_reg[54][2]  ( .D(n6004), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1730]), .Q(data_mem_out_wire[1730]) );
  DFF \memory_reg[54][1]  ( .D(n6003), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1729]), .Q(data_mem_out_wire[1729]) );
  DFF \memory_reg[54][0]  ( .D(n6002), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1728]), .Q(data_mem_out_wire[1728]) );
  DFF \memory_reg[55][31]  ( .D(n6001), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1791]), .Q(data_mem_out_wire[1791]) );
  DFF \memory_reg[55][30]  ( .D(n6000), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1790]), .Q(data_mem_out_wire[1790]) );
  DFF \memory_reg[55][29]  ( .D(n5999), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1789]), .Q(data_mem_out_wire[1789]) );
  DFF \memory_reg[55][28]  ( .D(n5998), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1788]), .Q(data_mem_out_wire[1788]) );
  DFF \memory_reg[55][27]  ( .D(n5997), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1787]), .Q(data_mem_out_wire[1787]) );
  DFF \memory_reg[55][26]  ( .D(n5996), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1786]), .Q(data_mem_out_wire[1786]) );
  DFF \memory_reg[55][25]  ( .D(n5995), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1785]), .Q(data_mem_out_wire[1785]) );
  DFF \memory_reg[55][24]  ( .D(n5994), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1784]), .Q(data_mem_out_wire[1784]) );
  DFF \memory_reg[55][23]  ( .D(n5993), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1783]), .Q(data_mem_out_wire[1783]) );
  DFF \memory_reg[55][22]  ( .D(n5992), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1782]), .Q(data_mem_out_wire[1782]) );
  DFF \memory_reg[55][21]  ( .D(n5991), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1781]), .Q(data_mem_out_wire[1781]) );
  DFF \memory_reg[55][20]  ( .D(n5990), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1780]), .Q(data_mem_out_wire[1780]) );
  DFF \memory_reg[55][19]  ( .D(n5989), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1779]), .Q(data_mem_out_wire[1779]) );
  DFF \memory_reg[55][18]  ( .D(n5988), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1778]), .Q(data_mem_out_wire[1778]) );
  DFF \memory_reg[55][17]  ( .D(n5987), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1777]), .Q(data_mem_out_wire[1777]) );
  DFF \memory_reg[55][16]  ( .D(n5986), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1776]), .Q(data_mem_out_wire[1776]) );
  DFF \memory_reg[55][15]  ( .D(n5985), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1775]), .Q(data_mem_out_wire[1775]) );
  DFF \memory_reg[55][14]  ( .D(n5984), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1774]), .Q(data_mem_out_wire[1774]) );
  DFF \memory_reg[55][13]  ( .D(n5983), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1773]), .Q(data_mem_out_wire[1773]) );
  DFF \memory_reg[55][12]  ( .D(n5982), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1772]), .Q(data_mem_out_wire[1772]) );
  DFF \memory_reg[55][11]  ( .D(n5981), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1771]), .Q(data_mem_out_wire[1771]) );
  DFF \memory_reg[55][10]  ( .D(n5980), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1770]), .Q(data_mem_out_wire[1770]) );
  DFF \memory_reg[55][9]  ( .D(n5979), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1769]), .Q(data_mem_out_wire[1769]) );
  DFF \memory_reg[55][8]  ( .D(n5978), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1768]), .Q(data_mem_out_wire[1768]) );
  DFF \memory_reg[55][7]  ( .D(n5977), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1767]), .Q(data_mem_out_wire[1767]) );
  DFF \memory_reg[55][6]  ( .D(n5976), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1766]), .Q(data_mem_out_wire[1766]) );
  DFF \memory_reg[55][5]  ( .D(n5975), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1765]), .Q(data_mem_out_wire[1765]) );
  DFF \memory_reg[55][4]  ( .D(n5974), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1764]), .Q(data_mem_out_wire[1764]) );
  DFF \memory_reg[55][3]  ( .D(n5973), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1763]), .Q(data_mem_out_wire[1763]) );
  DFF \memory_reg[55][2]  ( .D(n5972), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1762]), .Q(data_mem_out_wire[1762]) );
  DFF \memory_reg[55][1]  ( .D(n5971), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1761]), .Q(data_mem_out_wire[1761]) );
  DFF \memory_reg[55][0]  ( .D(n5970), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1760]), .Q(data_mem_out_wire[1760]) );
  DFF \memory_reg[56][31]  ( .D(n5969), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1823]), .Q(data_mem_out_wire[1823]) );
  DFF \memory_reg[56][30]  ( .D(n5968), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1822]), .Q(data_mem_out_wire[1822]) );
  DFF \memory_reg[56][29]  ( .D(n5967), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1821]), .Q(data_mem_out_wire[1821]) );
  DFF \memory_reg[56][28]  ( .D(n5966), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1820]), .Q(data_mem_out_wire[1820]) );
  DFF \memory_reg[56][27]  ( .D(n5965), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1819]), .Q(data_mem_out_wire[1819]) );
  DFF \memory_reg[56][26]  ( .D(n5964), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1818]), .Q(data_mem_out_wire[1818]) );
  DFF \memory_reg[56][25]  ( .D(n5963), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1817]), .Q(data_mem_out_wire[1817]) );
  DFF \memory_reg[56][24]  ( .D(n5962), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1816]), .Q(data_mem_out_wire[1816]) );
  DFF \memory_reg[56][23]  ( .D(n5961), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1815]), .Q(data_mem_out_wire[1815]) );
  DFF \memory_reg[56][22]  ( .D(n5960), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1814]), .Q(data_mem_out_wire[1814]) );
  DFF \memory_reg[56][21]  ( .D(n5959), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1813]), .Q(data_mem_out_wire[1813]) );
  DFF \memory_reg[56][20]  ( .D(n5958), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1812]), .Q(data_mem_out_wire[1812]) );
  DFF \memory_reg[56][19]  ( .D(n5957), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1811]), .Q(data_mem_out_wire[1811]) );
  DFF \memory_reg[56][18]  ( .D(n5956), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1810]), .Q(data_mem_out_wire[1810]) );
  DFF \memory_reg[56][17]  ( .D(n5955), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1809]), .Q(data_mem_out_wire[1809]) );
  DFF \memory_reg[56][16]  ( .D(n5954), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1808]), .Q(data_mem_out_wire[1808]) );
  DFF \memory_reg[56][15]  ( .D(n5953), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1807]), .Q(data_mem_out_wire[1807]) );
  DFF \memory_reg[56][14]  ( .D(n5952), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1806]), .Q(data_mem_out_wire[1806]) );
  DFF \memory_reg[56][13]  ( .D(n5951), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1805]), .Q(data_mem_out_wire[1805]) );
  DFF \memory_reg[56][12]  ( .D(n5950), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1804]), .Q(data_mem_out_wire[1804]) );
  DFF \memory_reg[56][11]  ( .D(n5949), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1803]), .Q(data_mem_out_wire[1803]) );
  DFF \memory_reg[56][10]  ( .D(n5948), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1802]), .Q(data_mem_out_wire[1802]) );
  DFF \memory_reg[56][9]  ( .D(n5947), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1801]), .Q(data_mem_out_wire[1801]) );
  DFF \memory_reg[56][8]  ( .D(n5946), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1800]), .Q(data_mem_out_wire[1800]) );
  DFF \memory_reg[56][7]  ( .D(n5945), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1799]), .Q(data_mem_out_wire[1799]) );
  DFF \memory_reg[56][6]  ( .D(n5944), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1798]), .Q(data_mem_out_wire[1798]) );
  DFF \memory_reg[56][5]  ( .D(n5943), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1797]), .Q(data_mem_out_wire[1797]) );
  DFF \memory_reg[56][4]  ( .D(n5942), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1796]), .Q(data_mem_out_wire[1796]) );
  DFF \memory_reg[56][3]  ( .D(n5941), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1795]), .Q(data_mem_out_wire[1795]) );
  DFF \memory_reg[56][2]  ( .D(n5940), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1794]), .Q(data_mem_out_wire[1794]) );
  DFF \memory_reg[56][1]  ( .D(n5939), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1793]), .Q(data_mem_out_wire[1793]) );
  DFF \memory_reg[56][0]  ( .D(n5938), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1792]), .Q(data_mem_out_wire[1792]) );
  DFF \memory_reg[57][31]  ( .D(n5937), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1855]), .Q(data_mem_out_wire[1855]) );
  DFF \memory_reg[57][30]  ( .D(n5936), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1854]), .Q(data_mem_out_wire[1854]) );
  DFF \memory_reg[57][29]  ( .D(n5935), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1853]), .Q(data_mem_out_wire[1853]) );
  DFF \memory_reg[57][28]  ( .D(n5934), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1852]), .Q(data_mem_out_wire[1852]) );
  DFF \memory_reg[57][27]  ( .D(n5933), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1851]), .Q(data_mem_out_wire[1851]) );
  DFF \memory_reg[57][26]  ( .D(n5932), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1850]), .Q(data_mem_out_wire[1850]) );
  DFF \memory_reg[57][25]  ( .D(n5931), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1849]), .Q(data_mem_out_wire[1849]) );
  DFF \memory_reg[57][24]  ( .D(n5930), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1848]), .Q(data_mem_out_wire[1848]) );
  DFF \memory_reg[57][23]  ( .D(n5929), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1847]), .Q(data_mem_out_wire[1847]) );
  DFF \memory_reg[57][22]  ( .D(n5928), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1846]), .Q(data_mem_out_wire[1846]) );
  DFF \memory_reg[57][21]  ( .D(n5927), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1845]), .Q(data_mem_out_wire[1845]) );
  DFF \memory_reg[57][20]  ( .D(n5926), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1844]), .Q(data_mem_out_wire[1844]) );
  DFF \memory_reg[57][19]  ( .D(n5925), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1843]), .Q(data_mem_out_wire[1843]) );
  DFF \memory_reg[57][18]  ( .D(n5924), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1842]), .Q(data_mem_out_wire[1842]) );
  DFF \memory_reg[57][17]  ( .D(n5923), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1841]), .Q(data_mem_out_wire[1841]) );
  DFF \memory_reg[57][16]  ( .D(n5922), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1840]), .Q(data_mem_out_wire[1840]) );
  DFF \memory_reg[57][15]  ( .D(n5921), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1839]), .Q(data_mem_out_wire[1839]) );
  DFF \memory_reg[57][14]  ( .D(n5920), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1838]), .Q(data_mem_out_wire[1838]) );
  DFF \memory_reg[57][13]  ( .D(n5919), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1837]), .Q(data_mem_out_wire[1837]) );
  DFF \memory_reg[57][12]  ( .D(n5918), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1836]), .Q(data_mem_out_wire[1836]) );
  DFF \memory_reg[57][11]  ( .D(n5917), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1835]), .Q(data_mem_out_wire[1835]) );
  DFF \memory_reg[57][10]  ( .D(n5916), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1834]), .Q(data_mem_out_wire[1834]) );
  DFF \memory_reg[57][9]  ( .D(n5915), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1833]), .Q(data_mem_out_wire[1833]) );
  DFF \memory_reg[57][8]  ( .D(n5914), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1832]), .Q(data_mem_out_wire[1832]) );
  DFF \memory_reg[57][7]  ( .D(n5913), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1831]), .Q(data_mem_out_wire[1831]) );
  DFF \memory_reg[57][6]  ( .D(n5912), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1830]), .Q(data_mem_out_wire[1830]) );
  DFF \memory_reg[57][5]  ( .D(n5911), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1829]), .Q(data_mem_out_wire[1829]) );
  DFF \memory_reg[57][4]  ( .D(n5910), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1828]), .Q(data_mem_out_wire[1828]) );
  DFF \memory_reg[57][3]  ( .D(n5909), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1827]), .Q(data_mem_out_wire[1827]) );
  DFF \memory_reg[57][2]  ( .D(n5908), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1826]), .Q(data_mem_out_wire[1826]) );
  DFF \memory_reg[57][1]  ( .D(n5907), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1825]), .Q(data_mem_out_wire[1825]) );
  DFF \memory_reg[57][0]  ( .D(n5906), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1824]), .Q(data_mem_out_wire[1824]) );
  DFF \memory_reg[58][31]  ( .D(n5905), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1887]), .Q(data_mem_out_wire[1887]) );
  DFF \memory_reg[58][30]  ( .D(n5904), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1886]), .Q(data_mem_out_wire[1886]) );
  DFF \memory_reg[58][29]  ( .D(n5903), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1885]), .Q(data_mem_out_wire[1885]) );
  DFF \memory_reg[58][28]  ( .D(n5902), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1884]), .Q(data_mem_out_wire[1884]) );
  DFF \memory_reg[58][27]  ( .D(n5901), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1883]), .Q(data_mem_out_wire[1883]) );
  DFF \memory_reg[58][26]  ( .D(n5900), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1882]), .Q(data_mem_out_wire[1882]) );
  DFF \memory_reg[58][25]  ( .D(n5899), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1881]), .Q(data_mem_out_wire[1881]) );
  DFF \memory_reg[58][24]  ( .D(n5898), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1880]), .Q(data_mem_out_wire[1880]) );
  DFF \memory_reg[58][23]  ( .D(n5897), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1879]), .Q(data_mem_out_wire[1879]) );
  DFF \memory_reg[58][22]  ( .D(n5896), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1878]), .Q(data_mem_out_wire[1878]) );
  DFF \memory_reg[58][21]  ( .D(n5895), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1877]), .Q(data_mem_out_wire[1877]) );
  DFF \memory_reg[58][20]  ( .D(n5894), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1876]), .Q(data_mem_out_wire[1876]) );
  DFF \memory_reg[58][19]  ( .D(n5893), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1875]), .Q(data_mem_out_wire[1875]) );
  DFF \memory_reg[58][18]  ( .D(n5892), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1874]), .Q(data_mem_out_wire[1874]) );
  DFF \memory_reg[58][17]  ( .D(n5891), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1873]), .Q(data_mem_out_wire[1873]) );
  DFF \memory_reg[58][16]  ( .D(n5890), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1872]), .Q(data_mem_out_wire[1872]) );
  DFF \memory_reg[58][15]  ( .D(n5889), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1871]), .Q(data_mem_out_wire[1871]) );
  DFF \memory_reg[58][14]  ( .D(n5888), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1870]), .Q(data_mem_out_wire[1870]) );
  DFF \memory_reg[58][13]  ( .D(n5887), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1869]), .Q(data_mem_out_wire[1869]) );
  DFF \memory_reg[58][12]  ( .D(n5886), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1868]), .Q(data_mem_out_wire[1868]) );
  DFF \memory_reg[58][11]  ( .D(n5885), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1867]), .Q(data_mem_out_wire[1867]) );
  DFF \memory_reg[58][10]  ( .D(n5884), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1866]), .Q(data_mem_out_wire[1866]) );
  DFF \memory_reg[58][9]  ( .D(n5883), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1865]), .Q(data_mem_out_wire[1865]) );
  DFF \memory_reg[58][8]  ( .D(n5882), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1864]), .Q(data_mem_out_wire[1864]) );
  DFF \memory_reg[58][7]  ( .D(n5881), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1863]), .Q(data_mem_out_wire[1863]) );
  DFF \memory_reg[58][6]  ( .D(n5880), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1862]), .Q(data_mem_out_wire[1862]) );
  DFF \memory_reg[58][5]  ( .D(n5879), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1861]), .Q(data_mem_out_wire[1861]) );
  DFF \memory_reg[58][4]  ( .D(n5878), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1860]), .Q(data_mem_out_wire[1860]) );
  DFF \memory_reg[58][3]  ( .D(n5877), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1859]), .Q(data_mem_out_wire[1859]) );
  DFF \memory_reg[58][2]  ( .D(n5876), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1858]), .Q(data_mem_out_wire[1858]) );
  DFF \memory_reg[58][1]  ( .D(n5875), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1857]), .Q(data_mem_out_wire[1857]) );
  DFF \memory_reg[58][0]  ( .D(n5874), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1856]), .Q(data_mem_out_wire[1856]) );
  DFF \memory_reg[59][31]  ( .D(n5873), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1919]), .Q(data_mem_out_wire[1919]) );
  DFF \memory_reg[59][30]  ( .D(n5872), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1918]), .Q(data_mem_out_wire[1918]) );
  DFF \memory_reg[59][29]  ( .D(n5871), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1917]), .Q(data_mem_out_wire[1917]) );
  DFF \memory_reg[59][28]  ( .D(n5870), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1916]), .Q(data_mem_out_wire[1916]) );
  DFF \memory_reg[59][27]  ( .D(n5869), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1915]), .Q(data_mem_out_wire[1915]) );
  DFF \memory_reg[59][26]  ( .D(n5868), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1914]), .Q(data_mem_out_wire[1914]) );
  DFF \memory_reg[59][25]  ( .D(n5867), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1913]), .Q(data_mem_out_wire[1913]) );
  DFF \memory_reg[59][24]  ( .D(n5866), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1912]), .Q(data_mem_out_wire[1912]) );
  DFF \memory_reg[59][23]  ( .D(n5865), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1911]), .Q(data_mem_out_wire[1911]) );
  DFF \memory_reg[59][22]  ( .D(n5864), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1910]), .Q(data_mem_out_wire[1910]) );
  DFF \memory_reg[59][21]  ( .D(n5863), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1909]), .Q(data_mem_out_wire[1909]) );
  DFF \memory_reg[59][20]  ( .D(n5862), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1908]), .Q(data_mem_out_wire[1908]) );
  DFF \memory_reg[59][19]  ( .D(n5861), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1907]), .Q(data_mem_out_wire[1907]) );
  DFF \memory_reg[59][18]  ( .D(n5860), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1906]), .Q(data_mem_out_wire[1906]) );
  DFF \memory_reg[59][17]  ( .D(n5859), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1905]), .Q(data_mem_out_wire[1905]) );
  DFF \memory_reg[59][16]  ( .D(n5858), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1904]), .Q(data_mem_out_wire[1904]) );
  DFF \memory_reg[59][15]  ( .D(n5857), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1903]), .Q(data_mem_out_wire[1903]) );
  DFF \memory_reg[59][14]  ( .D(n5856), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1902]), .Q(data_mem_out_wire[1902]) );
  DFF \memory_reg[59][13]  ( .D(n5855), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1901]), .Q(data_mem_out_wire[1901]) );
  DFF \memory_reg[59][12]  ( .D(n5854), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1900]), .Q(data_mem_out_wire[1900]) );
  DFF \memory_reg[59][11]  ( .D(n5853), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1899]), .Q(data_mem_out_wire[1899]) );
  DFF \memory_reg[59][10]  ( .D(n5852), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1898]), .Q(data_mem_out_wire[1898]) );
  DFF \memory_reg[59][9]  ( .D(n5851), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1897]), .Q(data_mem_out_wire[1897]) );
  DFF \memory_reg[59][8]  ( .D(n5850), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1896]), .Q(data_mem_out_wire[1896]) );
  DFF \memory_reg[59][7]  ( .D(n5849), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1895]), .Q(data_mem_out_wire[1895]) );
  DFF \memory_reg[59][6]  ( .D(n5848), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1894]), .Q(data_mem_out_wire[1894]) );
  DFF \memory_reg[59][5]  ( .D(n5847), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1893]), .Q(data_mem_out_wire[1893]) );
  DFF \memory_reg[59][4]  ( .D(n5846), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1892]), .Q(data_mem_out_wire[1892]) );
  DFF \memory_reg[59][3]  ( .D(n5845), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1891]), .Q(data_mem_out_wire[1891]) );
  DFF \memory_reg[59][2]  ( .D(n5844), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1890]), .Q(data_mem_out_wire[1890]) );
  DFF \memory_reg[59][1]  ( .D(n5843), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1889]), .Q(data_mem_out_wire[1889]) );
  DFF \memory_reg[59][0]  ( .D(n5842), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1888]), .Q(data_mem_out_wire[1888]) );
  DFF \memory_reg[60][31]  ( .D(n5841), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1951]), .Q(data_mem_out_wire[1951]) );
  DFF \memory_reg[60][30]  ( .D(n5840), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1950]), .Q(data_mem_out_wire[1950]) );
  DFF \memory_reg[60][29]  ( .D(n5839), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1949]), .Q(data_mem_out_wire[1949]) );
  DFF \memory_reg[60][28]  ( .D(n5838), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1948]), .Q(data_mem_out_wire[1948]) );
  DFF \memory_reg[60][27]  ( .D(n5837), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1947]), .Q(data_mem_out_wire[1947]) );
  DFF \memory_reg[60][26]  ( .D(n5836), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1946]), .Q(data_mem_out_wire[1946]) );
  DFF \memory_reg[60][25]  ( .D(n5835), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1945]), .Q(data_mem_out_wire[1945]) );
  DFF \memory_reg[60][24]  ( .D(n5834), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1944]), .Q(data_mem_out_wire[1944]) );
  DFF \memory_reg[60][23]  ( .D(n5833), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1943]), .Q(data_mem_out_wire[1943]) );
  DFF \memory_reg[60][22]  ( .D(n5832), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1942]), .Q(data_mem_out_wire[1942]) );
  DFF \memory_reg[60][21]  ( .D(n5831), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1941]), .Q(data_mem_out_wire[1941]) );
  DFF \memory_reg[60][20]  ( .D(n5830), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1940]), .Q(data_mem_out_wire[1940]) );
  DFF \memory_reg[60][19]  ( .D(n5829), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1939]), .Q(data_mem_out_wire[1939]) );
  DFF \memory_reg[60][18]  ( .D(n5828), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1938]), .Q(data_mem_out_wire[1938]) );
  DFF \memory_reg[60][17]  ( .D(n5827), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1937]), .Q(data_mem_out_wire[1937]) );
  DFF \memory_reg[60][16]  ( .D(n5826), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1936]), .Q(data_mem_out_wire[1936]) );
  DFF \memory_reg[60][15]  ( .D(n5825), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1935]), .Q(data_mem_out_wire[1935]) );
  DFF \memory_reg[60][14]  ( .D(n5824), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1934]), .Q(data_mem_out_wire[1934]) );
  DFF \memory_reg[60][13]  ( .D(n5823), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1933]), .Q(data_mem_out_wire[1933]) );
  DFF \memory_reg[60][12]  ( .D(n5822), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1932]), .Q(data_mem_out_wire[1932]) );
  DFF \memory_reg[60][11]  ( .D(n5821), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1931]), .Q(data_mem_out_wire[1931]) );
  DFF \memory_reg[60][10]  ( .D(n5820), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1930]), .Q(data_mem_out_wire[1930]) );
  DFF \memory_reg[60][9]  ( .D(n5819), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1929]), .Q(data_mem_out_wire[1929]) );
  DFF \memory_reg[60][8]  ( .D(n5818), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1928]), .Q(data_mem_out_wire[1928]) );
  DFF \memory_reg[60][7]  ( .D(n5817), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1927]), .Q(data_mem_out_wire[1927]) );
  DFF \memory_reg[60][6]  ( .D(n5816), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1926]), .Q(data_mem_out_wire[1926]) );
  DFF \memory_reg[60][5]  ( .D(n5815), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1925]), .Q(data_mem_out_wire[1925]) );
  DFF \memory_reg[60][4]  ( .D(n5814), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1924]), .Q(data_mem_out_wire[1924]) );
  DFF \memory_reg[60][3]  ( .D(n5813), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1923]), .Q(data_mem_out_wire[1923]) );
  DFF \memory_reg[60][2]  ( .D(n5812), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1922]), .Q(data_mem_out_wire[1922]) );
  DFF \memory_reg[60][1]  ( .D(n5811), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1921]), .Q(data_mem_out_wire[1921]) );
  DFF \memory_reg[60][0]  ( .D(n5810), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1920]), .Q(data_mem_out_wire[1920]) );
  DFF \memory_reg[61][31]  ( .D(n5809), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1983]), .Q(data_mem_out_wire[1983]) );
  DFF \memory_reg[61][30]  ( .D(n5808), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1982]), .Q(data_mem_out_wire[1982]) );
  DFF \memory_reg[61][29]  ( .D(n5807), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1981]), .Q(data_mem_out_wire[1981]) );
  DFF \memory_reg[61][28]  ( .D(n5806), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1980]), .Q(data_mem_out_wire[1980]) );
  DFF \memory_reg[61][27]  ( .D(n5805), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1979]), .Q(data_mem_out_wire[1979]) );
  DFF \memory_reg[61][26]  ( .D(n5804), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1978]), .Q(data_mem_out_wire[1978]) );
  DFF \memory_reg[61][25]  ( .D(n5803), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1977]), .Q(data_mem_out_wire[1977]) );
  DFF \memory_reg[61][24]  ( .D(n5802), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1976]), .Q(data_mem_out_wire[1976]) );
  DFF \memory_reg[61][23]  ( .D(n5801), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1975]), .Q(data_mem_out_wire[1975]) );
  DFF \memory_reg[61][22]  ( .D(n5800), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1974]), .Q(data_mem_out_wire[1974]) );
  DFF \memory_reg[61][21]  ( .D(n5799), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1973]), .Q(data_mem_out_wire[1973]) );
  DFF \memory_reg[61][20]  ( .D(n5798), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1972]), .Q(data_mem_out_wire[1972]) );
  DFF \memory_reg[61][19]  ( .D(n5797), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1971]), .Q(data_mem_out_wire[1971]) );
  DFF \memory_reg[61][18]  ( .D(n5796), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1970]), .Q(data_mem_out_wire[1970]) );
  DFF \memory_reg[61][17]  ( .D(n5795), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1969]), .Q(data_mem_out_wire[1969]) );
  DFF \memory_reg[61][16]  ( .D(n5794), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1968]), .Q(data_mem_out_wire[1968]) );
  DFF \memory_reg[61][15]  ( .D(n5793), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1967]), .Q(data_mem_out_wire[1967]) );
  DFF \memory_reg[61][14]  ( .D(n5792), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1966]), .Q(data_mem_out_wire[1966]) );
  DFF \memory_reg[61][13]  ( .D(n5791), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1965]), .Q(data_mem_out_wire[1965]) );
  DFF \memory_reg[61][12]  ( .D(n5790), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1964]), .Q(data_mem_out_wire[1964]) );
  DFF \memory_reg[61][11]  ( .D(n5789), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1963]), .Q(data_mem_out_wire[1963]) );
  DFF \memory_reg[61][10]  ( .D(n5788), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1962]), .Q(data_mem_out_wire[1962]) );
  DFF \memory_reg[61][9]  ( .D(n5787), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1961]), .Q(data_mem_out_wire[1961]) );
  DFF \memory_reg[61][8]  ( .D(n5786), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1960]), .Q(data_mem_out_wire[1960]) );
  DFF \memory_reg[61][7]  ( .D(n5785), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1959]), .Q(data_mem_out_wire[1959]) );
  DFF \memory_reg[61][6]  ( .D(n5784), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1958]), .Q(data_mem_out_wire[1958]) );
  DFF \memory_reg[61][5]  ( .D(n5783), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1957]), .Q(data_mem_out_wire[1957]) );
  DFF \memory_reg[61][4]  ( .D(n5782), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1956]), .Q(data_mem_out_wire[1956]) );
  DFF \memory_reg[61][3]  ( .D(n5781), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1955]), .Q(data_mem_out_wire[1955]) );
  DFF \memory_reg[61][2]  ( .D(n5780), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1954]), .Q(data_mem_out_wire[1954]) );
  DFF \memory_reg[61][1]  ( .D(n5779), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1953]), .Q(data_mem_out_wire[1953]) );
  DFF \memory_reg[61][0]  ( .D(n5778), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1952]), .Q(data_mem_out_wire[1952]) );
  DFF \memory_reg[62][31]  ( .D(n5777), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2015]), .Q(data_mem_out_wire[2015]) );
  DFF \memory_reg[62][30]  ( .D(n5776), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2014]), .Q(data_mem_out_wire[2014]) );
  DFF \memory_reg[62][29]  ( .D(n5775), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2013]), .Q(data_mem_out_wire[2013]) );
  DFF \memory_reg[62][28]  ( .D(n5774), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2012]), .Q(data_mem_out_wire[2012]) );
  DFF \memory_reg[62][27]  ( .D(n5773), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2011]), .Q(data_mem_out_wire[2011]) );
  DFF \memory_reg[62][26]  ( .D(n5772), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2010]), .Q(data_mem_out_wire[2010]) );
  DFF \memory_reg[62][25]  ( .D(n5771), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2009]), .Q(data_mem_out_wire[2009]) );
  DFF \memory_reg[62][24]  ( .D(n5770), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2008]), .Q(data_mem_out_wire[2008]) );
  DFF \memory_reg[62][23]  ( .D(n5769), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2007]), .Q(data_mem_out_wire[2007]) );
  DFF \memory_reg[62][22]  ( .D(n5768), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2006]), .Q(data_mem_out_wire[2006]) );
  DFF \memory_reg[62][21]  ( .D(n5767), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2005]), .Q(data_mem_out_wire[2005]) );
  DFF \memory_reg[62][20]  ( .D(n5766), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2004]), .Q(data_mem_out_wire[2004]) );
  DFF \memory_reg[62][19]  ( .D(n5765), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2003]), .Q(data_mem_out_wire[2003]) );
  DFF \memory_reg[62][18]  ( .D(n5764), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2002]), .Q(data_mem_out_wire[2002]) );
  DFF \memory_reg[62][17]  ( .D(n5763), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2001]), .Q(data_mem_out_wire[2001]) );
  DFF \memory_reg[62][16]  ( .D(n5762), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2000]), .Q(data_mem_out_wire[2000]) );
  DFF \memory_reg[62][15]  ( .D(n5761), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1999]), .Q(data_mem_out_wire[1999]) );
  DFF \memory_reg[62][14]  ( .D(n5760), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1998]), .Q(data_mem_out_wire[1998]) );
  DFF \memory_reg[62][13]  ( .D(n5759), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1997]), .Q(data_mem_out_wire[1997]) );
  DFF \memory_reg[62][12]  ( .D(n5758), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1996]), .Q(data_mem_out_wire[1996]) );
  DFF \memory_reg[62][11]  ( .D(n5757), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1995]), .Q(data_mem_out_wire[1995]) );
  DFF \memory_reg[62][10]  ( .D(n5756), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1994]), .Q(data_mem_out_wire[1994]) );
  DFF \memory_reg[62][9]  ( .D(n5755), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1993]), .Q(data_mem_out_wire[1993]) );
  DFF \memory_reg[62][8]  ( .D(n5754), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1992]), .Q(data_mem_out_wire[1992]) );
  DFF \memory_reg[62][7]  ( .D(n5753), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1991]), .Q(data_mem_out_wire[1991]) );
  DFF \memory_reg[62][6]  ( .D(n5752), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1990]), .Q(data_mem_out_wire[1990]) );
  DFF \memory_reg[62][5]  ( .D(n5751), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1989]), .Q(data_mem_out_wire[1989]) );
  DFF \memory_reg[62][4]  ( .D(n5750), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1988]), .Q(data_mem_out_wire[1988]) );
  DFF \memory_reg[62][3]  ( .D(n5749), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1987]), .Q(data_mem_out_wire[1987]) );
  DFF \memory_reg[62][2]  ( .D(n5748), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1986]), .Q(data_mem_out_wire[1986]) );
  DFF \memory_reg[62][1]  ( .D(n5747), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1985]), .Q(data_mem_out_wire[1985]) );
  DFF \memory_reg[62][0]  ( .D(n5746), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[1984]), .Q(data_mem_out_wire[1984]) );
  DFF \memory_reg[63][31]  ( .D(n5745), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2047]), .Q(data_mem_out_wire[2047]) );
  DFF \memory_reg[63][30]  ( .D(n5744), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2046]), .Q(data_mem_out_wire[2046]) );
  DFF \memory_reg[63][29]  ( .D(n5743), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2045]), .Q(data_mem_out_wire[2045]) );
  DFF \memory_reg[63][28]  ( .D(n5742), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2044]), .Q(data_mem_out_wire[2044]) );
  DFF \memory_reg[63][27]  ( .D(n5741), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2043]), .Q(data_mem_out_wire[2043]) );
  DFF \memory_reg[63][26]  ( .D(n5740), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2042]), .Q(data_mem_out_wire[2042]) );
  DFF \memory_reg[63][25]  ( .D(n5739), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2041]), .Q(data_mem_out_wire[2041]) );
  DFF \memory_reg[63][24]  ( .D(n5738), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2040]), .Q(data_mem_out_wire[2040]) );
  DFF \memory_reg[63][23]  ( .D(n5737), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2039]), .Q(data_mem_out_wire[2039]) );
  DFF \memory_reg[63][22]  ( .D(n5736), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2038]), .Q(data_mem_out_wire[2038]) );
  DFF \memory_reg[63][21]  ( .D(n5735), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2037]), .Q(data_mem_out_wire[2037]) );
  DFF \memory_reg[63][20]  ( .D(n5734), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2036]), .Q(data_mem_out_wire[2036]) );
  DFF \memory_reg[63][19]  ( .D(n5733), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2035]), .Q(data_mem_out_wire[2035]) );
  DFF \memory_reg[63][18]  ( .D(n5732), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2034]), .Q(data_mem_out_wire[2034]) );
  DFF \memory_reg[63][17]  ( .D(n5731), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2033]), .Q(data_mem_out_wire[2033]) );
  DFF \memory_reg[63][16]  ( .D(n5730), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2032]), .Q(data_mem_out_wire[2032]) );
  DFF \memory_reg[63][15]  ( .D(n5729), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2031]), .Q(data_mem_out_wire[2031]) );
  DFF \memory_reg[63][14]  ( .D(n5728), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2030]), .Q(data_mem_out_wire[2030]) );
  DFF \memory_reg[63][13]  ( .D(n5727), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2029]), .Q(data_mem_out_wire[2029]) );
  DFF \memory_reg[63][12]  ( .D(n5726), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2028]), .Q(data_mem_out_wire[2028]) );
  DFF \memory_reg[63][11]  ( .D(n5725), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2027]), .Q(data_mem_out_wire[2027]) );
  DFF \memory_reg[63][10]  ( .D(n5724), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2026]), .Q(data_mem_out_wire[2026]) );
  DFF \memory_reg[63][9]  ( .D(n5723), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2025]), .Q(data_mem_out_wire[2025]) );
  DFF \memory_reg[63][8]  ( .D(n5722), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2024]), .Q(data_mem_out_wire[2024]) );
  DFF \memory_reg[63][7]  ( .D(n5721), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2023]), .Q(data_mem_out_wire[2023]) );
  DFF \memory_reg[63][6]  ( .D(n5720), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2022]), .Q(data_mem_out_wire[2022]) );
  DFF \memory_reg[63][5]  ( .D(n5719), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2021]), .Q(data_mem_out_wire[2021]) );
  DFF \memory_reg[63][4]  ( .D(n5718), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2020]), .Q(data_mem_out_wire[2020]) );
  DFF \memory_reg[63][3]  ( .D(n5717), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2019]), .Q(data_mem_out_wire[2019]) );
  DFF \memory_reg[63][2]  ( .D(n5716), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2018]), .Q(data_mem_out_wire[2018]) );
  DFF \memory_reg[63][1]  ( .D(n5715), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2017]), .Q(data_mem_out_wire[2017]) );
  DFF \memory_reg[63][0]  ( .D(n5714), .CLK(clk), .RST(rst), .I(
        data_mem_in_wire[2016]), .Q(data_mem_out_wire[2016]) );
  MUX U7795 ( .IN0(data_mem_out_wire[1984]), .IN1(data_mem_out_wire[2016]), 
        .SEL(N37), .F(n7762) );
  MUX U7796 ( .IN0(data_mem_out_wire[1920]), .IN1(data_mem_out_wire[1952]), 
        .SEL(N37), .F(n7763) );
  MUX U7797 ( .IN0(n7763), .IN1(n7762), .SEL(N38), .F(n7764) );
  MUX U7798 ( .IN0(data_mem_out_wire[1856]), .IN1(data_mem_out_wire[1888]), 
        .SEL(N37), .F(n7765) );
  MUX U7799 ( .IN0(data_mem_out_wire[1792]), .IN1(data_mem_out_wire[1824]), 
        .SEL(N37), .F(n7766) );
  MUX U7800 ( .IN0(n7766), .IN1(n7765), .SEL(N38), .F(n7767) );
  MUX U7801 ( .IN0(n7767), .IN1(n7764), .SEL(N39), .F(n7768) );
  MUX U7802 ( .IN0(data_mem_out_wire[1728]), .IN1(data_mem_out_wire[1760]), 
        .SEL(N37), .F(n7769) );
  MUX U7803 ( .IN0(data_mem_out_wire[1664]), .IN1(data_mem_out_wire[1696]), 
        .SEL(N37), .F(n7770) );
  MUX U7804 ( .IN0(n7770), .IN1(n7769), .SEL(N38), .F(n7771) );
  MUX U7805 ( .IN0(data_mem_out_wire[1600]), .IN1(data_mem_out_wire[1632]), 
        .SEL(N37), .F(n7772) );
  MUX U7806 ( .IN0(data_mem_out_wire[1536]), .IN1(data_mem_out_wire[1568]), 
        .SEL(N37), .F(n7773) );
  MUX U7807 ( .IN0(n7773), .IN1(n7772), .SEL(N38), .F(n7774) );
  MUX U7808 ( .IN0(n7774), .IN1(n7771), .SEL(N39), .F(n7775) );
  MUX U7809 ( .IN0(n7775), .IN1(n7768), .SEL(N40), .F(n7776) );
  MUX U7810 ( .IN0(data_mem_out_wire[1472]), .IN1(data_mem_out_wire[1504]), 
        .SEL(N37), .F(n7777) );
  MUX U7811 ( .IN0(data_mem_out_wire[1408]), .IN1(data_mem_out_wire[1440]), 
        .SEL(N37), .F(n7778) );
  MUX U7812 ( .IN0(n7778), .IN1(n7777), .SEL(N38), .F(n7779) );
  MUX U7813 ( .IN0(data_mem_out_wire[1344]), .IN1(data_mem_out_wire[1376]), 
        .SEL(N37), .F(n7780) );
  MUX U7814 ( .IN0(data_mem_out_wire[1280]), .IN1(data_mem_out_wire[1312]), 
        .SEL(N37), .F(n7781) );
  MUX U7815 ( .IN0(n7781), .IN1(n7780), .SEL(N38), .F(n7782) );
  MUX U7816 ( .IN0(n7782), .IN1(n7779), .SEL(N39), .F(n7783) );
  MUX U7817 ( .IN0(data_mem_out_wire[1216]), .IN1(data_mem_out_wire[1248]), 
        .SEL(N37), .F(n7784) );
  MUX U7818 ( .IN0(data_mem_out_wire[1152]), .IN1(data_mem_out_wire[1184]), 
        .SEL(N37), .F(n7785) );
  MUX U7819 ( .IN0(n7785), .IN1(n7784), .SEL(N38), .F(n7786) );
  MUX U7820 ( .IN0(data_mem_out_wire[1088]), .IN1(data_mem_out_wire[1120]), 
        .SEL(N37), .F(n7787) );
  MUX U7821 ( .IN0(data_mem_out_wire[1024]), .IN1(data_mem_out_wire[1056]), 
        .SEL(N37), .F(n7788) );
  MUX U7822 ( .IN0(n7788), .IN1(n7787), .SEL(N38), .F(n7789) );
  MUX U7823 ( .IN0(n7789), .IN1(n7786), .SEL(N39), .F(n7790) );
  MUX U7824 ( .IN0(n7790), .IN1(n7783), .SEL(N40), .F(n7791) );
  MUX U7825 ( .IN0(n7791), .IN1(n7776), .SEL(N41), .F(n7792) );
  MUX U7826 ( .IN0(data_mem_out_wire[960]), .IN1(data_mem_out_wire[992]), 
        .SEL(N37), .F(n7793) );
  MUX U7827 ( .IN0(data_mem_out_wire[896]), .IN1(data_mem_out_wire[928]), 
        .SEL(N37), .F(n7794) );
  MUX U7828 ( .IN0(n7794), .IN1(n7793), .SEL(N38), .F(n7795) );
  MUX U7829 ( .IN0(data_mem_out_wire[832]), .IN1(data_mem_out_wire[864]), 
        .SEL(N37), .F(n7796) );
  MUX U7830 ( .IN0(data_mem_out_wire[768]), .IN1(data_mem_out_wire[800]), 
        .SEL(N37), .F(n7797) );
  MUX U7831 ( .IN0(n7797), .IN1(n7796), .SEL(N38), .F(n7798) );
  MUX U7832 ( .IN0(n7798), .IN1(n7795), .SEL(N39), .F(n7799) );
  MUX U7833 ( .IN0(data_mem_out_wire[704]), .IN1(data_mem_out_wire[736]), 
        .SEL(N37), .F(n7800) );
  MUX U7834 ( .IN0(data_mem_out_wire[640]), .IN1(data_mem_out_wire[672]), 
        .SEL(N37), .F(n7801) );
  MUX U7835 ( .IN0(n7801), .IN1(n7800), .SEL(N38), .F(n7802) );
  MUX U7836 ( .IN0(data_mem_out_wire[576]), .IN1(data_mem_out_wire[608]), 
        .SEL(N37), .F(n7803) );
  MUX U7837 ( .IN0(data_mem_out_wire[512]), .IN1(data_mem_out_wire[544]), 
        .SEL(N37), .F(n7804) );
  MUX U7838 ( .IN0(n7804), .IN1(n7803), .SEL(N38), .F(n7805) );
  MUX U7839 ( .IN0(n7805), .IN1(n7802), .SEL(N39), .F(n7806) );
  MUX U7840 ( .IN0(n7806), .IN1(n7799), .SEL(N40), .F(n7807) );
  MUX U7841 ( .IN0(data_mem_out_wire[448]), .IN1(data_mem_out_wire[480]), 
        .SEL(N37), .F(n7808) );
  MUX U7842 ( .IN0(data_mem_out_wire[384]), .IN1(data_mem_out_wire[416]), 
        .SEL(N37), .F(n7809) );
  MUX U7843 ( .IN0(n7809), .IN1(n7808), .SEL(N38), .F(n7810) );
  MUX U7844 ( .IN0(data_mem_out_wire[320]), .IN1(data_mem_out_wire[352]), 
        .SEL(N37), .F(n7811) );
  MUX U7845 ( .IN0(data_mem_out_wire[256]), .IN1(data_mem_out_wire[288]), 
        .SEL(N37), .F(n7812) );
  MUX U7846 ( .IN0(n7812), .IN1(n7811), .SEL(N38), .F(n7813) );
  MUX U7847 ( .IN0(n7813), .IN1(n7810), .SEL(N39), .F(n7814) );
  MUX U7848 ( .IN0(data_mem_out_wire[192]), .IN1(data_mem_out_wire[224]), 
        .SEL(N37), .F(n7815) );
  MUX U7849 ( .IN0(data_mem_out_wire[128]), .IN1(data_mem_out_wire[160]), 
        .SEL(N37), .F(n7816) );
  MUX U7850 ( .IN0(n7816), .IN1(n7815), .SEL(N38), .F(n7817) );
  MUX U7851 ( .IN0(data_mem_out_wire[64]), .IN1(data_mem_out_wire[96]), .SEL(
        N37), .F(n7818) );
  MUX U7852 ( .IN0(data_mem_out_wire[0]), .IN1(data_mem_out_wire[32]), .SEL(
        N37), .F(n7819) );
  MUX U7853 ( .IN0(n7819), .IN1(n7818), .SEL(N38), .F(n7820) );
  MUX U7854 ( .IN0(n7820), .IN1(n7817), .SEL(N39), .F(n7821) );
  MUX U7855 ( .IN0(n7821), .IN1(n7814), .SEL(N40), .F(n7822) );
  MUX U7856 ( .IN0(n7822), .IN1(n7807), .SEL(N41), .F(n7823) );
  MUX U7857 ( .IN0(n7823), .IN1(n7792), .SEL(N42), .F(N745) );
  MUX U7858 ( .IN0(data_mem_out_wire[1985]), .IN1(data_mem_out_wire[2017]), 
        .SEL(N37), .F(n7824) );
  MUX U7859 ( .IN0(data_mem_out_wire[1921]), .IN1(data_mem_out_wire[1953]), 
        .SEL(N37), .F(n7825) );
  MUX U7860 ( .IN0(n7825), .IN1(n7824), .SEL(N38), .F(n7826) );
  MUX U7861 ( .IN0(data_mem_out_wire[1857]), .IN1(data_mem_out_wire[1889]), 
        .SEL(N37), .F(n7827) );
  MUX U7862 ( .IN0(data_mem_out_wire[1793]), .IN1(data_mem_out_wire[1825]), 
        .SEL(N37), .F(n7828) );
  MUX U7863 ( .IN0(n7828), .IN1(n7827), .SEL(N38), .F(n7829) );
  MUX U7864 ( .IN0(n7829), .IN1(n7826), .SEL(N39), .F(n7830) );
  MUX U7865 ( .IN0(data_mem_out_wire[1729]), .IN1(data_mem_out_wire[1761]), 
        .SEL(N37), .F(n7831) );
  MUX U7866 ( .IN0(data_mem_out_wire[1665]), .IN1(data_mem_out_wire[1697]), 
        .SEL(N37), .F(n7832) );
  MUX U7867 ( .IN0(n7832), .IN1(n7831), .SEL(N38), .F(n7833) );
  MUX U7868 ( .IN0(data_mem_out_wire[1601]), .IN1(data_mem_out_wire[1633]), 
        .SEL(N37), .F(n7834) );
  MUX U7869 ( .IN0(data_mem_out_wire[1537]), .IN1(data_mem_out_wire[1569]), 
        .SEL(N37), .F(n7835) );
  MUX U7870 ( .IN0(n7835), .IN1(n7834), .SEL(N38), .F(n7836) );
  MUX U7871 ( .IN0(n7836), .IN1(n7833), .SEL(N39), .F(n7837) );
  MUX U7872 ( .IN0(n7837), .IN1(n7830), .SEL(N40), .F(n7838) );
  MUX U7873 ( .IN0(data_mem_out_wire[1473]), .IN1(data_mem_out_wire[1505]), 
        .SEL(N37), .F(n7839) );
  MUX U7874 ( .IN0(data_mem_out_wire[1409]), .IN1(data_mem_out_wire[1441]), 
        .SEL(N37), .F(n7840) );
  MUX U7875 ( .IN0(n7840), .IN1(n7839), .SEL(N38), .F(n7841) );
  MUX U7876 ( .IN0(data_mem_out_wire[1345]), .IN1(data_mem_out_wire[1377]), 
        .SEL(N37), .F(n7842) );
  MUX U7877 ( .IN0(data_mem_out_wire[1281]), .IN1(data_mem_out_wire[1313]), 
        .SEL(N37), .F(n7843) );
  MUX U7878 ( .IN0(n7843), .IN1(n7842), .SEL(N38), .F(n7844) );
  MUX U7879 ( .IN0(n7844), .IN1(n7841), .SEL(N39), .F(n7845) );
  MUX U7880 ( .IN0(data_mem_out_wire[1217]), .IN1(data_mem_out_wire[1249]), 
        .SEL(N37), .F(n7846) );
  MUX U7881 ( .IN0(data_mem_out_wire[1153]), .IN1(data_mem_out_wire[1185]), 
        .SEL(N37), .F(n7847) );
  MUX U7882 ( .IN0(n7847), .IN1(n7846), .SEL(N38), .F(n7848) );
  MUX U7883 ( .IN0(data_mem_out_wire[1089]), .IN1(data_mem_out_wire[1121]), 
        .SEL(N37), .F(n7849) );
  MUX U7884 ( .IN0(data_mem_out_wire[1025]), .IN1(data_mem_out_wire[1057]), 
        .SEL(N37), .F(n7850) );
  MUX U7885 ( .IN0(n7850), .IN1(n7849), .SEL(N38), .F(n7851) );
  MUX U7886 ( .IN0(n7851), .IN1(n7848), .SEL(N39), .F(n7852) );
  MUX U7887 ( .IN0(n7852), .IN1(n7845), .SEL(N40), .F(n7853) );
  MUX U7888 ( .IN0(n7853), .IN1(n7838), .SEL(N41), .F(n7854) );
  MUX U7889 ( .IN0(data_mem_out_wire[961]), .IN1(data_mem_out_wire[993]), 
        .SEL(N37), .F(n7855) );
  MUX U7890 ( .IN0(data_mem_out_wire[897]), .IN1(data_mem_out_wire[929]), 
        .SEL(N37), .F(n7856) );
  MUX U7891 ( .IN0(n7856), .IN1(n7855), .SEL(N38), .F(n7857) );
  MUX U7892 ( .IN0(data_mem_out_wire[833]), .IN1(data_mem_out_wire[865]), 
        .SEL(N37), .F(n7858) );
  MUX U7893 ( .IN0(data_mem_out_wire[769]), .IN1(data_mem_out_wire[801]), 
        .SEL(N37), .F(n7859) );
  MUX U7894 ( .IN0(n7859), .IN1(n7858), .SEL(N38), .F(n7860) );
  MUX U7895 ( .IN0(n7860), .IN1(n7857), .SEL(N39), .F(n7861) );
  MUX U7896 ( .IN0(data_mem_out_wire[705]), .IN1(data_mem_out_wire[737]), 
        .SEL(N37), .F(n7862) );
  MUX U7897 ( .IN0(data_mem_out_wire[641]), .IN1(data_mem_out_wire[673]), 
        .SEL(N37), .F(n7863) );
  MUX U7898 ( .IN0(n7863), .IN1(n7862), .SEL(N38), .F(n7864) );
  MUX U7899 ( .IN0(data_mem_out_wire[577]), .IN1(data_mem_out_wire[609]), 
        .SEL(N37), .F(n7865) );
  MUX U7900 ( .IN0(data_mem_out_wire[513]), .IN1(data_mem_out_wire[545]), 
        .SEL(N37), .F(n7866) );
  MUX U7901 ( .IN0(n7866), .IN1(n7865), .SEL(N38), .F(n7867) );
  MUX U7902 ( .IN0(n7867), .IN1(n7864), .SEL(N39), .F(n7868) );
  MUX U7903 ( .IN0(n7868), .IN1(n7861), .SEL(N40), .F(n7869) );
  MUX U7904 ( .IN0(data_mem_out_wire[449]), .IN1(data_mem_out_wire[481]), 
        .SEL(N37), .F(n7870) );
  MUX U7905 ( .IN0(data_mem_out_wire[385]), .IN1(data_mem_out_wire[417]), 
        .SEL(N37), .F(n7871) );
  MUX U7906 ( .IN0(n7871), .IN1(n7870), .SEL(N38), .F(n7872) );
  MUX U7907 ( .IN0(data_mem_out_wire[321]), .IN1(data_mem_out_wire[353]), 
        .SEL(N37), .F(n7873) );
  MUX U7908 ( .IN0(data_mem_out_wire[257]), .IN1(data_mem_out_wire[289]), 
        .SEL(N37), .F(n7874) );
  MUX U7909 ( .IN0(n7874), .IN1(n7873), .SEL(N38), .F(n7875) );
  MUX U7910 ( .IN0(n7875), .IN1(n7872), .SEL(N39), .F(n7876) );
  MUX U7911 ( .IN0(data_mem_out_wire[193]), .IN1(data_mem_out_wire[225]), 
        .SEL(N37), .F(n7877) );
  MUX U7912 ( .IN0(data_mem_out_wire[129]), .IN1(data_mem_out_wire[161]), 
        .SEL(N37), .F(n7878) );
  MUX U7913 ( .IN0(n7878), .IN1(n7877), .SEL(N38), .F(n7879) );
  MUX U7914 ( .IN0(data_mem_out_wire[65]), .IN1(data_mem_out_wire[97]), .SEL(
        N37), .F(n7880) );
  MUX U7915 ( .IN0(data_mem_out_wire[1]), .IN1(data_mem_out_wire[33]), .SEL(
        N37), .F(n7881) );
  MUX U7916 ( .IN0(n7881), .IN1(n7880), .SEL(N38), .F(n7882) );
  MUX U7917 ( .IN0(n7882), .IN1(n7879), .SEL(N39), .F(n7883) );
  MUX U7918 ( .IN0(n7883), .IN1(n7876), .SEL(N40), .F(n7884) );
  MUX U7919 ( .IN0(n7884), .IN1(n7869), .SEL(N41), .F(n7885) );
  MUX U7920 ( .IN0(n7885), .IN1(n7854), .SEL(N42), .F(N744) );
  MUX U7921 ( .IN0(data_mem_out_wire[1986]), .IN1(data_mem_out_wire[2018]), 
        .SEL(N37), .F(n7886) );
  MUX U7922 ( .IN0(data_mem_out_wire[1922]), .IN1(data_mem_out_wire[1954]), 
        .SEL(N37), .F(n7887) );
  MUX U7923 ( .IN0(n7887), .IN1(n7886), .SEL(N38), .F(n7888) );
  MUX U7924 ( .IN0(data_mem_out_wire[1858]), .IN1(data_mem_out_wire[1890]), 
        .SEL(N37), .F(n7889) );
  MUX U7925 ( .IN0(data_mem_out_wire[1794]), .IN1(data_mem_out_wire[1826]), 
        .SEL(N37), .F(n7890) );
  MUX U7926 ( .IN0(n7890), .IN1(n7889), .SEL(N38), .F(n7891) );
  MUX U7927 ( .IN0(n7891), .IN1(n7888), .SEL(N39), .F(n7892) );
  MUX U7928 ( .IN0(data_mem_out_wire[1730]), .IN1(data_mem_out_wire[1762]), 
        .SEL(N37), .F(n7893) );
  MUX U7929 ( .IN0(data_mem_out_wire[1666]), .IN1(data_mem_out_wire[1698]), 
        .SEL(N37), .F(n7894) );
  MUX U7930 ( .IN0(n7894), .IN1(n7893), .SEL(N38), .F(n7895) );
  MUX U7931 ( .IN0(data_mem_out_wire[1602]), .IN1(data_mem_out_wire[1634]), 
        .SEL(N37), .F(n7896) );
  MUX U7932 ( .IN0(data_mem_out_wire[1538]), .IN1(data_mem_out_wire[1570]), 
        .SEL(N37), .F(n7897) );
  MUX U7933 ( .IN0(n7897), .IN1(n7896), .SEL(N38), .F(n7898) );
  MUX U7934 ( .IN0(n7898), .IN1(n7895), .SEL(N39), .F(n7899) );
  MUX U7935 ( .IN0(n7899), .IN1(n7892), .SEL(N40), .F(n7900) );
  MUX U7936 ( .IN0(data_mem_out_wire[1474]), .IN1(data_mem_out_wire[1506]), 
        .SEL(N37), .F(n7901) );
  MUX U7937 ( .IN0(data_mem_out_wire[1410]), .IN1(data_mem_out_wire[1442]), 
        .SEL(N37), .F(n7902) );
  MUX U7938 ( .IN0(n7902), .IN1(n7901), .SEL(N38), .F(n7903) );
  MUX U7939 ( .IN0(data_mem_out_wire[1346]), .IN1(data_mem_out_wire[1378]), 
        .SEL(N37), .F(n7904) );
  MUX U7940 ( .IN0(data_mem_out_wire[1282]), .IN1(data_mem_out_wire[1314]), 
        .SEL(N37), .F(n7905) );
  MUX U7941 ( .IN0(n7905), .IN1(n7904), .SEL(N38), .F(n7906) );
  MUX U7942 ( .IN0(n7906), .IN1(n7903), .SEL(N39), .F(n7907) );
  MUX U7943 ( .IN0(data_mem_out_wire[1218]), .IN1(data_mem_out_wire[1250]), 
        .SEL(N37), .F(n7908) );
  MUX U7944 ( .IN0(data_mem_out_wire[1154]), .IN1(data_mem_out_wire[1186]), 
        .SEL(N37), .F(n7909) );
  MUX U7945 ( .IN0(n7909), .IN1(n7908), .SEL(N38), .F(n7910) );
  MUX U7946 ( .IN0(data_mem_out_wire[1090]), .IN1(data_mem_out_wire[1122]), 
        .SEL(N37), .F(n7911) );
  MUX U7947 ( .IN0(data_mem_out_wire[1026]), .IN1(data_mem_out_wire[1058]), 
        .SEL(N37), .F(n7912) );
  MUX U7948 ( .IN0(n7912), .IN1(n7911), .SEL(N38), .F(n7913) );
  MUX U7949 ( .IN0(n7913), .IN1(n7910), .SEL(N39), .F(n7914) );
  MUX U7950 ( .IN0(n7914), .IN1(n7907), .SEL(N40), .F(n7915) );
  MUX U7951 ( .IN0(n7915), .IN1(n7900), .SEL(N41), .F(n7916) );
  MUX U7952 ( .IN0(data_mem_out_wire[962]), .IN1(data_mem_out_wire[994]), 
        .SEL(N37), .F(n7917) );
  MUX U7953 ( .IN0(data_mem_out_wire[898]), .IN1(data_mem_out_wire[930]), 
        .SEL(N37), .F(n7918) );
  MUX U7954 ( .IN0(n7918), .IN1(n7917), .SEL(N38), .F(n7919) );
  MUX U7955 ( .IN0(data_mem_out_wire[834]), .IN1(data_mem_out_wire[866]), 
        .SEL(N37), .F(n7920) );
  MUX U7956 ( .IN0(data_mem_out_wire[770]), .IN1(data_mem_out_wire[802]), 
        .SEL(N37), .F(n7921) );
  MUX U7957 ( .IN0(n7921), .IN1(n7920), .SEL(N38), .F(n7922) );
  MUX U7958 ( .IN0(n7922), .IN1(n7919), .SEL(N39), .F(n7923) );
  MUX U7959 ( .IN0(data_mem_out_wire[706]), .IN1(data_mem_out_wire[738]), 
        .SEL(N37), .F(n7924) );
  MUX U7960 ( .IN0(data_mem_out_wire[642]), .IN1(data_mem_out_wire[674]), 
        .SEL(N37), .F(n7925) );
  MUX U7961 ( .IN0(n7925), .IN1(n7924), .SEL(N38), .F(n7926) );
  MUX U7962 ( .IN0(data_mem_out_wire[578]), .IN1(data_mem_out_wire[610]), 
        .SEL(N37), .F(n7927) );
  MUX U7963 ( .IN0(data_mem_out_wire[514]), .IN1(data_mem_out_wire[546]), 
        .SEL(N37), .F(n7928) );
  MUX U7964 ( .IN0(n7928), .IN1(n7927), .SEL(N38), .F(n7929) );
  MUX U7965 ( .IN0(n7929), .IN1(n7926), .SEL(N39), .F(n7930) );
  MUX U7966 ( .IN0(n7930), .IN1(n7923), .SEL(N40), .F(n7931) );
  MUX U7967 ( .IN0(data_mem_out_wire[450]), .IN1(data_mem_out_wire[482]), 
        .SEL(N37), .F(n7932) );
  MUX U7968 ( .IN0(data_mem_out_wire[386]), .IN1(data_mem_out_wire[418]), 
        .SEL(N37), .F(n7933) );
  MUX U7969 ( .IN0(n7933), .IN1(n7932), .SEL(N38), .F(n7934) );
  MUX U7970 ( .IN0(data_mem_out_wire[322]), .IN1(data_mem_out_wire[354]), 
        .SEL(N37), .F(n7935) );
  MUX U7971 ( .IN0(data_mem_out_wire[258]), .IN1(data_mem_out_wire[290]), 
        .SEL(N37), .F(n7936) );
  MUX U7972 ( .IN0(n7936), .IN1(n7935), .SEL(N38), .F(n7937) );
  MUX U7973 ( .IN0(n7937), .IN1(n7934), .SEL(N39), .F(n7938) );
  MUX U7974 ( .IN0(data_mem_out_wire[194]), .IN1(data_mem_out_wire[226]), 
        .SEL(N37), .F(n7939) );
  MUX U7975 ( .IN0(data_mem_out_wire[130]), .IN1(data_mem_out_wire[162]), 
        .SEL(N37), .F(n7940) );
  MUX U7976 ( .IN0(n7940), .IN1(n7939), .SEL(N38), .F(n7941) );
  MUX U7977 ( .IN0(data_mem_out_wire[66]), .IN1(data_mem_out_wire[98]), .SEL(
        N37), .F(n7942) );
  MUX U7978 ( .IN0(data_mem_out_wire[2]), .IN1(data_mem_out_wire[34]), .SEL(
        N37), .F(n7943) );
  MUX U7979 ( .IN0(n7943), .IN1(n7942), .SEL(N38), .F(n7944) );
  MUX U7980 ( .IN0(n7944), .IN1(n7941), .SEL(N39), .F(n7945) );
  MUX U7981 ( .IN0(n7945), .IN1(n7938), .SEL(N40), .F(n7946) );
  MUX U7982 ( .IN0(n7946), .IN1(n7931), .SEL(N41), .F(n7947) );
  MUX U7983 ( .IN0(n7947), .IN1(n7916), .SEL(N42), .F(N743) );
  MUX U7984 ( .IN0(data_mem_out_wire[1987]), .IN1(data_mem_out_wire[2019]), 
        .SEL(N37), .F(n7948) );
  MUX U7985 ( .IN0(data_mem_out_wire[1923]), .IN1(data_mem_out_wire[1955]), 
        .SEL(N37), .F(n7949) );
  MUX U7986 ( .IN0(n7949), .IN1(n7948), .SEL(N38), .F(n7950) );
  MUX U7987 ( .IN0(data_mem_out_wire[1859]), .IN1(data_mem_out_wire[1891]), 
        .SEL(N37), .F(n7951) );
  MUX U7988 ( .IN0(data_mem_out_wire[1795]), .IN1(data_mem_out_wire[1827]), 
        .SEL(N37), .F(n7952) );
  MUX U7989 ( .IN0(n7952), .IN1(n7951), .SEL(N38), .F(n7953) );
  MUX U7990 ( .IN0(n7953), .IN1(n7950), .SEL(N39), .F(n7954) );
  MUX U7991 ( .IN0(data_mem_out_wire[1731]), .IN1(data_mem_out_wire[1763]), 
        .SEL(N37), .F(n7955) );
  MUX U7992 ( .IN0(data_mem_out_wire[1667]), .IN1(data_mem_out_wire[1699]), 
        .SEL(N37), .F(n7956) );
  MUX U7993 ( .IN0(n7956), .IN1(n7955), .SEL(N38), .F(n7957) );
  MUX U7994 ( .IN0(data_mem_out_wire[1603]), .IN1(data_mem_out_wire[1635]), 
        .SEL(N37), .F(n7958) );
  MUX U7995 ( .IN0(data_mem_out_wire[1539]), .IN1(data_mem_out_wire[1571]), 
        .SEL(N37), .F(n7959) );
  MUX U7996 ( .IN0(n7959), .IN1(n7958), .SEL(N38), .F(n7960) );
  MUX U7997 ( .IN0(n7960), .IN1(n7957), .SEL(N39), .F(n7961) );
  MUX U7998 ( .IN0(n7961), .IN1(n7954), .SEL(N40), .F(n7962) );
  MUX U7999 ( .IN0(data_mem_out_wire[1475]), .IN1(data_mem_out_wire[1507]), 
        .SEL(N37), .F(n7963) );
  MUX U8000 ( .IN0(data_mem_out_wire[1411]), .IN1(data_mem_out_wire[1443]), 
        .SEL(N37), .F(n7964) );
  MUX U8001 ( .IN0(n7964), .IN1(n7963), .SEL(N38), .F(n7965) );
  MUX U8002 ( .IN0(data_mem_out_wire[1347]), .IN1(data_mem_out_wire[1379]), 
        .SEL(N37), .F(n7966) );
  MUX U8003 ( .IN0(data_mem_out_wire[1283]), .IN1(data_mem_out_wire[1315]), 
        .SEL(N37), .F(n7967) );
  MUX U8004 ( .IN0(n7967), .IN1(n7966), .SEL(N38), .F(n7968) );
  MUX U8005 ( .IN0(n7968), .IN1(n7965), .SEL(N39), .F(n7969) );
  MUX U8006 ( .IN0(data_mem_out_wire[1219]), .IN1(data_mem_out_wire[1251]), 
        .SEL(N37), .F(n7970) );
  MUX U8007 ( .IN0(data_mem_out_wire[1155]), .IN1(data_mem_out_wire[1187]), 
        .SEL(N37), .F(n7971) );
  MUX U8008 ( .IN0(n7971), .IN1(n7970), .SEL(N38), .F(n7972) );
  MUX U8009 ( .IN0(data_mem_out_wire[1091]), .IN1(data_mem_out_wire[1123]), 
        .SEL(N37), .F(n7973) );
  MUX U8010 ( .IN0(data_mem_out_wire[1027]), .IN1(data_mem_out_wire[1059]), 
        .SEL(N37), .F(n7974) );
  MUX U8011 ( .IN0(n7974), .IN1(n7973), .SEL(N38), .F(n7975) );
  MUX U8012 ( .IN0(n7975), .IN1(n7972), .SEL(N39), .F(n7976) );
  MUX U8013 ( .IN0(n7976), .IN1(n7969), .SEL(N40), .F(n7977) );
  MUX U8014 ( .IN0(n7977), .IN1(n7962), .SEL(N41), .F(n7978) );
  MUX U8015 ( .IN0(data_mem_out_wire[963]), .IN1(data_mem_out_wire[995]), 
        .SEL(N37), .F(n7979) );
  MUX U8016 ( .IN0(data_mem_out_wire[899]), .IN1(data_mem_out_wire[931]), 
        .SEL(N37), .F(n7980) );
  MUX U8017 ( .IN0(n7980), .IN1(n7979), .SEL(N38), .F(n7981) );
  MUX U8018 ( .IN0(data_mem_out_wire[835]), .IN1(data_mem_out_wire[867]), 
        .SEL(N37), .F(n7982) );
  MUX U8019 ( .IN0(data_mem_out_wire[771]), .IN1(data_mem_out_wire[803]), 
        .SEL(N37), .F(n7983) );
  MUX U8020 ( .IN0(n7983), .IN1(n7982), .SEL(N38), .F(n7984) );
  MUX U8021 ( .IN0(n7984), .IN1(n7981), .SEL(N39), .F(n7985) );
  MUX U8022 ( .IN0(data_mem_out_wire[707]), .IN1(data_mem_out_wire[739]), 
        .SEL(N37), .F(n7986) );
  MUX U8023 ( .IN0(data_mem_out_wire[643]), .IN1(data_mem_out_wire[675]), 
        .SEL(N37), .F(n7987) );
  MUX U8024 ( .IN0(n7987), .IN1(n7986), .SEL(N38), .F(n7988) );
  MUX U8025 ( .IN0(data_mem_out_wire[579]), .IN1(data_mem_out_wire[611]), 
        .SEL(N37), .F(n7989) );
  MUX U8026 ( .IN0(data_mem_out_wire[515]), .IN1(data_mem_out_wire[547]), 
        .SEL(N37), .F(n7990) );
  MUX U8027 ( .IN0(n7990), .IN1(n7989), .SEL(N38), .F(n7991) );
  MUX U8028 ( .IN0(n7991), .IN1(n7988), .SEL(N39), .F(n7992) );
  MUX U8029 ( .IN0(n7992), .IN1(n7985), .SEL(N40), .F(n7993) );
  MUX U8030 ( .IN0(data_mem_out_wire[451]), .IN1(data_mem_out_wire[483]), 
        .SEL(N37), .F(n7994) );
  MUX U8031 ( .IN0(data_mem_out_wire[387]), .IN1(data_mem_out_wire[419]), 
        .SEL(N37), .F(n7995) );
  MUX U8032 ( .IN0(n7995), .IN1(n7994), .SEL(N38), .F(n7996) );
  MUX U8033 ( .IN0(data_mem_out_wire[323]), .IN1(data_mem_out_wire[355]), 
        .SEL(N37), .F(n7997) );
  MUX U8034 ( .IN0(data_mem_out_wire[259]), .IN1(data_mem_out_wire[291]), 
        .SEL(N37), .F(n7998) );
  MUX U8035 ( .IN0(n7998), .IN1(n7997), .SEL(N38), .F(n7999) );
  MUX U8036 ( .IN0(n7999), .IN1(n7996), .SEL(N39), .F(n8000) );
  MUX U8037 ( .IN0(data_mem_out_wire[195]), .IN1(data_mem_out_wire[227]), 
        .SEL(N37), .F(n8001) );
  MUX U8038 ( .IN0(data_mem_out_wire[131]), .IN1(data_mem_out_wire[163]), 
        .SEL(N37), .F(n8002) );
  MUX U8039 ( .IN0(n8002), .IN1(n8001), .SEL(N38), .F(n8003) );
  MUX U8040 ( .IN0(data_mem_out_wire[67]), .IN1(data_mem_out_wire[99]), .SEL(
        N37), .F(n8004) );
  MUX U8041 ( .IN0(data_mem_out_wire[3]), .IN1(data_mem_out_wire[35]), .SEL(
        N37), .F(n8005) );
  MUX U8042 ( .IN0(n8005), .IN1(n8004), .SEL(N38), .F(n8006) );
  MUX U8043 ( .IN0(n8006), .IN1(n8003), .SEL(N39), .F(n8007) );
  MUX U8044 ( .IN0(n8007), .IN1(n8000), .SEL(N40), .F(n8008) );
  MUX U8045 ( .IN0(n8008), .IN1(n7993), .SEL(N41), .F(n8009) );
  MUX U8046 ( .IN0(n8009), .IN1(n7978), .SEL(N42), .F(N742) );
  MUX U8047 ( .IN0(data_mem_out_wire[1988]), .IN1(data_mem_out_wire[2020]), 
        .SEL(N37), .F(n8010) );
  MUX U8048 ( .IN0(data_mem_out_wire[1924]), .IN1(data_mem_out_wire[1956]), 
        .SEL(N37), .F(n8011) );
  MUX U8049 ( .IN0(n8011), .IN1(n8010), .SEL(N38), .F(n8012) );
  MUX U8050 ( .IN0(data_mem_out_wire[1860]), .IN1(data_mem_out_wire[1892]), 
        .SEL(N37), .F(n8013) );
  MUX U8051 ( .IN0(data_mem_out_wire[1796]), .IN1(data_mem_out_wire[1828]), 
        .SEL(N37), .F(n8014) );
  MUX U8052 ( .IN0(n8014), .IN1(n8013), .SEL(N38), .F(n8015) );
  MUX U8053 ( .IN0(n8015), .IN1(n8012), .SEL(N39), .F(n8016) );
  MUX U8054 ( .IN0(data_mem_out_wire[1732]), .IN1(data_mem_out_wire[1764]), 
        .SEL(N37), .F(n8017) );
  MUX U8055 ( .IN0(data_mem_out_wire[1668]), .IN1(data_mem_out_wire[1700]), 
        .SEL(N37), .F(n8018) );
  MUX U8056 ( .IN0(n8018), .IN1(n8017), .SEL(N38), .F(n8019) );
  MUX U8057 ( .IN0(data_mem_out_wire[1604]), .IN1(data_mem_out_wire[1636]), 
        .SEL(N37), .F(n8020) );
  MUX U8058 ( .IN0(data_mem_out_wire[1540]), .IN1(data_mem_out_wire[1572]), 
        .SEL(N37), .F(n8021) );
  MUX U8059 ( .IN0(n8021), .IN1(n8020), .SEL(N38), .F(n8022) );
  MUX U8060 ( .IN0(n8022), .IN1(n8019), .SEL(N39), .F(n8023) );
  MUX U8061 ( .IN0(n8023), .IN1(n8016), .SEL(N40), .F(n8024) );
  MUX U8062 ( .IN0(data_mem_out_wire[1476]), .IN1(data_mem_out_wire[1508]), 
        .SEL(N37), .F(n8025) );
  MUX U8063 ( .IN0(data_mem_out_wire[1412]), .IN1(data_mem_out_wire[1444]), 
        .SEL(N37), .F(n8026) );
  MUX U8064 ( .IN0(n8026), .IN1(n8025), .SEL(N38), .F(n8027) );
  MUX U8065 ( .IN0(data_mem_out_wire[1348]), .IN1(data_mem_out_wire[1380]), 
        .SEL(N37), .F(n8028) );
  MUX U8066 ( .IN0(data_mem_out_wire[1284]), .IN1(data_mem_out_wire[1316]), 
        .SEL(N37), .F(n8029) );
  MUX U8067 ( .IN0(n8029), .IN1(n8028), .SEL(N38), .F(n8030) );
  MUX U8068 ( .IN0(n8030), .IN1(n8027), .SEL(N39), .F(n8031) );
  MUX U8069 ( .IN0(data_mem_out_wire[1220]), .IN1(data_mem_out_wire[1252]), 
        .SEL(N37), .F(n8032) );
  MUX U8070 ( .IN0(data_mem_out_wire[1156]), .IN1(data_mem_out_wire[1188]), 
        .SEL(N37), .F(n8033) );
  MUX U8071 ( .IN0(n8033), .IN1(n8032), .SEL(N38), .F(n8034) );
  MUX U8072 ( .IN0(data_mem_out_wire[1092]), .IN1(data_mem_out_wire[1124]), 
        .SEL(N37), .F(n8035) );
  MUX U8073 ( .IN0(data_mem_out_wire[1028]), .IN1(data_mem_out_wire[1060]), 
        .SEL(N37), .F(n8036) );
  MUX U8074 ( .IN0(n8036), .IN1(n8035), .SEL(N38), .F(n8037) );
  MUX U8075 ( .IN0(n8037), .IN1(n8034), .SEL(N39), .F(n8038) );
  MUX U8076 ( .IN0(n8038), .IN1(n8031), .SEL(N40), .F(n8039) );
  MUX U8077 ( .IN0(n8039), .IN1(n8024), .SEL(N41), .F(n8040) );
  MUX U8078 ( .IN0(data_mem_out_wire[964]), .IN1(data_mem_out_wire[996]), 
        .SEL(N37), .F(n8041) );
  MUX U8079 ( .IN0(data_mem_out_wire[900]), .IN1(data_mem_out_wire[932]), 
        .SEL(N37), .F(n8042) );
  MUX U8080 ( .IN0(n8042), .IN1(n8041), .SEL(N38), .F(n8043) );
  MUX U8081 ( .IN0(data_mem_out_wire[836]), .IN1(data_mem_out_wire[868]), 
        .SEL(N37), .F(n8044) );
  MUX U8082 ( .IN0(data_mem_out_wire[772]), .IN1(data_mem_out_wire[804]), 
        .SEL(N37), .F(n8045) );
  MUX U8083 ( .IN0(n8045), .IN1(n8044), .SEL(N38), .F(n8046) );
  MUX U8084 ( .IN0(n8046), .IN1(n8043), .SEL(N39), .F(n8047) );
  MUX U8085 ( .IN0(data_mem_out_wire[708]), .IN1(data_mem_out_wire[740]), 
        .SEL(N37), .F(n8048) );
  MUX U8086 ( .IN0(data_mem_out_wire[644]), .IN1(data_mem_out_wire[676]), 
        .SEL(N37), .F(n8049) );
  MUX U8087 ( .IN0(n8049), .IN1(n8048), .SEL(N38), .F(n8050) );
  MUX U8088 ( .IN0(data_mem_out_wire[580]), .IN1(data_mem_out_wire[612]), 
        .SEL(N37), .F(n8051) );
  MUX U8089 ( .IN0(data_mem_out_wire[516]), .IN1(data_mem_out_wire[548]), 
        .SEL(N37), .F(n8052) );
  MUX U8090 ( .IN0(n8052), .IN1(n8051), .SEL(N38), .F(n8053) );
  MUX U8091 ( .IN0(n8053), .IN1(n8050), .SEL(N39), .F(n8054) );
  MUX U8092 ( .IN0(n8054), .IN1(n8047), .SEL(N40), .F(n8055) );
  MUX U8093 ( .IN0(data_mem_out_wire[452]), .IN1(data_mem_out_wire[484]), 
        .SEL(N37), .F(n8056) );
  MUX U8094 ( .IN0(data_mem_out_wire[388]), .IN1(data_mem_out_wire[420]), 
        .SEL(N37), .F(n8057) );
  MUX U8095 ( .IN0(n8057), .IN1(n8056), .SEL(N38), .F(n8058) );
  MUX U8096 ( .IN0(data_mem_out_wire[324]), .IN1(data_mem_out_wire[356]), 
        .SEL(N37), .F(n8059) );
  MUX U8097 ( .IN0(data_mem_out_wire[260]), .IN1(data_mem_out_wire[292]), 
        .SEL(N37), .F(n8060) );
  MUX U8098 ( .IN0(n8060), .IN1(n8059), .SEL(N38), .F(n8061) );
  MUX U8099 ( .IN0(n8061), .IN1(n8058), .SEL(N39), .F(n8062) );
  MUX U8100 ( .IN0(data_mem_out_wire[196]), .IN1(data_mem_out_wire[228]), 
        .SEL(N37), .F(n8063) );
  MUX U8101 ( .IN0(data_mem_out_wire[132]), .IN1(data_mem_out_wire[164]), 
        .SEL(N37), .F(n8064) );
  MUX U8102 ( .IN0(n8064), .IN1(n8063), .SEL(N38), .F(n8065) );
  MUX U8103 ( .IN0(data_mem_out_wire[68]), .IN1(data_mem_out_wire[100]), .SEL(
        N37), .F(n8066) );
  MUX U8104 ( .IN0(data_mem_out_wire[4]), .IN1(data_mem_out_wire[36]), .SEL(
        N37), .F(n8067) );
  MUX U8105 ( .IN0(n8067), .IN1(n8066), .SEL(N38), .F(n8068) );
  MUX U8106 ( .IN0(n8068), .IN1(n8065), .SEL(N39), .F(n8069) );
  MUX U8107 ( .IN0(n8069), .IN1(n8062), .SEL(N40), .F(n8070) );
  MUX U8108 ( .IN0(n8070), .IN1(n8055), .SEL(N41), .F(n8071) );
  MUX U8109 ( .IN0(n8071), .IN1(n8040), .SEL(N42), .F(N741) );
  MUX U8110 ( .IN0(data_mem_out_wire[1989]), .IN1(data_mem_out_wire[2021]), 
        .SEL(N37), .F(n8072) );
  MUX U8111 ( .IN0(data_mem_out_wire[1925]), .IN1(data_mem_out_wire[1957]), 
        .SEL(N37), .F(n8073) );
  MUX U8112 ( .IN0(n8073), .IN1(n8072), .SEL(N38), .F(n8074) );
  MUX U8113 ( .IN0(data_mem_out_wire[1861]), .IN1(data_mem_out_wire[1893]), 
        .SEL(N37), .F(n8075) );
  MUX U8114 ( .IN0(data_mem_out_wire[1797]), .IN1(data_mem_out_wire[1829]), 
        .SEL(N37), .F(n8076) );
  MUX U8115 ( .IN0(n8076), .IN1(n8075), .SEL(N38), .F(n8077) );
  MUX U8116 ( .IN0(n8077), .IN1(n8074), .SEL(N39), .F(n8078) );
  MUX U8117 ( .IN0(data_mem_out_wire[1733]), .IN1(data_mem_out_wire[1765]), 
        .SEL(N37), .F(n8079) );
  MUX U8118 ( .IN0(data_mem_out_wire[1669]), .IN1(data_mem_out_wire[1701]), 
        .SEL(N37), .F(n8080) );
  MUX U8119 ( .IN0(n8080), .IN1(n8079), .SEL(N38), .F(n8081) );
  MUX U8120 ( .IN0(data_mem_out_wire[1605]), .IN1(data_mem_out_wire[1637]), 
        .SEL(N37), .F(n8082) );
  MUX U8121 ( .IN0(data_mem_out_wire[1541]), .IN1(data_mem_out_wire[1573]), 
        .SEL(N37), .F(n8083) );
  MUX U8122 ( .IN0(n8083), .IN1(n8082), .SEL(N38), .F(n8084) );
  MUX U8123 ( .IN0(n8084), .IN1(n8081), .SEL(N39), .F(n8085) );
  MUX U8124 ( .IN0(n8085), .IN1(n8078), .SEL(N40), .F(n8086) );
  MUX U8125 ( .IN0(data_mem_out_wire[1477]), .IN1(data_mem_out_wire[1509]), 
        .SEL(N37), .F(n8087) );
  MUX U8126 ( .IN0(data_mem_out_wire[1413]), .IN1(data_mem_out_wire[1445]), 
        .SEL(N37), .F(n8088) );
  MUX U8127 ( .IN0(n8088), .IN1(n8087), .SEL(N38), .F(n8089) );
  MUX U8128 ( .IN0(data_mem_out_wire[1349]), .IN1(data_mem_out_wire[1381]), 
        .SEL(N37), .F(n8090) );
  MUX U8129 ( .IN0(data_mem_out_wire[1285]), .IN1(data_mem_out_wire[1317]), 
        .SEL(N37), .F(n8091) );
  MUX U8130 ( .IN0(n8091), .IN1(n8090), .SEL(N38), .F(n8092) );
  MUX U8131 ( .IN0(n8092), .IN1(n8089), .SEL(N39), .F(n8093) );
  MUX U8132 ( .IN0(data_mem_out_wire[1221]), .IN1(data_mem_out_wire[1253]), 
        .SEL(N37), .F(n8094) );
  MUX U8133 ( .IN0(data_mem_out_wire[1157]), .IN1(data_mem_out_wire[1189]), 
        .SEL(N37), .F(n8095) );
  MUX U8134 ( .IN0(n8095), .IN1(n8094), .SEL(N38), .F(n8096) );
  MUX U8135 ( .IN0(data_mem_out_wire[1093]), .IN1(data_mem_out_wire[1125]), 
        .SEL(N37), .F(n8097) );
  MUX U8136 ( .IN0(data_mem_out_wire[1029]), .IN1(data_mem_out_wire[1061]), 
        .SEL(N37), .F(n8098) );
  MUX U8137 ( .IN0(n8098), .IN1(n8097), .SEL(N38), .F(n8099) );
  MUX U8138 ( .IN0(n8099), .IN1(n8096), .SEL(N39), .F(n8100) );
  MUX U8139 ( .IN0(n8100), .IN1(n8093), .SEL(N40), .F(n8101) );
  MUX U8140 ( .IN0(n8101), .IN1(n8086), .SEL(N41), .F(n8102) );
  MUX U8141 ( .IN0(data_mem_out_wire[965]), .IN1(data_mem_out_wire[997]), 
        .SEL(N37), .F(n8103) );
  MUX U8142 ( .IN0(data_mem_out_wire[901]), .IN1(data_mem_out_wire[933]), 
        .SEL(N37), .F(n8104) );
  MUX U8143 ( .IN0(n8104), .IN1(n8103), .SEL(N38), .F(n8105) );
  MUX U8144 ( .IN0(data_mem_out_wire[837]), .IN1(data_mem_out_wire[869]), 
        .SEL(N37), .F(n8106) );
  MUX U8145 ( .IN0(data_mem_out_wire[773]), .IN1(data_mem_out_wire[805]), 
        .SEL(N37), .F(n8107) );
  MUX U8146 ( .IN0(n8107), .IN1(n8106), .SEL(N38), .F(n8108) );
  MUX U8147 ( .IN0(n8108), .IN1(n8105), .SEL(N39), .F(n8109) );
  MUX U8148 ( .IN0(data_mem_out_wire[709]), .IN1(data_mem_out_wire[741]), 
        .SEL(N37), .F(n8110) );
  MUX U8149 ( .IN0(data_mem_out_wire[645]), .IN1(data_mem_out_wire[677]), 
        .SEL(N37), .F(n8111) );
  MUX U8150 ( .IN0(n8111), .IN1(n8110), .SEL(N38), .F(n8112) );
  MUX U8151 ( .IN0(data_mem_out_wire[581]), .IN1(data_mem_out_wire[613]), 
        .SEL(N37), .F(n8113) );
  MUX U8152 ( .IN0(data_mem_out_wire[517]), .IN1(data_mem_out_wire[549]), 
        .SEL(N37), .F(n8114) );
  MUX U8153 ( .IN0(n8114), .IN1(n8113), .SEL(N38), .F(n8115) );
  MUX U8154 ( .IN0(n8115), .IN1(n8112), .SEL(N39), .F(n8116) );
  MUX U8155 ( .IN0(n8116), .IN1(n8109), .SEL(N40), .F(n8117) );
  MUX U8156 ( .IN0(data_mem_out_wire[453]), .IN1(data_mem_out_wire[485]), 
        .SEL(N37), .F(n8118) );
  MUX U8157 ( .IN0(data_mem_out_wire[389]), .IN1(data_mem_out_wire[421]), 
        .SEL(N37), .F(n8119) );
  MUX U8158 ( .IN0(n8119), .IN1(n8118), .SEL(N38), .F(n8120) );
  MUX U8159 ( .IN0(data_mem_out_wire[325]), .IN1(data_mem_out_wire[357]), 
        .SEL(N37), .F(n8121) );
  MUX U8160 ( .IN0(data_mem_out_wire[261]), .IN1(data_mem_out_wire[293]), 
        .SEL(N37), .F(n8122) );
  MUX U8161 ( .IN0(n8122), .IN1(n8121), .SEL(N38), .F(n8123) );
  MUX U8162 ( .IN0(n8123), .IN1(n8120), .SEL(N39), .F(n8124) );
  MUX U8163 ( .IN0(data_mem_out_wire[197]), .IN1(data_mem_out_wire[229]), 
        .SEL(N37), .F(n8125) );
  MUX U8164 ( .IN0(data_mem_out_wire[133]), .IN1(data_mem_out_wire[165]), 
        .SEL(N37), .F(n8126) );
  MUX U8165 ( .IN0(n8126), .IN1(n8125), .SEL(N38), .F(n8127) );
  MUX U8166 ( .IN0(data_mem_out_wire[69]), .IN1(data_mem_out_wire[101]), .SEL(
        N37), .F(n8128) );
  MUX U8167 ( .IN0(data_mem_out_wire[5]), .IN1(data_mem_out_wire[37]), .SEL(
        N37), .F(n8129) );
  MUX U8168 ( .IN0(n8129), .IN1(n8128), .SEL(N38), .F(n8130) );
  MUX U8169 ( .IN0(n8130), .IN1(n8127), .SEL(N39), .F(n8131) );
  MUX U8170 ( .IN0(n8131), .IN1(n8124), .SEL(N40), .F(n8132) );
  MUX U8171 ( .IN0(n8132), .IN1(n8117), .SEL(N41), .F(n8133) );
  MUX U8172 ( .IN0(n8133), .IN1(n8102), .SEL(N42), .F(N740) );
  MUX U8173 ( .IN0(data_mem_out_wire[1990]), .IN1(data_mem_out_wire[2022]), 
        .SEL(N37), .F(n8134) );
  MUX U8174 ( .IN0(data_mem_out_wire[1926]), .IN1(data_mem_out_wire[1958]), 
        .SEL(N37), .F(n8135) );
  MUX U8175 ( .IN0(n8135), .IN1(n8134), .SEL(N38), .F(n8136) );
  MUX U8176 ( .IN0(data_mem_out_wire[1862]), .IN1(data_mem_out_wire[1894]), 
        .SEL(N37), .F(n8137) );
  MUX U8177 ( .IN0(data_mem_out_wire[1798]), .IN1(data_mem_out_wire[1830]), 
        .SEL(N37), .F(n8138) );
  MUX U8178 ( .IN0(n8138), .IN1(n8137), .SEL(N38), .F(n8139) );
  MUX U8179 ( .IN0(n8139), .IN1(n8136), .SEL(N39), .F(n8140) );
  MUX U8180 ( .IN0(data_mem_out_wire[1734]), .IN1(data_mem_out_wire[1766]), 
        .SEL(N37), .F(n8141) );
  MUX U8181 ( .IN0(data_mem_out_wire[1670]), .IN1(data_mem_out_wire[1702]), 
        .SEL(N37), .F(n8142) );
  MUX U8182 ( .IN0(n8142), .IN1(n8141), .SEL(N38), .F(n8143) );
  MUX U8183 ( .IN0(data_mem_out_wire[1606]), .IN1(data_mem_out_wire[1638]), 
        .SEL(N37), .F(n8144) );
  MUX U8184 ( .IN0(data_mem_out_wire[1542]), .IN1(data_mem_out_wire[1574]), 
        .SEL(N37), .F(n8145) );
  MUX U8185 ( .IN0(n8145), .IN1(n8144), .SEL(N38), .F(n8146) );
  MUX U8186 ( .IN0(n8146), .IN1(n8143), .SEL(N39), .F(n8147) );
  MUX U8187 ( .IN0(n8147), .IN1(n8140), .SEL(N40), .F(n8148) );
  MUX U8188 ( .IN0(data_mem_out_wire[1478]), .IN1(data_mem_out_wire[1510]), 
        .SEL(N37), .F(n8149) );
  MUX U8189 ( .IN0(data_mem_out_wire[1414]), .IN1(data_mem_out_wire[1446]), 
        .SEL(N37), .F(n8150) );
  MUX U8190 ( .IN0(n8150), .IN1(n8149), .SEL(N38), .F(n8151) );
  MUX U8191 ( .IN0(data_mem_out_wire[1350]), .IN1(data_mem_out_wire[1382]), 
        .SEL(N37), .F(n8152) );
  MUX U8192 ( .IN0(data_mem_out_wire[1286]), .IN1(data_mem_out_wire[1318]), 
        .SEL(N37), .F(n8153) );
  MUX U8193 ( .IN0(n8153), .IN1(n8152), .SEL(N38), .F(n8154) );
  MUX U8194 ( .IN0(n8154), .IN1(n8151), .SEL(N39), .F(n8155) );
  MUX U8195 ( .IN0(data_mem_out_wire[1222]), .IN1(data_mem_out_wire[1254]), 
        .SEL(N37), .F(n8156) );
  MUX U8196 ( .IN0(data_mem_out_wire[1158]), .IN1(data_mem_out_wire[1190]), 
        .SEL(N37), .F(n8157) );
  MUX U8197 ( .IN0(n8157), .IN1(n8156), .SEL(N38), .F(n8158) );
  MUX U8198 ( .IN0(data_mem_out_wire[1094]), .IN1(data_mem_out_wire[1126]), 
        .SEL(N37), .F(n8159) );
  MUX U8199 ( .IN0(data_mem_out_wire[1030]), .IN1(data_mem_out_wire[1062]), 
        .SEL(N37), .F(n8160) );
  MUX U8200 ( .IN0(n8160), .IN1(n8159), .SEL(N38), .F(n8161) );
  MUX U8201 ( .IN0(n8161), .IN1(n8158), .SEL(N39), .F(n8162) );
  MUX U8202 ( .IN0(n8162), .IN1(n8155), .SEL(N40), .F(n8163) );
  MUX U8203 ( .IN0(n8163), .IN1(n8148), .SEL(N41), .F(n8164) );
  MUX U8204 ( .IN0(data_mem_out_wire[966]), .IN1(data_mem_out_wire[998]), 
        .SEL(N37), .F(n8165) );
  MUX U8205 ( .IN0(data_mem_out_wire[902]), .IN1(data_mem_out_wire[934]), 
        .SEL(N37), .F(n8166) );
  MUX U8206 ( .IN0(n8166), .IN1(n8165), .SEL(N38), .F(n8167) );
  MUX U8207 ( .IN0(data_mem_out_wire[838]), .IN1(data_mem_out_wire[870]), 
        .SEL(N37), .F(n8168) );
  MUX U8208 ( .IN0(data_mem_out_wire[774]), .IN1(data_mem_out_wire[806]), 
        .SEL(N37), .F(n8169) );
  MUX U8209 ( .IN0(n8169), .IN1(n8168), .SEL(N38), .F(n8170) );
  MUX U8210 ( .IN0(n8170), .IN1(n8167), .SEL(N39), .F(n8171) );
  MUX U8211 ( .IN0(data_mem_out_wire[710]), .IN1(data_mem_out_wire[742]), 
        .SEL(N37), .F(n8172) );
  MUX U8212 ( .IN0(data_mem_out_wire[646]), .IN1(data_mem_out_wire[678]), 
        .SEL(N37), .F(n8173) );
  MUX U8213 ( .IN0(n8173), .IN1(n8172), .SEL(N38), .F(n8174) );
  MUX U8214 ( .IN0(data_mem_out_wire[582]), .IN1(data_mem_out_wire[614]), 
        .SEL(N37), .F(n8175) );
  MUX U8215 ( .IN0(data_mem_out_wire[518]), .IN1(data_mem_out_wire[550]), 
        .SEL(N37), .F(n8176) );
  MUX U8216 ( .IN0(n8176), .IN1(n8175), .SEL(N38), .F(n8177) );
  MUX U8217 ( .IN0(n8177), .IN1(n8174), .SEL(N39), .F(n8178) );
  MUX U8218 ( .IN0(n8178), .IN1(n8171), .SEL(N40), .F(n8179) );
  MUX U8219 ( .IN0(data_mem_out_wire[454]), .IN1(data_mem_out_wire[486]), 
        .SEL(N37), .F(n8180) );
  MUX U8220 ( .IN0(data_mem_out_wire[390]), .IN1(data_mem_out_wire[422]), 
        .SEL(N37), .F(n8181) );
  MUX U8221 ( .IN0(n8181), .IN1(n8180), .SEL(N38), .F(n8182) );
  MUX U8222 ( .IN0(data_mem_out_wire[326]), .IN1(data_mem_out_wire[358]), 
        .SEL(N37), .F(n8183) );
  MUX U8223 ( .IN0(data_mem_out_wire[262]), .IN1(data_mem_out_wire[294]), 
        .SEL(N37), .F(n8184) );
  MUX U8224 ( .IN0(n8184), .IN1(n8183), .SEL(N38), .F(n8185) );
  MUX U8225 ( .IN0(n8185), .IN1(n8182), .SEL(N39), .F(n8186) );
  MUX U8226 ( .IN0(data_mem_out_wire[198]), .IN1(data_mem_out_wire[230]), 
        .SEL(N37), .F(n8187) );
  MUX U8227 ( .IN0(data_mem_out_wire[134]), .IN1(data_mem_out_wire[166]), 
        .SEL(N37), .F(n8188) );
  MUX U8228 ( .IN0(n8188), .IN1(n8187), .SEL(N38), .F(n8189) );
  MUX U8229 ( .IN0(data_mem_out_wire[70]), .IN1(data_mem_out_wire[102]), .SEL(
        N37), .F(n8190) );
  MUX U8230 ( .IN0(data_mem_out_wire[6]), .IN1(data_mem_out_wire[38]), .SEL(
        N37), .F(n8191) );
  MUX U8231 ( .IN0(n8191), .IN1(n8190), .SEL(N38), .F(n8192) );
  MUX U8232 ( .IN0(n8192), .IN1(n8189), .SEL(N39), .F(n8193) );
  MUX U8233 ( .IN0(n8193), .IN1(n8186), .SEL(N40), .F(n8194) );
  MUX U8234 ( .IN0(n8194), .IN1(n8179), .SEL(N41), .F(n8195) );
  MUX U8235 ( .IN0(n8195), .IN1(n8164), .SEL(N42), .F(N739) );
  MUX U8236 ( .IN0(data_mem_out_wire[1991]), .IN1(data_mem_out_wire[2023]), 
        .SEL(N37), .F(n8196) );
  MUX U8237 ( .IN0(data_mem_out_wire[1927]), .IN1(data_mem_out_wire[1959]), 
        .SEL(N37), .F(n8197) );
  MUX U8238 ( .IN0(n8197), .IN1(n8196), .SEL(N38), .F(n8198) );
  MUX U8239 ( .IN0(data_mem_out_wire[1863]), .IN1(data_mem_out_wire[1895]), 
        .SEL(N37), .F(n8199) );
  MUX U8240 ( .IN0(data_mem_out_wire[1799]), .IN1(data_mem_out_wire[1831]), 
        .SEL(N37), .F(n8200) );
  MUX U8241 ( .IN0(n8200), .IN1(n8199), .SEL(N38), .F(n8201) );
  MUX U8242 ( .IN0(n8201), .IN1(n8198), .SEL(N39), .F(n8202) );
  MUX U8243 ( .IN0(data_mem_out_wire[1735]), .IN1(data_mem_out_wire[1767]), 
        .SEL(N37), .F(n8203) );
  MUX U8244 ( .IN0(data_mem_out_wire[1671]), .IN1(data_mem_out_wire[1703]), 
        .SEL(N37), .F(n8204) );
  MUX U8245 ( .IN0(n8204), .IN1(n8203), .SEL(N38), .F(n8205) );
  MUX U8246 ( .IN0(data_mem_out_wire[1607]), .IN1(data_mem_out_wire[1639]), 
        .SEL(N37), .F(n8206) );
  MUX U8247 ( .IN0(data_mem_out_wire[1543]), .IN1(data_mem_out_wire[1575]), 
        .SEL(N37), .F(n8207) );
  MUX U8248 ( .IN0(n8207), .IN1(n8206), .SEL(N38), .F(n8208) );
  MUX U8249 ( .IN0(n8208), .IN1(n8205), .SEL(N39), .F(n8209) );
  MUX U8250 ( .IN0(n8209), .IN1(n8202), .SEL(N40), .F(n8210) );
  MUX U8251 ( .IN0(data_mem_out_wire[1479]), .IN1(data_mem_out_wire[1511]), 
        .SEL(N37), .F(n8211) );
  MUX U8252 ( .IN0(data_mem_out_wire[1415]), .IN1(data_mem_out_wire[1447]), 
        .SEL(N37), .F(n8212) );
  MUX U8253 ( .IN0(n8212), .IN1(n8211), .SEL(N38), .F(n8213) );
  MUX U8254 ( .IN0(data_mem_out_wire[1351]), .IN1(data_mem_out_wire[1383]), 
        .SEL(N37), .F(n8214) );
  MUX U8255 ( .IN0(data_mem_out_wire[1287]), .IN1(data_mem_out_wire[1319]), 
        .SEL(N37), .F(n8215) );
  MUX U8256 ( .IN0(n8215), .IN1(n8214), .SEL(N38), .F(n8216) );
  MUX U8257 ( .IN0(n8216), .IN1(n8213), .SEL(N39), .F(n8217) );
  MUX U8258 ( .IN0(data_mem_out_wire[1223]), .IN1(data_mem_out_wire[1255]), 
        .SEL(N37), .F(n8218) );
  MUX U8259 ( .IN0(data_mem_out_wire[1159]), .IN1(data_mem_out_wire[1191]), 
        .SEL(N37), .F(n8219) );
  MUX U8260 ( .IN0(n8219), .IN1(n8218), .SEL(N38), .F(n8220) );
  MUX U8261 ( .IN0(data_mem_out_wire[1095]), .IN1(data_mem_out_wire[1127]), 
        .SEL(N37), .F(n8221) );
  MUX U8262 ( .IN0(data_mem_out_wire[1031]), .IN1(data_mem_out_wire[1063]), 
        .SEL(N37), .F(n8222) );
  MUX U8263 ( .IN0(n8222), .IN1(n8221), .SEL(N38), .F(n8223) );
  MUX U8264 ( .IN0(n8223), .IN1(n8220), .SEL(N39), .F(n8224) );
  MUX U8265 ( .IN0(n8224), .IN1(n8217), .SEL(N40), .F(n8225) );
  MUX U8266 ( .IN0(n8225), .IN1(n8210), .SEL(N41), .F(n8226) );
  MUX U8267 ( .IN0(data_mem_out_wire[967]), .IN1(data_mem_out_wire[999]), 
        .SEL(N37), .F(n8227) );
  MUX U8268 ( .IN0(data_mem_out_wire[903]), .IN1(data_mem_out_wire[935]), 
        .SEL(N37), .F(n8228) );
  MUX U8269 ( .IN0(n8228), .IN1(n8227), .SEL(N38), .F(n8229) );
  MUX U8270 ( .IN0(data_mem_out_wire[839]), .IN1(data_mem_out_wire[871]), 
        .SEL(N37), .F(n8230) );
  MUX U8271 ( .IN0(data_mem_out_wire[775]), .IN1(data_mem_out_wire[807]), 
        .SEL(N37), .F(n8231) );
  MUX U8272 ( .IN0(n8231), .IN1(n8230), .SEL(N38), .F(n8232) );
  MUX U8273 ( .IN0(n8232), .IN1(n8229), .SEL(N39), .F(n8233) );
  MUX U8274 ( .IN0(data_mem_out_wire[711]), .IN1(data_mem_out_wire[743]), 
        .SEL(N37), .F(n8234) );
  MUX U8275 ( .IN0(data_mem_out_wire[647]), .IN1(data_mem_out_wire[679]), 
        .SEL(N37), .F(n8235) );
  MUX U8276 ( .IN0(n8235), .IN1(n8234), .SEL(N38), .F(n8236) );
  MUX U8277 ( .IN0(data_mem_out_wire[583]), .IN1(data_mem_out_wire[615]), 
        .SEL(N37), .F(n8237) );
  MUX U8278 ( .IN0(data_mem_out_wire[519]), .IN1(data_mem_out_wire[551]), 
        .SEL(N37), .F(n8238) );
  MUX U8279 ( .IN0(n8238), .IN1(n8237), .SEL(N38), .F(n8239) );
  MUX U8280 ( .IN0(n8239), .IN1(n8236), .SEL(N39), .F(n8240) );
  MUX U8281 ( .IN0(n8240), .IN1(n8233), .SEL(N40), .F(n8241) );
  MUX U8282 ( .IN0(data_mem_out_wire[455]), .IN1(data_mem_out_wire[487]), 
        .SEL(N37), .F(n8242) );
  MUX U8283 ( .IN0(data_mem_out_wire[391]), .IN1(data_mem_out_wire[423]), 
        .SEL(N37), .F(n8243) );
  MUX U8284 ( .IN0(n8243), .IN1(n8242), .SEL(N38), .F(n8244) );
  MUX U8285 ( .IN0(data_mem_out_wire[327]), .IN1(data_mem_out_wire[359]), 
        .SEL(N37), .F(n8245) );
  MUX U8286 ( .IN0(data_mem_out_wire[263]), .IN1(data_mem_out_wire[295]), 
        .SEL(N37), .F(n8246) );
  MUX U8287 ( .IN0(n8246), .IN1(n8245), .SEL(N38), .F(n8247) );
  MUX U8288 ( .IN0(n8247), .IN1(n8244), .SEL(N39), .F(n8248) );
  MUX U8289 ( .IN0(data_mem_out_wire[199]), .IN1(data_mem_out_wire[231]), 
        .SEL(N37), .F(n8249) );
  MUX U8290 ( .IN0(data_mem_out_wire[135]), .IN1(data_mem_out_wire[167]), 
        .SEL(N37), .F(n8250) );
  MUX U8291 ( .IN0(n8250), .IN1(n8249), .SEL(N38), .F(n8251) );
  MUX U8292 ( .IN0(data_mem_out_wire[71]), .IN1(data_mem_out_wire[103]), .SEL(
        N37), .F(n8252) );
  MUX U8293 ( .IN0(data_mem_out_wire[7]), .IN1(data_mem_out_wire[39]), .SEL(
        N37), .F(n8253) );
  MUX U8294 ( .IN0(n8253), .IN1(n8252), .SEL(N38), .F(n8254) );
  MUX U8295 ( .IN0(n8254), .IN1(n8251), .SEL(N39), .F(n8255) );
  MUX U8296 ( .IN0(n8255), .IN1(n8248), .SEL(N40), .F(n8256) );
  MUX U8297 ( .IN0(n8256), .IN1(n8241), .SEL(N41), .F(n8257) );
  MUX U8298 ( .IN0(n8257), .IN1(n8226), .SEL(N42), .F(N738) );
  MUX U8299 ( .IN0(data_mem_out_wire[1992]), .IN1(data_mem_out_wire[2024]), 
        .SEL(N37), .F(n8258) );
  MUX U8300 ( .IN0(data_mem_out_wire[1928]), .IN1(data_mem_out_wire[1960]), 
        .SEL(N37), .F(n8259) );
  MUX U8301 ( .IN0(n8259), .IN1(n8258), .SEL(N38), .F(n8260) );
  MUX U8302 ( .IN0(data_mem_out_wire[1864]), .IN1(data_mem_out_wire[1896]), 
        .SEL(N37), .F(n8261) );
  MUX U8303 ( .IN0(data_mem_out_wire[1800]), .IN1(data_mem_out_wire[1832]), 
        .SEL(N37), .F(n8262) );
  MUX U8304 ( .IN0(n8262), .IN1(n8261), .SEL(N38), .F(n8263) );
  MUX U8305 ( .IN0(n8263), .IN1(n8260), .SEL(N39), .F(n8264) );
  MUX U8306 ( .IN0(data_mem_out_wire[1736]), .IN1(data_mem_out_wire[1768]), 
        .SEL(N37), .F(n8265) );
  MUX U8307 ( .IN0(data_mem_out_wire[1672]), .IN1(data_mem_out_wire[1704]), 
        .SEL(N37), .F(n8266) );
  MUX U8308 ( .IN0(n8266), .IN1(n8265), .SEL(N38), .F(n8267) );
  MUX U8309 ( .IN0(data_mem_out_wire[1608]), .IN1(data_mem_out_wire[1640]), 
        .SEL(N37), .F(n8268) );
  MUX U8310 ( .IN0(data_mem_out_wire[1544]), .IN1(data_mem_out_wire[1576]), 
        .SEL(N37), .F(n8269) );
  MUX U8311 ( .IN0(n8269), .IN1(n8268), .SEL(N38), .F(n8270) );
  MUX U8312 ( .IN0(n8270), .IN1(n8267), .SEL(N39), .F(n8271) );
  MUX U8313 ( .IN0(n8271), .IN1(n8264), .SEL(N40), .F(n8272) );
  MUX U8314 ( .IN0(data_mem_out_wire[1480]), .IN1(data_mem_out_wire[1512]), 
        .SEL(N37), .F(n8273) );
  MUX U8315 ( .IN0(data_mem_out_wire[1416]), .IN1(data_mem_out_wire[1448]), 
        .SEL(N37), .F(n8274) );
  MUX U8316 ( .IN0(n8274), .IN1(n8273), .SEL(N38), .F(n8275) );
  MUX U8317 ( .IN0(data_mem_out_wire[1352]), .IN1(data_mem_out_wire[1384]), 
        .SEL(N37), .F(n8276) );
  MUX U8318 ( .IN0(data_mem_out_wire[1288]), .IN1(data_mem_out_wire[1320]), 
        .SEL(N37), .F(n8277) );
  MUX U8319 ( .IN0(n8277), .IN1(n8276), .SEL(N38), .F(n8278) );
  MUX U8320 ( .IN0(n8278), .IN1(n8275), .SEL(N39), .F(n8279) );
  MUX U8321 ( .IN0(data_mem_out_wire[1224]), .IN1(data_mem_out_wire[1256]), 
        .SEL(N37), .F(n8280) );
  MUX U8322 ( .IN0(data_mem_out_wire[1160]), .IN1(data_mem_out_wire[1192]), 
        .SEL(N37), .F(n8281) );
  MUX U8323 ( .IN0(n8281), .IN1(n8280), .SEL(N38), .F(n8282) );
  MUX U8324 ( .IN0(data_mem_out_wire[1096]), .IN1(data_mem_out_wire[1128]), 
        .SEL(N37), .F(n8283) );
  MUX U8325 ( .IN0(data_mem_out_wire[1032]), .IN1(data_mem_out_wire[1064]), 
        .SEL(N37), .F(n8284) );
  MUX U8326 ( .IN0(n8284), .IN1(n8283), .SEL(N38), .F(n8285) );
  MUX U8327 ( .IN0(n8285), .IN1(n8282), .SEL(N39), .F(n8286) );
  MUX U8328 ( .IN0(n8286), .IN1(n8279), .SEL(N40), .F(n8287) );
  MUX U8329 ( .IN0(n8287), .IN1(n8272), .SEL(N41), .F(n8288) );
  MUX U8330 ( .IN0(data_mem_out_wire[968]), .IN1(data_mem_out_wire[1000]), 
        .SEL(N37), .F(n8289) );
  MUX U8331 ( .IN0(data_mem_out_wire[904]), .IN1(data_mem_out_wire[936]), 
        .SEL(N37), .F(n8290) );
  MUX U8332 ( .IN0(n8290), .IN1(n8289), .SEL(N38), .F(n8291) );
  MUX U8333 ( .IN0(data_mem_out_wire[840]), .IN1(data_mem_out_wire[872]), 
        .SEL(N37), .F(n8292) );
  MUX U8334 ( .IN0(data_mem_out_wire[776]), .IN1(data_mem_out_wire[808]), 
        .SEL(N37), .F(n8293) );
  MUX U8335 ( .IN0(n8293), .IN1(n8292), .SEL(N38), .F(n8294) );
  MUX U8336 ( .IN0(n8294), .IN1(n8291), .SEL(N39), .F(n8295) );
  MUX U8337 ( .IN0(data_mem_out_wire[712]), .IN1(data_mem_out_wire[744]), 
        .SEL(N37), .F(n8296) );
  MUX U8338 ( .IN0(data_mem_out_wire[648]), .IN1(data_mem_out_wire[680]), 
        .SEL(N37), .F(n8297) );
  MUX U8339 ( .IN0(n8297), .IN1(n8296), .SEL(N38), .F(n8298) );
  MUX U8340 ( .IN0(data_mem_out_wire[584]), .IN1(data_mem_out_wire[616]), 
        .SEL(N37), .F(n8299) );
  MUX U8341 ( .IN0(data_mem_out_wire[520]), .IN1(data_mem_out_wire[552]), 
        .SEL(N37), .F(n8300) );
  MUX U8342 ( .IN0(n8300), .IN1(n8299), .SEL(N38), .F(n8301) );
  MUX U8343 ( .IN0(n8301), .IN1(n8298), .SEL(N39), .F(n8302) );
  MUX U8344 ( .IN0(n8302), .IN1(n8295), .SEL(N40), .F(n8303) );
  MUX U8345 ( .IN0(data_mem_out_wire[456]), .IN1(data_mem_out_wire[488]), 
        .SEL(N37), .F(n8304) );
  MUX U8346 ( .IN0(data_mem_out_wire[392]), .IN1(data_mem_out_wire[424]), 
        .SEL(N37), .F(n8305) );
  MUX U8347 ( .IN0(n8305), .IN1(n8304), .SEL(N38), .F(n8306) );
  MUX U8348 ( .IN0(data_mem_out_wire[328]), .IN1(data_mem_out_wire[360]), 
        .SEL(N37), .F(n8307) );
  MUX U8349 ( .IN0(data_mem_out_wire[264]), .IN1(data_mem_out_wire[296]), 
        .SEL(N37), .F(n8308) );
  MUX U8350 ( .IN0(n8308), .IN1(n8307), .SEL(N38), .F(n8309) );
  MUX U8351 ( .IN0(n8309), .IN1(n8306), .SEL(N39), .F(n8310) );
  MUX U8352 ( .IN0(data_mem_out_wire[200]), .IN1(data_mem_out_wire[232]), 
        .SEL(N37), .F(n8311) );
  MUX U8353 ( .IN0(data_mem_out_wire[136]), .IN1(data_mem_out_wire[168]), 
        .SEL(N37), .F(n8312) );
  MUX U8354 ( .IN0(n8312), .IN1(n8311), .SEL(N38), .F(n8313) );
  MUX U8355 ( .IN0(data_mem_out_wire[72]), .IN1(data_mem_out_wire[104]), .SEL(
        N37), .F(n8314) );
  MUX U8356 ( .IN0(data_mem_out_wire[8]), .IN1(data_mem_out_wire[40]), .SEL(
        N37), .F(n8315) );
  MUX U8357 ( .IN0(n8315), .IN1(n8314), .SEL(N38), .F(n8316) );
  MUX U8358 ( .IN0(n8316), .IN1(n8313), .SEL(N39), .F(n8317) );
  MUX U8359 ( .IN0(n8317), .IN1(n8310), .SEL(N40), .F(n8318) );
  MUX U8360 ( .IN0(n8318), .IN1(n8303), .SEL(N41), .F(n8319) );
  MUX U8361 ( .IN0(n8319), .IN1(n8288), .SEL(N42), .F(N737) );
  MUX U8362 ( .IN0(data_mem_out_wire[1993]), .IN1(data_mem_out_wire[2025]), 
        .SEL(N37), .F(n8320) );
  MUX U8363 ( .IN0(data_mem_out_wire[1929]), .IN1(data_mem_out_wire[1961]), 
        .SEL(N37), .F(n8321) );
  MUX U8364 ( .IN0(n8321), .IN1(n8320), .SEL(N38), .F(n8322) );
  MUX U8365 ( .IN0(data_mem_out_wire[1865]), .IN1(data_mem_out_wire[1897]), 
        .SEL(N37), .F(n8323) );
  MUX U8366 ( .IN0(data_mem_out_wire[1801]), .IN1(data_mem_out_wire[1833]), 
        .SEL(N37), .F(n8324) );
  MUX U8367 ( .IN0(n8324), .IN1(n8323), .SEL(N38), .F(n8325) );
  MUX U8368 ( .IN0(n8325), .IN1(n8322), .SEL(N39), .F(n8326) );
  MUX U8369 ( .IN0(data_mem_out_wire[1737]), .IN1(data_mem_out_wire[1769]), 
        .SEL(N37), .F(n8327) );
  MUX U8370 ( .IN0(data_mem_out_wire[1673]), .IN1(data_mem_out_wire[1705]), 
        .SEL(N37), .F(n8328) );
  MUX U8371 ( .IN0(n8328), .IN1(n8327), .SEL(N38), .F(n8329) );
  MUX U8372 ( .IN0(data_mem_out_wire[1609]), .IN1(data_mem_out_wire[1641]), 
        .SEL(N37), .F(n8330) );
  MUX U8373 ( .IN0(data_mem_out_wire[1545]), .IN1(data_mem_out_wire[1577]), 
        .SEL(N37), .F(n8331) );
  MUX U8374 ( .IN0(n8331), .IN1(n8330), .SEL(N38), .F(n8332) );
  MUX U8375 ( .IN0(n8332), .IN1(n8329), .SEL(N39), .F(n8333) );
  MUX U8376 ( .IN0(n8333), .IN1(n8326), .SEL(N40), .F(n8334) );
  MUX U8377 ( .IN0(data_mem_out_wire[1481]), .IN1(data_mem_out_wire[1513]), 
        .SEL(N37), .F(n8335) );
  MUX U8378 ( .IN0(data_mem_out_wire[1417]), .IN1(data_mem_out_wire[1449]), 
        .SEL(N37), .F(n8336) );
  MUX U8379 ( .IN0(n8336), .IN1(n8335), .SEL(N38), .F(n8337) );
  MUX U8380 ( .IN0(data_mem_out_wire[1353]), .IN1(data_mem_out_wire[1385]), 
        .SEL(N37), .F(n8338) );
  MUX U8381 ( .IN0(data_mem_out_wire[1289]), .IN1(data_mem_out_wire[1321]), 
        .SEL(N37), .F(n8339) );
  MUX U8382 ( .IN0(n8339), .IN1(n8338), .SEL(N38), .F(n8340) );
  MUX U8383 ( .IN0(n8340), .IN1(n8337), .SEL(N39), .F(n8341) );
  MUX U8384 ( .IN0(data_mem_out_wire[1225]), .IN1(data_mem_out_wire[1257]), 
        .SEL(N37), .F(n8342) );
  MUX U8385 ( .IN0(data_mem_out_wire[1161]), .IN1(data_mem_out_wire[1193]), 
        .SEL(N37), .F(n8343) );
  MUX U8386 ( .IN0(n8343), .IN1(n8342), .SEL(N38), .F(n8344) );
  MUX U8387 ( .IN0(data_mem_out_wire[1097]), .IN1(data_mem_out_wire[1129]), 
        .SEL(N37), .F(n8345) );
  MUX U8388 ( .IN0(data_mem_out_wire[1033]), .IN1(data_mem_out_wire[1065]), 
        .SEL(N37), .F(n8346) );
  MUX U8389 ( .IN0(n8346), .IN1(n8345), .SEL(N38), .F(n8347) );
  MUX U8390 ( .IN0(n8347), .IN1(n8344), .SEL(N39), .F(n8348) );
  MUX U8391 ( .IN0(n8348), .IN1(n8341), .SEL(N40), .F(n8349) );
  MUX U8392 ( .IN0(n8349), .IN1(n8334), .SEL(N41), .F(n8350) );
  MUX U8393 ( .IN0(data_mem_out_wire[969]), .IN1(data_mem_out_wire[1001]), 
        .SEL(N37), .F(n8351) );
  MUX U8394 ( .IN0(data_mem_out_wire[905]), .IN1(data_mem_out_wire[937]), 
        .SEL(N37), .F(n8352) );
  MUX U8395 ( .IN0(n8352), .IN1(n8351), .SEL(N38), .F(n8353) );
  MUX U8396 ( .IN0(data_mem_out_wire[841]), .IN1(data_mem_out_wire[873]), 
        .SEL(N37), .F(n8354) );
  MUX U8397 ( .IN0(data_mem_out_wire[777]), .IN1(data_mem_out_wire[809]), 
        .SEL(N37), .F(n8355) );
  MUX U8398 ( .IN0(n8355), .IN1(n8354), .SEL(N38), .F(n8356) );
  MUX U8399 ( .IN0(n8356), .IN1(n8353), .SEL(N39), .F(n8357) );
  MUX U8400 ( .IN0(data_mem_out_wire[713]), .IN1(data_mem_out_wire[745]), 
        .SEL(N37), .F(n8358) );
  MUX U8401 ( .IN0(data_mem_out_wire[649]), .IN1(data_mem_out_wire[681]), 
        .SEL(N37), .F(n8359) );
  MUX U8402 ( .IN0(n8359), .IN1(n8358), .SEL(N38), .F(n8360) );
  MUX U8403 ( .IN0(data_mem_out_wire[585]), .IN1(data_mem_out_wire[617]), 
        .SEL(N37), .F(n8361) );
  MUX U8404 ( .IN0(data_mem_out_wire[521]), .IN1(data_mem_out_wire[553]), 
        .SEL(N37), .F(n8362) );
  MUX U8405 ( .IN0(n8362), .IN1(n8361), .SEL(N38), .F(n8363) );
  MUX U8406 ( .IN0(n8363), .IN1(n8360), .SEL(N39), .F(n8364) );
  MUX U8407 ( .IN0(n8364), .IN1(n8357), .SEL(N40), .F(n8365) );
  MUX U8408 ( .IN0(data_mem_out_wire[457]), .IN1(data_mem_out_wire[489]), 
        .SEL(N37), .F(n8366) );
  MUX U8409 ( .IN0(data_mem_out_wire[393]), .IN1(data_mem_out_wire[425]), 
        .SEL(N37), .F(n8367) );
  MUX U8410 ( .IN0(n8367), .IN1(n8366), .SEL(N38), .F(n8368) );
  MUX U8411 ( .IN0(data_mem_out_wire[329]), .IN1(data_mem_out_wire[361]), 
        .SEL(N37), .F(n8369) );
  MUX U8412 ( .IN0(data_mem_out_wire[265]), .IN1(data_mem_out_wire[297]), 
        .SEL(N37), .F(n8370) );
  MUX U8413 ( .IN0(n8370), .IN1(n8369), .SEL(N38), .F(n8371) );
  MUX U8414 ( .IN0(n8371), .IN1(n8368), .SEL(N39), .F(n8372) );
  MUX U8415 ( .IN0(data_mem_out_wire[201]), .IN1(data_mem_out_wire[233]), 
        .SEL(N37), .F(n8373) );
  MUX U8416 ( .IN0(data_mem_out_wire[137]), .IN1(data_mem_out_wire[169]), 
        .SEL(N37), .F(n8374) );
  MUX U8417 ( .IN0(n8374), .IN1(n8373), .SEL(N38), .F(n8375) );
  MUX U8418 ( .IN0(data_mem_out_wire[73]), .IN1(data_mem_out_wire[105]), .SEL(
        N37), .F(n8376) );
  MUX U8419 ( .IN0(data_mem_out_wire[9]), .IN1(data_mem_out_wire[41]), .SEL(
        N37), .F(n8377) );
  MUX U8420 ( .IN0(n8377), .IN1(n8376), .SEL(N38), .F(n8378) );
  MUX U8421 ( .IN0(n8378), .IN1(n8375), .SEL(N39), .F(n8379) );
  MUX U8422 ( .IN0(n8379), .IN1(n8372), .SEL(N40), .F(n8380) );
  MUX U8423 ( .IN0(n8380), .IN1(n8365), .SEL(N41), .F(n8381) );
  MUX U8424 ( .IN0(n8381), .IN1(n8350), .SEL(N42), .F(N736) );
  MUX U8425 ( .IN0(data_mem_out_wire[1994]), .IN1(data_mem_out_wire[2026]), 
        .SEL(N37), .F(n8382) );
  MUX U8426 ( .IN0(data_mem_out_wire[1930]), .IN1(data_mem_out_wire[1962]), 
        .SEL(N37), .F(n8383) );
  MUX U8427 ( .IN0(n8383), .IN1(n8382), .SEL(N38), .F(n8384) );
  MUX U8428 ( .IN0(data_mem_out_wire[1866]), .IN1(data_mem_out_wire[1898]), 
        .SEL(N37), .F(n8385) );
  MUX U8429 ( .IN0(data_mem_out_wire[1802]), .IN1(data_mem_out_wire[1834]), 
        .SEL(N37), .F(n8386) );
  MUX U8430 ( .IN0(n8386), .IN1(n8385), .SEL(N38), .F(n8387) );
  MUX U8431 ( .IN0(n8387), .IN1(n8384), .SEL(N39), .F(n8388) );
  MUX U8432 ( .IN0(data_mem_out_wire[1738]), .IN1(data_mem_out_wire[1770]), 
        .SEL(N37), .F(n8389) );
  MUX U8433 ( .IN0(data_mem_out_wire[1674]), .IN1(data_mem_out_wire[1706]), 
        .SEL(N37), .F(n8390) );
  MUX U8434 ( .IN0(n8390), .IN1(n8389), .SEL(N38), .F(n8391) );
  MUX U8435 ( .IN0(data_mem_out_wire[1610]), .IN1(data_mem_out_wire[1642]), 
        .SEL(N37), .F(n8392) );
  MUX U8436 ( .IN0(data_mem_out_wire[1546]), .IN1(data_mem_out_wire[1578]), 
        .SEL(N37), .F(n8393) );
  MUX U8437 ( .IN0(n8393), .IN1(n8392), .SEL(N38), .F(n8394) );
  MUX U8438 ( .IN0(n8394), .IN1(n8391), .SEL(N39), .F(n8395) );
  MUX U8439 ( .IN0(n8395), .IN1(n8388), .SEL(N40), .F(n8396) );
  MUX U8440 ( .IN0(data_mem_out_wire[1482]), .IN1(data_mem_out_wire[1514]), 
        .SEL(N37), .F(n8397) );
  MUX U8441 ( .IN0(data_mem_out_wire[1418]), .IN1(data_mem_out_wire[1450]), 
        .SEL(N37), .F(n8398) );
  MUX U8442 ( .IN0(n8398), .IN1(n8397), .SEL(N38), .F(n8399) );
  MUX U8443 ( .IN0(data_mem_out_wire[1354]), .IN1(data_mem_out_wire[1386]), 
        .SEL(N37), .F(n8400) );
  MUX U8444 ( .IN0(data_mem_out_wire[1290]), .IN1(data_mem_out_wire[1322]), 
        .SEL(N37), .F(n8401) );
  MUX U8445 ( .IN0(n8401), .IN1(n8400), .SEL(N38), .F(n8402) );
  MUX U8446 ( .IN0(n8402), .IN1(n8399), .SEL(N39), .F(n8403) );
  MUX U8447 ( .IN0(data_mem_out_wire[1226]), .IN1(data_mem_out_wire[1258]), 
        .SEL(N37), .F(n8404) );
  MUX U8448 ( .IN0(data_mem_out_wire[1162]), .IN1(data_mem_out_wire[1194]), 
        .SEL(N37), .F(n8405) );
  MUX U8449 ( .IN0(n8405), .IN1(n8404), .SEL(N38), .F(n8406) );
  MUX U8450 ( .IN0(data_mem_out_wire[1098]), .IN1(data_mem_out_wire[1130]), 
        .SEL(N37), .F(n8407) );
  MUX U8451 ( .IN0(data_mem_out_wire[1034]), .IN1(data_mem_out_wire[1066]), 
        .SEL(N37), .F(n8408) );
  MUX U8452 ( .IN0(n8408), .IN1(n8407), .SEL(N38), .F(n8409) );
  MUX U8453 ( .IN0(n8409), .IN1(n8406), .SEL(N39), .F(n8410) );
  MUX U8454 ( .IN0(n8410), .IN1(n8403), .SEL(N40), .F(n8411) );
  MUX U8455 ( .IN0(n8411), .IN1(n8396), .SEL(N41), .F(n8412) );
  MUX U8456 ( .IN0(data_mem_out_wire[970]), .IN1(data_mem_out_wire[1002]), 
        .SEL(N37), .F(n8413) );
  MUX U8457 ( .IN0(data_mem_out_wire[906]), .IN1(data_mem_out_wire[938]), 
        .SEL(N37), .F(n8414) );
  MUX U8458 ( .IN0(n8414), .IN1(n8413), .SEL(N38), .F(n8415) );
  MUX U8459 ( .IN0(data_mem_out_wire[842]), .IN1(data_mem_out_wire[874]), 
        .SEL(N37), .F(n8416) );
  MUX U8460 ( .IN0(data_mem_out_wire[778]), .IN1(data_mem_out_wire[810]), 
        .SEL(N37), .F(n8417) );
  MUX U8461 ( .IN0(n8417), .IN1(n8416), .SEL(N38), .F(n8418) );
  MUX U8462 ( .IN0(n8418), .IN1(n8415), .SEL(N39), .F(n8419) );
  MUX U8463 ( .IN0(data_mem_out_wire[714]), .IN1(data_mem_out_wire[746]), 
        .SEL(N37), .F(n8420) );
  MUX U8464 ( .IN0(data_mem_out_wire[650]), .IN1(data_mem_out_wire[682]), 
        .SEL(N37), .F(n8421) );
  MUX U8465 ( .IN0(n8421), .IN1(n8420), .SEL(N38), .F(n8422) );
  MUX U8466 ( .IN0(data_mem_out_wire[586]), .IN1(data_mem_out_wire[618]), 
        .SEL(N37), .F(n8423) );
  MUX U8467 ( .IN0(data_mem_out_wire[522]), .IN1(data_mem_out_wire[554]), 
        .SEL(N37), .F(n8424) );
  MUX U8468 ( .IN0(n8424), .IN1(n8423), .SEL(N38), .F(n8425) );
  MUX U8469 ( .IN0(n8425), .IN1(n8422), .SEL(N39), .F(n8426) );
  MUX U8470 ( .IN0(n8426), .IN1(n8419), .SEL(N40), .F(n8427) );
  MUX U8471 ( .IN0(data_mem_out_wire[458]), .IN1(data_mem_out_wire[490]), 
        .SEL(N37), .F(n8428) );
  MUX U8472 ( .IN0(data_mem_out_wire[394]), .IN1(data_mem_out_wire[426]), 
        .SEL(N37), .F(n8429) );
  MUX U8473 ( .IN0(n8429), .IN1(n8428), .SEL(N38), .F(n8430) );
  MUX U8474 ( .IN0(data_mem_out_wire[330]), .IN1(data_mem_out_wire[362]), 
        .SEL(N37), .F(n8431) );
  MUX U8475 ( .IN0(data_mem_out_wire[266]), .IN1(data_mem_out_wire[298]), 
        .SEL(N37), .F(n8432) );
  MUX U8476 ( .IN0(n8432), .IN1(n8431), .SEL(N38), .F(n8433) );
  MUX U8477 ( .IN0(n8433), .IN1(n8430), .SEL(N39), .F(n8434) );
  MUX U8478 ( .IN0(data_mem_out_wire[202]), .IN1(data_mem_out_wire[234]), 
        .SEL(N37), .F(n8435) );
  MUX U8479 ( .IN0(data_mem_out_wire[138]), .IN1(data_mem_out_wire[170]), 
        .SEL(N37), .F(n8436) );
  MUX U8480 ( .IN0(n8436), .IN1(n8435), .SEL(N38), .F(n8437) );
  MUX U8481 ( .IN0(data_mem_out_wire[74]), .IN1(data_mem_out_wire[106]), .SEL(
        N37), .F(n8438) );
  MUX U8482 ( .IN0(data_mem_out_wire[10]), .IN1(data_mem_out_wire[42]), .SEL(
        N37), .F(n8439) );
  MUX U8483 ( .IN0(n8439), .IN1(n8438), .SEL(N38), .F(n8440) );
  MUX U8484 ( .IN0(n8440), .IN1(n8437), .SEL(N39), .F(n8441) );
  MUX U8485 ( .IN0(n8441), .IN1(n8434), .SEL(N40), .F(n8442) );
  MUX U8486 ( .IN0(n8442), .IN1(n8427), .SEL(N41), .F(n8443) );
  MUX U8487 ( .IN0(n8443), .IN1(n8412), .SEL(N42), .F(N735) );
  MUX U8488 ( .IN0(data_mem_out_wire[1995]), .IN1(data_mem_out_wire[2027]), 
        .SEL(N37), .F(n8444) );
  MUX U8489 ( .IN0(data_mem_out_wire[1931]), .IN1(data_mem_out_wire[1963]), 
        .SEL(N37), .F(n8445) );
  MUX U8490 ( .IN0(n8445), .IN1(n8444), .SEL(N38), .F(n8446) );
  MUX U8491 ( .IN0(data_mem_out_wire[1867]), .IN1(data_mem_out_wire[1899]), 
        .SEL(N37), .F(n8447) );
  MUX U8492 ( .IN0(data_mem_out_wire[1803]), .IN1(data_mem_out_wire[1835]), 
        .SEL(N37), .F(n8448) );
  MUX U8493 ( .IN0(n8448), .IN1(n8447), .SEL(N38), .F(n8449) );
  MUX U8494 ( .IN0(n8449), .IN1(n8446), .SEL(N39), .F(n8450) );
  MUX U8495 ( .IN0(data_mem_out_wire[1739]), .IN1(data_mem_out_wire[1771]), 
        .SEL(N37), .F(n8451) );
  MUX U8496 ( .IN0(data_mem_out_wire[1675]), .IN1(data_mem_out_wire[1707]), 
        .SEL(N37), .F(n8452) );
  MUX U8497 ( .IN0(n8452), .IN1(n8451), .SEL(N38), .F(n8453) );
  MUX U8498 ( .IN0(data_mem_out_wire[1611]), .IN1(data_mem_out_wire[1643]), 
        .SEL(N37), .F(n8454) );
  MUX U8499 ( .IN0(data_mem_out_wire[1547]), .IN1(data_mem_out_wire[1579]), 
        .SEL(N37), .F(n8455) );
  MUX U8500 ( .IN0(n8455), .IN1(n8454), .SEL(N38), .F(n8456) );
  MUX U8501 ( .IN0(n8456), .IN1(n8453), .SEL(N39), .F(n8457) );
  MUX U8502 ( .IN0(n8457), .IN1(n8450), .SEL(N40), .F(n8458) );
  MUX U8503 ( .IN0(data_mem_out_wire[1483]), .IN1(data_mem_out_wire[1515]), 
        .SEL(N37), .F(n8459) );
  MUX U8504 ( .IN0(data_mem_out_wire[1419]), .IN1(data_mem_out_wire[1451]), 
        .SEL(N37), .F(n8460) );
  MUX U8505 ( .IN0(n8460), .IN1(n8459), .SEL(N38), .F(n8461) );
  MUX U8506 ( .IN0(data_mem_out_wire[1355]), .IN1(data_mem_out_wire[1387]), 
        .SEL(N37), .F(n8462) );
  MUX U8507 ( .IN0(data_mem_out_wire[1291]), .IN1(data_mem_out_wire[1323]), 
        .SEL(N37), .F(n8463) );
  MUX U8508 ( .IN0(n8463), .IN1(n8462), .SEL(N38), .F(n8464) );
  MUX U8509 ( .IN0(n8464), .IN1(n8461), .SEL(N39), .F(n8465) );
  MUX U8510 ( .IN0(data_mem_out_wire[1227]), .IN1(data_mem_out_wire[1259]), 
        .SEL(N37), .F(n8466) );
  MUX U8511 ( .IN0(data_mem_out_wire[1163]), .IN1(data_mem_out_wire[1195]), 
        .SEL(N37), .F(n8467) );
  MUX U8512 ( .IN0(n8467), .IN1(n8466), .SEL(N38), .F(n8468) );
  MUX U8513 ( .IN0(data_mem_out_wire[1099]), .IN1(data_mem_out_wire[1131]), 
        .SEL(N37), .F(n8469) );
  MUX U8514 ( .IN0(data_mem_out_wire[1035]), .IN1(data_mem_out_wire[1067]), 
        .SEL(N37), .F(n8470) );
  MUX U8515 ( .IN0(n8470), .IN1(n8469), .SEL(N38), .F(n8471) );
  MUX U8516 ( .IN0(n8471), .IN1(n8468), .SEL(N39), .F(n8472) );
  MUX U8517 ( .IN0(n8472), .IN1(n8465), .SEL(N40), .F(n8473) );
  MUX U8518 ( .IN0(n8473), .IN1(n8458), .SEL(N41), .F(n8474) );
  MUX U8519 ( .IN0(data_mem_out_wire[971]), .IN1(data_mem_out_wire[1003]), 
        .SEL(N37), .F(n8475) );
  MUX U8520 ( .IN0(data_mem_out_wire[907]), .IN1(data_mem_out_wire[939]), 
        .SEL(N37), .F(n8476) );
  MUX U8521 ( .IN0(n8476), .IN1(n8475), .SEL(N38), .F(n8477) );
  MUX U8522 ( .IN0(data_mem_out_wire[843]), .IN1(data_mem_out_wire[875]), 
        .SEL(N37), .F(n8478) );
  MUX U8523 ( .IN0(data_mem_out_wire[779]), .IN1(data_mem_out_wire[811]), 
        .SEL(N37), .F(n8479) );
  MUX U8524 ( .IN0(n8479), .IN1(n8478), .SEL(N38), .F(n8480) );
  MUX U8525 ( .IN0(n8480), .IN1(n8477), .SEL(N39), .F(n8481) );
  MUX U8526 ( .IN0(data_mem_out_wire[715]), .IN1(data_mem_out_wire[747]), 
        .SEL(N37), .F(n8482) );
  MUX U8527 ( .IN0(data_mem_out_wire[651]), .IN1(data_mem_out_wire[683]), 
        .SEL(N37), .F(n8483) );
  MUX U8528 ( .IN0(n8483), .IN1(n8482), .SEL(N38), .F(n8484) );
  MUX U8529 ( .IN0(data_mem_out_wire[587]), .IN1(data_mem_out_wire[619]), 
        .SEL(N37), .F(n8485) );
  MUX U8530 ( .IN0(data_mem_out_wire[523]), .IN1(data_mem_out_wire[555]), 
        .SEL(N37), .F(n8486) );
  MUX U8531 ( .IN0(n8486), .IN1(n8485), .SEL(N38), .F(n8487) );
  MUX U8532 ( .IN0(n8487), .IN1(n8484), .SEL(N39), .F(n8488) );
  MUX U8533 ( .IN0(n8488), .IN1(n8481), .SEL(N40), .F(n8489) );
  MUX U8534 ( .IN0(data_mem_out_wire[459]), .IN1(data_mem_out_wire[491]), 
        .SEL(N37), .F(n8490) );
  MUX U8535 ( .IN0(data_mem_out_wire[395]), .IN1(data_mem_out_wire[427]), 
        .SEL(N37), .F(n8491) );
  MUX U8536 ( .IN0(n8491), .IN1(n8490), .SEL(N38), .F(n8492) );
  MUX U8537 ( .IN0(data_mem_out_wire[331]), .IN1(data_mem_out_wire[363]), 
        .SEL(N37), .F(n8493) );
  MUX U8538 ( .IN0(data_mem_out_wire[267]), .IN1(data_mem_out_wire[299]), 
        .SEL(N37), .F(n8494) );
  MUX U8539 ( .IN0(n8494), .IN1(n8493), .SEL(N38), .F(n8495) );
  MUX U8540 ( .IN0(n8495), .IN1(n8492), .SEL(N39), .F(n8496) );
  MUX U8541 ( .IN0(data_mem_out_wire[203]), .IN1(data_mem_out_wire[235]), 
        .SEL(N37), .F(n8497) );
  MUX U8542 ( .IN0(data_mem_out_wire[139]), .IN1(data_mem_out_wire[171]), 
        .SEL(N37), .F(n8498) );
  MUX U8543 ( .IN0(n8498), .IN1(n8497), .SEL(N38), .F(n8499) );
  MUX U8544 ( .IN0(data_mem_out_wire[75]), .IN1(data_mem_out_wire[107]), .SEL(
        N37), .F(n8500) );
  MUX U8545 ( .IN0(data_mem_out_wire[11]), .IN1(data_mem_out_wire[43]), .SEL(
        N37), .F(n8501) );
  MUX U8546 ( .IN0(n8501), .IN1(n8500), .SEL(N38), .F(n8502) );
  MUX U8547 ( .IN0(n8502), .IN1(n8499), .SEL(N39), .F(n8503) );
  MUX U8548 ( .IN0(n8503), .IN1(n8496), .SEL(N40), .F(n8504) );
  MUX U8549 ( .IN0(n8504), .IN1(n8489), .SEL(N41), .F(n8505) );
  MUX U8550 ( .IN0(n8505), .IN1(n8474), .SEL(N42), .F(N734) );
  MUX U8551 ( .IN0(data_mem_out_wire[1996]), .IN1(data_mem_out_wire[2028]), 
        .SEL(N37), .F(n8506) );
  MUX U8552 ( .IN0(data_mem_out_wire[1932]), .IN1(data_mem_out_wire[1964]), 
        .SEL(N37), .F(n8507) );
  MUX U8553 ( .IN0(n8507), .IN1(n8506), .SEL(N38), .F(n8508) );
  MUX U8554 ( .IN0(data_mem_out_wire[1868]), .IN1(data_mem_out_wire[1900]), 
        .SEL(N37), .F(n8509) );
  MUX U8555 ( .IN0(data_mem_out_wire[1804]), .IN1(data_mem_out_wire[1836]), 
        .SEL(N37), .F(n8510) );
  MUX U8556 ( .IN0(n8510), .IN1(n8509), .SEL(N38), .F(n8511) );
  MUX U8557 ( .IN0(n8511), .IN1(n8508), .SEL(N39), .F(n8512) );
  MUX U8558 ( .IN0(data_mem_out_wire[1740]), .IN1(data_mem_out_wire[1772]), 
        .SEL(N37), .F(n8513) );
  MUX U8559 ( .IN0(data_mem_out_wire[1676]), .IN1(data_mem_out_wire[1708]), 
        .SEL(N37), .F(n8514) );
  MUX U8560 ( .IN0(n8514), .IN1(n8513), .SEL(N38), .F(n8515) );
  MUX U8561 ( .IN0(data_mem_out_wire[1612]), .IN1(data_mem_out_wire[1644]), 
        .SEL(N37), .F(n8516) );
  MUX U8562 ( .IN0(data_mem_out_wire[1548]), .IN1(data_mem_out_wire[1580]), 
        .SEL(N37), .F(n8517) );
  MUX U8563 ( .IN0(n8517), .IN1(n8516), .SEL(N38), .F(n8518) );
  MUX U8564 ( .IN0(n8518), .IN1(n8515), .SEL(N39), .F(n8519) );
  MUX U8565 ( .IN0(n8519), .IN1(n8512), .SEL(N40), .F(n8520) );
  MUX U8566 ( .IN0(data_mem_out_wire[1484]), .IN1(data_mem_out_wire[1516]), 
        .SEL(N37), .F(n8521) );
  MUX U8567 ( .IN0(data_mem_out_wire[1420]), .IN1(data_mem_out_wire[1452]), 
        .SEL(N37), .F(n8522) );
  MUX U8568 ( .IN0(n8522), .IN1(n8521), .SEL(N38), .F(n8523) );
  MUX U8569 ( .IN0(data_mem_out_wire[1356]), .IN1(data_mem_out_wire[1388]), 
        .SEL(N37), .F(n8524) );
  MUX U8570 ( .IN0(data_mem_out_wire[1292]), .IN1(data_mem_out_wire[1324]), 
        .SEL(N37), .F(n8525) );
  MUX U8571 ( .IN0(n8525), .IN1(n8524), .SEL(N38), .F(n8526) );
  MUX U8572 ( .IN0(n8526), .IN1(n8523), .SEL(N39), .F(n8527) );
  MUX U8573 ( .IN0(data_mem_out_wire[1228]), .IN1(data_mem_out_wire[1260]), 
        .SEL(N37), .F(n8528) );
  MUX U8574 ( .IN0(data_mem_out_wire[1164]), .IN1(data_mem_out_wire[1196]), 
        .SEL(N37), .F(n8529) );
  MUX U8575 ( .IN0(n8529), .IN1(n8528), .SEL(N38), .F(n8530) );
  MUX U8576 ( .IN0(data_mem_out_wire[1100]), .IN1(data_mem_out_wire[1132]), 
        .SEL(N37), .F(n8531) );
  MUX U8577 ( .IN0(data_mem_out_wire[1036]), .IN1(data_mem_out_wire[1068]), 
        .SEL(N37), .F(n8532) );
  MUX U8578 ( .IN0(n8532), .IN1(n8531), .SEL(N38), .F(n8533) );
  MUX U8579 ( .IN0(n8533), .IN1(n8530), .SEL(N39), .F(n8534) );
  MUX U8580 ( .IN0(n8534), .IN1(n8527), .SEL(N40), .F(n8535) );
  MUX U8581 ( .IN0(n8535), .IN1(n8520), .SEL(N41), .F(n8536) );
  MUX U8582 ( .IN0(data_mem_out_wire[972]), .IN1(data_mem_out_wire[1004]), 
        .SEL(N37), .F(n8537) );
  MUX U8583 ( .IN0(data_mem_out_wire[908]), .IN1(data_mem_out_wire[940]), 
        .SEL(N37), .F(n8538) );
  MUX U8584 ( .IN0(n8538), .IN1(n8537), .SEL(N38), .F(n8539) );
  MUX U8585 ( .IN0(data_mem_out_wire[844]), .IN1(data_mem_out_wire[876]), 
        .SEL(N37), .F(n8540) );
  MUX U8586 ( .IN0(data_mem_out_wire[780]), .IN1(data_mem_out_wire[812]), 
        .SEL(N37), .F(n8541) );
  MUX U8587 ( .IN0(n8541), .IN1(n8540), .SEL(N38), .F(n8542) );
  MUX U8588 ( .IN0(n8542), .IN1(n8539), .SEL(N39), .F(n8543) );
  MUX U8589 ( .IN0(data_mem_out_wire[716]), .IN1(data_mem_out_wire[748]), 
        .SEL(N37), .F(n8544) );
  MUX U8590 ( .IN0(data_mem_out_wire[652]), .IN1(data_mem_out_wire[684]), 
        .SEL(N37), .F(n8545) );
  MUX U8591 ( .IN0(n8545), .IN1(n8544), .SEL(N38), .F(n8546) );
  MUX U8592 ( .IN0(data_mem_out_wire[588]), .IN1(data_mem_out_wire[620]), 
        .SEL(N37), .F(n8547) );
  MUX U8593 ( .IN0(data_mem_out_wire[524]), .IN1(data_mem_out_wire[556]), 
        .SEL(N37), .F(n8548) );
  MUX U8594 ( .IN0(n8548), .IN1(n8547), .SEL(N38), .F(n8549) );
  MUX U8595 ( .IN0(n8549), .IN1(n8546), .SEL(N39), .F(n8550) );
  MUX U8596 ( .IN0(n8550), .IN1(n8543), .SEL(N40), .F(n8551) );
  MUX U8597 ( .IN0(data_mem_out_wire[460]), .IN1(data_mem_out_wire[492]), 
        .SEL(N37), .F(n8552) );
  MUX U8598 ( .IN0(data_mem_out_wire[396]), .IN1(data_mem_out_wire[428]), 
        .SEL(N37), .F(n8553) );
  MUX U8599 ( .IN0(n8553), .IN1(n8552), .SEL(N38), .F(n8554) );
  MUX U8600 ( .IN0(data_mem_out_wire[332]), .IN1(data_mem_out_wire[364]), 
        .SEL(N37), .F(n8555) );
  MUX U8601 ( .IN0(data_mem_out_wire[268]), .IN1(data_mem_out_wire[300]), 
        .SEL(N37), .F(n8556) );
  MUX U8602 ( .IN0(n8556), .IN1(n8555), .SEL(N38), .F(n8557) );
  MUX U8603 ( .IN0(n8557), .IN1(n8554), .SEL(N39), .F(n8558) );
  MUX U8604 ( .IN0(data_mem_out_wire[204]), .IN1(data_mem_out_wire[236]), 
        .SEL(N37), .F(n8559) );
  MUX U8605 ( .IN0(data_mem_out_wire[140]), .IN1(data_mem_out_wire[172]), 
        .SEL(N37), .F(n8560) );
  MUX U8606 ( .IN0(n8560), .IN1(n8559), .SEL(N38), .F(n8561) );
  MUX U8607 ( .IN0(data_mem_out_wire[76]), .IN1(data_mem_out_wire[108]), .SEL(
        N37), .F(n8562) );
  MUX U8608 ( .IN0(data_mem_out_wire[12]), .IN1(data_mem_out_wire[44]), .SEL(
        N37), .F(n8563) );
  MUX U8609 ( .IN0(n8563), .IN1(n8562), .SEL(N38), .F(n8564) );
  MUX U8610 ( .IN0(n8564), .IN1(n8561), .SEL(N39), .F(n8565) );
  MUX U8611 ( .IN0(n8565), .IN1(n8558), .SEL(N40), .F(n8566) );
  MUX U8612 ( .IN0(n8566), .IN1(n8551), .SEL(N41), .F(n8567) );
  MUX U8613 ( .IN0(n8567), .IN1(n8536), .SEL(N42), .F(N733) );
  MUX U8614 ( .IN0(data_mem_out_wire[1997]), .IN1(data_mem_out_wire[2029]), 
        .SEL(N37), .F(n8568) );
  MUX U8615 ( .IN0(data_mem_out_wire[1933]), .IN1(data_mem_out_wire[1965]), 
        .SEL(N37), .F(n8569) );
  MUX U8616 ( .IN0(n8569), .IN1(n8568), .SEL(N38), .F(n8570) );
  MUX U8617 ( .IN0(data_mem_out_wire[1869]), .IN1(data_mem_out_wire[1901]), 
        .SEL(N37), .F(n8571) );
  MUX U8618 ( .IN0(data_mem_out_wire[1805]), .IN1(data_mem_out_wire[1837]), 
        .SEL(N37), .F(n8572) );
  MUX U8619 ( .IN0(n8572), .IN1(n8571), .SEL(N38), .F(n8573) );
  MUX U8620 ( .IN0(n8573), .IN1(n8570), .SEL(N39), .F(n8574) );
  MUX U8621 ( .IN0(data_mem_out_wire[1741]), .IN1(data_mem_out_wire[1773]), 
        .SEL(N37), .F(n8575) );
  MUX U8622 ( .IN0(data_mem_out_wire[1677]), .IN1(data_mem_out_wire[1709]), 
        .SEL(N37), .F(n8576) );
  MUX U8623 ( .IN0(n8576), .IN1(n8575), .SEL(N38), .F(n8577) );
  MUX U8624 ( .IN0(data_mem_out_wire[1613]), .IN1(data_mem_out_wire[1645]), 
        .SEL(N37), .F(n8578) );
  MUX U8625 ( .IN0(data_mem_out_wire[1549]), .IN1(data_mem_out_wire[1581]), 
        .SEL(N37), .F(n8579) );
  MUX U8626 ( .IN0(n8579), .IN1(n8578), .SEL(N38), .F(n8580) );
  MUX U8627 ( .IN0(n8580), .IN1(n8577), .SEL(N39), .F(n8581) );
  MUX U8628 ( .IN0(n8581), .IN1(n8574), .SEL(N40), .F(n8582) );
  MUX U8629 ( .IN0(data_mem_out_wire[1485]), .IN1(data_mem_out_wire[1517]), 
        .SEL(N37), .F(n8583) );
  MUX U8630 ( .IN0(data_mem_out_wire[1421]), .IN1(data_mem_out_wire[1453]), 
        .SEL(N37), .F(n8584) );
  MUX U8631 ( .IN0(n8584), .IN1(n8583), .SEL(N38), .F(n8585) );
  MUX U8632 ( .IN0(data_mem_out_wire[1357]), .IN1(data_mem_out_wire[1389]), 
        .SEL(N37), .F(n8586) );
  MUX U8633 ( .IN0(data_mem_out_wire[1293]), .IN1(data_mem_out_wire[1325]), 
        .SEL(N37), .F(n8587) );
  MUX U8634 ( .IN0(n8587), .IN1(n8586), .SEL(N38), .F(n8588) );
  MUX U8635 ( .IN0(n8588), .IN1(n8585), .SEL(N39), .F(n8589) );
  MUX U8636 ( .IN0(data_mem_out_wire[1229]), .IN1(data_mem_out_wire[1261]), 
        .SEL(N37), .F(n8590) );
  MUX U8637 ( .IN0(data_mem_out_wire[1165]), .IN1(data_mem_out_wire[1197]), 
        .SEL(N37), .F(n8591) );
  MUX U8638 ( .IN0(n8591), .IN1(n8590), .SEL(N38), .F(n8592) );
  MUX U8639 ( .IN0(data_mem_out_wire[1101]), .IN1(data_mem_out_wire[1133]), 
        .SEL(N37), .F(n8593) );
  MUX U8640 ( .IN0(data_mem_out_wire[1037]), .IN1(data_mem_out_wire[1069]), 
        .SEL(N37), .F(n8594) );
  MUX U8641 ( .IN0(n8594), .IN1(n8593), .SEL(N38), .F(n8595) );
  MUX U8642 ( .IN0(n8595), .IN1(n8592), .SEL(N39), .F(n8596) );
  MUX U8643 ( .IN0(n8596), .IN1(n8589), .SEL(N40), .F(n8597) );
  MUX U8644 ( .IN0(n8597), .IN1(n8582), .SEL(N41), .F(n8598) );
  MUX U8645 ( .IN0(data_mem_out_wire[973]), .IN1(data_mem_out_wire[1005]), 
        .SEL(N37), .F(n8599) );
  MUX U8646 ( .IN0(data_mem_out_wire[909]), .IN1(data_mem_out_wire[941]), 
        .SEL(N37), .F(n8600) );
  MUX U8647 ( .IN0(n8600), .IN1(n8599), .SEL(N38), .F(n8601) );
  MUX U8648 ( .IN0(data_mem_out_wire[845]), .IN1(data_mem_out_wire[877]), 
        .SEL(N37), .F(n8602) );
  MUX U8649 ( .IN0(data_mem_out_wire[781]), .IN1(data_mem_out_wire[813]), 
        .SEL(N37), .F(n8603) );
  MUX U8650 ( .IN0(n8603), .IN1(n8602), .SEL(N38), .F(n8604) );
  MUX U8651 ( .IN0(n8604), .IN1(n8601), .SEL(N39), .F(n8605) );
  MUX U8652 ( .IN0(data_mem_out_wire[717]), .IN1(data_mem_out_wire[749]), 
        .SEL(N37), .F(n8606) );
  MUX U8653 ( .IN0(data_mem_out_wire[653]), .IN1(data_mem_out_wire[685]), 
        .SEL(N37), .F(n8607) );
  MUX U8654 ( .IN0(n8607), .IN1(n8606), .SEL(N38), .F(n8608) );
  MUX U8655 ( .IN0(data_mem_out_wire[589]), .IN1(data_mem_out_wire[621]), 
        .SEL(N37), .F(n8609) );
  MUX U8656 ( .IN0(data_mem_out_wire[525]), .IN1(data_mem_out_wire[557]), 
        .SEL(N37), .F(n8610) );
  MUX U8657 ( .IN0(n8610), .IN1(n8609), .SEL(N38), .F(n8611) );
  MUX U8658 ( .IN0(n8611), .IN1(n8608), .SEL(N39), .F(n8612) );
  MUX U8659 ( .IN0(n8612), .IN1(n8605), .SEL(N40), .F(n8613) );
  MUX U8660 ( .IN0(data_mem_out_wire[461]), .IN1(data_mem_out_wire[493]), 
        .SEL(N37), .F(n8614) );
  MUX U8661 ( .IN0(data_mem_out_wire[397]), .IN1(data_mem_out_wire[429]), 
        .SEL(N37), .F(n8615) );
  MUX U8662 ( .IN0(n8615), .IN1(n8614), .SEL(N38), .F(n8616) );
  MUX U8663 ( .IN0(data_mem_out_wire[333]), .IN1(data_mem_out_wire[365]), 
        .SEL(N37), .F(n8617) );
  MUX U8664 ( .IN0(data_mem_out_wire[269]), .IN1(data_mem_out_wire[301]), 
        .SEL(N37), .F(n8618) );
  MUX U8665 ( .IN0(n8618), .IN1(n8617), .SEL(N38), .F(n8619) );
  MUX U8666 ( .IN0(n8619), .IN1(n8616), .SEL(N39), .F(n8620) );
  MUX U8667 ( .IN0(data_mem_out_wire[205]), .IN1(data_mem_out_wire[237]), 
        .SEL(N37), .F(n8621) );
  MUX U8668 ( .IN0(data_mem_out_wire[141]), .IN1(data_mem_out_wire[173]), 
        .SEL(N37), .F(n8622) );
  MUX U8669 ( .IN0(n8622), .IN1(n8621), .SEL(N38), .F(n8623) );
  MUX U8670 ( .IN0(data_mem_out_wire[77]), .IN1(data_mem_out_wire[109]), .SEL(
        N37), .F(n8624) );
  MUX U8671 ( .IN0(data_mem_out_wire[13]), .IN1(data_mem_out_wire[45]), .SEL(
        N37), .F(n8625) );
  MUX U8672 ( .IN0(n8625), .IN1(n8624), .SEL(N38), .F(n8626) );
  MUX U8673 ( .IN0(n8626), .IN1(n8623), .SEL(N39), .F(n8627) );
  MUX U8674 ( .IN0(n8627), .IN1(n8620), .SEL(N40), .F(n8628) );
  MUX U8675 ( .IN0(n8628), .IN1(n8613), .SEL(N41), .F(n8629) );
  MUX U8676 ( .IN0(n8629), .IN1(n8598), .SEL(N42), .F(N732) );
  MUX U8677 ( .IN0(data_mem_out_wire[1998]), .IN1(data_mem_out_wire[2030]), 
        .SEL(N37), .F(n8630) );
  MUX U8678 ( .IN0(data_mem_out_wire[1934]), .IN1(data_mem_out_wire[1966]), 
        .SEL(N37), .F(n8631) );
  MUX U8679 ( .IN0(n8631), .IN1(n8630), .SEL(N38), .F(n8632) );
  MUX U8680 ( .IN0(data_mem_out_wire[1870]), .IN1(data_mem_out_wire[1902]), 
        .SEL(N37), .F(n8633) );
  MUX U8681 ( .IN0(data_mem_out_wire[1806]), .IN1(data_mem_out_wire[1838]), 
        .SEL(N37), .F(n8634) );
  MUX U8682 ( .IN0(n8634), .IN1(n8633), .SEL(N38), .F(n8635) );
  MUX U8683 ( .IN0(n8635), .IN1(n8632), .SEL(N39), .F(n8636) );
  MUX U8684 ( .IN0(data_mem_out_wire[1742]), .IN1(data_mem_out_wire[1774]), 
        .SEL(N37), .F(n8637) );
  MUX U8685 ( .IN0(data_mem_out_wire[1678]), .IN1(data_mem_out_wire[1710]), 
        .SEL(N37), .F(n8638) );
  MUX U8686 ( .IN0(n8638), .IN1(n8637), .SEL(N38), .F(n8639) );
  MUX U8687 ( .IN0(data_mem_out_wire[1614]), .IN1(data_mem_out_wire[1646]), 
        .SEL(N37), .F(n8640) );
  MUX U8688 ( .IN0(data_mem_out_wire[1550]), .IN1(data_mem_out_wire[1582]), 
        .SEL(N37), .F(n8641) );
  MUX U8689 ( .IN0(n8641), .IN1(n8640), .SEL(N38), .F(n8642) );
  MUX U8690 ( .IN0(n8642), .IN1(n8639), .SEL(N39), .F(n8643) );
  MUX U8691 ( .IN0(n8643), .IN1(n8636), .SEL(N40), .F(n8644) );
  MUX U8692 ( .IN0(data_mem_out_wire[1486]), .IN1(data_mem_out_wire[1518]), 
        .SEL(N37), .F(n8645) );
  MUX U8693 ( .IN0(data_mem_out_wire[1422]), .IN1(data_mem_out_wire[1454]), 
        .SEL(N37), .F(n8646) );
  MUX U8694 ( .IN0(n8646), .IN1(n8645), .SEL(N38), .F(n8647) );
  MUX U8695 ( .IN0(data_mem_out_wire[1358]), .IN1(data_mem_out_wire[1390]), 
        .SEL(N37), .F(n8648) );
  MUX U8696 ( .IN0(data_mem_out_wire[1294]), .IN1(data_mem_out_wire[1326]), 
        .SEL(N37), .F(n8649) );
  MUX U8697 ( .IN0(n8649), .IN1(n8648), .SEL(N38), .F(n8650) );
  MUX U8698 ( .IN0(n8650), .IN1(n8647), .SEL(N39), .F(n8651) );
  MUX U8699 ( .IN0(data_mem_out_wire[1230]), .IN1(data_mem_out_wire[1262]), 
        .SEL(N37), .F(n8652) );
  MUX U8700 ( .IN0(data_mem_out_wire[1166]), .IN1(data_mem_out_wire[1198]), 
        .SEL(N37), .F(n8653) );
  MUX U8701 ( .IN0(n8653), .IN1(n8652), .SEL(N38), .F(n8654) );
  MUX U8702 ( .IN0(data_mem_out_wire[1102]), .IN1(data_mem_out_wire[1134]), 
        .SEL(N37), .F(n8655) );
  MUX U8703 ( .IN0(data_mem_out_wire[1038]), .IN1(data_mem_out_wire[1070]), 
        .SEL(N37), .F(n8656) );
  MUX U8704 ( .IN0(n8656), .IN1(n8655), .SEL(N38), .F(n8657) );
  MUX U8705 ( .IN0(n8657), .IN1(n8654), .SEL(N39), .F(n8658) );
  MUX U8706 ( .IN0(n8658), .IN1(n8651), .SEL(N40), .F(n8659) );
  MUX U8707 ( .IN0(n8659), .IN1(n8644), .SEL(N41), .F(n8660) );
  MUX U8708 ( .IN0(data_mem_out_wire[974]), .IN1(data_mem_out_wire[1006]), 
        .SEL(N37), .F(n8661) );
  MUX U8709 ( .IN0(data_mem_out_wire[910]), .IN1(data_mem_out_wire[942]), 
        .SEL(N37), .F(n8662) );
  MUX U8710 ( .IN0(n8662), .IN1(n8661), .SEL(N38), .F(n8663) );
  MUX U8711 ( .IN0(data_mem_out_wire[846]), .IN1(data_mem_out_wire[878]), 
        .SEL(N37), .F(n8664) );
  MUX U8712 ( .IN0(data_mem_out_wire[782]), .IN1(data_mem_out_wire[814]), 
        .SEL(N37), .F(n8665) );
  MUX U8713 ( .IN0(n8665), .IN1(n8664), .SEL(N38), .F(n8666) );
  MUX U8714 ( .IN0(n8666), .IN1(n8663), .SEL(N39), .F(n8667) );
  MUX U8715 ( .IN0(data_mem_out_wire[718]), .IN1(data_mem_out_wire[750]), 
        .SEL(N37), .F(n8668) );
  MUX U8716 ( .IN0(data_mem_out_wire[654]), .IN1(data_mem_out_wire[686]), 
        .SEL(N37), .F(n8669) );
  MUX U8717 ( .IN0(n8669), .IN1(n8668), .SEL(N38), .F(n8670) );
  MUX U8718 ( .IN0(data_mem_out_wire[590]), .IN1(data_mem_out_wire[622]), 
        .SEL(N37), .F(n8671) );
  MUX U8719 ( .IN0(data_mem_out_wire[526]), .IN1(data_mem_out_wire[558]), 
        .SEL(N37), .F(n8672) );
  MUX U8720 ( .IN0(n8672), .IN1(n8671), .SEL(N38), .F(n8673) );
  MUX U8721 ( .IN0(n8673), .IN1(n8670), .SEL(N39), .F(n8674) );
  MUX U8722 ( .IN0(n8674), .IN1(n8667), .SEL(N40), .F(n8675) );
  MUX U8723 ( .IN0(data_mem_out_wire[462]), .IN1(data_mem_out_wire[494]), 
        .SEL(N37), .F(n8676) );
  MUX U8724 ( .IN0(data_mem_out_wire[398]), .IN1(data_mem_out_wire[430]), 
        .SEL(N37), .F(n8677) );
  MUX U8725 ( .IN0(n8677), .IN1(n8676), .SEL(N38), .F(n8678) );
  MUX U8726 ( .IN0(data_mem_out_wire[334]), .IN1(data_mem_out_wire[366]), 
        .SEL(N37), .F(n8679) );
  MUX U8727 ( .IN0(data_mem_out_wire[270]), .IN1(data_mem_out_wire[302]), 
        .SEL(N37), .F(n8680) );
  MUX U8728 ( .IN0(n8680), .IN1(n8679), .SEL(N38), .F(n8681) );
  MUX U8729 ( .IN0(n8681), .IN1(n8678), .SEL(N39), .F(n8682) );
  MUX U8730 ( .IN0(data_mem_out_wire[206]), .IN1(data_mem_out_wire[238]), 
        .SEL(N37), .F(n8683) );
  MUX U8731 ( .IN0(data_mem_out_wire[142]), .IN1(data_mem_out_wire[174]), 
        .SEL(N37), .F(n8684) );
  MUX U8732 ( .IN0(n8684), .IN1(n8683), .SEL(N38), .F(n8685) );
  MUX U8733 ( .IN0(data_mem_out_wire[78]), .IN1(data_mem_out_wire[110]), .SEL(
        N37), .F(n8686) );
  MUX U8734 ( .IN0(data_mem_out_wire[14]), .IN1(data_mem_out_wire[46]), .SEL(
        N37), .F(n8687) );
  MUX U8735 ( .IN0(n8687), .IN1(n8686), .SEL(N38), .F(n8688) );
  MUX U8736 ( .IN0(n8688), .IN1(n8685), .SEL(N39), .F(n8689) );
  MUX U8737 ( .IN0(n8689), .IN1(n8682), .SEL(N40), .F(n8690) );
  MUX U8738 ( .IN0(n8690), .IN1(n8675), .SEL(N41), .F(n8691) );
  MUX U8739 ( .IN0(n8691), .IN1(n8660), .SEL(N42), .F(N731) );
  MUX U8740 ( .IN0(data_mem_out_wire[1999]), .IN1(data_mem_out_wire[2031]), 
        .SEL(N37), .F(n8692) );
  MUX U8741 ( .IN0(data_mem_out_wire[1935]), .IN1(data_mem_out_wire[1967]), 
        .SEL(N37), .F(n8693) );
  MUX U8742 ( .IN0(n8693), .IN1(n8692), .SEL(N38), .F(n8694) );
  MUX U8743 ( .IN0(data_mem_out_wire[1871]), .IN1(data_mem_out_wire[1903]), 
        .SEL(N37), .F(n8695) );
  MUX U8744 ( .IN0(data_mem_out_wire[1807]), .IN1(data_mem_out_wire[1839]), 
        .SEL(N37), .F(n8696) );
  MUX U8745 ( .IN0(n8696), .IN1(n8695), .SEL(N38), .F(n8697) );
  MUX U8746 ( .IN0(n8697), .IN1(n8694), .SEL(N39), .F(n8698) );
  MUX U8747 ( .IN0(data_mem_out_wire[1743]), .IN1(data_mem_out_wire[1775]), 
        .SEL(N37), .F(n8699) );
  MUX U8748 ( .IN0(data_mem_out_wire[1679]), .IN1(data_mem_out_wire[1711]), 
        .SEL(N37), .F(n8700) );
  MUX U8749 ( .IN0(n8700), .IN1(n8699), .SEL(N38), .F(n8701) );
  MUX U8750 ( .IN0(data_mem_out_wire[1615]), .IN1(data_mem_out_wire[1647]), 
        .SEL(N37), .F(n8702) );
  MUX U8751 ( .IN0(data_mem_out_wire[1551]), .IN1(data_mem_out_wire[1583]), 
        .SEL(N37), .F(n8703) );
  MUX U8752 ( .IN0(n8703), .IN1(n8702), .SEL(N38), .F(n8704) );
  MUX U8753 ( .IN0(n8704), .IN1(n8701), .SEL(N39), .F(n8705) );
  MUX U8754 ( .IN0(n8705), .IN1(n8698), .SEL(N40), .F(n8706) );
  MUX U8755 ( .IN0(data_mem_out_wire[1487]), .IN1(data_mem_out_wire[1519]), 
        .SEL(N37), .F(n8707) );
  MUX U8756 ( .IN0(data_mem_out_wire[1423]), .IN1(data_mem_out_wire[1455]), 
        .SEL(N37), .F(n8708) );
  MUX U8757 ( .IN0(n8708), .IN1(n8707), .SEL(N38), .F(n8709) );
  MUX U8758 ( .IN0(data_mem_out_wire[1359]), .IN1(data_mem_out_wire[1391]), 
        .SEL(N37), .F(n8710) );
  MUX U8759 ( .IN0(data_mem_out_wire[1295]), .IN1(data_mem_out_wire[1327]), 
        .SEL(N37), .F(n8711) );
  MUX U8760 ( .IN0(n8711), .IN1(n8710), .SEL(N38), .F(n8712) );
  MUX U8761 ( .IN0(n8712), .IN1(n8709), .SEL(N39), .F(n8713) );
  MUX U8762 ( .IN0(data_mem_out_wire[1231]), .IN1(data_mem_out_wire[1263]), 
        .SEL(N37), .F(n8714) );
  MUX U8763 ( .IN0(data_mem_out_wire[1167]), .IN1(data_mem_out_wire[1199]), 
        .SEL(N37), .F(n8715) );
  MUX U8764 ( .IN0(n8715), .IN1(n8714), .SEL(N38), .F(n8716) );
  MUX U8765 ( .IN0(data_mem_out_wire[1103]), .IN1(data_mem_out_wire[1135]), 
        .SEL(N37), .F(n8717) );
  MUX U8766 ( .IN0(data_mem_out_wire[1039]), .IN1(data_mem_out_wire[1071]), 
        .SEL(N37), .F(n8718) );
  MUX U8767 ( .IN0(n8718), .IN1(n8717), .SEL(N38), .F(n8719) );
  MUX U8768 ( .IN0(n8719), .IN1(n8716), .SEL(N39), .F(n8720) );
  MUX U8769 ( .IN0(n8720), .IN1(n8713), .SEL(N40), .F(n8721) );
  MUX U8770 ( .IN0(n8721), .IN1(n8706), .SEL(N41), .F(n8722) );
  MUX U8771 ( .IN0(data_mem_out_wire[975]), .IN1(data_mem_out_wire[1007]), 
        .SEL(N37), .F(n8723) );
  MUX U8772 ( .IN0(data_mem_out_wire[911]), .IN1(data_mem_out_wire[943]), 
        .SEL(N37), .F(n8724) );
  MUX U8773 ( .IN0(n8724), .IN1(n8723), .SEL(N38), .F(n8725) );
  MUX U8774 ( .IN0(data_mem_out_wire[847]), .IN1(data_mem_out_wire[879]), 
        .SEL(N37), .F(n8726) );
  MUX U8775 ( .IN0(data_mem_out_wire[783]), .IN1(data_mem_out_wire[815]), 
        .SEL(N37), .F(n8727) );
  MUX U8776 ( .IN0(n8727), .IN1(n8726), .SEL(N38), .F(n8728) );
  MUX U8777 ( .IN0(n8728), .IN1(n8725), .SEL(N39), .F(n8729) );
  MUX U8778 ( .IN0(data_mem_out_wire[719]), .IN1(data_mem_out_wire[751]), 
        .SEL(N37), .F(n8730) );
  MUX U8779 ( .IN0(data_mem_out_wire[655]), .IN1(data_mem_out_wire[687]), 
        .SEL(N37), .F(n8731) );
  MUX U8780 ( .IN0(n8731), .IN1(n8730), .SEL(N38), .F(n8732) );
  MUX U8781 ( .IN0(data_mem_out_wire[591]), .IN1(data_mem_out_wire[623]), 
        .SEL(N37), .F(n8733) );
  MUX U8782 ( .IN0(data_mem_out_wire[527]), .IN1(data_mem_out_wire[559]), 
        .SEL(N37), .F(n8734) );
  MUX U8783 ( .IN0(n8734), .IN1(n8733), .SEL(N38), .F(n8735) );
  MUX U8784 ( .IN0(n8735), .IN1(n8732), .SEL(N39), .F(n8736) );
  MUX U8785 ( .IN0(n8736), .IN1(n8729), .SEL(N40), .F(n8737) );
  MUX U8786 ( .IN0(data_mem_out_wire[463]), .IN1(data_mem_out_wire[495]), 
        .SEL(N37), .F(n8738) );
  MUX U8787 ( .IN0(data_mem_out_wire[399]), .IN1(data_mem_out_wire[431]), 
        .SEL(N37), .F(n8739) );
  MUX U8788 ( .IN0(n8739), .IN1(n8738), .SEL(N38), .F(n8740) );
  MUX U8789 ( .IN0(data_mem_out_wire[335]), .IN1(data_mem_out_wire[367]), 
        .SEL(N37), .F(n8741) );
  MUX U8790 ( .IN0(data_mem_out_wire[271]), .IN1(data_mem_out_wire[303]), 
        .SEL(N37), .F(n8742) );
  MUX U8791 ( .IN0(n8742), .IN1(n8741), .SEL(N38), .F(n8743) );
  MUX U8792 ( .IN0(n8743), .IN1(n8740), .SEL(N39), .F(n8744) );
  MUX U8793 ( .IN0(data_mem_out_wire[207]), .IN1(data_mem_out_wire[239]), 
        .SEL(N37), .F(n8745) );
  MUX U8794 ( .IN0(data_mem_out_wire[143]), .IN1(data_mem_out_wire[175]), 
        .SEL(N37), .F(n8746) );
  MUX U8795 ( .IN0(n8746), .IN1(n8745), .SEL(N38), .F(n8747) );
  MUX U8796 ( .IN0(data_mem_out_wire[79]), .IN1(data_mem_out_wire[111]), .SEL(
        N37), .F(n8748) );
  MUX U8797 ( .IN0(data_mem_out_wire[15]), .IN1(data_mem_out_wire[47]), .SEL(
        N37), .F(n8749) );
  MUX U8798 ( .IN0(n8749), .IN1(n8748), .SEL(N38), .F(n8750) );
  MUX U8799 ( .IN0(n8750), .IN1(n8747), .SEL(N39), .F(n8751) );
  MUX U8800 ( .IN0(n8751), .IN1(n8744), .SEL(N40), .F(n8752) );
  MUX U8801 ( .IN0(n8752), .IN1(n8737), .SEL(N41), .F(n8753) );
  MUX U8802 ( .IN0(n8753), .IN1(n8722), .SEL(N42), .F(N730) );
  MUX U8803 ( .IN0(data_mem_out_wire[2000]), .IN1(data_mem_out_wire[2032]), 
        .SEL(N37), .F(n8754) );
  MUX U8804 ( .IN0(data_mem_out_wire[1936]), .IN1(data_mem_out_wire[1968]), 
        .SEL(N37), .F(n8755) );
  MUX U8805 ( .IN0(n8755), .IN1(n8754), .SEL(N38), .F(n8756) );
  MUX U8806 ( .IN0(data_mem_out_wire[1872]), .IN1(data_mem_out_wire[1904]), 
        .SEL(N37), .F(n8757) );
  MUX U8807 ( .IN0(data_mem_out_wire[1808]), .IN1(data_mem_out_wire[1840]), 
        .SEL(N37), .F(n8758) );
  MUX U8808 ( .IN0(n8758), .IN1(n8757), .SEL(N38), .F(n8759) );
  MUX U8809 ( .IN0(n8759), .IN1(n8756), .SEL(N39), .F(n8760) );
  MUX U8810 ( .IN0(data_mem_out_wire[1744]), .IN1(data_mem_out_wire[1776]), 
        .SEL(N37), .F(n8761) );
  MUX U8811 ( .IN0(data_mem_out_wire[1680]), .IN1(data_mem_out_wire[1712]), 
        .SEL(N37), .F(n8762) );
  MUX U8812 ( .IN0(n8762), .IN1(n8761), .SEL(N38), .F(n8763) );
  MUX U8813 ( .IN0(data_mem_out_wire[1616]), .IN1(data_mem_out_wire[1648]), 
        .SEL(N37), .F(n8764) );
  MUX U8814 ( .IN0(data_mem_out_wire[1552]), .IN1(data_mem_out_wire[1584]), 
        .SEL(N37), .F(n8765) );
  MUX U8815 ( .IN0(n8765), .IN1(n8764), .SEL(N38), .F(n8766) );
  MUX U8816 ( .IN0(n8766), .IN1(n8763), .SEL(N39), .F(n8767) );
  MUX U8817 ( .IN0(n8767), .IN1(n8760), .SEL(N40), .F(n8768) );
  MUX U8818 ( .IN0(data_mem_out_wire[1488]), .IN1(data_mem_out_wire[1520]), 
        .SEL(N37), .F(n8769) );
  MUX U8819 ( .IN0(data_mem_out_wire[1424]), .IN1(data_mem_out_wire[1456]), 
        .SEL(N37), .F(n8770) );
  MUX U8820 ( .IN0(n8770), .IN1(n8769), .SEL(N38), .F(n8771) );
  MUX U8821 ( .IN0(data_mem_out_wire[1360]), .IN1(data_mem_out_wire[1392]), 
        .SEL(N37), .F(n8772) );
  MUX U8822 ( .IN0(data_mem_out_wire[1296]), .IN1(data_mem_out_wire[1328]), 
        .SEL(N37), .F(n8773) );
  MUX U8823 ( .IN0(n8773), .IN1(n8772), .SEL(N38), .F(n8774) );
  MUX U8824 ( .IN0(n8774), .IN1(n8771), .SEL(N39), .F(n8775) );
  MUX U8825 ( .IN0(data_mem_out_wire[1232]), .IN1(data_mem_out_wire[1264]), 
        .SEL(N37), .F(n8776) );
  MUX U8826 ( .IN0(data_mem_out_wire[1168]), .IN1(data_mem_out_wire[1200]), 
        .SEL(N37), .F(n8777) );
  MUX U8827 ( .IN0(n8777), .IN1(n8776), .SEL(N38), .F(n8778) );
  MUX U8828 ( .IN0(data_mem_out_wire[1104]), .IN1(data_mem_out_wire[1136]), 
        .SEL(N37), .F(n8779) );
  MUX U8829 ( .IN0(data_mem_out_wire[1040]), .IN1(data_mem_out_wire[1072]), 
        .SEL(N37), .F(n8780) );
  MUX U8830 ( .IN0(n8780), .IN1(n8779), .SEL(N38), .F(n8781) );
  MUX U8831 ( .IN0(n8781), .IN1(n8778), .SEL(N39), .F(n8782) );
  MUX U8832 ( .IN0(n8782), .IN1(n8775), .SEL(N40), .F(n8783) );
  MUX U8833 ( .IN0(n8783), .IN1(n8768), .SEL(N41), .F(n8784) );
  MUX U8834 ( .IN0(data_mem_out_wire[976]), .IN1(data_mem_out_wire[1008]), 
        .SEL(N37), .F(n8785) );
  MUX U8835 ( .IN0(data_mem_out_wire[912]), .IN1(data_mem_out_wire[944]), 
        .SEL(N37), .F(n8786) );
  MUX U8836 ( .IN0(n8786), .IN1(n8785), .SEL(N38), .F(n8787) );
  MUX U8837 ( .IN0(data_mem_out_wire[848]), .IN1(data_mem_out_wire[880]), 
        .SEL(N37), .F(n8788) );
  MUX U8838 ( .IN0(data_mem_out_wire[784]), .IN1(data_mem_out_wire[816]), 
        .SEL(N37), .F(n8789) );
  MUX U8839 ( .IN0(n8789), .IN1(n8788), .SEL(N38), .F(n8790) );
  MUX U8840 ( .IN0(n8790), .IN1(n8787), .SEL(N39), .F(n8791) );
  MUX U8841 ( .IN0(data_mem_out_wire[720]), .IN1(data_mem_out_wire[752]), 
        .SEL(N37), .F(n8792) );
  MUX U8842 ( .IN0(data_mem_out_wire[656]), .IN1(data_mem_out_wire[688]), 
        .SEL(N37), .F(n8793) );
  MUX U8843 ( .IN0(n8793), .IN1(n8792), .SEL(N38), .F(n8794) );
  MUX U8844 ( .IN0(data_mem_out_wire[592]), .IN1(data_mem_out_wire[624]), 
        .SEL(N37), .F(n8795) );
  MUX U8845 ( .IN0(data_mem_out_wire[528]), .IN1(data_mem_out_wire[560]), 
        .SEL(N37), .F(n8796) );
  MUX U8846 ( .IN0(n8796), .IN1(n8795), .SEL(N38), .F(n8797) );
  MUX U8847 ( .IN0(n8797), .IN1(n8794), .SEL(N39), .F(n8798) );
  MUX U8848 ( .IN0(n8798), .IN1(n8791), .SEL(N40), .F(n8799) );
  MUX U8849 ( .IN0(data_mem_out_wire[464]), .IN1(data_mem_out_wire[496]), 
        .SEL(N37), .F(n8800) );
  MUX U8850 ( .IN0(data_mem_out_wire[400]), .IN1(data_mem_out_wire[432]), 
        .SEL(N37), .F(n8801) );
  MUX U8851 ( .IN0(n8801), .IN1(n8800), .SEL(N38), .F(n8802) );
  MUX U8852 ( .IN0(data_mem_out_wire[336]), .IN1(data_mem_out_wire[368]), 
        .SEL(N37), .F(n8803) );
  MUX U8853 ( .IN0(data_mem_out_wire[272]), .IN1(data_mem_out_wire[304]), 
        .SEL(N37), .F(n8804) );
  MUX U8854 ( .IN0(n8804), .IN1(n8803), .SEL(N38), .F(n8805) );
  MUX U8855 ( .IN0(n8805), .IN1(n8802), .SEL(N39), .F(n8806) );
  MUX U8856 ( .IN0(data_mem_out_wire[208]), .IN1(data_mem_out_wire[240]), 
        .SEL(N37), .F(n8807) );
  MUX U8857 ( .IN0(data_mem_out_wire[144]), .IN1(data_mem_out_wire[176]), 
        .SEL(N37), .F(n8808) );
  MUX U8858 ( .IN0(n8808), .IN1(n8807), .SEL(N38), .F(n8809) );
  MUX U8859 ( .IN0(data_mem_out_wire[80]), .IN1(data_mem_out_wire[112]), .SEL(
        N37), .F(n8810) );
  MUX U8860 ( .IN0(data_mem_out_wire[16]), .IN1(data_mem_out_wire[48]), .SEL(
        N37), .F(n8811) );
  MUX U8861 ( .IN0(n8811), .IN1(n8810), .SEL(N38), .F(n8812) );
  MUX U8862 ( .IN0(n8812), .IN1(n8809), .SEL(N39), .F(n8813) );
  MUX U8863 ( .IN0(n8813), .IN1(n8806), .SEL(N40), .F(n8814) );
  MUX U8864 ( .IN0(n8814), .IN1(n8799), .SEL(N41), .F(n8815) );
  MUX U8865 ( .IN0(n8815), .IN1(n8784), .SEL(N42), .F(N729) );
  MUX U8866 ( .IN0(data_mem_out_wire[2001]), .IN1(data_mem_out_wire[2033]), 
        .SEL(N37), .F(n8816) );
  MUX U8867 ( .IN0(data_mem_out_wire[1937]), .IN1(data_mem_out_wire[1969]), 
        .SEL(N37), .F(n8817) );
  MUX U8868 ( .IN0(n8817), .IN1(n8816), .SEL(N38), .F(n8818) );
  MUX U8869 ( .IN0(data_mem_out_wire[1873]), .IN1(data_mem_out_wire[1905]), 
        .SEL(N37), .F(n8819) );
  MUX U8870 ( .IN0(data_mem_out_wire[1809]), .IN1(data_mem_out_wire[1841]), 
        .SEL(N37), .F(n8820) );
  MUX U8871 ( .IN0(n8820), .IN1(n8819), .SEL(N38), .F(n8821) );
  MUX U8872 ( .IN0(n8821), .IN1(n8818), .SEL(N39), .F(n8822) );
  MUX U8873 ( .IN0(data_mem_out_wire[1745]), .IN1(data_mem_out_wire[1777]), 
        .SEL(N37), .F(n8823) );
  MUX U8874 ( .IN0(data_mem_out_wire[1681]), .IN1(data_mem_out_wire[1713]), 
        .SEL(N37), .F(n8824) );
  MUX U8875 ( .IN0(n8824), .IN1(n8823), .SEL(N38), .F(n8825) );
  MUX U8876 ( .IN0(data_mem_out_wire[1617]), .IN1(data_mem_out_wire[1649]), 
        .SEL(N37), .F(n8826) );
  MUX U8877 ( .IN0(data_mem_out_wire[1553]), .IN1(data_mem_out_wire[1585]), 
        .SEL(N37), .F(n8827) );
  MUX U8878 ( .IN0(n8827), .IN1(n8826), .SEL(N38), .F(n8828) );
  MUX U8879 ( .IN0(n8828), .IN1(n8825), .SEL(N39), .F(n8829) );
  MUX U8880 ( .IN0(n8829), .IN1(n8822), .SEL(N40), .F(n8830) );
  MUX U8881 ( .IN0(data_mem_out_wire[1489]), .IN1(data_mem_out_wire[1521]), 
        .SEL(N37), .F(n8831) );
  MUX U8882 ( .IN0(data_mem_out_wire[1425]), .IN1(data_mem_out_wire[1457]), 
        .SEL(N37), .F(n8832) );
  MUX U8883 ( .IN0(n8832), .IN1(n8831), .SEL(N38), .F(n8833) );
  MUX U8884 ( .IN0(data_mem_out_wire[1361]), .IN1(data_mem_out_wire[1393]), 
        .SEL(N37), .F(n8834) );
  MUX U8885 ( .IN0(data_mem_out_wire[1297]), .IN1(data_mem_out_wire[1329]), 
        .SEL(N37), .F(n8835) );
  MUX U8886 ( .IN0(n8835), .IN1(n8834), .SEL(N38), .F(n8836) );
  MUX U8887 ( .IN0(n8836), .IN1(n8833), .SEL(N39), .F(n8837) );
  MUX U8888 ( .IN0(data_mem_out_wire[1233]), .IN1(data_mem_out_wire[1265]), 
        .SEL(N37), .F(n8838) );
  MUX U8889 ( .IN0(data_mem_out_wire[1169]), .IN1(data_mem_out_wire[1201]), 
        .SEL(N37), .F(n8839) );
  MUX U8890 ( .IN0(n8839), .IN1(n8838), .SEL(N38), .F(n8840) );
  MUX U8891 ( .IN0(data_mem_out_wire[1105]), .IN1(data_mem_out_wire[1137]), 
        .SEL(N37), .F(n8841) );
  MUX U8892 ( .IN0(data_mem_out_wire[1041]), .IN1(data_mem_out_wire[1073]), 
        .SEL(N37), .F(n8842) );
  MUX U8893 ( .IN0(n8842), .IN1(n8841), .SEL(N38), .F(n8843) );
  MUX U8894 ( .IN0(n8843), .IN1(n8840), .SEL(N39), .F(n8844) );
  MUX U8895 ( .IN0(n8844), .IN1(n8837), .SEL(N40), .F(n8845) );
  MUX U8896 ( .IN0(n8845), .IN1(n8830), .SEL(N41), .F(n8846) );
  MUX U8897 ( .IN0(data_mem_out_wire[977]), .IN1(data_mem_out_wire[1009]), 
        .SEL(N37), .F(n8847) );
  MUX U8898 ( .IN0(data_mem_out_wire[913]), .IN1(data_mem_out_wire[945]), 
        .SEL(N37), .F(n8848) );
  MUX U8899 ( .IN0(n8848), .IN1(n8847), .SEL(N38), .F(n8849) );
  MUX U8900 ( .IN0(data_mem_out_wire[849]), .IN1(data_mem_out_wire[881]), 
        .SEL(N37), .F(n8850) );
  MUX U8901 ( .IN0(data_mem_out_wire[785]), .IN1(data_mem_out_wire[817]), 
        .SEL(N37), .F(n8851) );
  MUX U8902 ( .IN0(n8851), .IN1(n8850), .SEL(N38), .F(n8852) );
  MUX U8903 ( .IN0(n8852), .IN1(n8849), .SEL(N39), .F(n8853) );
  MUX U8904 ( .IN0(data_mem_out_wire[721]), .IN1(data_mem_out_wire[753]), 
        .SEL(N37), .F(n8854) );
  MUX U8905 ( .IN0(data_mem_out_wire[657]), .IN1(data_mem_out_wire[689]), 
        .SEL(N37), .F(n8855) );
  MUX U8906 ( .IN0(n8855), .IN1(n8854), .SEL(N38), .F(n8856) );
  MUX U8907 ( .IN0(data_mem_out_wire[593]), .IN1(data_mem_out_wire[625]), 
        .SEL(N37), .F(n8857) );
  MUX U8908 ( .IN0(data_mem_out_wire[529]), .IN1(data_mem_out_wire[561]), 
        .SEL(N37), .F(n8858) );
  MUX U8909 ( .IN0(n8858), .IN1(n8857), .SEL(N38), .F(n8859) );
  MUX U8910 ( .IN0(n8859), .IN1(n8856), .SEL(N39), .F(n8860) );
  MUX U8911 ( .IN0(n8860), .IN1(n8853), .SEL(N40), .F(n8861) );
  MUX U8912 ( .IN0(data_mem_out_wire[465]), .IN1(data_mem_out_wire[497]), 
        .SEL(N37), .F(n8862) );
  MUX U8913 ( .IN0(data_mem_out_wire[401]), .IN1(data_mem_out_wire[433]), 
        .SEL(N37), .F(n8863) );
  MUX U8914 ( .IN0(n8863), .IN1(n8862), .SEL(N38), .F(n8864) );
  MUX U8915 ( .IN0(data_mem_out_wire[337]), .IN1(data_mem_out_wire[369]), 
        .SEL(N37), .F(n8865) );
  MUX U8916 ( .IN0(data_mem_out_wire[273]), .IN1(data_mem_out_wire[305]), 
        .SEL(N37), .F(n8866) );
  MUX U8917 ( .IN0(n8866), .IN1(n8865), .SEL(N38), .F(n8867) );
  MUX U8918 ( .IN0(n8867), .IN1(n8864), .SEL(N39), .F(n8868) );
  MUX U8919 ( .IN0(data_mem_out_wire[209]), .IN1(data_mem_out_wire[241]), 
        .SEL(N37), .F(n8869) );
  MUX U8920 ( .IN0(data_mem_out_wire[145]), .IN1(data_mem_out_wire[177]), 
        .SEL(N37), .F(n8870) );
  MUX U8921 ( .IN0(n8870), .IN1(n8869), .SEL(N38), .F(n8871) );
  MUX U8922 ( .IN0(data_mem_out_wire[81]), .IN1(data_mem_out_wire[113]), .SEL(
        N37), .F(n8872) );
  MUX U8923 ( .IN0(data_mem_out_wire[17]), .IN1(data_mem_out_wire[49]), .SEL(
        N37), .F(n8873) );
  MUX U8924 ( .IN0(n8873), .IN1(n8872), .SEL(N38), .F(n8874) );
  MUX U8925 ( .IN0(n8874), .IN1(n8871), .SEL(N39), .F(n8875) );
  MUX U8926 ( .IN0(n8875), .IN1(n8868), .SEL(N40), .F(n8876) );
  MUX U8927 ( .IN0(n8876), .IN1(n8861), .SEL(N41), .F(n8877) );
  MUX U8928 ( .IN0(n8877), .IN1(n8846), .SEL(N42), .F(N728) );
  MUX U8929 ( .IN0(data_mem_out_wire[2002]), .IN1(data_mem_out_wire[2034]), 
        .SEL(N37), .F(n8878) );
  MUX U8930 ( .IN0(data_mem_out_wire[1938]), .IN1(data_mem_out_wire[1970]), 
        .SEL(N37), .F(n8879) );
  MUX U8931 ( .IN0(n8879), .IN1(n8878), .SEL(N38), .F(n8880) );
  MUX U8932 ( .IN0(data_mem_out_wire[1874]), .IN1(data_mem_out_wire[1906]), 
        .SEL(N37), .F(n8881) );
  MUX U8933 ( .IN0(data_mem_out_wire[1810]), .IN1(data_mem_out_wire[1842]), 
        .SEL(N37), .F(n8882) );
  MUX U8934 ( .IN0(n8882), .IN1(n8881), .SEL(N38), .F(n8883) );
  MUX U8935 ( .IN0(n8883), .IN1(n8880), .SEL(N39), .F(n8884) );
  MUX U8936 ( .IN0(data_mem_out_wire[1746]), .IN1(data_mem_out_wire[1778]), 
        .SEL(N37), .F(n8885) );
  MUX U8937 ( .IN0(data_mem_out_wire[1682]), .IN1(data_mem_out_wire[1714]), 
        .SEL(N37), .F(n8886) );
  MUX U8938 ( .IN0(n8886), .IN1(n8885), .SEL(N38), .F(n8887) );
  MUX U8939 ( .IN0(data_mem_out_wire[1618]), .IN1(data_mem_out_wire[1650]), 
        .SEL(N37), .F(n8888) );
  MUX U8940 ( .IN0(data_mem_out_wire[1554]), .IN1(data_mem_out_wire[1586]), 
        .SEL(N37), .F(n8889) );
  MUX U8941 ( .IN0(n8889), .IN1(n8888), .SEL(N38), .F(n8890) );
  MUX U8942 ( .IN0(n8890), .IN1(n8887), .SEL(N39), .F(n8891) );
  MUX U8943 ( .IN0(n8891), .IN1(n8884), .SEL(N40), .F(n8892) );
  MUX U8944 ( .IN0(data_mem_out_wire[1490]), .IN1(data_mem_out_wire[1522]), 
        .SEL(N37), .F(n8893) );
  MUX U8945 ( .IN0(data_mem_out_wire[1426]), .IN1(data_mem_out_wire[1458]), 
        .SEL(N37), .F(n8894) );
  MUX U8946 ( .IN0(n8894), .IN1(n8893), .SEL(N38), .F(n8895) );
  MUX U8947 ( .IN0(data_mem_out_wire[1362]), .IN1(data_mem_out_wire[1394]), 
        .SEL(N37), .F(n8896) );
  MUX U8948 ( .IN0(data_mem_out_wire[1298]), .IN1(data_mem_out_wire[1330]), 
        .SEL(N37), .F(n8897) );
  MUX U8949 ( .IN0(n8897), .IN1(n8896), .SEL(N38), .F(n8898) );
  MUX U8950 ( .IN0(n8898), .IN1(n8895), .SEL(N39), .F(n8899) );
  MUX U8951 ( .IN0(data_mem_out_wire[1234]), .IN1(data_mem_out_wire[1266]), 
        .SEL(N37), .F(n8900) );
  MUX U8952 ( .IN0(data_mem_out_wire[1170]), .IN1(data_mem_out_wire[1202]), 
        .SEL(N37), .F(n8901) );
  MUX U8953 ( .IN0(n8901), .IN1(n8900), .SEL(N38), .F(n8902) );
  MUX U8954 ( .IN0(data_mem_out_wire[1106]), .IN1(data_mem_out_wire[1138]), 
        .SEL(N37), .F(n8903) );
  MUX U8955 ( .IN0(data_mem_out_wire[1042]), .IN1(data_mem_out_wire[1074]), 
        .SEL(N37), .F(n8904) );
  MUX U8956 ( .IN0(n8904), .IN1(n8903), .SEL(N38), .F(n8905) );
  MUX U8957 ( .IN0(n8905), .IN1(n8902), .SEL(N39), .F(n8906) );
  MUX U8958 ( .IN0(n8906), .IN1(n8899), .SEL(N40), .F(n8907) );
  MUX U8959 ( .IN0(n8907), .IN1(n8892), .SEL(N41), .F(n8908) );
  MUX U8960 ( .IN0(data_mem_out_wire[978]), .IN1(data_mem_out_wire[1010]), 
        .SEL(N37), .F(n8909) );
  MUX U8961 ( .IN0(data_mem_out_wire[914]), .IN1(data_mem_out_wire[946]), 
        .SEL(N37), .F(n8910) );
  MUX U8962 ( .IN0(n8910), .IN1(n8909), .SEL(N38), .F(n8911) );
  MUX U8963 ( .IN0(data_mem_out_wire[850]), .IN1(data_mem_out_wire[882]), 
        .SEL(N37), .F(n8912) );
  MUX U8964 ( .IN0(data_mem_out_wire[786]), .IN1(data_mem_out_wire[818]), 
        .SEL(N37), .F(n8913) );
  MUX U8965 ( .IN0(n8913), .IN1(n8912), .SEL(N38), .F(n8914) );
  MUX U8966 ( .IN0(n8914), .IN1(n8911), .SEL(N39), .F(n8915) );
  MUX U8967 ( .IN0(data_mem_out_wire[722]), .IN1(data_mem_out_wire[754]), 
        .SEL(N37), .F(n8916) );
  MUX U8968 ( .IN0(data_mem_out_wire[658]), .IN1(data_mem_out_wire[690]), 
        .SEL(N37), .F(n8917) );
  MUX U8969 ( .IN0(n8917), .IN1(n8916), .SEL(N38), .F(n8918) );
  MUX U8970 ( .IN0(data_mem_out_wire[594]), .IN1(data_mem_out_wire[626]), 
        .SEL(N37), .F(n8919) );
  MUX U8971 ( .IN0(data_mem_out_wire[530]), .IN1(data_mem_out_wire[562]), 
        .SEL(N37), .F(n8920) );
  MUX U8972 ( .IN0(n8920), .IN1(n8919), .SEL(N38), .F(n8921) );
  MUX U8973 ( .IN0(n8921), .IN1(n8918), .SEL(N39), .F(n8922) );
  MUX U8974 ( .IN0(n8922), .IN1(n8915), .SEL(N40), .F(n8923) );
  MUX U8975 ( .IN0(data_mem_out_wire[466]), .IN1(data_mem_out_wire[498]), 
        .SEL(N37), .F(n8924) );
  MUX U8976 ( .IN0(data_mem_out_wire[402]), .IN1(data_mem_out_wire[434]), 
        .SEL(N37), .F(n8925) );
  MUX U8977 ( .IN0(n8925), .IN1(n8924), .SEL(N38), .F(n8926) );
  MUX U8978 ( .IN0(data_mem_out_wire[338]), .IN1(data_mem_out_wire[370]), 
        .SEL(N37), .F(n8927) );
  MUX U8979 ( .IN0(data_mem_out_wire[274]), .IN1(data_mem_out_wire[306]), 
        .SEL(N37), .F(n8928) );
  MUX U8980 ( .IN0(n8928), .IN1(n8927), .SEL(N38), .F(n8929) );
  MUX U8981 ( .IN0(n8929), .IN1(n8926), .SEL(N39), .F(n8930) );
  MUX U8982 ( .IN0(data_mem_out_wire[210]), .IN1(data_mem_out_wire[242]), 
        .SEL(N37), .F(n8931) );
  MUX U8983 ( .IN0(data_mem_out_wire[146]), .IN1(data_mem_out_wire[178]), 
        .SEL(N37), .F(n8932) );
  MUX U8984 ( .IN0(n8932), .IN1(n8931), .SEL(N38), .F(n8933) );
  MUX U8985 ( .IN0(data_mem_out_wire[82]), .IN1(data_mem_out_wire[114]), .SEL(
        N37), .F(n8934) );
  MUX U8986 ( .IN0(data_mem_out_wire[18]), .IN1(data_mem_out_wire[50]), .SEL(
        N37), .F(n8935) );
  MUX U8987 ( .IN0(n8935), .IN1(n8934), .SEL(N38), .F(n8936) );
  MUX U8988 ( .IN0(n8936), .IN1(n8933), .SEL(N39), .F(n8937) );
  MUX U8989 ( .IN0(n8937), .IN1(n8930), .SEL(N40), .F(n8938) );
  MUX U8990 ( .IN0(n8938), .IN1(n8923), .SEL(N41), .F(n8939) );
  MUX U8991 ( .IN0(n8939), .IN1(n8908), .SEL(N42), .F(N727) );
  MUX U8992 ( .IN0(data_mem_out_wire[2003]), .IN1(data_mem_out_wire[2035]), 
        .SEL(N37), .F(n8940) );
  MUX U8993 ( .IN0(data_mem_out_wire[1939]), .IN1(data_mem_out_wire[1971]), 
        .SEL(N37), .F(n8941) );
  MUX U8994 ( .IN0(n8941), .IN1(n8940), .SEL(N38), .F(n8942) );
  MUX U8995 ( .IN0(data_mem_out_wire[1875]), .IN1(data_mem_out_wire[1907]), 
        .SEL(N37), .F(n8943) );
  MUX U8996 ( .IN0(data_mem_out_wire[1811]), .IN1(data_mem_out_wire[1843]), 
        .SEL(N37), .F(n8944) );
  MUX U8997 ( .IN0(n8944), .IN1(n8943), .SEL(N38), .F(n8945) );
  MUX U8998 ( .IN0(n8945), .IN1(n8942), .SEL(N39), .F(n8946) );
  MUX U8999 ( .IN0(data_mem_out_wire[1747]), .IN1(data_mem_out_wire[1779]), 
        .SEL(N37), .F(n8947) );
  MUX U9000 ( .IN0(data_mem_out_wire[1683]), .IN1(data_mem_out_wire[1715]), 
        .SEL(N37), .F(n8948) );
  MUX U9001 ( .IN0(n8948), .IN1(n8947), .SEL(N38), .F(n8949) );
  MUX U9002 ( .IN0(data_mem_out_wire[1619]), .IN1(data_mem_out_wire[1651]), 
        .SEL(N37), .F(n8950) );
  MUX U9003 ( .IN0(data_mem_out_wire[1555]), .IN1(data_mem_out_wire[1587]), 
        .SEL(N37), .F(n8951) );
  MUX U9004 ( .IN0(n8951), .IN1(n8950), .SEL(N38), .F(n8952) );
  MUX U9005 ( .IN0(n8952), .IN1(n8949), .SEL(N39), .F(n8953) );
  MUX U9006 ( .IN0(n8953), .IN1(n8946), .SEL(N40), .F(n8954) );
  MUX U9007 ( .IN0(data_mem_out_wire[1491]), .IN1(data_mem_out_wire[1523]), 
        .SEL(N37), .F(n8955) );
  MUX U9008 ( .IN0(data_mem_out_wire[1427]), .IN1(data_mem_out_wire[1459]), 
        .SEL(N37), .F(n8956) );
  MUX U9009 ( .IN0(n8956), .IN1(n8955), .SEL(N38), .F(n8957) );
  MUX U9010 ( .IN0(data_mem_out_wire[1363]), .IN1(data_mem_out_wire[1395]), 
        .SEL(N37), .F(n8958) );
  MUX U9011 ( .IN0(data_mem_out_wire[1299]), .IN1(data_mem_out_wire[1331]), 
        .SEL(N37), .F(n8959) );
  MUX U9012 ( .IN0(n8959), .IN1(n8958), .SEL(N38), .F(n8960) );
  MUX U9013 ( .IN0(n8960), .IN1(n8957), .SEL(N39), .F(n8961) );
  MUX U9014 ( .IN0(data_mem_out_wire[1235]), .IN1(data_mem_out_wire[1267]), 
        .SEL(N37), .F(n8962) );
  MUX U9015 ( .IN0(data_mem_out_wire[1171]), .IN1(data_mem_out_wire[1203]), 
        .SEL(N37), .F(n8963) );
  MUX U9016 ( .IN0(n8963), .IN1(n8962), .SEL(N38), .F(n8964) );
  MUX U9017 ( .IN0(data_mem_out_wire[1107]), .IN1(data_mem_out_wire[1139]), 
        .SEL(N37), .F(n8965) );
  MUX U9018 ( .IN0(data_mem_out_wire[1043]), .IN1(data_mem_out_wire[1075]), 
        .SEL(N37), .F(n8966) );
  MUX U9019 ( .IN0(n8966), .IN1(n8965), .SEL(N38), .F(n8967) );
  MUX U9020 ( .IN0(n8967), .IN1(n8964), .SEL(N39), .F(n8968) );
  MUX U9021 ( .IN0(n8968), .IN1(n8961), .SEL(N40), .F(n8969) );
  MUX U9022 ( .IN0(n8969), .IN1(n8954), .SEL(N41), .F(n8970) );
  MUX U9023 ( .IN0(data_mem_out_wire[979]), .IN1(data_mem_out_wire[1011]), 
        .SEL(N37), .F(n8971) );
  MUX U9024 ( .IN0(data_mem_out_wire[915]), .IN1(data_mem_out_wire[947]), 
        .SEL(N37), .F(n8972) );
  MUX U9025 ( .IN0(n8972), .IN1(n8971), .SEL(N38), .F(n8973) );
  MUX U9026 ( .IN0(data_mem_out_wire[851]), .IN1(data_mem_out_wire[883]), 
        .SEL(N37), .F(n8974) );
  MUX U9027 ( .IN0(data_mem_out_wire[787]), .IN1(data_mem_out_wire[819]), 
        .SEL(N37), .F(n8975) );
  MUX U9028 ( .IN0(n8975), .IN1(n8974), .SEL(N38), .F(n8976) );
  MUX U9029 ( .IN0(n8976), .IN1(n8973), .SEL(N39), .F(n8977) );
  MUX U9030 ( .IN0(data_mem_out_wire[723]), .IN1(data_mem_out_wire[755]), 
        .SEL(N37), .F(n8978) );
  MUX U9031 ( .IN0(data_mem_out_wire[659]), .IN1(data_mem_out_wire[691]), 
        .SEL(N37), .F(n8979) );
  MUX U9032 ( .IN0(n8979), .IN1(n8978), .SEL(N38), .F(n8980) );
  MUX U9033 ( .IN0(data_mem_out_wire[595]), .IN1(data_mem_out_wire[627]), 
        .SEL(N37), .F(n8981) );
  MUX U9034 ( .IN0(data_mem_out_wire[531]), .IN1(data_mem_out_wire[563]), 
        .SEL(N37), .F(n8982) );
  MUX U9035 ( .IN0(n8982), .IN1(n8981), .SEL(N38), .F(n8983) );
  MUX U9036 ( .IN0(n8983), .IN1(n8980), .SEL(N39), .F(n8984) );
  MUX U9037 ( .IN0(n8984), .IN1(n8977), .SEL(N40), .F(n8985) );
  MUX U9038 ( .IN0(data_mem_out_wire[467]), .IN1(data_mem_out_wire[499]), 
        .SEL(N37), .F(n8986) );
  MUX U9039 ( .IN0(data_mem_out_wire[403]), .IN1(data_mem_out_wire[435]), 
        .SEL(N37), .F(n8987) );
  MUX U9040 ( .IN0(n8987), .IN1(n8986), .SEL(N38), .F(n8988) );
  MUX U9041 ( .IN0(data_mem_out_wire[339]), .IN1(data_mem_out_wire[371]), 
        .SEL(N37), .F(n8989) );
  MUX U9042 ( .IN0(data_mem_out_wire[275]), .IN1(data_mem_out_wire[307]), 
        .SEL(N37), .F(n8990) );
  MUX U9043 ( .IN0(n8990), .IN1(n8989), .SEL(N38), .F(n8991) );
  MUX U9044 ( .IN0(n8991), .IN1(n8988), .SEL(N39), .F(n8992) );
  MUX U9045 ( .IN0(data_mem_out_wire[211]), .IN1(data_mem_out_wire[243]), 
        .SEL(N37), .F(n8993) );
  MUX U9046 ( .IN0(data_mem_out_wire[147]), .IN1(data_mem_out_wire[179]), 
        .SEL(N37), .F(n8994) );
  MUX U9047 ( .IN0(n8994), .IN1(n8993), .SEL(N38), .F(n8995) );
  MUX U9048 ( .IN0(data_mem_out_wire[83]), .IN1(data_mem_out_wire[115]), .SEL(
        N37), .F(n8996) );
  MUX U9049 ( .IN0(data_mem_out_wire[19]), .IN1(data_mem_out_wire[51]), .SEL(
        N37), .F(n8997) );
  MUX U9050 ( .IN0(n8997), .IN1(n8996), .SEL(N38), .F(n8998) );
  MUX U9051 ( .IN0(n8998), .IN1(n8995), .SEL(N39), .F(n8999) );
  MUX U9052 ( .IN0(n8999), .IN1(n8992), .SEL(N40), .F(n9000) );
  MUX U9053 ( .IN0(n9000), .IN1(n8985), .SEL(N41), .F(n9001) );
  MUX U9054 ( .IN0(n9001), .IN1(n8970), .SEL(N42), .F(N726) );
  MUX U9055 ( .IN0(data_mem_out_wire[2004]), .IN1(data_mem_out_wire[2036]), 
        .SEL(N37), .F(n9002) );
  MUX U9056 ( .IN0(data_mem_out_wire[1940]), .IN1(data_mem_out_wire[1972]), 
        .SEL(N37), .F(n9003) );
  MUX U9057 ( .IN0(n9003), .IN1(n9002), .SEL(N38), .F(n9004) );
  MUX U9058 ( .IN0(data_mem_out_wire[1876]), .IN1(data_mem_out_wire[1908]), 
        .SEL(N37), .F(n9005) );
  MUX U9059 ( .IN0(data_mem_out_wire[1812]), .IN1(data_mem_out_wire[1844]), 
        .SEL(N37), .F(n9006) );
  MUX U9060 ( .IN0(n9006), .IN1(n9005), .SEL(N38), .F(n9007) );
  MUX U9061 ( .IN0(n9007), .IN1(n9004), .SEL(N39), .F(n9008) );
  MUX U9062 ( .IN0(data_mem_out_wire[1748]), .IN1(data_mem_out_wire[1780]), 
        .SEL(N37), .F(n9009) );
  MUX U9063 ( .IN0(data_mem_out_wire[1684]), .IN1(data_mem_out_wire[1716]), 
        .SEL(N37), .F(n9010) );
  MUX U9064 ( .IN0(n9010), .IN1(n9009), .SEL(N38), .F(n9011) );
  MUX U9065 ( .IN0(data_mem_out_wire[1620]), .IN1(data_mem_out_wire[1652]), 
        .SEL(N37), .F(n9012) );
  MUX U9066 ( .IN0(data_mem_out_wire[1556]), .IN1(data_mem_out_wire[1588]), 
        .SEL(N37), .F(n9013) );
  MUX U9067 ( .IN0(n9013), .IN1(n9012), .SEL(N38), .F(n9014) );
  MUX U9068 ( .IN0(n9014), .IN1(n9011), .SEL(N39), .F(n9015) );
  MUX U9069 ( .IN0(n9015), .IN1(n9008), .SEL(N40), .F(n9016) );
  MUX U9070 ( .IN0(data_mem_out_wire[1492]), .IN1(data_mem_out_wire[1524]), 
        .SEL(N37), .F(n9017) );
  MUX U9071 ( .IN0(data_mem_out_wire[1428]), .IN1(data_mem_out_wire[1460]), 
        .SEL(N37), .F(n9018) );
  MUX U9072 ( .IN0(n9018), .IN1(n9017), .SEL(N38), .F(n9019) );
  MUX U9073 ( .IN0(data_mem_out_wire[1364]), .IN1(data_mem_out_wire[1396]), 
        .SEL(N37), .F(n9020) );
  MUX U9074 ( .IN0(data_mem_out_wire[1300]), .IN1(data_mem_out_wire[1332]), 
        .SEL(N37), .F(n9021) );
  MUX U9075 ( .IN0(n9021), .IN1(n9020), .SEL(N38), .F(n9022) );
  MUX U9076 ( .IN0(n9022), .IN1(n9019), .SEL(N39), .F(n9023) );
  MUX U9077 ( .IN0(data_mem_out_wire[1236]), .IN1(data_mem_out_wire[1268]), 
        .SEL(N37), .F(n9024) );
  MUX U9078 ( .IN0(data_mem_out_wire[1172]), .IN1(data_mem_out_wire[1204]), 
        .SEL(N37), .F(n9025) );
  MUX U9079 ( .IN0(n9025), .IN1(n9024), .SEL(N38), .F(n9026) );
  MUX U9080 ( .IN0(data_mem_out_wire[1108]), .IN1(data_mem_out_wire[1140]), 
        .SEL(N37), .F(n9027) );
  MUX U9081 ( .IN0(data_mem_out_wire[1044]), .IN1(data_mem_out_wire[1076]), 
        .SEL(N37), .F(n9028) );
  MUX U9082 ( .IN0(n9028), .IN1(n9027), .SEL(N38), .F(n9029) );
  MUX U9083 ( .IN0(n9029), .IN1(n9026), .SEL(N39), .F(n9030) );
  MUX U9084 ( .IN0(n9030), .IN1(n9023), .SEL(N40), .F(n9031) );
  MUX U9085 ( .IN0(n9031), .IN1(n9016), .SEL(N41), .F(n9032) );
  MUX U9086 ( .IN0(data_mem_out_wire[980]), .IN1(data_mem_out_wire[1012]), 
        .SEL(N37), .F(n9033) );
  MUX U9087 ( .IN0(data_mem_out_wire[916]), .IN1(data_mem_out_wire[948]), 
        .SEL(N37), .F(n9034) );
  MUX U9088 ( .IN0(n9034), .IN1(n9033), .SEL(N38), .F(n9035) );
  MUX U9089 ( .IN0(data_mem_out_wire[852]), .IN1(data_mem_out_wire[884]), 
        .SEL(N37), .F(n9036) );
  MUX U9090 ( .IN0(data_mem_out_wire[788]), .IN1(data_mem_out_wire[820]), 
        .SEL(N37), .F(n9037) );
  MUX U9091 ( .IN0(n9037), .IN1(n9036), .SEL(N38), .F(n9038) );
  MUX U9092 ( .IN0(n9038), .IN1(n9035), .SEL(N39), .F(n9039) );
  MUX U9093 ( .IN0(data_mem_out_wire[724]), .IN1(data_mem_out_wire[756]), 
        .SEL(N37), .F(n9040) );
  MUX U9094 ( .IN0(data_mem_out_wire[660]), .IN1(data_mem_out_wire[692]), 
        .SEL(N37), .F(n9041) );
  MUX U9095 ( .IN0(n9041), .IN1(n9040), .SEL(N38), .F(n9042) );
  MUX U9096 ( .IN0(data_mem_out_wire[596]), .IN1(data_mem_out_wire[628]), 
        .SEL(N37), .F(n9043) );
  MUX U9097 ( .IN0(data_mem_out_wire[532]), .IN1(data_mem_out_wire[564]), 
        .SEL(N37), .F(n9044) );
  MUX U9098 ( .IN0(n9044), .IN1(n9043), .SEL(N38), .F(n9045) );
  MUX U9099 ( .IN0(n9045), .IN1(n9042), .SEL(N39), .F(n9046) );
  MUX U9100 ( .IN0(n9046), .IN1(n9039), .SEL(N40), .F(n9047) );
  MUX U9101 ( .IN0(data_mem_out_wire[468]), .IN1(data_mem_out_wire[500]), 
        .SEL(N37), .F(n9048) );
  MUX U9102 ( .IN0(data_mem_out_wire[404]), .IN1(data_mem_out_wire[436]), 
        .SEL(N37), .F(n9049) );
  MUX U9103 ( .IN0(n9049), .IN1(n9048), .SEL(N38), .F(n9050) );
  MUX U9104 ( .IN0(data_mem_out_wire[340]), .IN1(data_mem_out_wire[372]), 
        .SEL(N37), .F(n9051) );
  MUX U9105 ( .IN0(data_mem_out_wire[276]), .IN1(data_mem_out_wire[308]), 
        .SEL(N37), .F(n9052) );
  MUX U9106 ( .IN0(n9052), .IN1(n9051), .SEL(N38), .F(n9053) );
  MUX U9107 ( .IN0(n9053), .IN1(n9050), .SEL(N39), .F(n9054) );
  MUX U9108 ( .IN0(data_mem_out_wire[212]), .IN1(data_mem_out_wire[244]), 
        .SEL(N37), .F(n9055) );
  MUX U9109 ( .IN0(data_mem_out_wire[148]), .IN1(data_mem_out_wire[180]), 
        .SEL(N37), .F(n9056) );
  MUX U9110 ( .IN0(n9056), .IN1(n9055), .SEL(N38), .F(n9057) );
  MUX U9111 ( .IN0(data_mem_out_wire[84]), .IN1(data_mem_out_wire[116]), .SEL(
        N37), .F(n9058) );
  MUX U9112 ( .IN0(data_mem_out_wire[20]), .IN1(data_mem_out_wire[52]), .SEL(
        N37), .F(n9059) );
  MUX U9113 ( .IN0(n9059), .IN1(n9058), .SEL(N38), .F(n9060) );
  MUX U9114 ( .IN0(n9060), .IN1(n9057), .SEL(N39), .F(n9061) );
  MUX U9115 ( .IN0(n9061), .IN1(n9054), .SEL(N40), .F(n9062) );
  MUX U9116 ( .IN0(n9062), .IN1(n9047), .SEL(N41), .F(n9063) );
  MUX U9117 ( .IN0(n9063), .IN1(n9032), .SEL(N42), .F(N725) );
  MUX U9118 ( .IN0(data_mem_out_wire[2005]), .IN1(data_mem_out_wire[2037]), 
        .SEL(N37), .F(n9064) );
  MUX U9119 ( .IN0(data_mem_out_wire[1941]), .IN1(data_mem_out_wire[1973]), 
        .SEL(N37), .F(n9065) );
  MUX U9120 ( .IN0(n9065), .IN1(n9064), .SEL(N38), .F(n9066) );
  MUX U9121 ( .IN0(data_mem_out_wire[1877]), .IN1(data_mem_out_wire[1909]), 
        .SEL(N37), .F(n9067) );
  MUX U9122 ( .IN0(data_mem_out_wire[1813]), .IN1(data_mem_out_wire[1845]), 
        .SEL(N37), .F(n9068) );
  MUX U9123 ( .IN0(n9068), .IN1(n9067), .SEL(N38), .F(n9069) );
  MUX U9124 ( .IN0(n9069), .IN1(n9066), .SEL(N39), .F(n9070) );
  MUX U9125 ( .IN0(data_mem_out_wire[1749]), .IN1(data_mem_out_wire[1781]), 
        .SEL(N37), .F(n9071) );
  MUX U9126 ( .IN0(data_mem_out_wire[1685]), .IN1(data_mem_out_wire[1717]), 
        .SEL(N37), .F(n9072) );
  MUX U9127 ( .IN0(n9072), .IN1(n9071), .SEL(N38), .F(n9073) );
  MUX U9128 ( .IN0(data_mem_out_wire[1621]), .IN1(data_mem_out_wire[1653]), 
        .SEL(N37), .F(n9074) );
  MUX U9129 ( .IN0(data_mem_out_wire[1557]), .IN1(data_mem_out_wire[1589]), 
        .SEL(N37), .F(n9075) );
  MUX U9130 ( .IN0(n9075), .IN1(n9074), .SEL(N38), .F(n9076) );
  MUX U9131 ( .IN0(n9076), .IN1(n9073), .SEL(N39), .F(n9077) );
  MUX U9132 ( .IN0(n9077), .IN1(n9070), .SEL(N40), .F(n9078) );
  MUX U9133 ( .IN0(data_mem_out_wire[1493]), .IN1(data_mem_out_wire[1525]), 
        .SEL(N37), .F(n9079) );
  MUX U9134 ( .IN0(data_mem_out_wire[1429]), .IN1(data_mem_out_wire[1461]), 
        .SEL(N37), .F(n9080) );
  MUX U9135 ( .IN0(n9080), .IN1(n9079), .SEL(N38), .F(n9081) );
  MUX U9136 ( .IN0(data_mem_out_wire[1365]), .IN1(data_mem_out_wire[1397]), 
        .SEL(N37), .F(n9082) );
  MUX U9137 ( .IN0(data_mem_out_wire[1301]), .IN1(data_mem_out_wire[1333]), 
        .SEL(N37), .F(n9083) );
  MUX U9138 ( .IN0(n9083), .IN1(n9082), .SEL(N38), .F(n9084) );
  MUX U9139 ( .IN0(n9084), .IN1(n9081), .SEL(N39), .F(n9085) );
  MUX U9140 ( .IN0(data_mem_out_wire[1237]), .IN1(data_mem_out_wire[1269]), 
        .SEL(N37), .F(n9086) );
  MUX U9141 ( .IN0(data_mem_out_wire[1173]), .IN1(data_mem_out_wire[1205]), 
        .SEL(N37), .F(n9087) );
  MUX U9142 ( .IN0(n9087), .IN1(n9086), .SEL(N38), .F(n9088) );
  MUX U9143 ( .IN0(data_mem_out_wire[1109]), .IN1(data_mem_out_wire[1141]), 
        .SEL(N37), .F(n9089) );
  MUX U9144 ( .IN0(data_mem_out_wire[1045]), .IN1(data_mem_out_wire[1077]), 
        .SEL(N37), .F(n9090) );
  MUX U9145 ( .IN0(n9090), .IN1(n9089), .SEL(N38), .F(n9091) );
  MUX U9146 ( .IN0(n9091), .IN1(n9088), .SEL(N39), .F(n9092) );
  MUX U9147 ( .IN0(n9092), .IN1(n9085), .SEL(N40), .F(n9093) );
  MUX U9148 ( .IN0(n9093), .IN1(n9078), .SEL(N41), .F(n9094) );
  MUX U9149 ( .IN0(data_mem_out_wire[981]), .IN1(data_mem_out_wire[1013]), 
        .SEL(N37), .F(n9095) );
  MUX U9150 ( .IN0(data_mem_out_wire[917]), .IN1(data_mem_out_wire[949]), 
        .SEL(N37), .F(n9096) );
  MUX U9151 ( .IN0(n9096), .IN1(n9095), .SEL(N38), .F(n9097) );
  MUX U9152 ( .IN0(data_mem_out_wire[853]), .IN1(data_mem_out_wire[885]), 
        .SEL(N37), .F(n9098) );
  MUX U9153 ( .IN0(data_mem_out_wire[789]), .IN1(data_mem_out_wire[821]), 
        .SEL(N37), .F(n9099) );
  MUX U9154 ( .IN0(n9099), .IN1(n9098), .SEL(N38), .F(n9100) );
  MUX U9155 ( .IN0(n9100), .IN1(n9097), .SEL(N39), .F(n9101) );
  MUX U9156 ( .IN0(data_mem_out_wire[725]), .IN1(data_mem_out_wire[757]), 
        .SEL(N37), .F(n9102) );
  MUX U9157 ( .IN0(data_mem_out_wire[661]), .IN1(data_mem_out_wire[693]), 
        .SEL(N37), .F(n9103) );
  MUX U9158 ( .IN0(n9103), .IN1(n9102), .SEL(N38), .F(n9104) );
  MUX U9159 ( .IN0(data_mem_out_wire[597]), .IN1(data_mem_out_wire[629]), 
        .SEL(N37), .F(n9105) );
  MUX U9160 ( .IN0(data_mem_out_wire[533]), .IN1(data_mem_out_wire[565]), 
        .SEL(N37), .F(n9106) );
  MUX U9161 ( .IN0(n9106), .IN1(n9105), .SEL(N38), .F(n9107) );
  MUX U9162 ( .IN0(n9107), .IN1(n9104), .SEL(N39), .F(n9108) );
  MUX U9163 ( .IN0(n9108), .IN1(n9101), .SEL(N40), .F(n9109) );
  MUX U9164 ( .IN0(data_mem_out_wire[469]), .IN1(data_mem_out_wire[501]), 
        .SEL(N37), .F(n9110) );
  MUX U9165 ( .IN0(data_mem_out_wire[405]), .IN1(data_mem_out_wire[437]), 
        .SEL(N37), .F(n9111) );
  MUX U9166 ( .IN0(n9111), .IN1(n9110), .SEL(N38), .F(n9112) );
  MUX U9167 ( .IN0(data_mem_out_wire[341]), .IN1(data_mem_out_wire[373]), 
        .SEL(N37), .F(n9113) );
  MUX U9168 ( .IN0(data_mem_out_wire[277]), .IN1(data_mem_out_wire[309]), 
        .SEL(N37), .F(n9114) );
  MUX U9169 ( .IN0(n9114), .IN1(n9113), .SEL(N38), .F(n9115) );
  MUX U9170 ( .IN0(n9115), .IN1(n9112), .SEL(N39), .F(n9116) );
  MUX U9171 ( .IN0(data_mem_out_wire[213]), .IN1(data_mem_out_wire[245]), 
        .SEL(N37), .F(n9117) );
  MUX U9172 ( .IN0(data_mem_out_wire[149]), .IN1(data_mem_out_wire[181]), 
        .SEL(N37), .F(n9118) );
  MUX U9173 ( .IN0(n9118), .IN1(n9117), .SEL(N38), .F(n9119) );
  MUX U9174 ( .IN0(data_mem_out_wire[85]), .IN1(data_mem_out_wire[117]), .SEL(
        N37), .F(n9120) );
  MUX U9175 ( .IN0(data_mem_out_wire[21]), .IN1(data_mem_out_wire[53]), .SEL(
        N37), .F(n9121) );
  MUX U9176 ( .IN0(n9121), .IN1(n9120), .SEL(N38), .F(n9122) );
  MUX U9177 ( .IN0(n9122), .IN1(n9119), .SEL(N39), .F(n9123) );
  MUX U9178 ( .IN0(n9123), .IN1(n9116), .SEL(N40), .F(n9124) );
  MUX U9179 ( .IN0(n9124), .IN1(n9109), .SEL(N41), .F(n9125) );
  MUX U9180 ( .IN0(n9125), .IN1(n9094), .SEL(N42), .F(N724) );
  MUX U9181 ( .IN0(data_mem_out_wire[2006]), .IN1(data_mem_out_wire[2038]), 
        .SEL(N37), .F(n9126) );
  MUX U9182 ( .IN0(data_mem_out_wire[1942]), .IN1(data_mem_out_wire[1974]), 
        .SEL(N37), .F(n9127) );
  MUX U9183 ( .IN0(n9127), .IN1(n9126), .SEL(N38), .F(n9128) );
  MUX U9184 ( .IN0(data_mem_out_wire[1878]), .IN1(data_mem_out_wire[1910]), 
        .SEL(N37), .F(n9129) );
  MUX U9185 ( .IN0(data_mem_out_wire[1814]), .IN1(data_mem_out_wire[1846]), 
        .SEL(N37), .F(n9130) );
  MUX U9186 ( .IN0(n9130), .IN1(n9129), .SEL(N38), .F(n9131) );
  MUX U9187 ( .IN0(n9131), .IN1(n9128), .SEL(N39), .F(n9132) );
  MUX U9188 ( .IN0(data_mem_out_wire[1750]), .IN1(data_mem_out_wire[1782]), 
        .SEL(N37), .F(n9133) );
  MUX U9189 ( .IN0(data_mem_out_wire[1686]), .IN1(data_mem_out_wire[1718]), 
        .SEL(N37), .F(n9134) );
  MUX U9190 ( .IN0(n9134), .IN1(n9133), .SEL(N38), .F(n9135) );
  MUX U9191 ( .IN0(data_mem_out_wire[1622]), .IN1(data_mem_out_wire[1654]), 
        .SEL(N37), .F(n9136) );
  MUX U9192 ( .IN0(data_mem_out_wire[1558]), .IN1(data_mem_out_wire[1590]), 
        .SEL(N37), .F(n9137) );
  MUX U9193 ( .IN0(n9137), .IN1(n9136), .SEL(N38), .F(n9138) );
  MUX U9194 ( .IN0(n9138), .IN1(n9135), .SEL(N39), .F(n9139) );
  MUX U9195 ( .IN0(n9139), .IN1(n9132), .SEL(N40), .F(n9140) );
  MUX U9196 ( .IN0(data_mem_out_wire[1494]), .IN1(data_mem_out_wire[1526]), 
        .SEL(N37), .F(n9141) );
  MUX U9197 ( .IN0(data_mem_out_wire[1430]), .IN1(data_mem_out_wire[1462]), 
        .SEL(N37), .F(n9142) );
  MUX U9198 ( .IN0(n9142), .IN1(n9141), .SEL(N38), .F(n9143) );
  MUX U9199 ( .IN0(data_mem_out_wire[1366]), .IN1(data_mem_out_wire[1398]), 
        .SEL(N37), .F(n9144) );
  MUX U9200 ( .IN0(data_mem_out_wire[1302]), .IN1(data_mem_out_wire[1334]), 
        .SEL(N37), .F(n9145) );
  MUX U9201 ( .IN0(n9145), .IN1(n9144), .SEL(N38), .F(n9146) );
  MUX U9202 ( .IN0(n9146), .IN1(n9143), .SEL(N39), .F(n9147) );
  MUX U9203 ( .IN0(data_mem_out_wire[1238]), .IN1(data_mem_out_wire[1270]), 
        .SEL(N37), .F(n9148) );
  MUX U9204 ( .IN0(data_mem_out_wire[1174]), .IN1(data_mem_out_wire[1206]), 
        .SEL(N37), .F(n9149) );
  MUX U9205 ( .IN0(n9149), .IN1(n9148), .SEL(N38), .F(n9150) );
  MUX U9206 ( .IN0(data_mem_out_wire[1110]), .IN1(data_mem_out_wire[1142]), 
        .SEL(N37), .F(n9151) );
  MUX U9207 ( .IN0(data_mem_out_wire[1046]), .IN1(data_mem_out_wire[1078]), 
        .SEL(N37), .F(n9152) );
  MUX U9208 ( .IN0(n9152), .IN1(n9151), .SEL(N38), .F(n9153) );
  MUX U9209 ( .IN0(n9153), .IN1(n9150), .SEL(N39), .F(n9154) );
  MUX U9210 ( .IN0(n9154), .IN1(n9147), .SEL(N40), .F(n9155) );
  MUX U9211 ( .IN0(n9155), .IN1(n9140), .SEL(N41), .F(n9156) );
  MUX U9212 ( .IN0(data_mem_out_wire[982]), .IN1(data_mem_out_wire[1014]), 
        .SEL(N37), .F(n9157) );
  MUX U9213 ( .IN0(data_mem_out_wire[918]), .IN1(data_mem_out_wire[950]), 
        .SEL(N37), .F(n9158) );
  MUX U9214 ( .IN0(n9158), .IN1(n9157), .SEL(N38), .F(n9159) );
  MUX U9215 ( .IN0(data_mem_out_wire[854]), .IN1(data_mem_out_wire[886]), 
        .SEL(N37), .F(n9160) );
  MUX U9216 ( .IN0(data_mem_out_wire[790]), .IN1(data_mem_out_wire[822]), 
        .SEL(N37), .F(n9161) );
  MUX U9217 ( .IN0(n9161), .IN1(n9160), .SEL(N38), .F(n9162) );
  MUX U9218 ( .IN0(n9162), .IN1(n9159), .SEL(N39), .F(n9163) );
  MUX U9219 ( .IN0(data_mem_out_wire[726]), .IN1(data_mem_out_wire[758]), 
        .SEL(N37), .F(n9164) );
  MUX U9220 ( .IN0(data_mem_out_wire[662]), .IN1(data_mem_out_wire[694]), 
        .SEL(N37), .F(n9165) );
  MUX U9221 ( .IN0(n9165), .IN1(n9164), .SEL(N38), .F(n9166) );
  MUX U9222 ( .IN0(data_mem_out_wire[598]), .IN1(data_mem_out_wire[630]), 
        .SEL(N37), .F(n9167) );
  MUX U9223 ( .IN0(data_mem_out_wire[534]), .IN1(data_mem_out_wire[566]), 
        .SEL(N37), .F(n9168) );
  MUX U9224 ( .IN0(n9168), .IN1(n9167), .SEL(N38), .F(n9169) );
  MUX U9225 ( .IN0(n9169), .IN1(n9166), .SEL(N39), .F(n9170) );
  MUX U9226 ( .IN0(n9170), .IN1(n9163), .SEL(N40), .F(n9171) );
  MUX U9227 ( .IN0(data_mem_out_wire[470]), .IN1(data_mem_out_wire[502]), 
        .SEL(N37), .F(n9172) );
  MUX U9228 ( .IN0(data_mem_out_wire[406]), .IN1(data_mem_out_wire[438]), 
        .SEL(N37), .F(n9173) );
  MUX U9229 ( .IN0(n9173), .IN1(n9172), .SEL(N38), .F(n9174) );
  MUX U9230 ( .IN0(data_mem_out_wire[342]), .IN1(data_mem_out_wire[374]), 
        .SEL(N37), .F(n9175) );
  MUX U9231 ( .IN0(data_mem_out_wire[278]), .IN1(data_mem_out_wire[310]), 
        .SEL(N37), .F(n9176) );
  MUX U9232 ( .IN0(n9176), .IN1(n9175), .SEL(N38), .F(n9177) );
  MUX U9233 ( .IN0(n9177), .IN1(n9174), .SEL(N39), .F(n9178) );
  MUX U9234 ( .IN0(data_mem_out_wire[214]), .IN1(data_mem_out_wire[246]), 
        .SEL(N37), .F(n9179) );
  MUX U9235 ( .IN0(data_mem_out_wire[150]), .IN1(data_mem_out_wire[182]), 
        .SEL(N37), .F(n9180) );
  MUX U9236 ( .IN0(n9180), .IN1(n9179), .SEL(N38), .F(n9181) );
  MUX U9237 ( .IN0(data_mem_out_wire[86]), .IN1(data_mem_out_wire[118]), .SEL(
        N37), .F(n9182) );
  MUX U9238 ( .IN0(data_mem_out_wire[22]), .IN1(data_mem_out_wire[54]), .SEL(
        N37), .F(n9183) );
  MUX U9239 ( .IN0(n9183), .IN1(n9182), .SEL(N38), .F(n9184) );
  MUX U9240 ( .IN0(n9184), .IN1(n9181), .SEL(N39), .F(n9185) );
  MUX U9241 ( .IN0(n9185), .IN1(n9178), .SEL(N40), .F(n9186) );
  MUX U9242 ( .IN0(n9186), .IN1(n9171), .SEL(N41), .F(n9187) );
  MUX U9243 ( .IN0(n9187), .IN1(n9156), .SEL(N42), .F(N723) );
  MUX U9244 ( .IN0(data_mem_out_wire[2007]), .IN1(data_mem_out_wire[2039]), 
        .SEL(N37), .F(n9188) );
  MUX U9245 ( .IN0(data_mem_out_wire[1943]), .IN1(data_mem_out_wire[1975]), 
        .SEL(N37), .F(n9189) );
  MUX U9246 ( .IN0(n9189), .IN1(n9188), .SEL(N38), .F(n9190) );
  MUX U9247 ( .IN0(data_mem_out_wire[1879]), .IN1(data_mem_out_wire[1911]), 
        .SEL(N37), .F(n9191) );
  MUX U9248 ( .IN0(data_mem_out_wire[1815]), .IN1(data_mem_out_wire[1847]), 
        .SEL(N37), .F(n9192) );
  MUX U9249 ( .IN0(n9192), .IN1(n9191), .SEL(N38), .F(n9193) );
  MUX U9250 ( .IN0(n9193), .IN1(n9190), .SEL(N39), .F(n9194) );
  MUX U9251 ( .IN0(data_mem_out_wire[1751]), .IN1(data_mem_out_wire[1783]), 
        .SEL(N37), .F(n9195) );
  MUX U9252 ( .IN0(data_mem_out_wire[1687]), .IN1(data_mem_out_wire[1719]), 
        .SEL(N37), .F(n9196) );
  MUX U9253 ( .IN0(n9196), .IN1(n9195), .SEL(N38), .F(n9197) );
  MUX U9254 ( .IN0(data_mem_out_wire[1623]), .IN1(data_mem_out_wire[1655]), 
        .SEL(N37), .F(n9198) );
  MUX U9255 ( .IN0(data_mem_out_wire[1559]), .IN1(data_mem_out_wire[1591]), 
        .SEL(N37), .F(n9199) );
  MUX U9256 ( .IN0(n9199), .IN1(n9198), .SEL(N38), .F(n9200) );
  MUX U9257 ( .IN0(n9200), .IN1(n9197), .SEL(N39), .F(n9201) );
  MUX U9258 ( .IN0(n9201), .IN1(n9194), .SEL(N40), .F(n9202) );
  MUX U9259 ( .IN0(data_mem_out_wire[1495]), .IN1(data_mem_out_wire[1527]), 
        .SEL(N37), .F(n9203) );
  MUX U9260 ( .IN0(data_mem_out_wire[1431]), .IN1(data_mem_out_wire[1463]), 
        .SEL(N37), .F(n9204) );
  MUX U9261 ( .IN0(n9204), .IN1(n9203), .SEL(N38), .F(n9205) );
  MUX U9262 ( .IN0(data_mem_out_wire[1367]), .IN1(data_mem_out_wire[1399]), 
        .SEL(N37), .F(n9206) );
  MUX U9263 ( .IN0(data_mem_out_wire[1303]), .IN1(data_mem_out_wire[1335]), 
        .SEL(N37), .F(n9207) );
  MUX U9264 ( .IN0(n9207), .IN1(n9206), .SEL(N38), .F(n9208) );
  MUX U9265 ( .IN0(n9208), .IN1(n9205), .SEL(N39), .F(n9209) );
  MUX U9266 ( .IN0(data_mem_out_wire[1239]), .IN1(data_mem_out_wire[1271]), 
        .SEL(N37), .F(n9210) );
  MUX U9267 ( .IN0(data_mem_out_wire[1175]), .IN1(data_mem_out_wire[1207]), 
        .SEL(N37), .F(n9211) );
  MUX U9268 ( .IN0(n9211), .IN1(n9210), .SEL(N38), .F(n9212) );
  MUX U9269 ( .IN0(data_mem_out_wire[1111]), .IN1(data_mem_out_wire[1143]), 
        .SEL(N37), .F(n9213) );
  MUX U9270 ( .IN0(data_mem_out_wire[1047]), .IN1(data_mem_out_wire[1079]), 
        .SEL(N37), .F(n9214) );
  MUX U9271 ( .IN0(n9214), .IN1(n9213), .SEL(N38), .F(n9215) );
  MUX U9272 ( .IN0(n9215), .IN1(n9212), .SEL(N39), .F(n9216) );
  MUX U9273 ( .IN0(n9216), .IN1(n9209), .SEL(N40), .F(n9217) );
  MUX U9274 ( .IN0(n9217), .IN1(n9202), .SEL(N41), .F(n9218) );
  MUX U9275 ( .IN0(data_mem_out_wire[983]), .IN1(data_mem_out_wire[1015]), 
        .SEL(N37), .F(n9219) );
  MUX U9276 ( .IN0(data_mem_out_wire[919]), .IN1(data_mem_out_wire[951]), 
        .SEL(N37), .F(n9220) );
  MUX U9277 ( .IN0(n9220), .IN1(n9219), .SEL(N38), .F(n9221) );
  MUX U9278 ( .IN0(data_mem_out_wire[855]), .IN1(data_mem_out_wire[887]), 
        .SEL(N37), .F(n9222) );
  MUX U9279 ( .IN0(data_mem_out_wire[791]), .IN1(data_mem_out_wire[823]), 
        .SEL(N37), .F(n9223) );
  MUX U9280 ( .IN0(n9223), .IN1(n9222), .SEL(N38), .F(n9224) );
  MUX U9281 ( .IN0(n9224), .IN1(n9221), .SEL(N39), .F(n9225) );
  MUX U9282 ( .IN0(data_mem_out_wire[727]), .IN1(data_mem_out_wire[759]), 
        .SEL(N37), .F(n9226) );
  MUX U9283 ( .IN0(data_mem_out_wire[663]), .IN1(data_mem_out_wire[695]), 
        .SEL(N37), .F(n9227) );
  MUX U9284 ( .IN0(n9227), .IN1(n9226), .SEL(N38), .F(n9228) );
  MUX U9285 ( .IN0(data_mem_out_wire[599]), .IN1(data_mem_out_wire[631]), 
        .SEL(N37), .F(n9229) );
  MUX U9286 ( .IN0(data_mem_out_wire[535]), .IN1(data_mem_out_wire[567]), 
        .SEL(N37), .F(n9230) );
  MUX U9287 ( .IN0(n9230), .IN1(n9229), .SEL(N38), .F(n9231) );
  MUX U9288 ( .IN0(n9231), .IN1(n9228), .SEL(N39), .F(n9232) );
  MUX U9289 ( .IN0(n9232), .IN1(n9225), .SEL(N40), .F(n9233) );
  MUX U9290 ( .IN0(data_mem_out_wire[471]), .IN1(data_mem_out_wire[503]), 
        .SEL(N37), .F(n9234) );
  MUX U9291 ( .IN0(data_mem_out_wire[407]), .IN1(data_mem_out_wire[439]), 
        .SEL(N37), .F(n9235) );
  MUX U9292 ( .IN0(n9235), .IN1(n9234), .SEL(N38), .F(n9236) );
  MUX U9293 ( .IN0(data_mem_out_wire[343]), .IN1(data_mem_out_wire[375]), 
        .SEL(N37), .F(n9237) );
  MUX U9294 ( .IN0(data_mem_out_wire[279]), .IN1(data_mem_out_wire[311]), 
        .SEL(N37), .F(n9238) );
  MUX U9295 ( .IN0(n9238), .IN1(n9237), .SEL(N38), .F(n9239) );
  MUX U9296 ( .IN0(n9239), .IN1(n9236), .SEL(N39), .F(n9240) );
  MUX U9297 ( .IN0(data_mem_out_wire[215]), .IN1(data_mem_out_wire[247]), 
        .SEL(N37), .F(n9241) );
  MUX U9298 ( .IN0(data_mem_out_wire[151]), .IN1(data_mem_out_wire[183]), 
        .SEL(N37), .F(n9242) );
  MUX U9299 ( .IN0(n9242), .IN1(n9241), .SEL(N38), .F(n9243) );
  MUX U9300 ( .IN0(data_mem_out_wire[87]), .IN1(data_mem_out_wire[119]), .SEL(
        N37), .F(n9244) );
  MUX U9301 ( .IN0(data_mem_out_wire[23]), .IN1(data_mem_out_wire[55]), .SEL(
        N37), .F(n9245) );
  MUX U9302 ( .IN0(n9245), .IN1(n9244), .SEL(N38), .F(n9246) );
  MUX U9303 ( .IN0(n9246), .IN1(n9243), .SEL(N39), .F(n9247) );
  MUX U9304 ( .IN0(n9247), .IN1(n9240), .SEL(N40), .F(n9248) );
  MUX U9305 ( .IN0(n9248), .IN1(n9233), .SEL(N41), .F(n9249) );
  MUX U9306 ( .IN0(n9249), .IN1(n9218), .SEL(N42), .F(N722) );
  MUX U9307 ( .IN0(data_mem_out_wire[2008]), .IN1(data_mem_out_wire[2040]), 
        .SEL(N37), .F(n9250) );
  MUX U9308 ( .IN0(data_mem_out_wire[1944]), .IN1(data_mem_out_wire[1976]), 
        .SEL(N37), .F(n9251) );
  MUX U9309 ( .IN0(n9251), .IN1(n9250), .SEL(N38), .F(n9252) );
  MUX U9310 ( .IN0(data_mem_out_wire[1880]), .IN1(data_mem_out_wire[1912]), 
        .SEL(N37), .F(n9253) );
  MUX U9311 ( .IN0(data_mem_out_wire[1816]), .IN1(data_mem_out_wire[1848]), 
        .SEL(N37), .F(n9254) );
  MUX U9312 ( .IN0(n9254), .IN1(n9253), .SEL(N38), .F(n9255) );
  MUX U9313 ( .IN0(n9255), .IN1(n9252), .SEL(N39), .F(n9256) );
  MUX U9314 ( .IN0(data_mem_out_wire[1752]), .IN1(data_mem_out_wire[1784]), 
        .SEL(N37), .F(n9257) );
  MUX U9315 ( .IN0(data_mem_out_wire[1688]), .IN1(data_mem_out_wire[1720]), 
        .SEL(N37), .F(n9258) );
  MUX U9316 ( .IN0(n9258), .IN1(n9257), .SEL(N38), .F(n9259) );
  MUX U9317 ( .IN0(data_mem_out_wire[1624]), .IN1(data_mem_out_wire[1656]), 
        .SEL(N37), .F(n9260) );
  MUX U9318 ( .IN0(data_mem_out_wire[1560]), .IN1(data_mem_out_wire[1592]), 
        .SEL(N37), .F(n9261) );
  MUX U9319 ( .IN0(n9261), .IN1(n9260), .SEL(N38), .F(n9262) );
  MUX U9320 ( .IN0(n9262), .IN1(n9259), .SEL(N39), .F(n9263) );
  MUX U9321 ( .IN0(n9263), .IN1(n9256), .SEL(N40), .F(n9264) );
  MUX U9322 ( .IN0(data_mem_out_wire[1496]), .IN1(data_mem_out_wire[1528]), 
        .SEL(N37), .F(n9265) );
  MUX U9323 ( .IN0(data_mem_out_wire[1432]), .IN1(data_mem_out_wire[1464]), 
        .SEL(N37), .F(n9266) );
  MUX U9324 ( .IN0(n9266), .IN1(n9265), .SEL(N38), .F(n9267) );
  MUX U9325 ( .IN0(data_mem_out_wire[1368]), .IN1(data_mem_out_wire[1400]), 
        .SEL(N37), .F(n9268) );
  MUX U9326 ( .IN0(data_mem_out_wire[1304]), .IN1(data_mem_out_wire[1336]), 
        .SEL(N37), .F(n9269) );
  MUX U9327 ( .IN0(n9269), .IN1(n9268), .SEL(N38), .F(n9270) );
  MUX U9328 ( .IN0(n9270), .IN1(n9267), .SEL(N39), .F(n9271) );
  MUX U9329 ( .IN0(data_mem_out_wire[1240]), .IN1(data_mem_out_wire[1272]), 
        .SEL(N37), .F(n9272) );
  MUX U9330 ( .IN0(data_mem_out_wire[1176]), .IN1(data_mem_out_wire[1208]), 
        .SEL(N37), .F(n9273) );
  MUX U9331 ( .IN0(n9273), .IN1(n9272), .SEL(N38), .F(n9274) );
  MUX U9332 ( .IN0(data_mem_out_wire[1112]), .IN1(data_mem_out_wire[1144]), 
        .SEL(N37), .F(n9275) );
  MUX U9333 ( .IN0(data_mem_out_wire[1048]), .IN1(data_mem_out_wire[1080]), 
        .SEL(N37), .F(n9276) );
  MUX U9334 ( .IN0(n9276), .IN1(n9275), .SEL(N38), .F(n9277) );
  MUX U9335 ( .IN0(n9277), .IN1(n9274), .SEL(N39), .F(n9278) );
  MUX U9336 ( .IN0(n9278), .IN1(n9271), .SEL(N40), .F(n9279) );
  MUX U9337 ( .IN0(n9279), .IN1(n9264), .SEL(N41), .F(n9280) );
  MUX U9338 ( .IN0(data_mem_out_wire[984]), .IN1(data_mem_out_wire[1016]), 
        .SEL(N37), .F(n9281) );
  MUX U9339 ( .IN0(data_mem_out_wire[920]), .IN1(data_mem_out_wire[952]), 
        .SEL(N37), .F(n9282) );
  MUX U9340 ( .IN0(n9282), .IN1(n9281), .SEL(N38), .F(n9283) );
  MUX U9341 ( .IN0(data_mem_out_wire[856]), .IN1(data_mem_out_wire[888]), 
        .SEL(N37), .F(n9284) );
  MUX U9342 ( .IN0(data_mem_out_wire[792]), .IN1(data_mem_out_wire[824]), 
        .SEL(N37), .F(n9285) );
  MUX U9343 ( .IN0(n9285), .IN1(n9284), .SEL(N38), .F(n9286) );
  MUX U9344 ( .IN0(n9286), .IN1(n9283), .SEL(N39), .F(n9287) );
  MUX U9345 ( .IN0(data_mem_out_wire[728]), .IN1(data_mem_out_wire[760]), 
        .SEL(N37), .F(n9288) );
  MUX U9346 ( .IN0(data_mem_out_wire[664]), .IN1(data_mem_out_wire[696]), 
        .SEL(N37), .F(n9289) );
  MUX U9347 ( .IN0(n9289), .IN1(n9288), .SEL(N38), .F(n9290) );
  MUX U9348 ( .IN0(data_mem_out_wire[600]), .IN1(data_mem_out_wire[632]), 
        .SEL(N37), .F(n9291) );
  MUX U9349 ( .IN0(data_mem_out_wire[536]), .IN1(data_mem_out_wire[568]), 
        .SEL(N37), .F(n9292) );
  MUX U9350 ( .IN0(n9292), .IN1(n9291), .SEL(N38), .F(n9293) );
  MUX U9351 ( .IN0(n9293), .IN1(n9290), .SEL(N39), .F(n9294) );
  MUX U9352 ( .IN0(n9294), .IN1(n9287), .SEL(N40), .F(n9295) );
  MUX U9353 ( .IN0(data_mem_out_wire[472]), .IN1(data_mem_out_wire[504]), 
        .SEL(N37), .F(n9296) );
  MUX U9354 ( .IN0(data_mem_out_wire[408]), .IN1(data_mem_out_wire[440]), 
        .SEL(N37), .F(n9297) );
  MUX U9355 ( .IN0(n9297), .IN1(n9296), .SEL(N38), .F(n9298) );
  MUX U9356 ( .IN0(data_mem_out_wire[344]), .IN1(data_mem_out_wire[376]), 
        .SEL(N37), .F(n9299) );
  MUX U9357 ( .IN0(data_mem_out_wire[280]), .IN1(data_mem_out_wire[312]), 
        .SEL(N37), .F(n9300) );
  MUX U9358 ( .IN0(n9300), .IN1(n9299), .SEL(N38), .F(n9301) );
  MUX U9359 ( .IN0(n9301), .IN1(n9298), .SEL(N39), .F(n9302) );
  MUX U9360 ( .IN0(data_mem_out_wire[216]), .IN1(data_mem_out_wire[248]), 
        .SEL(N37), .F(n9303) );
  MUX U9361 ( .IN0(data_mem_out_wire[152]), .IN1(data_mem_out_wire[184]), 
        .SEL(N37), .F(n9304) );
  MUX U9362 ( .IN0(n9304), .IN1(n9303), .SEL(N38), .F(n9305) );
  MUX U9363 ( .IN0(data_mem_out_wire[88]), .IN1(data_mem_out_wire[120]), .SEL(
        N37), .F(n9306) );
  MUX U9364 ( .IN0(data_mem_out_wire[24]), .IN1(data_mem_out_wire[56]), .SEL(
        N37), .F(n9307) );
  MUX U9365 ( .IN0(n9307), .IN1(n9306), .SEL(N38), .F(n9308) );
  MUX U9366 ( .IN0(n9308), .IN1(n9305), .SEL(N39), .F(n9309) );
  MUX U9367 ( .IN0(n9309), .IN1(n9302), .SEL(N40), .F(n9310) );
  MUX U9368 ( .IN0(n9310), .IN1(n9295), .SEL(N41), .F(n9311) );
  MUX U9369 ( .IN0(n9311), .IN1(n9280), .SEL(N42), .F(N721) );
  MUX U9370 ( .IN0(data_mem_out_wire[2009]), .IN1(data_mem_out_wire[2041]), 
        .SEL(N37), .F(n9312) );
  MUX U9371 ( .IN0(data_mem_out_wire[1945]), .IN1(data_mem_out_wire[1977]), 
        .SEL(N37), .F(n9313) );
  MUX U9372 ( .IN0(n9313), .IN1(n9312), .SEL(N38), .F(n9314) );
  MUX U9373 ( .IN0(data_mem_out_wire[1881]), .IN1(data_mem_out_wire[1913]), 
        .SEL(N37), .F(n9315) );
  MUX U9374 ( .IN0(data_mem_out_wire[1817]), .IN1(data_mem_out_wire[1849]), 
        .SEL(N37), .F(n9316) );
  MUX U9375 ( .IN0(n9316), .IN1(n9315), .SEL(N38), .F(n9317) );
  MUX U9376 ( .IN0(n9317), .IN1(n9314), .SEL(N39), .F(n9318) );
  MUX U9377 ( .IN0(data_mem_out_wire[1753]), .IN1(data_mem_out_wire[1785]), 
        .SEL(N37), .F(n9319) );
  MUX U9378 ( .IN0(data_mem_out_wire[1689]), .IN1(data_mem_out_wire[1721]), 
        .SEL(N37), .F(n9320) );
  MUX U9379 ( .IN0(n9320), .IN1(n9319), .SEL(N38), .F(n9321) );
  MUX U9380 ( .IN0(data_mem_out_wire[1625]), .IN1(data_mem_out_wire[1657]), 
        .SEL(N37), .F(n9322) );
  MUX U9381 ( .IN0(data_mem_out_wire[1561]), .IN1(data_mem_out_wire[1593]), 
        .SEL(N37), .F(n9323) );
  MUX U9382 ( .IN0(n9323), .IN1(n9322), .SEL(N38), .F(n9324) );
  MUX U9383 ( .IN0(n9324), .IN1(n9321), .SEL(N39), .F(n9325) );
  MUX U9384 ( .IN0(n9325), .IN1(n9318), .SEL(N40), .F(n9326) );
  MUX U9385 ( .IN0(data_mem_out_wire[1497]), .IN1(data_mem_out_wire[1529]), 
        .SEL(N37), .F(n9327) );
  MUX U9386 ( .IN0(data_mem_out_wire[1433]), .IN1(data_mem_out_wire[1465]), 
        .SEL(N37), .F(n9328) );
  MUX U9387 ( .IN0(n9328), .IN1(n9327), .SEL(N38), .F(n9329) );
  MUX U9388 ( .IN0(data_mem_out_wire[1369]), .IN1(data_mem_out_wire[1401]), 
        .SEL(N37), .F(n9330) );
  MUX U9389 ( .IN0(data_mem_out_wire[1305]), .IN1(data_mem_out_wire[1337]), 
        .SEL(N37), .F(n9331) );
  MUX U9390 ( .IN0(n9331), .IN1(n9330), .SEL(N38), .F(n9332) );
  MUX U9391 ( .IN0(n9332), .IN1(n9329), .SEL(N39), .F(n9333) );
  MUX U9392 ( .IN0(data_mem_out_wire[1241]), .IN1(data_mem_out_wire[1273]), 
        .SEL(N37), .F(n9334) );
  MUX U9393 ( .IN0(data_mem_out_wire[1177]), .IN1(data_mem_out_wire[1209]), 
        .SEL(N37), .F(n9335) );
  MUX U9394 ( .IN0(n9335), .IN1(n9334), .SEL(N38), .F(n9336) );
  MUX U9395 ( .IN0(data_mem_out_wire[1113]), .IN1(data_mem_out_wire[1145]), 
        .SEL(N37), .F(n9337) );
  MUX U9396 ( .IN0(data_mem_out_wire[1049]), .IN1(data_mem_out_wire[1081]), 
        .SEL(N37), .F(n9338) );
  MUX U9397 ( .IN0(n9338), .IN1(n9337), .SEL(N38), .F(n9339) );
  MUX U9398 ( .IN0(n9339), .IN1(n9336), .SEL(N39), .F(n9340) );
  MUX U9399 ( .IN0(n9340), .IN1(n9333), .SEL(N40), .F(n9341) );
  MUX U9400 ( .IN0(n9341), .IN1(n9326), .SEL(N41), .F(n9342) );
  MUX U9401 ( .IN0(data_mem_out_wire[985]), .IN1(data_mem_out_wire[1017]), 
        .SEL(N37), .F(n9343) );
  MUX U9402 ( .IN0(data_mem_out_wire[921]), .IN1(data_mem_out_wire[953]), 
        .SEL(N37), .F(n9344) );
  MUX U9403 ( .IN0(n9344), .IN1(n9343), .SEL(N38), .F(n9345) );
  MUX U9404 ( .IN0(data_mem_out_wire[857]), .IN1(data_mem_out_wire[889]), 
        .SEL(N37), .F(n9346) );
  MUX U9405 ( .IN0(data_mem_out_wire[793]), .IN1(data_mem_out_wire[825]), 
        .SEL(N37), .F(n9347) );
  MUX U9406 ( .IN0(n9347), .IN1(n9346), .SEL(N38), .F(n9348) );
  MUX U9407 ( .IN0(n9348), .IN1(n9345), .SEL(N39), .F(n9349) );
  MUX U9408 ( .IN0(data_mem_out_wire[729]), .IN1(data_mem_out_wire[761]), 
        .SEL(N37), .F(n9350) );
  MUX U9409 ( .IN0(data_mem_out_wire[665]), .IN1(data_mem_out_wire[697]), 
        .SEL(N37), .F(n9351) );
  MUX U9410 ( .IN0(n9351), .IN1(n9350), .SEL(N38), .F(n9352) );
  MUX U9411 ( .IN0(data_mem_out_wire[601]), .IN1(data_mem_out_wire[633]), 
        .SEL(N37), .F(n9353) );
  MUX U9412 ( .IN0(data_mem_out_wire[537]), .IN1(data_mem_out_wire[569]), 
        .SEL(N37), .F(n9354) );
  MUX U9413 ( .IN0(n9354), .IN1(n9353), .SEL(N38), .F(n9355) );
  MUX U9414 ( .IN0(n9355), .IN1(n9352), .SEL(N39), .F(n9356) );
  MUX U9415 ( .IN0(n9356), .IN1(n9349), .SEL(N40), .F(n9357) );
  MUX U9416 ( .IN0(data_mem_out_wire[473]), .IN1(data_mem_out_wire[505]), 
        .SEL(N37), .F(n9358) );
  MUX U9417 ( .IN0(data_mem_out_wire[409]), .IN1(data_mem_out_wire[441]), 
        .SEL(N37), .F(n9359) );
  MUX U9418 ( .IN0(n9359), .IN1(n9358), .SEL(N38), .F(n9360) );
  MUX U9419 ( .IN0(data_mem_out_wire[345]), .IN1(data_mem_out_wire[377]), 
        .SEL(N37), .F(n9361) );
  MUX U9420 ( .IN0(data_mem_out_wire[281]), .IN1(data_mem_out_wire[313]), 
        .SEL(N37), .F(n9362) );
  MUX U9421 ( .IN0(n9362), .IN1(n9361), .SEL(N38), .F(n9363) );
  MUX U9422 ( .IN0(n9363), .IN1(n9360), .SEL(N39), .F(n9364) );
  MUX U9423 ( .IN0(data_mem_out_wire[217]), .IN1(data_mem_out_wire[249]), 
        .SEL(N37), .F(n9365) );
  MUX U9424 ( .IN0(data_mem_out_wire[153]), .IN1(data_mem_out_wire[185]), 
        .SEL(N37), .F(n9366) );
  MUX U9425 ( .IN0(n9366), .IN1(n9365), .SEL(N38), .F(n9367) );
  MUX U9426 ( .IN0(data_mem_out_wire[89]), .IN1(data_mem_out_wire[121]), .SEL(
        N37), .F(n9368) );
  MUX U9427 ( .IN0(data_mem_out_wire[25]), .IN1(data_mem_out_wire[57]), .SEL(
        N37), .F(n9369) );
  MUX U9428 ( .IN0(n9369), .IN1(n9368), .SEL(N38), .F(n9370) );
  MUX U9429 ( .IN0(n9370), .IN1(n9367), .SEL(N39), .F(n9371) );
  MUX U9430 ( .IN0(n9371), .IN1(n9364), .SEL(N40), .F(n9372) );
  MUX U9431 ( .IN0(n9372), .IN1(n9357), .SEL(N41), .F(n9373) );
  MUX U9432 ( .IN0(n9373), .IN1(n9342), .SEL(N42), .F(N720) );
  MUX U9433 ( .IN0(data_mem_out_wire[2010]), .IN1(data_mem_out_wire[2042]), 
        .SEL(N37), .F(n9374) );
  MUX U9434 ( .IN0(data_mem_out_wire[1946]), .IN1(data_mem_out_wire[1978]), 
        .SEL(N37), .F(n9375) );
  MUX U9435 ( .IN0(n9375), .IN1(n9374), .SEL(N38), .F(n9376) );
  MUX U9436 ( .IN0(data_mem_out_wire[1882]), .IN1(data_mem_out_wire[1914]), 
        .SEL(N37), .F(n9377) );
  MUX U9437 ( .IN0(data_mem_out_wire[1818]), .IN1(data_mem_out_wire[1850]), 
        .SEL(N37), .F(n9378) );
  MUX U9438 ( .IN0(n9378), .IN1(n9377), .SEL(N38), .F(n9379) );
  MUX U9439 ( .IN0(n9379), .IN1(n9376), .SEL(N39), .F(n9380) );
  MUX U9440 ( .IN0(data_mem_out_wire[1754]), .IN1(data_mem_out_wire[1786]), 
        .SEL(N37), .F(n9381) );
  MUX U9441 ( .IN0(data_mem_out_wire[1690]), .IN1(data_mem_out_wire[1722]), 
        .SEL(N37), .F(n9382) );
  MUX U9442 ( .IN0(n9382), .IN1(n9381), .SEL(N38), .F(n9383) );
  MUX U9443 ( .IN0(data_mem_out_wire[1626]), .IN1(data_mem_out_wire[1658]), 
        .SEL(N37), .F(n9384) );
  MUX U9444 ( .IN0(data_mem_out_wire[1562]), .IN1(data_mem_out_wire[1594]), 
        .SEL(N37), .F(n9385) );
  MUX U9445 ( .IN0(n9385), .IN1(n9384), .SEL(N38), .F(n9386) );
  MUX U9446 ( .IN0(n9386), .IN1(n9383), .SEL(N39), .F(n9387) );
  MUX U9447 ( .IN0(n9387), .IN1(n9380), .SEL(N40), .F(n9388) );
  MUX U9448 ( .IN0(data_mem_out_wire[1498]), .IN1(data_mem_out_wire[1530]), 
        .SEL(N37), .F(n9389) );
  MUX U9449 ( .IN0(data_mem_out_wire[1434]), .IN1(data_mem_out_wire[1466]), 
        .SEL(N37), .F(n9390) );
  MUX U9450 ( .IN0(n9390), .IN1(n9389), .SEL(N38), .F(n9391) );
  MUX U9451 ( .IN0(data_mem_out_wire[1370]), .IN1(data_mem_out_wire[1402]), 
        .SEL(N37), .F(n9392) );
  MUX U9452 ( .IN0(data_mem_out_wire[1306]), .IN1(data_mem_out_wire[1338]), 
        .SEL(N37), .F(n9393) );
  MUX U9453 ( .IN0(n9393), .IN1(n9392), .SEL(N38), .F(n9394) );
  MUX U9454 ( .IN0(n9394), .IN1(n9391), .SEL(N39), .F(n9395) );
  MUX U9455 ( .IN0(data_mem_out_wire[1242]), .IN1(data_mem_out_wire[1274]), 
        .SEL(N37), .F(n9396) );
  MUX U9456 ( .IN0(data_mem_out_wire[1178]), .IN1(data_mem_out_wire[1210]), 
        .SEL(N37), .F(n9397) );
  MUX U9457 ( .IN0(n9397), .IN1(n9396), .SEL(N38), .F(n9398) );
  MUX U9458 ( .IN0(data_mem_out_wire[1114]), .IN1(data_mem_out_wire[1146]), 
        .SEL(N37), .F(n9399) );
  MUX U9459 ( .IN0(data_mem_out_wire[1050]), .IN1(data_mem_out_wire[1082]), 
        .SEL(N37), .F(n9400) );
  MUX U9460 ( .IN0(n9400), .IN1(n9399), .SEL(N38), .F(n9401) );
  MUX U9461 ( .IN0(n9401), .IN1(n9398), .SEL(N39), .F(n9402) );
  MUX U9462 ( .IN0(n9402), .IN1(n9395), .SEL(N40), .F(n9403) );
  MUX U9463 ( .IN0(n9403), .IN1(n9388), .SEL(N41), .F(n9404) );
  MUX U9464 ( .IN0(data_mem_out_wire[986]), .IN1(data_mem_out_wire[1018]), 
        .SEL(N37), .F(n9405) );
  MUX U9465 ( .IN0(data_mem_out_wire[922]), .IN1(data_mem_out_wire[954]), 
        .SEL(N37), .F(n9406) );
  MUX U9466 ( .IN0(n9406), .IN1(n9405), .SEL(N38), .F(n9407) );
  MUX U9467 ( .IN0(data_mem_out_wire[858]), .IN1(data_mem_out_wire[890]), 
        .SEL(N37), .F(n9408) );
  MUX U9468 ( .IN0(data_mem_out_wire[794]), .IN1(data_mem_out_wire[826]), 
        .SEL(N37), .F(n9409) );
  MUX U9469 ( .IN0(n9409), .IN1(n9408), .SEL(N38), .F(n9410) );
  MUX U9470 ( .IN0(n9410), .IN1(n9407), .SEL(N39), .F(n9411) );
  MUX U9471 ( .IN0(data_mem_out_wire[730]), .IN1(data_mem_out_wire[762]), 
        .SEL(N37), .F(n9412) );
  MUX U9472 ( .IN0(data_mem_out_wire[666]), .IN1(data_mem_out_wire[698]), 
        .SEL(N37), .F(n9413) );
  MUX U9473 ( .IN0(n9413), .IN1(n9412), .SEL(N38), .F(n9414) );
  MUX U9474 ( .IN0(data_mem_out_wire[602]), .IN1(data_mem_out_wire[634]), 
        .SEL(N37), .F(n9415) );
  MUX U9475 ( .IN0(data_mem_out_wire[538]), .IN1(data_mem_out_wire[570]), 
        .SEL(N37), .F(n9416) );
  MUX U9476 ( .IN0(n9416), .IN1(n9415), .SEL(N38), .F(n9417) );
  MUX U9477 ( .IN0(n9417), .IN1(n9414), .SEL(N39), .F(n9418) );
  MUX U9478 ( .IN0(n9418), .IN1(n9411), .SEL(N40), .F(n9419) );
  MUX U9479 ( .IN0(data_mem_out_wire[474]), .IN1(data_mem_out_wire[506]), 
        .SEL(N37), .F(n9420) );
  MUX U9480 ( .IN0(data_mem_out_wire[410]), .IN1(data_mem_out_wire[442]), 
        .SEL(N37), .F(n9421) );
  MUX U9481 ( .IN0(n9421), .IN1(n9420), .SEL(N38), .F(n9422) );
  MUX U9482 ( .IN0(data_mem_out_wire[346]), .IN1(data_mem_out_wire[378]), 
        .SEL(N37), .F(n9423) );
  MUX U9483 ( .IN0(data_mem_out_wire[282]), .IN1(data_mem_out_wire[314]), 
        .SEL(N37), .F(n9424) );
  MUX U9484 ( .IN0(n9424), .IN1(n9423), .SEL(N38), .F(n9425) );
  MUX U9485 ( .IN0(n9425), .IN1(n9422), .SEL(N39), .F(n9426) );
  MUX U9486 ( .IN0(data_mem_out_wire[218]), .IN1(data_mem_out_wire[250]), 
        .SEL(N37), .F(n9427) );
  MUX U9487 ( .IN0(data_mem_out_wire[154]), .IN1(data_mem_out_wire[186]), 
        .SEL(N37), .F(n9428) );
  MUX U9488 ( .IN0(n9428), .IN1(n9427), .SEL(N38), .F(n9429) );
  MUX U9489 ( .IN0(data_mem_out_wire[90]), .IN1(data_mem_out_wire[122]), .SEL(
        N37), .F(n9430) );
  MUX U9490 ( .IN0(data_mem_out_wire[26]), .IN1(data_mem_out_wire[58]), .SEL(
        N37), .F(n9431) );
  MUX U9491 ( .IN0(n9431), .IN1(n9430), .SEL(N38), .F(n9432) );
  MUX U9492 ( .IN0(n9432), .IN1(n9429), .SEL(N39), .F(n9433) );
  MUX U9493 ( .IN0(n9433), .IN1(n9426), .SEL(N40), .F(n9434) );
  MUX U9494 ( .IN0(n9434), .IN1(n9419), .SEL(N41), .F(n9435) );
  MUX U9495 ( .IN0(n9435), .IN1(n9404), .SEL(N42), .F(N719) );
  MUX U9496 ( .IN0(data_mem_out_wire[2011]), .IN1(data_mem_out_wire[2043]), 
        .SEL(N37), .F(n9436) );
  MUX U9497 ( .IN0(data_mem_out_wire[1947]), .IN1(data_mem_out_wire[1979]), 
        .SEL(N37), .F(n9437) );
  MUX U9498 ( .IN0(n9437), .IN1(n9436), .SEL(N38), .F(n9438) );
  MUX U9499 ( .IN0(data_mem_out_wire[1883]), .IN1(data_mem_out_wire[1915]), 
        .SEL(N37), .F(n9439) );
  MUX U9500 ( .IN0(data_mem_out_wire[1819]), .IN1(data_mem_out_wire[1851]), 
        .SEL(N37), .F(n9440) );
  MUX U9501 ( .IN0(n9440), .IN1(n9439), .SEL(N38), .F(n9441) );
  MUX U9502 ( .IN0(n9441), .IN1(n9438), .SEL(N39), .F(n9442) );
  MUX U9503 ( .IN0(data_mem_out_wire[1755]), .IN1(data_mem_out_wire[1787]), 
        .SEL(N37), .F(n9443) );
  MUX U9504 ( .IN0(data_mem_out_wire[1691]), .IN1(data_mem_out_wire[1723]), 
        .SEL(N37), .F(n9444) );
  MUX U9505 ( .IN0(n9444), .IN1(n9443), .SEL(N38), .F(n9445) );
  MUX U9506 ( .IN0(data_mem_out_wire[1627]), .IN1(data_mem_out_wire[1659]), 
        .SEL(N37), .F(n9446) );
  MUX U9507 ( .IN0(data_mem_out_wire[1563]), .IN1(data_mem_out_wire[1595]), 
        .SEL(N37), .F(n9447) );
  MUX U9508 ( .IN0(n9447), .IN1(n9446), .SEL(N38), .F(n9448) );
  MUX U9509 ( .IN0(n9448), .IN1(n9445), .SEL(N39), .F(n9449) );
  MUX U9510 ( .IN0(n9449), .IN1(n9442), .SEL(N40), .F(n9450) );
  MUX U9511 ( .IN0(data_mem_out_wire[1499]), .IN1(data_mem_out_wire[1531]), 
        .SEL(N37), .F(n9451) );
  MUX U9512 ( .IN0(data_mem_out_wire[1435]), .IN1(data_mem_out_wire[1467]), 
        .SEL(N37), .F(n9452) );
  MUX U9513 ( .IN0(n9452), .IN1(n9451), .SEL(N38), .F(n9453) );
  MUX U9514 ( .IN0(data_mem_out_wire[1371]), .IN1(data_mem_out_wire[1403]), 
        .SEL(N37), .F(n9454) );
  MUX U9515 ( .IN0(data_mem_out_wire[1307]), .IN1(data_mem_out_wire[1339]), 
        .SEL(N37), .F(n9455) );
  MUX U9516 ( .IN0(n9455), .IN1(n9454), .SEL(N38), .F(n9456) );
  MUX U9517 ( .IN0(n9456), .IN1(n9453), .SEL(N39), .F(n9457) );
  MUX U9518 ( .IN0(data_mem_out_wire[1243]), .IN1(data_mem_out_wire[1275]), 
        .SEL(N37), .F(n9458) );
  MUX U9519 ( .IN0(data_mem_out_wire[1179]), .IN1(data_mem_out_wire[1211]), 
        .SEL(N37), .F(n9459) );
  MUX U9520 ( .IN0(n9459), .IN1(n9458), .SEL(N38), .F(n9460) );
  MUX U9521 ( .IN0(data_mem_out_wire[1115]), .IN1(data_mem_out_wire[1147]), 
        .SEL(N37), .F(n9461) );
  MUX U9522 ( .IN0(data_mem_out_wire[1051]), .IN1(data_mem_out_wire[1083]), 
        .SEL(N37), .F(n9462) );
  MUX U9523 ( .IN0(n9462), .IN1(n9461), .SEL(N38), .F(n9463) );
  MUX U9524 ( .IN0(n9463), .IN1(n9460), .SEL(N39), .F(n9464) );
  MUX U9525 ( .IN0(n9464), .IN1(n9457), .SEL(N40), .F(n9465) );
  MUX U9526 ( .IN0(n9465), .IN1(n9450), .SEL(N41), .F(n9466) );
  MUX U9527 ( .IN0(data_mem_out_wire[987]), .IN1(data_mem_out_wire[1019]), 
        .SEL(N37), .F(n9467) );
  MUX U9528 ( .IN0(data_mem_out_wire[923]), .IN1(data_mem_out_wire[955]), 
        .SEL(N37), .F(n9468) );
  MUX U9529 ( .IN0(n9468), .IN1(n9467), .SEL(N38), .F(n9469) );
  MUX U9530 ( .IN0(data_mem_out_wire[859]), .IN1(data_mem_out_wire[891]), 
        .SEL(N37), .F(n9470) );
  MUX U9531 ( .IN0(data_mem_out_wire[795]), .IN1(data_mem_out_wire[827]), 
        .SEL(N37), .F(n9471) );
  MUX U9532 ( .IN0(n9471), .IN1(n9470), .SEL(N38), .F(n9472) );
  MUX U9533 ( .IN0(n9472), .IN1(n9469), .SEL(N39), .F(n9473) );
  MUX U9534 ( .IN0(data_mem_out_wire[731]), .IN1(data_mem_out_wire[763]), 
        .SEL(N37), .F(n9474) );
  MUX U9535 ( .IN0(data_mem_out_wire[667]), .IN1(data_mem_out_wire[699]), 
        .SEL(N37), .F(n9475) );
  MUX U9536 ( .IN0(n9475), .IN1(n9474), .SEL(N38), .F(n9476) );
  MUX U9537 ( .IN0(data_mem_out_wire[603]), .IN1(data_mem_out_wire[635]), 
        .SEL(N37), .F(n9477) );
  MUX U9538 ( .IN0(data_mem_out_wire[539]), .IN1(data_mem_out_wire[571]), 
        .SEL(N37), .F(n9478) );
  MUX U9539 ( .IN0(n9478), .IN1(n9477), .SEL(N38), .F(n9479) );
  MUX U9540 ( .IN0(n9479), .IN1(n9476), .SEL(N39), .F(n9480) );
  MUX U9541 ( .IN0(n9480), .IN1(n9473), .SEL(N40), .F(n9481) );
  MUX U9542 ( .IN0(data_mem_out_wire[475]), .IN1(data_mem_out_wire[507]), 
        .SEL(N37), .F(n9482) );
  MUX U9543 ( .IN0(data_mem_out_wire[411]), .IN1(data_mem_out_wire[443]), 
        .SEL(N37), .F(n9483) );
  MUX U9544 ( .IN0(n9483), .IN1(n9482), .SEL(N38), .F(n9484) );
  MUX U9545 ( .IN0(data_mem_out_wire[347]), .IN1(data_mem_out_wire[379]), 
        .SEL(N37), .F(n9485) );
  MUX U9546 ( .IN0(data_mem_out_wire[283]), .IN1(data_mem_out_wire[315]), 
        .SEL(N37), .F(n9486) );
  MUX U9547 ( .IN0(n9486), .IN1(n9485), .SEL(N38), .F(n9487) );
  MUX U9548 ( .IN0(n9487), .IN1(n9484), .SEL(N39), .F(n9488) );
  MUX U9549 ( .IN0(data_mem_out_wire[219]), .IN1(data_mem_out_wire[251]), 
        .SEL(N37), .F(n9489) );
  MUX U9550 ( .IN0(data_mem_out_wire[155]), .IN1(data_mem_out_wire[187]), 
        .SEL(N37), .F(n9490) );
  MUX U9551 ( .IN0(n9490), .IN1(n9489), .SEL(N38), .F(n9491) );
  MUX U9552 ( .IN0(data_mem_out_wire[91]), .IN1(data_mem_out_wire[123]), .SEL(
        N37), .F(n9492) );
  MUX U9553 ( .IN0(data_mem_out_wire[27]), .IN1(data_mem_out_wire[59]), .SEL(
        N37), .F(n9493) );
  MUX U9554 ( .IN0(n9493), .IN1(n9492), .SEL(N38), .F(n9494) );
  MUX U9555 ( .IN0(n9494), .IN1(n9491), .SEL(N39), .F(n9495) );
  MUX U9556 ( .IN0(n9495), .IN1(n9488), .SEL(N40), .F(n9496) );
  MUX U9557 ( .IN0(n9496), .IN1(n9481), .SEL(N41), .F(n9497) );
  MUX U9558 ( .IN0(n9497), .IN1(n9466), .SEL(N42), .F(N718) );
  MUX U9559 ( .IN0(data_mem_out_wire[2012]), .IN1(data_mem_out_wire[2044]), 
        .SEL(N37), .F(n9498) );
  MUX U9560 ( .IN0(data_mem_out_wire[1948]), .IN1(data_mem_out_wire[1980]), 
        .SEL(N37), .F(n9499) );
  MUX U9561 ( .IN0(n9499), .IN1(n9498), .SEL(N38), .F(n9500) );
  MUX U9562 ( .IN0(data_mem_out_wire[1884]), .IN1(data_mem_out_wire[1916]), 
        .SEL(N37), .F(n9501) );
  MUX U9563 ( .IN0(data_mem_out_wire[1820]), .IN1(data_mem_out_wire[1852]), 
        .SEL(N37), .F(n9502) );
  MUX U9564 ( .IN0(n9502), .IN1(n9501), .SEL(N38), .F(n9503) );
  MUX U9565 ( .IN0(n9503), .IN1(n9500), .SEL(N39), .F(n9504) );
  MUX U9566 ( .IN0(data_mem_out_wire[1756]), .IN1(data_mem_out_wire[1788]), 
        .SEL(N37), .F(n9505) );
  MUX U9567 ( .IN0(data_mem_out_wire[1692]), .IN1(data_mem_out_wire[1724]), 
        .SEL(N37), .F(n9506) );
  MUX U9568 ( .IN0(n9506), .IN1(n9505), .SEL(N38), .F(n9507) );
  MUX U9569 ( .IN0(data_mem_out_wire[1628]), .IN1(data_mem_out_wire[1660]), 
        .SEL(N37), .F(n9508) );
  MUX U9570 ( .IN0(data_mem_out_wire[1564]), .IN1(data_mem_out_wire[1596]), 
        .SEL(N37), .F(n9509) );
  MUX U9571 ( .IN0(n9509), .IN1(n9508), .SEL(N38), .F(n9510) );
  MUX U9572 ( .IN0(n9510), .IN1(n9507), .SEL(N39), .F(n9511) );
  MUX U9573 ( .IN0(n9511), .IN1(n9504), .SEL(N40), .F(n9512) );
  MUX U9574 ( .IN0(data_mem_out_wire[1500]), .IN1(data_mem_out_wire[1532]), 
        .SEL(N37), .F(n9513) );
  MUX U9575 ( .IN0(data_mem_out_wire[1436]), .IN1(data_mem_out_wire[1468]), 
        .SEL(N37), .F(n9514) );
  MUX U9576 ( .IN0(n9514), .IN1(n9513), .SEL(N38), .F(n9515) );
  MUX U9577 ( .IN0(data_mem_out_wire[1372]), .IN1(data_mem_out_wire[1404]), 
        .SEL(N37), .F(n9516) );
  MUX U9578 ( .IN0(data_mem_out_wire[1308]), .IN1(data_mem_out_wire[1340]), 
        .SEL(N37), .F(n9517) );
  MUX U9579 ( .IN0(n9517), .IN1(n9516), .SEL(N38), .F(n9518) );
  MUX U9580 ( .IN0(n9518), .IN1(n9515), .SEL(N39), .F(n9519) );
  MUX U9581 ( .IN0(data_mem_out_wire[1244]), .IN1(data_mem_out_wire[1276]), 
        .SEL(N37), .F(n9520) );
  MUX U9582 ( .IN0(data_mem_out_wire[1180]), .IN1(data_mem_out_wire[1212]), 
        .SEL(N37), .F(n9521) );
  MUX U9583 ( .IN0(n9521), .IN1(n9520), .SEL(N38), .F(n9522) );
  MUX U9584 ( .IN0(data_mem_out_wire[1116]), .IN1(data_mem_out_wire[1148]), 
        .SEL(N37), .F(n9523) );
  MUX U9585 ( .IN0(data_mem_out_wire[1052]), .IN1(data_mem_out_wire[1084]), 
        .SEL(N37), .F(n9524) );
  MUX U9586 ( .IN0(n9524), .IN1(n9523), .SEL(N38), .F(n9525) );
  MUX U9587 ( .IN0(n9525), .IN1(n9522), .SEL(N39), .F(n9526) );
  MUX U9588 ( .IN0(n9526), .IN1(n9519), .SEL(N40), .F(n9527) );
  MUX U9589 ( .IN0(n9527), .IN1(n9512), .SEL(N41), .F(n9528) );
  MUX U9590 ( .IN0(data_mem_out_wire[988]), .IN1(data_mem_out_wire[1020]), 
        .SEL(N37), .F(n9529) );
  MUX U9591 ( .IN0(data_mem_out_wire[924]), .IN1(data_mem_out_wire[956]), 
        .SEL(N37), .F(n9530) );
  MUX U9592 ( .IN0(n9530), .IN1(n9529), .SEL(N38), .F(n9531) );
  MUX U9593 ( .IN0(data_mem_out_wire[860]), .IN1(data_mem_out_wire[892]), 
        .SEL(N37), .F(n9532) );
  MUX U9594 ( .IN0(data_mem_out_wire[796]), .IN1(data_mem_out_wire[828]), 
        .SEL(N37), .F(n9533) );
  MUX U9595 ( .IN0(n9533), .IN1(n9532), .SEL(N38), .F(n9534) );
  MUX U9596 ( .IN0(n9534), .IN1(n9531), .SEL(N39), .F(n9535) );
  MUX U9597 ( .IN0(data_mem_out_wire[732]), .IN1(data_mem_out_wire[764]), 
        .SEL(N37), .F(n9536) );
  MUX U9598 ( .IN0(data_mem_out_wire[668]), .IN1(data_mem_out_wire[700]), 
        .SEL(N37), .F(n9537) );
  MUX U9599 ( .IN0(n9537), .IN1(n9536), .SEL(N38), .F(n9538) );
  MUX U9600 ( .IN0(data_mem_out_wire[604]), .IN1(data_mem_out_wire[636]), 
        .SEL(N37), .F(n9539) );
  MUX U9601 ( .IN0(data_mem_out_wire[540]), .IN1(data_mem_out_wire[572]), 
        .SEL(N37), .F(n9540) );
  MUX U9602 ( .IN0(n9540), .IN1(n9539), .SEL(N38), .F(n9541) );
  MUX U9603 ( .IN0(n9541), .IN1(n9538), .SEL(N39), .F(n9542) );
  MUX U9604 ( .IN0(n9542), .IN1(n9535), .SEL(N40), .F(n9543) );
  MUX U9605 ( .IN0(data_mem_out_wire[476]), .IN1(data_mem_out_wire[508]), 
        .SEL(N37), .F(n9544) );
  MUX U9606 ( .IN0(data_mem_out_wire[412]), .IN1(data_mem_out_wire[444]), 
        .SEL(N37), .F(n9545) );
  MUX U9607 ( .IN0(n9545), .IN1(n9544), .SEL(N38), .F(n9546) );
  MUX U9608 ( .IN0(data_mem_out_wire[348]), .IN1(data_mem_out_wire[380]), 
        .SEL(N37), .F(n9547) );
  MUX U9609 ( .IN0(data_mem_out_wire[284]), .IN1(data_mem_out_wire[316]), 
        .SEL(N37), .F(n9548) );
  MUX U9610 ( .IN0(n9548), .IN1(n9547), .SEL(N38), .F(n9549) );
  MUX U9611 ( .IN0(n9549), .IN1(n9546), .SEL(N39), .F(n9550) );
  MUX U9612 ( .IN0(data_mem_out_wire[220]), .IN1(data_mem_out_wire[252]), 
        .SEL(N37), .F(n9551) );
  MUX U9613 ( .IN0(data_mem_out_wire[156]), .IN1(data_mem_out_wire[188]), 
        .SEL(N37), .F(n9552) );
  MUX U9614 ( .IN0(n9552), .IN1(n9551), .SEL(N38), .F(n9553) );
  MUX U9615 ( .IN0(data_mem_out_wire[92]), .IN1(data_mem_out_wire[124]), .SEL(
        N37), .F(n9554) );
  MUX U9616 ( .IN0(data_mem_out_wire[28]), .IN1(data_mem_out_wire[60]), .SEL(
        N37), .F(n9555) );
  MUX U9617 ( .IN0(n9555), .IN1(n9554), .SEL(N38), .F(n9556) );
  MUX U9618 ( .IN0(n9556), .IN1(n9553), .SEL(N39), .F(n9557) );
  MUX U9619 ( .IN0(n9557), .IN1(n9550), .SEL(N40), .F(n9558) );
  MUX U9620 ( .IN0(n9558), .IN1(n9543), .SEL(N41), .F(n9559) );
  MUX U9621 ( .IN0(n9559), .IN1(n9528), .SEL(N42), .F(N717) );
  MUX U9622 ( .IN0(data_mem_out_wire[2013]), .IN1(data_mem_out_wire[2045]), 
        .SEL(N37), .F(n9560) );
  MUX U9623 ( .IN0(data_mem_out_wire[1949]), .IN1(data_mem_out_wire[1981]), 
        .SEL(N37), .F(n9561) );
  MUX U9624 ( .IN0(n9561), .IN1(n9560), .SEL(N38), .F(n9562) );
  MUX U9625 ( .IN0(data_mem_out_wire[1885]), .IN1(data_mem_out_wire[1917]), 
        .SEL(N37), .F(n9563) );
  MUX U9626 ( .IN0(data_mem_out_wire[1821]), .IN1(data_mem_out_wire[1853]), 
        .SEL(N37), .F(n9564) );
  MUX U9627 ( .IN0(n9564), .IN1(n9563), .SEL(N38), .F(n9565) );
  MUX U9628 ( .IN0(n9565), .IN1(n9562), .SEL(N39), .F(n9566) );
  MUX U9629 ( .IN0(data_mem_out_wire[1757]), .IN1(data_mem_out_wire[1789]), 
        .SEL(N37), .F(n9567) );
  MUX U9630 ( .IN0(data_mem_out_wire[1693]), .IN1(data_mem_out_wire[1725]), 
        .SEL(N37), .F(n9568) );
  MUX U9631 ( .IN0(n9568), .IN1(n9567), .SEL(N38), .F(n9569) );
  MUX U9632 ( .IN0(data_mem_out_wire[1629]), .IN1(data_mem_out_wire[1661]), 
        .SEL(N37), .F(n9570) );
  MUX U9633 ( .IN0(data_mem_out_wire[1565]), .IN1(data_mem_out_wire[1597]), 
        .SEL(N37), .F(n9571) );
  MUX U9634 ( .IN0(n9571), .IN1(n9570), .SEL(N38), .F(n9572) );
  MUX U9635 ( .IN0(n9572), .IN1(n9569), .SEL(N39), .F(n9573) );
  MUX U9636 ( .IN0(n9573), .IN1(n9566), .SEL(N40), .F(n9574) );
  MUX U9637 ( .IN0(data_mem_out_wire[1501]), .IN1(data_mem_out_wire[1533]), 
        .SEL(N37), .F(n9575) );
  MUX U9638 ( .IN0(data_mem_out_wire[1437]), .IN1(data_mem_out_wire[1469]), 
        .SEL(N37), .F(n9576) );
  MUX U9639 ( .IN0(n9576), .IN1(n9575), .SEL(N38), .F(n9577) );
  MUX U9640 ( .IN0(data_mem_out_wire[1373]), .IN1(data_mem_out_wire[1405]), 
        .SEL(N37), .F(n9578) );
  MUX U9641 ( .IN0(data_mem_out_wire[1309]), .IN1(data_mem_out_wire[1341]), 
        .SEL(N37), .F(n9579) );
  MUX U9642 ( .IN0(n9579), .IN1(n9578), .SEL(N38), .F(n9580) );
  MUX U9643 ( .IN0(n9580), .IN1(n9577), .SEL(N39), .F(n9581) );
  MUX U9644 ( .IN0(data_mem_out_wire[1245]), .IN1(data_mem_out_wire[1277]), 
        .SEL(N37), .F(n9582) );
  MUX U9645 ( .IN0(data_mem_out_wire[1181]), .IN1(data_mem_out_wire[1213]), 
        .SEL(N37), .F(n9583) );
  MUX U9646 ( .IN0(n9583), .IN1(n9582), .SEL(N38), .F(n9584) );
  MUX U9647 ( .IN0(data_mem_out_wire[1117]), .IN1(data_mem_out_wire[1149]), 
        .SEL(N37), .F(n9585) );
  MUX U9648 ( .IN0(data_mem_out_wire[1053]), .IN1(data_mem_out_wire[1085]), 
        .SEL(N37), .F(n9586) );
  MUX U9649 ( .IN0(n9586), .IN1(n9585), .SEL(N38), .F(n9587) );
  MUX U9650 ( .IN0(n9587), .IN1(n9584), .SEL(N39), .F(n9588) );
  MUX U9651 ( .IN0(n9588), .IN1(n9581), .SEL(N40), .F(n9589) );
  MUX U9652 ( .IN0(n9589), .IN1(n9574), .SEL(N41), .F(n9590) );
  MUX U9653 ( .IN0(data_mem_out_wire[989]), .IN1(data_mem_out_wire[1021]), 
        .SEL(N37), .F(n9591) );
  MUX U9654 ( .IN0(data_mem_out_wire[925]), .IN1(data_mem_out_wire[957]), 
        .SEL(N37), .F(n9592) );
  MUX U9655 ( .IN0(n9592), .IN1(n9591), .SEL(N38), .F(n9593) );
  MUX U9656 ( .IN0(data_mem_out_wire[861]), .IN1(data_mem_out_wire[893]), 
        .SEL(N37), .F(n9594) );
  MUX U9657 ( .IN0(data_mem_out_wire[797]), .IN1(data_mem_out_wire[829]), 
        .SEL(N37), .F(n9595) );
  MUX U9658 ( .IN0(n9595), .IN1(n9594), .SEL(N38), .F(n9596) );
  MUX U9659 ( .IN0(n9596), .IN1(n9593), .SEL(N39), .F(n9597) );
  MUX U9660 ( .IN0(data_mem_out_wire[733]), .IN1(data_mem_out_wire[765]), 
        .SEL(N37), .F(n9598) );
  MUX U9661 ( .IN0(data_mem_out_wire[669]), .IN1(data_mem_out_wire[701]), 
        .SEL(N37), .F(n9599) );
  MUX U9662 ( .IN0(n9599), .IN1(n9598), .SEL(N38), .F(n9600) );
  MUX U9663 ( .IN0(data_mem_out_wire[605]), .IN1(data_mem_out_wire[637]), 
        .SEL(N37), .F(n9601) );
  MUX U9664 ( .IN0(data_mem_out_wire[541]), .IN1(data_mem_out_wire[573]), 
        .SEL(N37), .F(n9602) );
  MUX U9665 ( .IN0(n9602), .IN1(n9601), .SEL(N38), .F(n9603) );
  MUX U9666 ( .IN0(n9603), .IN1(n9600), .SEL(N39), .F(n9604) );
  MUX U9667 ( .IN0(n9604), .IN1(n9597), .SEL(N40), .F(n9605) );
  MUX U9668 ( .IN0(data_mem_out_wire[477]), .IN1(data_mem_out_wire[509]), 
        .SEL(N37), .F(n9606) );
  MUX U9669 ( .IN0(data_mem_out_wire[413]), .IN1(data_mem_out_wire[445]), 
        .SEL(N37), .F(n9607) );
  MUX U9670 ( .IN0(n9607), .IN1(n9606), .SEL(N38), .F(n9608) );
  MUX U9671 ( .IN0(data_mem_out_wire[349]), .IN1(data_mem_out_wire[381]), 
        .SEL(N37), .F(n9609) );
  MUX U9672 ( .IN0(data_mem_out_wire[285]), .IN1(data_mem_out_wire[317]), 
        .SEL(N37), .F(n9610) );
  MUX U9673 ( .IN0(n9610), .IN1(n9609), .SEL(N38), .F(n9611) );
  MUX U9674 ( .IN0(n9611), .IN1(n9608), .SEL(N39), .F(n9612) );
  MUX U9675 ( .IN0(data_mem_out_wire[221]), .IN1(data_mem_out_wire[253]), 
        .SEL(N37), .F(n9613) );
  MUX U9676 ( .IN0(data_mem_out_wire[157]), .IN1(data_mem_out_wire[189]), 
        .SEL(N37), .F(n9614) );
  MUX U9677 ( .IN0(n9614), .IN1(n9613), .SEL(N38), .F(n9615) );
  MUX U9678 ( .IN0(data_mem_out_wire[93]), .IN1(data_mem_out_wire[125]), .SEL(
        N37), .F(n9616) );
  MUX U9679 ( .IN0(data_mem_out_wire[29]), .IN1(data_mem_out_wire[61]), .SEL(
        N37), .F(n9617) );
  MUX U9680 ( .IN0(n9617), .IN1(n9616), .SEL(N38), .F(n9618) );
  MUX U9681 ( .IN0(n9618), .IN1(n9615), .SEL(N39), .F(n9619) );
  MUX U9682 ( .IN0(n9619), .IN1(n9612), .SEL(N40), .F(n9620) );
  MUX U9683 ( .IN0(n9620), .IN1(n9605), .SEL(N41), .F(n9621) );
  MUX U9684 ( .IN0(n9621), .IN1(n9590), .SEL(N42), .F(N716) );
  MUX U9685 ( .IN0(data_mem_out_wire[2014]), .IN1(data_mem_out_wire[2046]), 
        .SEL(N37), .F(n9622) );
  MUX U9686 ( .IN0(data_mem_out_wire[1950]), .IN1(data_mem_out_wire[1982]), 
        .SEL(N37), .F(n9623) );
  MUX U9687 ( .IN0(n9623), .IN1(n9622), .SEL(N38), .F(n9624) );
  MUX U9688 ( .IN0(data_mem_out_wire[1886]), .IN1(data_mem_out_wire[1918]), 
        .SEL(N37), .F(n9625) );
  MUX U9689 ( .IN0(data_mem_out_wire[1822]), .IN1(data_mem_out_wire[1854]), 
        .SEL(N37), .F(n9626) );
  MUX U9690 ( .IN0(n9626), .IN1(n9625), .SEL(N38), .F(n9627) );
  MUX U9691 ( .IN0(n9627), .IN1(n9624), .SEL(N39), .F(n9628) );
  MUX U9692 ( .IN0(data_mem_out_wire[1758]), .IN1(data_mem_out_wire[1790]), 
        .SEL(N37), .F(n9629) );
  MUX U9693 ( .IN0(data_mem_out_wire[1694]), .IN1(data_mem_out_wire[1726]), 
        .SEL(N37), .F(n9630) );
  MUX U9694 ( .IN0(n9630), .IN1(n9629), .SEL(N38), .F(n9631) );
  MUX U9695 ( .IN0(data_mem_out_wire[1630]), .IN1(data_mem_out_wire[1662]), 
        .SEL(N37), .F(n9632) );
  MUX U9696 ( .IN0(data_mem_out_wire[1566]), .IN1(data_mem_out_wire[1598]), 
        .SEL(N37), .F(n9633) );
  MUX U9697 ( .IN0(n9633), .IN1(n9632), .SEL(N38), .F(n9634) );
  MUX U9698 ( .IN0(n9634), .IN1(n9631), .SEL(N39), .F(n9635) );
  MUX U9699 ( .IN0(n9635), .IN1(n9628), .SEL(N40), .F(n9636) );
  MUX U9700 ( .IN0(data_mem_out_wire[1502]), .IN1(data_mem_out_wire[1534]), 
        .SEL(N37), .F(n9637) );
  MUX U9701 ( .IN0(data_mem_out_wire[1438]), .IN1(data_mem_out_wire[1470]), 
        .SEL(N37), .F(n9638) );
  MUX U9702 ( .IN0(n9638), .IN1(n9637), .SEL(N38), .F(n9639) );
  MUX U9703 ( .IN0(data_mem_out_wire[1374]), .IN1(data_mem_out_wire[1406]), 
        .SEL(N37), .F(n9640) );
  MUX U9704 ( .IN0(data_mem_out_wire[1310]), .IN1(data_mem_out_wire[1342]), 
        .SEL(N37), .F(n9641) );
  MUX U9705 ( .IN0(n9641), .IN1(n9640), .SEL(N38), .F(n9642) );
  MUX U9706 ( .IN0(n9642), .IN1(n9639), .SEL(N39), .F(n9643) );
  MUX U9707 ( .IN0(data_mem_out_wire[1246]), .IN1(data_mem_out_wire[1278]), 
        .SEL(N37), .F(n9644) );
  MUX U9708 ( .IN0(data_mem_out_wire[1182]), .IN1(data_mem_out_wire[1214]), 
        .SEL(N37), .F(n9645) );
  MUX U9709 ( .IN0(n9645), .IN1(n9644), .SEL(N38), .F(n9646) );
  MUX U9710 ( .IN0(data_mem_out_wire[1118]), .IN1(data_mem_out_wire[1150]), 
        .SEL(N37), .F(n9647) );
  MUX U9711 ( .IN0(data_mem_out_wire[1054]), .IN1(data_mem_out_wire[1086]), 
        .SEL(N37), .F(n9648) );
  MUX U9712 ( .IN0(n9648), .IN1(n9647), .SEL(N38), .F(n9649) );
  MUX U9713 ( .IN0(n9649), .IN1(n9646), .SEL(N39), .F(n9650) );
  MUX U9714 ( .IN0(n9650), .IN1(n9643), .SEL(N40), .F(n9651) );
  MUX U9715 ( .IN0(n9651), .IN1(n9636), .SEL(N41), .F(n9652) );
  MUX U9716 ( .IN0(data_mem_out_wire[990]), .IN1(data_mem_out_wire[1022]), 
        .SEL(N37), .F(n9653) );
  MUX U9717 ( .IN0(data_mem_out_wire[926]), .IN1(data_mem_out_wire[958]), 
        .SEL(N37), .F(n9654) );
  MUX U9718 ( .IN0(n9654), .IN1(n9653), .SEL(N38), .F(n9655) );
  MUX U9719 ( .IN0(data_mem_out_wire[862]), .IN1(data_mem_out_wire[894]), 
        .SEL(N37), .F(n9656) );
  MUX U9720 ( .IN0(data_mem_out_wire[798]), .IN1(data_mem_out_wire[830]), 
        .SEL(N37), .F(n9657) );
  MUX U9721 ( .IN0(n9657), .IN1(n9656), .SEL(N38), .F(n9658) );
  MUX U9722 ( .IN0(n9658), .IN1(n9655), .SEL(N39), .F(n9659) );
  MUX U9723 ( .IN0(data_mem_out_wire[734]), .IN1(data_mem_out_wire[766]), 
        .SEL(N37), .F(n9660) );
  MUX U9724 ( .IN0(data_mem_out_wire[670]), .IN1(data_mem_out_wire[702]), 
        .SEL(N37), .F(n9661) );
  MUX U9725 ( .IN0(n9661), .IN1(n9660), .SEL(N38), .F(n9662) );
  MUX U9726 ( .IN0(data_mem_out_wire[606]), .IN1(data_mem_out_wire[638]), 
        .SEL(N37), .F(n9663) );
  MUX U9727 ( .IN0(data_mem_out_wire[542]), .IN1(data_mem_out_wire[574]), 
        .SEL(N37), .F(n9664) );
  MUX U9728 ( .IN0(n9664), .IN1(n9663), .SEL(N38), .F(n9665) );
  MUX U9729 ( .IN0(n9665), .IN1(n9662), .SEL(N39), .F(n9666) );
  MUX U9730 ( .IN0(n9666), .IN1(n9659), .SEL(N40), .F(n9667) );
  MUX U9731 ( .IN0(data_mem_out_wire[478]), .IN1(data_mem_out_wire[510]), 
        .SEL(N37), .F(n9668) );
  MUX U9732 ( .IN0(data_mem_out_wire[414]), .IN1(data_mem_out_wire[446]), 
        .SEL(N37), .F(n9669) );
  MUX U9733 ( .IN0(n9669), .IN1(n9668), .SEL(N38), .F(n9670) );
  MUX U9734 ( .IN0(data_mem_out_wire[350]), .IN1(data_mem_out_wire[382]), 
        .SEL(N37), .F(n9671) );
  MUX U9735 ( .IN0(data_mem_out_wire[286]), .IN1(data_mem_out_wire[318]), 
        .SEL(N37), .F(n9672) );
  MUX U9736 ( .IN0(n9672), .IN1(n9671), .SEL(N38), .F(n9673) );
  MUX U9737 ( .IN0(n9673), .IN1(n9670), .SEL(N39), .F(n9674) );
  MUX U9738 ( .IN0(data_mem_out_wire[222]), .IN1(data_mem_out_wire[254]), 
        .SEL(N37), .F(n9675) );
  MUX U9739 ( .IN0(data_mem_out_wire[158]), .IN1(data_mem_out_wire[190]), 
        .SEL(N37), .F(n9676) );
  MUX U9740 ( .IN0(n9676), .IN1(n9675), .SEL(N38), .F(n9677) );
  MUX U9741 ( .IN0(data_mem_out_wire[94]), .IN1(data_mem_out_wire[126]), .SEL(
        N37), .F(n9678) );
  MUX U9742 ( .IN0(data_mem_out_wire[30]), .IN1(data_mem_out_wire[62]), .SEL(
        N37), .F(n9679) );
  MUX U9743 ( .IN0(n9679), .IN1(n9678), .SEL(N38), .F(n9680) );
  MUX U9744 ( .IN0(n9680), .IN1(n9677), .SEL(N39), .F(n9681) );
  MUX U9745 ( .IN0(n9681), .IN1(n9674), .SEL(N40), .F(n9682) );
  MUX U9746 ( .IN0(n9682), .IN1(n9667), .SEL(N41), .F(n9683) );
  MUX U9747 ( .IN0(n9683), .IN1(n9652), .SEL(N42), .F(N715) );
  MUX U9748 ( .IN0(data_mem_out_wire[2015]), .IN1(data_mem_out_wire[2047]), 
        .SEL(N37), .F(n9684) );
  MUX U9749 ( .IN0(data_mem_out_wire[1951]), .IN1(data_mem_out_wire[1983]), 
        .SEL(N37), .F(n9685) );
  MUX U9750 ( .IN0(n9685), .IN1(n9684), .SEL(N38), .F(n9686) );
  MUX U9751 ( .IN0(data_mem_out_wire[1887]), .IN1(data_mem_out_wire[1919]), 
        .SEL(N37), .F(n9687) );
  MUX U9752 ( .IN0(data_mem_out_wire[1823]), .IN1(data_mem_out_wire[1855]), 
        .SEL(N37), .F(n9688) );
  MUX U9753 ( .IN0(n9688), .IN1(n9687), .SEL(N38), .F(n9689) );
  MUX U9754 ( .IN0(n9689), .IN1(n9686), .SEL(N39), .F(n9690) );
  MUX U9755 ( .IN0(data_mem_out_wire[1759]), .IN1(data_mem_out_wire[1791]), 
        .SEL(N37), .F(n9691) );
  MUX U9756 ( .IN0(data_mem_out_wire[1695]), .IN1(data_mem_out_wire[1727]), 
        .SEL(N37), .F(n9692) );
  MUX U9757 ( .IN0(n9692), .IN1(n9691), .SEL(N38), .F(n9693) );
  MUX U9758 ( .IN0(data_mem_out_wire[1631]), .IN1(data_mem_out_wire[1663]), 
        .SEL(N37), .F(n9694) );
  MUX U9759 ( .IN0(data_mem_out_wire[1567]), .IN1(data_mem_out_wire[1599]), 
        .SEL(N37), .F(n9695) );
  MUX U9760 ( .IN0(n9695), .IN1(n9694), .SEL(N38), .F(n9696) );
  MUX U9761 ( .IN0(n9696), .IN1(n9693), .SEL(N39), .F(n9697) );
  MUX U9762 ( .IN0(n9697), .IN1(n9690), .SEL(N40), .F(n9698) );
  MUX U9763 ( .IN0(data_mem_out_wire[1503]), .IN1(data_mem_out_wire[1535]), 
        .SEL(N37), .F(n9699) );
  MUX U9764 ( .IN0(data_mem_out_wire[1439]), .IN1(data_mem_out_wire[1471]), 
        .SEL(N37), .F(n9700) );
  MUX U9765 ( .IN0(n9700), .IN1(n9699), .SEL(N38), .F(n9701) );
  MUX U9766 ( .IN0(data_mem_out_wire[1375]), .IN1(data_mem_out_wire[1407]), 
        .SEL(N37), .F(n9702) );
  MUX U9767 ( .IN0(data_mem_out_wire[1311]), .IN1(data_mem_out_wire[1343]), 
        .SEL(N37), .F(n9703) );
  MUX U9768 ( .IN0(n9703), .IN1(n9702), .SEL(N38), .F(n9704) );
  MUX U9769 ( .IN0(n9704), .IN1(n9701), .SEL(N39), .F(n9705) );
  MUX U9770 ( .IN0(data_mem_out_wire[1247]), .IN1(data_mem_out_wire[1279]), 
        .SEL(N37), .F(n9706) );
  MUX U9771 ( .IN0(data_mem_out_wire[1183]), .IN1(data_mem_out_wire[1215]), 
        .SEL(N37), .F(n9707) );
  MUX U9772 ( .IN0(n9707), .IN1(n9706), .SEL(N38), .F(n9708) );
  MUX U9773 ( .IN0(data_mem_out_wire[1119]), .IN1(data_mem_out_wire[1151]), 
        .SEL(N37), .F(n9709) );
  MUX U9774 ( .IN0(data_mem_out_wire[1055]), .IN1(data_mem_out_wire[1087]), 
        .SEL(N37), .F(n9710) );
  MUX U9775 ( .IN0(n9710), .IN1(n9709), .SEL(N38), .F(n9711) );
  MUX U9776 ( .IN0(n9711), .IN1(n9708), .SEL(N39), .F(n9712) );
  MUX U9777 ( .IN0(n9712), .IN1(n9705), .SEL(N40), .F(n9713) );
  MUX U9778 ( .IN0(n9713), .IN1(n9698), .SEL(N41), .F(n9714) );
  MUX U9779 ( .IN0(data_mem_out_wire[991]), .IN1(data_mem_out_wire[1023]), 
        .SEL(N37), .F(n9715) );
  MUX U9780 ( .IN0(data_mem_out_wire[927]), .IN1(data_mem_out_wire[959]), 
        .SEL(N37), .F(n9716) );
  MUX U9781 ( .IN0(n9716), .IN1(n9715), .SEL(N38), .F(n9717) );
  MUX U9782 ( .IN0(data_mem_out_wire[863]), .IN1(data_mem_out_wire[895]), 
        .SEL(N37), .F(n9718) );
  MUX U9783 ( .IN0(data_mem_out_wire[799]), .IN1(data_mem_out_wire[831]), 
        .SEL(N37), .F(n9719) );
  MUX U9784 ( .IN0(n9719), .IN1(n9718), .SEL(N38), .F(n9720) );
  MUX U9785 ( .IN0(n9720), .IN1(n9717), .SEL(N39), .F(n9721) );
  MUX U9786 ( .IN0(data_mem_out_wire[735]), .IN1(data_mem_out_wire[767]), 
        .SEL(N37), .F(n9722) );
  MUX U9787 ( .IN0(data_mem_out_wire[671]), .IN1(data_mem_out_wire[703]), 
        .SEL(N37), .F(n9723) );
  MUX U9788 ( .IN0(n9723), .IN1(n9722), .SEL(N38), .F(n9724) );
  MUX U9789 ( .IN0(data_mem_out_wire[607]), .IN1(data_mem_out_wire[639]), 
        .SEL(N37), .F(n9725) );
  MUX U9790 ( .IN0(data_mem_out_wire[543]), .IN1(data_mem_out_wire[575]), 
        .SEL(N37), .F(n9726) );
  MUX U9791 ( .IN0(n9726), .IN1(n9725), .SEL(N38), .F(n9727) );
  MUX U9792 ( .IN0(n9727), .IN1(n9724), .SEL(N39), .F(n9728) );
  MUX U9793 ( .IN0(n9728), .IN1(n9721), .SEL(N40), .F(n9729) );
  MUX U9794 ( .IN0(data_mem_out_wire[479]), .IN1(data_mem_out_wire[511]), 
        .SEL(N37), .F(n9730) );
  MUX U9795 ( .IN0(data_mem_out_wire[415]), .IN1(data_mem_out_wire[447]), 
        .SEL(N37), .F(n9731) );
  MUX U9796 ( .IN0(n9731), .IN1(n9730), .SEL(N38), .F(n9732) );
  MUX U9797 ( .IN0(data_mem_out_wire[351]), .IN1(data_mem_out_wire[383]), 
        .SEL(N37), .F(n9733) );
  MUX U9798 ( .IN0(data_mem_out_wire[287]), .IN1(data_mem_out_wire[319]), 
        .SEL(N37), .F(n9734) );
  MUX U9799 ( .IN0(n9734), .IN1(n9733), .SEL(N38), .F(n9735) );
  MUX U9800 ( .IN0(n9735), .IN1(n9732), .SEL(N39), .F(n9736) );
  MUX U9801 ( .IN0(data_mem_out_wire[223]), .IN1(data_mem_out_wire[255]), 
        .SEL(N37), .F(n9737) );
  MUX U9802 ( .IN0(data_mem_out_wire[159]), .IN1(data_mem_out_wire[191]), 
        .SEL(N37), .F(n9738) );
  MUX U9803 ( .IN0(n9738), .IN1(n9737), .SEL(N38), .F(n9739) );
  MUX U9804 ( .IN0(data_mem_out_wire[95]), .IN1(data_mem_out_wire[127]), .SEL(
        N37), .F(n9740) );
  MUX U9805 ( .IN0(data_mem_out_wire[31]), .IN1(data_mem_out_wire[63]), .SEL(
        N37), .F(n9741) );
  MUX U9806 ( .IN0(n9741), .IN1(n9740), .SEL(N38), .F(n9742) );
  MUX U9807 ( .IN0(n9742), .IN1(n9739), .SEL(N39), .F(n9743) );
  MUX U9808 ( .IN0(n9743), .IN1(n9736), .SEL(N40), .F(n9744) );
  MUX U9809 ( .IN0(n9744), .IN1(n9729), .SEL(N41), .F(n9745) );
  MUX U9810 ( .IN0(n9745), .IN1(n9714), .SEL(N42), .F(N714) );
  MUX U9811 ( .IN0(n9746), .IN1(data_mem_out_wire[31]), .SEL(n9747), .F(n7761)
         );
  MUX U9812 ( .IN0(n9748), .IN1(data_mem_out_wire[30]), .SEL(n9747), .F(n7760)
         );
  MUX U9813 ( .IN0(n9749), .IN1(data_mem_out_wire[29]), .SEL(n9747), .F(n7759)
         );
  MUX U9814 ( .IN0(n9750), .IN1(data_mem_out_wire[28]), .SEL(n9747), .F(n7758)
         );
  MUX U9815 ( .IN0(n9751), .IN1(data_mem_out_wire[27]), .SEL(n9747), .F(n7757)
         );
  MUX U9816 ( .IN0(n9752), .IN1(data_mem_out_wire[26]), .SEL(n9747), .F(n7756)
         );
  MUX U9817 ( .IN0(n9753), .IN1(data_mem_out_wire[25]), .SEL(n9747), .F(n7755)
         );
  MUX U9818 ( .IN0(n9754), .IN1(data_mem_out_wire[24]), .SEL(n9747), .F(n7754)
         );
  AND U9819 ( .A(n9755), .B(n9756), .Z(n9747) );
  ANDN U9820 ( .B(n9757), .A(n9758), .Z(n9755) );
  OR U9821 ( .A(n9759), .B(n9760), .Z(n9757) );
  MUX U9822 ( .IN0(data_mem_out_wire[23]), .IN1(n9761), .SEL(n9762), .F(n7753)
         );
  MUX U9823 ( .IN0(data_mem_out_wire[22]), .IN1(n9763), .SEL(n9762), .F(n7752)
         );
  MUX U9824 ( .IN0(data_mem_out_wire[21]), .IN1(n9764), .SEL(n9762), .F(n7751)
         );
  MUX U9825 ( .IN0(data_mem_out_wire[20]), .IN1(n9765), .SEL(n9762), .F(n7750)
         );
  MUX U9826 ( .IN0(data_mem_out_wire[19]), .IN1(n9766), .SEL(n9762), .F(n7749)
         );
  IV U9827 ( .A(n9767), .Z(n9762) );
  MUX U9828 ( .IN0(n9768), .IN1(data_mem_out_wire[18]), .SEL(n9767), .F(n7748)
         );
  MUX U9829 ( .IN0(n9769), .IN1(data_mem_out_wire[17]), .SEL(n9767), .F(n7747)
         );
  MUX U9830 ( .IN0(n9770), .IN1(data_mem_out_wire[16]), .SEL(n9767), .F(n7746)
         );
  AND U9831 ( .A(n9771), .B(n9772), .Z(n9767) );
  OR U9832 ( .A(n9759), .B(n9773), .Z(n9772) );
  ANDN U9833 ( .B(n9756), .A(n9758), .Z(n9771) );
  AND U9834 ( .A(n9774), .B(addr[1]), .Z(n9758) );
  ANDN U9835 ( .B(n9775), .A(n9759), .Z(n9774) );
  MUX U9836 ( .IN0(data_mem_out_wire[15]), .IN1(n9776), .SEL(n9777), .F(n7745)
         );
  MUX U9837 ( .IN0(data_mem_out_wire[14]), .IN1(n9778), .SEL(n9777), .F(n7744)
         );
  MUX U9838 ( .IN0(data_mem_out_wire[13]), .IN1(n9779), .SEL(n9777), .F(n7743)
         );
  MUX U9839 ( .IN0(data_mem_out_wire[12]), .IN1(n9780), .SEL(n9777), .F(n7742)
         );
  MUX U9840 ( .IN0(data_mem_out_wire[11]), .IN1(n9781), .SEL(n9777), .F(n7741)
         );
  IV U9841 ( .A(n9782), .Z(n9777) );
  MUX U9842 ( .IN0(n9783), .IN1(data_mem_out_wire[10]), .SEL(n9782), .F(n7740)
         );
  MUX U9843 ( .IN0(n9784), .IN1(data_mem_out_wire[9]), .SEL(n9782), .F(n7739)
         );
  MUX U9844 ( .IN0(n9785), .IN1(data_mem_out_wire[8]), .SEL(n9782), .F(n7738)
         );
  AND U9845 ( .A(n9786), .B(n9787), .Z(n9782) );
  OR U9846 ( .A(n9759), .B(n9788), .Z(n9787) );
  MUX U9847 ( .IN0(data_mem_out_wire[7]), .IN1(data_in[7]), .SEL(n9789), .F(
        n7737) );
  MUX U9848 ( .IN0(data_mem_out_wire[6]), .IN1(data_in[6]), .SEL(n9789), .F(
        n7736) );
  MUX U9849 ( .IN0(data_mem_out_wire[5]), .IN1(data_in[5]), .SEL(n9789), .F(
        n7735) );
  MUX U9850 ( .IN0(data_mem_out_wire[4]), .IN1(data_in[4]), .SEL(n9789), .F(
        n7734) );
  MUX U9851 ( .IN0(data_mem_out_wire[3]), .IN1(data_in[3]), .SEL(n9789), .F(
        n7733) );
  IV U9852 ( .A(n9790), .Z(n9789) );
  MUX U9853 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[2]), .SEL(n9790), .F(
        n7732) );
  MUX U9854 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1]), .SEL(n9790), .F(
        n7731) );
  MUX U9855 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[0]), .SEL(n9790), .F(
        n7730) );
  AND U9856 ( .A(n9786), .B(n9791), .Z(n9790) );
  NANDN U9857 ( .A(n9759), .B(n9792), .Z(n9791) );
  ANDN U9858 ( .B(n9756), .A(n9793), .Z(n9786) );
  AND U9859 ( .A(n9794), .B(n9775), .Z(n9793) );
  ANDN U9860 ( .B(n9795), .A(n9759), .Z(n9794) );
  NANDN U9861 ( .A(n9759), .B(n9796), .Z(n9756) );
  NAND U9862 ( .A(n9797), .B(n9798), .Z(n9759) );
  MUX U9863 ( .IN0(n9746), .IN1(data_mem_out_wire[63]), .SEL(n9799), .F(n7729)
         );
  MUX U9864 ( .IN0(n9748), .IN1(data_mem_out_wire[62]), .SEL(n9799), .F(n7728)
         );
  MUX U9865 ( .IN0(n9749), .IN1(data_mem_out_wire[61]), .SEL(n9799), .F(n7727)
         );
  MUX U9866 ( .IN0(n9750), .IN1(data_mem_out_wire[60]), .SEL(n9799), .F(n7726)
         );
  MUX U9867 ( .IN0(n9751), .IN1(data_mem_out_wire[59]), .SEL(n9799), .F(n7725)
         );
  MUX U9868 ( .IN0(n9752), .IN1(data_mem_out_wire[58]), .SEL(n9799), .F(n7724)
         );
  MUX U9869 ( .IN0(n9753), .IN1(data_mem_out_wire[57]), .SEL(n9799), .F(n7723)
         );
  MUX U9870 ( .IN0(n9754), .IN1(data_mem_out_wire[56]), .SEL(n9799), .F(n7722)
         );
  AND U9871 ( .A(n9800), .B(n9801), .Z(n9799) );
  AND U9872 ( .A(n9802), .B(n9803), .Z(n9800) );
  OR U9873 ( .A(n9760), .B(n9804), .Z(n9803) );
  MUX U9874 ( .IN0(data_mem_out_wire[55]), .IN1(n9761), .SEL(n9805), .F(n7721)
         );
  MUX U9875 ( .IN0(data_mem_out_wire[54]), .IN1(n9763), .SEL(n9805), .F(n7720)
         );
  MUX U9876 ( .IN0(data_mem_out_wire[53]), .IN1(n9764), .SEL(n9805), .F(n7719)
         );
  MUX U9877 ( .IN0(data_mem_out_wire[52]), .IN1(n9765), .SEL(n9805), .F(n7718)
         );
  MUX U9878 ( .IN0(data_mem_out_wire[51]), .IN1(n9766), .SEL(n9805), .F(n7717)
         );
  IV U9879 ( .A(n9806), .Z(n9805) );
  MUX U9880 ( .IN0(n9768), .IN1(data_mem_out_wire[50]), .SEL(n9806), .F(n7716)
         );
  MUX U9881 ( .IN0(n9769), .IN1(data_mem_out_wire[49]), .SEL(n9806), .F(n7715)
         );
  MUX U9882 ( .IN0(n9770), .IN1(data_mem_out_wire[48]), .SEL(n9806), .F(n7714)
         );
  AND U9883 ( .A(n9807), .B(n9808), .Z(n9806) );
  OR U9884 ( .A(n9773), .B(n9804), .Z(n9808) );
  AND U9885 ( .A(n9802), .B(n9801), .Z(n9807) );
  NANDN U9886 ( .A(n9804), .B(n9809), .Z(n9802) );
  MUX U9887 ( .IN0(data_mem_out_wire[47]), .IN1(n9776), .SEL(n9810), .F(n7713)
         );
  MUX U9888 ( .IN0(data_mem_out_wire[46]), .IN1(n9778), .SEL(n9810), .F(n7712)
         );
  MUX U9889 ( .IN0(data_mem_out_wire[45]), .IN1(n9779), .SEL(n9810), .F(n7711)
         );
  MUX U9890 ( .IN0(data_mem_out_wire[44]), .IN1(n9780), .SEL(n9810), .F(n7710)
         );
  MUX U9891 ( .IN0(data_mem_out_wire[43]), .IN1(n9781), .SEL(n9810), .F(n7709)
         );
  IV U9892 ( .A(n9811), .Z(n9810) );
  MUX U9893 ( .IN0(n9783), .IN1(data_mem_out_wire[42]), .SEL(n9811), .F(n7708)
         );
  MUX U9894 ( .IN0(n9784), .IN1(data_mem_out_wire[41]), .SEL(n9811), .F(n7707)
         );
  MUX U9895 ( .IN0(n9785), .IN1(data_mem_out_wire[40]), .SEL(n9811), .F(n7706)
         );
  AND U9896 ( .A(n9812), .B(n9813), .Z(n9811) );
  OR U9897 ( .A(n9788), .B(n9804), .Z(n9813) );
  MUX U9898 ( .IN0(data_mem_out_wire[39]), .IN1(data_in[7]), .SEL(n9814), .F(
        n7705) );
  MUX U9899 ( .IN0(data_mem_out_wire[38]), .IN1(data_in[6]), .SEL(n9814), .F(
        n7704) );
  MUX U9900 ( .IN0(data_mem_out_wire[37]), .IN1(data_in[5]), .SEL(n9814), .F(
        n7703) );
  MUX U9901 ( .IN0(data_mem_out_wire[36]), .IN1(data_in[4]), .SEL(n9814), .F(
        n7702) );
  MUX U9902 ( .IN0(data_mem_out_wire[35]), .IN1(data_in[3]), .SEL(n9814), .F(
        n7701) );
  IV U9903 ( .A(n9815), .Z(n9814) );
  MUX U9904 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[34]), .SEL(n9815), .F(
        n7700) );
  MUX U9905 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[33]), .SEL(n9815), .F(
        n7699) );
  MUX U9906 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[32]), .SEL(n9815), .F(
        n7698) );
  AND U9907 ( .A(n9812), .B(n9816), .Z(n9815) );
  NANDN U9908 ( .A(n9804), .B(n9792), .Z(n9816) );
  AND U9909 ( .A(n9817), .B(n9801), .Z(n9812) );
  NANDN U9910 ( .A(n9804), .B(n9796), .Z(n9801) );
  NANDN U9911 ( .A(n9804), .B(n9818), .Z(n9817) );
  NAND U9912 ( .A(n9797), .B(n9819), .Z(n9804) );
  MUX U9913 ( .IN0(n9746), .IN1(data_mem_out_wire[95]), .SEL(n9820), .F(n7697)
         );
  MUX U9914 ( .IN0(n9748), .IN1(data_mem_out_wire[94]), .SEL(n9820), .F(n7696)
         );
  MUX U9915 ( .IN0(n9749), .IN1(data_mem_out_wire[93]), .SEL(n9820), .F(n7695)
         );
  MUX U9916 ( .IN0(n9750), .IN1(data_mem_out_wire[92]), .SEL(n9820), .F(n7694)
         );
  MUX U9917 ( .IN0(n9751), .IN1(data_mem_out_wire[91]), .SEL(n9820), .F(n7693)
         );
  MUX U9918 ( .IN0(n9752), .IN1(data_mem_out_wire[90]), .SEL(n9820), .F(n7692)
         );
  MUX U9919 ( .IN0(n9753), .IN1(data_mem_out_wire[89]), .SEL(n9820), .F(n7691)
         );
  MUX U9920 ( .IN0(n9754), .IN1(data_mem_out_wire[88]), .SEL(n9820), .F(n7690)
         );
  AND U9921 ( .A(n9821), .B(n9822), .Z(n9820) );
  AND U9922 ( .A(n9823), .B(n9824), .Z(n9821) );
  OR U9923 ( .A(n9760), .B(n9825), .Z(n9824) );
  MUX U9924 ( .IN0(data_mem_out_wire[87]), .IN1(n9761), .SEL(n9826), .F(n7689)
         );
  MUX U9925 ( .IN0(data_mem_out_wire[86]), .IN1(n9763), .SEL(n9826), .F(n7688)
         );
  MUX U9926 ( .IN0(data_mem_out_wire[85]), .IN1(n9764), .SEL(n9826), .F(n7687)
         );
  MUX U9927 ( .IN0(data_mem_out_wire[84]), .IN1(n9765), .SEL(n9826), .F(n7686)
         );
  MUX U9928 ( .IN0(data_mem_out_wire[83]), .IN1(n9766), .SEL(n9826), .F(n7685)
         );
  IV U9929 ( .A(n9827), .Z(n9826) );
  MUX U9930 ( .IN0(n9768), .IN1(data_mem_out_wire[82]), .SEL(n9827), .F(n7684)
         );
  MUX U9931 ( .IN0(n9769), .IN1(data_mem_out_wire[81]), .SEL(n9827), .F(n7683)
         );
  MUX U9932 ( .IN0(n9770), .IN1(data_mem_out_wire[80]), .SEL(n9827), .F(n7682)
         );
  AND U9933 ( .A(n9828), .B(n9829), .Z(n9827) );
  OR U9934 ( .A(n9773), .B(n9825), .Z(n9829) );
  AND U9935 ( .A(n9823), .B(n9822), .Z(n9828) );
  NANDN U9936 ( .A(n9825), .B(n9809), .Z(n9823) );
  MUX U9937 ( .IN0(data_mem_out_wire[79]), .IN1(n9776), .SEL(n9830), .F(n7681)
         );
  MUX U9938 ( .IN0(data_mem_out_wire[78]), .IN1(n9778), .SEL(n9830), .F(n7680)
         );
  MUX U9939 ( .IN0(data_mem_out_wire[77]), .IN1(n9779), .SEL(n9830), .F(n7679)
         );
  MUX U9940 ( .IN0(data_mem_out_wire[76]), .IN1(n9780), .SEL(n9830), .F(n7678)
         );
  MUX U9941 ( .IN0(data_mem_out_wire[75]), .IN1(n9781), .SEL(n9830), .F(n7677)
         );
  IV U9942 ( .A(n9831), .Z(n9830) );
  MUX U9943 ( .IN0(n9783), .IN1(data_mem_out_wire[74]), .SEL(n9831), .F(n7676)
         );
  MUX U9944 ( .IN0(n9784), .IN1(data_mem_out_wire[73]), .SEL(n9831), .F(n7675)
         );
  MUX U9945 ( .IN0(n9785), .IN1(data_mem_out_wire[72]), .SEL(n9831), .F(n7674)
         );
  AND U9946 ( .A(n9832), .B(n9833), .Z(n9831) );
  OR U9947 ( .A(n9788), .B(n9825), .Z(n9833) );
  MUX U9948 ( .IN0(data_mem_out_wire[71]), .IN1(data_in[7]), .SEL(n9834), .F(
        n7673) );
  MUX U9949 ( .IN0(data_mem_out_wire[70]), .IN1(data_in[6]), .SEL(n9834), .F(
        n7672) );
  MUX U9950 ( .IN0(data_mem_out_wire[69]), .IN1(data_in[5]), .SEL(n9834), .F(
        n7671) );
  MUX U9951 ( .IN0(data_mem_out_wire[68]), .IN1(data_in[4]), .SEL(n9834), .F(
        n7670) );
  MUX U9952 ( .IN0(data_mem_out_wire[67]), .IN1(data_in[3]), .SEL(n9834), .F(
        n7669) );
  IV U9953 ( .A(n9835), .Z(n9834) );
  MUX U9954 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[66]), .SEL(n9835), .F(
        n7668) );
  MUX U9955 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[65]), .SEL(n9835), .F(
        n7667) );
  MUX U9956 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[64]), .SEL(n9835), .F(
        n7666) );
  AND U9957 ( .A(n9832), .B(n9836), .Z(n9835) );
  NANDN U9958 ( .A(n9825), .B(n9792), .Z(n9836) );
  AND U9959 ( .A(n9837), .B(n9822), .Z(n9832) );
  NANDN U9960 ( .A(n9825), .B(n9796), .Z(n9822) );
  NANDN U9961 ( .A(n9825), .B(n9818), .Z(n9837) );
  NAND U9962 ( .A(n9797), .B(n9838), .Z(n9825) );
  MUX U9963 ( .IN0(n9746), .IN1(data_mem_out_wire[127]), .SEL(n9839), .F(n7665) );
  MUX U9964 ( .IN0(n9748), .IN1(data_mem_out_wire[126]), .SEL(n9839), .F(n7664) );
  MUX U9965 ( .IN0(n9749), .IN1(data_mem_out_wire[125]), .SEL(n9839), .F(n7663) );
  MUX U9966 ( .IN0(n9750), .IN1(data_mem_out_wire[124]), .SEL(n9839), .F(n7662) );
  MUX U9967 ( .IN0(n9751), .IN1(data_mem_out_wire[123]), .SEL(n9839), .F(n7661) );
  MUX U9968 ( .IN0(n9752), .IN1(data_mem_out_wire[122]), .SEL(n9839), .F(n7660) );
  MUX U9969 ( .IN0(n9753), .IN1(data_mem_out_wire[121]), .SEL(n9839), .F(n7659) );
  MUX U9970 ( .IN0(n9754), .IN1(data_mem_out_wire[120]), .SEL(n9839), .F(n7658) );
  AND U9971 ( .A(n9840), .B(n9841), .Z(n9839) );
  AND U9972 ( .A(n9842), .B(n9843), .Z(n9840) );
  OR U9973 ( .A(n9844), .B(n9845), .Z(n9843) );
  MUX U9974 ( .IN0(data_mem_out_wire[119]), .IN1(n9761), .SEL(n9846), .F(n7657) );
  MUX U9975 ( .IN0(data_mem_out_wire[118]), .IN1(n9763), .SEL(n9846), .F(n7656) );
  MUX U9976 ( .IN0(data_mem_out_wire[117]), .IN1(n9764), .SEL(n9846), .F(n7655) );
  MUX U9977 ( .IN0(data_mem_out_wire[116]), .IN1(n9765), .SEL(n9846), .F(n7654) );
  MUX U9978 ( .IN0(data_mem_out_wire[115]), .IN1(n9766), .SEL(n9846), .F(n7653) );
  IV U9979 ( .A(n9847), .Z(n9846) );
  MUX U9980 ( .IN0(n9768), .IN1(data_mem_out_wire[114]), .SEL(n9847), .F(n7652) );
  MUX U9981 ( .IN0(n9769), .IN1(data_mem_out_wire[113]), .SEL(n9847), .F(n7651) );
  MUX U9982 ( .IN0(n9770), .IN1(data_mem_out_wire[112]), .SEL(n9847), .F(n7650) );
  AND U9983 ( .A(n9848), .B(n9849), .Z(n9847) );
  OR U9984 ( .A(n9850), .B(n9845), .Z(n9849) );
  AND U9985 ( .A(n9842), .B(n9841), .Z(n9848) );
  NANDN U9986 ( .A(n9851), .B(n9809), .Z(n9842) );
  MUX U9987 ( .IN0(data_mem_out_wire[111]), .IN1(n9776), .SEL(n9852), .F(n7649) );
  MUX U9988 ( .IN0(data_mem_out_wire[110]), .IN1(n9778), .SEL(n9852), .F(n7648) );
  MUX U9989 ( .IN0(data_mem_out_wire[109]), .IN1(n9779), .SEL(n9852), .F(n7647) );
  MUX U9990 ( .IN0(data_mem_out_wire[108]), .IN1(n9780), .SEL(n9852), .F(n7646) );
  MUX U9991 ( .IN0(data_mem_out_wire[107]), .IN1(n9781), .SEL(n9852), .F(n7645) );
  IV U9992 ( .A(n9853), .Z(n9852) );
  MUX U9993 ( .IN0(n9783), .IN1(data_mem_out_wire[106]), .SEL(n9853), .F(n7644) );
  MUX U9994 ( .IN0(n9784), .IN1(data_mem_out_wire[105]), .SEL(n9853), .F(n7643) );
  MUX U9995 ( .IN0(n9785), .IN1(data_mem_out_wire[104]), .SEL(n9853), .F(n7642) );
  AND U9996 ( .A(n9854), .B(n9855), .Z(n9853) );
  NANDN U9997 ( .A(n9845), .B(n9856), .Z(n9855) );
  NANDN U9998 ( .A(n9851), .B(n9857), .Z(n9845) );
  MUX U9999 ( .IN0(data_mem_out_wire[103]), .IN1(data_in[7]), .SEL(n9858), .F(
        n7641) );
  MUX U10000 ( .IN0(data_mem_out_wire[102]), .IN1(data_in[6]), .SEL(n9858), 
        .F(n7640) );
  MUX U10001 ( .IN0(data_mem_out_wire[101]), .IN1(data_in[5]), .SEL(n9858), 
        .F(n7639) );
  MUX U10002 ( .IN0(data_mem_out_wire[100]), .IN1(data_in[4]), .SEL(n9858), 
        .F(n7638) );
  MUX U10003 ( .IN0(data_mem_out_wire[99]), .IN1(data_in[3]), .SEL(n9858), .F(
        n7637) );
  IV U10004 ( .A(n9859), .Z(n9858) );
  MUX U10005 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[98]), .SEL(n9859), .F(
        n7636) );
  MUX U10006 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[97]), .SEL(n9859), .F(
        n7635) );
  MUX U10007 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[96]), .SEL(n9859), .F(
        n7634) );
  AND U10008 ( .A(n9854), .B(n9860), .Z(n9859) );
  NANDN U10009 ( .A(n9851), .B(n9792), .Z(n9860) );
  AND U10010 ( .A(n9861), .B(n9841), .Z(n9854) );
  NANDN U10011 ( .A(n9851), .B(n9796), .Z(n9841) );
  NANDN U10012 ( .A(n9851), .B(n9818), .Z(n9861) );
  NAND U10013 ( .A(n9797), .B(n9862), .Z(n9851) );
  MUX U10014 ( .IN0(n9746), .IN1(data_mem_out_wire[159]), .SEL(n9863), .F(
        n7633) );
  MUX U10015 ( .IN0(n9748), .IN1(data_mem_out_wire[158]), .SEL(n9863), .F(
        n7632) );
  MUX U10016 ( .IN0(n9749), .IN1(data_mem_out_wire[157]), .SEL(n9863), .F(
        n7631) );
  MUX U10017 ( .IN0(n9750), .IN1(data_mem_out_wire[156]), .SEL(n9863), .F(
        n7630) );
  MUX U10018 ( .IN0(n9751), .IN1(data_mem_out_wire[155]), .SEL(n9863), .F(
        n7629) );
  MUX U10019 ( .IN0(n9752), .IN1(data_mem_out_wire[154]), .SEL(n9863), .F(
        n7628) );
  MUX U10020 ( .IN0(n9753), .IN1(data_mem_out_wire[153]), .SEL(n9863), .F(
        n7627) );
  MUX U10021 ( .IN0(n9754), .IN1(data_mem_out_wire[152]), .SEL(n9863), .F(
        n7626) );
  AND U10022 ( .A(n9864), .B(n9865), .Z(n9863) );
  AND U10023 ( .A(n9866), .B(n9867), .Z(n9864) );
  OR U10024 ( .A(n9760), .B(n9868), .Z(n9867) );
  MUX U10025 ( .IN0(data_mem_out_wire[151]), .IN1(n9761), .SEL(n9869), .F(
        n7625) );
  MUX U10026 ( .IN0(data_mem_out_wire[150]), .IN1(n9763), .SEL(n9869), .F(
        n7624) );
  MUX U10027 ( .IN0(data_mem_out_wire[149]), .IN1(n9764), .SEL(n9869), .F(
        n7623) );
  MUX U10028 ( .IN0(data_mem_out_wire[148]), .IN1(n9765), .SEL(n9869), .F(
        n7622) );
  MUX U10029 ( .IN0(data_mem_out_wire[147]), .IN1(n9766), .SEL(n9869), .F(
        n7621) );
  IV U10030 ( .A(n9870), .Z(n9869) );
  MUX U10031 ( .IN0(n9768), .IN1(data_mem_out_wire[146]), .SEL(n9870), .F(
        n7620) );
  MUX U10032 ( .IN0(n9769), .IN1(data_mem_out_wire[145]), .SEL(n9870), .F(
        n7619) );
  MUX U10033 ( .IN0(n9770), .IN1(data_mem_out_wire[144]), .SEL(n9870), .F(
        n7618) );
  AND U10034 ( .A(n9871), .B(n9872), .Z(n9870) );
  OR U10035 ( .A(n9773), .B(n9868), .Z(n9872) );
  AND U10036 ( .A(n9866), .B(n9865), .Z(n9871) );
  NANDN U10037 ( .A(n9868), .B(n9809), .Z(n9866) );
  MUX U10038 ( .IN0(data_mem_out_wire[143]), .IN1(n9776), .SEL(n9873), .F(
        n7617) );
  MUX U10039 ( .IN0(data_mem_out_wire[142]), .IN1(n9778), .SEL(n9873), .F(
        n7616) );
  MUX U10040 ( .IN0(data_mem_out_wire[141]), .IN1(n9779), .SEL(n9873), .F(
        n7615) );
  MUX U10041 ( .IN0(data_mem_out_wire[140]), .IN1(n9780), .SEL(n9873), .F(
        n7614) );
  MUX U10042 ( .IN0(data_mem_out_wire[139]), .IN1(n9781), .SEL(n9873), .F(
        n7613) );
  IV U10043 ( .A(n9874), .Z(n9873) );
  MUX U10044 ( .IN0(n9783), .IN1(data_mem_out_wire[138]), .SEL(n9874), .F(
        n7612) );
  MUX U10045 ( .IN0(n9784), .IN1(data_mem_out_wire[137]), .SEL(n9874), .F(
        n7611) );
  MUX U10046 ( .IN0(n9785), .IN1(data_mem_out_wire[136]), .SEL(n9874), .F(
        n7610) );
  AND U10047 ( .A(n9875), .B(n9876), .Z(n9874) );
  OR U10048 ( .A(n9788), .B(n9868), .Z(n9876) );
  MUX U10049 ( .IN0(data_mem_out_wire[135]), .IN1(data_in[7]), .SEL(n9877), 
        .F(n7609) );
  MUX U10050 ( .IN0(data_mem_out_wire[134]), .IN1(data_in[6]), .SEL(n9877), 
        .F(n7608) );
  MUX U10051 ( .IN0(data_mem_out_wire[133]), .IN1(data_in[5]), .SEL(n9877), 
        .F(n7607) );
  MUX U10052 ( .IN0(data_mem_out_wire[132]), .IN1(data_in[4]), .SEL(n9877), 
        .F(n7606) );
  MUX U10053 ( .IN0(data_mem_out_wire[131]), .IN1(data_in[3]), .SEL(n9877), 
        .F(n7605) );
  IV U10054 ( .A(n9878), .Z(n9877) );
  MUX U10055 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[130]), .SEL(n9878), 
        .F(n7604) );
  MUX U10056 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[129]), .SEL(n9878), 
        .F(n7603) );
  MUX U10057 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[128]), .SEL(n9878), 
        .F(n7602) );
  AND U10058 ( .A(n9875), .B(n9879), .Z(n9878) );
  NANDN U10059 ( .A(n9868), .B(n9792), .Z(n9879) );
  AND U10060 ( .A(n9880), .B(n9865), .Z(n9875) );
  NANDN U10061 ( .A(n9868), .B(n9796), .Z(n9865) );
  NANDN U10062 ( .A(n9868), .B(n9818), .Z(n9880) );
  NAND U10063 ( .A(n9797), .B(n9881), .Z(n9868) );
  MUX U10064 ( .IN0(n9746), .IN1(data_mem_out_wire[191]), .SEL(n9882), .F(
        n7601) );
  MUX U10065 ( .IN0(n9748), .IN1(data_mem_out_wire[190]), .SEL(n9882), .F(
        n7600) );
  MUX U10066 ( .IN0(n9749), .IN1(data_mem_out_wire[189]), .SEL(n9882), .F(
        n7599) );
  MUX U10067 ( .IN0(n9750), .IN1(data_mem_out_wire[188]), .SEL(n9882), .F(
        n7598) );
  MUX U10068 ( .IN0(n9751), .IN1(data_mem_out_wire[187]), .SEL(n9882), .F(
        n7597) );
  MUX U10069 ( .IN0(n9752), .IN1(data_mem_out_wire[186]), .SEL(n9882), .F(
        n7596) );
  MUX U10070 ( .IN0(n9753), .IN1(data_mem_out_wire[185]), .SEL(n9882), .F(
        n7595) );
  MUX U10071 ( .IN0(n9754), .IN1(data_mem_out_wire[184]), .SEL(n9882), .F(
        n7594) );
  AND U10072 ( .A(n9883), .B(n9884), .Z(n9882) );
  AND U10073 ( .A(n9885), .B(n9886), .Z(n9883) );
  OR U10074 ( .A(n9760), .B(n9887), .Z(n9886) );
  MUX U10075 ( .IN0(data_mem_out_wire[183]), .IN1(n9761), .SEL(n9888), .F(
        n7593) );
  MUX U10076 ( .IN0(data_mem_out_wire[182]), .IN1(n9763), .SEL(n9888), .F(
        n7592) );
  MUX U10077 ( .IN0(data_mem_out_wire[181]), .IN1(n9764), .SEL(n9888), .F(
        n7591) );
  MUX U10078 ( .IN0(data_mem_out_wire[180]), .IN1(n9765), .SEL(n9888), .F(
        n7590) );
  MUX U10079 ( .IN0(data_mem_out_wire[179]), .IN1(n9766), .SEL(n9888), .F(
        n7589) );
  IV U10080 ( .A(n9889), .Z(n9888) );
  MUX U10081 ( .IN0(n9768), .IN1(data_mem_out_wire[178]), .SEL(n9889), .F(
        n7588) );
  MUX U10082 ( .IN0(n9769), .IN1(data_mem_out_wire[177]), .SEL(n9889), .F(
        n7587) );
  MUX U10083 ( .IN0(n9770), .IN1(data_mem_out_wire[176]), .SEL(n9889), .F(
        n7586) );
  AND U10084 ( .A(n9890), .B(n9891), .Z(n9889) );
  OR U10085 ( .A(n9773), .B(n9887), .Z(n9891) );
  AND U10086 ( .A(n9885), .B(n9884), .Z(n9890) );
  NANDN U10087 ( .A(n9887), .B(n9809), .Z(n9885) );
  MUX U10088 ( .IN0(data_mem_out_wire[175]), .IN1(n9776), .SEL(n9892), .F(
        n7585) );
  MUX U10089 ( .IN0(data_mem_out_wire[174]), .IN1(n9778), .SEL(n9892), .F(
        n7584) );
  MUX U10090 ( .IN0(data_mem_out_wire[173]), .IN1(n9779), .SEL(n9892), .F(
        n7583) );
  MUX U10091 ( .IN0(data_mem_out_wire[172]), .IN1(n9780), .SEL(n9892), .F(
        n7582) );
  MUX U10092 ( .IN0(data_mem_out_wire[171]), .IN1(n9781), .SEL(n9892), .F(
        n7581) );
  IV U10093 ( .A(n9893), .Z(n9892) );
  MUX U10094 ( .IN0(n9783), .IN1(data_mem_out_wire[170]), .SEL(n9893), .F(
        n7580) );
  MUX U10095 ( .IN0(n9784), .IN1(data_mem_out_wire[169]), .SEL(n9893), .F(
        n7579) );
  MUX U10096 ( .IN0(n9785), .IN1(data_mem_out_wire[168]), .SEL(n9893), .F(
        n7578) );
  AND U10097 ( .A(n9894), .B(n9895), .Z(n9893) );
  OR U10098 ( .A(n9788), .B(n9887), .Z(n9895) );
  MUX U10099 ( .IN0(data_mem_out_wire[167]), .IN1(data_in[7]), .SEL(n9896), 
        .F(n7577) );
  MUX U10100 ( .IN0(data_mem_out_wire[166]), .IN1(data_in[6]), .SEL(n9896), 
        .F(n7576) );
  MUX U10101 ( .IN0(data_mem_out_wire[165]), .IN1(data_in[5]), .SEL(n9896), 
        .F(n7575) );
  MUX U10102 ( .IN0(data_mem_out_wire[164]), .IN1(data_in[4]), .SEL(n9896), 
        .F(n7574) );
  MUX U10103 ( .IN0(data_mem_out_wire[163]), .IN1(data_in[3]), .SEL(n9896), 
        .F(n7573) );
  IV U10104 ( .A(n9897), .Z(n9896) );
  MUX U10105 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[162]), .SEL(n9897), 
        .F(n7572) );
  MUX U10106 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[161]), .SEL(n9897), 
        .F(n7571) );
  MUX U10107 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[160]), .SEL(n9897), 
        .F(n7570) );
  AND U10108 ( .A(n9894), .B(n9898), .Z(n9897) );
  NANDN U10109 ( .A(n9887), .B(n9792), .Z(n9898) );
  AND U10110 ( .A(n9899), .B(n9884), .Z(n9894) );
  NANDN U10111 ( .A(n9887), .B(n9796), .Z(n9884) );
  NANDN U10112 ( .A(n9887), .B(n9818), .Z(n9899) );
  NAND U10113 ( .A(n9797), .B(n9900), .Z(n9887) );
  MUX U10114 ( .IN0(n9746), .IN1(data_mem_out_wire[223]), .SEL(n9901), .F(
        n7569) );
  MUX U10115 ( .IN0(n9748), .IN1(data_mem_out_wire[222]), .SEL(n9901), .F(
        n7568) );
  MUX U10116 ( .IN0(n9749), .IN1(data_mem_out_wire[221]), .SEL(n9901), .F(
        n7567) );
  MUX U10117 ( .IN0(n9750), .IN1(data_mem_out_wire[220]), .SEL(n9901), .F(
        n7566) );
  MUX U10118 ( .IN0(n9751), .IN1(data_mem_out_wire[219]), .SEL(n9901), .F(
        n7565) );
  MUX U10119 ( .IN0(n9752), .IN1(data_mem_out_wire[218]), .SEL(n9901), .F(
        n7564) );
  MUX U10120 ( .IN0(n9753), .IN1(data_mem_out_wire[217]), .SEL(n9901), .F(
        n7563) );
  MUX U10121 ( .IN0(n9754), .IN1(data_mem_out_wire[216]), .SEL(n9901), .F(
        n7562) );
  AND U10122 ( .A(n9902), .B(n9903), .Z(n9901) );
  AND U10123 ( .A(n9904), .B(n9905), .Z(n9902) );
  OR U10124 ( .A(n9760), .B(n9906), .Z(n9905) );
  MUX U10125 ( .IN0(data_mem_out_wire[215]), .IN1(n9761), .SEL(n9907), .F(
        n7561) );
  MUX U10126 ( .IN0(data_mem_out_wire[214]), .IN1(n9763), .SEL(n9907), .F(
        n7560) );
  MUX U10127 ( .IN0(data_mem_out_wire[213]), .IN1(n9764), .SEL(n9907), .F(
        n7559) );
  MUX U10128 ( .IN0(data_mem_out_wire[212]), .IN1(n9765), .SEL(n9907), .F(
        n7558) );
  MUX U10129 ( .IN0(data_mem_out_wire[211]), .IN1(n9766), .SEL(n9907), .F(
        n7557) );
  IV U10130 ( .A(n9908), .Z(n9907) );
  MUX U10131 ( .IN0(n9768), .IN1(data_mem_out_wire[210]), .SEL(n9908), .F(
        n7556) );
  MUX U10132 ( .IN0(n9769), .IN1(data_mem_out_wire[209]), .SEL(n9908), .F(
        n7555) );
  MUX U10133 ( .IN0(n9770), .IN1(data_mem_out_wire[208]), .SEL(n9908), .F(
        n7554) );
  AND U10134 ( .A(n9909), .B(n9910), .Z(n9908) );
  OR U10135 ( .A(n9773), .B(n9906), .Z(n9910) );
  AND U10136 ( .A(n9904), .B(n9903), .Z(n9909) );
  NANDN U10137 ( .A(n9906), .B(n9809), .Z(n9904) );
  MUX U10138 ( .IN0(data_mem_out_wire[207]), .IN1(n9776), .SEL(n9911), .F(
        n7553) );
  MUX U10139 ( .IN0(data_mem_out_wire[206]), .IN1(n9778), .SEL(n9911), .F(
        n7552) );
  MUX U10140 ( .IN0(data_mem_out_wire[205]), .IN1(n9779), .SEL(n9911), .F(
        n7551) );
  MUX U10141 ( .IN0(data_mem_out_wire[204]), .IN1(n9780), .SEL(n9911), .F(
        n7550) );
  MUX U10142 ( .IN0(data_mem_out_wire[203]), .IN1(n9781), .SEL(n9911), .F(
        n7549) );
  IV U10143 ( .A(n9912), .Z(n9911) );
  MUX U10144 ( .IN0(n9783), .IN1(data_mem_out_wire[202]), .SEL(n9912), .F(
        n7548) );
  MUX U10145 ( .IN0(n9784), .IN1(data_mem_out_wire[201]), .SEL(n9912), .F(
        n7547) );
  MUX U10146 ( .IN0(n9785), .IN1(data_mem_out_wire[200]), .SEL(n9912), .F(
        n7546) );
  AND U10147 ( .A(n9913), .B(n9914), .Z(n9912) );
  OR U10148 ( .A(n9788), .B(n9906), .Z(n9914) );
  MUX U10149 ( .IN0(data_mem_out_wire[199]), .IN1(data_in[7]), .SEL(n9915), 
        .F(n7545) );
  MUX U10150 ( .IN0(data_mem_out_wire[198]), .IN1(data_in[6]), .SEL(n9915), 
        .F(n7544) );
  MUX U10151 ( .IN0(data_mem_out_wire[197]), .IN1(data_in[5]), .SEL(n9915), 
        .F(n7543) );
  MUX U10152 ( .IN0(data_mem_out_wire[196]), .IN1(data_in[4]), .SEL(n9915), 
        .F(n7542) );
  MUX U10153 ( .IN0(data_mem_out_wire[195]), .IN1(data_in[3]), .SEL(n9915), 
        .F(n7541) );
  IV U10154 ( .A(n9916), .Z(n9915) );
  MUX U10155 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[194]), .SEL(n9916), 
        .F(n7540) );
  MUX U10156 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[193]), .SEL(n9916), 
        .F(n7539) );
  MUX U10157 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[192]), .SEL(n9916), 
        .F(n7538) );
  AND U10158 ( .A(n9913), .B(n9917), .Z(n9916) );
  NANDN U10159 ( .A(n9906), .B(n9792), .Z(n9917) );
  AND U10160 ( .A(n9918), .B(n9903), .Z(n9913) );
  NANDN U10161 ( .A(n9906), .B(n9796), .Z(n9903) );
  NANDN U10162 ( .A(n9906), .B(n9818), .Z(n9918) );
  NAND U10163 ( .A(n9797), .B(n9919), .Z(n9906) );
  MUX U10164 ( .IN0(n9746), .IN1(data_mem_out_wire[255]), .SEL(n9920), .F(
        n7537) );
  MUX U10165 ( .IN0(n9748), .IN1(data_mem_out_wire[254]), .SEL(n9920), .F(
        n7536) );
  MUX U10166 ( .IN0(n9749), .IN1(data_mem_out_wire[253]), .SEL(n9920), .F(
        n7535) );
  MUX U10167 ( .IN0(n9750), .IN1(data_mem_out_wire[252]), .SEL(n9920), .F(
        n7534) );
  MUX U10168 ( .IN0(n9751), .IN1(data_mem_out_wire[251]), .SEL(n9920), .F(
        n7533) );
  MUX U10169 ( .IN0(n9752), .IN1(data_mem_out_wire[250]), .SEL(n9920), .F(
        n7532) );
  MUX U10170 ( .IN0(n9753), .IN1(data_mem_out_wire[249]), .SEL(n9920), .F(
        n7531) );
  MUX U10171 ( .IN0(n9754), .IN1(data_mem_out_wire[248]), .SEL(n9920), .F(
        n7530) );
  AND U10172 ( .A(n9921), .B(n9922), .Z(n9920) );
  AND U10173 ( .A(n9923), .B(n9924), .Z(n9921) );
  OR U10174 ( .A(n9760), .B(n9925), .Z(n9924) );
  MUX U10175 ( .IN0(data_mem_out_wire[247]), .IN1(n9761), .SEL(n9926), .F(
        n7529) );
  MUX U10176 ( .IN0(data_mem_out_wire[246]), .IN1(n9763), .SEL(n9926), .F(
        n7528) );
  MUX U10177 ( .IN0(data_mem_out_wire[245]), .IN1(n9764), .SEL(n9926), .F(
        n7527) );
  MUX U10178 ( .IN0(data_mem_out_wire[244]), .IN1(n9765), .SEL(n9926), .F(
        n7526) );
  MUX U10179 ( .IN0(data_mem_out_wire[243]), .IN1(n9766), .SEL(n9926), .F(
        n7525) );
  IV U10180 ( .A(n9927), .Z(n9926) );
  MUX U10181 ( .IN0(n9768), .IN1(data_mem_out_wire[242]), .SEL(n9927), .F(
        n7524) );
  MUX U10182 ( .IN0(n9769), .IN1(data_mem_out_wire[241]), .SEL(n9927), .F(
        n7523) );
  MUX U10183 ( .IN0(n9770), .IN1(data_mem_out_wire[240]), .SEL(n9927), .F(
        n7522) );
  AND U10184 ( .A(n9928), .B(n9929), .Z(n9927) );
  OR U10185 ( .A(n9773), .B(n9925), .Z(n9929) );
  AND U10186 ( .A(n9923), .B(n9922), .Z(n9928) );
  NANDN U10187 ( .A(n9925), .B(n9809), .Z(n9923) );
  MUX U10188 ( .IN0(data_mem_out_wire[239]), .IN1(n9776), .SEL(n9930), .F(
        n7521) );
  MUX U10189 ( .IN0(data_mem_out_wire[238]), .IN1(n9778), .SEL(n9930), .F(
        n7520) );
  MUX U10190 ( .IN0(data_mem_out_wire[237]), .IN1(n9779), .SEL(n9930), .F(
        n7519) );
  MUX U10191 ( .IN0(data_mem_out_wire[236]), .IN1(n9780), .SEL(n9930), .F(
        n7518) );
  MUX U10192 ( .IN0(data_mem_out_wire[235]), .IN1(n9781), .SEL(n9930), .F(
        n7517) );
  IV U10193 ( .A(n9931), .Z(n9930) );
  MUX U10194 ( .IN0(n9783), .IN1(data_mem_out_wire[234]), .SEL(n9931), .F(
        n7516) );
  MUX U10195 ( .IN0(n9784), .IN1(data_mem_out_wire[233]), .SEL(n9931), .F(
        n7515) );
  MUX U10196 ( .IN0(n9785), .IN1(data_mem_out_wire[232]), .SEL(n9931), .F(
        n7514) );
  AND U10197 ( .A(n9932), .B(n9933), .Z(n9931) );
  OR U10198 ( .A(n9788), .B(n9925), .Z(n9933) );
  MUX U10199 ( .IN0(data_mem_out_wire[231]), .IN1(data_in[7]), .SEL(n9934), 
        .F(n7513) );
  MUX U10200 ( .IN0(data_mem_out_wire[230]), .IN1(data_in[6]), .SEL(n9934), 
        .F(n7512) );
  MUX U10201 ( .IN0(data_mem_out_wire[229]), .IN1(data_in[5]), .SEL(n9934), 
        .F(n7511) );
  MUX U10202 ( .IN0(data_mem_out_wire[228]), .IN1(data_in[4]), .SEL(n9934), 
        .F(n7510) );
  MUX U10203 ( .IN0(data_mem_out_wire[227]), .IN1(data_in[3]), .SEL(n9934), 
        .F(n7509) );
  IV U10204 ( .A(n9935), .Z(n9934) );
  MUX U10205 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[226]), .SEL(n9935), 
        .F(n7508) );
  MUX U10206 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[225]), .SEL(n9935), 
        .F(n7507) );
  MUX U10207 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[224]), .SEL(n9935), 
        .F(n7506) );
  AND U10208 ( .A(n9932), .B(n9936), .Z(n9935) );
  NANDN U10209 ( .A(n9925), .B(n9792), .Z(n9936) );
  AND U10210 ( .A(n9937), .B(n9922), .Z(n9932) );
  NANDN U10211 ( .A(n9925), .B(n9796), .Z(n9922) );
  NANDN U10212 ( .A(n9925), .B(n9818), .Z(n9937) );
  NAND U10213 ( .A(n9938), .B(n9797), .Z(n9925) );
  ANDN U10214 ( .B(n9939), .A(N42), .Z(n9797) );
  MUX U10215 ( .IN0(n9746), .IN1(data_mem_out_wire[287]), .SEL(n9940), .F(
        n7505) );
  MUX U10216 ( .IN0(n9748), .IN1(data_mem_out_wire[286]), .SEL(n9940), .F(
        n7504) );
  MUX U10217 ( .IN0(n9749), .IN1(data_mem_out_wire[285]), .SEL(n9940), .F(
        n7503) );
  MUX U10218 ( .IN0(n9750), .IN1(data_mem_out_wire[284]), .SEL(n9940), .F(
        n7502) );
  MUX U10219 ( .IN0(n9751), .IN1(data_mem_out_wire[283]), .SEL(n9940), .F(
        n7501) );
  MUX U10220 ( .IN0(n9752), .IN1(data_mem_out_wire[282]), .SEL(n9940), .F(
        n7500) );
  MUX U10221 ( .IN0(n9753), .IN1(data_mem_out_wire[281]), .SEL(n9940), .F(
        n7499) );
  MUX U10222 ( .IN0(n9754), .IN1(data_mem_out_wire[280]), .SEL(n9940), .F(
        n7498) );
  AND U10223 ( .A(n9941), .B(n9942), .Z(n9940) );
  AND U10224 ( .A(n9943), .B(n9944), .Z(n9941) );
  OR U10225 ( .A(n9760), .B(n9945), .Z(n9944) );
  MUX U10226 ( .IN0(data_mem_out_wire[279]), .IN1(n9761), .SEL(n9946), .F(
        n7497) );
  MUX U10227 ( .IN0(data_mem_out_wire[278]), .IN1(n9763), .SEL(n9946), .F(
        n7496) );
  MUX U10228 ( .IN0(data_mem_out_wire[277]), .IN1(n9764), .SEL(n9946), .F(
        n7495) );
  MUX U10229 ( .IN0(data_mem_out_wire[276]), .IN1(n9765), .SEL(n9946), .F(
        n7494) );
  MUX U10230 ( .IN0(data_mem_out_wire[275]), .IN1(n9766), .SEL(n9946), .F(
        n7493) );
  IV U10231 ( .A(n9947), .Z(n9946) );
  MUX U10232 ( .IN0(n9768), .IN1(data_mem_out_wire[274]), .SEL(n9947), .F(
        n7492) );
  MUX U10233 ( .IN0(n9769), .IN1(data_mem_out_wire[273]), .SEL(n9947), .F(
        n7491) );
  MUX U10234 ( .IN0(n9770), .IN1(data_mem_out_wire[272]), .SEL(n9947), .F(
        n7490) );
  AND U10235 ( .A(n9948), .B(n9949), .Z(n9947) );
  OR U10236 ( .A(n9773), .B(n9945), .Z(n9949) );
  AND U10237 ( .A(n9943), .B(n9942), .Z(n9948) );
  NANDN U10238 ( .A(n9945), .B(n9809), .Z(n9943) );
  MUX U10239 ( .IN0(data_mem_out_wire[271]), .IN1(n9776), .SEL(n9950), .F(
        n7489) );
  MUX U10240 ( .IN0(data_mem_out_wire[270]), .IN1(n9778), .SEL(n9950), .F(
        n7488) );
  MUX U10241 ( .IN0(data_mem_out_wire[269]), .IN1(n9779), .SEL(n9950), .F(
        n7487) );
  MUX U10242 ( .IN0(data_mem_out_wire[268]), .IN1(n9780), .SEL(n9950), .F(
        n7486) );
  MUX U10243 ( .IN0(data_mem_out_wire[267]), .IN1(n9781), .SEL(n9950), .F(
        n7485) );
  IV U10244 ( .A(n9951), .Z(n9950) );
  MUX U10245 ( .IN0(n9783), .IN1(data_mem_out_wire[266]), .SEL(n9951), .F(
        n7484) );
  MUX U10246 ( .IN0(n9784), .IN1(data_mem_out_wire[265]), .SEL(n9951), .F(
        n7483) );
  MUX U10247 ( .IN0(n9785), .IN1(data_mem_out_wire[264]), .SEL(n9951), .F(
        n7482) );
  AND U10248 ( .A(n9952), .B(n9953), .Z(n9951) );
  OR U10249 ( .A(n9788), .B(n9945), .Z(n9953) );
  MUX U10250 ( .IN0(data_mem_out_wire[263]), .IN1(data_in[7]), .SEL(n9954), 
        .F(n7481) );
  MUX U10251 ( .IN0(data_mem_out_wire[262]), .IN1(data_in[6]), .SEL(n9954), 
        .F(n7480) );
  MUX U10252 ( .IN0(data_mem_out_wire[261]), .IN1(data_in[5]), .SEL(n9954), 
        .F(n7479) );
  MUX U10253 ( .IN0(data_mem_out_wire[260]), .IN1(data_in[4]), .SEL(n9954), 
        .F(n7478) );
  MUX U10254 ( .IN0(data_mem_out_wire[259]), .IN1(data_in[3]), .SEL(n9954), 
        .F(n7477) );
  IV U10255 ( .A(n9955), .Z(n9954) );
  MUX U10256 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[258]), .SEL(n9955), 
        .F(n7476) );
  MUX U10257 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[257]), .SEL(n9955), 
        .F(n7475) );
  MUX U10258 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[256]), .SEL(n9955), 
        .F(n7474) );
  AND U10259 ( .A(n9952), .B(n9956), .Z(n9955) );
  NANDN U10260 ( .A(n9945), .B(n9792), .Z(n9956) );
  AND U10261 ( .A(n9957), .B(n9942), .Z(n9952) );
  NANDN U10262 ( .A(n9945), .B(n9796), .Z(n9942) );
  NANDN U10263 ( .A(n9945), .B(n9818), .Z(n9957) );
  NAND U10264 ( .A(n9798), .B(n9958), .Z(n9945) );
  MUX U10265 ( .IN0(n9746), .IN1(data_mem_out_wire[319]), .SEL(n9959), .F(
        n7473) );
  MUX U10266 ( .IN0(n9748), .IN1(data_mem_out_wire[318]), .SEL(n9959), .F(
        n7472) );
  MUX U10267 ( .IN0(n9749), .IN1(data_mem_out_wire[317]), .SEL(n9959), .F(
        n7471) );
  MUX U10268 ( .IN0(n9750), .IN1(data_mem_out_wire[316]), .SEL(n9959), .F(
        n7470) );
  MUX U10269 ( .IN0(n9751), .IN1(data_mem_out_wire[315]), .SEL(n9959), .F(
        n7469) );
  MUX U10270 ( .IN0(n9752), .IN1(data_mem_out_wire[314]), .SEL(n9959), .F(
        n7468) );
  MUX U10271 ( .IN0(n9753), .IN1(data_mem_out_wire[313]), .SEL(n9959), .F(
        n7467) );
  MUX U10272 ( .IN0(n9754), .IN1(data_mem_out_wire[312]), .SEL(n9959), .F(
        n7466) );
  AND U10273 ( .A(n9960), .B(n9961), .Z(n9959) );
  AND U10274 ( .A(n9962), .B(n9963), .Z(n9960) );
  OR U10275 ( .A(n9760), .B(n9964), .Z(n9963) );
  MUX U10276 ( .IN0(data_mem_out_wire[311]), .IN1(n9761), .SEL(n9965), .F(
        n7465) );
  MUX U10277 ( .IN0(data_mem_out_wire[310]), .IN1(n9763), .SEL(n9965), .F(
        n7464) );
  MUX U10278 ( .IN0(data_mem_out_wire[309]), .IN1(n9764), .SEL(n9965), .F(
        n7463) );
  MUX U10279 ( .IN0(data_mem_out_wire[308]), .IN1(n9765), .SEL(n9965), .F(
        n7462) );
  MUX U10280 ( .IN0(data_mem_out_wire[307]), .IN1(n9766), .SEL(n9965), .F(
        n7461) );
  IV U10281 ( .A(n9966), .Z(n9965) );
  MUX U10282 ( .IN0(n9768), .IN1(data_mem_out_wire[306]), .SEL(n9966), .F(
        n7460) );
  MUX U10283 ( .IN0(n9769), .IN1(data_mem_out_wire[305]), .SEL(n9966), .F(
        n7459) );
  MUX U10284 ( .IN0(n9770), .IN1(data_mem_out_wire[304]), .SEL(n9966), .F(
        n7458) );
  AND U10285 ( .A(n9967), .B(n9968), .Z(n9966) );
  OR U10286 ( .A(n9773), .B(n9964), .Z(n9968) );
  AND U10287 ( .A(n9962), .B(n9961), .Z(n9967) );
  NANDN U10288 ( .A(n9964), .B(n9809), .Z(n9962) );
  MUX U10289 ( .IN0(data_mem_out_wire[303]), .IN1(n9776), .SEL(n9969), .F(
        n7457) );
  MUX U10290 ( .IN0(data_mem_out_wire[302]), .IN1(n9778), .SEL(n9969), .F(
        n7456) );
  MUX U10291 ( .IN0(data_mem_out_wire[301]), .IN1(n9779), .SEL(n9969), .F(
        n7455) );
  MUX U10292 ( .IN0(data_mem_out_wire[300]), .IN1(n9780), .SEL(n9969), .F(
        n7454) );
  MUX U10293 ( .IN0(data_mem_out_wire[299]), .IN1(n9781), .SEL(n9969), .F(
        n7453) );
  IV U10294 ( .A(n9970), .Z(n9969) );
  MUX U10295 ( .IN0(n9783), .IN1(data_mem_out_wire[298]), .SEL(n9970), .F(
        n7452) );
  MUX U10296 ( .IN0(n9784), .IN1(data_mem_out_wire[297]), .SEL(n9970), .F(
        n7451) );
  MUX U10297 ( .IN0(n9785), .IN1(data_mem_out_wire[296]), .SEL(n9970), .F(
        n7450) );
  AND U10298 ( .A(n9971), .B(n9972), .Z(n9970) );
  OR U10299 ( .A(n9788), .B(n9964), .Z(n9972) );
  MUX U10300 ( .IN0(data_mem_out_wire[295]), .IN1(data_in[7]), .SEL(n9973), 
        .F(n7449) );
  MUX U10301 ( .IN0(data_mem_out_wire[294]), .IN1(data_in[6]), .SEL(n9973), 
        .F(n7448) );
  MUX U10302 ( .IN0(data_mem_out_wire[293]), .IN1(data_in[5]), .SEL(n9973), 
        .F(n7447) );
  MUX U10303 ( .IN0(data_mem_out_wire[292]), .IN1(data_in[4]), .SEL(n9973), 
        .F(n7446) );
  MUX U10304 ( .IN0(data_mem_out_wire[291]), .IN1(data_in[3]), .SEL(n9973), 
        .F(n7445) );
  IV U10305 ( .A(n9974), .Z(n9973) );
  MUX U10306 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[290]), .SEL(n9974), 
        .F(n7444) );
  MUX U10307 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[289]), .SEL(n9974), 
        .F(n7443) );
  MUX U10308 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[288]), .SEL(n9974), 
        .F(n7442) );
  AND U10309 ( .A(n9971), .B(n9975), .Z(n9974) );
  NANDN U10310 ( .A(n9964), .B(n9792), .Z(n9975) );
  AND U10311 ( .A(n9976), .B(n9961), .Z(n9971) );
  NANDN U10312 ( .A(n9964), .B(n9796), .Z(n9961) );
  NANDN U10313 ( .A(n9964), .B(n9818), .Z(n9976) );
  NAND U10314 ( .A(n9819), .B(n9958), .Z(n9964) );
  MUX U10315 ( .IN0(n9746), .IN1(data_mem_out_wire[351]), .SEL(n9977), .F(
        n7441) );
  MUX U10316 ( .IN0(n9748), .IN1(data_mem_out_wire[350]), .SEL(n9977), .F(
        n7440) );
  MUX U10317 ( .IN0(n9749), .IN1(data_mem_out_wire[349]), .SEL(n9977), .F(
        n7439) );
  MUX U10318 ( .IN0(n9750), .IN1(data_mem_out_wire[348]), .SEL(n9977), .F(
        n7438) );
  MUX U10319 ( .IN0(n9751), .IN1(data_mem_out_wire[347]), .SEL(n9977), .F(
        n7437) );
  MUX U10320 ( .IN0(n9752), .IN1(data_mem_out_wire[346]), .SEL(n9977), .F(
        n7436) );
  MUX U10321 ( .IN0(n9753), .IN1(data_mem_out_wire[345]), .SEL(n9977), .F(
        n7435) );
  MUX U10322 ( .IN0(n9754), .IN1(data_mem_out_wire[344]), .SEL(n9977), .F(
        n7434) );
  AND U10323 ( .A(n9978), .B(n9979), .Z(n9977) );
  AND U10324 ( .A(n9980), .B(n9981), .Z(n9978) );
  OR U10325 ( .A(n9760), .B(n9982), .Z(n9981) );
  MUX U10326 ( .IN0(data_mem_out_wire[343]), .IN1(n9761), .SEL(n9983), .F(
        n7433) );
  MUX U10327 ( .IN0(data_mem_out_wire[342]), .IN1(n9763), .SEL(n9983), .F(
        n7432) );
  MUX U10328 ( .IN0(data_mem_out_wire[341]), .IN1(n9764), .SEL(n9983), .F(
        n7431) );
  MUX U10329 ( .IN0(data_mem_out_wire[340]), .IN1(n9765), .SEL(n9983), .F(
        n7430) );
  MUX U10330 ( .IN0(data_mem_out_wire[339]), .IN1(n9766), .SEL(n9983), .F(
        n7429) );
  IV U10331 ( .A(n9984), .Z(n9983) );
  MUX U10332 ( .IN0(n9768), .IN1(data_mem_out_wire[338]), .SEL(n9984), .F(
        n7428) );
  MUX U10333 ( .IN0(n9769), .IN1(data_mem_out_wire[337]), .SEL(n9984), .F(
        n7427) );
  MUX U10334 ( .IN0(n9770), .IN1(data_mem_out_wire[336]), .SEL(n9984), .F(
        n7426) );
  AND U10335 ( .A(n9985), .B(n9986), .Z(n9984) );
  OR U10336 ( .A(n9773), .B(n9982), .Z(n9986) );
  AND U10337 ( .A(n9980), .B(n9979), .Z(n9985) );
  NANDN U10338 ( .A(n9982), .B(n9809), .Z(n9980) );
  MUX U10339 ( .IN0(data_mem_out_wire[335]), .IN1(n9776), .SEL(n9987), .F(
        n7425) );
  MUX U10340 ( .IN0(data_mem_out_wire[334]), .IN1(n9778), .SEL(n9987), .F(
        n7424) );
  MUX U10341 ( .IN0(data_mem_out_wire[333]), .IN1(n9779), .SEL(n9987), .F(
        n7423) );
  MUX U10342 ( .IN0(data_mem_out_wire[332]), .IN1(n9780), .SEL(n9987), .F(
        n7422) );
  MUX U10343 ( .IN0(data_mem_out_wire[331]), .IN1(n9781), .SEL(n9987), .F(
        n7421) );
  IV U10344 ( .A(n9988), .Z(n9987) );
  MUX U10345 ( .IN0(n9783), .IN1(data_mem_out_wire[330]), .SEL(n9988), .F(
        n7420) );
  MUX U10346 ( .IN0(n9784), .IN1(data_mem_out_wire[329]), .SEL(n9988), .F(
        n7419) );
  MUX U10347 ( .IN0(n9785), .IN1(data_mem_out_wire[328]), .SEL(n9988), .F(
        n7418) );
  AND U10348 ( .A(n9989), .B(n9990), .Z(n9988) );
  OR U10349 ( .A(n9788), .B(n9982), .Z(n9990) );
  MUX U10350 ( .IN0(data_mem_out_wire[327]), .IN1(data_in[7]), .SEL(n9991), 
        .F(n7417) );
  MUX U10351 ( .IN0(data_mem_out_wire[326]), .IN1(data_in[6]), .SEL(n9991), 
        .F(n7416) );
  MUX U10352 ( .IN0(data_mem_out_wire[325]), .IN1(data_in[5]), .SEL(n9991), 
        .F(n7415) );
  MUX U10353 ( .IN0(data_mem_out_wire[324]), .IN1(data_in[4]), .SEL(n9991), 
        .F(n7414) );
  MUX U10354 ( .IN0(data_mem_out_wire[323]), .IN1(data_in[3]), .SEL(n9991), 
        .F(n7413) );
  IV U10355 ( .A(n9992), .Z(n9991) );
  MUX U10356 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[322]), .SEL(n9992), 
        .F(n7412) );
  MUX U10357 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[321]), .SEL(n9992), 
        .F(n7411) );
  MUX U10358 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[320]), .SEL(n9992), 
        .F(n7410) );
  AND U10359 ( .A(n9989), .B(n9993), .Z(n9992) );
  NANDN U10360 ( .A(n9982), .B(n9792), .Z(n9993) );
  AND U10361 ( .A(n9994), .B(n9979), .Z(n9989) );
  NANDN U10362 ( .A(n9982), .B(n9796), .Z(n9979) );
  NANDN U10363 ( .A(n9982), .B(n9818), .Z(n9994) );
  NAND U10364 ( .A(n9838), .B(n9958), .Z(n9982) );
  MUX U10365 ( .IN0(n9746), .IN1(data_mem_out_wire[383]), .SEL(n9995), .F(
        n7409) );
  MUX U10366 ( .IN0(n9748), .IN1(data_mem_out_wire[382]), .SEL(n9995), .F(
        n7408) );
  MUX U10367 ( .IN0(n9749), .IN1(data_mem_out_wire[381]), .SEL(n9995), .F(
        n7407) );
  MUX U10368 ( .IN0(n9750), .IN1(data_mem_out_wire[380]), .SEL(n9995), .F(
        n7406) );
  MUX U10369 ( .IN0(n9751), .IN1(data_mem_out_wire[379]), .SEL(n9995), .F(
        n7405) );
  MUX U10370 ( .IN0(n9752), .IN1(data_mem_out_wire[378]), .SEL(n9995), .F(
        n7404) );
  MUX U10371 ( .IN0(n9753), .IN1(data_mem_out_wire[377]), .SEL(n9995), .F(
        n7403) );
  MUX U10372 ( .IN0(n9754), .IN1(data_mem_out_wire[376]), .SEL(n9995), .F(
        n7402) );
  AND U10373 ( .A(n9996), .B(n9997), .Z(n9995) );
  AND U10374 ( .A(n9998), .B(n9999), .Z(n9996) );
  OR U10375 ( .A(n9760), .B(n10000), .Z(n9999) );
  MUX U10376 ( .IN0(data_mem_out_wire[375]), .IN1(n9761), .SEL(n10001), .F(
        n7401) );
  MUX U10377 ( .IN0(data_mem_out_wire[374]), .IN1(n9763), .SEL(n10001), .F(
        n7400) );
  MUX U10378 ( .IN0(data_mem_out_wire[373]), .IN1(n9764), .SEL(n10001), .F(
        n7399) );
  MUX U10379 ( .IN0(data_mem_out_wire[372]), .IN1(n9765), .SEL(n10001), .F(
        n7398) );
  MUX U10380 ( .IN0(data_mem_out_wire[371]), .IN1(n9766), .SEL(n10001), .F(
        n7397) );
  IV U10381 ( .A(n10002), .Z(n10001) );
  MUX U10382 ( .IN0(n9768), .IN1(data_mem_out_wire[370]), .SEL(n10002), .F(
        n7396) );
  MUX U10383 ( .IN0(n9769), .IN1(data_mem_out_wire[369]), .SEL(n10002), .F(
        n7395) );
  MUX U10384 ( .IN0(n9770), .IN1(data_mem_out_wire[368]), .SEL(n10002), .F(
        n7394) );
  AND U10385 ( .A(n10003), .B(n10004), .Z(n10002) );
  OR U10386 ( .A(n9773), .B(n10000), .Z(n10004) );
  AND U10387 ( .A(n9998), .B(n9997), .Z(n10003) );
  NANDN U10388 ( .A(n10000), .B(n9809), .Z(n9998) );
  MUX U10389 ( .IN0(data_mem_out_wire[367]), .IN1(n9776), .SEL(n10005), .F(
        n7393) );
  MUX U10390 ( .IN0(data_mem_out_wire[366]), .IN1(n9778), .SEL(n10005), .F(
        n7392) );
  MUX U10391 ( .IN0(data_mem_out_wire[365]), .IN1(n9779), .SEL(n10005), .F(
        n7391) );
  MUX U10392 ( .IN0(data_mem_out_wire[364]), .IN1(n9780), .SEL(n10005), .F(
        n7390) );
  MUX U10393 ( .IN0(data_mem_out_wire[363]), .IN1(n9781), .SEL(n10005), .F(
        n7389) );
  IV U10394 ( .A(n10006), .Z(n10005) );
  MUX U10395 ( .IN0(n9783), .IN1(data_mem_out_wire[362]), .SEL(n10006), .F(
        n7388) );
  MUX U10396 ( .IN0(n9784), .IN1(data_mem_out_wire[361]), .SEL(n10006), .F(
        n7387) );
  MUX U10397 ( .IN0(n9785), .IN1(data_mem_out_wire[360]), .SEL(n10006), .F(
        n7386) );
  AND U10398 ( .A(n10007), .B(n10008), .Z(n10006) );
  OR U10399 ( .A(n9788), .B(n10000), .Z(n10008) );
  MUX U10400 ( .IN0(data_mem_out_wire[359]), .IN1(data_in[7]), .SEL(n10009), 
        .F(n7385) );
  MUX U10401 ( .IN0(data_mem_out_wire[358]), .IN1(data_in[6]), .SEL(n10009), 
        .F(n7384) );
  MUX U10402 ( .IN0(data_mem_out_wire[357]), .IN1(data_in[5]), .SEL(n10009), 
        .F(n7383) );
  MUX U10403 ( .IN0(data_mem_out_wire[356]), .IN1(data_in[4]), .SEL(n10009), 
        .F(n7382) );
  MUX U10404 ( .IN0(data_mem_out_wire[355]), .IN1(data_in[3]), .SEL(n10009), 
        .F(n7381) );
  IV U10405 ( .A(n10010), .Z(n10009) );
  MUX U10406 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[354]), .SEL(n10010), 
        .F(n7380) );
  MUX U10407 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[353]), .SEL(n10010), 
        .F(n7379) );
  MUX U10408 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[352]), .SEL(n10010), 
        .F(n7378) );
  AND U10409 ( .A(n10007), .B(n10011), .Z(n10010) );
  NANDN U10410 ( .A(n10000), .B(n9792), .Z(n10011) );
  AND U10411 ( .A(n10012), .B(n9997), .Z(n10007) );
  NANDN U10412 ( .A(n10000), .B(n9796), .Z(n9997) );
  NANDN U10413 ( .A(n10000), .B(n9818), .Z(n10012) );
  NAND U10414 ( .A(n9862), .B(n9958), .Z(n10000) );
  MUX U10415 ( .IN0(n9746), .IN1(data_mem_out_wire[415]), .SEL(n10013), .F(
        n7377) );
  MUX U10416 ( .IN0(n9748), .IN1(data_mem_out_wire[414]), .SEL(n10013), .F(
        n7376) );
  MUX U10417 ( .IN0(n9749), .IN1(data_mem_out_wire[413]), .SEL(n10013), .F(
        n7375) );
  MUX U10418 ( .IN0(n9750), .IN1(data_mem_out_wire[412]), .SEL(n10013), .F(
        n7374) );
  MUX U10419 ( .IN0(n9751), .IN1(data_mem_out_wire[411]), .SEL(n10013), .F(
        n7373) );
  MUX U10420 ( .IN0(n9752), .IN1(data_mem_out_wire[410]), .SEL(n10013), .F(
        n7372) );
  MUX U10421 ( .IN0(n9753), .IN1(data_mem_out_wire[409]), .SEL(n10013), .F(
        n7371) );
  MUX U10422 ( .IN0(n9754), .IN1(data_mem_out_wire[408]), .SEL(n10013), .F(
        n7370) );
  AND U10423 ( .A(n10014), .B(n10015), .Z(n10013) );
  AND U10424 ( .A(n10016), .B(n10017), .Z(n10014) );
  OR U10425 ( .A(n9760), .B(n10018), .Z(n10017) );
  MUX U10426 ( .IN0(data_mem_out_wire[407]), .IN1(n9761), .SEL(n10019), .F(
        n7369) );
  MUX U10427 ( .IN0(data_mem_out_wire[406]), .IN1(n9763), .SEL(n10019), .F(
        n7368) );
  MUX U10428 ( .IN0(data_mem_out_wire[405]), .IN1(n9764), .SEL(n10019), .F(
        n7367) );
  MUX U10429 ( .IN0(data_mem_out_wire[404]), .IN1(n9765), .SEL(n10019), .F(
        n7366) );
  MUX U10430 ( .IN0(data_mem_out_wire[403]), .IN1(n9766), .SEL(n10019), .F(
        n7365) );
  IV U10431 ( .A(n10020), .Z(n10019) );
  MUX U10432 ( .IN0(n9768), .IN1(data_mem_out_wire[402]), .SEL(n10020), .F(
        n7364) );
  MUX U10433 ( .IN0(n9769), .IN1(data_mem_out_wire[401]), .SEL(n10020), .F(
        n7363) );
  MUX U10434 ( .IN0(n9770), .IN1(data_mem_out_wire[400]), .SEL(n10020), .F(
        n7362) );
  AND U10435 ( .A(n10021), .B(n10022), .Z(n10020) );
  OR U10436 ( .A(n9773), .B(n10018), .Z(n10022) );
  AND U10437 ( .A(n10016), .B(n10015), .Z(n10021) );
  NANDN U10438 ( .A(n10018), .B(n9809), .Z(n10016) );
  MUX U10439 ( .IN0(data_mem_out_wire[399]), .IN1(n9776), .SEL(n10023), .F(
        n7361) );
  MUX U10440 ( .IN0(data_mem_out_wire[398]), .IN1(n9778), .SEL(n10023), .F(
        n7360) );
  MUX U10441 ( .IN0(data_mem_out_wire[397]), .IN1(n9779), .SEL(n10023), .F(
        n7359) );
  MUX U10442 ( .IN0(data_mem_out_wire[396]), .IN1(n9780), .SEL(n10023), .F(
        n7358) );
  MUX U10443 ( .IN0(data_mem_out_wire[395]), .IN1(n9781), .SEL(n10023), .F(
        n7357) );
  IV U10444 ( .A(n10024), .Z(n10023) );
  MUX U10445 ( .IN0(n9783), .IN1(data_mem_out_wire[394]), .SEL(n10024), .F(
        n7356) );
  MUX U10446 ( .IN0(n9784), .IN1(data_mem_out_wire[393]), .SEL(n10024), .F(
        n7355) );
  MUX U10447 ( .IN0(n9785), .IN1(data_mem_out_wire[392]), .SEL(n10024), .F(
        n7354) );
  AND U10448 ( .A(n10025), .B(n10026), .Z(n10024) );
  OR U10449 ( .A(n9788), .B(n10018), .Z(n10026) );
  MUX U10450 ( .IN0(data_mem_out_wire[391]), .IN1(data_in[7]), .SEL(n10027), 
        .F(n7353) );
  MUX U10451 ( .IN0(data_mem_out_wire[390]), .IN1(data_in[6]), .SEL(n10027), 
        .F(n7352) );
  MUX U10452 ( .IN0(data_mem_out_wire[389]), .IN1(data_in[5]), .SEL(n10027), 
        .F(n7351) );
  MUX U10453 ( .IN0(data_mem_out_wire[388]), .IN1(data_in[4]), .SEL(n10027), 
        .F(n7350) );
  MUX U10454 ( .IN0(data_mem_out_wire[387]), .IN1(data_in[3]), .SEL(n10027), 
        .F(n7349) );
  IV U10455 ( .A(n10028), .Z(n10027) );
  MUX U10456 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[386]), .SEL(n10028), 
        .F(n7348) );
  MUX U10457 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[385]), .SEL(n10028), 
        .F(n7347) );
  MUX U10458 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[384]), .SEL(n10028), 
        .F(n7346) );
  AND U10459 ( .A(n10025), .B(n10029), .Z(n10028) );
  NANDN U10460 ( .A(n10018), .B(n9792), .Z(n10029) );
  AND U10461 ( .A(n10030), .B(n10015), .Z(n10025) );
  NANDN U10462 ( .A(n10018), .B(n9796), .Z(n10015) );
  NANDN U10463 ( .A(n10018), .B(n9818), .Z(n10030) );
  NAND U10464 ( .A(n9881), .B(n9958), .Z(n10018) );
  MUX U10465 ( .IN0(n9746), .IN1(data_mem_out_wire[447]), .SEL(n10031), .F(
        n7345) );
  MUX U10466 ( .IN0(n9748), .IN1(data_mem_out_wire[446]), .SEL(n10031), .F(
        n7344) );
  MUX U10467 ( .IN0(n9749), .IN1(data_mem_out_wire[445]), .SEL(n10031), .F(
        n7343) );
  MUX U10468 ( .IN0(n9750), .IN1(data_mem_out_wire[444]), .SEL(n10031), .F(
        n7342) );
  MUX U10469 ( .IN0(n9751), .IN1(data_mem_out_wire[443]), .SEL(n10031), .F(
        n7341) );
  MUX U10470 ( .IN0(n9752), .IN1(data_mem_out_wire[442]), .SEL(n10031), .F(
        n7340) );
  MUX U10471 ( .IN0(n9753), .IN1(data_mem_out_wire[441]), .SEL(n10031), .F(
        n7339) );
  MUX U10472 ( .IN0(n9754), .IN1(data_mem_out_wire[440]), .SEL(n10031), .F(
        n7338) );
  AND U10473 ( .A(n10032), .B(n10033), .Z(n10031) );
  AND U10474 ( .A(n10034), .B(n10035), .Z(n10032) );
  OR U10475 ( .A(n9760), .B(n10036), .Z(n10035) );
  MUX U10476 ( .IN0(data_mem_out_wire[439]), .IN1(n9761), .SEL(n10037), .F(
        n7337) );
  MUX U10477 ( .IN0(data_mem_out_wire[438]), .IN1(n9763), .SEL(n10037), .F(
        n7336) );
  MUX U10478 ( .IN0(data_mem_out_wire[437]), .IN1(n9764), .SEL(n10037), .F(
        n7335) );
  MUX U10479 ( .IN0(data_mem_out_wire[436]), .IN1(n9765), .SEL(n10037), .F(
        n7334) );
  MUX U10480 ( .IN0(data_mem_out_wire[435]), .IN1(n9766), .SEL(n10037), .F(
        n7333) );
  IV U10481 ( .A(n10038), .Z(n10037) );
  MUX U10482 ( .IN0(n9768), .IN1(data_mem_out_wire[434]), .SEL(n10038), .F(
        n7332) );
  MUX U10483 ( .IN0(n9769), .IN1(data_mem_out_wire[433]), .SEL(n10038), .F(
        n7331) );
  MUX U10484 ( .IN0(n9770), .IN1(data_mem_out_wire[432]), .SEL(n10038), .F(
        n7330) );
  AND U10485 ( .A(n10039), .B(n10040), .Z(n10038) );
  OR U10486 ( .A(n9773), .B(n10036), .Z(n10040) );
  AND U10487 ( .A(n10034), .B(n10033), .Z(n10039) );
  NANDN U10488 ( .A(n10036), .B(n9809), .Z(n10034) );
  MUX U10489 ( .IN0(data_mem_out_wire[431]), .IN1(n9776), .SEL(n10041), .F(
        n7329) );
  MUX U10490 ( .IN0(data_mem_out_wire[430]), .IN1(n9778), .SEL(n10041), .F(
        n7328) );
  MUX U10491 ( .IN0(data_mem_out_wire[429]), .IN1(n9779), .SEL(n10041), .F(
        n7327) );
  MUX U10492 ( .IN0(data_mem_out_wire[428]), .IN1(n9780), .SEL(n10041), .F(
        n7326) );
  MUX U10493 ( .IN0(data_mem_out_wire[427]), .IN1(n9781), .SEL(n10041), .F(
        n7325) );
  IV U10494 ( .A(n10042), .Z(n10041) );
  MUX U10495 ( .IN0(n9783), .IN1(data_mem_out_wire[426]), .SEL(n10042), .F(
        n7324) );
  MUX U10496 ( .IN0(n9784), .IN1(data_mem_out_wire[425]), .SEL(n10042), .F(
        n7323) );
  MUX U10497 ( .IN0(n9785), .IN1(data_mem_out_wire[424]), .SEL(n10042), .F(
        n7322) );
  AND U10498 ( .A(n10043), .B(n10044), .Z(n10042) );
  OR U10499 ( .A(n9788), .B(n10036), .Z(n10044) );
  MUX U10500 ( .IN0(data_mem_out_wire[423]), .IN1(data_in[7]), .SEL(n10045), 
        .F(n7321) );
  MUX U10501 ( .IN0(data_mem_out_wire[422]), .IN1(data_in[6]), .SEL(n10045), 
        .F(n7320) );
  MUX U10502 ( .IN0(data_mem_out_wire[421]), .IN1(data_in[5]), .SEL(n10045), 
        .F(n7319) );
  MUX U10503 ( .IN0(data_mem_out_wire[420]), .IN1(data_in[4]), .SEL(n10045), 
        .F(n7318) );
  MUX U10504 ( .IN0(data_mem_out_wire[419]), .IN1(data_in[3]), .SEL(n10045), 
        .F(n7317) );
  IV U10505 ( .A(n10046), .Z(n10045) );
  MUX U10506 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[418]), .SEL(n10046), 
        .F(n7316) );
  MUX U10507 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[417]), .SEL(n10046), 
        .F(n7315) );
  MUX U10508 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[416]), .SEL(n10046), 
        .F(n7314) );
  AND U10509 ( .A(n10043), .B(n10047), .Z(n10046) );
  NANDN U10510 ( .A(n10036), .B(n9792), .Z(n10047) );
  AND U10511 ( .A(n10048), .B(n10033), .Z(n10043) );
  NANDN U10512 ( .A(n10036), .B(n9796), .Z(n10033) );
  NANDN U10513 ( .A(n10036), .B(n9818), .Z(n10048) );
  NAND U10514 ( .A(n9900), .B(n9958), .Z(n10036) );
  MUX U10515 ( .IN0(n9746), .IN1(data_mem_out_wire[479]), .SEL(n10049), .F(
        n7313) );
  MUX U10516 ( .IN0(n9748), .IN1(data_mem_out_wire[478]), .SEL(n10049), .F(
        n7312) );
  MUX U10517 ( .IN0(n9749), .IN1(data_mem_out_wire[477]), .SEL(n10049), .F(
        n7311) );
  MUX U10518 ( .IN0(n9750), .IN1(data_mem_out_wire[476]), .SEL(n10049), .F(
        n7310) );
  MUX U10519 ( .IN0(n9751), .IN1(data_mem_out_wire[475]), .SEL(n10049), .F(
        n7309) );
  MUX U10520 ( .IN0(n9752), .IN1(data_mem_out_wire[474]), .SEL(n10049), .F(
        n7308) );
  MUX U10521 ( .IN0(n9753), .IN1(data_mem_out_wire[473]), .SEL(n10049), .F(
        n7307) );
  MUX U10522 ( .IN0(n9754), .IN1(data_mem_out_wire[472]), .SEL(n10049), .F(
        n7306) );
  AND U10523 ( .A(n10050), .B(n10051), .Z(n10049) );
  AND U10524 ( .A(n10052), .B(n10053), .Z(n10050) );
  OR U10525 ( .A(n9760), .B(n10054), .Z(n10053) );
  MUX U10526 ( .IN0(data_mem_out_wire[471]), .IN1(n9761), .SEL(n10055), .F(
        n7305) );
  MUX U10527 ( .IN0(data_mem_out_wire[470]), .IN1(n9763), .SEL(n10055), .F(
        n7304) );
  MUX U10528 ( .IN0(data_mem_out_wire[469]), .IN1(n9764), .SEL(n10055), .F(
        n7303) );
  MUX U10529 ( .IN0(data_mem_out_wire[468]), .IN1(n9765), .SEL(n10055), .F(
        n7302) );
  MUX U10530 ( .IN0(data_mem_out_wire[467]), .IN1(n9766), .SEL(n10055), .F(
        n7301) );
  IV U10531 ( .A(n10056), .Z(n10055) );
  MUX U10532 ( .IN0(n9768), .IN1(data_mem_out_wire[466]), .SEL(n10056), .F(
        n7300) );
  MUX U10533 ( .IN0(n9769), .IN1(data_mem_out_wire[465]), .SEL(n10056), .F(
        n7299) );
  MUX U10534 ( .IN0(n9770), .IN1(data_mem_out_wire[464]), .SEL(n10056), .F(
        n7298) );
  AND U10535 ( .A(n10057), .B(n10058), .Z(n10056) );
  OR U10536 ( .A(n9773), .B(n10054), .Z(n10058) );
  AND U10537 ( .A(n10052), .B(n10051), .Z(n10057) );
  NANDN U10538 ( .A(n10054), .B(n9809), .Z(n10052) );
  MUX U10539 ( .IN0(data_mem_out_wire[463]), .IN1(n9776), .SEL(n10059), .F(
        n7297) );
  MUX U10540 ( .IN0(data_mem_out_wire[462]), .IN1(n9778), .SEL(n10059), .F(
        n7296) );
  MUX U10541 ( .IN0(data_mem_out_wire[461]), .IN1(n9779), .SEL(n10059), .F(
        n7295) );
  MUX U10542 ( .IN0(data_mem_out_wire[460]), .IN1(n9780), .SEL(n10059), .F(
        n7294) );
  MUX U10543 ( .IN0(data_mem_out_wire[459]), .IN1(n9781), .SEL(n10059), .F(
        n7293) );
  IV U10544 ( .A(n10060), .Z(n10059) );
  MUX U10545 ( .IN0(n9783), .IN1(data_mem_out_wire[458]), .SEL(n10060), .F(
        n7292) );
  MUX U10546 ( .IN0(n9784), .IN1(data_mem_out_wire[457]), .SEL(n10060), .F(
        n7291) );
  MUX U10547 ( .IN0(n9785), .IN1(data_mem_out_wire[456]), .SEL(n10060), .F(
        n7290) );
  AND U10548 ( .A(n10061), .B(n10062), .Z(n10060) );
  OR U10549 ( .A(n9788), .B(n10054), .Z(n10062) );
  MUX U10550 ( .IN0(data_mem_out_wire[455]), .IN1(data_in[7]), .SEL(n10063), 
        .F(n7289) );
  MUX U10551 ( .IN0(data_mem_out_wire[454]), .IN1(data_in[6]), .SEL(n10063), 
        .F(n7288) );
  MUX U10552 ( .IN0(data_mem_out_wire[453]), .IN1(data_in[5]), .SEL(n10063), 
        .F(n7287) );
  MUX U10553 ( .IN0(data_mem_out_wire[452]), .IN1(data_in[4]), .SEL(n10063), 
        .F(n7286) );
  MUX U10554 ( .IN0(data_mem_out_wire[451]), .IN1(data_in[3]), .SEL(n10063), 
        .F(n7285) );
  IV U10555 ( .A(n10064), .Z(n10063) );
  MUX U10556 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[450]), .SEL(n10064), 
        .F(n7284) );
  MUX U10557 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[449]), .SEL(n10064), 
        .F(n7283) );
  MUX U10558 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[448]), .SEL(n10064), 
        .F(n7282) );
  AND U10559 ( .A(n10061), .B(n10065), .Z(n10064) );
  NANDN U10560 ( .A(n10054), .B(n9792), .Z(n10065) );
  AND U10561 ( .A(n10066), .B(n10051), .Z(n10061) );
  NANDN U10562 ( .A(n10054), .B(n9796), .Z(n10051) );
  NANDN U10563 ( .A(n10054), .B(n9818), .Z(n10066) );
  NAND U10564 ( .A(n9919), .B(n9958), .Z(n10054) );
  MUX U10565 ( .IN0(n9746), .IN1(data_mem_out_wire[511]), .SEL(n10067), .F(
        n7281) );
  MUX U10566 ( .IN0(n9748), .IN1(data_mem_out_wire[510]), .SEL(n10067), .F(
        n7280) );
  MUX U10567 ( .IN0(n9749), .IN1(data_mem_out_wire[509]), .SEL(n10067), .F(
        n7279) );
  MUX U10568 ( .IN0(n9750), .IN1(data_mem_out_wire[508]), .SEL(n10067), .F(
        n7278) );
  MUX U10569 ( .IN0(n9751), .IN1(data_mem_out_wire[507]), .SEL(n10067), .F(
        n7277) );
  MUX U10570 ( .IN0(n9752), .IN1(data_mem_out_wire[506]), .SEL(n10067), .F(
        n7276) );
  MUX U10571 ( .IN0(n9753), .IN1(data_mem_out_wire[505]), .SEL(n10067), .F(
        n7275) );
  MUX U10572 ( .IN0(n9754), .IN1(data_mem_out_wire[504]), .SEL(n10067), .F(
        n7274) );
  AND U10573 ( .A(n10068), .B(n10069), .Z(n10067) );
  AND U10574 ( .A(n10070), .B(n10071), .Z(n10068) );
  OR U10575 ( .A(n9760), .B(n10072), .Z(n10071) );
  MUX U10576 ( .IN0(data_mem_out_wire[503]), .IN1(n9761), .SEL(n10073), .F(
        n7273) );
  MUX U10577 ( .IN0(data_mem_out_wire[502]), .IN1(n9763), .SEL(n10073), .F(
        n7272) );
  MUX U10578 ( .IN0(data_mem_out_wire[501]), .IN1(n9764), .SEL(n10073), .F(
        n7271) );
  MUX U10579 ( .IN0(data_mem_out_wire[500]), .IN1(n9765), .SEL(n10073), .F(
        n7270) );
  MUX U10580 ( .IN0(data_mem_out_wire[499]), .IN1(n9766), .SEL(n10073), .F(
        n7269) );
  IV U10581 ( .A(n10074), .Z(n10073) );
  MUX U10582 ( .IN0(n9768), .IN1(data_mem_out_wire[498]), .SEL(n10074), .F(
        n7268) );
  MUX U10583 ( .IN0(n9769), .IN1(data_mem_out_wire[497]), .SEL(n10074), .F(
        n7267) );
  MUX U10584 ( .IN0(n9770), .IN1(data_mem_out_wire[496]), .SEL(n10074), .F(
        n7266) );
  AND U10585 ( .A(n10075), .B(n10076), .Z(n10074) );
  OR U10586 ( .A(n9773), .B(n10072), .Z(n10076) );
  AND U10587 ( .A(n10070), .B(n10069), .Z(n10075) );
  NANDN U10588 ( .A(n10072), .B(n9809), .Z(n10070) );
  MUX U10589 ( .IN0(data_mem_out_wire[495]), .IN1(n9776), .SEL(n10077), .F(
        n7265) );
  MUX U10590 ( .IN0(data_mem_out_wire[494]), .IN1(n9778), .SEL(n10077), .F(
        n7264) );
  MUX U10591 ( .IN0(data_mem_out_wire[493]), .IN1(n9779), .SEL(n10077), .F(
        n7263) );
  MUX U10592 ( .IN0(data_mem_out_wire[492]), .IN1(n9780), .SEL(n10077), .F(
        n7262) );
  MUX U10593 ( .IN0(data_mem_out_wire[491]), .IN1(n9781), .SEL(n10077), .F(
        n7261) );
  IV U10594 ( .A(n10078), .Z(n10077) );
  MUX U10595 ( .IN0(n9783), .IN1(data_mem_out_wire[490]), .SEL(n10078), .F(
        n7260) );
  MUX U10596 ( .IN0(n9784), .IN1(data_mem_out_wire[489]), .SEL(n10078), .F(
        n7259) );
  MUX U10597 ( .IN0(n9785), .IN1(data_mem_out_wire[488]), .SEL(n10078), .F(
        n7258) );
  AND U10598 ( .A(n10079), .B(n10080), .Z(n10078) );
  OR U10599 ( .A(n9788), .B(n10072), .Z(n10080) );
  MUX U10600 ( .IN0(data_mem_out_wire[487]), .IN1(data_in[7]), .SEL(n10081), 
        .F(n7257) );
  MUX U10601 ( .IN0(data_mem_out_wire[486]), .IN1(data_in[6]), .SEL(n10081), 
        .F(n7256) );
  MUX U10602 ( .IN0(data_mem_out_wire[485]), .IN1(data_in[5]), .SEL(n10081), 
        .F(n7255) );
  MUX U10603 ( .IN0(data_mem_out_wire[484]), .IN1(data_in[4]), .SEL(n10081), 
        .F(n7254) );
  MUX U10604 ( .IN0(data_mem_out_wire[483]), .IN1(data_in[3]), .SEL(n10081), 
        .F(n7253) );
  IV U10605 ( .A(n10082), .Z(n10081) );
  MUX U10606 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[482]), .SEL(n10082), 
        .F(n7252) );
  MUX U10607 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[481]), .SEL(n10082), 
        .F(n7251) );
  MUX U10608 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[480]), .SEL(n10082), 
        .F(n7250) );
  AND U10609 ( .A(n10079), .B(n10083), .Z(n10082) );
  NANDN U10610 ( .A(n10072), .B(n9792), .Z(n10083) );
  AND U10611 ( .A(n10084), .B(n10069), .Z(n10079) );
  NANDN U10612 ( .A(n10072), .B(n9796), .Z(n10069) );
  NANDN U10613 ( .A(n10072), .B(n9818), .Z(n10084) );
  NAND U10614 ( .A(n9958), .B(n9938), .Z(n10072) );
  ANDN U10615 ( .B(n10085), .A(N42), .Z(n9958) );
  MUX U10616 ( .IN0(n9746), .IN1(data_mem_out_wire[543]), .SEL(n10086), .F(
        n7249) );
  MUX U10617 ( .IN0(n9748), .IN1(data_mem_out_wire[542]), .SEL(n10086), .F(
        n7248) );
  MUX U10618 ( .IN0(n9749), .IN1(data_mem_out_wire[541]), .SEL(n10086), .F(
        n7247) );
  MUX U10619 ( .IN0(n9750), .IN1(data_mem_out_wire[540]), .SEL(n10086), .F(
        n7246) );
  MUX U10620 ( .IN0(n9751), .IN1(data_mem_out_wire[539]), .SEL(n10086), .F(
        n7245) );
  MUX U10621 ( .IN0(n9752), .IN1(data_mem_out_wire[538]), .SEL(n10086), .F(
        n7244) );
  MUX U10622 ( .IN0(n9753), .IN1(data_mem_out_wire[537]), .SEL(n10086), .F(
        n7243) );
  MUX U10623 ( .IN0(n9754), .IN1(data_mem_out_wire[536]), .SEL(n10086), .F(
        n7242) );
  AND U10624 ( .A(n10087), .B(n10088), .Z(n10086) );
  AND U10625 ( .A(n10089), .B(n10090), .Z(n10087) );
  OR U10626 ( .A(n9760), .B(n10091), .Z(n10090) );
  MUX U10627 ( .IN0(data_mem_out_wire[535]), .IN1(n9761), .SEL(n10092), .F(
        n7241) );
  MUX U10628 ( .IN0(data_mem_out_wire[534]), .IN1(n9763), .SEL(n10092), .F(
        n7240) );
  MUX U10629 ( .IN0(data_mem_out_wire[533]), .IN1(n9764), .SEL(n10092), .F(
        n7239) );
  MUX U10630 ( .IN0(data_mem_out_wire[532]), .IN1(n9765), .SEL(n10092), .F(
        n7238) );
  MUX U10631 ( .IN0(data_mem_out_wire[531]), .IN1(n9766), .SEL(n10092), .F(
        n7237) );
  IV U10632 ( .A(n10093), .Z(n10092) );
  MUX U10633 ( .IN0(n9768), .IN1(data_mem_out_wire[530]), .SEL(n10093), .F(
        n7236) );
  MUX U10634 ( .IN0(n9769), .IN1(data_mem_out_wire[529]), .SEL(n10093), .F(
        n7235) );
  MUX U10635 ( .IN0(n9770), .IN1(data_mem_out_wire[528]), .SEL(n10093), .F(
        n7234) );
  AND U10636 ( .A(n10094), .B(n10095), .Z(n10093) );
  OR U10637 ( .A(n9773), .B(n10091), .Z(n10095) );
  AND U10638 ( .A(n10089), .B(n10088), .Z(n10094) );
  NANDN U10639 ( .A(n10091), .B(n9809), .Z(n10089) );
  MUX U10640 ( .IN0(data_mem_out_wire[527]), .IN1(n9776), .SEL(n10096), .F(
        n7233) );
  MUX U10641 ( .IN0(data_mem_out_wire[526]), .IN1(n9778), .SEL(n10096), .F(
        n7232) );
  MUX U10642 ( .IN0(data_mem_out_wire[525]), .IN1(n9779), .SEL(n10096), .F(
        n7231) );
  MUX U10643 ( .IN0(data_mem_out_wire[524]), .IN1(n9780), .SEL(n10096), .F(
        n7230) );
  MUX U10644 ( .IN0(data_mem_out_wire[523]), .IN1(n9781), .SEL(n10096), .F(
        n7229) );
  IV U10645 ( .A(n10097), .Z(n10096) );
  MUX U10646 ( .IN0(n9783), .IN1(data_mem_out_wire[522]), .SEL(n10097), .F(
        n7228) );
  MUX U10647 ( .IN0(n9784), .IN1(data_mem_out_wire[521]), .SEL(n10097), .F(
        n7227) );
  MUX U10648 ( .IN0(n9785), .IN1(data_mem_out_wire[520]), .SEL(n10097), .F(
        n7226) );
  AND U10649 ( .A(n10098), .B(n10099), .Z(n10097) );
  OR U10650 ( .A(n9788), .B(n10091), .Z(n10099) );
  MUX U10651 ( .IN0(data_mem_out_wire[519]), .IN1(data_in[7]), .SEL(n10100), 
        .F(n7225) );
  MUX U10652 ( .IN0(data_mem_out_wire[518]), .IN1(data_in[6]), .SEL(n10100), 
        .F(n7224) );
  MUX U10653 ( .IN0(data_mem_out_wire[517]), .IN1(data_in[5]), .SEL(n10100), 
        .F(n7223) );
  MUX U10654 ( .IN0(data_mem_out_wire[516]), .IN1(data_in[4]), .SEL(n10100), 
        .F(n7222) );
  MUX U10655 ( .IN0(data_mem_out_wire[515]), .IN1(data_in[3]), .SEL(n10100), 
        .F(n7221) );
  IV U10656 ( .A(n10101), .Z(n10100) );
  MUX U10657 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[514]), .SEL(n10101), 
        .F(n7220) );
  MUX U10658 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[513]), .SEL(n10101), 
        .F(n7219) );
  MUX U10659 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[512]), .SEL(n10101), 
        .F(n7218) );
  AND U10660 ( .A(n10098), .B(n10102), .Z(n10101) );
  NANDN U10661 ( .A(n10091), .B(n9792), .Z(n10102) );
  AND U10662 ( .A(n10103), .B(n10088), .Z(n10098) );
  NANDN U10663 ( .A(n10091), .B(n9796), .Z(n10088) );
  NANDN U10664 ( .A(n10091), .B(n9818), .Z(n10103) );
  NAND U10665 ( .A(n9798), .B(n10104), .Z(n10091) );
  MUX U10666 ( .IN0(n9746), .IN1(data_mem_out_wire[575]), .SEL(n10105), .F(
        n7217) );
  MUX U10667 ( .IN0(n9748), .IN1(data_mem_out_wire[574]), .SEL(n10105), .F(
        n7216) );
  MUX U10668 ( .IN0(n9749), .IN1(data_mem_out_wire[573]), .SEL(n10105), .F(
        n7215) );
  MUX U10669 ( .IN0(n9750), .IN1(data_mem_out_wire[572]), .SEL(n10105), .F(
        n7214) );
  MUX U10670 ( .IN0(n9751), .IN1(data_mem_out_wire[571]), .SEL(n10105), .F(
        n7213) );
  MUX U10671 ( .IN0(n9752), .IN1(data_mem_out_wire[570]), .SEL(n10105), .F(
        n7212) );
  MUX U10672 ( .IN0(n9753), .IN1(data_mem_out_wire[569]), .SEL(n10105), .F(
        n7211) );
  MUX U10673 ( .IN0(n9754), .IN1(data_mem_out_wire[568]), .SEL(n10105), .F(
        n7210) );
  AND U10674 ( .A(n10106), .B(n10107), .Z(n10105) );
  AND U10675 ( .A(n10108), .B(n10109), .Z(n10106) );
  OR U10676 ( .A(n9760), .B(n10110), .Z(n10109) );
  MUX U10677 ( .IN0(data_mem_out_wire[567]), .IN1(n9761), .SEL(n10111), .F(
        n7209) );
  MUX U10678 ( .IN0(data_mem_out_wire[566]), .IN1(n9763), .SEL(n10111), .F(
        n7208) );
  MUX U10679 ( .IN0(data_mem_out_wire[565]), .IN1(n9764), .SEL(n10111), .F(
        n7207) );
  MUX U10680 ( .IN0(data_mem_out_wire[564]), .IN1(n9765), .SEL(n10111), .F(
        n7206) );
  MUX U10681 ( .IN0(data_mem_out_wire[563]), .IN1(n9766), .SEL(n10111), .F(
        n7205) );
  IV U10682 ( .A(n10112), .Z(n10111) );
  MUX U10683 ( .IN0(n9768), .IN1(data_mem_out_wire[562]), .SEL(n10112), .F(
        n7204) );
  MUX U10684 ( .IN0(n9769), .IN1(data_mem_out_wire[561]), .SEL(n10112), .F(
        n7203) );
  MUX U10685 ( .IN0(n9770), .IN1(data_mem_out_wire[560]), .SEL(n10112), .F(
        n7202) );
  AND U10686 ( .A(n10113), .B(n10114), .Z(n10112) );
  OR U10687 ( .A(n9773), .B(n10110), .Z(n10114) );
  AND U10688 ( .A(n10108), .B(n10107), .Z(n10113) );
  NANDN U10689 ( .A(n10110), .B(n9809), .Z(n10108) );
  MUX U10690 ( .IN0(data_mem_out_wire[559]), .IN1(n9776), .SEL(n10115), .F(
        n7201) );
  MUX U10691 ( .IN0(data_mem_out_wire[558]), .IN1(n9778), .SEL(n10115), .F(
        n7200) );
  MUX U10692 ( .IN0(data_mem_out_wire[557]), .IN1(n9779), .SEL(n10115), .F(
        n7199) );
  MUX U10693 ( .IN0(data_mem_out_wire[556]), .IN1(n9780), .SEL(n10115), .F(
        n7198) );
  MUX U10694 ( .IN0(data_mem_out_wire[555]), .IN1(n9781), .SEL(n10115), .F(
        n7197) );
  IV U10695 ( .A(n10116), .Z(n10115) );
  MUX U10696 ( .IN0(n9783), .IN1(data_mem_out_wire[554]), .SEL(n10116), .F(
        n7196) );
  MUX U10697 ( .IN0(n9784), .IN1(data_mem_out_wire[553]), .SEL(n10116), .F(
        n7195) );
  MUX U10698 ( .IN0(n9785), .IN1(data_mem_out_wire[552]), .SEL(n10116), .F(
        n7194) );
  AND U10699 ( .A(n10117), .B(n10118), .Z(n10116) );
  OR U10700 ( .A(n9788), .B(n10110), .Z(n10118) );
  MUX U10701 ( .IN0(data_mem_out_wire[551]), .IN1(data_in[7]), .SEL(n10119), 
        .F(n7193) );
  MUX U10702 ( .IN0(data_mem_out_wire[550]), .IN1(data_in[6]), .SEL(n10119), 
        .F(n7192) );
  MUX U10703 ( .IN0(data_mem_out_wire[549]), .IN1(data_in[5]), .SEL(n10119), 
        .F(n7191) );
  MUX U10704 ( .IN0(data_mem_out_wire[548]), .IN1(data_in[4]), .SEL(n10119), 
        .F(n7190) );
  MUX U10705 ( .IN0(data_mem_out_wire[547]), .IN1(data_in[3]), .SEL(n10119), 
        .F(n7189) );
  IV U10706 ( .A(n10120), .Z(n10119) );
  MUX U10707 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[546]), .SEL(n10120), 
        .F(n7188) );
  MUX U10708 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[545]), .SEL(n10120), 
        .F(n7187) );
  MUX U10709 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[544]), .SEL(n10120), 
        .F(n7186) );
  AND U10710 ( .A(n10117), .B(n10121), .Z(n10120) );
  NANDN U10711 ( .A(n10110), .B(n9792), .Z(n10121) );
  AND U10712 ( .A(n10122), .B(n10107), .Z(n10117) );
  NANDN U10713 ( .A(n10110), .B(n9796), .Z(n10107) );
  NANDN U10714 ( .A(n10110), .B(n9818), .Z(n10122) );
  NAND U10715 ( .A(n9819), .B(n10104), .Z(n10110) );
  MUX U10716 ( .IN0(n9746), .IN1(data_mem_out_wire[607]), .SEL(n10123), .F(
        n7185) );
  MUX U10717 ( .IN0(n9748), .IN1(data_mem_out_wire[606]), .SEL(n10123), .F(
        n7184) );
  MUX U10718 ( .IN0(n9749), .IN1(data_mem_out_wire[605]), .SEL(n10123), .F(
        n7183) );
  MUX U10719 ( .IN0(n9750), .IN1(data_mem_out_wire[604]), .SEL(n10123), .F(
        n7182) );
  MUX U10720 ( .IN0(n9751), .IN1(data_mem_out_wire[603]), .SEL(n10123), .F(
        n7181) );
  MUX U10721 ( .IN0(n9752), .IN1(data_mem_out_wire[602]), .SEL(n10123), .F(
        n7180) );
  MUX U10722 ( .IN0(n9753), .IN1(data_mem_out_wire[601]), .SEL(n10123), .F(
        n7179) );
  MUX U10723 ( .IN0(n9754), .IN1(data_mem_out_wire[600]), .SEL(n10123), .F(
        n7178) );
  AND U10724 ( .A(n10124), .B(n10125), .Z(n10123) );
  AND U10725 ( .A(n10126), .B(n10127), .Z(n10124) );
  OR U10726 ( .A(n9760), .B(n10128), .Z(n10127) );
  MUX U10727 ( .IN0(data_mem_out_wire[599]), .IN1(n9761), .SEL(n10129), .F(
        n7177) );
  MUX U10728 ( .IN0(data_mem_out_wire[598]), .IN1(n9763), .SEL(n10129), .F(
        n7176) );
  MUX U10729 ( .IN0(data_mem_out_wire[597]), .IN1(n9764), .SEL(n10129), .F(
        n7175) );
  MUX U10730 ( .IN0(data_mem_out_wire[596]), .IN1(n9765), .SEL(n10129), .F(
        n7174) );
  MUX U10731 ( .IN0(data_mem_out_wire[595]), .IN1(n9766), .SEL(n10129), .F(
        n7173) );
  IV U10732 ( .A(n10130), .Z(n10129) );
  MUX U10733 ( .IN0(n9768), .IN1(data_mem_out_wire[594]), .SEL(n10130), .F(
        n7172) );
  MUX U10734 ( .IN0(n9769), .IN1(data_mem_out_wire[593]), .SEL(n10130), .F(
        n7171) );
  MUX U10735 ( .IN0(n9770), .IN1(data_mem_out_wire[592]), .SEL(n10130), .F(
        n7170) );
  AND U10736 ( .A(n10131), .B(n10132), .Z(n10130) );
  OR U10737 ( .A(n9773), .B(n10128), .Z(n10132) );
  AND U10738 ( .A(n10126), .B(n10125), .Z(n10131) );
  NANDN U10739 ( .A(n10128), .B(n9809), .Z(n10126) );
  MUX U10740 ( .IN0(data_mem_out_wire[591]), .IN1(n9776), .SEL(n10133), .F(
        n7169) );
  MUX U10741 ( .IN0(data_mem_out_wire[590]), .IN1(n9778), .SEL(n10133), .F(
        n7168) );
  MUX U10742 ( .IN0(data_mem_out_wire[589]), .IN1(n9779), .SEL(n10133), .F(
        n7167) );
  MUX U10743 ( .IN0(data_mem_out_wire[588]), .IN1(n9780), .SEL(n10133), .F(
        n7166) );
  MUX U10744 ( .IN0(data_mem_out_wire[587]), .IN1(n9781), .SEL(n10133), .F(
        n7165) );
  IV U10745 ( .A(n10134), .Z(n10133) );
  MUX U10746 ( .IN0(n9783), .IN1(data_mem_out_wire[586]), .SEL(n10134), .F(
        n7164) );
  MUX U10747 ( .IN0(n9784), .IN1(data_mem_out_wire[585]), .SEL(n10134), .F(
        n7163) );
  MUX U10748 ( .IN0(n9785), .IN1(data_mem_out_wire[584]), .SEL(n10134), .F(
        n7162) );
  AND U10749 ( .A(n10135), .B(n10136), .Z(n10134) );
  OR U10750 ( .A(n9788), .B(n10128), .Z(n10136) );
  MUX U10751 ( .IN0(data_mem_out_wire[583]), .IN1(data_in[7]), .SEL(n10137), 
        .F(n7161) );
  MUX U10752 ( .IN0(data_mem_out_wire[582]), .IN1(data_in[6]), .SEL(n10137), 
        .F(n7160) );
  MUX U10753 ( .IN0(data_mem_out_wire[581]), .IN1(data_in[5]), .SEL(n10137), 
        .F(n7159) );
  MUX U10754 ( .IN0(data_mem_out_wire[580]), .IN1(data_in[4]), .SEL(n10137), 
        .F(n7158) );
  MUX U10755 ( .IN0(data_mem_out_wire[579]), .IN1(data_in[3]), .SEL(n10137), 
        .F(n7157) );
  IV U10756 ( .A(n10138), .Z(n10137) );
  MUX U10757 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[578]), .SEL(n10138), 
        .F(n7156) );
  MUX U10758 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[577]), .SEL(n10138), 
        .F(n7155) );
  MUX U10759 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[576]), .SEL(n10138), 
        .F(n7154) );
  AND U10760 ( .A(n10135), .B(n10139), .Z(n10138) );
  NANDN U10761 ( .A(n10128), .B(n9792), .Z(n10139) );
  AND U10762 ( .A(n10140), .B(n10125), .Z(n10135) );
  NANDN U10763 ( .A(n10128), .B(n9796), .Z(n10125) );
  NANDN U10764 ( .A(n10128), .B(n9818), .Z(n10140) );
  NAND U10765 ( .A(n9838), .B(n10104), .Z(n10128) );
  MUX U10766 ( .IN0(n9746), .IN1(data_mem_out_wire[639]), .SEL(n10141), .F(
        n7153) );
  MUX U10767 ( .IN0(n9748), .IN1(data_mem_out_wire[638]), .SEL(n10141), .F(
        n7152) );
  MUX U10768 ( .IN0(n9749), .IN1(data_mem_out_wire[637]), .SEL(n10141), .F(
        n7151) );
  MUX U10769 ( .IN0(n9750), .IN1(data_mem_out_wire[636]), .SEL(n10141), .F(
        n7150) );
  MUX U10770 ( .IN0(n9751), .IN1(data_mem_out_wire[635]), .SEL(n10141), .F(
        n7149) );
  MUX U10771 ( .IN0(n9752), .IN1(data_mem_out_wire[634]), .SEL(n10141), .F(
        n7148) );
  MUX U10772 ( .IN0(n9753), .IN1(data_mem_out_wire[633]), .SEL(n10141), .F(
        n7147) );
  MUX U10773 ( .IN0(n9754), .IN1(data_mem_out_wire[632]), .SEL(n10141), .F(
        n7146) );
  AND U10774 ( .A(n10142), .B(n10143), .Z(n10141) );
  AND U10775 ( .A(n10144), .B(n10145), .Z(n10142) );
  OR U10776 ( .A(n9760), .B(n10146), .Z(n10145) );
  MUX U10777 ( .IN0(data_mem_out_wire[631]), .IN1(n9761), .SEL(n10147), .F(
        n7145) );
  MUX U10778 ( .IN0(data_mem_out_wire[630]), .IN1(n9763), .SEL(n10147), .F(
        n7144) );
  MUX U10779 ( .IN0(data_mem_out_wire[629]), .IN1(n9764), .SEL(n10147), .F(
        n7143) );
  MUX U10780 ( .IN0(data_mem_out_wire[628]), .IN1(n9765), .SEL(n10147), .F(
        n7142) );
  MUX U10781 ( .IN0(data_mem_out_wire[627]), .IN1(n9766), .SEL(n10147), .F(
        n7141) );
  IV U10782 ( .A(n10148), .Z(n10147) );
  MUX U10783 ( .IN0(n9768), .IN1(data_mem_out_wire[626]), .SEL(n10148), .F(
        n7140) );
  MUX U10784 ( .IN0(n9769), .IN1(data_mem_out_wire[625]), .SEL(n10148), .F(
        n7139) );
  MUX U10785 ( .IN0(n9770), .IN1(data_mem_out_wire[624]), .SEL(n10148), .F(
        n7138) );
  AND U10786 ( .A(n10149), .B(n10150), .Z(n10148) );
  OR U10787 ( .A(n9773), .B(n10146), .Z(n10150) );
  AND U10788 ( .A(n10144), .B(n10143), .Z(n10149) );
  NANDN U10789 ( .A(n10146), .B(n9809), .Z(n10144) );
  MUX U10790 ( .IN0(data_mem_out_wire[623]), .IN1(n9776), .SEL(n10151), .F(
        n7137) );
  MUX U10791 ( .IN0(data_mem_out_wire[622]), .IN1(n9778), .SEL(n10151), .F(
        n7136) );
  MUX U10792 ( .IN0(data_mem_out_wire[621]), .IN1(n9779), .SEL(n10151), .F(
        n7135) );
  MUX U10793 ( .IN0(data_mem_out_wire[620]), .IN1(n9780), .SEL(n10151), .F(
        n7134) );
  MUX U10794 ( .IN0(data_mem_out_wire[619]), .IN1(n9781), .SEL(n10151), .F(
        n7133) );
  IV U10795 ( .A(n10152), .Z(n10151) );
  MUX U10796 ( .IN0(n9783), .IN1(data_mem_out_wire[618]), .SEL(n10152), .F(
        n7132) );
  MUX U10797 ( .IN0(n9784), .IN1(data_mem_out_wire[617]), .SEL(n10152), .F(
        n7131) );
  MUX U10798 ( .IN0(n9785), .IN1(data_mem_out_wire[616]), .SEL(n10152), .F(
        n7130) );
  AND U10799 ( .A(n10153), .B(n10154), .Z(n10152) );
  OR U10800 ( .A(n9788), .B(n10146), .Z(n10154) );
  MUX U10801 ( .IN0(data_mem_out_wire[615]), .IN1(data_in[7]), .SEL(n10155), 
        .F(n7129) );
  MUX U10802 ( .IN0(data_mem_out_wire[614]), .IN1(data_in[6]), .SEL(n10155), 
        .F(n7128) );
  MUX U10803 ( .IN0(data_mem_out_wire[613]), .IN1(data_in[5]), .SEL(n10155), 
        .F(n7127) );
  MUX U10804 ( .IN0(data_mem_out_wire[612]), .IN1(data_in[4]), .SEL(n10155), 
        .F(n7126) );
  MUX U10805 ( .IN0(data_mem_out_wire[611]), .IN1(data_in[3]), .SEL(n10155), 
        .F(n7125) );
  IV U10806 ( .A(n10156), .Z(n10155) );
  MUX U10807 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[610]), .SEL(n10156), 
        .F(n7124) );
  MUX U10808 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[609]), .SEL(n10156), 
        .F(n7123) );
  MUX U10809 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[608]), .SEL(n10156), 
        .F(n7122) );
  AND U10810 ( .A(n10153), .B(n10157), .Z(n10156) );
  NANDN U10811 ( .A(n10146), .B(n9792), .Z(n10157) );
  AND U10812 ( .A(n10158), .B(n10143), .Z(n10153) );
  NANDN U10813 ( .A(n10146), .B(n9796), .Z(n10143) );
  NANDN U10814 ( .A(n10146), .B(n9818), .Z(n10158) );
  NAND U10815 ( .A(n9862), .B(n10104), .Z(n10146) );
  MUX U10816 ( .IN0(n9746), .IN1(data_mem_out_wire[671]), .SEL(n10159), .F(
        n7121) );
  MUX U10817 ( .IN0(n9748), .IN1(data_mem_out_wire[670]), .SEL(n10159), .F(
        n7120) );
  MUX U10818 ( .IN0(n9749), .IN1(data_mem_out_wire[669]), .SEL(n10159), .F(
        n7119) );
  MUX U10819 ( .IN0(n9750), .IN1(data_mem_out_wire[668]), .SEL(n10159), .F(
        n7118) );
  MUX U10820 ( .IN0(n9751), .IN1(data_mem_out_wire[667]), .SEL(n10159), .F(
        n7117) );
  MUX U10821 ( .IN0(n9752), .IN1(data_mem_out_wire[666]), .SEL(n10159), .F(
        n7116) );
  MUX U10822 ( .IN0(n9753), .IN1(data_mem_out_wire[665]), .SEL(n10159), .F(
        n7115) );
  MUX U10823 ( .IN0(n9754), .IN1(data_mem_out_wire[664]), .SEL(n10159), .F(
        n7114) );
  AND U10824 ( .A(n10160), .B(n10161), .Z(n10159) );
  AND U10825 ( .A(n10162), .B(n10163), .Z(n10160) );
  OR U10826 ( .A(n9760), .B(n10164), .Z(n10163) );
  MUX U10827 ( .IN0(data_mem_out_wire[663]), .IN1(n9761), .SEL(n10165), .F(
        n7113) );
  MUX U10828 ( .IN0(data_mem_out_wire[662]), .IN1(n9763), .SEL(n10165), .F(
        n7112) );
  MUX U10829 ( .IN0(data_mem_out_wire[661]), .IN1(n9764), .SEL(n10165), .F(
        n7111) );
  MUX U10830 ( .IN0(data_mem_out_wire[660]), .IN1(n9765), .SEL(n10165), .F(
        n7110) );
  MUX U10831 ( .IN0(data_mem_out_wire[659]), .IN1(n9766), .SEL(n10165), .F(
        n7109) );
  IV U10832 ( .A(n10166), .Z(n10165) );
  MUX U10833 ( .IN0(n9768), .IN1(data_mem_out_wire[658]), .SEL(n10166), .F(
        n7108) );
  MUX U10834 ( .IN0(n9769), .IN1(data_mem_out_wire[657]), .SEL(n10166), .F(
        n7107) );
  MUX U10835 ( .IN0(n9770), .IN1(data_mem_out_wire[656]), .SEL(n10166), .F(
        n7106) );
  AND U10836 ( .A(n10167), .B(n10168), .Z(n10166) );
  OR U10837 ( .A(n9773), .B(n10164), .Z(n10168) );
  AND U10838 ( .A(n10162), .B(n10161), .Z(n10167) );
  NANDN U10839 ( .A(n10164), .B(n9809), .Z(n10162) );
  MUX U10840 ( .IN0(data_mem_out_wire[655]), .IN1(n9776), .SEL(n10169), .F(
        n7105) );
  MUX U10841 ( .IN0(data_mem_out_wire[654]), .IN1(n9778), .SEL(n10169), .F(
        n7104) );
  MUX U10842 ( .IN0(data_mem_out_wire[653]), .IN1(n9779), .SEL(n10169), .F(
        n7103) );
  MUX U10843 ( .IN0(data_mem_out_wire[652]), .IN1(n9780), .SEL(n10169), .F(
        n7102) );
  MUX U10844 ( .IN0(data_mem_out_wire[651]), .IN1(n9781), .SEL(n10169), .F(
        n7101) );
  IV U10845 ( .A(n10170), .Z(n10169) );
  MUX U10846 ( .IN0(n9783), .IN1(data_mem_out_wire[650]), .SEL(n10170), .F(
        n7100) );
  MUX U10847 ( .IN0(n9784), .IN1(data_mem_out_wire[649]), .SEL(n10170), .F(
        n7099) );
  MUX U10848 ( .IN0(n9785), .IN1(data_mem_out_wire[648]), .SEL(n10170), .F(
        n7098) );
  AND U10849 ( .A(n10171), .B(n10172), .Z(n10170) );
  OR U10850 ( .A(n9788), .B(n10164), .Z(n10172) );
  MUX U10851 ( .IN0(data_mem_out_wire[647]), .IN1(data_in[7]), .SEL(n10173), 
        .F(n7097) );
  MUX U10852 ( .IN0(data_mem_out_wire[646]), .IN1(data_in[6]), .SEL(n10173), 
        .F(n7096) );
  MUX U10853 ( .IN0(data_mem_out_wire[645]), .IN1(data_in[5]), .SEL(n10173), 
        .F(n7095) );
  MUX U10854 ( .IN0(data_mem_out_wire[644]), .IN1(data_in[4]), .SEL(n10173), 
        .F(n7094) );
  MUX U10855 ( .IN0(data_mem_out_wire[643]), .IN1(data_in[3]), .SEL(n10173), 
        .F(n7093) );
  IV U10856 ( .A(n10174), .Z(n10173) );
  MUX U10857 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[642]), .SEL(n10174), 
        .F(n7092) );
  MUX U10858 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[641]), .SEL(n10174), 
        .F(n7091) );
  MUX U10859 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[640]), .SEL(n10174), 
        .F(n7090) );
  AND U10860 ( .A(n10171), .B(n10175), .Z(n10174) );
  NANDN U10861 ( .A(n10164), .B(n9792), .Z(n10175) );
  AND U10862 ( .A(n10176), .B(n10161), .Z(n10171) );
  NANDN U10863 ( .A(n10164), .B(n9796), .Z(n10161) );
  NANDN U10864 ( .A(n10164), .B(n9818), .Z(n10176) );
  NAND U10865 ( .A(n9881), .B(n10104), .Z(n10164) );
  MUX U10866 ( .IN0(n9746), .IN1(data_mem_out_wire[703]), .SEL(n10177), .F(
        n7089) );
  MUX U10867 ( .IN0(n9748), .IN1(data_mem_out_wire[702]), .SEL(n10177), .F(
        n7088) );
  MUX U10868 ( .IN0(n9749), .IN1(data_mem_out_wire[701]), .SEL(n10177), .F(
        n7087) );
  MUX U10869 ( .IN0(n9750), .IN1(data_mem_out_wire[700]), .SEL(n10177), .F(
        n7086) );
  MUX U10870 ( .IN0(n9751), .IN1(data_mem_out_wire[699]), .SEL(n10177), .F(
        n7085) );
  MUX U10871 ( .IN0(n9752), .IN1(data_mem_out_wire[698]), .SEL(n10177), .F(
        n7084) );
  MUX U10872 ( .IN0(n9753), .IN1(data_mem_out_wire[697]), .SEL(n10177), .F(
        n7083) );
  MUX U10873 ( .IN0(n9754), .IN1(data_mem_out_wire[696]), .SEL(n10177), .F(
        n7082) );
  AND U10874 ( .A(n10178), .B(n10179), .Z(n10177) );
  AND U10875 ( .A(n10180), .B(n10181), .Z(n10178) );
  OR U10876 ( .A(n9760), .B(n10182), .Z(n10181) );
  MUX U10877 ( .IN0(data_mem_out_wire[695]), .IN1(n9761), .SEL(n10183), .F(
        n7081) );
  MUX U10878 ( .IN0(data_mem_out_wire[694]), .IN1(n9763), .SEL(n10183), .F(
        n7080) );
  MUX U10879 ( .IN0(data_mem_out_wire[693]), .IN1(n9764), .SEL(n10183), .F(
        n7079) );
  MUX U10880 ( .IN0(data_mem_out_wire[692]), .IN1(n9765), .SEL(n10183), .F(
        n7078) );
  MUX U10881 ( .IN0(data_mem_out_wire[691]), .IN1(n9766), .SEL(n10183), .F(
        n7077) );
  IV U10882 ( .A(n10184), .Z(n10183) );
  MUX U10883 ( .IN0(n9768), .IN1(data_mem_out_wire[690]), .SEL(n10184), .F(
        n7076) );
  MUX U10884 ( .IN0(n9769), .IN1(data_mem_out_wire[689]), .SEL(n10184), .F(
        n7075) );
  MUX U10885 ( .IN0(n9770), .IN1(data_mem_out_wire[688]), .SEL(n10184), .F(
        n7074) );
  AND U10886 ( .A(n10185), .B(n10186), .Z(n10184) );
  OR U10887 ( .A(n9773), .B(n10182), .Z(n10186) );
  AND U10888 ( .A(n10180), .B(n10179), .Z(n10185) );
  NANDN U10889 ( .A(n10182), .B(n9809), .Z(n10180) );
  MUX U10890 ( .IN0(data_mem_out_wire[687]), .IN1(n9776), .SEL(n10187), .F(
        n7073) );
  MUX U10891 ( .IN0(data_mem_out_wire[686]), .IN1(n9778), .SEL(n10187), .F(
        n7072) );
  MUX U10892 ( .IN0(data_mem_out_wire[685]), .IN1(n9779), .SEL(n10187), .F(
        n7071) );
  MUX U10893 ( .IN0(data_mem_out_wire[684]), .IN1(n9780), .SEL(n10187), .F(
        n7070) );
  MUX U10894 ( .IN0(data_mem_out_wire[683]), .IN1(n9781), .SEL(n10187), .F(
        n7069) );
  IV U10895 ( .A(n10188), .Z(n10187) );
  MUX U10896 ( .IN0(n9783), .IN1(data_mem_out_wire[682]), .SEL(n10188), .F(
        n7068) );
  MUX U10897 ( .IN0(n9784), .IN1(data_mem_out_wire[681]), .SEL(n10188), .F(
        n7067) );
  MUX U10898 ( .IN0(n9785), .IN1(data_mem_out_wire[680]), .SEL(n10188), .F(
        n7066) );
  AND U10899 ( .A(n10189), .B(n10190), .Z(n10188) );
  OR U10900 ( .A(n9788), .B(n10182), .Z(n10190) );
  MUX U10901 ( .IN0(data_mem_out_wire[679]), .IN1(data_in[7]), .SEL(n10191), 
        .F(n7065) );
  MUX U10902 ( .IN0(data_mem_out_wire[678]), .IN1(data_in[6]), .SEL(n10191), 
        .F(n7064) );
  MUX U10903 ( .IN0(data_mem_out_wire[677]), .IN1(data_in[5]), .SEL(n10191), 
        .F(n7063) );
  MUX U10904 ( .IN0(data_mem_out_wire[676]), .IN1(data_in[4]), .SEL(n10191), 
        .F(n7062) );
  MUX U10905 ( .IN0(data_mem_out_wire[675]), .IN1(data_in[3]), .SEL(n10191), 
        .F(n7061) );
  IV U10906 ( .A(n10192), .Z(n10191) );
  MUX U10907 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[674]), .SEL(n10192), 
        .F(n7060) );
  MUX U10908 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[673]), .SEL(n10192), 
        .F(n7059) );
  MUX U10909 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[672]), .SEL(n10192), 
        .F(n7058) );
  AND U10910 ( .A(n10189), .B(n10193), .Z(n10192) );
  NANDN U10911 ( .A(n10182), .B(n9792), .Z(n10193) );
  AND U10912 ( .A(n10194), .B(n10179), .Z(n10189) );
  NANDN U10913 ( .A(n10182), .B(n9796), .Z(n10179) );
  NANDN U10914 ( .A(n10182), .B(n9818), .Z(n10194) );
  NAND U10915 ( .A(n9900), .B(n10104), .Z(n10182) );
  MUX U10916 ( .IN0(n9746), .IN1(data_mem_out_wire[735]), .SEL(n10195), .F(
        n7057) );
  MUX U10917 ( .IN0(n9748), .IN1(data_mem_out_wire[734]), .SEL(n10195), .F(
        n7056) );
  MUX U10918 ( .IN0(n9749), .IN1(data_mem_out_wire[733]), .SEL(n10195), .F(
        n7055) );
  MUX U10919 ( .IN0(n9750), .IN1(data_mem_out_wire[732]), .SEL(n10195), .F(
        n7054) );
  MUX U10920 ( .IN0(n9751), .IN1(data_mem_out_wire[731]), .SEL(n10195), .F(
        n7053) );
  MUX U10921 ( .IN0(n9752), .IN1(data_mem_out_wire[730]), .SEL(n10195), .F(
        n7052) );
  MUX U10922 ( .IN0(n9753), .IN1(data_mem_out_wire[729]), .SEL(n10195), .F(
        n7051) );
  MUX U10923 ( .IN0(n9754), .IN1(data_mem_out_wire[728]), .SEL(n10195), .F(
        n7050) );
  AND U10924 ( .A(n10196), .B(n10197), .Z(n10195) );
  AND U10925 ( .A(n10198), .B(n10199), .Z(n10196) );
  OR U10926 ( .A(n9760), .B(n10200), .Z(n10199) );
  MUX U10927 ( .IN0(data_mem_out_wire[727]), .IN1(n9761), .SEL(n10201), .F(
        n7049) );
  MUX U10928 ( .IN0(data_mem_out_wire[726]), .IN1(n9763), .SEL(n10201), .F(
        n7048) );
  MUX U10929 ( .IN0(data_mem_out_wire[725]), .IN1(n9764), .SEL(n10201), .F(
        n7047) );
  MUX U10930 ( .IN0(data_mem_out_wire[724]), .IN1(n9765), .SEL(n10201), .F(
        n7046) );
  MUX U10931 ( .IN0(data_mem_out_wire[723]), .IN1(n9766), .SEL(n10201), .F(
        n7045) );
  IV U10932 ( .A(n10202), .Z(n10201) );
  MUX U10933 ( .IN0(n9768), .IN1(data_mem_out_wire[722]), .SEL(n10202), .F(
        n7044) );
  MUX U10934 ( .IN0(n9769), .IN1(data_mem_out_wire[721]), .SEL(n10202), .F(
        n7043) );
  MUX U10935 ( .IN0(n9770), .IN1(data_mem_out_wire[720]), .SEL(n10202), .F(
        n7042) );
  AND U10936 ( .A(n10203), .B(n10204), .Z(n10202) );
  OR U10937 ( .A(n9773), .B(n10200), .Z(n10204) );
  AND U10938 ( .A(n10198), .B(n10197), .Z(n10203) );
  NANDN U10939 ( .A(n10200), .B(n9809), .Z(n10198) );
  MUX U10940 ( .IN0(data_mem_out_wire[719]), .IN1(n9776), .SEL(n10205), .F(
        n7041) );
  MUX U10941 ( .IN0(data_mem_out_wire[718]), .IN1(n9778), .SEL(n10205), .F(
        n7040) );
  MUX U10942 ( .IN0(data_mem_out_wire[717]), .IN1(n9779), .SEL(n10205), .F(
        n7039) );
  MUX U10943 ( .IN0(data_mem_out_wire[716]), .IN1(n9780), .SEL(n10205), .F(
        n7038) );
  MUX U10944 ( .IN0(data_mem_out_wire[715]), .IN1(n9781), .SEL(n10205), .F(
        n7037) );
  IV U10945 ( .A(n10206), .Z(n10205) );
  MUX U10946 ( .IN0(n9783), .IN1(data_mem_out_wire[714]), .SEL(n10206), .F(
        n7036) );
  MUX U10947 ( .IN0(n9784), .IN1(data_mem_out_wire[713]), .SEL(n10206), .F(
        n7035) );
  MUX U10948 ( .IN0(n9785), .IN1(data_mem_out_wire[712]), .SEL(n10206), .F(
        n7034) );
  AND U10949 ( .A(n10207), .B(n10208), .Z(n10206) );
  OR U10950 ( .A(n9788), .B(n10200), .Z(n10208) );
  MUX U10951 ( .IN0(data_mem_out_wire[711]), .IN1(data_in[7]), .SEL(n10209), 
        .F(n7033) );
  MUX U10952 ( .IN0(data_mem_out_wire[710]), .IN1(data_in[6]), .SEL(n10209), 
        .F(n7032) );
  MUX U10953 ( .IN0(data_mem_out_wire[709]), .IN1(data_in[5]), .SEL(n10209), 
        .F(n7031) );
  MUX U10954 ( .IN0(data_mem_out_wire[708]), .IN1(data_in[4]), .SEL(n10209), 
        .F(n7030) );
  MUX U10955 ( .IN0(data_mem_out_wire[707]), .IN1(data_in[3]), .SEL(n10209), 
        .F(n7029) );
  IV U10956 ( .A(n10210), .Z(n10209) );
  MUX U10957 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[706]), .SEL(n10210), 
        .F(n7028) );
  MUX U10958 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[705]), .SEL(n10210), 
        .F(n7027) );
  MUX U10959 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[704]), .SEL(n10210), 
        .F(n7026) );
  AND U10960 ( .A(n10207), .B(n10211), .Z(n10210) );
  NANDN U10961 ( .A(n10200), .B(n9792), .Z(n10211) );
  AND U10962 ( .A(n10212), .B(n10197), .Z(n10207) );
  NANDN U10963 ( .A(n10200), .B(n9796), .Z(n10197) );
  NANDN U10964 ( .A(n10200), .B(n9818), .Z(n10212) );
  NAND U10965 ( .A(n9919), .B(n10104), .Z(n10200) );
  MUX U10966 ( .IN0(n9746), .IN1(data_mem_out_wire[767]), .SEL(n10213), .F(
        n7025) );
  MUX U10967 ( .IN0(n9748), .IN1(data_mem_out_wire[766]), .SEL(n10213), .F(
        n7024) );
  MUX U10968 ( .IN0(n9749), .IN1(data_mem_out_wire[765]), .SEL(n10213), .F(
        n7023) );
  MUX U10969 ( .IN0(n9750), .IN1(data_mem_out_wire[764]), .SEL(n10213), .F(
        n7022) );
  MUX U10970 ( .IN0(n9751), .IN1(data_mem_out_wire[763]), .SEL(n10213), .F(
        n7021) );
  MUX U10971 ( .IN0(n9752), .IN1(data_mem_out_wire[762]), .SEL(n10213), .F(
        n7020) );
  MUX U10972 ( .IN0(n9753), .IN1(data_mem_out_wire[761]), .SEL(n10213), .F(
        n7019) );
  MUX U10973 ( .IN0(n9754), .IN1(data_mem_out_wire[760]), .SEL(n10213), .F(
        n7018) );
  AND U10974 ( .A(n10214), .B(n10215), .Z(n10213) );
  AND U10975 ( .A(n10216), .B(n10217), .Z(n10214) );
  OR U10976 ( .A(n9760), .B(n10218), .Z(n10217) );
  MUX U10977 ( .IN0(data_mem_out_wire[759]), .IN1(n9761), .SEL(n10219), .F(
        n7017) );
  MUX U10978 ( .IN0(data_mem_out_wire[758]), .IN1(n9763), .SEL(n10219), .F(
        n7016) );
  MUX U10979 ( .IN0(data_mem_out_wire[757]), .IN1(n9764), .SEL(n10219), .F(
        n7015) );
  MUX U10980 ( .IN0(data_mem_out_wire[756]), .IN1(n9765), .SEL(n10219), .F(
        n7014) );
  MUX U10981 ( .IN0(data_mem_out_wire[755]), .IN1(n9766), .SEL(n10219), .F(
        n7013) );
  IV U10982 ( .A(n10220), .Z(n10219) );
  MUX U10983 ( .IN0(n9768), .IN1(data_mem_out_wire[754]), .SEL(n10220), .F(
        n7012) );
  MUX U10984 ( .IN0(n9769), .IN1(data_mem_out_wire[753]), .SEL(n10220), .F(
        n7011) );
  MUX U10985 ( .IN0(n9770), .IN1(data_mem_out_wire[752]), .SEL(n10220), .F(
        n7010) );
  AND U10986 ( .A(n10221), .B(n10222), .Z(n10220) );
  OR U10987 ( .A(n9773), .B(n10218), .Z(n10222) );
  AND U10988 ( .A(n10216), .B(n10215), .Z(n10221) );
  NANDN U10989 ( .A(n10218), .B(n9809), .Z(n10216) );
  MUX U10990 ( .IN0(data_mem_out_wire[751]), .IN1(n9776), .SEL(n10223), .F(
        n7009) );
  MUX U10991 ( .IN0(data_mem_out_wire[750]), .IN1(n9778), .SEL(n10223), .F(
        n7008) );
  MUX U10992 ( .IN0(data_mem_out_wire[749]), .IN1(n9779), .SEL(n10223), .F(
        n7007) );
  MUX U10993 ( .IN0(data_mem_out_wire[748]), .IN1(n9780), .SEL(n10223), .F(
        n7006) );
  MUX U10994 ( .IN0(data_mem_out_wire[747]), .IN1(n9781), .SEL(n10223), .F(
        n7005) );
  IV U10995 ( .A(n10224), .Z(n10223) );
  MUX U10996 ( .IN0(n9783), .IN1(data_mem_out_wire[746]), .SEL(n10224), .F(
        n7004) );
  MUX U10997 ( .IN0(n9784), .IN1(data_mem_out_wire[745]), .SEL(n10224), .F(
        n7003) );
  MUX U10998 ( .IN0(n9785), .IN1(data_mem_out_wire[744]), .SEL(n10224), .F(
        n7002) );
  AND U10999 ( .A(n10225), .B(n10226), .Z(n10224) );
  OR U11000 ( .A(n9788), .B(n10218), .Z(n10226) );
  MUX U11001 ( .IN0(data_mem_out_wire[743]), .IN1(data_in[7]), .SEL(n10227), 
        .F(n7001) );
  MUX U11002 ( .IN0(data_mem_out_wire[742]), .IN1(data_in[6]), .SEL(n10227), 
        .F(n7000) );
  MUX U11003 ( .IN0(data_mem_out_wire[741]), .IN1(data_in[5]), .SEL(n10227), 
        .F(n6999) );
  MUX U11004 ( .IN0(data_mem_out_wire[740]), .IN1(data_in[4]), .SEL(n10227), 
        .F(n6998) );
  MUX U11005 ( .IN0(data_mem_out_wire[739]), .IN1(data_in[3]), .SEL(n10227), 
        .F(n6997) );
  IV U11006 ( .A(n10228), .Z(n10227) );
  MUX U11007 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[738]), .SEL(n10228), 
        .F(n6996) );
  MUX U11008 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[737]), .SEL(n10228), 
        .F(n6995) );
  MUX U11009 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[736]), .SEL(n10228), 
        .F(n6994) );
  AND U11010 ( .A(n10225), .B(n10229), .Z(n10228) );
  NANDN U11011 ( .A(n10218), .B(n9792), .Z(n10229) );
  AND U11012 ( .A(n10230), .B(n10215), .Z(n10225) );
  NANDN U11013 ( .A(n10218), .B(n9796), .Z(n10215) );
  NANDN U11014 ( .A(n10218), .B(n9818), .Z(n10230) );
  NAND U11015 ( .A(n10104), .B(n9938), .Z(n10218) );
  ANDN U11016 ( .B(n10231), .A(N42), .Z(n10104) );
  MUX U11017 ( .IN0(n9746), .IN1(data_mem_out_wire[799]), .SEL(n10232), .F(
        n6993) );
  MUX U11018 ( .IN0(n9748), .IN1(data_mem_out_wire[798]), .SEL(n10232), .F(
        n6992) );
  MUX U11019 ( .IN0(n9749), .IN1(data_mem_out_wire[797]), .SEL(n10232), .F(
        n6991) );
  MUX U11020 ( .IN0(n9750), .IN1(data_mem_out_wire[796]), .SEL(n10232), .F(
        n6990) );
  MUX U11021 ( .IN0(n9751), .IN1(data_mem_out_wire[795]), .SEL(n10232), .F(
        n6989) );
  MUX U11022 ( .IN0(n9752), .IN1(data_mem_out_wire[794]), .SEL(n10232), .F(
        n6988) );
  MUX U11023 ( .IN0(n9753), .IN1(data_mem_out_wire[793]), .SEL(n10232), .F(
        n6987) );
  MUX U11024 ( .IN0(n9754), .IN1(data_mem_out_wire[792]), .SEL(n10232), .F(
        n6986) );
  AND U11025 ( .A(n10233), .B(n10234), .Z(n10232) );
  AND U11026 ( .A(n10235), .B(n10236), .Z(n10233) );
  OR U11027 ( .A(n9760), .B(n10237), .Z(n10236) );
  MUX U11028 ( .IN0(data_mem_out_wire[791]), .IN1(n9761), .SEL(n10238), .F(
        n6985) );
  MUX U11029 ( .IN0(data_mem_out_wire[790]), .IN1(n9763), .SEL(n10238), .F(
        n6984) );
  MUX U11030 ( .IN0(data_mem_out_wire[789]), .IN1(n9764), .SEL(n10238), .F(
        n6983) );
  MUX U11031 ( .IN0(data_mem_out_wire[788]), .IN1(n9765), .SEL(n10238), .F(
        n6982) );
  MUX U11032 ( .IN0(data_mem_out_wire[787]), .IN1(n9766), .SEL(n10238), .F(
        n6981) );
  IV U11033 ( .A(n10239), .Z(n10238) );
  MUX U11034 ( .IN0(n9768), .IN1(data_mem_out_wire[786]), .SEL(n10239), .F(
        n6980) );
  MUX U11035 ( .IN0(n9769), .IN1(data_mem_out_wire[785]), .SEL(n10239), .F(
        n6979) );
  MUX U11036 ( .IN0(n9770), .IN1(data_mem_out_wire[784]), .SEL(n10239), .F(
        n6978) );
  AND U11037 ( .A(n10240), .B(n10241), .Z(n10239) );
  OR U11038 ( .A(n9773), .B(n10237), .Z(n10241) );
  AND U11039 ( .A(n10235), .B(n10234), .Z(n10240) );
  NANDN U11040 ( .A(n10237), .B(n9809), .Z(n10235) );
  MUX U11041 ( .IN0(data_mem_out_wire[783]), .IN1(n9776), .SEL(n10242), .F(
        n6977) );
  MUX U11042 ( .IN0(data_mem_out_wire[782]), .IN1(n9778), .SEL(n10242), .F(
        n6976) );
  MUX U11043 ( .IN0(data_mem_out_wire[781]), .IN1(n9779), .SEL(n10242), .F(
        n6975) );
  MUX U11044 ( .IN0(data_mem_out_wire[780]), .IN1(n9780), .SEL(n10242), .F(
        n6974) );
  MUX U11045 ( .IN0(data_mem_out_wire[779]), .IN1(n9781), .SEL(n10242), .F(
        n6973) );
  IV U11046 ( .A(n10243), .Z(n10242) );
  MUX U11047 ( .IN0(n9783), .IN1(data_mem_out_wire[778]), .SEL(n10243), .F(
        n6972) );
  MUX U11048 ( .IN0(n9784), .IN1(data_mem_out_wire[777]), .SEL(n10243), .F(
        n6971) );
  MUX U11049 ( .IN0(n9785), .IN1(data_mem_out_wire[776]), .SEL(n10243), .F(
        n6970) );
  AND U11050 ( .A(n10244), .B(n10245), .Z(n10243) );
  OR U11051 ( .A(n9788), .B(n10237), .Z(n10245) );
  MUX U11052 ( .IN0(data_mem_out_wire[775]), .IN1(data_in[7]), .SEL(n10246), 
        .F(n6969) );
  MUX U11053 ( .IN0(data_mem_out_wire[774]), .IN1(data_in[6]), .SEL(n10246), 
        .F(n6968) );
  MUX U11054 ( .IN0(data_mem_out_wire[773]), .IN1(data_in[5]), .SEL(n10246), 
        .F(n6967) );
  MUX U11055 ( .IN0(data_mem_out_wire[772]), .IN1(data_in[4]), .SEL(n10246), 
        .F(n6966) );
  MUX U11056 ( .IN0(data_mem_out_wire[771]), .IN1(data_in[3]), .SEL(n10246), 
        .F(n6965) );
  IV U11057 ( .A(n10247), .Z(n10246) );
  MUX U11058 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[770]), .SEL(n10247), 
        .F(n6964) );
  MUX U11059 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[769]), .SEL(n10247), 
        .F(n6963) );
  MUX U11060 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[768]), .SEL(n10247), 
        .F(n6962) );
  AND U11061 ( .A(n10244), .B(n10248), .Z(n10247) );
  NANDN U11062 ( .A(n10237), .B(n9792), .Z(n10248) );
  AND U11063 ( .A(n10249), .B(n10234), .Z(n10244) );
  NANDN U11064 ( .A(n10237), .B(n9796), .Z(n10234) );
  NANDN U11065 ( .A(n10237), .B(n9818), .Z(n10249) );
  NAND U11066 ( .A(n9798), .B(n10250), .Z(n10237) );
  MUX U11067 ( .IN0(n9746), .IN1(data_mem_out_wire[831]), .SEL(n10251), .F(
        n6961) );
  MUX U11068 ( .IN0(n9748), .IN1(data_mem_out_wire[830]), .SEL(n10251), .F(
        n6960) );
  MUX U11069 ( .IN0(n9749), .IN1(data_mem_out_wire[829]), .SEL(n10251), .F(
        n6959) );
  MUX U11070 ( .IN0(n9750), .IN1(data_mem_out_wire[828]), .SEL(n10251), .F(
        n6958) );
  MUX U11071 ( .IN0(n9751), .IN1(data_mem_out_wire[827]), .SEL(n10251), .F(
        n6957) );
  MUX U11072 ( .IN0(n9752), .IN1(data_mem_out_wire[826]), .SEL(n10251), .F(
        n6956) );
  MUX U11073 ( .IN0(n9753), .IN1(data_mem_out_wire[825]), .SEL(n10251), .F(
        n6955) );
  MUX U11074 ( .IN0(n9754), .IN1(data_mem_out_wire[824]), .SEL(n10251), .F(
        n6954) );
  AND U11075 ( .A(n10252), .B(n10253), .Z(n10251) );
  AND U11076 ( .A(n10254), .B(n10255), .Z(n10252) );
  OR U11077 ( .A(n9760), .B(n10256), .Z(n10255) );
  MUX U11078 ( .IN0(data_mem_out_wire[823]), .IN1(n9761), .SEL(n10257), .F(
        n6953) );
  MUX U11079 ( .IN0(data_mem_out_wire[822]), .IN1(n9763), .SEL(n10257), .F(
        n6952) );
  MUX U11080 ( .IN0(data_mem_out_wire[821]), .IN1(n9764), .SEL(n10257), .F(
        n6951) );
  MUX U11081 ( .IN0(data_mem_out_wire[820]), .IN1(n9765), .SEL(n10257), .F(
        n6950) );
  MUX U11082 ( .IN0(data_mem_out_wire[819]), .IN1(n9766), .SEL(n10257), .F(
        n6949) );
  IV U11083 ( .A(n10258), .Z(n10257) );
  MUX U11084 ( .IN0(n9768), .IN1(data_mem_out_wire[818]), .SEL(n10258), .F(
        n6948) );
  MUX U11085 ( .IN0(n9769), .IN1(data_mem_out_wire[817]), .SEL(n10258), .F(
        n6947) );
  MUX U11086 ( .IN0(n9770), .IN1(data_mem_out_wire[816]), .SEL(n10258), .F(
        n6946) );
  AND U11087 ( .A(n10259), .B(n10260), .Z(n10258) );
  OR U11088 ( .A(n9773), .B(n10256), .Z(n10260) );
  AND U11089 ( .A(n10254), .B(n10253), .Z(n10259) );
  NANDN U11090 ( .A(n10256), .B(n9809), .Z(n10254) );
  MUX U11091 ( .IN0(data_mem_out_wire[815]), .IN1(n9776), .SEL(n10261), .F(
        n6945) );
  MUX U11092 ( .IN0(data_mem_out_wire[814]), .IN1(n9778), .SEL(n10261), .F(
        n6944) );
  MUX U11093 ( .IN0(data_mem_out_wire[813]), .IN1(n9779), .SEL(n10261), .F(
        n6943) );
  MUX U11094 ( .IN0(data_mem_out_wire[812]), .IN1(n9780), .SEL(n10261), .F(
        n6942) );
  MUX U11095 ( .IN0(data_mem_out_wire[811]), .IN1(n9781), .SEL(n10261), .F(
        n6941) );
  IV U11096 ( .A(n10262), .Z(n10261) );
  MUX U11097 ( .IN0(n9783), .IN1(data_mem_out_wire[810]), .SEL(n10262), .F(
        n6940) );
  MUX U11098 ( .IN0(n9784), .IN1(data_mem_out_wire[809]), .SEL(n10262), .F(
        n6939) );
  MUX U11099 ( .IN0(n9785), .IN1(data_mem_out_wire[808]), .SEL(n10262), .F(
        n6938) );
  AND U11100 ( .A(n10263), .B(n10264), .Z(n10262) );
  OR U11101 ( .A(n9788), .B(n10256), .Z(n10264) );
  MUX U11102 ( .IN0(data_mem_out_wire[807]), .IN1(data_in[7]), .SEL(n10265), 
        .F(n6937) );
  MUX U11103 ( .IN0(data_mem_out_wire[806]), .IN1(data_in[6]), .SEL(n10265), 
        .F(n6936) );
  MUX U11104 ( .IN0(data_mem_out_wire[805]), .IN1(data_in[5]), .SEL(n10265), 
        .F(n6935) );
  MUX U11105 ( .IN0(data_mem_out_wire[804]), .IN1(data_in[4]), .SEL(n10265), 
        .F(n6934) );
  MUX U11106 ( .IN0(data_mem_out_wire[803]), .IN1(data_in[3]), .SEL(n10265), 
        .F(n6933) );
  IV U11107 ( .A(n10266), .Z(n10265) );
  MUX U11108 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[802]), .SEL(n10266), 
        .F(n6932) );
  MUX U11109 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[801]), .SEL(n10266), 
        .F(n6931) );
  MUX U11110 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[800]), .SEL(n10266), 
        .F(n6930) );
  AND U11111 ( .A(n10263), .B(n10267), .Z(n10266) );
  NANDN U11112 ( .A(n10256), .B(n9792), .Z(n10267) );
  AND U11113 ( .A(n10268), .B(n10253), .Z(n10263) );
  NANDN U11114 ( .A(n10256), .B(n9796), .Z(n10253) );
  NANDN U11115 ( .A(n10256), .B(n9818), .Z(n10268) );
  NAND U11116 ( .A(n9819), .B(n10250), .Z(n10256) );
  MUX U11117 ( .IN0(n9746), .IN1(data_mem_out_wire[863]), .SEL(n10269), .F(
        n6929) );
  MUX U11118 ( .IN0(n9748), .IN1(data_mem_out_wire[862]), .SEL(n10269), .F(
        n6928) );
  MUX U11119 ( .IN0(n9749), .IN1(data_mem_out_wire[861]), .SEL(n10269), .F(
        n6927) );
  MUX U11120 ( .IN0(n9750), .IN1(data_mem_out_wire[860]), .SEL(n10269), .F(
        n6926) );
  MUX U11121 ( .IN0(n9751), .IN1(data_mem_out_wire[859]), .SEL(n10269), .F(
        n6925) );
  MUX U11122 ( .IN0(n9752), .IN1(data_mem_out_wire[858]), .SEL(n10269), .F(
        n6924) );
  MUX U11123 ( .IN0(n9753), .IN1(data_mem_out_wire[857]), .SEL(n10269), .F(
        n6923) );
  MUX U11124 ( .IN0(n9754), .IN1(data_mem_out_wire[856]), .SEL(n10269), .F(
        n6922) );
  AND U11125 ( .A(n10270), .B(n10271), .Z(n10269) );
  AND U11126 ( .A(n10272), .B(n10273), .Z(n10270) );
  OR U11127 ( .A(n9760), .B(n10274), .Z(n10273) );
  MUX U11128 ( .IN0(data_mem_out_wire[855]), .IN1(n9761), .SEL(n10275), .F(
        n6921) );
  MUX U11129 ( .IN0(data_mem_out_wire[854]), .IN1(n9763), .SEL(n10275), .F(
        n6920) );
  MUX U11130 ( .IN0(data_mem_out_wire[853]), .IN1(n9764), .SEL(n10275), .F(
        n6919) );
  MUX U11131 ( .IN0(data_mem_out_wire[852]), .IN1(n9765), .SEL(n10275), .F(
        n6918) );
  MUX U11132 ( .IN0(data_mem_out_wire[851]), .IN1(n9766), .SEL(n10275), .F(
        n6917) );
  IV U11133 ( .A(n10276), .Z(n10275) );
  MUX U11134 ( .IN0(n9768), .IN1(data_mem_out_wire[850]), .SEL(n10276), .F(
        n6916) );
  MUX U11135 ( .IN0(n9769), .IN1(data_mem_out_wire[849]), .SEL(n10276), .F(
        n6915) );
  MUX U11136 ( .IN0(n9770), .IN1(data_mem_out_wire[848]), .SEL(n10276), .F(
        n6914) );
  AND U11137 ( .A(n10277), .B(n10278), .Z(n10276) );
  OR U11138 ( .A(n9773), .B(n10274), .Z(n10278) );
  AND U11139 ( .A(n10272), .B(n10271), .Z(n10277) );
  NANDN U11140 ( .A(n10274), .B(n9809), .Z(n10272) );
  MUX U11141 ( .IN0(data_mem_out_wire[847]), .IN1(n9776), .SEL(n10279), .F(
        n6913) );
  MUX U11142 ( .IN0(data_mem_out_wire[846]), .IN1(n9778), .SEL(n10279), .F(
        n6912) );
  MUX U11143 ( .IN0(data_mem_out_wire[845]), .IN1(n9779), .SEL(n10279), .F(
        n6911) );
  MUX U11144 ( .IN0(data_mem_out_wire[844]), .IN1(n9780), .SEL(n10279), .F(
        n6910) );
  MUX U11145 ( .IN0(data_mem_out_wire[843]), .IN1(n9781), .SEL(n10279), .F(
        n6909) );
  IV U11146 ( .A(n10280), .Z(n10279) );
  MUX U11147 ( .IN0(n9783), .IN1(data_mem_out_wire[842]), .SEL(n10280), .F(
        n6908) );
  MUX U11148 ( .IN0(n9784), .IN1(data_mem_out_wire[841]), .SEL(n10280), .F(
        n6907) );
  MUX U11149 ( .IN0(n9785), .IN1(data_mem_out_wire[840]), .SEL(n10280), .F(
        n6906) );
  AND U11150 ( .A(n10281), .B(n10282), .Z(n10280) );
  OR U11151 ( .A(n9788), .B(n10274), .Z(n10282) );
  MUX U11152 ( .IN0(data_mem_out_wire[839]), .IN1(data_in[7]), .SEL(n10283), 
        .F(n6905) );
  MUX U11153 ( .IN0(data_mem_out_wire[838]), .IN1(data_in[6]), .SEL(n10283), 
        .F(n6904) );
  MUX U11154 ( .IN0(data_mem_out_wire[837]), .IN1(data_in[5]), .SEL(n10283), 
        .F(n6903) );
  MUX U11155 ( .IN0(data_mem_out_wire[836]), .IN1(data_in[4]), .SEL(n10283), 
        .F(n6902) );
  MUX U11156 ( .IN0(data_mem_out_wire[835]), .IN1(data_in[3]), .SEL(n10283), 
        .F(n6901) );
  IV U11157 ( .A(n10284), .Z(n10283) );
  MUX U11158 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[834]), .SEL(n10284), 
        .F(n6900) );
  MUX U11159 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[833]), .SEL(n10284), 
        .F(n6899) );
  MUX U11160 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[832]), .SEL(n10284), 
        .F(n6898) );
  AND U11161 ( .A(n10281), .B(n10285), .Z(n10284) );
  NANDN U11162 ( .A(n10274), .B(n9792), .Z(n10285) );
  AND U11163 ( .A(n10286), .B(n10271), .Z(n10281) );
  NANDN U11164 ( .A(n10274), .B(n9796), .Z(n10271) );
  NANDN U11165 ( .A(n10274), .B(n9818), .Z(n10286) );
  NAND U11166 ( .A(n9838), .B(n10250), .Z(n10274) );
  MUX U11167 ( .IN0(n9746), .IN1(data_mem_out_wire[895]), .SEL(n10287), .F(
        n6897) );
  MUX U11168 ( .IN0(n9748), .IN1(data_mem_out_wire[894]), .SEL(n10287), .F(
        n6896) );
  MUX U11169 ( .IN0(n9749), .IN1(data_mem_out_wire[893]), .SEL(n10287), .F(
        n6895) );
  MUX U11170 ( .IN0(n9750), .IN1(data_mem_out_wire[892]), .SEL(n10287), .F(
        n6894) );
  MUX U11171 ( .IN0(n9751), .IN1(data_mem_out_wire[891]), .SEL(n10287), .F(
        n6893) );
  MUX U11172 ( .IN0(n9752), .IN1(data_mem_out_wire[890]), .SEL(n10287), .F(
        n6892) );
  MUX U11173 ( .IN0(n9753), .IN1(data_mem_out_wire[889]), .SEL(n10287), .F(
        n6891) );
  MUX U11174 ( .IN0(n9754), .IN1(data_mem_out_wire[888]), .SEL(n10287), .F(
        n6890) );
  AND U11175 ( .A(n10288), .B(n10289), .Z(n10287) );
  AND U11176 ( .A(n10290), .B(n10291), .Z(n10288) );
  OR U11177 ( .A(n9760), .B(n10292), .Z(n10291) );
  MUX U11178 ( .IN0(data_mem_out_wire[887]), .IN1(n9761), .SEL(n10293), .F(
        n6889) );
  MUX U11179 ( .IN0(data_mem_out_wire[886]), .IN1(n9763), .SEL(n10293), .F(
        n6888) );
  MUX U11180 ( .IN0(data_mem_out_wire[885]), .IN1(n9764), .SEL(n10293), .F(
        n6887) );
  MUX U11181 ( .IN0(data_mem_out_wire[884]), .IN1(n9765), .SEL(n10293), .F(
        n6886) );
  MUX U11182 ( .IN0(data_mem_out_wire[883]), .IN1(n9766), .SEL(n10293), .F(
        n6885) );
  IV U11183 ( .A(n10294), .Z(n10293) );
  MUX U11184 ( .IN0(n9768), .IN1(data_mem_out_wire[882]), .SEL(n10294), .F(
        n6884) );
  MUX U11185 ( .IN0(n9769), .IN1(data_mem_out_wire[881]), .SEL(n10294), .F(
        n6883) );
  MUX U11186 ( .IN0(n9770), .IN1(data_mem_out_wire[880]), .SEL(n10294), .F(
        n6882) );
  AND U11187 ( .A(n10295), .B(n10296), .Z(n10294) );
  OR U11188 ( .A(n9773), .B(n10292), .Z(n10296) );
  AND U11189 ( .A(n10290), .B(n10289), .Z(n10295) );
  NANDN U11190 ( .A(n10292), .B(n9809), .Z(n10290) );
  MUX U11191 ( .IN0(data_mem_out_wire[879]), .IN1(n9776), .SEL(n10297), .F(
        n6881) );
  MUX U11192 ( .IN0(data_mem_out_wire[878]), .IN1(n9778), .SEL(n10297), .F(
        n6880) );
  MUX U11193 ( .IN0(data_mem_out_wire[877]), .IN1(n9779), .SEL(n10297), .F(
        n6879) );
  MUX U11194 ( .IN0(data_mem_out_wire[876]), .IN1(n9780), .SEL(n10297), .F(
        n6878) );
  MUX U11195 ( .IN0(data_mem_out_wire[875]), .IN1(n9781), .SEL(n10297), .F(
        n6877) );
  IV U11196 ( .A(n10298), .Z(n10297) );
  MUX U11197 ( .IN0(n9783), .IN1(data_mem_out_wire[874]), .SEL(n10298), .F(
        n6876) );
  MUX U11198 ( .IN0(n9784), .IN1(data_mem_out_wire[873]), .SEL(n10298), .F(
        n6875) );
  MUX U11199 ( .IN0(n9785), .IN1(data_mem_out_wire[872]), .SEL(n10298), .F(
        n6874) );
  AND U11200 ( .A(n10299), .B(n10300), .Z(n10298) );
  OR U11201 ( .A(n9788), .B(n10292), .Z(n10300) );
  MUX U11202 ( .IN0(data_mem_out_wire[871]), .IN1(data_in[7]), .SEL(n10301), 
        .F(n6873) );
  MUX U11203 ( .IN0(data_mem_out_wire[870]), .IN1(data_in[6]), .SEL(n10301), 
        .F(n6872) );
  MUX U11204 ( .IN0(data_mem_out_wire[869]), .IN1(data_in[5]), .SEL(n10301), 
        .F(n6871) );
  MUX U11205 ( .IN0(data_mem_out_wire[868]), .IN1(data_in[4]), .SEL(n10301), 
        .F(n6870) );
  MUX U11206 ( .IN0(data_mem_out_wire[867]), .IN1(data_in[3]), .SEL(n10301), 
        .F(n6869) );
  IV U11207 ( .A(n10302), .Z(n10301) );
  MUX U11208 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[866]), .SEL(n10302), 
        .F(n6868) );
  MUX U11209 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[865]), .SEL(n10302), 
        .F(n6867) );
  MUX U11210 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[864]), .SEL(n10302), 
        .F(n6866) );
  AND U11211 ( .A(n10299), .B(n10303), .Z(n10302) );
  NANDN U11212 ( .A(n10292), .B(n9792), .Z(n10303) );
  AND U11213 ( .A(n10304), .B(n10289), .Z(n10299) );
  NANDN U11214 ( .A(n10292), .B(n9796), .Z(n10289) );
  NANDN U11215 ( .A(n10292), .B(n9818), .Z(n10304) );
  NAND U11216 ( .A(n9862), .B(n10250), .Z(n10292) );
  MUX U11217 ( .IN0(n9746), .IN1(data_mem_out_wire[927]), .SEL(n10305), .F(
        n6865) );
  MUX U11218 ( .IN0(n9748), .IN1(data_mem_out_wire[926]), .SEL(n10305), .F(
        n6864) );
  MUX U11219 ( .IN0(n9749), .IN1(data_mem_out_wire[925]), .SEL(n10305), .F(
        n6863) );
  MUX U11220 ( .IN0(n9750), .IN1(data_mem_out_wire[924]), .SEL(n10305), .F(
        n6862) );
  MUX U11221 ( .IN0(n9751), .IN1(data_mem_out_wire[923]), .SEL(n10305), .F(
        n6861) );
  MUX U11222 ( .IN0(n9752), .IN1(data_mem_out_wire[922]), .SEL(n10305), .F(
        n6860) );
  MUX U11223 ( .IN0(n9753), .IN1(data_mem_out_wire[921]), .SEL(n10305), .F(
        n6859) );
  MUX U11224 ( .IN0(n9754), .IN1(data_mem_out_wire[920]), .SEL(n10305), .F(
        n6858) );
  AND U11225 ( .A(n10306), .B(n10307), .Z(n10305) );
  AND U11226 ( .A(n10308), .B(n10309), .Z(n10306) );
  OR U11227 ( .A(n9760), .B(n10310), .Z(n10309) );
  MUX U11228 ( .IN0(data_mem_out_wire[919]), .IN1(n9761), .SEL(n10311), .F(
        n6857) );
  MUX U11229 ( .IN0(data_mem_out_wire[918]), .IN1(n9763), .SEL(n10311), .F(
        n6856) );
  MUX U11230 ( .IN0(data_mem_out_wire[917]), .IN1(n9764), .SEL(n10311), .F(
        n6855) );
  MUX U11231 ( .IN0(data_mem_out_wire[916]), .IN1(n9765), .SEL(n10311), .F(
        n6854) );
  MUX U11232 ( .IN0(data_mem_out_wire[915]), .IN1(n9766), .SEL(n10311), .F(
        n6853) );
  IV U11233 ( .A(n10312), .Z(n10311) );
  MUX U11234 ( .IN0(n9768), .IN1(data_mem_out_wire[914]), .SEL(n10312), .F(
        n6852) );
  MUX U11235 ( .IN0(n9769), .IN1(data_mem_out_wire[913]), .SEL(n10312), .F(
        n6851) );
  MUX U11236 ( .IN0(n9770), .IN1(data_mem_out_wire[912]), .SEL(n10312), .F(
        n6850) );
  AND U11237 ( .A(n10313), .B(n10314), .Z(n10312) );
  OR U11238 ( .A(n9773), .B(n10310), .Z(n10314) );
  AND U11239 ( .A(n10308), .B(n10307), .Z(n10313) );
  NANDN U11240 ( .A(n10310), .B(n9809), .Z(n10308) );
  MUX U11241 ( .IN0(data_mem_out_wire[911]), .IN1(n9776), .SEL(n10315), .F(
        n6849) );
  MUX U11242 ( .IN0(data_mem_out_wire[910]), .IN1(n9778), .SEL(n10315), .F(
        n6848) );
  MUX U11243 ( .IN0(data_mem_out_wire[909]), .IN1(n9779), .SEL(n10315), .F(
        n6847) );
  MUX U11244 ( .IN0(data_mem_out_wire[908]), .IN1(n9780), .SEL(n10315), .F(
        n6846) );
  MUX U11245 ( .IN0(data_mem_out_wire[907]), .IN1(n9781), .SEL(n10315), .F(
        n6845) );
  IV U11246 ( .A(n10316), .Z(n10315) );
  MUX U11247 ( .IN0(n9783), .IN1(data_mem_out_wire[906]), .SEL(n10316), .F(
        n6844) );
  MUX U11248 ( .IN0(n9784), .IN1(data_mem_out_wire[905]), .SEL(n10316), .F(
        n6843) );
  MUX U11249 ( .IN0(n9785), .IN1(data_mem_out_wire[904]), .SEL(n10316), .F(
        n6842) );
  AND U11250 ( .A(n10317), .B(n10318), .Z(n10316) );
  OR U11251 ( .A(n9788), .B(n10310), .Z(n10318) );
  MUX U11252 ( .IN0(data_mem_out_wire[903]), .IN1(data_in[7]), .SEL(n10319), 
        .F(n6841) );
  MUX U11253 ( .IN0(data_mem_out_wire[902]), .IN1(data_in[6]), .SEL(n10319), 
        .F(n6840) );
  MUX U11254 ( .IN0(data_mem_out_wire[901]), .IN1(data_in[5]), .SEL(n10319), 
        .F(n6839) );
  MUX U11255 ( .IN0(data_mem_out_wire[900]), .IN1(data_in[4]), .SEL(n10319), 
        .F(n6838) );
  MUX U11256 ( .IN0(data_mem_out_wire[899]), .IN1(data_in[3]), .SEL(n10319), 
        .F(n6837) );
  IV U11257 ( .A(n10320), .Z(n10319) );
  MUX U11258 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[898]), .SEL(n10320), 
        .F(n6836) );
  MUX U11259 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[897]), .SEL(n10320), 
        .F(n6835) );
  MUX U11260 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[896]), .SEL(n10320), 
        .F(n6834) );
  AND U11261 ( .A(n10317), .B(n10321), .Z(n10320) );
  NANDN U11262 ( .A(n10310), .B(n9792), .Z(n10321) );
  AND U11263 ( .A(n10322), .B(n10307), .Z(n10317) );
  NANDN U11264 ( .A(n10310), .B(n9796), .Z(n10307) );
  NANDN U11265 ( .A(n10310), .B(n9818), .Z(n10322) );
  NAND U11266 ( .A(n9881), .B(n10250), .Z(n10310) );
  MUX U11267 ( .IN0(n9746), .IN1(data_mem_out_wire[959]), .SEL(n10323), .F(
        n6833) );
  MUX U11268 ( .IN0(n9748), .IN1(data_mem_out_wire[958]), .SEL(n10323), .F(
        n6832) );
  MUX U11269 ( .IN0(n9749), .IN1(data_mem_out_wire[957]), .SEL(n10323), .F(
        n6831) );
  MUX U11270 ( .IN0(n9750), .IN1(data_mem_out_wire[956]), .SEL(n10323), .F(
        n6830) );
  MUX U11271 ( .IN0(n9751), .IN1(data_mem_out_wire[955]), .SEL(n10323), .F(
        n6829) );
  MUX U11272 ( .IN0(n9752), .IN1(data_mem_out_wire[954]), .SEL(n10323), .F(
        n6828) );
  MUX U11273 ( .IN0(n9753), .IN1(data_mem_out_wire[953]), .SEL(n10323), .F(
        n6827) );
  MUX U11274 ( .IN0(n9754), .IN1(data_mem_out_wire[952]), .SEL(n10323), .F(
        n6826) );
  AND U11275 ( .A(n10324), .B(n10325), .Z(n10323) );
  AND U11276 ( .A(n10326), .B(n10327), .Z(n10324) );
  OR U11277 ( .A(n9760), .B(n10328), .Z(n10327) );
  MUX U11278 ( .IN0(data_mem_out_wire[951]), .IN1(n9761), .SEL(n10329), .F(
        n6825) );
  MUX U11279 ( .IN0(data_mem_out_wire[950]), .IN1(n9763), .SEL(n10329), .F(
        n6824) );
  MUX U11280 ( .IN0(data_mem_out_wire[949]), .IN1(n9764), .SEL(n10329), .F(
        n6823) );
  MUX U11281 ( .IN0(data_mem_out_wire[948]), .IN1(n9765), .SEL(n10329), .F(
        n6822) );
  MUX U11282 ( .IN0(data_mem_out_wire[947]), .IN1(n9766), .SEL(n10329), .F(
        n6821) );
  IV U11283 ( .A(n10330), .Z(n10329) );
  MUX U11284 ( .IN0(n9768), .IN1(data_mem_out_wire[946]), .SEL(n10330), .F(
        n6820) );
  MUX U11285 ( .IN0(n9769), .IN1(data_mem_out_wire[945]), .SEL(n10330), .F(
        n6819) );
  MUX U11286 ( .IN0(n9770), .IN1(data_mem_out_wire[944]), .SEL(n10330), .F(
        n6818) );
  AND U11287 ( .A(n10331), .B(n10332), .Z(n10330) );
  OR U11288 ( .A(n9773), .B(n10328), .Z(n10332) );
  AND U11289 ( .A(n10326), .B(n10325), .Z(n10331) );
  NANDN U11290 ( .A(n10328), .B(n9809), .Z(n10326) );
  MUX U11291 ( .IN0(data_mem_out_wire[943]), .IN1(n9776), .SEL(n10333), .F(
        n6817) );
  MUX U11292 ( .IN0(data_mem_out_wire[942]), .IN1(n9778), .SEL(n10333), .F(
        n6816) );
  MUX U11293 ( .IN0(data_mem_out_wire[941]), .IN1(n9779), .SEL(n10333), .F(
        n6815) );
  MUX U11294 ( .IN0(data_mem_out_wire[940]), .IN1(n9780), .SEL(n10333), .F(
        n6814) );
  MUX U11295 ( .IN0(data_mem_out_wire[939]), .IN1(n9781), .SEL(n10333), .F(
        n6813) );
  IV U11296 ( .A(n10334), .Z(n10333) );
  MUX U11297 ( .IN0(n9783), .IN1(data_mem_out_wire[938]), .SEL(n10334), .F(
        n6812) );
  MUX U11298 ( .IN0(n9784), .IN1(data_mem_out_wire[937]), .SEL(n10334), .F(
        n6811) );
  MUX U11299 ( .IN0(n9785), .IN1(data_mem_out_wire[936]), .SEL(n10334), .F(
        n6810) );
  AND U11300 ( .A(n10335), .B(n10336), .Z(n10334) );
  OR U11301 ( .A(n9788), .B(n10328), .Z(n10336) );
  MUX U11302 ( .IN0(data_mem_out_wire[935]), .IN1(data_in[7]), .SEL(n10337), 
        .F(n6809) );
  MUX U11303 ( .IN0(data_mem_out_wire[934]), .IN1(data_in[6]), .SEL(n10337), 
        .F(n6808) );
  MUX U11304 ( .IN0(data_mem_out_wire[933]), .IN1(data_in[5]), .SEL(n10337), 
        .F(n6807) );
  MUX U11305 ( .IN0(data_mem_out_wire[932]), .IN1(data_in[4]), .SEL(n10337), 
        .F(n6806) );
  MUX U11306 ( .IN0(data_mem_out_wire[931]), .IN1(data_in[3]), .SEL(n10337), 
        .F(n6805) );
  IV U11307 ( .A(n10338), .Z(n10337) );
  MUX U11308 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[930]), .SEL(n10338), 
        .F(n6804) );
  MUX U11309 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[929]), .SEL(n10338), 
        .F(n6803) );
  MUX U11310 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[928]), .SEL(n10338), 
        .F(n6802) );
  AND U11311 ( .A(n10335), .B(n10339), .Z(n10338) );
  NANDN U11312 ( .A(n10328), .B(n9792), .Z(n10339) );
  AND U11313 ( .A(n10340), .B(n10325), .Z(n10335) );
  NANDN U11314 ( .A(n10328), .B(n9796), .Z(n10325) );
  NANDN U11315 ( .A(n10328), .B(n9818), .Z(n10340) );
  NAND U11316 ( .A(n9900), .B(n10250), .Z(n10328) );
  MUX U11317 ( .IN0(n9746), .IN1(data_mem_out_wire[991]), .SEL(n10341), .F(
        n6801) );
  MUX U11318 ( .IN0(n9748), .IN1(data_mem_out_wire[990]), .SEL(n10341), .F(
        n6800) );
  MUX U11319 ( .IN0(n9749), .IN1(data_mem_out_wire[989]), .SEL(n10341), .F(
        n6799) );
  MUX U11320 ( .IN0(n9750), .IN1(data_mem_out_wire[988]), .SEL(n10341), .F(
        n6798) );
  MUX U11321 ( .IN0(n9751), .IN1(data_mem_out_wire[987]), .SEL(n10341), .F(
        n6797) );
  MUX U11322 ( .IN0(n9752), .IN1(data_mem_out_wire[986]), .SEL(n10341), .F(
        n6796) );
  MUX U11323 ( .IN0(n9753), .IN1(data_mem_out_wire[985]), .SEL(n10341), .F(
        n6795) );
  MUX U11324 ( .IN0(n9754), .IN1(data_mem_out_wire[984]), .SEL(n10341), .F(
        n6794) );
  AND U11325 ( .A(n10342), .B(n10343), .Z(n10341) );
  AND U11326 ( .A(n10344), .B(n10345), .Z(n10342) );
  OR U11327 ( .A(n9760), .B(n10346), .Z(n10345) );
  MUX U11328 ( .IN0(data_mem_out_wire[983]), .IN1(n9761), .SEL(n10347), .F(
        n6793) );
  MUX U11329 ( .IN0(data_mem_out_wire[982]), .IN1(n9763), .SEL(n10347), .F(
        n6792) );
  MUX U11330 ( .IN0(data_mem_out_wire[981]), .IN1(n9764), .SEL(n10347), .F(
        n6791) );
  MUX U11331 ( .IN0(data_mem_out_wire[980]), .IN1(n9765), .SEL(n10347), .F(
        n6790) );
  MUX U11332 ( .IN0(data_mem_out_wire[979]), .IN1(n9766), .SEL(n10347), .F(
        n6789) );
  IV U11333 ( .A(n10348), .Z(n10347) );
  MUX U11334 ( .IN0(n9768), .IN1(data_mem_out_wire[978]), .SEL(n10348), .F(
        n6788) );
  MUX U11335 ( .IN0(n9769), .IN1(data_mem_out_wire[977]), .SEL(n10348), .F(
        n6787) );
  MUX U11336 ( .IN0(n9770), .IN1(data_mem_out_wire[976]), .SEL(n10348), .F(
        n6786) );
  AND U11337 ( .A(n10349), .B(n10350), .Z(n10348) );
  OR U11338 ( .A(n9773), .B(n10346), .Z(n10350) );
  AND U11339 ( .A(n10344), .B(n10343), .Z(n10349) );
  NANDN U11340 ( .A(n10346), .B(n9809), .Z(n10344) );
  MUX U11341 ( .IN0(data_mem_out_wire[975]), .IN1(n9776), .SEL(n10351), .F(
        n6785) );
  MUX U11342 ( .IN0(data_mem_out_wire[974]), .IN1(n9778), .SEL(n10351), .F(
        n6784) );
  MUX U11343 ( .IN0(data_mem_out_wire[973]), .IN1(n9779), .SEL(n10351), .F(
        n6783) );
  MUX U11344 ( .IN0(data_mem_out_wire[972]), .IN1(n9780), .SEL(n10351), .F(
        n6782) );
  MUX U11345 ( .IN0(data_mem_out_wire[971]), .IN1(n9781), .SEL(n10351), .F(
        n6781) );
  IV U11346 ( .A(n10352), .Z(n10351) );
  MUX U11347 ( .IN0(n9783), .IN1(data_mem_out_wire[970]), .SEL(n10352), .F(
        n6780) );
  MUX U11348 ( .IN0(n9784), .IN1(data_mem_out_wire[969]), .SEL(n10352), .F(
        n6779) );
  MUX U11349 ( .IN0(n9785), .IN1(data_mem_out_wire[968]), .SEL(n10352), .F(
        n6778) );
  AND U11350 ( .A(n10353), .B(n10354), .Z(n10352) );
  OR U11351 ( .A(n9788), .B(n10346), .Z(n10354) );
  MUX U11352 ( .IN0(data_mem_out_wire[967]), .IN1(data_in[7]), .SEL(n10355), 
        .F(n6777) );
  MUX U11353 ( .IN0(data_mem_out_wire[966]), .IN1(data_in[6]), .SEL(n10355), 
        .F(n6776) );
  MUX U11354 ( .IN0(data_mem_out_wire[965]), .IN1(data_in[5]), .SEL(n10355), 
        .F(n6775) );
  MUX U11355 ( .IN0(data_mem_out_wire[964]), .IN1(data_in[4]), .SEL(n10355), 
        .F(n6774) );
  MUX U11356 ( .IN0(data_mem_out_wire[963]), .IN1(data_in[3]), .SEL(n10355), 
        .F(n6773) );
  IV U11357 ( .A(n10356), .Z(n10355) );
  MUX U11358 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[962]), .SEL(n10356), 
        .F(n6772) );
  MUX U11359 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[961]), .SEL(n10356), 
        .F(n6771) );
  MUX U11360 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[960]), .SEL(n10356), 
        .F(n6770) );
  AND U11361 ( .A(n10353), .B(n10357), .Z(n10356) );
  NANDN U11362 ( .A(n10346), .B(n9792), .Z(n10357) );
  AND U11363 ( .A(n10358), .B(n10343), .Z(n10353) );
  NANDN U11364 ( .A(n10346), .B(n9796), .Z(n10343) );
  NANDN U11365 ( .A(n10346), .B(n9818), .Z(n10358) );
  NAND U11366 ( .A(n9919), .B(n10250), .Z(n10346) );
  MUX U11367 ( .IN0(n9746), .IN1(data_mem_out_wire[1023]), .SEL(n10359), .F(
        n6769) );
  MUX U11368 ( .IN0(n9748), .IN1(data_mem_out_wire[1022]), .SEL(n10359), .F(
        n6768) );
  MUX U11369 ( .IN0(n9749), .IN1(data_mem_out_wire[1021]), .SEL(n10359), .F(
        n6767) );
  MUX U11370 ( .IN0(n9750), .IN1(data_mem_out_wire[1020]), .SEL(n10359), .F(
        n6766) );
  MUX U11371 ( .IN0(n9751), .IN1(data_mem_out_wire[1019]), .SEL(n10359), .F(
        n6765) );
  MUX U11372 ( .IN0(n9752), .IN1(data_mem_out_wire[1018]), .SEL(n10359), .F(
        n6764) );
  MUX U11373 ( .IN0(n9753), .IN1(data_mem_out_wire[1017]), .SEL(n10359), .F(
        n6763) );
  MUX U11374 ( .IN0(n9754), .IN1(data_mem_out_wire[1016]), .SEL(n10359), .F(
        n6762) );
  AND U11375 ( .A(n10360), .B(n10361), .Z(n10359) );
  AND U11376 ( .A(n10362), .B(n10363), .Z(n10360) );
  OR U11377 ( .A(n9760), .B(n10364), .Z(n10363) );
  MUX U11378 ( .IN0(data_mem_out_wire[1015]), .IN1(n9761), .SEL(n10365), .F(
        n6761) );
  MUX U11379 ( .IN0(data_mem_out_wire[1014]), .IN1(n9763), .SEL(n10365), .F(
        n6760) );
  MUX U11380 ( .IN0(data_mem_out_wire[1013]), .IN1(n9764), .SEL(n10365), .F(
        n6759) );
  MUX U11381 ( .IN0(data_mem_out_wire[1012]), .IN1(n9765), .SEL(n10365), .F(
        n6758) );
  MUX U11382 ( .IN0(data_mem_out_wire[1011]), .IN1(n9766), .SEL(n10365), .F(
        n6757) );
  IV U11383 ( .A(n10366), .Z(n10365) );
  MUX U11384 ( .IN0(n9768), .IN1(data_mem_out_wire[1010]), .SEL(n10366), .F(
        n6756) );
  MUX U11385 ( .IN0(n9769), .IN1(data_mem_out_wire[1009]), .SEL(n10366), .F(
        n6755) );
  MUX U11386 ( .IN0(n9770), .IN1(data_mem_out_wire[1008]), .SEL(n10366), .F(
        n6754) );
  AND U11387 ( .A(n10367), .B(n10368), .Z(n10366) );
  OR U11388 ( .A(n9773), .B(n10364), .Z(n10368) );
  AND U11389 ( .A(n10362), .B(n10361), .Z(n10367) );
  NANDN U11390 ( .A(n10364), .B(n9809), .Z(n10362) );
  MUX U11391 ( .IN0(data_mem_out_wire[1007]), .IN1(n9776), .SEL(n10369), .F(
        n6753) );
  MUX U11392 ( .IN0(data_mem_out_wire[1006]), .IN1(n9778), .SEL(n10369), .F(
        n6752) );
  MUX U11393 ( .IN0(data_mem_out_wire[1005]), .IN1(n9779), .SEL(n10369), .F(
        n6751) );
  MUX U11394 ( .IN0(data_mem_out_wire[1004]), .IN1(n9780), .SEL(n10369), .F(
        n6750) );
  MUX U11395 ( .IN0(data_mem_out_wire[1003]), .IN1(n9781), .SEL(n10369), .F(
        n6749) );
  IV U11396 ( .A(n10370), .Z(n10369) );
  MUX U11397 ( .IN0(n9783), .IN1(data_mem_out_wire[1002]), .SEL(n10370), .F(
        n6748) );
  MUX U11398 ( .IN0(n9784), .IN1(data_mem_out_wire[1001]), .SEL(n10370), .F(
        n6747) );
  MUX U11399 ( .IN0(n9785), .IN1(data_mem_out_wire[1000]), .SEL(n10370), .F(
        n6746) );
  AND U11400 ( .A(n10371), .B(n10372), .Z(n10370) );
  OR U11401 ( .A(n9788), .B(n10364), .Z(n10372) );
  MUX U11402 ( .IN0(data_mem_out_wire[999]), .IN1(data_in[7]), .SEL(n10373), 
        .F(n6745) );
  MUX U11403 ( .IN0(data_mem_out_wire[998]), .IN1(data_in[6]), .SEL(n10373), 
        .F(n6744) );
  MUX U11404 ( .IN0(data_mem_out_wire[997]), .IN1(data_in[5]), .SEL(n10373), 
        .F(n6743) );
  MUX U11405 ( .IN0(data_mem_out_wire[996]), .IN1(data_in[4]), .SEL(n10373), 
        .F(n6742) );
  MUX U11406 ( .IN0(data_mem_out_wire[995]), .IN1(data_in[3]), .SEL(n10373), 
        .F(n6741) );
  IV U11407 ( .A(n10374), .Z(n10373) );
  MUX U11408 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[994]), .SEL(n10374), 
        .F(n6740) );
  MUX U11409 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[993]), .SEL(n10374), 
        .F(n6739) );
  MUX U11410 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[992]), .SEL(n10374), 
        .F(n6738) );
  AND U11411 ( .A(n10371), .B(n10375), .Z(n10374) );
  NANDN U11412 ( .A(n10364), .B(n9792), .Z(n10375) );
  AND U11413 ( .A(n10376), .B(n10361), .Z(n10371) );
  NANDN U11414 ( .A(n10364), .B(n9796), .Z(n10361) );
  NANDN U11415 ( .A(n10364), .B(n9818), .Z(n10376) );
  NAND U11416 ( .A(n10250), .B(n9938), .Z(n10364) );
  ANDN U11417 ( .B(n10377), .A(N42), .Z(n10250) );
  MUX U11418 ( .IN0(n9746), .IN1(data_mem_out_wire[1055]), .SEL(n10378), .F(
        n6737) );
  MUX U11419 ( .IN0(n9748), .IN1(data_mem_out_wire[1054]), .SEL(n10378), .F(
        n6736) );
  MUX U11420 ( .IN0(n9749), .IN1(data_mem_out_wire[1053]), .SEL(n10378), .F(
        n6735) );
  MUX U11421 ( .IN0(n9750), .IN1(data_mem_out_wire[1052]), .SEL(n10378), .F(
        n6734) );
  MUX U11422 ( .IN0(n9751), .IN1(data_mem_out_wire[1051]), .SEL(n10378), .F(
        n6733) );
  MUX U11423 ( .IN0(n9752), .IN1(data_mem_out_wire[1050]), .SEL(n10378), .F(
        n6732) );
  MUX U11424 ( .IN0(n9753), .IN1(data_mem_out_wire[1049]), .SEL(n10378), .F(
        n6731) );
  MUX U11425 ( .IN0(n9754), .IN1(data_mem_out_wire[1048]), .SEL(n10378), .F(
        n6730) );
  AND U11426 ( .A(n10379), .B(n10380), .Z(n10378) );
  AND U11427 ( .A(n10381), .B(n10382), .Z(n10379) );
  OR U11428 ( .A(n9760), .B(n10383), .Z(n10382) );
  MUX U11429 ( .IN0(data_mem_out_wire[1047]), .IN1(n9761), .SEL(n10384), .F(
        n6729) );
  MUX U11430 ( .IN0(data_mem_out_wire[1046]), .IN1(n9763), .SEL(n10384), .F(
        n6728) );
  MUX U11431 ( .IN0(data_mem_out_wire[1045]), .IN1(n9764), .SEL(n10384), .F(
        n6727) );
  MUX U11432 ( .IN0(data_mem_out_wire[1044]), .IN1(n9765), .SEL(n10384), .F(
        n6726) );
  MUX U11433 ( .IN0(data_mem_out_wire[1043]), .IN1(n9766), .SEL(n10384), .F(
        n6725) );
  IV U11434 ( .A(n10385), .Z(n10384) );
  MUX U11435 ( .IN0(n9768), .IN1(data_mem_out_wire[1042]), .SEL(n10385), .F(
        n6724) );
  MUX U11436 ( .IN0(n9769), .IN1(data_mem_out_wire[1041]), .SEL(n10385), .F(
        n6723) );
  MUX U11437 ( .IN0(n9770), .IN1(data_mem_out_wire[1040]), .SEL(n10385), .F(
        n6722) );
  AND U11438 ( .A(n10386), .B(n10387), .Z(n10385) );
  OR U11439 ( .A(n9773), .B(n10383), .Z(n10387) );
  AND U11440 ( .A(n10381), .B(n10380), .Z(n10386) );
  NANDN U11441 ( .A(n10383), .B(n9809), .Z(n10381) );
  MUX U11442 ( .IN0(data_mem_out_wire[1039]), .IN1(n9776), .SEL(n10388), .F(
        n6721) );
  MUX U11443 ( .IN0(data_mem_out_wire[1038]), .IN1(n9778), .SEL(n10388), .F(
        n6720) );
  MUX U11444 ( .IN0(data_mem_out_wire[1037]), .IN1(n9779), .SEL(n10388), .F(
        n6719) );
  MUX U11445 ( .IN0(data_mem_out_wire[1036]), .IN1(n9780), .SEL(n10388), .F(
        n6718) );
  MUX U11446 ( .IN0(data_mem_out_wire[1035]), .IN1(n9781), .SEL(n10388), .F(
        n6717) );
  IV U11447 ( .A(n10389), .Z(n10388) );
  MUX U11448 ( .IN0(n9783), .IN1(data_mem_out_wire[1034]), .SEL(n10389), .F(
        n6716) );
  MUX U11449 ( .IN0(n9784), .IN1(data_mem_out_wire[1033]), .SEL(n10389), .F(
        n6715) );
  MUX U11450 ( .IN0(n9785), .IN1(data_mem_out_wire[1032]), .SEL(n10389), .F(
        n6714) );
  AND U11451 ( .A(n10390), .B(n10391), .Z(n10389) );
  OR U11452 ( .A(n9788), .B(n10383), .Z(n10391) );
  MUX U11453 ( .IN0(data_mem_out_wire[1031]), .IN1(data_in[7]), .SEL(n10392), 
        .F(n6713) );
  MUX U11454 ( .IN0(data_mem_out_wire[1030]), .IN1(data_in[6]), .SEL(n10392), 
        .F(n6712) );
  MUX U11455 ( .IN0(data_mem_out_wire[1029]), .IN1(data_in[5]), .SEL(n10392), 
        .F(n6711) );
  MUX U11456 ( .IN0(data_mem_out_wire[1028]), .IN1(data_in[4]), .SEL(n10392), 
        .F(n6710) );
  MUX U11457 ( .IN0(data_mem_out_wire[1027]), .IN1(data_in[3]), .SEL(n10392), 
        .F(n6709) );
  IV U11458 ( .A(n10393), .Z(n10392) );
  MUX U11459 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1026]), .SEL(n10393), 
        .F(n6708) );
  MUX U11460 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1025]), .SEL(n10393), 
        .F(n6707) );
  MUX U11461 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1024]), .SEL(n10393), 
        .F(n6706) );
  AND U11462 ( .A(n10390), .B(n10394), .Z(n10393) );
  NANDN U11463 ( .A(n10383), .B(n9792), .Z(n10394) );
  AND U11464 ( .A(n10395), .B(n10380), .Z(n10390) );
  NANDN U11465 ( .A(n10383), .B(n9796), .Z(n10380) );
  NANDN U11466 ( .A(n10383), .B(n9818), .Z(n10395) );
  NAND U11467 ( .A(n9798), .B(n10396), .Z(n10383) );
  MUX U11468 ( .IN0(n9746), .IN1(data_mem_out_wire[1087]), .SEL(n10397), .F(
        n6705) );
  MUX U11469 ( .IN0(n9748), .IN1(data_mem_out_wire[1086]), .SEL(n10397), .F(
        n6704) );
  MUX U11470 ( .IN0(n9749), .IN1(data_mem_out_wire[1085]), .SEL(n10397), .F(
        n6703) );
  MUX U11471 ( .IN0(n9750), .IN1(data_mem_out_wire[1084]), .SEL(n10397), .F(
        n6702) );
  MUX U11472 ( .IN0(n9751), .IN1(data_mem_out_wire[1083]), .SEL(n10397), .F(
        n6701) );
  MUX U11473 ( .IN0(n9752), .IN1(data_mem_out_wire[1082]), .SEL(n10397), .F(
        n6700) );
  MUX U11474 ( .IN0(n9753), .IN1(data_mem_out_wire[1081]), .SEL(n10397), .F(
        n6699) );
  MUX U11475 ( .IN0(n9754), .IN1(data_mem_out_wire[1080]), .SEL(n10397), .F(
        n6698) );
  AND U11476 ( .A(n10398), .B(n10399), .Z(n10397) );
  AND U11477 ( .A(n10400), .B(n10401), .Z(n10398) );
  OR U11478 ( .A(n9760), .B(n10402), .Z(n10401) );
  MUX U11479 ( .IN0(data_mem_out_wire[1079]), .IN1(n9761), .SEL(n10403), .F(
        n6697) );
  MUX U11480 ( .IN0(data_mem_out_wire[1078]), .IN1(n9763), .SEL(n10403), .F(
        n6696) );
  MUX U11481 ( .IN0(data_mem_out_wire[1077]), .IN1(n9764), .SEL(n10403), .F(
        n6695) );
  MUX U11482 ( .IN0(data_mem_out_wire[1076]), .IN1(n9765), .SEL(n10403), .F(
        n6694) );
  MUX U11483 ( .IN0(data_mem_out_wire[1075]), .IN1(n9766), .SEL(n10403), .F(
        n6693) );
  IV U11484 ( .A(n10404), .Z(n10403) );
  MUX U11485 ( .IN0(n9768), .IN1(data_mem_out_wire[1074]), .SEL(n10404), .F(
        n6692) );
  MUX U11486 ( .IN0(n9769), .IN1(data_mem_out_wire[1073]), .SEL(n10404), .F(
        n6691) );
  MUX U11487 ( .IN0(n9770), .IN1(data_mem_out_wire[1072]), .SEL(n10404), .F(
        n6690) );
  AND U11488 ( .A(n10405), .B(n10406), .Z(n10404) );
  OR U11489 ( .A(n9773), .B(n10402), .Z(n10406) );
  AND U11490 ( .A(n10400), .B(n10399), .Z(n10405) );
  NANDN U11491 ( .A(n10402), .B(n9809), .Z(n10400) );
  MUX U11492 ( .IN0(data_mem_out_wire[1071]), .IN1(n9776), .SEL(n10407), .F(
        n6689) );
  MUX U11493 ( .IN0(data_mem_out_wire[1070]), .IN1(n9778), .SEL(n10407), .F(
        n6688) );
  MUX U11494 ( .IN0(data_mem_out_wire[1069]), .IN1(n9779), .SEL(n10407), .F(
        n6687) );
  MUX U11495 ( .IN0(data_mem_out_wire[1068]), .IN1(n9780), .SEL(n10407), .F(
        n6686) );
  MUX U11496 ( .IN0(data_mem_out_wire[1067]), .IN1(n9781), .SEL(n10407), .F(
        n6685) );
  IV U11497 ( .A(n10408), .Z(n10407) );
  MUX U11498 ( .IN0(n9783), .IN1(data_mem_out_wire[1066]), .SEL(n10408), .F(
        n6684) );
  MUX U11499 ( .IN0(n9784), .IN1(data_mem_out_wire[1065]), .SEL(n10408), .F(
        n6683) );
  MUX U11500 ( .IN0(n9785), .IN1(data_mem_out_wire[1064]), .SEL(n10408), .F(
        n6682) );
  AND U11501 ( .A(n10409), .B(n10410), .Z(n10408) );
  OR U11502 ( .A(n9788), .B(n10402), .Z(n10410) );
  MUX U11503 ( .IN0(data_mem_out_wire[1063]), .IN1(data_in[7]), .SEL(n10411), 
        .F(n6681) );
  MUX U11504 ( .IN0(data_mem_out_wire[1062]), .IN1(data_in[6]), .SEL(n10411), 
        .F(n6680) );
  MUX U11505 ( .IN0(data_mem_out_wire[1061]), .IN1(data_in[5]), .SEL(n10411), 
        .F(n6679) );
  MUX U11506 ( .IN0(data_mem_out_wire[1060]), .IN1(data_in[4]), .SEL(n10411), 
        .F(n6678) );
  MUX U11507 ( .IN0(data_mem_out_wire[1059]), .IN1(data_in[3]), .SEL(n10411), 
        .F(n6677) );
  IV U11508 ( .A(n10412), .Z(n10411) );
  MUX U11509 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1058]), .SEL(n10412), 
        .F(n6676) );
  MUX U11510 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1057]), .SEL(n10412), 
        .F(n6675) );
  MUX U11511 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1056]), .SEL(n10412), 
        .F(n6674) );
  AND U11512 ( .A(n10409), .B(n10413), .Z(n10412) );
  NANDN U11513 ( .A(n10402), .B(n9792), .Z(n10413) );
  AND U11514 ( .A(n10414), .B(n10399), .Z(n10409) );
  NANDN U11515 ( .A(n10402), .B(n9796), .Z(n10399) );
  NANDN U11516 ( .A(n10402), .B(n9818), .Z(n10414) );
  NAND U11517 ( .A(n9819), .B(n10396), .Z(n10402) );
  MUX U11518 ( .IN0(n9746), .IN1(data_mem_out_wire[1119]), .SEL(n10415), .F(
        n6673) );
  MUX U11519 ( .IN0(n9748), .IN1(data_mem_out_wire[1118]), .SEL(n10415), .F(
        n6672) );
  MUX U11520 ( .IN0(n9749), .IN1(data_mem_out_wire[1117]), .SEL(n10415), .F(
        n6671) );
  MUX U11521 ( .IN0(n9750), .IN1(data_mem_out_wire[1116]), .SEL(n10415), .F(
        n6670) );
  MUX U11522 ( .IN0(n9751), .IN1(data_mem_out_wire[1115]), .SEL(n10415), .F(
        n6669) );
  MUX U11523 ( .IN0(n9752), .IN1(data_mem_out_wire[1114]), .SEL(n10415), .F(
        n6668) );
  MUX U11524 ( .IN0(n9753), .IN1(data_mem_out_wire[1113]), .SEL(n10415), .F(
        n6667) );
  MUX U11525 ( .IN0(n9754), .IN1(data_mem_out_wire[1112]), .SEL(n10415), .F(
        n6666) );
  AND U11526 ( .A(n10416), .B(n10417), .Z(n10415) );
  AND U11527 ( .A(n10418), .B(n10419), .Z(n10416) );
  OR U11528 ( .A(n9760), .B(n10420), .Z(n10419) );
  MUX U11529 ( .IN0(data_mem_out_wire[1111]), .IN1(n9761), .SEL(n10421), .F(
        n6665) );
  MUX U11530 ( .IN0(data_mem_out_wire[1110]), .IN1(n9763), .SEL(n10421), .F(
        n6664) );
  MUX U11531 ( .IN0(data_mem_out_wire[1109]), .IN1(n9764), .SEL(n10421), .F(
        n6663) );
  MUX U11532 ( .IN0(data_mem_out_wire[1108]), .IN1(n9765), .SEL(n10421), .F(
        n6662) );
  MUX U11533 ( .IN0(data_mem_out_wire[1107]), .IN1(n9766), .SEL(n10421), .F(
        n6661) );
  IV U11534 ( .A(n10422), .Z(n10421) );
  MUX U11535 ( .IN0(n9768), .IN1(data_mem_out_wire[1106]), .SEL(n10422), .F(
        n6660) );
  MUX U11536 ( .IN0(n9769), .IN1(data_mem_out_wire[1105]), .SEL(n10422), .F(
        n6659) );
  MUX U11537 ( .IN0(n9770), .IN1(data_mem_out_wire[1104]), .SEL(n10422), .F(
        n6658) );
  AND U11538 ( .A(n10423), .B(n10424), .Z(n10422) );
  OR U11539 ( .A(n9773), .B(n10420), .Z(n10424) );
  AND U11540 ( .A(n10418), .B(n10417), .Z(n10423) );
  NANDN U11541 ( .A(n10420), .B(n9809), .Z(n10418) );
  MUX U11542 ( .IN0(data_mem_out_wire[1103]), .IN1(n9776), .SEL(n10425), .F(
        n6657) );
  MUX U11543 ( .IN0(data_mem_out_wire[1102]), .IN1(n9778), .SEL(n10425), .F(
        n6656) );
  MUX U11544 ( .IN0(data_mem_out_wire[1101]), .IN1(n9779), .SEL(n10425), .F(
        n6655) );
  MUX U11545 ( .IN0(data_mem_out_wire[1100]), .IN1(n9780), .SEL(n10425), .F(
        n6654) );
  MUX U11546 ( .IN0(data_mem_out_wire[1099]), .IN1(n9781), .SEL(n10425), .F(
        n6653) );
  IV U11547 ( .A(n10426), .Z(n10425) );
  MUX U11548 ( .IN0(n9783), .IN1(data_mem_out_wire[1098]), .SEL(n10426), .F(
        n6652) );
  MUX U11549 ( .IN0(n9784), .IN1(data_mem_out_wire[1097]), .SEL(n10426), .F(
        n6651) );
  MUX U11550 ( .IN0(n9785), .IN1(data_mem_out_wire[1096]), .SEL(n10426), .F(
        n6650) );
  AND U11551 ( .A(n10427), .B(n10428), .Z(n10426) );
  OR U11552 ( .A(n9788), .B(n10420), .Z(n10428) );
  MUX U11553 ( .IN0(data_mem_out_wire[1095]), .IN1(data_in[7]), .SEL(n10429), 
        .F(n6649) );
  MUX U11554 ( .IN0(data_mem_out_wire[1094]), .IN1(data_in[6]), .SEL(n10429), 
        .F(n6648) );
  MUX U11555 ( .IN0(data_mem_out_wire[1093]), .IN1(data_in[5]), .SEL(n10429), 
        .F(n6647) );
  MUX U11556 ( .IN0(data_mem_out_wire[1092]), .IN1(data_in[4]), .SEL(n10429), 
        .F(n6646) );
  MUX U11557 ( .IN0(data_mem_out_wire[1091]), .IN1(data_in[3]), .SEL(n10429), 
        .F(n6645) );
  IV U11558 ( .A(n10430), .Z(n10429) );
  MUX U11559 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1090]), .SEL(n10430), 
        .F(n6644) );
  MUX U11560 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1089]), .SEL(n10430), 
        .F(n6643) );
  MUX U11561 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1088]), .SEL(n10430), 
        .F(n6642) );
  AND U11562 ( .A(n10427), .B(n10431), .Z(n10430) );
  NANDN U11563 ( .A(n10420), .B(n9792), .Z(n10431) );
  AND U11564 ( .A(n10432), .B(n10417), .Z(n10427) );
  NANDN U11565 ( .A(n10420), .B(n9796), .Z(n10417) );
  NANDN U11566 ( .A(n10420), .B(n9818), .Z(n10432) );
  NAND U11567 ( .A(n9838), .B(n10396), .Z(n10420) );
  MUX U11568 ( .IN0(n9746), .IN1(data_mem_out_wire[1151]), .SEL(n10433), .F(
        n6641) );
  MUX U11569 ( .IN0(n9748), .IN1(data_mem_out_wire[1150]), .SEL(n10433), .F(
        n6640) );
  MUX U11570 ( .IN0(n9749), .IN1(data_mem_out_wire[1149]), .SEL(n10433), .F(
        n6639) );
  MUX U11571 ( .IN0(n9750), .IN1(data_mem_out_wire[1148]), .SEL(n10433), .F(
        n6638) );
  MUX U11572 ( .IN0(n9751), .IN1(data_mem_out_wire[1147]), .SEL(n10433), .F(
        n6637) );
  MUX U11573 ( .IN0(n9752), .IN1(data_mem_out_wire[1146]), .SEL(n10433), .F(
        n6636) );
  MUX U11574 ( .IN0(n9753), .IN1(data_mem_out_wire[1145]), .SEL(n10433), .F(
        n6635) );
  MUX U11575 ( .IN0(n9754), .IN1(data_mem_out_wire[1144]), .SEL(n10433), .F(
        n6634) );
  AND U11576 ( .A(n10434), .B(n10435), .Z(n10433) );
  AND U11577 ( .A(n10436), .B(n10437), .Z(n10434) );
  OR U11578 ( .A(n9760), .B(n10438), .Z(n10437) );
  MUX U11579 ( .IN0(data_mem_out_wire[1143]), .IN1(n9761), .SEL(n10439), .F(
        n6633) );
  MUX U11580 ( .IN0(data_mem_out_wire[1142]), .IN1(n9763), .SEL(n10439), .F(
        n6632) );
  MUX U11581 ( .IN0(data_mem_out_wire[1141]), .IN1(n9764), .SEL(n10439), .F(
        n6631) );
  MUX U11582 ( .IN0(data_mem_out_wire[1140]), .IN1(n9765), .SEL(n10439), .F(
        n6630) );
  MUX U11583 ( .IN0(data_mem_out_wire[1139]), .IN1(n9766), .SEL(n10439), .F(
        n6629) );
  IV U11584 ( .A(n10440), .Z(n10439) );
  MUX U11585 ( .IN0(n9768), .IN1(data_mem_out_wire[1138]), .SEL(n10440), .F(
        n6628) );
  MUX U11586 ( .IN0(n9769), .IN1(data_mem_out_wire[1137]), .SEL(n10440), .F(
        n6627) );
  MUX U11587 ( .IN0(n9770), .IN1(data_mem_out_wire[1136]), .SEL(n10440), .F(
        n6626) );
  AND U11588 ( .A(n10441), .B(n10442), .Z(n10440) );
  OR U11589 ( .A(n9773), .B(n10438), .Z(n10442) );
  AND U11590 ( .A(n10436), .B(n10435), .Z(n10441) );
  NANDN U11591 ( .A(n10438), .B(n9809), .Z(n10436) );
  MUX U11592 ( .IN0(data_mem_out_wire[1135]), .IN1(n9776), .SEL(n10443), .F(
        n6625) );
  MUX U11593 ( .IN0(data_mem_out_wire[1134]), .IN1(n9778), .SEL(n10443), .F(
        n6624) );
  MUX U11594 ( .IN0(data_mem_out_wire[1133]), .IN1(n9779), .SEL(n10443), .F(
        n6623) );
  MUX U11595 ( .IN0(data_mem_out_wire[1132]), .IN1(n9780), .SEL(n10443), .F(
        n6622) );
  MUX U11596 ( .IN0(data_mem_out_wire[1131]), .IN1(n9781), .SEL(n10443), .F(
        n6621) );
  IV U11597 ( .A(n10444), .Z(n10443) );
  MUX U11598 ( .IN0(n9783), .IN1(data_mem_out_wire[1130]), .SEL(n10444), .F(
        n6620) );
  MUX U11599 ( .IN0(n9784), .IN1(data_mem_out_wire[1129]), .SEL(n10444), .F(
        n6619) );
  MUX U11600 ( .IN0(n9785), .IN1(data_mem_out_wire[1128]), .SEL(n10444), .F(
        n6618) );
  AND U11601 ( .A(n10445), .B(n10446), .Z(n10444) );
  OR U11602 ( .A(n9788), .B(n10438), .Z(n10446) );
  MUX U11603 ( .IN0(data_mem_out_wire[1127]), .IN1(data_in[7]), .SEL(n10447), 
        .F(n6617) );
  MUX U11604 ( .IN0(data_mem_out_wire[1126]), .IN1(data_in[6]), .SEL(n10447), 
        .F(n6616) );
  MUX U11605 ( .IN0(data_mem_out_wire[1125]), .IN1(data_in[5]), .SEL(n10447), 
        .F(n6615) );
  MUX U11606 ( .IN0(data_mem_out_wire[1124]), .IN1(data_in[4]), .SEL(n10447), 
        .F(n6614) );
  MUX U11607 ( .IN0(data_mem_out_wire[1123]), .IN1(data_in[3]), .SEL(n10447), 
        .F(n6613) );
  IV U11608 ( .A(n10448), .Z(n10447) );
  MUX U11609 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1122]), .SEL(n10448), 
        .F(n6612) );
  MUX U11610 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1121]), .SEL(n10448), 
        .F(n6611) );
  MUX U11611 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1120]), .SEL(n10448), 
        .F(n6610) );
  AND U11612 ( .A(n10445), .B(n10449), .Z(n10448) );
  NANDN U11613 ( .A(n10438), .B(n9792), .Z(n10449) );
  AND U11614 ( .A(n10450), .B(n10435), .Z(n10445) );
  NANDN U11615 ( .A(n10438), .B(n9796), .Z(n10435) );
  NANDN U11616 ( .A(n10438), .B(n9818), .Z(n10450) );
  NAND U11617 ( .A(n9862), .B(n10396), .Z(n10438) );
  MUX U11618 ( .IN0(n9746), .IN1(data_mem_out_wire[1183]), .SEL(n10451), .F(
        n6609) );
  MUX U11619 ( .IN0(n9748), .IN1(data_mem_out_wire[1182]), .SEL(n10451), .F(
        n6608) );
  MUX U11620 ( .IN0(n9749), .IN1(data_mem_out_wire[1181]), .SEL(n10451), .F(
        n6607) );
  MUX U11621 ( .IN0(n9750), .IN1(data_mem_out_wire[1180]), .SEL(n10451), .F(
        n6606) );
  MUX U11622 ( .IN0(n9751), .IN1(data_mem_out_wire[1179]), .SEL(n10451), .F(
        n6605) );
  MUX U11623 ( .IN0(n9752), .IN1(data_mem_out_wire[1178]), .SEL(n10451), .F(
        n6604) );
  MUX U11624 ( .IN0(n9753), .IN1(data_mem_out_wire[1177]), .SEL(n10451), .F(
        n6603) );
  MUX U11625 ( .IN0(n9754), .IN1(data_mem_out_wire[1176]), .SEL(n10451), .F(
        n6602) );
  AND U11626 ( .A(n10452), .B(n10453), .Z(n10451) );
  AND U11627 ( .A(n10454), .B(n10455), .Z(n10452) );
  OR U11628 ( .A(n9760), .B(n10456), .Z(n10455) );
  MUX U11629 ( .IN0(data_mem_out_wire[1175]), .IN1(n9761), .SEL(n10457), .F(
        n6601) );
  MUX U11630 ( .IN0(data_mem_out_wire[1174]), .IN1(n9763), .SEL(n10457), .F(
        n6600) );
  MUX U11631 ( .IN0(data_mem_out_wire[1173]), .IN1(n9764), .SEL(n10457), .F(
        n6599) );
  MUX U11632 ( .IN0(data_mem_out_wire[1172]), .IN1(n9765), .SEL(n10457), .F(
        n6598) );
  MUX U11633 ( .IN0(data_mem_out_wire[1171]), .IN1(n9766), .SEL(n10457), .F(
        n6597) );
  IV U11634 ( .A(n10458), .Z(n10457) );
  MUX U11635 ( .IN0(n9768), .IN1(data_mem_out_wire[1170]), .SEL(n10458), .F(
        n6596) );
  MUX U11636 ( .IN0(n9769), .IN1(data_mem_out_wire[1169]), .SEL(n10458), .F(
        n6595) );
  MUX U11637 ( .IN0(n9770), .IN1(data_mem_out_wire[1168]), .SEL(n10458), .F(
        n6594) );
  AND U11638 ( .A(n10459), .B(n10460), .Z(n10458) );
  OR U11639 ( .A(n9773), .B(n10456), .Z(n10460) );
  AND U11640 ( .A(n10454), .B(n10453), .Z(n10459) );
  NANDN U11641 ( .A(n10456), .B(n9809), .Z(n10454) );
  MUX U11642 ( .IN0(data_mem_out_wire[1167]), .IN1(n9776), .SEL(n10461), .F(
        n6593) );
  MUX U11643 ( .IN0(data_mem_out_wire[1166]), .IN1(n9778), .SEL(n10461), .F(
        n6592) );
  MUX U11644 ( .IN0(data_mem_out_wire[1165]), .IN1(n9779), .SEL(n10461), .F(
        n6591) );
  MUX U11645 ( .IN0(data_mem_out_wire[1164]), .IN1(n9780), .SEL(n10461), .F(
        n6590) );
  MUX U11646 ( .IN0(data_mem_out_wire[1163]), .IN1(n9781), .SEL(n10461), .F(
        n6589) );
  IV U11647 ( .A(n10462), .Z(n10461) );
  MUX U11648 ( .IN0(n9783), .IN1(data_mem_out_wire[1162]), .SEL(n10462), .F(
        n6588) );
  MUX U11649 ( .IN0(n9784), .IN1(data_mem_out_wire[1161]), .SEL(n10462), .F(
        n6587) );
  MUX U11650 ( .IN0(n9785), .IN1(data_mem_out_wire[1160]), .SEL(n10462), .F(
        n6586) );
  AND U11651 ( .A(n10463), .B(n10464), .Z(n10462) );
  OR U11652 ( .A(n9788), .B(n10456), .Z(n10464) );
  MUX U11653 ( .IN0(data_mem_out_wire[1159]), .IN1(data_in[7]), .SEL(n10465), 
        .F(n6585) );
  MUX U11654 ( .IN0(data_mem_out_wire[1158]), .IN1(data_in[6]), .SEL(n10465), 
        .F(n6584) );
  MUX U11655 ( .IN0(data_mem_out_wire[1157]), .IN1(data_in[5]), .SEL(n10465), 
        .F(n6583) );
  MUX U11656 ( .IN0(data_mem_out_wire[1156]), .IN1(data_in[4]), .SEL(n10465), 
        .F(n6582) );
  MUX U11657 ( .IN0(data_mem_out_wire[1155]), .IN1(data_in[3]), .SEL(n10465), 
        .F(n6581) );
  IV U11658 ( .A(n10466), .Z(n10465) );
  MUX U11659 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1154]), .SEL(n10466), 
        .F(n6580) );
  MUX U11660 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1153]), .SEL(n10466), 
        .F(n6579) );
  MUX U11661 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1152]), .SEL(n10466), 
        .F(n6578) );
  AND U11662 ( .A(n10463), .B(n10467), .Z(n10466) );
  NANDN U11663 ( .A(n10456), .B(n9792), .Z(n10467) );
  AND U11664 ( .A(n10468), .B(n10453), .Z(n10463) );
  NANDN U11665 ( .A(n10456), .B(n9796), .Z(n10453) );
  NANDN U11666 ( .A(n10456), .B(n9818), .Z(n10468) );
  NAND U11667 ( .A(n9881), .B(n10396), .Z(n10456) );
  MUX U11668 ( .IN0(n9746), .IN1(data_mem_out_wire[1215]), .SEL(n10469), .F(
        n6577) );
  MUX U11669 ( .IN0(n9748), .IN1(data_mem_out_wire[1214]), .SEL(n10469), .F(
        n6576) );
  MUX U11670 ( .IN0(n9749), .IN1(data_mem_out_wire[1213]), .SEL(n10469), .F(
        n6575) );
  MUX U11671 ( .IN0(n9750), .IN1(data_mem_out_wire[1212]), .SEL(n10469), .F(
        n6574) );
  MUX U11672 ( .IN0(n9751), .IN1(data_mem_out_wire[1211]), .SEL(n10469), .F(
        n6573) );
  MUX U11673 ( .IN0(n9752), .IN1(data_mem_out_wire[1210]), .SEL(n10469), .F(
        n6572) );
  MUX U11674 ( .IN0(n9753), .IN1(data_mem_out_wire[1209]), .SEL(n10469), .F(
        n6571) );
  MUX U11675 ( .IN0(n9754), .IN1(data_mem_out_wire[1208]), .SEL(n10469), .F(
        n6570) );
  AND U11676 ( .A(n10470), .B(n10471), .Z(n10469) );
  AND U11677 ( .A(n10472), .B(n10473), .Z(n10470) );
  OR U11678 ( .A(n9760), .B(n10474), .Z(n10473) );
  MUX U11679 ( .IN0(data_mem_out_wire[1207]), .IN1(n9761), .SEL(n10475), .F(
        n6569) );
  MUX U11680 ( .IN0(data_mem_out_wire[1206]), .IN1(n9763), .SEL(n10475), .F(
        n6568) );
  MUX U11681 ( .IN0(data_mem_out_wire[1205]), .IN1(n9764), .SEL(n10475), .F(
        n6567) );
  MUX U11682 ( .IN0(data_mem_out_wire[1204]), .IN1(n9765), .SEL(n10475), .F(
        n6566) );
  MUX U11683 ( .IN0(data_mem_out_wire[1203]), .IN1(n9766), .SEL(n10475), .F(
        n6565) );
  IV U11684 ( .A(n10476), .Z(n10475) );
  MUX U11685 ( .IN0(n9768), .IN1(data_mem_out_wire[1202]), .SEL(n10476), .F(
        n6564) );
  MUX U11686 ( .IN0(n9769), .IN1(data_mem_out_wire[1201]), .SEL(n10476), .F(
        n6563) );
  MUX U11687 ( .IN0(n9770), .IN1(data_mem_out_wire[1200]), .SEL(n10476), .F(
        n6562) );
  AND U11688 ( .A(n10477), .B(n10478), .Z(n10476) );
  OR U11689 ( .A(n9773), .B(n10474), .Z(n10478) );
  AND U11690 ( .A(n10472), .B(n10471), .Z(n10477) );
  NANDN U11691 ( .A(n10474), .B(n9809), .Z(n10472) );
  MUX U11692 ( .IN0(data_mem_out_wire[1199]), .IN1(n9776), .SEL(n10479), .F(
        n6561) );
  MUX U11693 ( .IN0(data_mem_out_wire[1198]), .IN1(n9778), .SEL(n10479), .F(
        n6560) );
  MUX U11694 ( .IN0(data_mem_out_wire[1197]), .IN1(n9779), .SEL(n10479), .F(
        n6559) );
  MUX U11695 ( .IN0(data_mem_out_wire[1196]), .IN1(n9780), .SEL(n10479), .F(
        n6558) );
  MUX U11696 ( .IN0(data_mem_out_wire[1195]), .IN1(n9781), .SEL(n10479), .F(
        n6557) );
  IV U11697 ( .A(n10480), .Z(n10479) );
  MUX U11698 ( .IN0(n9783), .IN1(data_mem_out_wire[1194]), .SEL(n10480), .F(
        n6556) );
  MUX U11699 ( .IN0(n9784), .IN1(data_mem_out_wire[1193]), .SEL(n10480), .F(
        n6555) );
  MUX U11700 ( .IN0(n9785), .IN1(data_mem_out_wire[1192]), .SEL(n10480), .F(
        n6554) );
  AND U11701 ( .A(n10481), .B(n10482), .Z(n10480) );
  OR U11702 ( .A(n9788), .B(n10474), .Z(n10482) );
  MUX U11703 ( .IN0(data_mem_out_wire[1191]), .IN1(data_in[7]), .SEL(n10483), 
        .F(n6553) );
  MUX U11704 ( .IN0(data_mem_out_wire[1190]), .IN1(data_in[6]), .SEL(n10483), 
        .F(n6552) );
  MUX U11705 ( .IN0(data_mem_out_wire[1189]), .IN1(data_in[5]), .SEL(n10483), 
        .F(n6551) );
  MUX U11706 ( .IN0(data_mem_out_wire[1188]), .IN1(data_in[4]), .SEL(n10483), 
        .F(n6550) );
  MUX U11707 ( .IN0(data_mem_out_wire[1187]), .IN1(data_in[3]), .SEL(n10483), 
        .F(n6549) );
  IV U11708 ( .A(n10484), .Z(n10483) );
  MUX U11709 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1186]), .SEL(n10484), 
        .F(n6548) );
  MUX U11710 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1185]), .SEL(n10484), 
        .F(n6547) );
  MUX U11711 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1184]), .SEL(n10484), 
        .F(n6546) );
  AND U11712 ( .A(n10481), .B(n10485), .Z(n10484) );
  NANDN U11713 ( .A(n10474), .B(n9792), .Z(n10485) );
  AND U11714 ( .A(n10486), .B(n10471), .Z(n10481) );
  NANDN U11715 ( .A(n10474), .B(n9796), .Z(n10471) );
  NANDN U11716 ( .A(n10474), .B(n9818), .Z(n10486) );
  NAND U11717 ( .A(n9900), .B(n10396), .Z(n10474) );
  MUX U11718 ( .IN0(n9746), .IN1(data_mem_out_wire[1247]), .SEL(n10487), .F(
        n6545) );
  MUX U11719 ( .IN0(n9748), .IN1(data_mem_out_wire[1246]), .SEL(n10487), .F(
        n6544) );
  MUX U11720 ( .IN0(n9749), .IN1(data_mem_out_wire[1245]), .SEL(n10487), .F(
        n6543) );
  MUX U11721 ( .IN0(n9750), .IN1(data_mem_out_wire[1244]), .SEL(n10487), .F(
        n6542) );
  MUX U11722 ( .IN0(n9751), .IN1(data_mem_out_wire[1243]), .SEL(n10487), .F(
        n6541) );
  MUX U11723 ( .IN0(n9752), .IN1(data_mem_out_wire[1242]), .SEL(n10487), .F(
        n6540) );
  MUX U11724 ( .IN0(n9753), .IN1(data_mem_out_wire[1241]), .SEL(n10487), .F(
        n6539) );
  MUX U11725 ( .IN0(n9754), .IN1(data_mem_out_wire[1240]), .SEL(n10487), .F(
        n6538) );
  AND U11726 ( .A(n10488), .B(n10489), .Z(n10487) );
  AND U11727 ( .A(n10490), .B(n10491), .Z(n10488) );
  OR U11728 ( .A(n9760), .B(n10492), .Z(n10491) );
  MUX U11729 ( .IN0(data_mem_out_wire[1239]), .IN1(n9761), .SEL(n10493), .F(
        n6537) );
  MUX U11730 ( .IN0(data_mem_out_wire[1238]), .IN1(n9763), .SEL(n10493), .F(
        n6536) );
  MUX U11731 ( .IN0(data_mem_out_wire[1237]), .IN1(n9764), .SEL(n10493), .F(
        n6535) );
  MUX U11732 ( .IN0(data_mem_out_wire[1236]), .IN1(n9765), .SEL(n10493), .F(
        n6534) );
  MUX U11733 ( .IN0(data_mem_out_wire[1235]), .IN1(n9766), .SEL(n10493), .F(
        n6533) );
  IV U11734 ( .A(n10494), .Z(n10493) );
  MUX U11735 ( .IN0(n9768), .IN1(data_mem_out_wire[1234]), .SEL(n10494), .F(
        n6532) );
  MUX U11736 ( .IN0(n9769), .IN1(data_mem_out_wire[1233]), .SEL(n10494), .F(
        n6531) );
  MUX U11737 ( .IN0(n9770), .IN1(data_mem_out_wire[1232]), .SEL(n10494), .F(
        n6530) );
  AND U11738 ( .A(n10495), .B(n10496), .Z(n10494) );
  OR U11739 ( .A(n9773), .B(n10492), .Z(n10496) );
  AND U11740 ( .A(n10490), .B(n10489), .Z(n10495) );
  NANDN U11741 ( .A(n10492), .B(n9809), .Z(n10490) );
  MUX U11742 ( .IN0(data_mem_out_wire[1231]), .IN1(n9776), .SEL(n10497), .F(
        n6529) );
  MUX U11743 ( .IN0(data_mem_out_wire[1230]), .IN1(n9778), .SEL(n10497), .F(
        n6528) );
  MUX U11744 ( .IN0(data_mem_out_wire[1229]), .IN1(n9779), .SEL(n10497), .F(
        n6527) );
  MUX U11745 ( .IN0(data_mem_out_wire[1228]), .IN1(n9780), .SEL(n10497), .F(
        n6526) );
  MUX U11746 ( .IN0(data_mem_out_wire[1227]), .IN1(n9781), .SEL(n10497), .F(
        n6525) );
  IV U11747 ( .A(n10498), .Z(n10497) );
  MUX U11748 ( .IN0(n9783), .IN1(data_mem_out_wire[1226]), .SEL(n10498), .F(
        n6524) );
  MUX U11749 ( .IN0(n9784), .IN1(data_mem_out_wire[1225]), .SEL(n10498), .F(
        n6523) );
  MUX U11750 ( .IN0(n9785), .IN1(data_mem_out_wire[1224]), .SEL(n10498), .F(
        n6522) );
  AND U11751 ( .A(n10499), .B(n10500), .Z(n10498) );
  OR U11752 ( .A(n9788), .B(n10492), .Z(n10500) );
  MUX U11753 ( .IN0(data_mem_out_wire[1223]), .IN1(data_in[7]), .SEL(n10501), 
        .F(n6521) );
  MUX U11754 ( .IN0(data_mem_out_wire[1222]), .IN1(data_in[6]), .SEL(n10501), 
        .F(n6520) );
  MUX U11755 ( .IN0(data_mem_out_wire[1221]), .IN1(data_in[5]), .SEL(n10501), 
        .F(n6519) );
  MUX U11756 ( .IN0(data_mem_out_wire[1220]), .IN1(data_in[4]), .SEL(n10501), 
        .F(n6518) );
  MUX U11757 ( .IN0(data_mem_out_wire[1219]), .IN1(data_in[3]), .SEL(n10501), 
        .F(n6517) );
  IV U11758 ( .A(n10502), .Z(n10501) );
  MUX U11759 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1218]), .SEL(n10502), 
        .F(n6516) );
  MUX U11760 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1217]), .SEL(n10502), 
        .F(n6515) );
  MUX U11761 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1216]), .SEL(n10502), 
        .F(n6514) );
  AND U11762 ( .A(n10499), .B(n10503), .Z(n10502) );
  NANDN U11763 ( .A(n10492), .B(n9792), .Z(n10503) );
  AND U11764 ( .A(n10504), .B(n10489), .Z(n10499) );
  NANDN U11765 ( .A(n10492), .B(n9796), .Z(n10489) );
  NANDN U11766 ( .A(n10492), .B(n9818), .Z(n10504) );
  NAND U11767 ( .A(n9919), .B(n10396), .Z(n10492) );
  MUX U11768 ( .IN0(n9746), .IN1(data_mem_out_wire[1279]), .SEL(n10505), .F(
        n6513) );
  MUX U11769 ( .IN0(n9748), .IN1(data_mem_out_wire[1278]), .SEL(n10505), .F(
        n6512) );
  MUX U11770 ( .IN0(n9749), .IN1(data_mem_out_wire[1277]), .SEL(n10505), .F(
        n6511) );
  MUX U11771 ( .IN0(n9750), .IN1(data_mem_out_wire[1276]), .SEL(n10505), .F(
        n6510) );
  MUX U11772 ( .IN0(n9751), .IN1(data_mem_out_wire[1275]), .SEL(n10505), .F(
        n6509) );
  MUX U11773 ( .IN0(n9752), .IN1(data_mem_out_wire[1274]), .SEL(n10505), .F(
        n6508) );
  MUX U11774 ( .IN0(n9753), .IN1(data_mem_out_wire[1273]), .SEL(n10505), .F(
        n6507) );
  MUX U11775 ( .IN0(n9754), .IN1(data_mem_out_wire[1272]), .SEL(n10505), .F(
        n6506) );
  AND U11776 ( .A(n10506), .B(n10507), .Z(n10505) );
  AND U11777 ( .A(n10508), .B(n10509), .Z(n10506) );
  OR U11778 ( .A(n9760), .B(n10510), .Z(n10509) );
  MUX U11779 ( .IN0(data_mem_out_wire[1271]), .IN1(n9761), .SEL(n10511), .F(
        n6505) );
  MUX U11780 ( .IN0(data_mem_out_wire[1270]), .IN1(n9763), .SEL(n10511), .F(
        n6504) );
  MUX U11781 ( .IN0(data_mem_out_wire[1269]), .IN1(n9764), .SEL(n10511), .F(
        n6503) );
  MUX U11782 ( .IN0(data_mem_out_wire[1268]), .IN1(n9765), .SEL(n10511), .F(
        n6502) );
  MUX U11783 ( .IN0(data_mem_out_wire[1267]), .IN1(n9766), .SEL(n10511), .F(
        n6501) );
  IV U11784 ( .A(n10512), .Z(n10511) );
  MUX U11785 ( .IN0(n9768), .IN1(data_mem_out_wire[1266]), .SEL(n10512), .F(
        n6500) );
  MUX U11786 ( .IN0(n9769), .IN1(data_mem_out_wire[1265]), .SEL(n10512), .F(
        n6499) );
  MUX U11787 ( .IN0(n9770), .IN1(data_mem_out_wire[1264]), .SEL(n10512), .F(
        n6498) );
  AND U11788 ( .A(n10513), .B(n10514), .Z(n10512) );
  OR U11789 ( .A(n9773), .B(n10510), .Z(n10514) );
  AND U11790 ( .A(n10508), .B(n10507), .Z(n10513) );
  NANDN U11791 ( .A(n10510), .B(n9809), .Z(n10508) );
  MUX U11792 ( .IN0(data_mem_out_wire[1263]), .IN1(n9776), .SEL(n10515), .F(
        n6497) );
  MUX U11793 ( .IN0(data_mem_out_wire[1262]), .IN1(n9778), .SEL(n10515), .F(
        n6496) );
  MUX U11794 ( .IN0(data_mem_out_wire[1261]), .IN1(n9779), .SEL(n10515), .F(
        n6495) );
  MUX U11795 ( .IN0(data_mem_out_wire[1260]), .IN1(n9780), .SEL(n10515), .F(
        n6494) );
  MUX U11796 ( .IN0(data_mem_out_wire[1259]), .IN1(n9781), .SEL(n10515), .F(
        n6493) );
  IV U11797 ( .A(n10516), .Z(n10515) );
  MUX U11798 ( .IN0(n9783), .IN1(data_mem_out_wire[1258]), .SEL(n10516), .F(
        n6492) );
  MUX U11799 ( .IN0(n9784), .IN1(data_mem_out_wire[1257]), .SEL(n10516), .F(
        n6491) );
  MUX U11800 ( .IN0(n9785), .IN1(data_mem_out_wire[1256]), .SEL(n10516), .F(
        n6490) );
  AND U11801 ( .A(n10517), .B(n10518), .Z(n10516) );
  OR U11802 ( .A(n9788), .B(n10510), .Z(n10518) );
  MUX U11803 ( .IN0(data_mem_out_wire[1255]), .IN1(data_in[7]), .SEL(n10519), 
        .F(n6489) );
  MUX U11804 ( .IN0(data_mem_out_wire[1254]), .IN1(data_in[6]), .SEL(n10519), 
        .F(n6488) );
  MUX U11805 ( .IN0(data_mem_out_wire[1253]), .IN1(data_in[5]), .SEL(n10519), 
        .F(n6487) );
  MUX U11806 ( .IN0(data_mem_out_wire[1252]), .IN1(data_in[4]), .SEL(n10519), 
        .F(n6486) );
  MUX U11807 ( .IN0(data_mem_out_wire[1251]), .IN1(data_in[3]), .SEL(n10519), 
        .F(n6485) );
  IV U11808 ( .A(n10520), .Z(n10519) );
  MUX U11809 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1250]), .SEL(n10520), 
        .F(n6484) );
  MUX U11810 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1249]), .SEL(n10520), 
        .F(n6483) );
  MUX U11811 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1248]), .SEL(n10520), 
        .F(n6482) );
  AND U11812 ( .A(n10517), .B(n10521), .Z(n10520) );
  NANDN U11813 ( .A(n10510), .B(n9792), .Z(n10521) );
  AND U11814 ( .A(n10522), .B(n10507), .Z(n10517) );
  NANDN U11815 ( .A(n10510), .B(n9796), .Z(n10507) );
  NANDN U11816 ( .A(n10510), .B(n9818), .Z(n10522) );
  NAND U11817 ( .A(n10396), .B(n9938), .Z(n10510) );
  AND U11818 ( .A(n9939), .B(N42), .Z(n10396) );
  NOR U11819 ( .A(N41), .B(N40), .Z(n9939) );
  MUX U11820 ( .IN0(n9746), .IN1(data_mem_out_wire[1311]), .SEL(n10523), .F(
        n6481) );
  MUX U11821 ( .IN0(n9748), .IN1(data_mem_out_wire[1310]), .SEL(n10523), .F(
        n6480) );
  MUX U11822 ( .IN0(n9749), .IN1(data_mem_out_wire[1309]), .SEL(n10523), .F(
        n6479) );
  MUX U11823 ( .IN0(n9750), .IN1(data_mem_out_wire[1308]), .SEL(n10523), .F(
        n6478) );
  MUX U11824 ( .IN0(n9751), .IN1(data_mem_out_wire[1307]), .SEL(n10523), .F(
        n6477) );
  MUX U11825 ( .IN0(n9752), .IN1(data_mem_out_wire[1306]), .SEL(n10523), .F(
        n6476) );
  MUX U11826 ( .IN0(n9753), .IN1(data_mem_out_wire[1305]), .SEL(n10523), .F(
        n6475) );
  MUX U11827 ( .IN0(n9754), .IN1(data_mem_out_wire[1304]), .SEL(n10523), .F(
        n6474) );
  AND U11828 ( .A(n10524), .B(n10525), .Z(n10523) );
  AND U11829 ( .A(n10526), .B(n10527), .Z(n10524) );
  OR U11830 ( .A(n9760), .B(n10528), .Z(n10527) );
  MUX U11831 ( .IN0(data_mem_out_wire[1303]), .IN1(n9761), .SEL(n10529), .F(
        n6473) );
  MUX U11832 ( .IN0(data_mem_out_wire[1302]), .IN1(n9763), .SEL(n10529), .F(
        n6472) );
  MUX U11833 ( .IN0(data_mem_out_wire[1301]), .IN1(n9764), .SEL(n10529), .F(
        n6471) );
  MUX U11834 ( .IN0(data_mem_out_wire[1300]), .IN1(n9765), .SEL(n10529), .F(
        n6470) );
  MUX U11835 ( .IN0(data_mem_out_wire[1299]), .IN1(n9766), .SEL(n10529), .F(
        n6469) );
  IV U11836 ( .A(n10530), .Z(n10529) );
  MUX U11837 ( .IN0(n9768), .IN1(data_mem_out_wire[1298]), .SEL(n10530), .F(
        n6468) );
  MUX U11838 ( .IN0(n9769), .IN1(data_mem_out_wire[1297]), .SEL(n10530), .F(
        n6467) );
  MUX U11839 ( .IN0(n9770), .IN1(data_mem_out_wire[1296]), .SEL(n10530), .F(
        n6466) );
  AND U11840 ( .A(n10531), .B(n10532), .Z(n10530) );
  OR U11841 ( .A(n9773), .B(n10528), .Z(n10532) );
  AND U11842 ( .A(n10526), .B(n10525), .Z(n10531) );
  NANDN U11843 ( .A(n10528), .B(n9809), .Z(n10526) );
  MUX U11844 ( .IN0(data_mem_out_wire[1295]), .IN1(n9776), .SEL(n10533), .F(
        n6465) );
  MUX U11845 ( .IN0(data_mem_out_wire[1294]), .IN1(n9778), .SEL(n10533), .F(
        n6464) );
  MUX U11846 ( .IN0(data_mem_out_wire[1293]), .IN1(n9779), .SEL(n10533), .F(
        n6463) );
  MUX U11847 ( .IN0(data_mem_out_wire[1292]), .IN1(n9780), .SEL(n10533), .F(
        n6462) );
  MUX U11848 ( .IN0(data_mem_out_wire[1291]), .IN1(n9781), .SEL(n10533), .F(
        n6461) );
  IV U11849 ( .A(n10534), .Z(n10533) );
  MUX U11850 ( .IN0(n9783), .IN1(data_mem_out_wire[1290]), .SEL(n10534), .F(
        n6460) );
  MUX U11851 ( .IN0(n9784), .IN1(data_mem_out_wire[1289]), .SEL(n10534), .F(
        n6459) );
  MUX U11852 ( .IN0(n9785), .IN1(data_mem_out_wire[1288]), .SEL(n10534), .F(
        n6458) );
  AND U11853 ( .A(n10535), .B(n10536), .Z(n10534) );
  OR U11854 ( .A(n9788), .B(n10528), .Z(n10536) );
  MUX U11855 ( .IN0(data_mem_out_wire[1287]), .IN1(data_in[7]), .SEL(n10537), 
        .F(n6457) );
  MUX U11856 ( .IN0(data_mem_out_wire[1286]), .IN1(data_in[6]), .SEL(n10537), 
        .F(n6456) );
  MUX U11857 ( .IN0(data_mem_out_wire[1285]), .IN1(data_in[5]), .SEL(n10537), 
        .F(n6455) );
  MUX U11858 ( .IN0(data_mem_out_wire[1284]), .IN1(data_in[4]), .SEL(n10537), 
        .F(n6454) );
  MUX U11859 ( .IN0(data_mem_out_wire[1283]), .IN1(data_in[3]), .SEL(n10537), 
        .F(n6453) );
  IV U11860 ( .A(n10538), .Z(n10537) );
  MUX U11861 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1282]), .SEL(n10538), 
        .F(n6452) );
  MUX U11862 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1281]), .SEL(n10538), 
        .F(n6451) );
  MUX U11863 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1280]), .SEL(n10538), 
        .F(n6450) );
  AND U11864 ( .A(n10535), .B(n10539), .Z(n10538) );
  NANDN U11865 ( .A(n10528), .B(n9792), .Z(n10539) );
  AND U11866 ( .A(n10540), .B(n10525), .Z(n10535) );
  NANDN U11867 ( .A(n10528), .B(n9796), .Z(n10525) );
  NANDN U11868 ( .A(n10528), .B(n9818), .Z(n10540) );
  NAND U11869 ( .A(n9798), .B(n10541), .Z(n10528) );
  MUX U11870 ( .IN0(n9746), .IN1(data_mem_out_wire[1343]), .SEL(n10542), .F(
        n6449) );
  MUX U11871 ( .IN0(n9748), .IN1(data_mem_out_wire[1342]), .SEL(n10542), .F(
        n6448) );
  MUX U11872 ( .IN0(n9749), .IN1(data_mem_out_wire[1341]), .SEL(n10542), .F(
        n6447) );
  MUX U11873 ( .IN0(n9750), .IN1(data_mem_out_wire[1340]), .SEL(n10542), .F(
        n6446) );
  MUX U11874 ( .IN0(n9751), .IN1(data_mem_out_wire[1339]), .SEL(n10542), .F(
        n6445) );
  MUX U11875 ( .IN0(n9752), .IN1(data_mem_out_wire[1338]), .SEL(n10542), .F(
        n6444) );
  MUX U11876 ( .IN0(n9753), .IN1(data_mem_out_wire[1337]), .SEL(n10542), .F(
        n6443) );
  MUX U11877 ( .IN0(n9754), .IN1(data_mem_out_wire[1336]), .SEL(n10542), .F(
        n6442) );
  AND U11878 ( .A(n10543), .B(n10544), .Z(n10542) );
  AND U11879 ( .A(n10545), .B(n10546), .Z(n10543) );
  OR U11880 ( .A(n9760), .B(n10547), .Z(n10546) );
  MUX U11881 ( .IN0(data_mem_out_wire[1335]), .IN1(n9761), .SEL(n10548), .F(
        n6441) );
  MUX U11882 ( .IN0(data_mem_out_wire[1334]), .IN1(n9763), .SEL(n10548), .F(
        n6440) );
  MUX U11883 ( .IN0(data_mem_out_wire[1333]), .IN1(n9764), .SEL(n10548), .F(
        n6439) );
  MUX U11884 ( .IN0(data_mem_out_wire[1332]), .IN1(n9765), .SEL(n10548), .F(
        n6438) );
  MUX U11885 ( .IN0(data_mem_out_wire[1331]), .IN1(n9766), .SEL(n10548), .F(
        n6437) );
  IV U11886 ( .A(n10549), .Z(n10548) );
  MUX U11887 ( .IN0(n9768), .IN1(data_mem_out_wire[1330]), .SEL(n10549), .F(
        n6436) );
  MUX U11888 ( .IN0(n9769), .IN1(data_mem_out_wire[1329]), .SEL(n10549), .F(
        n6435) );
  MUX U11889 ( .IN0(n9770), .IN1(data_mem_out_wire[1328]), .SEL(n10549), .F(
        n6434) );
  AND U11890 ( .A(n10550), .B(n10551), .Z(n10549) );
  OR U11891 ( .A(n9773), .B(n10547), .Z(n10551) );
  AND U11892 ( .A(n10545), .B(n10544), .Z(n10550) );
  NANDN U11893 ( .A(n10547), .B(n9809), .Z(n10545) );
  MUX U11894 ( .IN0(data_mem_out_wire[1327]), .IN1(n9776), .SEL(n10552), .F(
        n6433) );
  MUX U11895 ( .IN0(data_mem_out_wire[1326]), .IN1(n9778), .SEL(n10552), .F(
        n6432) );
  MUX U11896 ( .IN0(data_mem_out_wire[1325]), .IN1(n9779), .SEL(n10552), .F(
        n6431) );
  MUX U11897 ( .IN0(data_mem_out_wire[1324]), .IN1(n9780), .SEL(n10552), .F(
        n6430) );
  MUX U11898 ( .IN0(data_mem_out_wire[1323]), .IN1(n9781), .SEL(n10552), .F(
        n6429) );
  IV U11899 ( .A(n10553), .Z(n10552) );
  MUX U11900 ( .IN0(n9783), .IN1(data_mem_out_wire[1322]), .SEL(n10553), .F(
        n6428) );
  MUX U11901 ( .IN0(n9784), .IN1(data_mem_out_wire[1321]), .SEL(n10553), .F(
        n6427) );
  MUX U11902 ( .IN0(n9785), .IN1(data_mem_out_wire[1320]), .SEL(n10553), .F(
        n6426) );
  AND U11903 ( .A(n10554), .B(n10555), .Z(n10553) );
  OR U11904 ( .A(n9788), .B(n10547), .Z(n10555) );
  MUX U11905 ( .IN0(data_mem_out_wire[1319]), .IN1(data_in[7]), .SEL(n10556), 
        .F(n6425) );
  MUX U11906 ( .IN0(data_mem_out_wire[1318]), .IN1(data_in[6]), .SEL(n10556), 
        .F(n6424) );
  MUX U11907 ( .IN0(data_mem_out_wire[1317]), .IN1(data_in[5]), .SEL(n10556), 
        .F(n6423) );
  MUX U11908 ( .IN0(data_mem_out_wire[1316]), .IN1(data_in[4]), .SEL(n10556), 
        .F(n6422) );
  MUX U11909 ( .IN0(data_mem_out_wire[1315]), .IN1(data_in[3]), .SEL(n10556), 
        .F(n6421) );
  IV U11910 ( .A(n10557), .Z(n10556) );
  MUX U11911 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1314]), .SEL(n10557), 
        .F(n6420) );
  MUX U11912 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1313]), .SEL(n10557), 
        .F(n6419) );
  MUX U11913 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1312]), .SEL(n10557), 
        .F(n6418) );
  AND U11914 ( .A(n10554), .B(n10558), .Z(n10557) );
  NANDN U11915 ( .A(n10547), .B(n9792), .Z(n10558) );
  AND U11916 ( .A(n10559), .B(n10544), .Z(n10554) );
  NANDN U11917 ( .A(n10547), .B(n9796), .Z(n10544) );
  NANDN U11918 ( .A(n10547), .B(n9818), .Z(n10559) );
  NAND U11919 ( .A(n9819), .B(n10541), .Z(n10547) );
  MUX U11920 ( .IN0(n9746), .IN1(data_mem_out_wire[1375]), .SEL(n10560), .F(
        n6417) );
  MUX U11921 ( .IN0(n9748), .IN1(data_mem_out_wire[1374]), .SEL(n10560), .F(
        n6416) );
  MUX U11922 ( .IN0(n9749), .IN1(data_mem_out_wire[1373]), .SEL(n10560), .F(
        n6415) );
  MUX U11923 ( .IN0(n9750), .IN1(data_mem_out_wire[1372]), .SEL(n10560), .F(
        n6414) );
  MUX U11924 ( .IN0(n9751), .IN1(data_mem_out_wire[1371]), .SEL(n10560), .F(
        n6413) );
  MUX U11925 ( .IN0(n9752), .IN1(data_mem_out_wire[1370]), .SEL(n10560), .F(
        n6412) );
  MUX U11926 ( .IN0(n9753), .IN1(data_mem_out_wire[1369]), .SEL(n10560), .F(
        n6411) );
  MUX U11927 ( .IN0(n9754), .IN1(data_mem_out_wire[1368]), .SEL(n10560), .F(
        n6410) );
  AND U11928 ( .A(n10561), .B(n10562), .Z(n10560) );
  AND U11929 ( .A(n10563), .B(n10564), .Z(n10561) );
  OR U11930 ( .A(n9760), .B(n10565), .Z(n10564) );
  MUX U11931 ( .IN0(data_mem_out_wire[1367]), .IN1(n9761), .SEL(n10566), .F(
        n6409) );
  MUX U11932 ( .IN0(data_mem_out_wire[1366]), .IN1(n9763), .SEL(n10566), .F(
        n6408) );
  MUX U11933 ( .IN0(data_mem_out_wire[1365]), .IN1(n9764), .SEL(n10566), .F(
        n6407) );
  MUX U11934 ( .IN0(data_mem_out_wire[1364]), .IN1(n9765), .SEL(n10566), .F(
        n6406) );
  MUX U11935 ( .IN0(data_mem_out_wire[1363]), .IN1(n9766), .SEL(n10566), .F(
        n6405) );
  IV U11936 ( .A(n10567), .Z(n10566) );
  MUX U11937 ( .IN0(n9768), .IN1(data_mem_out_wire[1362]), .SEL(n10567), .F(
        n6404) );
  MUX U11938 ( .IN0(n9769), .IN1(data_mem_out_wire[1361]), .SEL(n10567), .F(
        n6403) );
  MUX U11939 ( .IN0(n9770), .IN1(data_mem_out_wire[1360]), .SEL(n10567), .F(
        n6402) );
  AND U11940 ( .A(n10568), .B(n10569), .Z(n10567) );
  OR U11941 ( .A(n9773), .B(n10565), .Z(n10569) );
  AND U11942 ( .A(n10563), .B(n10562), .Z(n10568) );
  NANDN U11943 ( .A(n10565), .B(n9809), .Z(n10563) );
  MUX U11944 ( .IN0(data_mem_out_wire[1359]), .IN1(n9776), .SEL(n10570), .F(
        n6401) );
  MUX U11945 ( .IN0(data_mem_out_wire[1358]), .IN1(n9778), .SEL(n10570), .F(
        n6400) );
  MUX U11946 ( .IN0(data_mem_out_wire[1357]), .IN1(n9779), .SEL(n10570), .F(
        n6399) );
  MUX U11947 ( .IN0(data_mem_out_wire[1356]), .IN1(n9780), .SEL(n10570), .F(
        n6398) );
  MUX U11948 ( .IN0(data_mem_out_wire[1355]), .IN1(n9781), .SEL(n10570), .F(
        n6397) );
  IV U11949 ( .A(n10571), .Z(n10570) );
  MUX U11950 ( .IN0(n9783), .IN1(data_mem_out_wire[1354]), .SEL(n10571), .F(
        n6396) );
  MUX U11951 ( .IN0(n9784), .IN1(data_mem_out_wire[1353]), .SEL(n10571), .F(
        n6395) );
  MUX U11952 ( .IN0(n9785), .IN1(data_mem_out_wire[1352]), .SEL(n10571), .F(
        n6394) );
  AND U11953 ( .A(n10572), .B(n10573), .Z(n10571) );
  OR U11954 ( .A(n9788), .B(n10565), .Z(n10573) );
  MUX U11955 ( .IN0(data_mem_out_wire[1351]), .IN1(data_in[7]), .SEL(n10574), 
        .F(n6393) );
  MUX U11956 ( .IN0(data_mem_out_wire[1350]), .IN1(data_in[6]), .SEL(n10574), 
        .F(n6392) );
  MUX U11957 ( .IN0(data_mem_out_wire[1349]), .IN1(data_in[5]), .SEL(n10574), 
        .F(n6391) );
  MUX U11958 ( .IN0(data_mem_out_wire[1348]), .IN1(data_in[4]), .SEL(n10574), 
        .F(n6390) );
  MUX U11959 ( .IN0(data_mem_out_wire[1347]), .IN1(data_in[3]), .SEL(n10574), 
        .F(n6389) );
  IV U11960 ( .A(n10575), .Z(n10574) );
  MUX U11961 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1346]), .SEL(n10575), 
        .F(n6388) );
  MUX U11962 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1345]), .SEL(n10575), 
        .F(n6387) );
  MUX U11963 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1344]), .SEL(n10575), 
        .F(n6386) );
  AND U11964 ( .A(n10572), .B(n10576), .Z(n10575) );
  NANDN U11965 ( .A(n10565), .B(n9792), .Z(n10576) );
  AND U11966 ( .A(n10577), .B(n10562), .Z(n10572) );
  NANDN U11967 ( .A(n10565), .B(n9796), .Z(n10562) );
  NANDN U11968 ( .A(n10565), .B(n9818), .Z(n10577) );
  NAND U11969 ( .A(n9838), .B(n10541), .Z(n10565) );
  MUX U11970 ( .IN0(n9746), .IN1(data_mem_out_wire[1407]), .SEL(n10578), .F(
        n6385) );
  MUX U11971 ( .IN0(n9748), .IN1(data_mem_out_wire[1406]), .SEL(n10578), .F(
        n6384) );
  MUX U11972 ( .IN0(n9749), .IN1(data_mem_out_wire[1405]), .SEL(n10578), .F(
        n6383) );
  MUX U11973 ( .IN0(n9750), .IN1(data_mem_out_wire[1404]), .SEL(n10578), .F(
        n6382) );
  MUX U11974 ( .IN0(n9751), .IN1(data_mem_out_wire[1403]), .SEL(n10578), .F(
        n6381) );
  MUX U11975 ( .IN0(n9752), .IN1(data_mem_out_wire[1402]), .SEL(n10578), .F(
        n6380) );
  MUX U11976 ( .IN0(n9753), .IN1(data_mem_out_wire[1401]), .SEL(n10578), .F(
        n6379) );
  MUX U11977 ( .IN0(n9754), .IN1(data_mem_out_wire[1400]), .SEL(n10578), .F(
        n6378) );
  AND U11978 ( .A(n10579), .B(n10580), .Z(n10578) );
  AND U11979 ( .A(n10581), .B(n10582), .Z(n10579) );
  OR U11980 ( .A(n9760), .B(n10583), .Z(n10582) );
  MUX U11981 ( .IN0(data_mem_out_wire[1399]), .IN1(n9761), .SEL(n10584), .F(
        n6377) );
  MUX U11982 ( .IN0(data_mem_out_wire[1398]), .IN1(n9763), .SEL(n10584), .F(
        n6376) );
  MUX U11983 ( .IN0(data_mem_out_wire[1397]), .IN1(n9764), .SEL(n10584), .F(
        n6375) );
  MUX U11984 ( .IN0(data_mem_out_wire[1396]), .IN1(n9765), .SEL(n10584), .F(
        n6374) );
  MUX U11985 ( .IN0(data_mem_out_wire[1395]), .IN1(n9766), .SEL(n10584), .F(
        n6373) );
  IV U11986 ( .A(n10585), .Z(n10584) );
  MUX U11987 ( .IN0(n9768), .IN1(data_mem_out_wire[1394]), .SEL(n10585), .F(
        n6372) );
  MUX U11988 ( .IN0(n9769), .IN1(data_mem_out_wire[1393]), .SEL(n10585), .F(
        n6371) );
  MUX U11989 ( .IN0(n9770), .IN1(data_mem_out_wire[1392]), .SEL(n10585), .F(
        n6370) );
  AND U11990 ( .A(n10586), .B(n10587), .Z(n10585) );
  OR U11991 ( .A(n9773), .B(n10583), .Z(n10587) );
  AND U11992 ( .A(n10581), .B(n10580), .Z(n10586) );
  NANDN U11993 ( .A(n10583), .B(n9809), .Z(n10581) );
  MUX U11994 ( .IN0(data_mem_out_wire[1391]), .IN1(n9776), .SEL(n10588), .F(
        n6369) );
  MUX U11995 ( .IN0(data_mem_out_wire[1390]), .IN1(n9778), .SEL(n10588), .F(
        n6368) );
  MUX U11996 ( .IN0(data_mem_out_wire[1389]), .IN1(n9779), .SEL(n10588), .F(
        n6367) );
  MUX U11997 ( .IN0(data_mem_out_wire[1388]), .IN1(n9780), .SEL(n10588), .F(
        n6366) );
  MUX U11998 ( .IN0(data_mem_out_wire[1387]), .IN1(n9781), .SEL(n10588), .F(
        n6365) );
  IV U11999 ( .A(n10589), .Z(n10588) );
  MUX U12000 ( .IN0(n9783), .IN1(data_mem_out_wire[1386]), .SEL(n10589), .F(
        n6364) );
  MUX U12001 ( .IN0(n9784), .IN1(data_mem_out_wire[1385]), .SEL(n10589), .F(
        n6363) );
  MUX U12002 ( .IN0(n9785), .IN1(data_mem_out_wire[1384]), .SEL(n10589), .F(
        n6362) );
  AND U12003 ( .A(n10590), .B(n10591), .Z(n10589) );
  OR U12004 ( .A(n9788), .B(n10583), .Z(n10591) );
  MUX U12005 ( .IN0(data_mem_out_wire[1383]), .IN1(data_in[7]), .SEL(n10592), 
        .F(n6361) );
  MUX U12006 ( .IN0(data_mem_out_wire[1382]), .IN1(data_in[6]), .SEL(n10592), 
        .F(n6360) );
  MUX U12007 ( .IN0(data_mem_out_wire[1381]), .IN1(data_in[5]), .SEL(n10592), 
        .F(n6359) );
  MUX U12008 ( .IN0(data_mem_out_wire[1380]), .IN1(data_in[4]), .SEL(n10592), 
        .F(n6358) );
  MUX U12009 ( .IN0(data_mem_out_wire[1379]), .IN1(data_in[3]), .SEL(n10592), 
        .F(n6357) );
  IV U12010 ( .A(n10593), .Z(n10592) );
  MUX U12011 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1378]), .SEL(n10593), 
        .F(n6356) );
  MUX U12012 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1377]), .SEL(n10593), 
        .F(n6355) );
  MUX U12013 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1376]), .SEL(n10593), 
        .F(n6354) );
  AND U12014 ( .A(n10590), .B(n10594), .Z(n10593) );
  NANDN U12015 ( .A(n10583), .B(n9792), .Z(n10594) );
  AND U12016 ( .A(n10595), .B(n10580), .Z(n10590) );
  NANDN U12017 ( .A(n10583), .B(n9796), .Z(n10580) );
  NANDN U12018 ( .A(n10583), .B(n9818), .Z(n10595) );
  NAND U12019 ( .A(n9862), .B(n10541), .Z(n10583) );
  MUX U12020 ( .IN0(n9746), .IN1(data_mem_out_wire[1439]), .SEL(n10596), .F(
        n6353) );
  MUX U12021 ( .IN0(n9748), .IN1(data_mem_out_wire[1438]), .SEL(n10596), .F(
        n6352) );
  MUX U12022 ( .IN0(n9749), .IN1(data_mem_out_wire[1437]), .SEL(n10596), .F(
        n6351) );
  MUX U12023 ( .IN0(n9750), .IN1(data_mem_out_wire[1436]), .SEL(n10596), .F(
        n6350) );
  MUX U12024 ( .IN0(n9751), .IN1(data_mem_out_wire[1435]), .SEL(n10596), .F(
        n6349) );
  MUX U12025 ( .IN0(n9752), .IN1(data_mem_out_wire[1434]), .SEL(n10596), .F(
        n6348) );
  MUX U12026 ( .IN0(n9753), .IN1(data_mem_out_wire[1433]), .SEL(n10596), .F(
        n6347) );
  MUX U12027 ( .IN0(n9754), .IN1(data_mem_out_wire[1432]), .SEL(n10596), .F(
        n6346) );
  AND U12028 ( .A(n10597), .B(n10598), .Z(n10596) );
  AND U12029 ( .A(n10599), .B(n10600), .Z(n10597) );
  OR U12030 ( .A(n9760), .B(n10601), .Z(n10600) );
  MUX U12031 ( .IN0(data_mem_out_wire[1431]), .IN1(n9761), .SEL(n10602), .F(
        n6345) );
  MUX U12032 ( .IN0(data_mem_out_wire[1430]), .IN1(n9763), .SEL(n10602), .F(
        n6344) );
  MUX U12033 ( .IN0(data_mem_out_wire[1429]), .IN1(n9764), .SEL(n10602), .F(
        n6343) );
  MUX U12034 ( .IN0(data_mem_out_wire[1428]), .IN1(n9765), .SEL(n10602), .F(
        n6342) );
  MUX U12035 ( .IN0(data_mem_out_wire[1427]), .IN1(n9766), .SEL(n10602), .F(
        n6341) );
  IV U12036 ( .A(n10603), .Z(n10602) );
  MUX U12037 ( .IN0(n9768), .IN1(data_mem_out_wire[1426]), .SEL(n10603), .F(
        n6340) );
  MUX U12038 ( .IN0(n9769), .IN1(data_mem_out_wire[1425]), .SEL(n10603), .F(
        n6339) );
  MUX U12039 ( .IN0(n9770), .IN1(data_mem_out_wire[1424]), .SEL(n10603), .F(
        n6338) );
  AND U12040 ( .A(n10604), .B(n10605), .Z(n10603) );
  OR U12041 ( .A(n9773), .B(n10601), .Z(n10605) );
  AND U12042 ( .A(n10599), .B(n10598), .Z(n10604) );
  NANDN U12043 ( .A(n10601), .B(n9809), .Z(n10599) );
  MUX U12044 ( .IN0(data_mem_out_wire[1423]), .IN1(n9776), .SEL(n10606), .F(
        n6337) );
  MUX U12045 ( .IN0(data_mem_out_wire[1422]), .IN1(n9778), .SEL(n10606), .F(
        n6336) );
  MUX U12046 ( .IN0(data_mem_out_wire[1421]), .IN1(n9779), .SEL(n10606), .F(
        n6335) );
  MUX U12047 ( .IN0(data_mem_out_wire[1420]), .IN1(n9780), .SEL(n10606), .F(
        n6334) );
  MUX U12048 ( .IN0(data_mem_out_wire[1419]), .IN1(n9781), .SEL(n10606), .F(
        n6333) );
  IV U12049 ( .A(n10607), .Z(n10606) );
  MUX U12050 ( .IN0(n9783), .IN1(data_mem_out_wire[1418]), .SEL(n10607), .F(
        n6332) );
  MUX U12051 ( .IN0(n9784), .IN1(data_mem_out_wire[1417]), .SEL(n10607), .F(
        n6331) );
  MUX U12052 ( .IN0(n9785), .IN1(data_mem_out_wire[1416]), .SEL(n10607), .F(
        n6330) );
  AND U12053 ( .A(n10608), .B(n10609), .Z(n10607) );
  OR U12054 ( .A(n9788), .B(n10601), .Z(n10609) );
  MUX U12055 ( .IN0(data_mem_out_wire[1415]), .IN1(data_in[7]), .SEL(n10610), 
        .F(n6329) );
  MUX U12056 ( .IN0(data_mem_out_wire[1414]), .IN1(data_in[6]), .SEL(n10610), 
        .F(n6328) );
  MUX U12057 ( .IN0(data_mem_out_wire[1413]), .IN1(data_in[5]), .SEL(n10610), 
        .F(n6327) );
  MUX U12058 ( .IN0(data_mem_out_wire[1412]), .IN1(data_in[4]), .SEL(n10610), 
        .F(n6326) );
  MUX U12059 ( .IN0(data_mem_out_wire[1411]), .IN1(data_in[3]), .SEL(n10610), 
        .F(n6325) );
  IV U12060 ( .A(n10611), .Z(n10610) );
  MUX U12061 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1410]), .SEL(n10611), 
        .F(n6324) );
  MUX U12062 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1409]), .SEL(n10611), 
        .F(n6323) );
  MUX U12063 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1408]), .SEL(n10611), 
        .F(n6322) );
  AND U12064 ( .A(n10608), .B(n10612), .Z(n10611) );
  NANDN U12065 ( .A(n10601), .B(n9792), .Z(n10612) );
  AND U12066 ( .A(n10613), .B(n10598), .Z(n10608) );
  NANDN U12067 ( .A(n10601), .B(n9796), .Z(n10598) );
  NANDN U12068 ( .A(n10601), .B(n9818), .Z(n10613) );
  NAND U12069 ( .A(n9881), .B(n10541), .Z(n10601) );
  MUX U12070 ( .IN0(n9746), .IN1(data_mem_out_wire[1471]), .SEL(n10614), .F(
        n6321) );
  MUX U12071 ( .IN0(n9748), .IN1(data_mem_out_wire[1470]), .SEL(n10614), .F(
        n6320) );
  MUX U12072 ( .IN0(n9749), .IN1(data_mem_out_wire[1469]), .SEL(n10614), .F(
        n6319) );
  MUX U12073 ( .IN0(n9750), .IN1(data_mem_out_wire[1468]), .SEL(n10614), .F(
        n6318) );
  MUX U12074 ( .IN0(n9751), .IN1(data_mem_out_wire[1467]), .SEL(n10614), .F(
        n6317) );
  MUX U12075 ( .IN0(n9752), .IN1(data_mem_out_wire[1466]), .SEL(n10614), .F(
        n6316) );
  MUX U12076 ( .IN0(n9753), .IN1(data_mem_out_wire[1465]), .SEL(n10614), .F(
        n6315) );
  MUX U12077 ( .IN0(n9754), .IN1(data_mem_out_wire[1464]), .SEL(n10614), .F(
        n6314) );
  AND U12078 ( .A(n10615), .B(n10616), .Z(n10614) );
  AND U12079 ( .A(n10617), .B(n10618), .Z(n10615) );
  OR U12080 ( .A(n9760), .B(n10619), .Z(n10618) );
  MUX U12081 ( .IN0(data_mem_out_wire[1463]), .IN1(n9761), .SEL(n10620), .F(
        n6313) );
  MUX U12082 ( .IN0(data_mem_out_wire[1462]), .IN1(n9763), .SEL(n10620), .F(
        n6312) );
  MUX U12083 ( .IN0(data_mem_out_wire[1461]), .IN1(n9764), .SEL(n10620), .F(
        n6311) );
  MUX U12084 ( .IN0(data_mem_out_wire[1460]), .IN1(n9765), .SEL(n10620), .F(
        n6310) );
  MUX U12085 ( .IN0(data_mem_out_wire[1459]), .IN1(n9766), .SEL(n10620), .F(
        n6309) );
  IV U12086 ( .A(n10621), .Z(n10620) );
  MUX U12087 ( .IN0(n9768), .IN1(data_mem_out_wire[1458]), .SEL(n10621), .F(
        n6308) );
  MUX U12088 ( .IN0(n9769), .IN1(data_mem_out_wire[1457]), .SEL(n10621), .F(
        n6307) );
  MUX U12089 ( .IN0(n9770), .IN1(data_mem_out_wire[1456]), .SEL(n10621), .F(
        n6306) );
  AND U12090 ( .A(n10622), .B(n10623), .Z(n10621) );
  OR U12091 ( .A(n9773), .B(n10619), .Z(n10623) );
  AND U12092 ( .A(n10617), .B(n10616), .Z(n10622) );
  NANDN U12093 ( .A(n10619), .B(n9809), .Z(n10617) );
  MUX U12094 ( .IN0(data_mem_out_wire[1455]), .IN1(n9776), .SEL(n10624), .F(
        n6305) );
  MUX U12095 ( .IN0(data_mem_out_wire[1454]), .IN1(n9778), .SEL(n10624), .F(
        n6304) );
  MUX U12096 ( .IN0(data_mem_out_wire[1453]), .IN1(n9779), .SEL(n10624), .F(
        n6303) );
  MUX U12097 ( .IN0(data_mem_out_wire[1452]), .IN1(n9780), .SEL(n10624), .F(
        n6302) );
  MUX U12098 ( .IN0(data_mem_out_wire[1451]), .IN1(n9781), .SEL(n10624), .F(
        n6301) );
  IV U12099 ( .A(n10625), .Z(n10624) );
  MUX U12100 ( .IN0(n9783), .IN1(data_mem_out_wire[1450]), .SEL(n10625), .F(
        n6300) );
  MUX U12101 ( .IN0(n9784), .IN1(data_mem_out_wire[1449]), .SEL(n10625), .F(
        n6299) );
  MUX U12102 ( .IN0(n9785), .IN1(data_mem_out_wire[1448]), .SEL(n10625), .F(
        n6298) );
  AND U12103 ( .A(n10626), .B(n10627), .Z(n10625) );
  OR U12104 ( .A(n9788), .B(n10619), .Z(n10627) );
  MUX U12105 ( .IN0(data_mem_out_wire[1447]), .IN1(data_in[7]), .SEL(n10628), 
        .F(n6297) );
  MUX U12106 ( .IN0(data_mem_out_wire[1446]), .IN1(data_in[6]), .SEL(n10628), 
        .F(n6296) );
  MUX U12107 ( .IN0(data_mem_out_wire[1445]), .IN1(data_in[5]), .SEL(n10628), 
        .F(n6295) );
  MUX U12108 ( .IN0(data_mem_out_wire[1444]), .IN1(data_in[4]), .SEL(n10628), 
        .F(n6294) );
  MUX U12109 ( .IN0(data_mem_out_wire[1443]), .IN1(data_in[3]), .SEL(n10628), 
        .F(n6293) );
  IV U12110 ( .A(n10629), .Z(n10628) );
  MUX U12111 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1442]), .SEL(n10629), 
        .F(n6292) );
  MUX U12112 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1441]), .SEL(n10629), 
        .F(n6291) );
  MUX U12113 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1440]), .SEL(n10629), 
        .F(n6290) );
  AND U12114 ( .A(n10626), .B(n10630), .Z(n10629) );
  NANDN U12115 ( .A(n10619), .B(n9792), .Z(n10630) );
  AND U12116 ( .A(n10631), .B(n10616), .Z(n10626) );
  NANDN U12117 ( .A(n10619), .B(n9796), .Z(n10616) );
  NANDN U12118 ( .A(n10619), .B(n9818), .Z(n10631) );
  NAND U12119 ( .A(n9900), .B(n10541), .Z(n10619) );
  MUX U12120 ( .IN0(n9746), .IN1(data_mem_out_wire[1503]), .SEL(n10632), .F(
        n6289) );
  MUX U12121 ( .IN0(n9748), .IN1(data_mem_out_wire[1502]), .SEL(n10632), .F(
        n6288) );
  MUX U12122 ( .IN0(n9749), .IN1(data_mem_out_wire[1501]), .SEL(n10632), .F(
        n6287) );
  MUX U12123 ( .IN0(n9750), .IN1(data_mem_out_wire[1500]), .SEL(n10632), .F(
        n6286) );
  MUX U12124 ( .IN0(n9751), .IN1(data_mem_out_wire[1499]), .SEL(n10632), .F(
        n6285) );
  MUX U12125 ( .IN0(n9752), .IN1(data_mem_out_wire[1498]), .SEL(n10632), .F(
        n6284) );
  MUX U12126 ( .IN0(n9753), .IN1(data_mem_out_wire[1497]), .SEL(n10632), .F(
        n6283) );
  MUX U12127 ( .IN0(n9754), .IN1(data_mem_out_wire[1496]), .SEL(n10632), .F(
        n6282) );
  AND U12128 ( .A(n10633), .B(n10634), .Z(n10632) );
  AND U12129 ( .A(n10635), .B(n10636), .Z(n10633) );
  OR U12130 ( .A(n9760), .B(n10637), .Z(n10636) );
  MUX U12131 ( .IN0(data_mem_out_wire[1495]), .IN1(n9761), .SEL(n10638), .F(
        n6281) );
  MUX U12132 ( .IN0(data_mem_out_wire[1494]), .IN1(n9763), .SEL(n10638), .F(
        n6280) );
  MUX U12133 ( .IN0(data_mem_out_wire[1493]), .IN1(n9764), .SEL(n10638), .F(
        n6279) );
  MUX U12134 ( .IN0(data_mem_out_wire[1492]), .IN1(n9765), .SEL(n10638), .F(
        n6278) );
  MUX U12135 ( .IN0(data_mem_out_wire[1491]), .IN1(n9766), .SEL(n10638), .F(
        n6277) );
  IV U12136 ( .A(n10639), .Z(n10638) );
  MUX U12137 ( .IN0(n9768), .IN1(data_mem_out_wire[1490]), .SEL(n10639), .F(
        n6276) );
  MUX U12138 ( .IN0(n9769), .IN1(data_mem_out_wire[1489]), .SEL(n10639), .F(
        n6275) );
  MUX U12139 ( .IN0(n9770), .IN1(data_mem_out_wire[1488]), .SEL(n10639), .F(
        n6274) );
  AND U12140 ( .A(n10640), .B(n10641), .Z(n10639) );
  OR U12141 ( .A(n9773), .B(n10637), .Z(n10641) );
  AND U12142 ( .A(n10635), .B(n10634), .Z(n10640) );
  NANDN U12143 ( .A(n10637), .B(n9809), .Z(n10635) );
  MUX U12144 ( .IN0(data_mem_out_wire[1487]), .IN1(n9776), .SEL(n10642), .F(
        n6273) );
  MUX U12145 ( .IN0(data_mem_out_wire[1486]), .IN1(n9778), .SEL(n10642), .F(
        n6272) );
  MUX U12146 ( .IN0(data_mem_out_wire[1485]), .IN1(n9779), .SEL(n10642), .F(
        n6271) );
  MUX U12147 ( .IN0(data_mem_out_wire[1484]), .IN1(n9780), .SEL(n10642), .F(
        n6270) );
  MUX U12148 ( .IN0(data_mem_out_wire[1483]), .IN1(n9781), .SEL(n10642), .F(
        n6269) );
  IV U12149 ( .A(n10643), .Z(n10642) );
  MUX U12150 ( .IN0(n9783), .IN1(data_mem_out_wire[1482]), .SEL(n10643), .F(
        n6268) );
  MUX U12151 ( .IN0(n9784), .IN1(data_mem_out_wire[1481]), .SEL(n10643), .F(
        n6267) );
  MUX U12152 ( .IN0(n9785), .IN1(data_mem_out_wire[1480]), .SEL(n10643), .F(
        n6266) );
  AND U12153 ( .A(n10644), .B(n10645), .Z(n10643) );
  OR U12154 ( .A(n9788), .B(n10637), .Z(n10645) );
  MUX U12155 ( .IN0(data_mem_out_wire[1479]), .IN1(data_in[7]), .SEL(n10646), 
        .F(n6265) );
  MUX U12156 ( .IN0(data_mem_out_wire[1478]), .IN1(data_in[6]), .SEL(n10646), 
        .F(n6264) );
  MUX U12157 ( .IN0(data_mem_out_wire[1477]), .IN1(data_in[5]), .SEL(n10646), 
        .F(n6263) );
  MUX U12158 ( .IN0(data_mem_out_wire[1476]), .IN1(data_in[4]), .SEL(n10646), 
        .F(n6262) );
  MUX U12159 ( .IN0(data_mem_out_wire[1475]), .IN1(data_in[3]), .SEL(n10646), 
        .F(n6261) );
  IV U12160 ( .A(n10647), .Z(n10646) );
  MUX U12161 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1474]), .SEL(n10647), 
        .F(n6260) );
  MUX U12162 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1473]), .SEL(n10647), 
        .F(n6259) );
  MUX U12163 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1472]), .SEL(n10647), 
        .F(n6258) );
  AND U12164 ( .A(n10644), .B(n10648), .Z(n10647) );
  NANDN U12165 ( .A(n10637), .B(n9792), .Z(n10648) );
  AND U12166 ( .A(n10649), .B(n10634), .Z(n10644) );
  NANDN U12167 ( .A(n10637), .B(n9796), .Z(n10634) );
  NANDN U12168 ( .A(n10637), .B(n9818), .Z(n10649) );
  NAND U12169 ( .A(n9919), .B(n10541), .Z(n10637) );
  MUX U12170 ( .IN0(n9746), .IN1(data_mem_out_wire[1535]), .SEL(n10650), .F(
        n6257) );
  MUX U12171 ( .IN0(n9748), .IN1(data_mem_out_wire[1534]), .SEL(n10650), .F(
        n6256) );
  MUX U12172 ( .IN0(n9749), .IN1(data_mem_out_wire[1533]), .SEL(n10650), .F(
        n6255) );
  MUX U12173 ( .IN0(n9750), .IN1(data_mem_out_wire[1532]), .SEL(n10650), .F(
        n6254) );
  MUX U12174 ( .IN0(n9751), .IN1(data_mem_out_wire[1531]), .SEL(n10650), .F(
        n6253) );
  MUX U12175 ( .IN0(n9752), .IN1(data_mem_out_wire[1530]), .SEL(n10650), .F(
        n6252) );
  MUX U12176 ( .IN0(n9753), .IN1(data_mem_out_wire[1529]), .SEL(n10650), .F(
        n6251) );
  MUX U12177 ( .IN0(n9754), .IN1(data_mem_out_wire[1528]), .SEL(n10650), .F(
        n6250) );
  AND U12178 ( .A(n10651), .B(n10652), .Z(n10650) );
  AND U12179 ( .A(n10653), .B(n10654), .Z(n10651) );
  OR U12180 ( .A(n9760), .B(n10655), .Z(n10654) );
  MUX U12181 ( .IN0(data_mem_out_wire[1527]), .IN1(n9761), .SEL(n10656), .F(
        n6249) );
  MUX U12182 ( .IN0(data_mem_out_wire[1526]), .IN1(n9763), .SEL(n10656), .F(
        n6248) );
  MUX U12183 ( .IN0(data_mem_out_wire[1525]), .IN1(n9764), .SEL(n10656), .F(
        n6247) );
  MUX U12184 ( .IN0(data_mem_out_wire[1524]), .IN1(n9765), .SEL(n10656), .F(
        n6246) );
  MUX U12185 ( .IN0(data_mem_out_wire[1523]), .IN1(n9766), .SEL(n10656), .F(
        n6245) );
  IV U12186 ( .A(n10657), .Z(n10656) );
  MUX U12187 ( .IN0(n9768), .IN1(data_mem_out_wire[1522]), .SEL(n10657), .F(
        n6244) );
  MUX U12188 ( .IN0(n9769), .IN1(data_mem_out_wire[1521]), .SEL(n10657), .F(
        n6243) );
  MUX U12189 ( .IN0(n9770), .IN1(data_mem_out_wire[1520]), .SEL(n10657), .F(
        n6242) );
  AND U12190 ( .A(n10658), .B(n10659), .Z(n10657) );
  OR U12191 ( .A(n9773), .B(n10655), .Z(n10659) );
  AND U12192 ( .A(n10653), .B(n10652), .Z(n10658) );
  NANDN U12193 ( .A(n10655), .B(n9809), .Z(n10653) );
  MUX U12194 ( .IN0(data_mem_out_wire[1519]), .IN1(n9776), .SEL(n10660), .F(
        n6241) );
  MUX U12195 ( .IN0(data_mem_out_wire[1518]), .IN1(n9778), .SEL(n10660), .F(
        n6240) );
  MUX U12196 ( .IN0(data_mem_out_wire[1517]), .IN1(n9779), .SEL(n10660), .F(
        n6239) );
  MUX U12197 ( .IN0(data_mem_out_wire[1516]), .IN1(n9780), .SEL(n10660), .F(
        n6238) );
  MUX U12198 ( .IN0(data_mem_out_wire[1515]), .IN1(n9781), .SEL(n10660), .F(
        n6237) );
  IV U12199 ( .A(n10661), .Z(n10660) );
  MUX U12200 ( .IN0(n9783), .IN1(data_mem_out_wire[1514]), .SEL(n10661), .F(
        n6236) );
  MUX U12201 ( .IN0(n9784), .IN1(data_mem_out_wire[1513]), .SEL(n10661), .F(
        n6235) );
  MUX U12202 ( .IN0(n9785), .IN1(data_mem_out_wire[1512]), .SEL(n10661), .F(
        n6234) );
  AND U12203 ( .A(n10662), .B(n10663), .Z(n10661) );
  OR U12204 ( .A(n9788), .B(n10655), .Z(n10663) );
  MUX U12205 ( .IN0(data_mem_out_wire[1511]), .IN1(data_in[7]), .SEL(n10664), 
        .F(n6233) );
  MUX U12206 ( .IN0(data_mem_out_wire[1510]), .IN1(data_in[6]), .SEL(n10664), 
        .F(n6232) );
  MUX U12207 ( .IN0(data_mem_out_wire[1509]), .IN1(data_in[5]), .SEL(n10664), 
        .F(n6231) );
  MUX U12208 ( .IN0(data_mem_out_wire[1508]), .IN1(data_in[4]), .SEL(n10664), 
        .F(n6230) );
  MUX U12209 ( .IN0(data_mem_out_wire[1507]), .IN1(data_in[3]), .SEL(n10664), 
        .F(n6229) );
  IV U12210 ( .A(n10665), .Z(n10664) );
  MUX U12211 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1506]), .SEL(n10665), 
        .F(n6228) );
  MUX U12212 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1505]), .SEL(n10665), 
        .F(n6227) );
  MUX U12213 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1504]), .SEL(n10665), 
        .F(n6226) );
  AND U12214 ( .A(n10662), .B(n10666), .Z(n10665) );
  NANDN U12215 ( .A(n10655), .B(n9792), .Z(n10666) );
  AND U12216 ( .A(n10667), .B(n10652), .Z(n10662) );
  NANDN U12217 ( .A(n10655), .B(n9796), .Z(n10652) );
  NANDN U12218 ( .A(n10655), .B(n9818), .Z(n10667) );
  NAND U12219 ( .A(n10541), .B(n9938), .Z(n10655) );
  AND U12220 ( .A(n10085), .B(N42), .Z(n10541) );
  AND U12221 ( .A(N40), .B(n10668), .Z(n10085) );
  MUX U12222 ( .IN0(n9746), .IN1(data_mem_out_wire[1567]), .SEL(n10669), .F(
        n6225) );
  MUX U12223 ( .IN0(n9748), .IN1(data_mem_out_wire[1566]), .SEL(n10669), .F(
        n6224) );
  MUX U12224 ( .IN0(n9749), .IN1(data_mem_out_wire[1565]), .SEL(n10669), .F(
        n6223) );
  MUX U12225 ( .IN0(n9750), .IN1(data_mem_out_wire[1564]), .SEL(n10669), .F(
        n6222) );
  MUX U12226 ( .IN0(n9751), .IN1(data_mem_out_wire[1563]), .SEL(n10669), .F(
        n6221) );
  MUX U12227 ( .IN0(n9752), .IN1(data_mem_out_wire[1562]), .SEL(n10669), .F(
        n6220) );
  MUX U12228 ( .IN0(n9753), .IN1(data_mem_out_wire[1561]), .SEL(n10669), .F(
        n6219) );
  MUX U12229 ( .IN0(n9754), .IN1(data_mem_out_wire[1560]), .SEL(n10669), .F(
        n6218) );
  AND U12230 ( .A(n10670), .B(n10671), .Z(n10669) );
  AND U12231 ( .A(n10672), .B(n10673), .Z(n10670) );
  OR U12232 ( .A(n9760), .B(n10674), .Z(n10673) );
  MUX U12233 ( .IN0(data_mem_out_wire[1559]), .IN1(n9761), .SEL(n10675), .F(
        n6217) );
  MUX U12234 ( .IN0(data_mem_out_wire[1558]), .IN1(n9763), .SEL(n10675), .F(
        n6216) );
  MUX U12235 ( .IN0(data_mem_out_wire[1557]), .IN1(n9764), .SEL(n10675), .F(
        n6215) );
  MUX U12236 ( .IN0(data_mem_out_wire[1556]), .IN1(n9765), .SEL(n10675), .F(
        n6214) );
  MUX U12237 ( .IN0(data_mem_out_wire[1555]), .IN1(n9766), .SEL(n10675), .F(
        n6213) );
  IV U12238 ( .A(n10676), .Z(n10675) );
  MUX U12239 ( .IN0(n9768), .IN1(data_mem_out_wire[1554]), .SEL(n10676), .F(
        n6212) );
  MUX U12240 ( .IN0(n9769), .IN1(data_mem_out_wire[1553]), .SEL(n10676), .F(
        n6211) );
  MUX U12241 ( .IN0(n9770), .IN1(data_mem_out_wire[1552]), .SEL(n10676), .F(
        n6210) );
  AND U12242 ( .A(n10677), .B(n10678), .Z(n10676) );
  OR U12243 ( .A(n9773), .B(n10674), .Z(n10678) );
  AND U12244 ( .A(n10672), .B(n10671), .Z(n10677) );
  NANDN U12245 ( .A(n10674), .B(n9809), .Z(n10672) );
  MUX U12246 ( .IN0(data_mem_out_wire[1551]), .IN1(n9776), .SEL(n10679), .F(
        n6209) );
  MUX U12247 ( .IN0(data_mem_out_wire[1550]), .IN1(n9778), .SEL(n10679), .F(
        n6208) );
  MUX U12248 ( .IN0(data_mem_out_wire[1549]), .IN1(n9779), .SEL(n10679), .F(
        n6207) );
  MUX U12249 ( .IN0(data_mem_out_wire[1548]), .IN1(n9780), .SEL(n10679), .F(
        n6206) );
  MUX U12250 ( .IN0(data_mem_out_wire[1547]), .IN1(n9781), .SEL(n10679), .F(
        n6205) );
  IV U12251 ( .A(n10680), .Z(n10679) );
  MUX U12252 ( .IN0(n9783), .IN1(data_mem_out_wire[1546]), .SEL(n10680), .F(
        n6204) );
  MUX U12253 ( .IN0(n9784), .IN1(data_mem_out_wire[1545]), .SEL(n10680), .F(
        n6203) );
  MUX U12254 ( .IN0(n9785), .IN1(data_mem_out_wire[1544]), .SEL(n10680), .F(
        n6202) );
  AND U12255 ( .A(n10681), .B(n10682), .Z(n10680) );
  OR U12256 ( .A(n9788), .B(n10674), .Z(n10682) );
  MUX U12257 ( .IN0(data_mem_out_wire[1543]), .IN1(data_in[7]), .SEL(n10683), 
        .F(n6201) );
  MUX U12258 ( .IN0(data_mem_out_wire[1542]), .IN1(data_in[6]), .SEL(n10683), 
        .F(n6200) );
  MUX U12259 ( .IN0(data_mem_out_wire[1541]), .IN1(data_in[5]), .SEL(n10683), 
        .F(n6199) );
  MUX U12260 ( .IN0(data_mem_out_wire[1540]), .IN1(data_in[4]), .SEL(n10683), 
        .F(n6198) );
  MUX U12261 ( .IN0(data_mem_out_wire[1539]), .IN1(data_in[3]), .SEL(n10683), 
        .F(n6197) );
  IV U12262 ( .A(n10684), .Z(n10683) );
  MUX U12263 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1538]), .SEL(n10684), 
        .F(n6196) );
  MUX U12264 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1537]), .SEL(n10684), 
        .F(n6195) );
  MUX U12265 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1536]), .SEL(n10684), 
        .F(n6194) );
  AND U12266 ( .A(n10681), .B(n10685), .Z(n10684) );
  NANDN U12267 ( .A(n10674), .B(n9792), .Z(n10685) );
  AND U12268 ( .A(n10686), .B(n10671), .Z(n10681) );
  NANDN U12269 ( .A(n10674), .B(n9796), .Z(n10671) );
  NANDN U12270 ( .A(n10674), .B(n9818), .Z(n10686) );
  NAND U12271 ( .A(n9798), .B(n10687), .Z(n10674) );
  MUX U12272 ( .IN0(n9746), .IN1(data_mem_out_wire[1599]), .SEL(n10688), .F(
        n6193) );
  MUX U12273 ( .IN0(n9748), .IN1(data_mem_out_wire[1598]), .SEL(n10688), .F(
        n6192) );
  MUX U12274 ( .IN0(n9749), .IN1(data_mem_out_wire[1597]), .SEL(n10688), .F(
        n6191) );
  MUX U12275 ( .IN0(n9750), .IN1(data_mem_out_wire[1596]), .SEL(n10688), .F(
        n6190) );
  MUX U12276 ( .IN0(n9751), .IN1(data_mem_out_wire[1595]), .SEL(n10688), .F(
        n6189) );
  MUX U12277 ( .IN0(n9752), .IN1(data_mem_out_wire[1594]), .SEL(n10688), .F(
        n6188) );
  MUX U12278 ( .IN0(n9753), .IN1(data_mem_out_wire[1593]), .SEL(n10688), .F(
        n6187) );
  MUX U12279 ( .IN0(n9754), .IN1(data_mem_out_wire[1592]), .SEL(n10688), .F(
        n6186) );
  AND U12280 ( .A(n10689), .B(n10690), .Z(n10688) );
  AND U12281 ( .A(n10691), .B(n10692), .Z(n10689) );
  OR U12282 ( .A(n9760), .B(n10693), .Z(n10692) );
  MUX U12283 ( .IN0(data_mem_out_wire[1591]), .IN1(n9761), .SEL(n10694), .F(
        n6185) );
  MUX U12284 ( .IN0(data_mem_out_wire[1590]), .IN1(n9763), .SEL(n10694), .F(
        n6184) );
  MUX U12285 ( .IN0(data_mem_out_wire[1589]), .IN1(n9764), .SEL(n10694), .F(
        n6183) );
  MUX U12286 ( .IN0(data_mem_out_wire[1588]), .IN1(n9765), .SEL(n10694), .F(
        n6182) );
  MUX U12287 ( .IN0(data_mem_out_wire[1587]), .IN1(n9766), .SEL(n10694), .F(
        n6181) );
  IV U12288 ( .A(n10695), .Z(n10694) );
  MUX U12289 ( .IN0(n9768), .IN1(data_mem_out_wire[1586]), .SEL(n10695), .F(
        n6180) );
  MUX U12290 ( .IN0(n9769), .IN1(data_mem_out_wire[1585]), .SEL(n10695), .F(
        n6179) );
  MUX U12291 ( .IN0(n9770), .IN1(data_mem_out_wire[1584]), .SEL(n10695), .F(
        n6178) );
  AND U12292 ( .A(n10696), .B(n10697), .Z(n10695) );
  OR U12293 ( .A(n9773), .B(n10693), .Z(n10697) );
  AND U12294 ( .A(n10691), .B(n10690), .Z(n10696) );
  NANDN U12295 ( .A(n10693), .B(n9809), .Z(n10691) );
  MUX U12296 ( .IN0(data_mem_out_wire[1583]), .IN1(n9776), .SEL(n10698), .F(
        n6177) );
  MUX U12297 ( .IN0(data_mem_out_wire[1582]), .IN1(n9778), .SEL(n10698), .F(
        n6176) );
  MUX U12298 ( .IN0(data_mem_out_wire[1581]), .IN1(n9779), .SEL(n10698), .F(
        n6175) );
  MUX U12299 ( .IN0(data_mem_out_wire[1580]), .IN1(n9780), .SEL(n10698), .F(
        n6174) );
  MUX U12300 ( .IN0(data_mem_out_wire[1579]), .IN1(n9781), .SEL(n10698), .F(
        n6173) );
  IV U12301 ( .A(n10699), .Z(n10698) );
  MUX U12302 ( .IN0(n9783), .IN1(data_mem_out_wire[1578]), .SEL(n10699), .F(
        n6172) );
  MUX U12303 ( .IN0(n9784), .IN1(data_mem_out_wire[1577]), .SEL(n10699), .F(
        n6171) );
  MUX U12304 ( .IN0(n9785), .IN1(data_mem_out_wire[1576]), .SEL(n10699), .F(
        n6170) );
  AND U12305 ( .A(n10700), .B(n10701), .Z(n10699) );
  OR U12306 ( .A(n9788), .B(n10693), .Z(n10701) );
  MUX U12307 ( .IN0(data_mem_out_wire[1575]), .IN1(data_in[7]), .SEL(n10702), 
        .F(n6169) );
  MUX U12308 ( .IN0(data_mem_out_wire[1574]), .IN1(data_in[6]), .SEL(n10702), 
        .F(n6168) );
  MUX U12309 ( .IN0(data_mem_out_wire[1573]), .IN1(data_in[5]), .SEL(n10702), 
        .F(n6167) );
  MUX U12310 ( .IN0(data_mem_out_wire[1572]), .IN1(data_in[4]), .SEL(n10702), 
        .F(n6166) );
  MUX U12311 ( .IN0(data_mem_out_wire[1571]), .IN1(data_in[3]), .SEL(n10702), 
        .F(n6165) );
  IV U12312 ( .A(n10703), .Z(n10702) );
  MUX U12313 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1570]), .SEL(n10703), 
        .F(n6164) );
  MUX U12314 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1569]), .SEL(n10703), 
        .F(n6163) );
  MUX U12315 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1568]), .SEL(n10703), 
        .F(n6162) );
  AND U12316 ( .A(n10700), .B(n10704), .Z(n10703) );
  NANDN U12317 ( .A(n10693), .B(n9792), .Z(n10704) );
  AND U12318 ( .A(n10705), .B(n10690), .Z(n10700) );
  NANDN U12319 ( .A(n10693), .B(n9796), .Z(n10690) );
  NANDN U12320 ( .A(n10693), .B(n9818), .Z(n10705) );
  NAND U12321 ( .A(n9819), .B(n10687), .Z(n10693) );
  MUX U12322 ( .IN0(n9746), .IN1(data_mem_out_wire[1631]), .SEL(n10706), .F(
        n6161) );
  MUX U12323 ( .IN0(n9748), .IN1(data_mem_out_wire[1630]), .SEL(n10706), .F(
        n6160) );
  MUX U12324 ( .IN0(n9749), .IN1(data_mem_out_wire[1629]), .SEL(n10706), .F(
        n6159) );
  MUX U12325 ( .IN0(n9750), .IN1(data_mem_out_wire[1628]), .SEL(n10706), .F(
        n6158) );
  MUX U12326 ( .IN0(n9751), .IN1(data_mem_out_wire[1627]), .SEL(n10706), .F(
        n6157) );
  MUX U12327 ( .IN0(n9752), .IN1(data_mem_out_wire[1626]), .SEL(n10706), .F(
        n6156) );
  MUX U12328 ( .IN0(n9753), .IN1(data_mem_out_wire[1625]), .SEL(n10706), .F(
        n6155) );
  MUX U12329 ( .IN0(n9754), .IN1(data_mem_out_wire[1624]), .SEL(n10706), .F(
        n6154) );
  AND U12330 ( .A(n10707), .B(n10708), .Z(n10706) );
  AND U12331 ( .A(n10709), .B(n10710), .Z(n10707) );
  OR U12332 ( .A(n9760), .B(n10711), .Z(n10710) );
  MUX U12333 ( .IN0(data_mem_out_wire[1623]), .IN1(n9761), .SEL(n10712), .F(
        n6153) );
  MUX U12334 ( .IN0(data_mem_out_wire[1622]), .IN1(n9763), .SEL(n10712), .F(
        n6152) );
  MUX U12335 ( .IN0(data_mem_out_wire[1621]), .IN1(n9764), .SEL(n10712), .F(
        n6151) );
  MUX U12336 ( .IN0(data_mem_out_wire[1620]), .IN1(n9765), .SEL(n10712), .F(
        n6150) );
  MUX U12337 ( .IN0(data_mem_out_wire[1619]), .IN1(n9766), .SEL(n10712), .F(
        n6149) );
  IV U12338 ( .A(n10713), .Z(n10712) );
  MUX U12339 ( .IN0(n9768), .IN1(data_mem_out_wire[1618]), .SEL(n10713), .F(
        n6148) );
  MUX U12340 ( .IN0(n9769), .IN1(data_mem_out_wire[1617]), .SEL(n10713), .F(
        n6147) );
  MUX U12341 ( .IN0(n9770), .IN1(data_mem_out_wire[1616]), .SEL(n10713), .F(
        n6146) );
  AND U12342 ( .A(n10714), .B(n10715), .Z(n10713) );
  OR U12343 ( .A(n9773), .B(n10711), .Z(n10715) );
  AND U12344 ( .A(n10709), .B(n10708), .Z(n10714) );
  NANDN U12345 ( .A(n10711), .B(n9809), .Z(n10709) );
  MUX U12346 ( .IN0(data_mem_out_wire[1615]), .IN1(n9776), .SEL(n10716), .F(
        n6145) );
  MUX U12347 ( .IN0(data_mem_out_wire[1614]), .IN1(n9778), .SEL(n10716), .F(
        n6144) );
  MUX U12348 ( .IN0(data_mem_out_wire[1613]), .IN1(n9779), .SEL(n10716), .F(
        n6143) );
  MUX U12349 ( .IN0(data_mem_out_wire[1612]), .IN1(n9780), .SEL(n10716), .F(
        n6142) );
  MUX U12350 ( .IN0(data_mem_out_wire[1611]), .IN1(n9781), .SEL(n10716), .F(
        n6141) );
  IV U12351 ( .A(n10717), .Z(n10716) );
  MUX U12352 ( .IN0(n9783), .IN1(data_mem_out_wire[1610]), .SEL(n10717), .F(
        n6140) );
  MUX U12353 ( .IN0(n9784), .IN1(data_mem_out_wire[1609]), .SEL(n10717), .F(
        n6139) );
  MUX U12354 ( .IN0(n9785), .IN1(data_mem_out_wire[1608]), .SEL(n10717), .F(
        n6138) );
  AND U12355 ( .A(n10718), .B(n10719), .Z(n10717) );
  OR U12356 ( .A(n9788), .B(n10711), .Z(n10719) );
  MUX U12357 ( .IN0(data_mem_out_wire[1607]), .IN1(data_in[7]), .SEL(n10720), 
        .F(n6137) );
  MUX U12358 ( .IN0(data_mem_out_wire[1606]), .IN1(data_in[6]), .SEL(n10720), 
        .F(n6136) );
  MUX U12359 ( .IN0(data_mem_out_wire[1605]), .IN1(data_in[5]), .SEL(n10720), 
        .F(n6135) );
  MUX U12360 ( .IN0(data_mem_out_wire[1604]), .IN1(data_in[4]), .SEL(n10720), 
        .F(n6134) );
  MUX U12361 ( .IN0(data_mem_out_wire[1603]), .IN1(data_in[3]), .SEL(n10720), 
        .F(n6133) );
  IV U12362 ( .A(n10721), .Z(n10720) );
  MUX U12363 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1602]), .SEL(n10721), 
        .F(n6132) );
  MUX U12364 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1601]), .SEL(n10721), 
        .F(n6131) );
  MUX U12365 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1600]), .SEL(n10721), 
        .F(n6130) );
  AND U12366 ( .A(n10718), .B(n10722), .Z(n10721) );
  NANDN U12367 ( .A(n10711), .B(n9792), .Z(n10722) );
  AND U12368 ( .A(n10723), .B(n10708), .Z(n10718) );
  NANDN U12369 ( .A(n10711), .B(n9796), .Z(n10708) );
  NANDN U12370 ( .A(n10711), .B(n9818), .Z(n10723) );
  NAND U12371 ( .A(n9838), .B(n10687), .Z(n10711) );
  MUX U12372 ( .IN0(n9746), .IN1(data_mem_out_wire[1663]), .SEL(n10724), .F(
        n6129) );
  MUX U12373 ( .IN0(n9748), .IN1(data_mem_out_wire[1662]), .SEL(n10724), .F(
        n6128) );
  MUX U12374 ( .IN0(n9749), .IN1(data_mem_out_wire[1661]), .SEL(n10724), .F(
        n6127) );
  MUX U12375 ( .IN0(n9750), .IN1(data_mem_out_wire[1660]), .SEL(n10724), .F(
        n6126) );
  MUX U12376 ( .IN0(n9751), .IN1(data_mem_out_wire[1659]), .SEL(n10724), .F(
        n6125) );
  MUX U12377 ( .IN0(n9752), .IN1(data_mem_out_wire[1658]), .SEL(n10724), .F(
        n6124) );
  MUX U12378 ( .IN0(n9753), .IN1(data_mem_out_wire[1657]), .SEL(n10724), .F(
        n6123) );
  MUX U12379 ( .IN0(n9754), .IN1(data_mem_out_wire[1656]), .SEL(n10724), .F(
        n6122) );
  AND U12380 ( .A(n10725), .B(n10726), .Z(n10724) );
  AND U12381 ( .A(n10727), .B(n10728), .Z(n10725) );
  OR U12382 ( .A(n9760), .B(n10729), .Z(n10728) );
  MUX U12383 ( .IN0(data_mem_out_wire[1655]), .IN1(n9761), .SEL(n10730), .F(
        n6121) );
  MUX U12384 ( .IN0(data_mem_out_wire[1654]), .IN1(n9763), .SEL(n10730), .F(
        n6120) );
  MUX U12385 ( .IN0(data_mem_out_wire[1653]), .IN1(n9764), .SEL(n10730), .F(
        n6119) );
  MUX U12386 ( .IN0(data_mem_out_wire[1652]), .IN1(n9765), .SEL(n10730), .F(
        n6118) );
  MUX U12387 ( .IN0(data_mem_out_wire[1651]), .IN1(n9766), .SEL(n10730), .F(
        n6117) );
  IV U12388 ( .A(n10731), .Z(n10730) );
  MUX U12389 ( .IN0(n9768), .IN1(data_mem_out_wire[1650]), .SEL(n10731), .F(
        n6116) );
  MUX U12390 ( .IN0(n9769), .IN1(data_mem_out_wire[1649]), .SEL(n10731), .F(
        n6115) );
  MUX U12391 ( .IN0(n9770), .IN1(data_mem_out_wire[1648]), .SEL(n10731), .F(
        n6114) );
  AND U12392 ( .A(n10732), .B(n10733), .Z(n10731) );
  OR U12393 ( .A(n9773), .B(n10729), .Z(n10733) );
  AND U12394 ( .A(n10727), .B(n10726), .Z(n10732) );
  NANDN U12395 ( .A(n10729), .B(n9809), .Z(n10727) );
  MUX U12396 ( .IN0(data_mem_out_wire[1647]), .IN1(n9776), .SEL(n10734), .F(
        n6113) );
  MUX U12397 ( .IN0(data_mem_out_wire[1646]), .IN1(n9778), .SEL(n10734), .F(
        n6112) );
  MUX U12398 ( .IN0(data_mem_out_wire[1645]), .IN1(n9779), .SEL(n10734), .F(
        n6111) );
  MUX U12399 ( .IN0(data_mem_out_wire[1644]), .IN1(n9780), .SEL(n10734), .F(
        n6110) );
  MUX U12400 ( .IN0(data_mem_out_wire[1643]), .IN1(n9781), .SEL(n10734), .F(
        n6109) );
  IV U12401 ( .A(n10735), .Z(n10734) );
  MUX U12402 ( .IN0(n9783), .IN1(data_mem_out_wire[1642]), .SEL(n10735), .F(
        n6108) );
  MUX U12403 ( .IN0(n9784), .IN1(data_mem_out_wire[1641]), .SEL(n10735), .F(
        n6107) );
  MUX U12404 ( .IN0(n9785), .IN1(data_mem_out_wire[1640]), .SEL(n10735), .F(
        n6106) );
  AND U12405 ( .A(n10736), .B(n10737), .Z(n10735) );
  OR U12406 ( .A(n9788), .B(n10729), .Z(n10737) );
  MUX U12407 ( .IN0(data_mem_out_wire[1639]), .IN1(data_in[7]), .SEL(n10738), 
        .F(n6105) );
  MUX U12408 ( .IN0(data_mem_out_wire[1638]), .IN1(data_in[6]), .SEL(n10738), 
        .F(n6104) );
  MUX U12409 ( .IN0(data_mem_out_wire[1637]), .IN1(data_in[5]), .SEL(n10738), 
        .F(n6103) );
  MUX U12410 ( .IN0(data_mem_out_wire[1636]), .IN1(data_in[4]), .SEL(n10738), 
        .F(n6102) );
  MUX U12411 ( .IN0(data_mem_out_wire[1635]), .IN1(data_in[3]), .SEL(n10738), 
        .F(n6101) );
  IV U12412 ( .A(n10739), .Z(n10738) );
  MUX U12413 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1634]), .SEL(n10739), 
        .F(n6100) );
  MUX U12414 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1633]), .SEL(n10739), 
        .F(n6099) );
  MUX U12415 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1632]), .SEL(n10739), 
        .F(n6098) );
  AND U12416 ( .A(n10736), .B(n10740), .Z(n10739) );
  NANDN U12417 ( .A(n10729), .B(n9792), .Z(n10740) );
  AND U12418 ( .A(n10741), .B(n10726), .Z(n10736) );
  NANDN U12419 ( .A(n10729), .B(n9796), .Z(n10726) );
  NANDN U12420 ( .A(n10729), .B(n9818), .Z(n10741) );
  NAND U12421 ( .A(n9862), .B(n10687), .Z(n10729) );
  MUX U12422 ( .IN0(n9746), .IN1(data_mem_out_wire[1695]), .SEL(n10742), .F(
        n6097) );
  MUX U12423 ( .IN0(n9748), .IN1(data_mem_out_wire[1694]), .SEL(n10742), .F(
        n6096) );
  MUX U12424 ( .IN0(n9749), .IN1(data_mem_out_wire[1693]), .SEL(n10742), .F(
        n6095) );
  MUX U12425 ( .IN0(n9750), .IN1(data_mem_out_wire[1692]), .SEL(n10742), .F(
        n6094) );
  MUX U12426 ( .IN0(n9751), .IN1(data_mem_out_wire[1691]), .SEL(n10742), .F(
        n6093) );
  MUX U12427 ( .IN0(n9752), .IN1(data_mem_out_wire[1690]), .SEL(n10742), .F(
        n6092) );
  MUX U12428 ( .IN0(n9753), .IN1(data_mem_out_wire[1689]), .SEL(n10742), .F(
        n6091) );
  MUX U12429 ( .IN0(n9754), .IN1(data_mem_out_wire[1688]), .SEL(n10742), .F(
        n6090) );
  AND U12430 ( .A(n10743), .B(n10744), .Z(n10742) );
  AND U12431 ( .A(n10745), .B(n10746), .Z(n10743) );
  OR U12432 ( .A(n9760), .B(n10747), .Z(n10746) );
  MUX U12433 ( .IN0(data_mem_out_wire[1687]), .IN1(n9761), .SEL(n10748), .F(
        n6089) );
  MUX U12434 ( .IN0(data_mem_out_wire[1686]), .IN1(n9763), .SEL(n10748), .F(
        n6088) );
  MUX U12435 ( .IN0(data_mem_out_wire[1685]), .IN1(n9764), .SEL(n10748), .F(
        n6087) );
  MUX U12436 ( .IN0(data_mem_out_wire[1684]), .IN1(n9765), .SEL(n10748), .F(
        n6086) );
  MUX U12437 ( .IN0(data_mem_out_wire[1683]), .IN1(n9766), .SEL(n10748), .F(
        n6085) );
  IV U12438 ( .A(n10749), .Z(n10748) );
  MUX U12439 ( .IN0(n9768), .IN1(data_mem_out_wire[1682]), .SEL(n10749), .F(
        n6084) );
  MUX U12440 ( .IN0(n9769), .IN1(data_mem_out_wire[1681]), .SEL(n10749), .F(
        n6083) );
  MUX U12441 ( .IN0(n9770), .IN1(data_mem_out_wire[1680]), .SEL(n10749), .F(
        n6082) );
  AND U12442 ( .A(n10750), .B(n10751), .Z(n10749) );
  OR U12443 ( .A(n9773), .B(n10747), .Z(n10751) );
  AND U12444 ( .A(n10745), .B(n10744), .Z(n10750) );
  NANDN U12445 ( .A(n10747), .B(n9809), .Z(n10745) );
  MUX U12446 ( .IN0(data_mem_out_wire[1679]), .IN1(n9776), .SEL(n10752), .F(
        n6081) );
  MUX U12447 ( .IN0(data_mem_out_wire[1678]), .IN1(n9778), .SEL(n10752), .F(
        n6080) );
  MUX U12448 ( .IN0(data_mem_out_wire[1677]), .IN1(n9779), .SEL(n10752), .F(
        n6079) );
  MUX U12449 ( .IN0(data_mem_out_wire[1676]), .IN1(n9780), .SEL(n10752), .F(
        n6078) );
  MUX U12450 ( .IN0(data_mem_out_wire[1675]), .IN1(n9781), .SEL(n10752), .F(
        n6077) );
  IV U12451 ( .A(n10753), .Z(n10752) );
  MUX U12452 ( .IN0(n9783), .IN1(data_mem_out_wire[1674]), .SEL(n10753), .F(
        n6076) );
  MUX U12453 ( .IN0(n9784), .IN1(data_mem_out_wire[1673]), .SEL(n10753), .F(
        n6075) );
  MUX U12454 ( .IN0(n9785), .IN1(data_mem_out_wire[1672]), .SEL(n10753), .F(
        n6074) );
  AND U12455 ( .A(n10754), .B(n10755), .Z(n10753) );
  OR U12456 ( .A(n9788), .B(n10747), .Z(n10755) );
  MUX U12457 ( .IN0(data_mem_out_wire[1671]), .IN1(data_in[7]), .SEL(n10756), 
        .F(n6073) );
  MUX U12458 ( .IN0(data_mem_out_wire[1670]), .IN1(data_in[6]), .SEL(n10756), 
        .F(n6072) );
  MUX U12459 ( .IN0(data_mem_out_wire[1669]), .IN1(data_in[5]), .SEL(n10756), 
        .F(n6071) );
  MUX U12460 ( .IN0(data_mem_out_wire[1668]), .IN1(data_in[4]), .SEL(n10756), 
        .F(n6070) );
  MUX U12461 ( .IN0(data_mem_out_wire[1667]), .IN1(data_in[3]), .SEL(n10756), 
        .F(n6069) );
  IV U12462 ( .A(n10757), .Z(n10756) );
  MUX U12463 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1666]), .SEL(n10757), 
        .F(n6068) );
  MUX U12464 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1665]), .SEL(n10757), 
        .F(n6067) );
  MUX U12465 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1664]), .SEL(n10757), 
        .F(n6066) );
  AND U12466 ( .A(n10754), .B(n10758), .Z(n10757) );
  NANDN U12467 ( .A(n10747), .B(n9792), .Z(n10758) );
  AND U12468 ( .A(n10759), .B(n10744), .Z(n10754) );
  NANDN U12469 ( .A(n10747), .B(n9796), .Z(n10744) );
  NANDN U12470 ( .A(n10747), .B(n9818), .Z(n10759) );
  NAND U12471 ( .A(n9881), .B(n10687), .Z(n10747) );
  MUX U12472 ( .IN0(n9746), .IN1(data_mem_out_wire[1727]), .SEL(n10760), .F(
        n6065) );
  MUX U12473 ( .IN0(n9748), .IN1(data_mem_out_wire[1726]), .SEL(n10760), .F(
        n6064) );
  MUX U12474 ( .IN0(n9749), .IN1(data_mem_out_wire[1725]), .SEL(n10760), .F(
        n6063) );
  MUX U12475 ( .IN0(n9750), .IN1(data_mem_out_wire[1724]), .SEL(n10760), .F(
        n6062) );
  MUX U12476 ( .IN0(n9751), .IN1(data_mem_out_wire[1723]), .SEL(n10760), .F(
        n6061) );
  MUX U12477 ( .IN0(n9752), .IN1(data_mem_out_wire[1722]), .SEL(n10760), .F(
        n6060) );
  MUX U12478 ( .IN0(n9753), .IN1(data_mem_out_wire[1721]), .SEL(n10760), .F(
        n6059) );
  MUX U12479 ( .IN0(n9754), .IN1(data_mem_out_wire[1720]), .SEL(n10760), .F(
        n6058) );
  AND U12480 ( .A(n10761), .B(n10762), .Z(n10760) );
  AND U12481 ( .A(n10763), .B(n10764), .Z(n10761) );
  OR U12482 ( .A(n9760), .B(n10765), .Z(n10764) );
  MUX U12483 ( .IN0(data_mem_out_wire[1719]), .IN1(n9761), .SEL(n10766), .F(
        n6057) );
  MUX U12484 ( .IN0(data_mem_out_wire[1718]), .IN1(n9763), .SEL(n10766), .F(
        n6056) );
  MUX U12485 ( .IN0(data_mem_out_wire[1717]), .IN1(n9764), .SEL(n10766), .F(
        n6055) );
  MUX U12486 ( .IN0(data_mem_out_wire[1716]), .IN1(n9765), .SEL(n10766), .F(
        n6054) );
  MUX U12487 ( .IN0(data_mem_out_wire[1715]), .IN1(n9766), .SEL(n10766), .F(
        n6053) );
  IV U12488 ( .A(n10767), .Z(n10766) );
  MUX U12489 ( .IN0(n9768), .IN1(data_mem_out_wire[1714]), .SEL(n10767), .F(
        n6052) );
  MUX U12490 ( .IN0(n9769), .IN1(data_mem_out_wire[1713]), .SEL(n10767), .F(
        n6051) );
  MUX U12491 ( .IN0(n9770), .IN1(data_mem_out_wire[1712]), .SEL(n10767), .F(
        n6050) );
  AND U12492 ( .A(n10768), .B(n10769), .Z(n10767) );
  OR U12493 ( .A(n9773), .B(n10765), .Z(n10769) );
  AND U12494 ( .A(n10763), .B(n10762), .Z(n10768) );
  NANDN U12495 ( .A(n10765), .B(n9809), .Z(n10763) );
  MUX U12496 ( .IN0(data_mem_out_wire[1711]), .IN1(n9776), .SEL(n10770), .F(
        n6049) );
  MUX U12497 ( .IN0(data_mem_out_wire[1710]), .IN1(n9778), .SEL(n10770), .F(
        n6048) );
  MUX U12498 ( .IN0(data_mem_out_wire[1709]), .IN1(n9779), .SEL(n10770), .F(
        n6047) );
  MUX U12499 ( .IN0(data_mem_out_wire[1708]), .IN1(n9780), .SEL(n10770), .F(
        n6046) );
  MUX U12500 ( .IN0(data_mem_out_wire[1707]), .IN1(n9781), .SEL(n10770), .F(
        n6045) );
  IV U12501 ( .A(n10771), .Z(n10770) );
  MUX U12502 ( .IN0(n9783), .IN1(data_mem_out_wire[1706]), .SEL(n10771), .F(
        n6044) );
  MUX U12503 ( .IN0(n9784), .IN1(data_mem_out_wire[1705]), .SEL(n10771), .F(
        n6043) );
  MUX U12504 ( .IN0(n9785), .IN1(data_mem_out_wire[1704]), .SEL(n10771), .F(
        n6042) );
  AND U12505 ( .A(n10772), .B(n10773), .Z(n10771) );
  OR U12506 ( .A(n9788), .B(n10765), .Z(n10773) );
  MUX U12507 ( .IN0(data_mem_out_wire[1703]), .IN1(data_in[7]), .SEL(n10774), 
        .F(n6041) );
  MUX U12508 ( .IN0(data_mem_out_wire[1702]), .IN1(data_in[6]), .SEL(n10774), 
        .F(n6040) );
  MUX U12509 ( .IN0(data_mem_out_wire[1701]), .IN1(data_in[5]), .SEL(n10774), 
        .F(n6039) );
  MUX U12510 ( .IN0(data_mem_out_wire[1700]), .IN1(data_in[4]), .SEL(n10774), 
        .F(n6038) );
  MUX U12511 ( .IN0(data_mem_out_wire[1699]), .IN1(data_in[3]), .SEL(n10774), 
        .F(n6037) );
  IV U12512 ( .A(n10775), .Z(n10774) );
  MUX U12513 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1698]), .SEL(n10775), 
        .F(n6036) );
  MUX U12514 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1697]), .SEL(n10775), 
        .F(n6035) );
  MUX U12515 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1696]), .SEL(n10775), 
        .F(n6034) );
  AND U12516 ( .A(n10772), .B(n10776), .Z(n10775) );
  NANDN U12517 ( .A(n10765), .B(n9792), .Z(n10776) );
  AND U12518 ( .A(n10777), .B(n10762), .Z(n10772) );
  NANDN U12519 ( .A(n10765), .B(n9796), .Z(n10762) );
  NANDN U12520 ( .A(n10765), .B(n9818), .Z(n10777) );
  NAND U12521 ( .A(n9900), .B(n10687), .Z(n10765) );
  MUX U12522 ( .IN0(n9746), .IN1(data_mem_out_wire[1759]), .SEL(n10778), .F(
        n6033) );
  MUX U12523 ( .IN0(n9748), .IN1(data_mem_out_wire[1758]), .SEL(n10778), .F(
        n6032) );
  MUX U12524 ( .IN0(n9749), .IN1(data_mem_out_wire[1757]), .SEL(n10778), .F(
        n6031) );
  MUX U12525 ( .IN0(n9750), .IN1(data_mem_out_wire[1756]), .SEL(n10778), .F(
        n6030) );
  MUX U12526 ( .IN0(n9751), .IN1(data_mem_out_wire[1755]), .SEL(n10778), .F(
        n6029) );
  MUX U12527 ( .IN0(n9752), .IN1(data_mem_out_wire[1754]), .SEL(n10778), .F(
        n6028) );
  MUX U12528 ( .IN0(n9753), .IN1(data_mem_out_wire[1753]), .SEL(n10778), .F(
        n6027) );
  MUX U12529 ( .IN0(n9754), .IN1(data_mem_out_wire[1752]), .SEL(n10778), .F(
        n6026) );
  AND U12530 ( .A(n10779), .B(n10780), .Z(n10778) );
  AND U12531 ( .A(n10781), .B(n10782), .Z(n10779) );
  OR U12532 ( .A(n9760), .B(n10783), .Z(n10782) );
  MUX U12533 ( .IN0(data_mem_out_wire[1751]), .IN1(n9761), .SEL(n10784), .F(
        n6025) );
  MUX U12534 ( .IN0(data_mem_out_wire[1750]), .IN1(n9763), .SEL(n10784), .F(
        n6024) );
  MUX U12535 ( .IN0(data_mem_out_wire[1749]), .IN1(n9764), .SEL(n10784), .F(
        n6023) );
  MUX U12536 ( .IN0(data_mem_out_wire[1748]), .IN1(n9765), .SEL(n10784), .F(
        n6022) );
  MUX U12537 ( .IN0(data_mem_out_wire[1747]), .IN1(n9766), .SEL(n10784), .F(
        n6021) );
  IV U12538 ( .A(n10785), .Z(n10784) );
  MUX U12539 ( .IN0(n9768), .IN1(data_mem_out_wire[1746]), .SEL(n10785), .F(
        n6020) );
  MUX U12540 ( .IN0(n9769), .IN1(data_mem_out_wire[1745]), .SEL(n10785), .F(
        n6019) );
  MUX U12541 ( .IN0(n9770), .IN1(data_mem_out_wire[1744]), .SEL(n10785), .F(
        n6018) );
  AND U12542 ( .A(n10786), .B(n10787), .Z(n10785) );
  OR U12543 ( .A(n9773), .B(n10783), .Z(n10787) );
  AND U12544 ( .A(n10781), .B(n10780), .Z(n10786) );
  NANDN U12545 ( .A(n10783), .B(n9809), .Z(n10781) );
  MUX U12546 ( .IN0(data_mem_out_wire[1743]), .IN1(n9776), .SEL(n10788), .F(
        n6017) );
  MUX U12547 ( .IN0(data_mem_out_wire[1742]), .IN1(n9778), .SEL(n10788), .F(
        n6016) );
  MUX U12548 ( .IN0(data_mem_out_wire[1741]), .IN1(n9779), .SEL(n10788), .F(
        n6015) );
  MUX U12549 ( .IN0(data_mem_out_wire[1740]), .IN1(n9780), .SEL(n10788), .F(
        n6014) );
  MUX U12550 ( .IN0(data_mem_out_wire[1739]), .IN1(n9781), .SEL(n10788), .F(
        n6013) );
  IV U12551 ( .A(n10789), .Z(n10788) );
  MUX U12552 ( .IN0(n9783), .IN1(data_mem_out_wire[1738]), .SEL(n10789), .F(
        n6012) );
  MUX U12553 ( .IN0(n9784), .IN1(data_mem_out_wire[1737]), .SEL(n10789), .F(
        n6011) );
  MUX U12554 ( .IN0(n9785), .IN1(data_mem_out_wire[1736]), .SEL(n10789), .F(
        n6010) );
  AND U12555 ( .A(n10790), .B(n10791), .Z(n10789) );
  OR U12556 ( .A(n9788), .B(n10783), .Z(n10791) );
  MUX U12557 ( .IN0(data_mem_out_wire[1735]), .IN1(data_in[7]), .SEL(n10792), 
        .F(n6009) );
  MUX U12558 ( .IN0(data_mem_out_wire[1734]), .IN1(data_in[6]), .SEL(n10792), 
        .F(n6008) );
  MUX U12559 ( .IN0(data_mem_out_wire[1733]), .IN1(data_in[5]), .SEL(n10792), 
        .F(n6007) );
  MUX U12560 ( .IN0(data_mem_out_wire[1732]), .IN1(data_in[4]), .SEL(n10792), 
        .F(n6006) );
  MUX U12561 ( .IN0(data_mem_out_wire[1731]), .IN1(data_in[3]), .SEL(n10792), 
        .F(n6005) );
  IV U12562 ( .A(n10793), .Z(n10792) );
  MUX U12563 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1730]), .SEL(n10793), 
        .F(n6004) );
  MUX U12564 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1729]), .SEL(n10793), 
        .F(n6003) );
  MUX U12565 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1728]), .SEL(n10793), 
        .F(n6002) );
  AND U12566 ( .A(n10790), .B(n10794), .Z(n10793) );
  NANDN U12567 ( .A(n10783), .B(n9792), .Z(n10794) );
  AND U12568 ( .A(n10795), .B(n10780), .Z(n10790) );
  NANDN U12569 ( .A(n10783), .B(n9796), .Z(n10780) );
  NANDN U12570 ( .A(n10783), .B(n9818), .Z(n10795) );
  NAND U12571 ( .A(n9919), .B(n10687), .Z(n10783) );
  MUX U12572 ( .IN0(n9746), .IN1(data_mem_out_wire[1791]), .SEL(n10796), .F(
        n6001) );
  MUX U12573 ( .IN0(n9748), .IN1(data_mem_out_wire[1790]), .SEL(n10796), .F(
        n6000) );
  MUX U12574 ( .IN0(n9749), .IN1(data_mem_out_wire[1789]), .SEL(n10796), .F(
        n5999) );
  MUX U12575 ( .IN0(n9750), .IN1(data_mem_out_wire[1788]), .SEL(n10796), .F(
        n5998) );
  MUX U12576 ( .IN0(n9751), .IN1(data_mem_out_wire[1787]), .SEL(n10796), .F(
        n5997) );
  MUX U12577 ( .IN0(n9752), .IN1(data_mem_out_wire[1786]), .SEL(n10796), .F(
        n5996) );
  MUX U12578 ( .IN0(n9753), .IN1(data_mem_out_wire[1785]), .SEL(n10796), .F(
        n5995) );
  MUX U12579 ( .IN0(n9754), .IN1(data_mem_out_wire[1784]), .SEL(n10796), .F(
        n5994) );
  AND U12580 ( .A(n10797), .B(n10798), .Z(n10796) );
  AND U12581 ( .A(n10799), .B(n10800), .Z(n10797) );
  OR U12582 ( .A(n9760), .B(n10801), .Z(n10800) );
  MUX U12583 ( .IN0(data_mem_out_wire[1783]), .IN1(n9761), .SEL(n10802), .F(
        n5993) );
  MUX U12584 ( .IN0(data_mem_out_wire[1782]), .IN1(n9763), .SEL(n10802), .F(
        n5992) );
  MUX U12585 ( .IN0(data_mem_out_wire[1781]), .IN1(n9764), .SEL(n10802), .F(
        n5991) );
  MUX U12586 ( .IN0(data_mem_out_wire[1780]), .IN1(n9765), .SEL(n10802), .F(
        n5990) );
  MUX U12587 ( .IN0(data_mem_out_wire[1779]), .IN1(n9766), .SEL(n10802), .F(
        n5989) );
  IV U12588 ( .A(n10803), .Z(n10802) );
  MUX U12589 ( .IN0(n9768), .IN1(data_mem_out_wire[1778]), .SEL(n10803), .F(
        n5988) );
  MUX U12590 ( .IN0(n9769), .IN1(data_mem_out_wire[1777]), .SEL(n10803), .F(
        n5987) );
  MUX U12591 ( .IN0(n9770), .IN1(data_mem_out_wire[1776]), .SEL(n10803), .F(
        n5986) );
  AND U12592 ( .A(n10804), .B(n10805), .Z(n10803) );
  OR U12593 ( .A(n9773), .B(n10801), .Z(n10805) );
  AND U12594 ( .A(n10799), .B(n10798), .Z(n10804) );
  NANDN U12595 ( .A(n10801), .B(n9809), .Z(n10799) );
  MUX U12596 ( .IN0(data_mem_out_wire[1775]), .IN1(n9776), .SEL(n10806), .F(
        n5985) );
  MUX U12597 ( .IN0(data_mem_out_wire[1774]), .IN1(n9778), .SEL(n10806), .F(
        n5984) );
  MUX U12598 ( .IN0(data_mem_out_wire[1773]), .IN1(n9779), .SEL(n10806), .F(
        n5983) );
  MUX U12599 ( .IN0(data_mem_out_wire[1772]), .IN1(n9780), .SEL(n10806), .F(
        n5982) );
  MUX U12600 ( .IN0(data_mem_out_wire[1771]), .IN1(n9781), .SEL(n10806), .F(
        n5981) );
  IV U12601 ( .A(n10807), .Z(n10806) );
  MUX U12602 ( .IN0(n9783), .IN1(data_mem_out_wire[1770]), .SEL(n10807), .F(
        n5980) );
  MUX U12603 ( .IN0(n9784), .IN1(data_mem_out_wire[1769]), .SEL(n10807), .F(
        n5979) );
  MUX U12604 ( .IN0(n9785), .IN1(data_mem_out_wire[1768]), .SEL(n10807), .F(
        n5978) );
  AND U12605 ( .A(n10808), .B(n10809), .Z(n10807) );
  OR U12606 ( .A(n9788), .B(n10801), .Z(n10809) );
  MUX U12607 ( .IN0(data_mem_out_wire[1767]), .IN1(data_in[7]), .SEL(n10810), 
        .F(n5977) );
  MUX U12608 ( .IN0(data_mem_out_wire[1766]), .IN1(data_in[6]), .SEL(n10810), 
        .F(n5976) );
  MUX U12609 ( .IN0(data_mem_out_wire[1765]), .IN1(data_in[5]), .SEL(n10810), 
        .F(n5975) );
  MUX U12610 ( .IN0(data_mem_out_wire[1764]), .IN1(data_in[4]), .SEL(n10810), 
        .F(n5974) );
  MUX U12611 ( .IN0(data_mem_out_wire[1763]), .IN1(data_in[3]), .SEL(n10810), 
        .F(n5973) );
  IV U12612 ( .A(n10811), .Z(n10810) );
  MUX U12613 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1762]), .SEL(n10811), 
        .F(n5972) );
  MUX U12614 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1761]), .SEL(n10811), 
        .F(n5971) );
  MUX U12615 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1760]), .SEL(n10811), 
        .F(n5970) );
  AND U12616 ( .A(n10808), .B(n10812), .Z(n10811) );
  NANDN U12617 ( .A(n10801), .B(n9792), .Z(n10812) );
  AND U12618 ( .A(n10813), .B(n10798), .Z(n10808) );
  NANDN U12619 ( .A(n10801), .B(n9796), .Z(n10798) );
  NANDN U12620 ( .A(n10801), .B(n9818), .Z(n10813) );
  NAND U12621 ( .A(n10687), .B(n9938), .Z(n10801) );
  AND U12622 ( .A(n10231), .B(N42), .Z(n10687) );
  NOR U12623 ( .A(n10668), .B(N40), .Z(n10231) );
  IV U12624 ( .A(N41), .Z(n10668) );
  MUX U12625 ( .IN0(n9746), .IN1(data_mem_out_wire[1823]), .SEL(n10814), .F(
        n5969) );
  MUX U12626 ( .IN0(n9748), .IN1(data_mem_out_wire[1822]), .SEL(n10814), .F(
        n5968) );
  MUX U12627 ( .IN0(n9749), .IN1(data_mem_out_wire[1821]), .SEL(n10814), .F(
        n5967) );
  MUX U12628 ( .IN0(n9750), .IN1(data_mem_out_wire[1820]), .SEL(n10814), .F(
        n5966) );
  MUX U12629 ( .IN0(n9751), .IN1(data_mem_out_wire[1819]), .SEL(n10814), .F(
        n5965) );
  MUX U12630 ( .IN0(n9752), .IN1(data_mem_out_wire[1818]), .SEL(n10814), .F(
        n5964) );
  MUX U12631 ( .IN0(n9753), .IN1(data_mem_out_wire[1817]), .SEL(n10814), .F(
        n5963) );
  MUX U12632 ( .IN0(n9754), .IN1(data_mem_out_wire[1816]), .SEL(n10814), .F(
        n5962) );
  AND U12633 ( .A(n10815), .B(n10816), .Z(n10814) );
  AND U12634 ( .A(n10817), .B(n10818), .Z(n10815) );
  OR U12635 ( .A(n9760), .B(n10819), .Z(n10818) );
  MUX U12636 ( .IN0(data_mem_out_wire[1815]), .IN1(n9761), .SEL(n10820), .F(
        n5961) );
  MUX U12637 ( .IN0(data_mem_out_wire[1814]), .IN1(n9763), .SEL(n10820), .F(
        n5960) );
  MUX U12638 ( .IN0(data_mem_out_wire[1813]), .IN1(n9764), .SEL(n10820), .F(
        n5959) );
  MUX U12639 ( .IN0(data_mem_out_wire[1812]), .IN1(n9765), .SEL(n10820), .F(
        n5958) );
  MUX U12640 ( .IN0(data_mem_out_wire[1811]), .IN1(n9766), .SEL(n10820), .F(
        n5957) );
  IV U12641 ( .A(n10821), .Z(n10820) );
  MUX U12642 ( .IN0(n9768), .IN1(data_mem_out_wire[1810]), .SEL(n10821), .F(
        n5956) );
  MUX U12643 ( .IN0(n9769), .IN1(data_mem_out_wire[1809]), .SEL(n10821), .F(
        n5955) );
  MUX U12644 ( .IN0(n9770), .IN1(data_mem_out_wire[1808]), .SEL(n10821), .F(
        n5954) );
  AND U12645 ( .A(n10822), .B(n10823), .Z(n10821) );
  OR U12646 ( .A(n9773), .B(n10819), .Z(n10823) );
  AND U12647 ( .A(n10817), .B(n10816), .Z(n10822) );
  NANDN U12648 ( .A(n10819), .B(n9809), .Z(n10817) );
  MUX U12649 ( .IN0(data_mem_out_wire[1807]), .IN1(n9776), .SEL(n10824), .F(
        n5953) );
  MUX U12650 ( .IN0(data_mem_out_wire[1806]), .IN1(n9778), .SEL(n10824), .F(
        n5952) );
  MUX U12651 ( .IN0(data_mem_out_wire[1805]), .IN1(n9779), .SEL(n10824), .F(
        n5951) );
  MUX U12652 ( .IN0(data_mem_out_wire[1804]), .IN1(n9780), .SEL(n10824), .F(
        n5950) );
  MUX U12653 ( .IN0(data_mem_out_wire[1803]), .IN1(n9781), .SEL(n10824), .F(
        n5949) );
  IV U12654 ( .A(n10825), .Z(n10824) );
  MUX U12655 ( .IN0(n9783), .IN1(data_mem_out_wire[1802]), .SEL(n10825), .F(
        n5948) );
  MUX U12656 ( .IN0(n9784), .IN1(data_mem_out_wire[1801]), .SEL(n10825), .F(
        n5947) );
  MUX U12657 ( .IN0(n9785), .IN1(data_mem_out_wire[1800]), .SEL(n10825), .F(
        n5946) );
  AND U12658 ( .A(n10826), .B(n10827), .Z(n10825) );
  OR U12659 ( .A(n9788), .B(n10819), .Z(n10827) );
  MUX U12660 ( .IN0(data_mem_out_wire[1799]), .IN1(data_in[7]), .SEL(n10828), 
        .F(n5945) );
  MUX U12661 ( .IN0(data_mem_out_wire[1798]), .IN1(data_in[6]), .SEL(n10828), 
        .F(n5944) );
  MUX U12662 ( .IN0(data_mem_out_wire[1797]), .IN1(data_in[5]), .SEL(n10828), 
        .F(n5943) );
  MUX U12663 ( .IN0(data_mem_out_wire[1796]), .IN1(data_in[4]), .SEL(n10828), 
        .F(n5942) );
  MUX U12664 ( .IN0(data_mem_out_wire[1795]), .IN1(data_in[3]), .SEL(n10828), 
        .F(n5941) );
  IV U12665 ( .A(n10829), .Z(n10828) );
  MUX U12666 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1794]), .SEL(n10829), 
        .F(n5940) );
  MUX U12667 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1793]), .SEL(n10829), 
        .F(n5939) );
  MUX U12668 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1792]), .SEL(n10829), 
        .F(n5938) );
  AND U12669 ( .A(n10826), .B(n10830), .Z(n10829) );
  NANDN U12670 ( .A(n10819), .B(n9792), .Z(n10830) );
  AND U12671 ( .A(n10831), .B(n10816), .Z(n10826) );
  NANDN U12672 ( .A(n10819), .B(n9796), .Z(n10816) );
  NANDN U12673 ( .A(n10819), .B(n9818), .Z(n10831) );
  NANDN U12674 ( .A(n10832), .B(n9798), .Z(n10819) );
  ANDN U12675 ( .B(n10833), .A(N39), .Z(n9798) );
  MUX U12676 ( .IN0(n9746), .IN1(data_mem_out_wire[1855]), .SEL(n10834), .F(
        n5937) );
  MUX U12677 ( .IN0(n9748), .IN1(data_mem_out_wire[1854]), .SEL(n10834), .F(
        n5936) );
  MUX U12678 ( .IN0(n9749), .IN1(data_mem_out_wire[1853]), .SEL(n10834), .F(
        n5935) );
  MUX U12679 ( .IN0(n9750), .IN1(data_mem_out_wire[1852]), .SEL(n10834), .F(
        n5934) );
  MUX U12680 ( .IN0(n9751), .IN1(data_mem_out_wire[1851]), .SEL(n10834), .F(
        n5933) );
  MUX U12681 ( .IN0(n9752), .IN1(data_mem_out_wire[1850]), .SEL(n10834), .F(
        n5932) );
  MUX U12682 ( .IN0(n9753), .IN1(data_mem_out_wire[1849]), .SEL(n10834), .F(
        n5931) );
  MUX U12683 ( .IN0(n9754), .IN1(data_mem_out_wire[1848]), .SEL(n10834), .F(
        n5930) );
  AND U12684 ( .A(n10835), .B(n10836), .Z(n10834) );
  AND U12685 ( .A(n10837), .B(n10838), .Z(n10835) );
  OR U12686 ( .A(n9760), .B(n10839), .Z(n10838) );
  MUX U12687 ( .IN0(data_mem_out_wire[1847]), .IN1(n9761), .SEL(n10840), .F(
        n5929) );
  MUX U12688 ( .IN0(data_mem_out_wire[1846]), .IN1(n9763), .SEL(n10840), .F(
        n5928) );
  MUX U12689 ( .IN0(data_mem_out_wire[1845]), .IN1(n9764), .SEL(n10840), .F(
        n5927) );
  MUX U12690 ( .IN0(data_mem_out_wire[1844]), .IN1(n9765), .SEL(n10840), .F(
        n5926) );
  MUX U12691 ( .IN0(data_mem_out_wire[1843]), .IN1(n9766), .SEL(n10840), .F(
        n5925) );
  IV U12692 ( .A(n10841), .Z(n10840) );
  MUX U12693 ( .IN0(n9768), .IN1(data_mem_out_wire[1842]), .SEL(n10841), .F(
        n5924) );
  MUX U12694 ( .IN0(n9769), .IN1(data_mem_out_wire[1841]), .SEL(n10841), .F(
        n5923) );
  MUX U12695 ( .IN0(n9770), .IN1(data_mem_out_wire[1840]), .SEL(n10841), .F(
        n5922) );
  AND U12696 ( .A(n10842), .B(n10843), .Z(n10841) );
  OR U12697 ( .A(n9773), .B(n10839), .Z(n10843) );
  AND U12698 ( .A(n10837), .B(n10836), .Z(n10842) );
  NANDN U12699 ( .A(n10839), .B(n9809), .Z(n10837) );
  MUX U12700 ( .IN0(data_mem_out_wire[1839]), .IN1(n9776), .SEL(n10844), .F(
        n5921) );
  MUX U12701 ( .IN0(data_mem_out_wire[1838]), .IN1(n9778), .SEL(n10844), .F(
        n5920) );
  MUX U12702 ( .IN0(data_mem_out_wire[1837]), .IN1(n9779), .SEL(n10844), .F(
        n5919) );
  MUX U12703 ( .IN0(data_mem_out_wire[1836]), .IN1(n9780), .SEL(n10844), .F(
        n5918) );
  MUX U12704 ( .IN0(data_mem_out_wire[1835]), .IN1(n9781), .SEL(n10844), .F(
        n5917) );
  IV U12705 ( .A(n10845), .Z(n10844) );
  MUX U12706 ( .IN0(n9783), .IN1(data_mem_out_wire[1834]), .SEL(n10845), .F(
        n5916) );
  MUX U12707 ( .IN0(n9784), .IN1(data_mem_out_wire[1833]), .SEL(n10845), .F(
        n5915) );
  MUX U12708 ( .IN0(n9785), .IN1(data_mem_out_wire[1832]), .SEL(n10845), .F(
        n5914) );
  AND U12709 ( .A(n10846), .B(n10847), .Z(n10845) );
  OR U12710 ( .A(n9788), .B(n10839), .Z(n10847) );
  MUX U12711 ( .IN0(data_mem_out_wire[1831]), .IN1(data_in[7]), .SEL(n10848), 
        .F(n5913) );
  MUX U12712 ( .IN0(data_mem_out_wire[1830]), .IN1(data_in[6]), .SEL(n10848), 
        .F(n5912) );
  MUX U12713 ( .IN0(data_mem_out_wire[1829]), .IN1(data_in[5]), .SEL(n10848), 
        .F(n5911) );
  MUX U12714 ( .IN0(data_mem_out_wire[1828]), .IN1(data_in[4]), .SEL(n10848), 
        .F(n5910) );
  MUX U12715 ( .IN0(data_mem_out_wire[1827]), .IN1(data_in[3]), .SEL(n10848), 
        .F(n5909) );
  IV U12716 ( .A(n10849), .Z(n10848) );
  MUX U12717 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1826]), .SEL(n10849), 
        .F(n5908) );
  MUX U12718 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1825]), .SEL(n10849), 
        .F(n5907) );
  MUX U12719 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1824]), .SEL(n10849), 
        .F(n5906) );
  AND U12720 ( .A(n10846), .B(n10850), .Z(n10849) );
  NANDN U12721 ( .A(n10839), .B(n9792), .Z(n10850) );
  AND U12722 ( .A(n10851), .B(n10836), .Z(n10846) );
  NANDN U12723 ( .A(n10839), .B(n9796), .Z(n10836) );
  NANDN U12724 ( .A(n10839), .B(n9818), .Z(n10851) );
  NANDN U12725 ( .A(n10832), .B(n9819), .Z(n10839) );
  ANDN U12726 ( .B(n10852), .A(N39), .Z(n9819) );
  MUX U12727 ( .IN0(n9746), .IN1(data_mem_out_wire[1887]), .SEL(n10853), .F(
        n5905) );
  MUX U12728 ( .IN0(n9748), .IN1(data_mem_out_wire[1886]), .SEL(n10853), .F(
        n5904) );
  MUX U12729 ( .IN0(n9749), .IN1(data_mem_out_wire[1885]), .SEL(n10853), .F(
        n5903) );
  MUX U12730 ( .IN0(n9750), .IN1(data_mem_out_wire[1884]), .SEL(n10853), .F(
        n5902) );
  MUX U12731 ( .IN0(n9751), .IN1(data_mem_out_wire[1883]), .SEL(n10853), .F(
        n5901) );
  MUX U12732 ( .IN0(n9752), .IN1(data_mem_out_wire[1882]), .SEL(n10853), .F(
        n5900) );
  MUX U12733 ( .IN0(n9753), .IN1(data_mem_out_wire[1881]), .SEL(n10853), .F(
        n5899) );
  MUX U12734 ( .IN0(n9754), .IN1(data_mem_out_wire[1880]), .SEL(n10853), .F(
        n5898) );
  AND U12735 ( .A(n10854), .B(n10855), .Z(n10853) );
  AND U12736 ( .A(n10856), .B(n10857), .Z(n10854) );
  OR U12737 ( .A(n9760), .B(n10858), .Z(n10857) );
  MUX U12738 ( .IN0(data_mem_out_wire[1879]), .IN1(n9761), .SEL(n10859), .F(
        n5897) );
  MUX U12739 ( .IN0(data_mem_out_wire[1878]), .IN1(n9763), .SEL(n10859), .F(
        n5896) );
  MUX U12740 ( .IN0(data_mem_out_wire[1877]), .IN1(n9764), .SEL(n10859), .F(
        n5895) );
  MUX U12741 ( .IN0(data_mem_out_wire[1876]), .IN1(n9765), .SEL(n10859), .F(
        n5894) );
  MUX U12742 ( .IN0(data_mem_out_wire[1875]), .IN1(n9766), .SEL(n10859), .F(
        n5893) );
  IV U12743 ( .A(n10860), .Z(n10859) );
  MUX U12744 ( .IN0(n9768), .IN1(data_mem_out_wire[1874]), .SEL(n10860), .F(
        n5892) );
  MUX U12745 ( .IN0(n9769), .IN1(data_mem_out_wire[1873]), .SEL(n10860), .F(
        n5891) );
  MUX U12746 ( .IN0(n9770), .IN1(data_mem_out_wire[1872]), .SEL(n10860), .F(
        n5890) );
  AND U12747 ( .A(n10861), .B(n10862), .Z(n10860) );
  OR U12748 ( .A(n9773), .B(n10858), .Z(n10862) );
  AND U12749 ( .A(n10856), .B(n10855), .Z(n10861) );
  NANDN U12750 ( .A(n10858), .B(n9809), .Z(n10856) );
  MUX U12751 ( .IN0(data_mem_out_wire[1871]), .IN1(n9776), .SEL(n10863), .F(
        n5889) );
  MUX U12752 ( .IN0(data_mem_out_wire[1870]), .IN1(n9778), .SEL(n10863), .F(
        n5888) );
  MUX U12753 ( .IN0(data_mem_out_wire[1869]), .IN1(n9779), .SEL(n10863), .F(
        n5887) );
  MUX U12754 ( .IN0(data_mem_out_wire[1868]), .IN1(n9780), .SEL(n10863), .F(
        n5886) );
  MUX U12755 ( .IN0(data_mem_out_wire[1867]), .IN1(n9781), .SEL(n10863), .F(
        n5885) );
  IV U12756 ( .A(n10864), .Z(n10863) );
  MUX U12757 ( .IN0(n9783), .IN1(data_mem_out_wire[1866]), .SEL(n10864), .F(
        n5884) );
  MUX U12758 ( .IN0(n9784), .IN1(data_mem_out_wire[1865]), .SEL(n10864), .F(
        n5883) );
  MUX U12759 ( .IN0(n9785), .IN1(data_mem_out_wire[1864]), .SEL(n10864), .F(
        n5882) );
  AND U12760 ( .A(n10865), .B(n10866), .Z(n10864) );
  OR U12761 ( .A(n9788), .B(n10858), .Z(n10866) );
  MUX U12762 ( .IN0(data_mem_out_wire[1863]), .IN1(data_in[7]), .SEL(n10867), 
        .F(n5881) );
  MUX U12763 ( .IN0(data_mem_out_wire[1862]), .IN1(data_in[6]), .SEL(n10867), 
        .F(n5880) );
  MUX U12764 ( .IN0(data_mem_out_wire[1861]), .IN1(data_in[5]), .SEL(n10867), 
        .F(n5879) );
  MUX U12765 ( .IN0(data_mem_out_wire[1860]), .IN1(data_in[4]), .SEL(n10867), 
        .F(n5878) );
  MUX U12766 ( .IN0(data_mem_out_wire[1859]), .IN1(data_in[3]), .SEL(n10867), 
        .F(n5877) );
  IV U12767 ( .A(n10868), .Z(n10867) );
  MUX U12768 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1858]), .SEL(n10868), 
        .F(n5876) );
  MUX U12769 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1857]), .SEL(n10868), 
        .F(n5875) );
  MUX U12770 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1856]), .SEL(n10868), 
        .F(n5874) );
  AND U12771 ( .A(n10865), .B(n10869), .Z(n10868) );
  NANDN U12772 ( .A(n10858), .B(n9792), .Z(n10869) );
  AND U12773 ( .A(n10870), .B(n10855), .Z(n10865) );
  NANDN U12774 ( .A(n10858), .B(n9796), .Z(n10855) );
  NANDN U12775 ( .A(n10858), .B(n9818), .Z(n10870) );
  NANDN U12776 ( .A(n10832), .B(n9838), .Z(n10858) );
  ANDN U12777 ( .B(n10871), .A(N39), .Z(n9838) );
  MUX U12778 ( .IN0(n9746), .IN1(data_mem_out_wire[1919]), .SEL(n10872), .F(
        n5873) );
  MUX U12779 ( .IN0(n9748), .IN1(data_mem_out_wire[1918]), .SEL(n10872), .F(
        n5872) );
  MUX U12780 ( .IN0(n9749), .IN1(data_mem_out_wire[1917]), .SEL(n10872), .F(
        n5871) );
  MUX U12781 ( .IN0(n9750), .IN1(data_mem_out_wire[1916]), .SEL(n10872), .F(
        n5870) );
  MUX U12782 ( .IN0(n9751), .IN1(data_mem_out_wire[1915]), .SEL(n10872), .F(
        n5869) );
  MUX U12783 ( .IN0(n9752), .IN1(data_mem_out_wire[1914]), .SEL(n10872), .F(
        n5868) );
  MUX U12784 ( .IN0(n9753), .IN1(data_mem_out_wire[1913]), .SEL(n10872), .F(
        n5867) );
  MUX U12785 ( .IN0(n9754), .IN1(data_mem_out_wire[1912]), .SEL(n10872), .F(
        n5866) );
  AND U12786 ( .A(n10873), .B(n10874), .Z(n10872) );
  AND U12787 ( .A(n10875), .B(n10876), .Z(n10873) );
  OR U12788 ( .A(n9760), .B(n10877), .Z(n10876) );
  MUX U12789 ( .IN0(data_mem_out_wire[1911]), .IN1(n9761), .SEL(n10878), .F(
        n5865) );
  MUX U12790 ( .IN0(data_mem_out_wire[1910]), .IN1(n9763), .SEL(n10878), .F(
        n5864) );
  MUX U12791 ( .IN0(data_mem_out_wire[1909]), .IN1(n9764), .SEL(n10878), .F(
        n5863) );
  MUX U12792 ( .IN0(data_mem_out_wire[1908]), .IN1(n9765), .SEL(n10878), .F(
        n5862) );
  MUX U12793 ( .IN0(data_mem_out_wire[1907]), .IN1(n9766), .SEL(n10878), .F(
        n5861) );
  IV U12794 ( .A(n10879), .Z(n10878) );
  MUX U12795 ( .IN0(n9768), .IN1(data_mem_out_wire[1906]), .SEL(n10879), .F(
        n5860) );
  MUX U12796 ( .IN0(n9769), .IN1(data_mem_out_wire[1905]), .SEL(n10879), .F(
        n5859) );
  MUX U12797 ( .IN0(n9770), .IN1(data_mem_out_wire[1904]), .SEL(n10879), .F(
        n5858) );
  AND U12798 ( .A(n10880), .B(n10881), .Z(n10879) );
  OR U12799 ( .A(n9773), .B(n10877), .Z(n10881) );
  AND U12800 ( .A(n10875), .B(n10874), .Z(n10880) );
  NANDN U12801 ( .A(n10877), .B(n9809), .Z(n10875) );
  MUX U12802 ( .IN0(data_mem_out_wire[1903]), .IN1(n9776), .SEL(n10882), .F(
        n5857) );
  MUX U12803 ( .IN0(data_mem_out_wire[1902]), .IN1(n9778), .SEL(n10882), .F(
        n5856) );
  MUX U12804 ( .IN0(data_mem_out_wire[1901]), .IN1(n9779), .SEL(n10882), .F(
        n5855) );
  MUX U12805 ( .IN0(data_mem_out_wire[1900]), .IN1(n9780), .SEL(n10882), .F(
        n5854) );
  MUX U12806 ( .IN0(data_mem_out_wire[1899]), .IN1(n9781), .SEL(n10882), .F(
        n5853) );
  IV U12807 ( .A(n10883), .Z(n10882) );
  MUX U12808 ( .IN0(n9783), .IN1(data_mem_out_wire[1898]), .SEL(n10883), .F(
        n5852) );
  MUX U12809 ( .IN0(n9784), .IN1(data_mem_out_wire[1897]), .SEL(n10883), .F(
        n5851) );
  MUX U12810 ( .IN0(n9785), .IN1(data_mem_out_wire[1896]), .SEL(n10883), .F(
        n5850) );
  AND U12811 ( .A(n10884), .B(n10885), .Z(n10883) );
  OR U12812 ( .A(n9788), .B(n10877), .Z(n10885) );
  MUX U12813 ( .IN0(data_mem_out_wire[1895]), .IN1(data_in[7]), .SEL(n10886), 
        .F(n5849) );
  MUX U12814 ( .IN0(data_mem_out_wire[1894]), .IN1(data_in[6]), .SEL(n10886), 
        .F(n5848) );
  MUX U12815 ( .IN0(data_mem_out_wire[1893]), .IN1(data_in[5]), .SEL(n10886), 
        .F(n5847) );
  MUX U12816 ( .IN0(data_mem_out_wire[1892]), .IN1(data_in[4]), .SEL(n10886), 
        .F(n5846) );
  MUX U12817 ( .IN0(data_mem_out_wire[1891]), .IN1(data_in[3]), .SEL(n10886), 
        .F(n5845) );
  IV U12818 ( .A(n10887), .Z(n10886) );
  MUX U12819 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1890]), .SEL(n10887), 
        .F(n5844) );
  MUX U12820 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1889]), .SEL(n10887), 
        .F(n5843) );
  MUX U12821 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1888]), .SEL(n10887), 
        .F(n5842) );
  AND U12822 ( .A(n10884), .B(n10888), .Z(n10887) );
  NANDN U12823 ( .A(n10877), .B(n9792), .Z(n10888) );
  AND U12824 ( .A(n10889), .B(n10874), .Z(n10884) );
  NANDN U12825 ( .A(n10877), .B(n9796), .Z(n10874) );
  NANDN U12826 ( .A(n10877), .B(n9818), .Z(n10889) );
  NANDN U12827 ( .A(n10832), .B(n9862), .Z(n10877) );
  ANDN U12828 ( .B(n10890), .A(N39), .Z(n9862) );
  MUX U12829 ( .IN0(n9746), .IN1(data_mem_out_wire[1951]), .SEL(n10891), .F(
        n5841) );
  MUX U12830 ( .IN0(n9748), .IN1(data_mem_out_wire[1950]), .SEL(n10891), .F(
        n5840) );
  MUX U12831 ( .IN0(n9749), .IN1(data_mem_out_wire[1949]), .SEL(n10891), .F(
        n5839) );
  MUX U12832 ( .IN0(n9750), .IN1(data_mem_out_wire[1948]), .SEL(n10891), .F(
        n5838) );
  MUX U12833 ( .IN0(n9751), .IN1(data_mem_out_wire[1947]), .SEL(n10891), .F(
        n5837) );
  MUX U12834 ( .IN0(n9752), .IN1(data_mem_out_wire[1946]), .SEL(n10891), .F(
        n5836) );
  MUX U12835 ( .IN0(n9753), .IN1(data_mem_out_wire[1945]), .SEL(n10891), .F(
        n5835) );
  MUX U12836 ( .IN0(n9754), .IN1(data_mem_out_wire[1944]), .SEL(n10891), .F(
        n5834) );
  AND U12837 ( .A(n10892), .B(n10893), .Z(n10891) );
  AND U12838 ( .A(n10894), .B(n10895), .Z(n10892) );
  OR U12839 ( .A(n9760), .B(n10896), .Z(n10895) );
  MUX U12840 ( .IN0(data_mem_out_wire[1943]), .IN1(n9761), .SEL(n10897), .F(
        n5833) );
  MUX U12841 ( .IN0(data_mem_out_wire[1942]), .IN1(n9763), .SEL(n10897), .F(
        n5832) );
  MUX U12842 ( .IN0(data_mem_out_wire[1941]), .IN1(n9764), .SEL(n10897), .F(
        n5831) );
  MUX U12843 ( .IN0(data_mem_out_wire[1940]), .IN1(n9765), .SEL(n10897), .F(
        n5830) );
  MUX U12844 ( .IN0(data_mem_out_wire[1939]), .IN1(n9766), .SEL(n10897), .F(
        n5829) );
  IV U12845 ( .A(n10898), .Z(n10897) );
  MUX U12846 ( .IN0(n9768), .IN1(data_mem_out_wire[1938]), .SEL(n10898), .F(
        n5828) );
  MUX U12847 ( .IN0(n9769), .IN1(data_mem_out_wire[1937]), .SEL(n10898), .F(
        n5827) );
  MUX U12848 ( .IN0(n9770), .IN1(data_mem_out_wire[1936]), .SEL(n10898), .F(
        n5826) );
  AND U12849 ( .A(n10899), .B(n10900), .Z(n10898) );
  OR U12850 ( .A(n9773), .B(n10896), .Z(n10900) );
  AND U12851 ( .A(n10894), .B(n10893), .Z(n10899) );
  NANDN U12852 ( .A(n10896), .B(n9809), .Z(n10894) );
  MUX U12853 ( .IN0(data_mem_out_wire[1935]), .IN1(n9776), .SEL(n10901), .F(
        n5825) );
  MUX U12854 ( .IN0(data_mem_out_wire[1934]), .IN1(n9778), .SEL(n10901), .F(
        n5824) );
  MUX U12855 ( .IN0(data_mem_out_wire[1933]), .IN1(n9779), .SEL(n10901), .F(
        n5823) );
  MUX U12856 ( .IN0(data_mem_out_wire[1932]), .IN1(n9780), .SEL(n10901), .F(
        n5822) );
  MUX U12857 ( .IN0(data_mem_out_wire[1931]), .IN1(n9781), .SEL(n10901), .F(
        n5821) );
  IV U12858 ( .A(n10902), .Z(n10901) );
  MUX U12859 ( .IN0(n9783), .IN1(data_mem_out_wire[1930]), .SEL(n10902), .F(
        n5820) );
  MUX U12860 ( .IN0(n9784), .IN1(data_mem_out_wire[1929]), .SEL(n10902), .F(
        n5819) );
  MUX U12861 ( .IN0(n9785), .IN1(data_mem_out_wire[1928]), .SEL(n10902), .F(
        n5818) );
  AND U12862 ( .A(n10903), .B(n10904), .Z(n10902) );
  OR U12863 ( .A(n9788), .B(n10896), .Z(n10904) );
  MUX U12864 ( .IN0(data_mem_out_wire[1927]), .IN1(data_in[7]), .SEL(n10905), 
        .F(n5817) );
  MUX U12865 ( .IN0(data_mem_out_wire[1926]), .IN1(data_in[6]), .SEL(n10905), 
        .F(n5816) );
  MUX U12866 ( .IN0(data_mem_out_wire[1925]), .IN1(data_in[5]), .SEL(n10905), 
        .F(n5815) );
  MUX U12867 ( .IN0(data_mem_out_wire[1924]), .IN1(data_in[4]), .SEL(n10905), 
        .F(n5814) );
  MUX U12868 ( .IN0(data_mem_out_wire[1923]), .IN1(data_in[3]), .SEL(n10905), 
        .F(n5813) );
  IV U12869 ( .A(n10906), .Z(n10905) );
  MUX U12870 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1922]), .SEL(n10906), 
        .F(n5812) );
  MUX U12871 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1921]), .SEL(n10906), 
        .F(n5811) );
  MUX U12872 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1920]), .SEL(n10906), 
        .F(n5810) );
  AND U12873 ( .A(n10903), .B(n10907), .Z(n10906) );
  NANDN U12874 ( .A(n10896), .B(n9792), .Z(n10907) );
  AND U12875 ( .A(n10908), .B(n10893), .Z(n10903) );
  NANDN U12876 ( .A(n10896), .B(n9796), .Z(n10893) );
  NANDN U12877 ( .A(n10896), .B(n9818), .Z(n10908) );
  NANDN U12878 ( .A(n10832), .B(n9881), .Z(n10896) );
  AND U12879 ( .A(n10833), .B(N39), .Z(n9881) );
  NOR U12880 ( .A(N37), .B(N38), .Z(n10833) );
  MUX U12881 ( .IN0(n9746), .IN1(data_mem_out_wire[1983]), .SEL(n10909), .F(
        n5809) );
  MUX U12882 ( .IN0(n9748), .IN1(data_mem_out_wire[1982]), .SEL(n10909), .F(
        n5808) );
  MUX U12883 ( .IN0(n9749), .IN1(data_mem_out_wire[1981]), .SEL(n10909), .F(
        n5807) );
  MUX U12884 ( .IN0(n9750), .IN1(data_mem_out_wire[1980]), .SEL(n10909), .F(
        n5806) );
  MUX U12885 ( .IN0(n9751), .IN1(data_mem_out_wire[1979]), .SEL(n10909), .F(
        n5805) );
  MUX U12886 ( .IN0(n9752), .IN1(data_mem_out_wire[1978]), .SEL(n10909), .F(
        n5804) );
  MUX U12887 ( .IN0(n9753), .IN1(data_mem_out_wire[1977]), .SEL(n10909), .F(
        n5803) );
  MUX U12888 ( .IN0(n9754), .IN1(data_mem_out_wire[1976]), .SEL(n10909), .F(
        n5802) );
  AND U12889 ( .A(n10910), .B(n10911), .Z(n10909) );
  AND U12890 ( .A(n10912), .B(n10913), .Z(n10910) );
  OR U12891 ( .A(n9760), .B(n10914), .Z(n10913) );
  MUX U12892 ( .IN0(data_mem_out_wire[1975]), .IN1(n9761), .SEL(n10915), .F(
        n5801) );
  MUX U12893 ( .IN0(data_mem_out_wire[1974]), .IN1(n9763), .SEL(n10915), .F(
        n5800) );
  MUX U12894 ( .IN0(data_mem_out_wire[1973]), .IN1(n9764), .SEL(n10915), .F(
        n5799) );
  MUX U12895 ( .IN0(data_mem_out_wire[1972]), .IN1(n9765), .SEL(n10915), .F(
        n5798) );
  MUX U12896 ( .IN0(data_mem_out_wire[1971]), .IN1(n9766), .SEL(n10915), .F(
        n5797) );
  IV U12897 ( .A(n10916), .Z(n10915) );
  MUX U12898 ( .IN0(n9768), .IN1(data_mem_out_wire[1970]), .SEL(n10916), .F(
        n5796) );
  MUX U12899 ( .IN0(n9769), .IN1(data_mem_out_wire[1969]), .SEL(n10916), .F(
        n5795) );
  MUX U12900 ( .IN0(n9770), .IN1(data_mem_out_wire[1968]), .SEL(n10916), .F(
        n5794) );
  AND U12901 ( .A(n10917), .B(n10918), .Z(n10916) );
  OR U12902 ( .A(n9773), .B(n10914), .Z(n10918) );
  AND U12903 ( .A(n10912), .B(n10911), .Z(n10917) );
  NANDN U12904 ( .A(n10914), .B(n9809), .Z(n10912) );
  MUX U12905 ( .IN0(data_mem_out_wire[1967]), .IN1(n9776), .SEL(n10919), .F(
        n5793) );
  MUX U12906 ( .IN0(data_mem_out_wire[1966]), .IN1(n9778), .SEL(n10919), .F(
        n5792) );
  MUX U12907 ( .IN0(data_mem_out_wire[1965]), .IN1(n9779), .SEL(n10919), .F(
        n5791) );
  MUX U12908 ( .IN0(data_mem_out_wire[1964]), .IN1(n9780), .SEL(n10919), .F(
        n5790) );
  MUX U12909 ( .IN0(data_mem_out_wire[1963]), .IN1(n9781), .SEL(n10919), .F(
        n5789) );
  IV U12910 ( .A(n10920), .Z(n10919) );
  MUX U12911 ( .IN0(n9783), .IN1(data_mem_out_wire[1962]), .SEL(n10920), .F(
        n5788) );
  MUX U12912 ( .IN0(n9784), .IN1(data_mem_out_wire[1961]), .SEL(n10920), .F(
        n5787) );
  MUX U12913 ( .IN0(n9785), .IN1(data_mem_out_wire[1960]), .SEL(n10920), .F(
        n5786) );
  AND U12914 ( .A(n10921), .B(n10922), .Z(n10920) );
  OR U12915 ( .A(n9788), .B(n10914), .Z(n10922) );
  MUX U12916 ( .IN0(data_mem_out_wire[1959]), .IN1(data_in[7]), .SEL(n10923), 
        .F(n5785) );
  MUX U12917 ( .IN0(data_mem_out_wire[1958]), .IN1(data_in[6]), .SEL(n10923), 
        .F(n5784) );
  MUX U12918 ( .IN0(data_mem_out_wire[1957]), .IN1(data_in[5]), .SEL(n10923), 
        .F(n5783) );
  MUX U12919 ( .IN0(data_mem_out_wire[1956]), .IN1(data_in[4]), .SEL(n10923), 
        .F(n5782) );
  MUX U12920 ( .IN0(data_mem_out_wire[1955]), .IN1(data_in[3]), .SEL(n10923), 
        .F(n5781) );
  IV U12921 ( .A(n10924), .Z(n10923) );
  MUX U12922 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1954]), .SEL(n10924), 
        .F(n5780) );
  MUX U12923 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1953]), .SEL(n10924), 
        .F(n5779) );
  MUX U12924 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1952]), .SEL(n10924), 
        .F(n5778) );
  AND U12925 ( .A(n10921), .B(n10925), .Z(n10924) );
  NANDN U12926 ( .A(n10914), .B(n9792), .Z(n10925) );
  AND U12927 ( .A(n10926), .B(n10911), .Z(n10921) );
  NANDN U12928 ( .A(n10914), .B(n9796), .Z(n10911) );
  NANDN U12929 ( .A(n10914), .B(n9818), .Z(n10926) );
  NANDN U12930 ( .A(n10832), .B(n9900), .Z(n10914) );
  AND U12931 ( .A(n10852), .B(N39), .Z(n9900) );
  NOR U12932 ( .A(n10927), .B(N38), .Z(n10852) );
  MUX U12933 ( .IN0(n9746), .IN1(data_mem_out_wire[2015]), .SEL(n10928), .F(
        n5777) );
  MUX U12934 ( .IN0(n9748), .IN1(data_mem_out_wire[2014]), .SEL(n10928), .F(
        n5776) );
  MUX U12935 ( .IN0(n9749), .IN1(data_mem_out_wire[2013]), .SEL(n10928), .F(
        n5775) );
  MUX U12936 ( .IN0(n9750), .IN1(data_mem_out_wire[2012]), .SEL(n10928), .F(
        n5774) );
  MUX U12937 ( .IN0(n9751), .IN1(data_mem_out_wire[2011]), .SEL(n10928), .F(
        n5773) );
  MUX U12938 ( .IN0(n9752), .IN1(data_mem_out_wire[2010]), .SEL(n10928), .F(
        n5772) );
  MUX U12939 ( .IN0(n9753), .IN1(data_mem_out_wire[2009]), .SEL(n10928), .F(
        n5771) );
  MUX U12940 ( .IN0(n9754), .IN1(data_mem_out_wire[2008]), .SEL(n10928), .F(
        n5770) );
  AND U12941 ( .A(n10929), .B(n10930), .Z(n10928) );
  AND U12942 ( .A(n10931), .B(n10932), .Z(n10929) );
  OR U12943 ( .A(n9760), .B(n10933), .Z(n10932) );
  MUX U12944 ( .IN0(data_mem_out_wire[2007]), .IN1(n9761), .SEL(n10934), .F(
        n5769) );
  MUX U12945 ( .IN0(data_mem_out_wire[2006]), .IN1(n9763), .SEL(n10934), .F(
        n5768) );
  MUX U12946 ( .IN0(data_mem_out_wire[2005]), .IN1(n9764), .SEL(n10934), .F(
        n5767) );
  MUX U12947 ( .IN0(data_mem_out_wire[2004]), .IN1(n9765), .SEL(n10934), .F(
        n5766) );
  MUX U12948 ( .IN0(data_mem_out_wire[2003]), .IN1(n9766), .SEL(n10934), .F(
        n5765) );
  IV U12949 ( .A(n10935), .Z(n10934) );
  MUX U12950 ( .IN0(n9768), .IN1(data_mem_out_wire[2002]), .SEL(n10935), .F(
        n5764) );
  MUX U12951 ( .IN0(n9769), .IN1(data_mem_out_wire[2001]), .SEL(n10935), .F(
        n5763) );
  MUX U12952 ( .IN0(n9770), .IN1(data_mem_out_wire[2000]), .SEL(n10935), .F(
        n5762) );
  AND U12953 ( .A(n10936), .B(n10937), .Z(n10935) );
  OR U12954 ( .A(n9773), .B(n10933), .Z(n10937) );
  AND U12955 ( .A(n10931), .B(n10930), .Z(n10936) );
  NANDN U12956 ( .A(n10933), .B(n9809), .Z(n10931) );
  MUX U12957 ( .IN0(data_mem_out_wire[1999]), .IN1(n9776), .SEL(n10938), .F(
        n5761) );
  MUX U12958 ( .IN0(data_mem_out_wire[1998]), .IN1(n9778), .SEL(n10938), .F(
        n5760) );
  MUX U12959 ( .IN0(data_mem_out_wire[1997]), .IN1(n9779), .SEL(n10938), .F(
        n5759) );
  MUX U12960 ( .IN0(data_mem_out_wire[1996]), .IN1(n9780), .SEL(n10938), .F(
        n5758) );
  MUX U12961 ( .IN0(data_mem_out_wire[1995]), .IN1(n9781), .SEL(n10938), .F(
        n5757) );
  IV U12962 ( .A(n10939), .Z(n10938) );
  MUX U12963 ( .IN0(n9783), .IN1(data_mem_out_wire[1994]), .SEL(n10939), .F(
        n5756) );
  MUX U12964 ( .IN0(n9784), .IN1(data_mem_out_wire[1993]), .SEL(n10939), .F(
        n5755) );
  MUX U12965 ( .IN0(n9785), .IN1(data_mem_out_wire[1992]), .SEL(n10939), .F(
        n5754) );
  AND U12966 ( .A(n10940), .B(n10941), .Z(n10939) );
  OR U12967 ( .A(n9788), .B(n10933), .Z(n10941) );
  MUX U12968 ( .IN0(data_mem_out_wire[1991]), .IN1(data_in[7]), .SEL(n10942), 
        .F(n5753) );
  MUX U12969 ( .IN0(data_mem_out_wire[1990]), .IN1(data_in[6]), .SEL(n10942), 
        .F(n5752) );
  MUX U12970 ( .IN0(data_mem_out_wire[1989]), .IN1(data_in[5]), .SEL(n10942), 
        .F(n5751) );
  MUX U12971 ( .IN0(data_mem_out_wire[1988]), .IN1(data_in[4]), .SEL(n10942), 
        .F(n5750) );
  MUX U12972 ( .IN0(data_mem_out_wire[1987]), .IN1(data_in[3]), .SEL(n10942), 
        .F(n5749) );
  IV U12973 ( .A(n10943), .Z(n10942) );
  MUX U12974 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[1986]), .SEL(n10943), 
        .F(n5748) );
  MUX U12975 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[1985]), .SEL(n10943), 
        .F(n5747) );
  MUX U12976 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[1984]), .SEL(n10943), 
        .F(n5746) );
  AND U12977 ( .A(n10940), .B(n10944), .Z(n10943) );
  NANDN U12978 ( .A(n10933), .B(n9792), .Z(n10944) );
  AND U12979 ( .A(n10945), .B(n10930), .Z(n10940) );
  NANDN U12980 ( .A(n10933), .B(n9796), .Z(n10930) );
  NANDN U12981 ( .A(n10933), .B(n9818), .Z(n10945) );
  NANDN U12982 ( .A(n10832), .B(n9919), .Z(n10933) );
  AND U12983 ( .A(n10871), .B(N39), .Z(n9919) );
  AND U12984 ( .A(N38), .B(n10927), .Z(n10871) );
  IV U12985 ( .A(N37), .Z(n10927) );
  MUX U12986 ( .IN0(n9746), .IN1(data_mem_out_wire[2047]), .SEL(n10946), .F(
        n5745) );
  NAND U12987 ( .A(n10947), .B(n10948), .Z(n9746) );
  NAND U12988 ( .A(n9796), .B(data_in[31]), .Z(n10948) );
  AND U12989 ( .A(n10949), .B(n10950), .Z(n10947) );
  NAND U12990 ( .A(n9775), .B(data_in[15]), .Z(n10950) );
  MUX U12991 ( .IN0(n9748), .IN1(data_mem_out_wire[2046]), .SEL(n10946), .F(
        n5744) );
  NAND U12992 ( .A(n10951), .B(n10952), .Z(n9748) );
  NAND U12993 ( .A(n9796), .B(data_in[30]), .Z(n10952) );
  AND U12994 ( .A(n10953), .B(n10954), .Z(n10951) );
  NAND U12995 ( .A(n9775), .B(data_in[14]), .Z(n10954) );
  MUX U12996 ( .IN0(n9749), .IN1(data_mem_out_wire[2045]), .SEL(n10946), .F(
        n5743) );
  NAND U12997 ( .A(n10955), .B(n10956), .Z(n9749) );
  NAND U12998 ( .A(n9796), .B(data_in[29]), .Z(n10956) );
  AND U12999 ( .A(n10957), .B(n10958), .Z(n10955) );
  NAND U13000 ( .A(n9775), .B(data_in[13]), .Z(n10958) );
  MUX U13001 ( .IN0(n9750), .IN1(data_mem_out_wire[2044]), .SEL(n10946), .F(
        n5742) );
  NAND U13002 ( .A(n10959), .B(n10960), .Z(n9750) );
  NAND U13003 ( .A(n9796), .B(data_in[28]), .Z(n10960) );
  AND U13004 ( .A(n10961), .B(n10962), .Z(n10959) );
  NAND U13005 ( .A(n9775), .B(data_in[12]), .Z(n10962) );
  MUX U13006 ( .IN0(n9751), .IN1(data_mem_out_wire[2043]), .SEL(n10946), .F(
        n5741) );
  NAND U13007 ( .A(n10963), .B(n10964), .Z(n9751) );
  NAND U13008 ( .A(n9796), .B(data_in[27]), .Z(n10964) );
  AND U13009 ( .A(n10965), .B(n10966), .Z(n10963) );
  NAND U13010 ( .A(n9775), .B(data_in[11]), .Z(n10966) );
  MUX U13011 ( .IN0(n9752), .IN1(data_mem_out_wire[2042]), .SEL(n10946), .F(
        n5740) );
  NAND U13012 ( .A(n10967), .B(n10968), .Z(n9752) );
  NAND U13013 ( .A(n9796), .B(data_in[26]), .Z(n10968) );
  AND U13014 ( .A(n10969), .B(n10970), .Z(n10967) );
  NAND U13015 ( .A(n9775), .B(data_in[10]), .Z(n10970) );
  MUX U13016 ( .IN0(n9753), .IN1(data_mem_out_wire[2041]), .SEL(n10946), .F(
        n5739) );
  NAND U13017 ( .A(n10971), .B(n10972), .Z(n9753) );
  NAND U13018 ( .A(n9796), .B(data_in[25]), .Z(n10972) );
  AND U13019 ( .A(n10973), .B(n10974), .Z(n10971) );
  NAND U13020 ( .A(n9775), .B(data_in[9]), .Z(n10974) );
  MUX U13021 ( .IN0(n9754), .IN1(data_mem_out_wire[2040]), .SEL(n10946), .F(
        n5738) );
  ANDN U13022 ( .B(n10975), .A(n10976), .Z(n10946) );
  ANDN U13023 ( .B(n10977), .A(n10978), .Z(n10975) );
  NANDN U13024 ( .A(n9760), .B(n10979), .Z(n10977) );
  NANDN U13025 ( .A(n9844), .B(n9857), .Z(n9760) );
  NAND U13026 ( .A(n10980), .B(n10981), .Z(n9754) );
  NAND U13027 ( .A(n9796), .B(data_in[24]), .Z(n10981) );
  AND U13028 ( .A(n10982), .B(n10983), .Z(n10980) );
  NAND U13029 ( .A(n9775), .B(data_in[8]), .Z(n10983) );
  MUX U13030 ( .IN0(data_mem_out_wire[2039]), .IN1(n9761), .SEL(n10984), .F(
        n5737) );
  NAND U13031 ( .A(n10985), .B(n10986), .Z(n9761) );
  NAND U13032 ( .A(n10987), .B(data_in[7]), .Z(n10986) );
  NAND U13033 ( .A(n9796), .B(data_in[23]), .Z(n10985) );
  MUX U13034 ( .IN0(data_mem_out_wire[2038]), .IN1(n9763), .SEL(n10984), .F(
        n5736) );
  NAND U13035 ( .A(n10988), .B(n10989), .Z(n9763) );
  NAND U13036 ( .A(n10987), .B(data_in[6]), .Z(n10989) );
  NAND U13037 ( .A(n9796), .B(data_in[22]), .Z(n10988) );
  MUX U13038 ( .IN0(data_mem_out_wire[2037]), .IN1(n9764), .SEL(n10984), .F(
        n5735) );
  NAND U13039 ( .A(n10990), .B(n10991), .Z(n9764) );
  NAND U13040 ( .A(n10987), .B(data_in[5]), .Z(n10991) );
  NAND U13041 ( .A(n9796), .B(data_in[21]), .Z(n10990) );
  MUX U13042 ( .IN0(data_mem_out_wire[2036]), .IN1(n9765), .SEL(n10984), .F(
        n5734) );
  NAND U13043 ( .A(n10992), .B(n10993), .Z(n9765) );
  NAND U13044 ( .A(n10987), .B(data_in[4]), .Z(n10993) );
  NAND U13045 ( .A(n9796), .B(data_in[20]), .Z(n10992) );
  MUX U13046 ( .IN0(data_mem_out_wire[2035]), .IN1(n9766), .SEL(n10984), .F(
        n5733) );
  IV U13047 ( .A(n10994), .Z(n10984) );
  NAND U13048 ( .A(n10995), .B(n10996), .Z(n9766) );
  NAND U13049 ( .A(n10987), .B(data_in[3]), .Z(n10996) );
  NAND U13050 ( .A(n9796), .B(data_in[19]), .Z(n10995) );
  MUX U13051 ( .IN0(n9768), .IN1(data_mem_out_wire[2034]), .SEL(n10994), .F(
        n5732) );
  NAND U13052 ( .A(n10997), .B(n10998), .Z(n9768) );
  NAND U13053 ( .A(n10987), .B(data_in[2]), .Z(n10998) );
  NAND U13054 ( .A(n9796), .B(data_in[18]), .Z(n10997) );
  MUX U13055 ( .IN0(n9769), .IN1(data_mem_out_wire[2033]), .SEL(n10994), .F(
        n5731) );
  NAND U13056 ( .A(n10999), .B(n11000), .Z(n9769) );
  NAND U13057 ( .A(n10987), .B(data_in[1]), .Z(n11000) );
  NAND U13058 ( .A(n9796), .B(data_in[17]), .Z(n10999) );
  MUX U13059 ( .IN0(n9770), .IN1(data_mem_out_wire[2032]), .SEL(n10994), .F(
        n5730) );
  AND U13060 ( .A(n11001), .B(n11002), .Z(n10994) );
  NANDN U13061 ( .A(n9773), .B(n10979), .Z(n11002) );
  NANDN U13062 ( .A(n9850), .B(n9857), .Z(n9773) );
  NOR U13063 ( .A(n10976), .B(n10978), .Z(n11001) );
  AND U13064 ( .A(n9809), .B(n10979), .Z(n10978) );
  AND U13065 ( .A(n9775), .B(addr[1]), .Z(n9809) );
  NAND U13066 ( .A(n11003), .B(n11004), .Z(n9770) );
  NAND U13067 ( .A(data_in[0]), .B(n10987), .Z(n11004) );
  OR U13068 ( .A(n9857), .B(n9775), .Z(n10987) );
  NAND U13069 ( .A(n9796), .B(data_in[16]), .Z(n11003) );
  MUX U13070 ( .IN0(data_mem_out_wire[2031]), .IN1(n9776), .SEL(n11005), .F(
        n5729) );
  NAND U13071 ( .A(n10949), .B(n11006), .Z(n9776) );
  NAND U13072 ( .A(n11007), .B(data_in[15]), .Z(n11006) );
  NAND U13073 ( .A(n9857), .B(data_in[7]), .Z(n10949) );
  MUX U13074 ( .IN0(data_mem_out_wire[2030]), .IN1(n9778), .SEL(n11005), .F(
        n5728) );
  NAND U13075 ( .A(n10953), .B(n11008), .Z(n9778) );
  NAND U13076 ( .A(n11007), .B(data_in[14]), .Z(n11008) );
  NAND U13077 ( .A(n9857), .B(data_in[6]), .Z(n10953) );
  MUX U13078 ( .IN0(data_mem_out_wire[2029]), .IN1(n9779), .SEL(n11005), .F(
        n5727) );
  NAND U13079 ( .A(n10957), .B(n11009), .Z(n9779) );
  NAND U13080 ( .A(n11007), .B(data_in[13]), .Z(n11009) );
  NAND U13081 ( .A(n9857), .B(data_in[5]), .Z(n10957) );
  MUX U13082 ( .IN0(data_mem_out_wire[2028]), .IN1(n9780), .SEL(n11005), .F(
        n5726) );
  NAND U13083 ( .A(n10961), .B(n11010), .Z(n9780) );
  NAND U13084 ( .A(n11007), .B(data_in[12]), .Z(n11010) );
  NAND U13085 ( .A(n9857), .B(data_in[4]), .Z(n10961) );
  MUX U13086 ( .IN0(data_mem_out_wire[2027]), .IN1(n9781), .SEL(n11005), .F(
        n5725) );
  IV U13087 ( .A(n11011), .Z(n11005) );
  NAND U13088 ( .A(n10965), .B(n11012), .Z(n9781) );
  NAND U13089 ( .A(n11007), .B(data_in[11]), .Z(n11012) );
  NAND U13090 ( .A(n9857), .B(data_in[3]), .Z(n10965) );
  MUX U13091 ( .IN0(n9783), .IN1(data_mem_out_wire[2026]), .SEL(n11011), .F(
        n5724) );
  NAND U13092 ( .A(n10969), .B(n11013), .Z(n9783) );
  NAND U13093 ( .A(n11007), .B(data_in[10]), .Z(n11013) );
  NAND U13094 ( .A(n9857), .B(data_in[2]), .Z(n10969) );
  MUX U13095 ( .IN0(n9784), .IN1(data_mem_out_wire[2025]), .SEL(n11011), .F(
        n5723) );
  NAND U13096 ( .A(n10973), .B(n11014), .Z(n9784) );
  NAND U13097 ( .A(n11007), .B(data_in[9]), .Z(n11014) );
  NAND U13098 ( .A(n9857), .B(data_in[1]), .Z(n10973) );
  MUX U13099 ( .IN0(n9785), .IN1(data_mem_out_wire[2024]), .SEL(n11011), .F(
        n5722) );
  AND U13100 ( .A(n11015), .B(n11016), .Z(n11011) );
  NANDN U13101 ( .A(n9788), .B(n10979), .Z(n11016) );
  NAND U13102 ( .A(n9857), .B(n9856), .Z(n9788) );
  NAND U13103 ( .A(n10982), .B(n11017), .Z(n9785) );
  NAND U13104 ( .A(data_in[8]), .B(n11007), .Z(n11017) );
  OR U13105 ( .A(n9796), .B(n9775), .Z(n11007) );
  NAND U13106 ( .A(n9857), .B(data_in[0]), .Z(n10982) );
  MUX U13107 ( .IN0(data_mem_out_wire[2023]), .IN1(data_in[7]), .SEL(n11018), 
        .F(n5721) );
  MUX U13108 ( .IN0(data_mem_out_wire[2022]), .IN1(data_in[6]), .SEL(n11018), 
        .F(n5720) );
  MUX U13109 ( .IN0(data_mem_out_wire[2021]), .IN1(data_in[5]), .SEL(n11018), 
        .F(n5719) );
  MUX U13110 ( .IN0(data_mem_out_wire[2020]), .IN1(data_in[4]), .SEL(n11018), 
        .F(n5718) );
  MUX U13111 ( .IN0(data_mem_out_wire[2019]), .IN1(data_in[3]), .SEL(n11018), 
        .F(n5717) );
  IV U13112 ( .A(n11019), .Z(n11018) );
  MUX U13113 ( .IN0(data_in[2]), .IN1(data_mem_out_wire[2018]), .SEL(n11019), 
        .F(n5716) );
  MUX U13114 ( .IN0(data_in[1]), .IN1(data_mem_out_wire[2017]), .SEL(n11019), 
        .F(n5715) );
  MUX U13115 ( .IN0(data_in[0]), .IN1(data_mem_out_wire[2016]), .SEL(n11019), 
        .F(n5714) );
  AND U13116 ( .A(n11015), .B(n11020), .Z(n11019) );
  NAND U13117 ( .A(n10979), .B(n9792), .Z(n11020) );
  ANDN U13118 ( .B(n9857), .A(n11021), .Z(n9792) );
  AND U13119 ( .A(n11022), .B(n11023), .Z(n9857) );
  AND U13120 ( .A(mem_source[0]), .B(n11024), .Z(n11022) );
  NOR U13121 ( .A(n10976), .B(n11025), .Z(n11015) );
  AND U13122 ( .A(n9818), .B(n10979), .Z(n11025) );
  IV U13123 ( .A(n11026), .Z(n10979) );
  AND U13124 ( .A(n9775), .B(n9795), .Z(n9818) );
  AND U13125 ( .A(n11027), .B(n11028), .Z(n9775) );
  NOR U13126 ( .A(mem_source[1]), .B(mem_source[2]), .Z(n11028) );
  AND U13127 ( .A(mem_source[0]), .B(mem_source[3]), .Z(n11027) );
  ANDN U13128 ( .B(n9796), .A(n11026), .Z(n10976) );
  NANDN U13129 ( .A(n10832), .B(n9938), .Z(n11026) );
  AND U13130 ( .A(n10890), .B(N39), .Z(n9938) );
  AND U13131 ( .A(N38), .B(N37), .Z(n10890) );
  NAND U13132 ( .A(n10377), .B(N42), .Z(n10832) );
  AND U13133 ( .A(N40), .B(N41), .Z(n10377) );
  AND U13134 ( .A(n11029), .B(n11030), .Z(n9796) );
  AND U13135 ( .A(mem_source[0]), .B(mem_source[2]), .Z(n11029) );
  ANDN U13136 ( .B(n11031), .A(mem_source[0]), .Z(data_out[9]) );
  NAND U13137 ( .A(n11032), .B(n11033), .Z(n11031) );
  AND U13138 ( .A(n11034), .B(n11035), .Z(n11033) );
  NANDN U13139 ( .A(n11036), .B(N736), .Z(n11034) );
  AND U13140 ( .A(n11037), .B(n11038), .Z(n11032) );
  NAND U13141 ( .A(n11039), .B(n11040), .Z(n11038) );
  NAND U13142 ( .A(n11039), .B(n11041), .Z(n11037) );
  MUX U13143 ( .IN0(N736), .IN1(N720), .SEL(addr[1]), .F(n11039) );
  ANDN U13144 ( .B(n11042), .A(mem_source[0]), .Z(data_out[8]) );
  NAND U13145 ( .A(n11043), .B(n11044), .Z(n11042) );
  AND U13146 ( .A(n11045), .B(n11035), .Z(n11044) );
  NANDN U13147 ( .A(n11036), .B(N737), .Z(n11045) );
  AND U13148 ( .A(n11046), .B(n11047), .Z(n11043) );
  NAND U13149 ( .A(n11048), .B(n11040), .Z(n11047) );
  NAND U13150 ( .A(n11048), .B(n11041), .Z(n11046) );
  MUX U13151 ( .IN0(N737), .IN1(N721), .SEL(addr[1]), .F(n11048) );
  ANDN U13152 ( .B(n11049), .A(mem_source[0]), .Z(data_out[7]) );
  NAND U13153 ( .A(n11050), .B(n11051), .Z(n11049) );
  AND U13154 ( .A(n11052), .B(n11053), .Z(n11051) );
  NANDN U13155 ( .A(n11054), .B(n11055), .Z(n11053) );
  AND U13156 ( .A(n11056), .B(n11057), .Z(n11052) );
  NANDN U13157 ( .A(n11036), .B(N738), .Z(n11057) );
  NAND U13158 ( .A(n11058), .B(n11040), .Z(n11056) );
  AND U13159 ( .A(n11059), .B(n11060), .Z(n11050) );
  OR U13160 ( .A(n11061), .B(n11054), .Z(n11060) );
  AND U13161 ( .A(n11062), .B(n11063), .Z(n11054) );
  AND U13162 ( .A(n11064), .B(n11065), .Z(n11063) );
  NANDN U13163 ( .A(n11021), .B(N738), .Z(n11065) );
  NAND U13164 ( .A(N730), .B(n9856), .Z(n11064) );
  AND U13165 ( .A(n11066), .B(n11067), .Z(n11062) );
  NANDN U13166 ( .A(n9850), .B(N722), .Z(n11067) );
  NANDN U13167 ( .A(n9844), .B(N714), .Z(n11066) );
  NAND U13168 ( .A(n11058), .B(n11041), .Z(n11059) );
  MUX U13169 ( .IN0(N738), .IN1(N722), .SEL(addr[1]), .F(n11058) );
  ANDN U13170 ( .B(n11068), .A(mem_source[0]), .Z(data_out[6]) );
  NAND U13171 ( .A(n11069), .B(n11070), .Z(n11068) );
  AND U13172 ( .A(n11071), .B(n11072), .Z(n11070) );
  NANDN U13173 ( .A(n11073), .B(n11055), .Z(n11072) );
  AND U13174 ( .A(n11074), .B(n11075), .Z(n11071) );
  NANDN U13175 ( .A(n11036), .B(N739), .Z(n11075) );
  NAND U13176 ( .A(n11076), .B(n11040), .Z(n11074) );
  AND U13177 ( .A(n11077), .B(n11078), .Z(n11069) );
  OR U13178 ( .A(n11061), .B(n11073), .Z(n11078) );
  AND U13179 ( .A(n11079), .B(n11080), .Z(n11073) );
  AND U13180 ( .A(n11081), .B(n11082), .Z(n11080) );
  NANDN U13181 ( .A(n11021), .B(N739), .Z(n11082) );
  NAND U13182 ( .A(n9856), .B(N731), .Z(n11081) );
  AND U13183 ( .A(n11083), .B(n11084), .Z(n11079) );
  NANDN U13184 ( .A(n9850), .B(N723), .Z(n11084) );
  NANDN U13185 ( .A(n9844), .B(N715), .Z(n11083) );
  NAND U13186 ( .A(n11076), .B(n11041), .Z(n11077) );
  MUX U13187 ( .IN0(N739), .IN1(N723), .SEL(addr[1]), .F(n11076) );
  ANDN U13188 ( .B(n11085), .A(mem_source[0]), .Z(data_out[5]) );
  NAND U13189 ( .A(n11086), .B(n11087), .Z(n11085) );
  AND U13190 ( .A(n11088), .B(n11089), .Z(n11087) );
  NANDN U13191 ( .A(n11090), .B(n11055), .Z(n11089) );
  AND U13192 ( .A(n11091), .B(n11092), .Z(n11088) );
  NANDN U13193 ( .A(n11036), .B(N740), .Z(n11092) );
  NAND U13194 ( .A(n11093), .B(n11040), .Z(n11091) );
  AND U13195 ( .A(n11094), .B(n11095), .Z(n11086) );
  OR U13196 ( .A(n11061), .B(n11090), .Z(n11095) );
  AND U13197 ( .A(n11096), .B(n11097), .Z(n11090) );
  AND U13198 ( .A(n11098), .B(n11099), .Z(n11097) );
  NANDN U13199 ( .A(n11021), .B(N740), .Z(n11099) );
  NAND U13200 ( .A(n9856), .B(N732), .Z(n11098) );
  AND U13201 ( .A(n11100), .B(n11101), .Z(n11096) );
  NANDN U13202 ( .A(n9850), .B(N724), .Z(n11101) );
  NANDN U13203 ( .A(n9844), .B(N716), .Z(n11100) );
  NAND U13204 ( .A(n11093), .B(n11041), .Z(n11094) );
  MUX U13205 ( .IN0(N740), .IN1(N724), .SEL(addr[1]), .F(n11093) );
  ANDN U13206 ( .B(n11102), .A(mem_source[0]), .Z(data_out[4]) );
  NAND U13207 ( .A(n11103), .B(n11104), .Z(n11102) );
  AND U13208 ( .A(n11105), .B(n11106), .Z(n11104) );
  NANDN U13209 ( .A(n11107), .B(n11055), .Z(n11106) );
  AND U13210 ( .A(n11108), .B(n11109), .Z(n11105) );
  NANDN U13211 ( .A(n11036), .B(N741), .Z(n11109) );
  NAND U13212 ( .A(n11110), .B(n11040), .Z(n11108) );
  AND U13213 ( .A(n11111), .B(n11112), .Z(n11103) );
  OR U13214 ( .A(n11061), .B(n11107), .Z(n11112) );
  AND U13215 ( .A(n11113), .B(n11114), .Z(n11107) );
  AND U13216 ( .A(n11115), .B(n11116), .Z(n11114) );
  NANDN U13217 ( .A(n11021), .B(N741), .Z(n11116) );
  NAND U13218 ( .A(n9856), .B(N733), .Z(n11115) );
  AND U13219 ( .A(n11117), .B(n11118), .Z(n11113) );
  NANDN U13220 ( .A(n9850), .B(N725), .Z(n11118) );
  NANDN U13221 ( .A(n9844), .B(N717), .Z(n11117) );
  NAND U13222 ( .A(n11110), .B(n11041), .Z(n11111) );
  MUX U13223 ( .IN0(N741), .IN1(N725), .SEL(addr[1]), .F(n11110) );
  ANDN U13224 ( .B(n11119), .A(mem_source[0]), .Z(data_out[3]) );
  NAND U13225 ( .A(n11120), .B(n11121), .Z(n11119) );
  AND U13226 ( .A(n11122), .B(n11123), .Z(n11121) );
  NANDN U13227 ( .A(n11124), .B(n11055), .Z(n11123) );
  AND U13228 ( .A(n11125), .B(n11126), .Z(n11122) );
  NANDN U13229 ( .A(n11036), .B(N742), .Z(n11126) );
  NAND U13230 ( .A(n11127), .B(n11040), .Z(n11125) );
  AND U13231 ( .A(n11128), .B(n11129), .Z(n11120) );
  OR U13232 ( .A(n11061), .B(n11124), .Z(n11129) );
  AND U13233 ( .A(n11130), .B(n11131), .Z(n11124) );
  AND U13234 ( .A(n11132), .B(n11133), .Z(n11131) );
  NANDN U13235 ( .A(n11021), .B(N742), .Z(n11133) );
  NAND U13236 ( .A(n9856), .B(N734), .Z(n11132) );
  AND U13237 ( .A(n11134), .B(n11135), .Z(n11130) );
  NANDN U13238 ( .A(n9850), .B(N726), .Z(n11135) );
  NANDN U13239 ( .A(n9844), .B(N718), .Z(n11134) );
  NAND U13240 ( .A(n11127), .B(n11041), .Z(n11128) );
  MUX U13241 ( .IN0(N742), .IN1(N726), .SEL(addr[1]), .F(n11127) );
  ANDN U13242 ( .B(n11136), .A(mem_source[0]), .Z(data_out[31]) );
  NAND U13243 ( .A(n11137), .B(n11138), .Z(n11136) );
  NANDN U13244 ( .A(n11036), .B(N714), .Z(n11137) );
  ANDN U13245 ( .B(n11139), .A(mem_source[0]), .Z(data_out[30]) );
  NAND U13246 ( .A(n11140), .B(n11138), .Z(n11139) );
  NANDN U13247 ( .A(n11036), .B(N715), .Z(n11140) );
  ANDN U13248 ( .B(n11141), .A(mem_source[0]), .Z(data_out[2]) );
  NAND U13249 ( .A(n11142), .B(n11143), .Z(n11141) );
  AND U13250 ( .A(n11144), .B(n11145), .Z(n11143) );
  NANDN U13251 ( .A(n11146), .B(n11055), .Z(n11145) );
  AND U13252 ( .A(n11147), .B(n11148), .Z(n11144) );
  NANDN U13253 ( .A(n11036), .B(N743), .Z(n11148) );
  NAND U13254 ( .A(n11149), .B(n11040), .Z(n11147) );
  AND U13255 ( .A(n11150), .B(n11151), .Z(n11142) );
  OR U13256 ( .A(n11061), .B(n11146), .Z(n11151) );
  AND U13257 ( .A(n11152), .B(n11153), .Z(n11146) );
  AND U13258 ( .A(n11154), .B(n11155), .Z(n11153) );
  NANDN U13259 ( .A(n11021), .B(N743), .Z(n11155) );
  NAND U13260 ( .A(n9856), .B(N735), .Z(n11154) );
  AND U13261 ( .A(n11156), .B(n11157), .Z(n11152) );
  NANDN U13262 ( .A(n9850), .B(N727), .Z(n11157) );
  NANDN U13263 ( .A(n9844), .B(N719), .Z(n11156) );
  NAND U13264 ( .A(n11149), .B(n11041), .Z(n11150) );
  MUX U13265 ( .IN0(N743), .IN1(N727), .SEL(addr[1]), .F(n11149) );
  ANDN U13266 ( .B(n11158), .A(mem_source[0]), .Z(data_out[29]) );
  NAND U13267 ( .A(n11159), .B(n11138), .Z(n11158) );
  NANDN U13268 ( .A(n11036), .B(N716), .Z(n11159) );
  ANDN U13269 ( .B(n11160), .A(mem_source[0]), .Z(data_out[28]) );
  NAND U13270 ( .A(n11161), .B(n11138), .Z(n11160) );
  NANDN U13271 ( .A(n11036), .B(N717), .Z(n11161) );
  ANDN U13272 ( .B(n11162), .A(mem_source[0]), .Z(data_out[27]) );
  NAND U13273 ( .A(n11163), .B(n11138), .Z(n11162) );
  NANDN U13274 ( .A(n11036), .B(N718), .Z(n11163) );
  ANDN U13275 ( .B(n11164), .A(mem_source[0]), .Z(data_out[26]) );
  NAND U13276 ( .A(n11165), .B(n11138), .Z(n11164) );
  NANDN U13277 ( .A(n11036), .B(N719), .Z(n11165) );
  ANDN U13278 ( .B(n11166), .A(mem_source[0]), .Z(data_out[25]) );
  NAND U13279 ( .A(n11167), .B(n11138), .Z(n11166) );
  NANDN U13280 ( .A(n11036), .B(N720), .Z(n11167) );
  ANDN U13281 ( .B(n11168), .A(mem_source[0]), .Z(data_out[24]) );
  NAND U13282 ( .A(n11169), .B(n11138), .Z(n11168) );
  NANDN U13283 ( .A(n11036), .B(N721), .Z(n11169) );
  ANDN U13284 ( .B(n11170), .A(mem_source[0]), .Z(data_out[23]) );
  NAND U13285 ( .A(n11171), .B(n11138), .Z(n11170) );
  NANDN U13286 ( .A(n11036), .B(N722), .Z(n11171) );
  ANDN U13287 ( .B(n11172), .A(mem_source[0]), .Z(data_out[22]) );
  NAND U13288 ( .A(n11173), .B(n11138), .Z(n11172) );
  NANDN U13289 ( .A(n11036), .B(N723), .Z(n11173) );
  ANDN U13290 ( .B(n11174), .A(mem_source[0]), .Z(data_out[21]) );
  NAND U13291 ( .A(n11175), .B(n11138), .Z(n11174) );
  NANDN U13292 ( .A(n11036), .B(N724), .Z(n11175) );
  ANDN U13293 ( .B(n11176), .A(mem_source[0]), .Z(data_out[20]) );
  NAND U13294 ( .A(n11177), .B(n11138), .Z(n11176) );
  NANDN U13295 ( .A(n11036), .B(N725), .Z(n11177) );
  ANDN U13296 ( .B(n11178), .A(mem_source[0]), .Z(data_out[1]) );
  NAND U13297 ( .A(n11179), .B(n11180), .Z(n11178) );
  AND U13298 ( .A(n11181), .B(n11182), .Z(n11180) );
  NANDN U13299 ( .A(n11183), .B(n11055), .Z(n11182) );
  AND U13300 ( .A(n11184), .B(n11185), .Z(n11181) );
  NANDN U13301 ( .A(n11036), .B(N744), .Z(n11185) );
  NAND U13302 ( .A(n11186), .B(n11040), .Z(n11184) );
  AND U13303 ( .A(n11187), .B(n11188), .Z(n11179) );
  OR U13304 ( .A(n11183), .B(n11061), .Z(n11188) );
  AND U13305 ( .A(n11189), .B(n11190), .Z(n11183) );
  AND U13306 ( .A(n11191), .B(n11192), .Z(n11190) );
  NANDN U13307 ( .A(n11021), .B(N744), .Z(n11192) );
  NAND U13308 ( .A(n9856), .B(N736), .Z(n11191) );
  AND U13309 ( .A(n11193), .B(n11194), .Z(n11189) );
  NANDN U13310 ( .A(n9850), .B(N728), .Z(n11194) );
  NANDN U13311 ( .A(n9844), .B(N720), .Z(n11193) );
  NAND U13312 ( .A(n11186), .B(n11041), .Z(n11187) );
  MUX U13313 ( .IN0(N744), .IN1(N728), .SEL(addr[1]), .F(n11186) );
  ANDN U13314 ( .B(n11195), .A(mem_source[0]), .Z(data_out[19]) );
  NAND U13315 ( .A(n11196), .B(n11138), .Z(n11195) );
  NANDN U13316 ( .A(n11036), .B(N726), .Z(n11196) );
  ANDN U13317 ( .B(n11197), .A(mem_source[0]), .Z(data_out[18]) );
  NAND U13318 ( .A(n11198), .B(n11138), .Z(n11197) );
  NANDN U13319 ( .A(n11036), .B(N727), .Z(n11198) );
  ANDN U13320 ( .B(n11199), .A(mem_source[0]), .Z(data_out[17]) );
  NAND U13321 ( .A(n11200), .B(n11138), .Z(n11199) );
  NANDN U13322 ( .A(n11036), .B(N728), .Z(n11200) );
  ANDN U13323 ( .B(n11201), .A(mem_source[0]), .Z(data_out[16]) );
  NAND U13324 ( .A(n11202), .B(n11138), .Z(n11201) );
  ANDN U13325 ( .B(n11203), .A(n11204), .Z(n11138) );
  IV U13326 ( .A(n11035), .Z(n11204) );
  NAND U13327 ( .A(n11205), .B(n11040), .Z(n11203) );
  NANDN U13328 ( .A(n11206), .B(n11207), .Z(n11205) );
  NANDN U13329 ( .A(n11036), .B(N729), .Z(n11202) );
  ANDN U13330 ( .B(n11208), .A(mem_source[0]), .Z(data_out[15]) );
  NAND U13331 ( .A(n11209), .B(n11210), .Z(n11208) );
  AND U13332 ( .A(n11211), .B(n11035), .Z(n11210) );
  NANDN U13333 ( .A(n11036), .B(N730), .Z(n11211) );
  AND U13334 ( .A(n11212), .B(n11213), .Z(n11209) );
  NANDN U13335 ( .A(n11214), .B(n11040), .Z(n11213) );
  NANDN U13336 ( .A(n11214), .B(n11041), .Z(n11212) );
  ANDN U13337 ( .B(n11215), .A(n11206), .Z(n11214) );
  ANDN U13338 ( .B(n9795), .A(n11216), .Z(n11206) );
  IV U13339 ( .A(N730), .Z(n11216) );
  NAND U13340 ( .A(addr[1]), .B(N714), .Z(n11215) );
  ANDN U13341 ( .B(n11217), .A(mem_source[0]), .Z(data_out[14]) );
  NAND U13342 ( .A(n11218), .B(n11219), .Z(n11217) );
  AND U13343 ( .A(n11220), .B(n11035), .Z(n11219) );
  NANDN U13344 ( .A(n11036), .B(N731), .Z(n11220) );
  AND U13345 ( .A(n11221), .B(n11222), .Z(n11218) );
  NAND U13346 ( .A(n11040), .B(n11223), .Z(n11222) );
  NAND U13347 ( .A(n11223), .B(n11041), .Z(n11221) );
  MUX U13348 ( .IN0(N731), .IN1(N715), .SEL(addr[1]), .F(n11223) );
  ANDN U13349 ( .B(n11224), .A(mem_source[0]), .Z(data_out[13]) );
  NAND U13350 ( .A(n11225), .B(n11226), .Z(n11224) );
  AND U13351 ( .A(n11227), .B(n11035), .Z(n11226) );
  NANDN U13352 ( .A(n11036), .B(N732), .Z(n11227) );
  AND U13353 ( .A(n11228), .B(n11229), .Z(n11225) );
  NAND U13354 ( .A(n11040), .B(n11230), .Z(n11229) );
  NAND U13355 ( .A(n11230), .B(n11041), .Z(n11228) );
  MUX U13356 ( .IN0(N732), .IN1(N716), .SEL(addr[1]), .F(n11230) );
  ANDN U13357 ( .B(n11231), .A(mem_source[0]), .Z(data_out[12]) );
  NAND U13358 ( .A(n11232), .B(n11233), .Z(n11231) );
  AND U13359 ( .A(n11234), .B(n11035), .Z(n11233) );
  NANDN U13360 ( .A(n11036), .B(N733), .Z(n11234) );
  AND U13361 ( .A(n11235), .B(n11236), .Z(n11232) );
  NAND U13362 ( .A(n11040), .B(n11237), .Z(n11236) );
  NAND U13363 ( .A(n11237), .B(n11041), .Z(n11235) );
  MUX U13364 ( .IN0(N733), .IN1(N717), .SEL(addr[1]), .F(n11237) );
  ANDN U13365 ( .B(n11238), .A(mem_source[0]), .Z(data_out[11]) );
  NAND U13366 ( .A(n11239), .B(n11240), .Z(n11238) );
  AND U13367 ( .A(n11241), .B(n11035), .Z(n11240) );
  NANDN U13368 ( .A(n11036), .B(N734), .Z(n11241) );
  AND U13369 ( .A(n11242), .B(n11243), .Z(n11239) );
  NAND U13370 ( .A(n11040), .B(n11244), .Z(n11243) );
  NAND U13371 ( .A(n11244), .B(n11041), .Z(n11242) );
  MUX U13372 ( .IN0(N734), .IN1(N718), .SEL(addr[1]), .F(n11244) );
  ANDN U13373 ( .B(n11245), .A(mem_source[0]), .Z(data_out[10]) );
  NAND U13374 ( .A(n11246), .B(n11247), .Z(n11245) );
  AND U13375 ( .A(n11248), .B(n11035), .Z(n11247) );
  NAND U13376 ( .A(n11055), .B(N738), .Z(n11035) );
  NANDN U13377 ( .A(n11036), .B(N735), .Z(n11248) );
  AND U13378 ( .A(n11249), .B(n11250), .Z(n11246) );
  NAND U13379 ( .A(n11040), .B(n11251), .Z(n11250) );
  NAND U13380 ( .A(n11251), .B(n11041), .Z(n11249) );
  MUX U13381 ( .IN0(N735), .IN1(N719), .SEL(addr[1]), .F(n11251) );
  ANDN U13382 ( .B(n11252), .A(mem_source[0]), .Z(data_out[0]) );
  NAND U13383 ( .A(n11253), .B(n11254), .Z(n11252) );
  AND U13384 ( .A(n11255), .B(n11256), .Z(n11254) );
  NANDN U13385 ( .A(n11257), .B(n11055), .Z(n11256) );
  AND U13386 ( .A(n11023), .B(mem_source[1]), .Z(n11055) );
  ANDN U13387 ( .B(mem_source[2]), .A(n11258), .Z(n11023) );
  AND U13388 ( .A(n11259), .B(n11260), .Z(n11255) );
  NANDN U13389 ( .A(n11036), .B(N745), .Z(n11260) );
  NAND U13390 ( .A(n11030), .B(mem_source[2]), .Z(n11036) );
  ANDN U13391 ( .B(n11258), .A(mem_source[1]), .Z(n11030) );
  NAND U13392 ( .A(n11261), .B(n11040), .Z(n11259) );
  AND U13393 ( .A(n11262), .B(mem_source[1]), .Z(n11040) );
  AND U13394 ( .A(n11263), .B(n11264), .Z(n11253) );
  OR U13395 ( .A(n11257), .B(n11061), .Z(n11264) );
  NAND U13396 ( .A(n11265), .B(mem_source[2]), .Z(n11061) );
  AND U13397 ( .A(n11024), .B(mem_source[3]), .Z(n11265) );
  IV U13398 ( .A(mem_source[1]), .Z(n11024) );
  AND U13399 ( .A(n11266), .B(n11267), .Z(n11257) );
  AND U13400 ( .A(n11268), .B(n11269), .Z(n11267) );
  NANDN U13401 ( .A(n11021), .B(N745), .Z(n11269) );
  NANDN U13402 ( .A(addr[0]), .B(n9795), .Z(n11021) );
  NAND U13403 ( .A(N737), .B(n9856), .Z(n11268) );
  AND U13404 ( .A(addr[0]), .B(n9795), .Z(n9856) );
  AND U13405 ( .A(n11270), .B(n11271), .Z(n11266) );
  NANDN U13406 ( .A(n9850), .B(N729), .Z(n11271) );
  NANDN U13407 ( .A(addr[0]), .B(addr[1]), .Z(n9850) );
  NANDN U13408 ( .A(n9844), .B(N721), .Z(n11270) );
  NAND U13409 ( .A(addr[1]), .B(addr[0]), .Z(n9844) );
  NAND U13410 ( .A(n11261), .B(n11041), .Z(n11263) );
  ANDN U13411 ( .B(n11262), .A(mem_source[1]), .Z(n11041) );
  NOR U13412 ( .A(n11258), .B(mem_source[2]), .Z(n11262) );
  IV U13413 ( .A(mem_source[3]), .Z(n11258) );
  NAND U13414 ( .A(n11272), .B(n11207), .Z(n11261) );
  NAND U13415 ( .A(addr[1]), .B(N729), .Z(n11207) );
  NAND U13416 ( .A(n9795), .B(N745), .Z(n11272) );
  IV U13417 ( .A(addr[1]), .Z(n9795) );
endmodule

