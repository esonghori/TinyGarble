
module sum_N1024_CC64 ( clk, rst, a, b, c );
  input [15:0] a;
  input [15:0] b;
  output [15:0] c;
  input clk, rst;
  wire   N34, N35, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232;
  wire   [1:0] carry_on;

  DFF \carry_on_reg[1]  ( .D(N35), .CLK(clk), .RST(rst), .Q(carry_on[1]) );
  DFF \carry_on_reg[0]  ( .D(N34), .CLK(clk), .RST(rst), .Q(carry_on[0]) );
  DFF \rc_reg[15]  ( .D(n64), .CLK(clk), .RST(1'b0), .Q(c[15]) );
  DFF \rc_reg[14]  ( .D(n63), .CLK(clk), .RST(1'b0), .Q(c[14]) );
  DFF \rc_reg[13]  ( .D(n62), .CLK(clk), .RST(1'b0), .Q(c[13]) );
  DFF \rc_reg[12]  ( .D(n61), .CLK(clk), .RST(1'b0), .Q(c[12]) );
  DFF \rc_reg[11]  ( .D(n60), .CLK(clk), .RST(1'b0), .Q(c[11]) );
  DFF \rc_reg[10]  ( .D(n59), .CLK(clk), .RST(1'b0), .Q(c[10]) );
  DFF \rc_reg[9]  ( .D(n58), .CLK(clk), .RST(1'b0), .Q(c[9]) );
  DFF \rc_reg[8]  ( .D(n57), .CLK(clk), .RST(1'b0), .Q(c[8]) );
  DFF \rc_reg[7]  ( .D(n56), .CLK(clk), .RST(1'b0), .Q(c[7]) );
  DFF \rc_reg[6]  ( .D(n55), .CLK(clk), .RST(1'b0), .Q(c[6]) );
  DFF \rc_reg[5]  ( .D(n54), .CLK(clk), .RST(1'b0), .Q(c[5]) );
  DFF \rc_reg[4]  ( .D(n53), .CLK(clk), .RST(1'b0), .Q(c[4]) );
  DFF \rc_reg[3]  ( .D(n52), .CLK(clk), .RST(1'b0), .Q(c[3]) );
  DFF \rc_reg[2]  ( .D(n51), .CLK(clk), .RST(1'b0), .Q(c[2]) );
  DFF \rc_reg[1]  ( .D(n50), .CLK(clk), .RST(1'b0), .Q(c[1]) );
  DFF \rc_reg[0]  ( .D(n49), .CLK(clk), .RST(1'b0), .Q(c[0]) );
  NANDN U67 ( .A(n145), .B(n146), .Z(n65) );
  NANDN U68 ( .A(n219), .B(n218), .Z(n66) );
  AND U69 ( .A(n65), .B(n66), .Z(n67) );
  NAND U70 ( .A(n224), .B(n223), .Z(n68) );
  NANDN U71 ( .A(n67), .B(n147), .Z(n69) );
  AND U72 ( .A(n68), .B(n69), .Z(n148) );
  XOR U73 ( .A(n124), .B(n123), .Z(n198) );
  XOR U74 ( .A(n87), .B(n86), .Z(n168) );
  XOR U75 ( .A(n112), .B(n111), .Z(n188) );
  XOR U76 ( .A(n136), .B(n135), .Z(n208) );
  AND U77 ( .A(b[15]), .B(a[15]), .Z(n153) );
  NAND U78 ( .A(a[13]), .B(b[13]), .Z(n147) );
  AND U79 ( .A(a[12]), .B(b[12]), .Z(n145) );
  XNOR U80 ( .A(a[1]), .B(b[1]), .Z(n72) );
  XNOR U81 ( .A(carry_on[1]), .B(n72), .Z(n159) );
  NAND U82 ( .A(a[0]), .B(b[0]), .Z(n71) );
  XOR U83 ( .A(a[0]), .B(b[0]), .Z(n154) );
  NAND U84 ( .A(n154), .B(carry_on[0]), .Z(n70) );
  NAND U85 ( .A(n71), .B(n70), .Z(n158) );
  NAND U86 ( .A(n159), .B(n158), .Z(n74) );
  ANDN U87 ( .B(carry_on[1]), .A(n72), .Z(n75) );
  ANDN U88 ( .B(n74), .A(n75), .Z(n73) );
  NAND U89 ( .A(a[1]), .B(b[1]), .Z(n76) );
  NAND U90 ( .A(n73), .B(n76), .Z(n80) );
  XNOR U91 ( .A(n76), .B(n74), .Z(n78) );
  NAND U92 ( .A(n76), .B(n75), .Z(n77) );
  NAND U93 ( .A(n78), .B(n77), .Z(n164) );
  XNOR U94 ( .A(a[2]), .B(b[2]), .Z(n163) );
  NAND U95 ( .A(n164), .B(n163), .Z(n79) );
  NAND U96 ( .A(n80), .B(n79), .Z(n86) );
  NAND U97 ( .A(a[2]), .B(b[2]), .Z(n87) );
  AND U98 ( .A(n86), .B(n87), .Z(n82) );
  XOR U99 ( .A(a[3]), .B(b[3]), .Z(n169) );
  ANDN U100 ( .B(n168), .A(n169), .Z(n81) );
  OR U101 ( .A(n82), .B(n81), .Z(n83) );
  AND U102 ( .A(a[3]), .B(b[3]), .Z(n85) );
  ANDN U103 ( .B(n83), .A(n85), .Z(n92) );
  NOR U104 ( .A(n87), .B(n86), .Z(n84) );
  XNOR U105 ( .A(n85), .B(n84), .Z(n90) );
  XOR U106 ( .A(n87), .B(n86), .Z(n88) );
  NAND U107 ( .A(n88), .B(n169), .Z(n89) );
  NAND U108 ( .A(n90), .B(n89), .Z(n174) );
  XNOR U109 ( .A(a[4]), .B(b[4]), .Z(n173) );
  NAND U110 ( .A(n174), .B(n173), .Z(n91) );
  NANDN U111 ( .A(n92), .B(n91), .Z(n99) );
  AND U112 ( .A(a[4]), .B(b[4]), .Z(n93) );
  IV U113 ( .A(n93), .Z(n100) );
  AND U114 ( .A(n99), .B(n100), .Z(n95) );
  XOR U115 ( .A(a[5]), .B(b[5]), .Z(n179) );
  XNOR U116 ( .A(n93), .B(n99), .Z(n178) );
  NANDN U117 ( .A(n179), .B(n178), .Z(n94) );
  NANDN U118 ( .A(n95), .B(n94), .Z(n96) );
  AND U119 ( .A(a[5]), .B(b[5]), .Z(n98) );
  ANDN U120 ( .B(n96), .A(n98), .Z(n105) );
  NOR U121 ( .A(n100), .B(n99), .Z(n97) );
  XNOR U122 ( .A(n98), .B(n97), .Z(n103) );
  XOR U123 ( .A(n100), .B(n99), .Z(n101) );
  NAND U124 ( .A(n101), .B(n179), .Z(n102) );
  NAND U125 ( .A(n103), .B(n102), .Z(n184) );
  XNOR U126 ( .A(a[6]), .B(b[6]), .Z(n183) );
  NAND U127 ( .A(n184), .B(n183), .Z(n104) );
  NANDN U128 ( .A(n105), .B(n104), .Z(n111) );
  NAND U129 ( .A(a[6]), .B(b[6]), .Z(n112) );
  AND U130 ( .A(n111), .B(n112), .Z(n107) );
  XOR U131 ( .A(a[7]), .B(b[7]), .Z(n189) );
  ANDN U132 ( .B(n188), .A(n189), .Z(n106) );
  OR U133 ( .A(n107), .B(n106), .Z(n108) );
  AND U134 ( .A(a[7]), .B(b[7]), .Z(n110) );
  ANDN U135 ( .B(n108), .A(n110), .Z(n117) );
  NOR U136 ( .A(n112), .B(n111), .Z(n109) );
  XNOR U137 ( .A(n110), .B(n109), .Z(n115) );
  XOR U138 ( .A(n112), .B(n111), .Z(n113) );
  NAND U139 ( .A(n113), .B(n189), .Z(n114) );
  NAND U140 ( .A(n115), .B(n114), .Z(n194) );
  XNOR U141 ( .A(a[8]), .B(b[8]), .Z(n193) );
  NAND U142 ( .A(n194), .B(n193), .Z(n116) );
  NANDN U143 ( .A(n117), .B(n116), .Z(n123) );
  NAND U144 ( .A(a[8]), .B(b[8]), .Z(n124) );
  AND U145 ( .A(n123), .B(n124), .Z(n119) );
  XOR U146 ( .A(a[9]), .B(b[9]), .Z(n199) );
  ANDN U147 ( .B(n198), .A(n199), .Z(n118) );
  OR U148 ( .A(n119), .B(n118), .Z(n120) );
  AND U149 ( .A(a[9]), .B(b[9]), .Z(n122) );
  ANDN U150 ( .B(n120), .A(n122), .Z(n129) );
  NOR U151 ( .A(n124), .B(n123), .Z(n121) );
  XNOR U152 ( .A(n122), .B(n121), .Z(n127) );
  XOR U153 ( .A(n124), .B(n123), .Z(n125) );
  NAND U154 ( .A(n125), .B(n199), .Z(n126) );
  NAND U155 ( .A(n127), .B(n126), .Z(n204) );
  XNOR U156 ( .A(a[10]), .B(b[10]), .Z(n203) );
  NAND U157 ( .A(n204), .B(n203), .Z(n128) );
  NANDN U158 ( .A(n129), .B(n128), .Z(n135) );
  NAND U159 ( .A(a[10]), .B(b[10]), .Z(n136) );
  AND U160 ( .A(n135), .B(n136), .Z(n131) );
  XOR U161 ( .A(a[11]), .B(b[11]), .Z(n209) );
  ANDN U162 ( .B(n208), .A(n209), .Z(n130) );
  OR U163 ( .A(n131), .B(n130), .Z(n132) );
  AND U164 ( .A(a[11]), .B(b[11]), .Z(n134) );
  ANDN U165 ( .B(n132), .A(n134), .Z(n141) );
  NOR U166 ( .A(n136), .B(n135), .Z(n133) );
  XNOR U167 ( .A(n134), .B(n133), .Z(n139) );
  XOR U168 ( .A(n136), .B(n135), .Z(n137) );
  NAND U169 ( .A(n137), .B(n209), .Z(n138) );
  NAND U170 ( .A(n139), .B(n138), .Z(n214) );
  XNOR U171 ( .A(a[12]), .B(b[12]), .Z(n213) );
  NAND U172 ( .A(n214), .B(n213), .Z(n140) );
  NANDN U173 ( .A(n141), .B(n140), .Z(n146) );
  ANDN U174 ( .B(n145), .A(n146), .Z(n142) );
  XOR U175 ( .A(n147), .B(n142), .Z(n144) );
  XOR U176 ( .A(a[13]), .B(b[13]), .Z(n219) );
  XNOR U177 ( .A(n145), .B(n146), .Z(n218) );
  NAND U178 ( .A(n219), .B(n218), .Z(n143) );
  NAND U179 ( .A(n144), .B(n143), .Z(n224) );
  XNOR U180 ( .A(a[14]), .B(b[14]), .Z(n223) );
  NAND U181 ( .A(a[14]), .B(b[14]), .Z(n149) );
  ANDN U182 ( .B(n148), .A(n149), .Z(n152) );
  XNOR U183 ( .A(n153), .B(n152), .Z(n151) );
  XNOR U184 ( .A(n149), .B(n148), .Z(n228) );
  XOR U185 ( .A(b[15]), .B(a[15]), .Z(n229) );
  NAND U186 ( .A(n228), .B(n229), .Z(n150) );
  NAND U187 ( .A(n151), .B(n150), .Z(N34) );
  AND U188 ( .A(n153), .B(n152), .Z(N35) );
  NAND U190 ( .A(c[0]), .B(rst), .Z(n157) );
  XOR U191 ( .A(n154), .B(carry_on[0]), .Z(n155) );
  NANDN U192 ( .A(rst), .B(n155), .Z(n156) );
  NAND U193 ( .A(n157), .B(n156), .Z(n49) );
  NAND U194 ( .A(c[1]), .B(rst), .Z(n162) );
  XOR U195 ( .A(n159), .B(n158), .Z(n160) );
  NANDN U196 ( .A(rst), .B(n160), .Z(n161) );
  NAND U197 ( .A(n162), .B(n161), .Z(n50) );
  NAND U198 ( .A(c[2]), .B(rst), .Z(n167) );
  XNOR U199 ( .A(n164), .B(n163), .Z(n165) );
  NANDN U200 ( .A(rst), .B(n165), .Z(n166) );
  NAND U201 ( .A(n167), .B(n166), .Z(n51) );
  NAND U202 ( .A(c[3]), .B(rst), .Z(n172) );
  XOR U203 ( .A(n169), .B(n168), .Z(n170) );
  NANDN U204 ( .A(rst), .B(n170), .Z(n171) );
  NAND U205 ( .A(n172), .B(n171), .Z(n52) );
  NAND U206 ( .A(c[4]), .B(rst), .Z(n177) );
  XNOR U207 ( .A(n174), .B(n173), .Z(n175) );
  NANDN U208 ( .A(rst), .B(n175), .Z(n176) );
  NAND U209 ( .A(n177), .B(n176), .Z(n53) );
  NAND U210 ( .A(c[5]), .B(rst), .Z(n182) );
  XOR U211 ( .A(n179), .B(n178), .Z(n180) );
  NANDN U212 ( .A(rst), .B(n180), .Z(n181) );
  NAND U213 ( .A(n182), .B(n181), .Z(n54) );
  NAND U214 ( .A(c[6]), .B(rst), .Z(n187) );
  XNOR U215 ( .A(n184), .B(n183), .Z(n185) );
  NANDN U216 ( .A(rst), .B(n185), .Z(n186) );
  NAND U217 ( .A(n187), .B(n186), .Z(n55) );
  NAND U218 ( .A(c[7]), .B(rst), .Z(n192) );
  XOR U219 ( .A(n189), .B(n188), .Z(n190) );
  NANDN U220 ( .A(rst), .B(n190), .Z(n191) );
  NAND U221 ( .A(n192), .B(n191), .Z(n56) );
  NAND U222 ( .A(c[8]), .B(rst), .Z(n197) );
  XNOR U223 ( .A(n194), .B(n193), .Z(n195) );
  NANDN U224 ( .A(rst), .B(n195), .Z(n196) );
  NAND U225 ( .A(n197), .B(n196), .Z(n57) );
  NAND U226 ( .A(c[9]), .B(rst), .Z(n202) );
  XOR U227 ( .A(n199), .B(n198), .Z(n200) );
  NANDN U228 ( .A(rst), .B(n200), .Z(n201) );
  NAND U229 ( .A(n202), .B(n201), .Z(n58) );
  NAND U230 ( .A(c[10]), .B(rst), .Z(n207) );
  XNOR U231 ( .A(n204), .B(n203), .Z(n205) );
  NANDN U232 ( .A(rst), .B(n205), .Z(n206) );
  NAND U233 ( .A(n207), .B(n206), .Z(n59) );
  NAND U234 ( .A(c[11]), .B(rst), .Z(n212) );
  XOR U235 ( .A(n209), .B(n208), .Z(n210) );
  NANDN U236 ( .A(rst), .B(n210), .Z(n211) );
  NAND U237 ( .A(n212), .B(n211), .Z(n60) );
  NAND U238 ( .A(c[12]), .B(rst), .Z(n217) );
  XNOR U239 ( .A(n214), .B(n213), .Z(n215) );
  NANDN U240 ( .A(rst), .B(n215), .Z(n216) );
  NAND U241 ( .A(n217), .B(n216), .Z(n61) );
  NAND U242 ( .A(c[13]), .B(rst), .Z(n222) );
  XOR U243 ( .A(n219), .B(n218), .Z(n220) );
  NANDN U244 ( .A(rst), .B(n220), .Z(n221) );
  NAND U245 ( .A(n222), .B(n221), .Z(n62) );
  NAND U246 ( .A(c[14]), .B(rst), .Z(n227) );
  XNOR U247 ( .A(n224), .B(n223), .Z(n225) );
  NANDN U248 ( .A(rst), .B(n225), .Z(n226) );
  NAND U249 ( .A(n227), .B(n226), .Z(n63) );
  NAND U250 ( .A(c[15]), .B(rst), .Z(n232) );
  XOR U251 ( .A(n229), .B(n228), .Z(n230) );
  NANDN U252 ( .A(rst), .B(n230), .Z(n231) );
  NAND U253 ( .A(n232), .B(n231), .Z(n64) );
endmodule

