
module hamming_N16000_CC640 ( clk, rst, x, y, o );
  input [24:0] x;
  input [24:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U28 ( .A(n123), .B(n124), .Z(n1) );
  XOR U29 ( .A(n123), .B(n124), .Z(n2) );
  NANDN U30 ( .A(n122), .B(n2), .Z(n3) );
  NAND U31 ( .A(n1), .B(n3), .Z(n134) );
  NAND U32 ( .A(n72), .B(n73), .Z(n4) );
  XOR U33 ( .A(n72), .B(n73), .Z(n5) );
  NANDN U34 ( .A(n71), .B(n5), .Z(n6) );
  NAND U35 ( .A(n4), .B(n6), .Z(n110) );
  NAND U36 ( .A(n98), .B(n96), .Z(n7) );
  XOR U37 ( .A(n98), .B(n96), .Z(n8) );
  NANDN U38 ( .A(n97), .B(n8), .Z(n9) );
  NAND U39 ( .A(n7), .B(n9), .Z(n104) );
  NAND U40 ( .A(n133), .B(n134), .Z(n10) );
  XOR U41 ( .A(n133), .B(n134), .Z(n11) );
  NAND U42 ( .A(n11), .B(n132), .Z(n12) );
  NAND U43 ( .A(n10), .B(n12), .Z(n154) );
  NANDN U44 ( .A(n82), .B(n83), .Z(n13) );
  NANDN U45 ( .A(n81), .B(n80), .Z(n14) );
  AND U46 ( .A(n13), .B(n14), .Z(n117) );
  NAND U47 ( .A(n100), .B(n101), .Z(n15) );
  XOR U48 ( .A(n100), .B(n101), .Z(n16) );
  NANDN U49 ( .A(n99), .B(n16), .Z(n17) );
  NAND U50 ( .A(n15), .B(n17), .Z(n127) );
  NAND U51 ( .A(n150), .B(n152), .Z(n18) );
  XOR U52 ( .A(n150), .B(n152), .Z(n19) );
  NAND U53 ( .A(n19), .B(n151), .Z(n20) );
  NAND U54 ( .A(n18), .B(n20), .Z(n160) );
  NAND U55 ( .A(n120), .B(n121), .Z(n21) );
  XOR U56 ( .A(n120), .B(n121), .Z(n22) );
  NANDN U57 ( .A(n119), .B(n22), .Z(n23) );
  NAND U58 ( .A(n21), .B(n23), .Z(n132) );
  NAND U59 ( .A(n117), .B(n115), .Z(n24) );
  XOR U60 ( .A(n117), .B(n115), .Z(n25) );
  NANDN U61 ( .A(n116), .B(n25), .Z(n26) );
  NAND U62 ( .A(n24), .B(n26), .Z(n137) );
  NAND U63 ( .A(n128), .B(n129), .Z(n27) );
  XOR U64 ( .A(n128), .B(n129), .Z(n28) );
  NANDN U65 ( .A(n127), .B(n28), .Z(n29) );
  NAND U66 ( .A(n27), .B(n29), .Z(n144) );
  NAND U67 ( .A(n160), .B(n159), .Z(n30) );
  XOR U68 ( .A(n160), .B(n159), .Z(n31) );
  NANDN U69 ( .A(oglobal[4]), .B(n31), .Z(n32) );
  NAND U70 ( .A(n30), .B(n32), .Z(n161) );
  NANDN U71 ( .A(n168), .B(oglobal[12]), .Z(n33) );
  XNOR U72 ( .A(oglobal[13]), .B(n33), .Z(o[13]) );
  XOR U73 ( .A(x[17]), .B(y[17]), .Z(n80) );
  XNOR U74 ( .A(x[13]), .B(y[13]), .Z(n81) );
  XNOR U75 ( .A(n80), .B(n81), .Z(n83) );
  XOR U76 ( .A(x[21]), .B(y[21]), .Z(n38) );
  XOR U77 ( .A(x[23]), .B(y[23]), .Z(n37) );
  XNOR U78 ( .A(n38), .B(n37), .Z(n82) );
  XNOR U79 ( .A(n83), .B(n82), .Z(n73) );
  XOR U80 ( .A(x[15]), .B(y[15]), .Z(n85) );
  XNOR U81 ( .A(x[19]), .B(y[19]), .Z(n84) );
  XOR U82 ( .A(oglobal[0]), .B(n84), .Z(n86) );
  XNOR U83 ( .A(n85), .B(n86), .Z(n72) );
  XOR U84 ( .A(x[7]), .B(y[7]), .Z(n76) );
  XOR U85 ( .A(x[11]), .B(y[11]), .Z(n74) );
  XNOR U86 ( .A(x[9]), .B(y[9]), .Z(n75) );
  XOR U87 ( .A(n74), .B(n75), .Z(n77) );
  XOR U88 ( .A(n76), .B(n77), .Z(n71) );
  XOR U89 ( .A(n72), .B(n71), .Z(n34) );
  XNOR U90 ( .A(n73), .B(n34), .Z(n101) );
  XOR U91 ( .A(x[4]), .B(y[4]), .Z(n66) );
  XOR U92 ( .A(x[2]), .B(y[2]), .Z(n64) );
  XNOR U93 ( .A(x[0]), .B(y[0]), .Z(n65) );
  XOR U94 ( .A(n64), .B(n65), .Z(n67) );
  XOR U95 ( .A(n66), .B(n67), .Z(n97) );
  XOR U96 ( .A(x[1]), .B(y[1]), .Z(n60) );
  XOR U97 ( .A(x[5]), .B(y[5]), .Z(n58) );
  XNOR U98 ( .A(x[3]), .B(y[3]), .Z(n59) );
  XOR U99 ( .A(n58), .B(n59), .Z(n61) );
  XNOR U100 ( .A(n60), .B(n61), .Z(n98) );
  XOR U101 ( .A(x[20]), .B(y[20]), .Z(n41) );
  XOR U102 ( .A(x[24]), .B(y[24]), .Z(n39) );
  XNOR U103 ( .A(x[18]), .B(y[18]), .Z(n40) );
  XOR U104 ( .A(n39), .B(n40), .Z(n42) );
  XNOR U105 ( .A(n41), .B(n42), .Z(n96) );
  XNOR U106 ( .A(n98), .B(n96), .Z(n35) );
  XOR U107 ( .A(n97), .B(n35), .Z(n100) );
  XOR U108 ( .A(x[10]), .B(y[10]), .Z(n54) );
  XOR U109 ( .A(x[8]), .B(y[8]), .Z(n52) );
  XNOR U110 ( .A(x[6]), .B(y[6]), .Z(n53) );
  XOR U111 ( .A(n52), .B(n53), .Z(n55) );
  XNOR U112 ( .A(n54), .B(n55), .Z(n92) );
  XOR U113 ( .A(x[22]), .B(y[22]), .Z(n90) );
  XOR U114 ( .A(x[16]), .B(y[16]), .Z(n47) );
  XOR U115 ( .A(x[14]), .B(y[14]), .Z(n45) );
  XNOR U116 ( .A(x[12]), .B(y[12]), .Z(n46) );
  XOR U117 ( .A(n45), .B(n46), .Z(n48) );
  XOR U118 ( .A(n47), .B(n48), .Z(n91) );
  XOR U119 ( .A(n90), .B(n91), .Z(n93) );
  XOR U120 ( .A(n92), .B(n93), .Z(n99) );
  XOR U121 ( .A(n100), .B(n99), .Z(n36) );
  XNOR U122 ( .A(n101), .B(n36), .Z(o[0]) );
  AND U123 ( .A(n38), .B(n37), .Z(n125) );
  XOR U124 ( .A(n125), .B(oglobal[1]), .Z(n120) );
  NANDN U125 ( .A(n40), .B(n39), .Z(n44) );
  NANDN U126 ( .A(n42), .B(n41), .Z(n43) );
  NAND U127 ( .A(n44), .B(n43), .Z(n121) );
  NANDN U128 ( .A(n46), .B(n45), .Z(n50) );
  NANDN U129 ( .A(n48), .B(n47), .Z(n49) );
  AND U130 ( .A(n50), .B(n49), .Z(n119) );
  XOR U131 ( .A(n121), .B(n119), .Z(n51) );
  XOR U132 ( .A(n120), .B(n51), .Z(n111) );
  NANDN U133 ( .A(n53), .B(n52), .Z(n57) );
  NANDN U134 ( .A(n55), .B(n54), .Z(n56) );
  NAND U135 ( .A(n57), .B(n56), .Z(n123) );
  NANDN U136 ( .A(n59), .B(n58), .Z(n63) );
  NANDN U137 ( .A(n61), .B(n60), .Z(n62) );
  NAND U138 ( .A(n63), .B(n62), .Z(n124) );
  NANDN U139 ( .A(n65), .B(n64), .Z(n69) );
  NANDN U140 ( .A(n67), .B(n66), .Z(n68) );
  AND U141 ( .A(n69), .B(n68), .Z(n122) );
  XOR U142 ( .A(n124), .B(n122), .Z(n70) );
  XOR U143 ( .A(n123), .B(n70), .Z(n109) );
  XOR U144 ( .A(n109), .B(n110), .Z(n112) );
  XNOR U145 ( .A(n111), .B(n112), .Z(n128) );
  NANDN U146 ( .A(n75), .B(n74), .Z(n79) );
  NANDN U147 ( .A(n77), .B(n76), .Z(n78) );
  NAND U148 ( .A(n79), .B(n78), .Z(n116) );
  NANDN U149 ( .A(n84), .B(oglobal[0]), .Z(n88) );
  NANDN U150 ( .A(n86), .B(n85), .Z(n87) );
  AND U151 ( .A(n88), .B(n87), .Z(n115) );
  XNOR U152 ( .A(n117), .B(n115), .Z(n89) );
  XOR U153 ( .A(n116), .B(n89), .Z(n105) );
  NANDN U154 ( .A(n91), .B(n90), .Z(n95) );
  NANDN U155 ( .A(n93), .B(n92), .Z(n94) );
  AND U156 ( .A(n95), .B(n94), .Z(n103) );
  XOR U157 ( .A(n103), .B(n104), .Z(n106) );
  XNOR U158 ( .A(n105), .B(n106), .Z(n129) );
  XNOR U159 ( .A(n129), .B(n127), .Z(n102) );
  XNOR U160 ( .A(n128), .B(n102), .Z(o[1]) );
  NANDN U161 ( .A(n104), .B(n103), .Z(n108) );
  NANDN U162 ( .A(n106), .B(n105), .Z(n107) );
  AND U163 ( .A(n108), .B(n107), .Z(n138) );
  NANDN U164 ( .A(n110), .B(n109), .Z(n114) );
  NANDN U165 ( .A(n112), .B(n111), .Z(n113) );
  NAND U166 ( .A(n114), .B(n113), .Z(n136) );
  IV U167 ( .A(n136), .Z(n135) );
  XNOR U168 ( .A(n135), .B(n137), .Z(n118) );
  XNOR U169 ( .A(n138), .B(n118), .Z(n145) );
  AND U170 ( .A(n125), .B(oglobal[1]), .Z(n131) );
  XOR U171 ( .A(n131), .B(oglobal[2]), .Z(n133) );
  XOR U172 ( .A(n134), .B(n133), .Z(n126) );
  XNOR U173 ( .A(n132), .B(n126), .Z(n143) );
  IV U174 ( .A(n143), .Z(n142) );
  XNOR U175 ( .A(n142), .B(n144), .Z(n130) );
  XNOR U176 ( .A(n145), .B(n130), .Z(o[2]) );
  AND U177 ( .A(n131), .B(oglobal[2]), .Z(n153) );
  XOR U178 ( .A(oglobal[3]), .B(n153), .Z(n155) );
  XNOR U179 ( .A(n155), .B(n154), .Z(n152) );
  NANDN U180 ( .A(n137), .B(n135), .Z(n141) );
  AND U181 ( .A(n137), .B(n136), .Z(n139) );
  NANDN U182 ( .A(n139), .B(n138), .Z(n140) );
  AND U183 ( .A(n141), .B(n140), .Z(n151) );
  NANDN U184 ( .A(n144), .B(n142), .Z(n148) );
  AND U185 ( .A(n144), .B(n143), .Z(n146) );
  OR U186 ( .A(n146), .B(n145), .Z(n147) );
  AND U187 ( .A(n148), .B(n147), .Z(n150) );
  XOR U188 ( .A(n151), .B(n150), .Z(n149) );
  XNOR U189 ( .A(n152), .B(n149), .Z(o[3]) );
  NAND U190 ( .A(n153), .B(oglobal[3]), .Z(n157) );
  NAND U191 ( .A(n155), .B(n154), .Z(n156) );
  AND U192 ( .A(n157), .B(n156), .Z(n159) );
  XNOR U193 ( .A(n160), .B(n159), .Z(n158) );
  XNOR U194 ( .A(oglobal[4]), .B(n158), .Z(o[4]) );
  XNOR U195 ( .A(n161), .B(oglobal[5]), .Z(o[5]) );
  ANDN U196 ( .B(oglobal[5]), .A(n161), .Z(n162) );
  XOR U197 ( .A(n162), .B(oglobal[6]), .Z(o[6]) );
  AND U198 ( .A(n162), .B(oglobal[6]), .Z(n163) );
  XOR U199 ( .A(n163), .B(oglobal[7]), .Z(o[7]) );
  AND U200 ( .A(n163), .B(oglobal[7]), .Z(n164) );
  XOR U201 ( .A(n164), .B(oglobal[8]), .Z(o[8]) );
  AND U202 ( .A(n164), .B(oglobal[8]), .Z(n165) );
  XOR U203 ( .A(n165), .B(oglobal[9]), .Z(o[9]) );
  AND U204 ( .A(n165), .B(oglobal[9]), .Z(n166) );
  XOR U205 ( .A(n166), .B(oglobal[10]), .Z(o[10]) );
  AND U206 ( .A(n166), .B(oglobal[10]), .Z(n167) );
  XOR U207 ( .A(n167), .B(oglobal[11]), .Z(o[11]) );
  NAND U208 ( .A(n167), .B(oglobal[11]), .Z(n168) );
  XNOR U209 ( .A(oglobal[12]), .B(n168), .Z(o[12]) );
endmodule

