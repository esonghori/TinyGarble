
module sum_N1024_CC8 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[0]), .B(b[0]), .Z(n1) );
  XOR U4 ( .A(n1), .B(carry_on), .Z(c[0]) );
  XOR U5 ( .A(a[1]), .B(b[1]), .Z(n4) );
  NAND U6 ( .A(b[0]), .B(a[0]), .Z(n3) );
  NAND U7 ( .A(carry_on), .B(n1), .Z(n2) );
  AND U8 ( .A(n3), .B(n2), .Z(n5) );
  XNOR U9 ( .A(n4), .B(n5), .Z(c[1]) );
  XOR U10 ( .A(a[2]), .B(b[2]), .Z(n8) );
  NAND U11 ( .A(b[1]), .B(a[1]), .Z(n7) );
  NANDN U12 ( .A(n5), .B(n4), .Z(n6) );
  AND U13 ( .A(n7), .B(n6), .Z(n9) );
  XNOR U14 ( .A(n8), .B(n9), .Z(c[2]) );
  XOR U15 ( .A(a[3]), .B(b[3]), .Z(n12) );
  NAND U16 ( .A(b[2]), .B(a[2]), .Z(n11) );
  NANDN U17 ( .A(n9), .B(n8), .Z(n10) );
  AND U18 ( .A(n11), .B(n10), .Z(n13) );
  XNOR U19 ( .A(n12), .B(n13), .Z(c[3]) );
  XOR U20 ( .A(a[4]), .B(b[4]), .Z(n16) );
  NAND U21 ( .A(b[3]), .B(a[3]), .Z(n15) );
  NANDN U22 ( .A(n13), .B(n12), .Z(n14) );
  AND U23 ( .A(n15), .B(n14), .Z(n17) );
  XNOR U24 ( .A(n16), .B(n17), .Z(c[4]) );
  XOR U25 ( .A(a[5]), .B(b[5]), .Z(n20) );
  NAND U26 ( .A(b[4]), .B(a[4]), .Z(n19) );
  NANDN U27 ( .A(n17), .B(n16), .Z(n18) );
  AND U28 ( .A(n19), .B(n18), .Z(n21) );
  XNOR U29 ( .A(n20), .B(n21), .Z(c[5]) );
  XOR U30 ( .A(a[6]), .B(b[6]), .Z(n24) );
  NAND U31 ( .A(b[5]), .B(a[5]), .Z(n23) );
  NANDN U32 ( .A(n21), .B(n20), .Z(n22) );
  AND U33 ( .A(n23), .B(n22), .Z(n25) );
  XNOR U34 ( .A(n24), .B(n25), .Z(c[6]) );
  XOR U35 ( .A(a[7]), .B(b[7]), .Z(n28) );
  NAND U36 ( .A(b[6]), .B(a[6]), .Z(n27) );
  NANDN U37 ( .A(n25), .B(n24), .Z(n26) );
  AND U38 ( .A(n27), .B(n26), .Z(n29) );
  XNOR U39 ( .A(n28), .B(n29), .Z(c[7]) );
  XOR U40 ( .A(a[8]), .B(b[8]), .Z(n32) );
  NAND U41 ( .A(b[7]), .B(a[7]), .Z(n31) );
  NANDN U42 ( .A(n29), .B(n28), .Z(n30) );
  AND U43 ( .A(n31), .B(n30), .Z(n33) );
  XNOR U44 ( .A(n32), .B(n33), .Z(c[8]) );
  XOR U45 ( .A(a[9]), .B(b[9]), .Z(n36) );
  NAND U46 ( .A(b[8]), .B(a[8]), .Z(n35) );
  NANDN U47 ( .A(n33), .B(n32), .Z(n34) );
  AND U48 ( .A(n35), .B(n34), .Z(n37) );
  XNOR U49 ( .A(n36), .B(n37), .Z(c[9]) );
  XOR U50 ( .A(a[10]), .B(b[10]), .Z(n40) );
  NAND U51 ( .A(b[9]), .B(a[9]), .Z(n39) );
  NANDN U52 ( .A(n37), .B(n36), .Z(n38) );
  AND U53 ( .A(n39), .B(n38), .Z(n41) );
  XNOR U54 ( .A(n40), .B(n41), .Z(c[10]) );
  XOR U55 ( .A(a[11]), .B(b[11]), .Z(n44) );
  NAND U56 ( .A(b[10]), .B(a[10]), .Z(n43) );
  NANDN U57 ( .A(n41), .B(n40), .Z(n42) );
  AND U58 ( .A(n43), .B(n42), .Z(n45) );
  XNOR U59 ( .A(n44), .B(n45), .Z(c[11]) );
  XOR U60 ( .A(a[12]), .B(b[12]), .Z(n48) );
  NAND U61 ( .A(b[11]), .B(a[11]), .Z(n47) );
  NANDN U62 ( .A(n45), .B(n44), .Z(n46) );
  AND U63 ( .A(n47), .B(n46), .Z(n49) );
  XNOR U64 ( .A(n48), .B(n49), .Z(c[12]) );
  XOR U65 ( .A(a[13]), .B(b[13]), .Z(n52) );
  NAND U66 ( .A(b[12]), .B(a[12]), .Z(n51) );
  NANDN U67 ( .A(n49), .B(n48), .Z(n50) );
  AND U68 ( .A(n51), .B(n50), .Z(n53) );
  XNOR U69 ( .A(n52), .B(n53), .Z(c[13]) );
  XOR U70 ( .A(a[14]), .B(b[14]), .Z(n56) );
  NAND U71 ( .A(b[13]), .B(a[13]), .Z(n55) );
  NANDN U72 ( .A(n53), .B(n52), .Z(n54) );
  AND U73 ( .A(n55), .B(n54), .Z(n57) );
  XNOR U74 ( .A(n56), .B(n57), .Z(c[14]) );
  XOR U75 ( .A(a[15]), .B(b[15]), .Z(n60) );
  NAND U76 ( .A(b[14]), .B(a[14]), .Z(n59) );
  NANDN U77 ( .A(n57), .B(n56), .Z(n58) );
  AND U78 ( .A(n59), .B(n58), .Z(n61) );
  XNOR U79 ( .A(n60), .B(n61), .Z(c[15]) );
  XOR U80 ( .A(a[16]), .B(b[16]), .Z(n64) );
  NAND U81 ( .A(b[15]), .B(a[15]), .Z(n63) );
  NANDN U82 ( .A(n61), .B(n60), .Z(n62) );
  AND U83 ( .A(n63), .B(n62), .Z(n65) );
  XNOR U84 ( .A(n64), .B(n65), .Z(c[16]) );
  XOR U85 ( .A(a[17]), .B(b[17]), .Z(n68) );
  NAND U86 ( .A(b[16]), .B(a[16]), .Z(n67) );
  NANDN U87 ( .A(n65), .B(n64), .Z(n66) );
  AND U88 ( .A(n67), .B(n66), .Z(n69) );
  XNOR U89 ( .A(n68), .B(n69), .Z(c[17]) );
  XOR U90 ( .A(a[18]), .B(b[18]), .Z(n72) );
  NAND U91 ( .A(b[17]), .B(a[17]), .Z(n71) );
  NANDN U92 ( .A(n69), .B(n68), .Z(n70) );
  AND U93 ( .A(n71), .B(n70), .Z(n73) );
  XNOR U94 ( .A(n72), .B(n73), .Z(c[18]) );
  XOR U95 ( .A(a[19]), .B(b[19]), .Z(n76) );
  NAND U96 ( .A(b[18]), .B(a[18]), .Z(n75) );
  NANDN U97 ( .A(n73), .B(n72), .Z(n74) );
  AND U98 ( .A(n75), .B(n74), .Z(n77) );
  XNOR U99 ( .A(n76), .B(n77), .Z(c[19]) );
  XOR U100 ( .A(a[20]), .B(b[20]), .Z(n80) );
  NAND U101 ( .A(b[19]), .B(a[19]), .Z(n79) );
  NANDN U102 ( .A(n77), .B(n76), .Z(n78) );
  AND U103 ( .A(n79), .B(n78), .Z(n81) );
  XNOR U104 ( .A(n80), .B(n81), .Z(c[20]) );
  XOR U105 ( .A(a[21]), .B(b[21]), .Z(n84) );
  NAND U106 ( .A(b[20]), .B(a[20]), .Z(n83) );
  NANDN U107 ( .A(n81), .B(n80), .Z(n82) );
  AND U108 ( .A(n83), .B(n82), .Z(n85) );
  XNOR U109 ( .A(n84), .B(n85), .Z(c[21]) );
  XOR U110 ( .A(a[22]), .B(b[22]), .Z(n88) );
  NAND U111 ( .A(b[21]), .B(a[21]), .Z(n87) );
  NANDN U112 ( .A(n85), .B(n84), .Z(n86) );
  AND U113 ( .A(n87), .B(n86), .Z(n89) );
  XNOR U114 ( .A(n88), .B(n89), .Z(c[22]) );
  XOR U115 ( .A(a[23]), .B(b[23]), .Z(n92) );
  NAND U116 ( .A(b[22]), .B(a[22]), .Z(n91) );
  NANDN U117 ( .A(n89), .B(n88), .Z(n90) );
  AND U118 ( .A(n91), .B(n90), .Z(n93) );
  XNOR U119 ( .A(n92), .B(n93), .Z(c[23]) );
  XOR U120 ( .A(a[24]), .B(b[24]), .Z(n96) );
  NAND U121 ( .A(b[23]), .B(a[23]), .Z(n95) );
  NANDN U122 ( .A(n93), .B(n92), .Z(n94) );
  AND U123 ( .A(n95), .B(n94), .Z(n97) );
  XNOR U124 ( .A(n96), .B(n97), .Z(c[24]) );
  XOR U125 ( .A(a[25]), .B(b[25]), .Z(n100) );
  NAND U126 ( .A(b[24]), .B(a[24]), .Z(n99) );
  NANDN U127 ( .A(n97), .B(n96), .Z(n98) );
  AND U128 ( .A(n99), .B(n98), .Z(n101) );
  XNOR U129 ( .A(n100), .B(n101), .Z(c[25]) );
  XOR U130 ( .A(a[26]), .B(b[26]), .Z(n104) );
  NAND U131 ( .A(b[25]), .B(a[25]), .Z(n103) );
  NANDN U132 ( .A(n101), .B(n100), .Z(n102) );
  AND U133 ( .A(n103), .B(n102), .Z(n105) );
  XNOR U134 ( .A(n104), .B(n105), .Z(c[26]) );
  XOR U135 ( .A(a[27]), .B(b[27]), .Z(n108) );
  NAND U136 ( .A(b[26]), .B(a[26]), .Z(n107) );
  NANDN U137 ( .A(n105), .B(n104), .Z(n106) );
  AND U138 ( .A(n107), .B(n106), .Z(n109) );
  XNOR U139 ( .A(n108), .B(n109), .Z(c[27]) );
  XOR U140 ( .A(a[28]), .B(b[28]), .Z(n112) );
  NAND U141 ( .A(b[27]), .B(a[27]), .Z(n111) );
  NANDN U142 ( .A(n109), .B(n108), .Z(n110) );
  AND U143 ( .A(n111), .B(n110), .Z(n113) );
  XNOR U144 ( .A(n112), .B(n113), .Z(c[28]) );
  XOR U145 ( .A(a[29]), .B(b[29]), .Z(n116) );
  NAND U146 ( .A(b[28]), .B(a[28]), .Z(n115) );
  NANDN U147 ( .A(n113), .B(n112), .Z(n114) );
  AND U148 ( .A(n115), .B(n114), .Z(n117) );
  XNOR U149 ( .A(n116), .B(n117), .Z(c[29]) );
  XOR U150 ( .A(a[30]), .B(b[30]), .Z(n120) );
  NAND U151 ( .A(b[29]), .B(a[29]), .Z(n119) );
  NANDN U152 ( .A(n117), .B(n116), .Z(n118) );
  AND U153 ( .A(n119), .B(n118), .Z(n121) );
  XNOR U154 ( .A(n120), .B(n121), .Z(c[30]) );
  XOR U155 ( .A(a[31]), .B(b[31]), .Z(n124) );
  NAND U156 ( .A(b[30]), .B(a[30]), .Z(n123) );
  NANDN U157 ( .A(n121), .B(n120), .Z(n122) );
  AND U158 ( .A(n123), .B(n122), .Z(n125) );
  XNOR U159 ( .A(n124), .B(n125), .Z(c[31]) );
  XOR U160 ( .A(a[32]), .B(b[32]), .Z(n128) );
  NAND U161 ( .A(b[31]), .B(a[31]), .Z(n127) );
  NANDN U162 ( .A(n125), .B(n124), .Z(n126) );
  AND U163 ( .A(n127), .B(n126), .Z(n129) );
  XNOR U164 ( .A(n128), .B(n129), .Z(c[32]) );
  XOR U165 ( .A(a[33]), .B(b[33]), .Z(n132) );
  NAND U166 ( .A(b[32]), .B(a[32]), .Z(n131) );
  NANDN U167 ( .A(n129), .B(n128), .Z(n130) );
  AND U168 ( .A(n131), .B(n130), .Z(n133) );
  XNOR U169 ( .A(n132), .B(n133), .Z(c[33]) );
  XOR U170 ( .A(a[34]), .B(b[34]), .Z(n136) );
  NAND U171 ( .A(b[33]), .B(a[33]), .Z(n135) );
  NANDN U172 ( .A(n133), .B(n132), .Z(n134) );
  AND U173 ( .A(n135), .B(n134), .Z(n137) );
  XNOR U174 ( .A(n136), .B(n137), .Z(c[34]) );
  XOR U175 ( .A(a[35]), .B(b[35]), .Z(n140) );
  NAND U176 ( .A(b[34]), .B(a[34]), .Z(n139) );
  NANDN U177 ( .A(n137), .B(n136), .Z(n138) );
  AND U178 ( .A(n139), .B(n138), .Z(n141) );
  XNOR U179 ( .A(n140), .B(n141), .Z(c[35]) );
  XOR U180 ( .A(a[36]), .B(b[36]), .Z(n144) );
  NAND U181 ( .A(b[35]), .B(a[35]), .Z(n143) );
  NANDN U182 ( .A(n141), .B(n140), .Z(n142) );
  AND U183 ( .A(n143), .B(n142), .Z(n145) );
  XNOR U184 ( .A(n144), .B(n145), .Z(c[36]) );
  XOR U185 ( .A(a[37]), .B(b[37]), .Z(n148) );
  NAND U186 ( .A(b[36]), .B(a[36]), .Z(n147) );
  NANDN U187 ( .A(n145), .B(n144), .Z(n146) );
  AND U188 ( .A(n147), .B(n146), .Z(n149) );
  XNOR U189 ( .A(n148), .B(n149), .Z(c[37]) );
  XOR U190 ( .A(a[38]), .B(b[38]), .Z(n152) );
  NAND U191 ( .A(b[37]), .B(a[37]), .Z(n151) );
  NANDN U192 ( .A(n149), .B(n148), .Z(n150) );
  AND U193 ( .A(n151), .B(n150), .Z(n153) );
  XNOR U194 ( .A(n152), .B(n153), .Z(c[38]) );
  XOR U195 ( .A(a[39]), .B(b[39]), .Z(n156) );
  NAND U196 ( .A(b[38]), .B(a[38]), .Z(n155) );
  NANDN U197 ( .A(n153), .B(n152), .Z(n154) );
  AND U198 ( .A(n155), .B(n154), .Z(n157) );
  XNOR U199 ( .A(n156), .B(n157), .Z(c[39]) );
  XOR U200 ( .A(a[40]), .B(b[40]), .Z(n160) );
  NAND U201 ( .A(b[39]), .B(a[39]), .Z(n159) );
  NANDN U202 ( .A(n157), .B(n156), .Z(n158) );
  AND U203 ( .A(n159), .B(n158), .Z(n161) );
  XNOR U204 ( .A(n160), .B(n161), .Z(c[40]) );
  XOR U205 ( .A(a[41]), .B(b[41]), .Z(n164) );
  NAND U206 ( .A(b[40]), .B(a[40]), .Z(n163) );
  NANDN U207 ( .A(n161), .B(n160), .Z(n162) );
  AND U208 ( .A(n163), .B(n162), .Z(n165) );
  XNOR U209 ( .A(n164), .B(n165), .Z(c[41]) );
  XOR U210 ( .A(a[42]), .B(b[42]), .Z(n168) );
  NAND U211 ( .A(b[41]), .B(a[41]), .Z(n167) );
  NANDN U212 ( .A(n165), .B(n164), .Z(n166) );
  AND U213 ( .A(n167), .B(n166), .Z(n169) );
  XNOR U214 ( .A(n168), .B(n169), .Z(c[42]) );
  XOR U215 ( .A(a[43]), .B(b[43]), .Z(n172) );
  NAND U216 ( .A(b[42]), .B(a[42]), .Z(n171) );
  NANDN U217 ( .A(n169), .B(n168), .Z(n170) );
  AND U218 ( .A(n171), .B(n170), .Z(n173) );
  XNOR U219 ( .A(n172), .B(n173), .Z(c[43]) );
  XOR U220 ( .A(a[44]), .B(b[44]), .Z(n176) );
  NAND U221 ( .A(b[43]), .B(a[43]), .Z(n175) );
  NANDN U222 ( .A(n173), .B(n172), .Z(n174) );
  AND U223 ( .A(n175), .B(n174), .Z(n177) );
  XNOR U224 ( .A(n176), .B(n177), .Z(c[44]) );
  XOR U225 ( .A(a[45]), .B(b[45]), .Z(n180) );
  NAND U226 ( .A(b[44]), .B(a[44]), .Z(n179) );
  NANDN U227 ( .A(n177), .B(n176), .Z(n178) );
  AND U228 ( .A(n179), .B(n178), .Z(n181) );
  XNOR U229 ( .A(n180), .B(n181), .Z(c[45]) );
  XOR U230 ( .A(a[46]), .B(b[46]), .Z(n184) );
  NAND U231 ( .A(b[45]), .B(a[45]), .Z(n183) );
  NANDN U232 ( .A(n181), .B(n180), .Z(n182) );
  AND U233 ( .A(n183), .B(n182), .Z(n185) );
  XNOR U234 ( .A(n184), .B(n185), .Z(c[46]) );
  XOR U235 ( .A(a[47]), .B(b[47]), .Z(n188) );
  NAND U236 ( .A(b[46]), .B(a[46]), .Z(n187) );
  NANDN U237 ( .A(n185), .B(n184), .Z(n186) );
  AND U238 ( .A(n187), .B(n186), .Z(n189) );
  XNOR U239 ( .A(n188), .B(n189), .Z(c[47]) );
  XOR U240 ( .A(a[48]), .B(b[48]), .Z(n192) );
  NAND U241 ( .A(b[47]), .B(a[47]), .Z(n191) );
  NANDN U242 ( .A(n189), .B(n188), .Z(n190) );
  AND U243 ( .A(n191), .B(n190), .Z(n193) );
  XNOR U244 ( .A(n192), .B(n193), .Z(c[48]) );
  XOR U245 ( .A(a[49]), .B(b[49]), .Z(n196) );
  NAND U246 ( .A(b[48]), .B(a[48]), .Z(n195) );
  NANDN U247 ( .A(n193), .B(n192), .Z(n194) );
  AND U248 ( .A(n195), .B(n194), .Z(n197) );
  XNOR U249 ( .A(n196), .B(n197), .Z(c[49]) );
  XOR U250 ( .A(a[50]), .B(b[50]), .Z(n200) );
  NAND U251 ( .A(b[49]), .B(a[49]), .Z(n199) );
  NANDN U252 ( .A(n197), .B(n196), .Z(n198) );
  AND U253 ( .A(n199), .B(n198), .Z(n201) );
  XNOR U254 ( .A(n200), .B(n201), .Z(c[50]) );
  XOR U255 ( .A(a[51]), .B(b[51]), .Z(n204) );
  NAND U256 ( .A(b[50]), .B(a[50]), .Z(n203) );
  NANDN U257 ( .A(n201), .B(n200), .Z(n202) );
  AND U258 ( .A(n203), .B(n202), .Z(n205) );
  XNOR U259 ( .A(n204), .B(n205), .Z(c[51]) );
  XOR U260 ( .A(a[52]), .B(b[52]), .Z(n208) );
  NAND U261 ( .A(b[51]), .B(a[51]), .Z(n207) );
  NANDN U262 ( .A(n205), .B(n204), .Z(n206) );
  AND U263 ( .A(n207), .B(n206), .Z(n209) );
  XNOR U264 ( .A(n208), .B(n209), .Z(c[52]) );
  XOR U265 ( .A(a[53]), .B(b[53]), .Z(n212) );
  NAND U266 ( .A(b[52]), .B(a[52]), .Z(n211) );
  NANDN U267 ( .A(n209), .B(n208), .Z(n210) );
  AND U268 ( .A(n211), .B(n210), .Z(n213) );
  XNOR U269 ( .A(n212), .B(n213), .Z(c[53]) );
  XOR U270 ( .A(a[54]), .B(b[54]), .Z(n216) );
  NAND U271 ( .A(b[53]), .B(a[53]), .Z(n215) );
  NANDN U272 ( .A(n213), .B(n212), .Z(n214) );
  AND U273 ( .A(n215), .B(n214), .Z(n217) );
  XNOR U274 ( .A(n216), .B(n217), .Z(c[54]) );
  XOR U275 ( .A(a[55]), .B(b[55]), .Z(n220) );
  NAND U276 ( .A(b[54]), .B(a[54]), .Z(n219) );
  NANDN U277 ( .A(n217), .B(n216), .Z(n218) );
  AND U278 ( .A(n219), .B(n218), .Z(n221) );
  XNOR U279 ( .A(n220), .B(n221), .Z(c[55]) );
  XOR U280 ( .A(a[56]), .B(b[56]), .Z(n224) );
  NAND U281 ( .A(b[55]), .B(a[55]), .Z(n223) );
  NANDN U282 ( .A(n221), .B(n220), .Z(n222) );
  AND U283 ( .A(n223), .B(n222), .Z(n225) );
  XNOR U284 ( .A(n224), .B(n225), .Z(c[56]) );
  XOR U285 ( .A(a[57]), .B(b[57]), .Z(n228) );
  NAND U286 ( .A(b[56]), .B(a[56]), .Z(n227) );
  NANDN U287 ( .A(n225), .B(n224), .Z(n226) );
  AND U288 ( .A(n227), .B(n226), .Z(n229) );
  XNOR U289 ( .A(n228), .B(n229), .Z(c[57]) );
  XOR U290 ( .A(a[58]), .B(b[58]), .Z(n232) );
  NAND U291 ( .A(b[57]), .B(a[57]), .Z(n231) );
  NANDN U292 ( .A(n229), .B(n228), .Z(n230) );
  AND U293 ( .A(n231), .B(n230), .Z(n233) );
  XNOR U294 ( .A(n232), .B(n233), .Z(c[58]) );
  XOR U295 ( .A(a[59]), .B(b[59]), .Z(n236) );
  NAND U296 ( .A(b[58]), .B(a[58]), .Z(n235) );
  NANDN U297 ( .A(n233), .B(n232), .Z(n234) );
  AND U298 ( .A(n235), .B(n234), .Z(n237) );
  XNOR U299 ( .A(n236), .B(n237), .Z(c[59]) );
  XOR U300 ( .A(a[60]), .B(b[60]), .Z(n240) );
  NAND U301 ( .A(b[59]), .B(a[59]), .Z(n239) );
  NANDN U302 ( .A(n237), .B(n236), .Z(n238) );
  AND U303 ( .A(n239), .B(n238), .Z(n241) );
  XNOR U304 ( .A(n240), .B(n241), .Z(c[60]) );
  XOR U305 ( .A(a[61]), .B(b[61]), .Z(n244) );
  NAND U306 ( .A(b[60]), .B(a[60]), .Z(n243) );
  NANDN U307 ( .A(n241), .B(n240), .Z(n242) );
  AND U308 ( .A(n243), .B(n242), .Z(n245) );
  XNOR U309 ( .A(n244), .B(n245), .Z(c[61]) );
  XOR U310 ( .A(a[62]), .B(b[62]), .Z(n248) );
  NAND U311 ( .A(b[61]), .B(a[61]), .Z(n247) );
  NANDN U312 ( .A(n245), .B(n244), .Z(n246) );
  AND U313 ( .A(n247), .B(n246), .Z(n249) );
  XNOR U314 ( .A(n248), .B(n249), .Z(c[62]) );
  XOR U315 ( .A(a[63]), .B(b[63]), .Z(n252) );
  NAND U316 ( .A(b[62]), .B(a[62]), .Z(n251) );
  NANDN U317 ( .A(n249), .B(n248), .Z(n250) );
  AND U318 ( .A(n251), .B(n250), .Z(n253) );
  XNOR U319 ( .A(n252), .B(n253), .Z(c[63]) );
  XOR U320 ( .A(a[64]), .B(b[64]), .Z(n256) );
  NAND U321 ( .A(b[63]), .B(a[63]), .Z(n255) );
  NANDN U322 ( .A(n253), .B(n252), .Z(n254) );
  AND U323 ( .A(n255), .B(n254), .Z(n257) );
  XNOR U324 ( .A(n256), .B(n257), .Z(c[64]) );
  XOR U325 ( .A(a[65]), .B(b[65]), .Z(n260) );
  NAND U326 ( .A(b[64]), .B(a[64]), .Z(n259) );
  NANDN U327 ( .A(n257), .B(n256), .Z(n258) );
  AND U328 ( .A(n259), .B(n258), .Z(n261) );
  XNOR U329 ( .A(n260), .B(n261), .Z(c[65]) );
  XOR U330 ( .A(a[66]), .B(b[66]), .Z(n264) );
  NAND U331 ( .A(b[65]), .B(a[65]), .Z(n263) );
  NANDN U332 ( .A(n261), .B(n260), .Z(n262) );
  AND U333 ( .A(n263), .B(n262), .Z(n265) );
  XNOR U334 ( .A(n264), .B(n265), .Z(c[66]) );
  XOR U335 ( .A(a[67]), .B(b[67]), .Z(n268) );
  NAND U336 ( .A(b[66]), .B(a[66]), .Z(n267) );
  NANDN U337 ( .A(n265), .B(n264), .Z(n266) );
  AND U338 ( .A(n267), .B(n266), .Z(n269) );
  XNOR U339 ( .A(n268), .B(n269), .Z(c[67]) );
  XOR U340 ( .A(a[68]), .B(b[68]), .Z(n272) );
  NAND U341 ( .A(b[67]), .B(a[67]), .Z(n271) );
  NANDN U342 ( .A(n269), .B(n268), .Z(n270) );
  AND U343 ( .A(n271), .B(n270), .Z(n273) );
  XNOR U344 ( .A(n272), .B(n273), .Z(c[68]) );
  XOR U345 ( .A(a[69]), .B(b[69]), .Z(n276) );
  NAND U346 ( .A(b[68]), .B(a[68]), .Z(n275) );
  NANDN U347 ( .A(n273), .B(n272), .Z(n274) );
  AND U348 ( .A(n275), .B(n274), .Z(n277) );
  XNOR U349 ( .A(n276), .B(n277), .Z(c[69]) );
  XOR U350 ( .A(a[70]), .B(b[70]), .Z(n280) );
  NAND U351 ( .A(b[69]), .B(a[69]), .Z(n279) );
  NANDN U352 ( .A(n277), .B(n276), .Z(n278) );
  AND U353 ( .A(n279), .B(n278), .Z(n281) );
  XNOR U354 ( .A(n280), .B(n281), .Z(c[70]) );
  XOR U355 ( .A(a[71]), .B(b[71]), .Z(n284) );
  NAND U356 ( .A(b[70]), .B(a[70]), .Z(n283) );
  NANDN U357 ( .A(n281), .B(n280), .Z(n282) );
  AND U358 ( .A(n283), .B(n282), .Z(n285) );
  XNOR U359 ( .A(n284), .B(n285), .Z(c[71]) );
  XOR U360 ( .A(a[72]), .B(b[72]), .Z(n288) );
  NAND U361 ( .A(b[71]), .B(a[71]), .Z(n287) );
  NANDN U362 ( .A(n285), .B(n284), .Z(n286) );
  AND U363 ( .A(n287), .B(n286), .Z(n289) );
  XNOR U364 ( .A(n288), .B(n289), .Z(c[72]) );
  XOR U365 ( .A(a[73]), .B(b[73]), .Z(n292) );
  NAND U366 ( .A(b[72]), .B(a[72]), .Z(n291) );
  NANDN U367 ( .A(n289), .B(n288), .Z(n290) );
  AND U368 ( .A(n291), .B(n290), .Z(n293) );
  XNOR U369 ( .A(n292), .B(n293), .Z(c[73]) );
  XOR U370 ( .A(a[74]), .B(b[74]), .Z(n296) );
  NAND U371 ( .A(b[73]), .B(a[73]), .Z(n295) );
  NANDN U372 ( .A(n293), .B(n292), .Z(n294) );
  AND U373 ( .A(n295), .B(n294), .Z(n297) );
  XNOR U374 ( .A(n296), .B(n297), .Z(c[74]) );
  XOR U375 ( .A(a[75]), .B(b[75]), .Z(n300) );
  NAND U376 ( .A(b[74]), .B(a[74]), .Z(n299) );
  NANDN U377 ( .A(n297), .B(n296), .Z(n298) );
  AND U378 ( .A(n299), .B(n298), .Z(n301) );
  XNOR U379 ( .A(n300), .B(n301), .Z(c[75]) );
  XOR U380 ( .A(a[76]), .B(b[76]), .Z(n304) );
  NAND U381 ( .A(b[75]), .B(a[75]), .Z(n303) );
  NANDN U382 ( .A(n301), .B(n300), .Z(n302) );
  AND U383 ( .A(n303), .B(n302), .Z(n305) );
  XNOR U384 ( .A(n304), .B(n305), .Z(c[76]) );
  XOR U385 ( .A(a[77]), .B(b[77]), .Z(n308) );
  NAND U386 ( .A(b[76]), .B(a[76]), .Z(n307) );
  NANDN U387 ( .A(n305), .B(n304), .Z(n306) );
  AND U388 ( .A(n307), .B(n306), .Z(n309) );
  XNOR U389 ( .A(n308), .B(n309), .Z(c[77]) );
  XOR U390 ( .A(a[78]), .B(b[78]), .Z(n312) );
  NAND U391 ( .A(b[77]), .B(a[77]), .Z(n311) );
  NANDN U392 ( .A(n309), .B(n308), .Z(n310) );
  AND U393 ( .A(n311), .B(n310), .Z(n313) );
  XNOR U394 ( .A(n312), .B(n313), .Z(c[78]) );
  XOR U395 ( .A(a[79]), .B(b[79]), .Z(n316) );
  NAND U396 ( .A(b[78]), .B(a[78]), .Z(n315) );
  NANDN U397 ( .A(n313), .B(n312), .Z(n314) );
  AND U398 ( .A(n315), .B(n314), .Z(n317) );
  XNOR U399 ( .A(n316), .B(n317), .Z(c[79]) );
  XOR U400 ( .A(a[80]), .B(b[80]), .Z(n320) );
  NAND U401 ( .A(b[79]), .B(a[79]), .Z(n319) );
  NANDN U402 ( .A(n317), .B(n316), .Z(n318) );
  AND U403 ( .A(n319), .B(n318), .Z(n321) );
  XNOR U404 ( .A(n320), .B(n321), .Z(c[80]) );
  XOR U405 ( .A(a[81]), .B(b[81]), .Z(n324) );
  NAND U406 ( .A(b[80]), .B(a[80]), .Z(n323) );
  NANDN U407 ( .A(n321), .B(n320), .Z(n322) );
  AND U408 ( .A(n323), .B(n322), .Z(n325) );
  XNOR U409 ( .A(n324), .B(n325), .Z(c[81]) );
  XOR U410 ( .A(a[82]), .B(b[82]), .Z(n328) );
  NAND U411 ( .A(b[81]), .B(a[81]), .Z(n327) );
  NANDN U412 ( .A(n325), .B(n324), .Z(n326) );
  AND U413 ( .A(n327), .B(n326), .Z(n329) );
  XNOR U414 ( .A(n328), .B(n329), .Z(c[82]) );
  XOR U415 ( .A(a[83]), .B(b[83]), .Z(n332) );
  NAND U416 ( .A(b[82]), .B(a[82]), .Z(n331) );
  NANDN U417 ( .A(n329), .B(n328), .Z(n330) );
  AND U418 ( .A(n331), .B(n330), .Z(n333) );
  XNOR U419 ( .A(n332), .B(n333), .Z(c[83]) );
  XOR U420 ( .A(a[84]), .B(b[84]), .Z(n336) );
  NAND U421 ( .A(b[83]), .B(a[83]), .Z(n335) );
  NANDN U422 ( .A(n333), .B(n332), .Z(n334) );
  AND U423 ( .A(n335), .B(n334), .Z(n337) );
  XNOR U424 ( .A(n336), .B(n337), .Z(c[84]) );
  XOR U425 ( .A(a[85]), .B(b[85]), .Z(n340) );
  NAND U426 ( .A(b[84]), .B(a[84]), .Z(n339) );
  NANDN U427 ( .A(n337), .B(n336), .Z(n338) );
  AND U428 ( .A(n339), .B(n338), .Z(n341) );
  XNOR U429 ( .A(n340), .B(n341), .Z(c[85]) );
  XOR U430 ( .A(a[86]), .B(b[86]), .Z(n344) );
  NAND U431 ( .A(b[85]), .B(a[85]), .Z(n343) );
  NANDN U432 ( .A(n341), .B(n340), .Z(n342) );
  AND U433 ( .A(n343), .B(n342), .Z(n345) );
  XNOR U434 ( .A(n344), .B(n345), .Z(c[86]) );
  XOR U435 ( .A(a[87]), .B(b[87]), .Z(n348) );
  NAND U436 ( .A(b[86]), .B(a[86]), .Z(n347) );
  NANDN U437 ( .A(n345), .B(n344), .Z(n346) );
  AND U438 ( .A(n347), .B(n346), .Z(n349) );
  XNOR U439 ( .A(n348), .B(n349), .Z(c[87]) );
  XOR U440 ( .A(a[88]), .B(b[88]), .Z(n352) );
  NAND U441 ( .A(b[87]), .B(a[87]), .Z(n351) );
  NANDN U442 ( .A(n349), .B(n348), .Z(n350) );
  AND U443 ( .A(n351), .B(n350), .Z(n353) );
  XNOR U444 ( .A(n352), .B(n353), .Z(c[88]) );
  XOR U445 ( .A(a[89]), .B(b[89]), .Z(n356) );
  NAND U446 ( .A(b[88]), .B(a[88]), .Z(n355) );
  NANDN U447 ( .A(n353), .B(n352), .Z(n354) );
  AND U448 ( .A(n355), .B(n354), .Z(n357) );
  XNOR U449 ( .A(n356), .B(n357), .Z(c[89]) );
  XOR U450 ( .A(a[90]), .B(b[90]), .Z(n360) );
  NAND U451 ( .A(b[89]), .B(a[89]), .Z(n359) );
  NANDN U452 ( .A(n357), .B(n356), .Z(n358) );
  AND U453 ( .A(n359), .B(n358), .Z(n361) );
  XNOR U454 ( .A(n360), .B(n361), .Z(c[90]) );
  XOR U455 ( .A(a[91]), .B(b[91]), .Z(n364) );
  NAND U456 ( .A(b[90]), .B(a[90]), .Z(n363) );
  NANDN U457 ( .A(n361), .B(n360), .Z(n362) );
  AND U458 ( .A(n363), .B(n362), .Z(n365) );
  XNOR U459 ( .A(n364), .B(n365), .Z(c[91]) );
  XOR U460 ( .A(a[92]), .B(b[92]), .Z(n368) );
  NAND U461 ( .A(b[91]), .B(a[91]), .Z(n367) );
  NANDN U462 ( .A(n365), .B(n364), .Z(n366) );
  AND U463 ( .A(n367), .B(n366), .Z(n369) );
  XNOR U464 ( .A(n368), .B(n369), .Z(c[92]) );
  XOR U465 ( .A(a[93]), .B(b[93]), .Z(n372) );
  NAND U466 ( .A(b[92]), .B(a[92]), .Z(n371) );
  NANDN U467 ( .A(n369), .B(n368), .Z(n370) );
  AND U468 ( .A(n371), .B(n370), .Z(n373) );
  XNOR U469 ( .A(n372), .B(n373), .Z(c[93]) );
  XOR U470 ( .A(a[94]), .B(b[94]), .Z(n376) );
  NAND U471 ( .A(b[93]), .B(a[93]), .Z(n375) );
  NANDN U472 ( .A(n373), .B(n372), .Z(n374) );
  AND U473 ( .A(n375), .B(n374), .Z(n377) );
  XNOR U474 ( .A(n376), .B(n377), .Z(c[94]) );
  XOR U475 ( .A(a[95]), .B(b[95]), .Z(n380) );
  NAND U476 ( .A(b[94]), .B(a[94]), .Z(n379) );
  NANDN U477 ( .A(n377), .B(n376), .Z(n378) );
  AND U478 ( .A(n379), .B(n378), .Z(n381) );
  XNOR U479 ( .A(n380), .B(n381), .Z(c[95]) );
  XOR U480 ( .A(a[96]), .B(b[96]), .Z(n384) );
  NAND U481 ( .A(b[95]), .B(a[95]), .Z(n383) );
  NANDN U482 ( .A(n381), .B(n380), .Z(n382) );
  AND U483 ( .A(n383), .B(n382), .Z(n385) );
  XNOR U484 ( .A(n384), .B(n385), .Z(c[96]) );
  XOR U485 ( .A(a[97]), .B(b[97]), .Z(n388) );
  NAND U486 ( .A(b[96]), .B(a[96]), .Z(n387) );
  NANDN U487 ( .A(n385), .B(n384), .Z(n386) );
  AND U488 ( .A(n387), .B(n386), .Z(n389) );
  XNOR U489 ( .A(n388), .B(n389), .Z(c[97]) );
  XOR U490 ( .A(a[98]), .B(b[98]), .Z(n392) );
  NAND U491 ( .A(b[97]), .B(a[97]), .Z(n391) );
  NANDN U492 ( .A(n389), .B(n388), .Z(n390) );
  AND U493 ( .A(n391), .B(n390), .Z(n393) );
  XNOR U494 ( .A(n392), .B(n393), .Z(c[98]) );
  XOR U495 ( .A(a[99]), .B(b[99]), .Z(n396) );
  NAND U496 ( .A(b[98]), .B(a[98]), .Z(n395) );
  NANDN U497 ( .A(n393), .B(n392), .Z(n394) );
  AND U498 ( .A(n395), .B(n394), .Z(n397) );
  XNOR U499 ( .A(n396), .B(n397), .Z(c[99]) );
  XOR U500 ( .A(a[100]), .B(b[100]), .Z(n400) );
  NAND U501 ( .A(b[99]), .B(a[99]), .Z(n399) );
  NANDN U502 ( .A(n397), .B(n396), .Z(n398) );
  AND U503 ( .A(n399), .B(n398), .Z(n401) );
  XNOR U504 ( .A(n400), .B(n401), .Z(c[100]) );
  XOR U505 ( .A(a[101]), .B(b[101]), .Z(n404) );
  NAND U506 ( .A(b[100]), .B(a[100]), .Z(n403) );
  NANDN U507 ( .A(n401), .B(n400), .Z(n402) );
  AND U508 ( .A(n403), .B(n402), .Z(n405) );
  XNOR U509 ( .A(n404), .B(n405), .Z(c[101]) );
  XOR U510 ( .A(a[102]), .B(b[102]), .Z(n408) );
  NAND U511 ( .A(b[101]), .B(a[101]), .Z(n407) );
  NANDN U512 ( .A(n405), .B(n404), .Z(n406) );
  AND U513 ( .A(n407), .B(n406), .Z(n409) );
  XNOR U514 ( .A(n408), .B(n409), .Z(c[102]) );
  XOR U515 ( .A(a[103]), .B(b[103]), .Z(n412) );
  NAND U516 ( .A(b[102]), .B(a[102]), .Z(n411) );
  NANDN U517 ( .A(n409), .B(n408), .Z(n410) );
  AND U518 ( .A(n411), .B(n410), .Z(n413) );
  XNOR U519 ( .A(n412), .B(n413), .Z(c[103]) );
  XOR U520 ( .A(a[104]), .B(b[104]), .Z(n416) );
  NAND U521 ( .A(b[103]), .B(a[103]), .Z(n415) );
  NANDN U522 ( .A(n413), .B(n412), .Z(n414) );
  AND U523 ( .A(n415), .B(n414), .Z(n417) );
  XNOR U524 ( .A(n416), .B(n417), .Z(c[104]) );
  XOR U525 ( .A(a[105]), .B(b[105]), .Z(n420) );
  NAND U526 ( .A(b[104]), .B(a[104]), .Z(n419) );
  NANDN U527 ( .A(n417), .B(n416), .Z(n418) );
  AND U528 ( .A(n419), .B(n418), .Z(n421) );
  XNOR U529 ( .A(n420), .B(n421), .Z(c[105]) );
  XOR U530 ( .A(a[106]), .B(b[106]), .Z(n424) );
  NAND U531 ( .A(b[105]), .B(a[105]), .Z(n423) );
  NANDN U532 ( .A(n421), .B(n420), .Z(n422) );
  AND U533 ( .A(n423), .B(n422), .Z(n425) );
  XNOR U534 ( .A(n424), .B(n425), .Z(c[106]) );
  XOR U535 ( .A(a[107]), .B(b[107]), .Z(n428) );
  NAND U536 ( .A(b[106]), .B(a[106]), .Z(n427) );
  NANDN U537 ( .A(n425), .B(n424), .Z(n426) );
  AND U538 ( .A(n427), .B(n426), .Z(n429) );
  XNOR U539 ( .A(n428), .B(n429), .Z(c[107]) );
  XOR U540 ( .A(a[108]), .B(b[108]), .Z(n432) );
  NAND U541 ( .A(b[107]), .B(a[107]), .Z(n431) );
  NANDN U542 ( .A(n429), .B(n428), .Z(n430) );
  AND U543 ( .A(n431), .B(n430), .Z(n433) );
  XNOR U544 ( .A(n432), .B(n433), .Z(c[108]) );
  XOR U545 ( .A(a[109]), .B(b[109]), .Z(n436) );
  NAND U546 ( .A(b[108]), .B(a[108]), .Z(n435) );
  NANDN U547 ( .A(n433), .B(n432), .Z(n434) );
  AND U548 ( .A(n435), .B(n434), .Z(n437) );
  XNOR U549 ( .A(n436), .B(n437), .Z(c[109]) );
  XOR U550 ( .A(a[110]), .B(b[110]), .Z(n440) );
  NAND U551 ( .A(b[109]), .B(a[109]), .Z(n439) );
  NANDN U552 ( .A(n437), .B(n436), .Z(n438) );
  AND U553 ( .A(n439), .B(n438), .Z(n441) );
  XNOR U554 ( .A(n440), .B(n441), .Z(c[110]) );
  XOR U555 ( .A(a[111]), .B(b[111]), .Z(n444) );
  NAND U556 ( .A(b[110]), .B(a[110]), .Z(n443) );
  NANDN U557 ( .A(n441), .B(n440), .Z(n442) );
  AND U558 ( .A(n443), .B(n442), .Z(n445) );
  XNOR U559 ( .A(n444), .B(n445), .Z(c[111]) );
  XOR U560 ( .A(a[112]), .B(b[112]), .Z(n448) );
  NAND U561 ( .A(b[111]), .B(a[111]), .Z(n447) );
  NANDN U562 ( .A(n445), .B(n444), .Z(n446) );
  AND U563 ( .A(n447), .B(n446), .Z(n449) );
  XNOR U564 ( .A(n448), .B(n449), .Z(c[112]) );
  XOR U565 ( .A(a[113]), .B(b[113]), .Z(n452) );
  NAND U566 ( .A(b[112]), .B(a[112]), .Z(n451) );
  NANDN U567 ( .A(n449), .B(n448), .Z(n450) );
  AND U568 ( .A(n451), .B(n450), .Z(n453) );
  XNOR U569 ( .A(n452), .B(n453), .Z(c[113]) );
  XOR U570 ( .A(a[114]), .B(b[114]), .Z(n456) );
  NAND U571 ( .A(b[113]), .B(a[113]), .Z(n455) );
  NANDN U572 ( .A(n453), .B(n452), .Z(n454) );
  AND U573 ( .A(n455), .B(n454), .Z(n457) );
  XNOR U574 ( .A(n456), .B(n457), .Z(c[114]) );
  XOR U575 ( .A(a[115]), .B(b[115]), .Z(n460) );
  NAND U576 ( .A(b[114]), .B(a[114]), .Z(n459) );
  NANDN U577 ( .A(n457), .B(n456), .Z(n458) );
  AND U578 ( .A(n459), .B(n458), .Z(n461) );
  XNOR U579 ( .A(n460), .B(n461), .Z(c[115]) );
  XOR U580 ( .A(a[116]), .B(b[116]), .Z(n464) );
  NAND U581 ( .A(b[115]), .B(a[115]), .Z(n463) );
  NANDN U582 ( .A(n461), .B(n460), .Z(n462) );
  AND U583 ( .A(n463), .B(n462), .Z(n465) );
  XNOR U584 ( .A(n464), .B(n465), .Z(c[116]) );
  XOR U585 ( .A(a[117]), .B(b[117]), .Z(n468) );
  NAND U586 ( .A(b[116]), .B(a[116]), .Z(n467) );
  NANDN U587 ( .A(n465), .B(n464), .Z(n466) );
  AND U588 ( .A(n467), .B(n466), .Z(n469) );
  XNOR U589 ( .A(n468), .B(n469), .Z(c[117]) );
  XOR U590 ( .A(a[118]), .B(b[118]), .Z(n472) );
  NAND U591 ( .A(b[117]), .B(a[117]), .Z(n471) );
  NANDN U592 ( .A(n469), .B(n468), .Z(n470) );
  AND U593 ( .A(n471), .B(n470), .Z(n473) );
  XNOR U594 ( .A(n472), .B(n473), .Z(c[118]) );
  XOR U595 ( .A(a[119]), .B(b[119]), .Z(n476) );
  NAND U596 ( .A(b[118]), .B(a[118]), .Z(n475) );
  NANDN U597 ( .A(n473), .B(n472), .Z(n474) );
  AND U598 ( .A(n475), .B(n474), .Z(n477) );
  XNOR U599 ( .A(n476), .B(n477), .Z(c[119]) );
  XOR U600 ( .A(a[120]), .B(b[120]), .Z(n480) );
  NAND U601 ( .A(b[119]), .B(a[119]), .Z(n479) );
  NANDN U602 ( .A(n477), .B(n476), .Z(n478) );
  AND U603 ( .A(n479), .B(n478), .Z(n481) );
  XNOR U604 ( .A(n480), .B(n481), .Z(c[120]) );
  XOR U605 ( .A(a[121]), .B(b[121]), .Z(n484) );
  NAND U606 ( .A(b[120]), .B(a[120]), .Z(n483) );
  NANDN U607 ( .A(n481), .B(n480), .Z(n482) );
  AND U608 ( .A(n483), .B(n482), .Z(n485) );
  XNOR U609 ( .A(n484), .B(n485), .Z(c[121]) );
  XOR U610 ( .A(a[122]), .B(b[122]), .Z(n488) );
  NAND U611 ( .A(b[121]), .B(a[121]), .Z(n487) );
  NANDN U612 ( .A(n485), .B(n484), .Z(n486) );
  AND U613 ( .A(n487), .B(n486), .Z(n489) );
  XNOR U614 ( .A(n488), .B(n489), .Z(c[122]) );
  XOR U615 ( .A(a[123]), .B(b[123]), .Z(n492) );
  NAND U616 ( .A(b[122]), .B(a[122]), .Z(n491) );
  NANDN U617 ( .A(n489), .B(n488), .Z(n490) );
  AND U618 ( .A(n491), .B(n490), .Z(n493) );
  XNOR U619 ( .A(n492), .B(n493), .Z(c[123]) );
  XOR U620 ( .A(a[124]), .B(b[124]), .Z(n496) );
  NAND U621 ( .A(b[123]), .B(a[123]), .Z(n495) );
  NANDN U622 ( .A(n493), .B(n492), .Z(n494) );
  AND U623 ( .A(n495), .B(n494), .Z(n497) );
  XNOR U624 ( .A(n496), .B(n497), .Z(c[124]) );
  XOR U625 ( .A(a[125]), .B(b[125]), .Z(n500) );
  NAND U626 ( .A(b[124]), .B(a[124]), .Z(n499) );
  NANDN U627 ( .A(n497), .B(n496), .Z(n498) );
  AND U628 ( .A(n499), .B(n498), .Z(n501) );
  XNOR U629 ( .A(n500), .B(n501), .Z(c[125]) );
  XOR U630 ( .A(a[126]), .B(b[126]), .Z(n504) );
  NAND U631 ( .A(b[125]), .B(a[125]), .Z(n503) );
  NANDN U632 ( .A(n501), .B(n500), .Z(n502) );
  AND U633 ( .A(n503), .B(n502), .Z(n505) );
  XNOR U634 ( .A(n504), .B(n505), .Z(c[126]) );
  NAND U635 ( .A(b[126]), .B(a[126]), .Z(n507) );
  NANDN U636 ( .A(n505), .B(n504), .Z(n506) );
  NAND U637 ( .A(n507), .B(n506), .Z(n508) );
  XOR U638 ( .A(a[127]), .B(b[127]), .Z(n509) );
  XOR U639 ( .A(n508), .B(n509), .Z(c[127]) );
  NAND U640 ( .A(b[127]), .B(a[127]), .Z(n511) );
  NAND U641 ( .A(n509), .B(n508), .Z(n510) );
  NAND U642 ( .A(n511), .B(n510), .Z(carry_on_d) );
endmodule

