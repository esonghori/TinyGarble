
module sum_N1024_CC2 ( clk, rst, a, b, c );
  input [511:0] a;
  input [511:0] b;
  output [511:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(carry_on), .B(a[0]), .Z(n1) );
  NAND U4 ( .A(n1), .B(b[0]), .Z(n2) );
  NAND U5 ( .A(carry_on), .B(a[0]), .Z(n3) );
  AND U6 ( .A(n2), .B(n3), .Z(n12) );
  NAND U7 ( .A(a[502]), .B(n2016), .Z(n4) );
  XOR U8 ( .A(a[502]), .B(n2016), .Z(n5) );
  NAND U9 ( .A(n5), .B(b[502]), .Z(n6) );
  NAND U10 ( .A(n4), .B(n6), .Z(n2018) );
  NAND U11 ( .A(b[511]), .B(n2050), .Z(n7) );
  XOR U12 ( .A(b[511]), .B(n2050), .Z(n8) );
  NAND U13 ( .A(n8), .B(a[511]), .Z(n9) );
  NAND U14 ( .A(n7), .B(n9), .Z(carry_on_d) );
  XNOR U15 ( .A(b[0]), .B(a[0]), .Z(n10) );
  XNOR U16 ( .A(carry_on), .B(n10), .Z(c[0]) );
  XOR U17 ( .A(a[1]), .B(b[1]), .Z(n11) );
  XNOR U18 ( .A(n12), .B(n11), .Z(c[1]) );
  XOR U19 ( .A(a[2]), .B(b[2]), .Z(n16) );
  NAND U20 ( .A(a[1]), .B(b[1]), .Z(n14) );
  NANDN U21 ( .A(n12), .B(n11), .Z(n13) );
  NAND U22 ( .A(n14), .B(n13), .Z(n15) );
  XOR U23 ( .A(n16), .B(n15), .Z(c[2]) );
  XOR U24 ( .A(a[3]), .B(b[3]), .Z(n20) );
  NAND U25 ( .A(a[2]), .B(b[2]), .Z(n18) );
  NAND U26 ( .A(n16), .B(n15), .Z(n17) );
  NAND U27 ( .A(n18), .B(n17), .Z(n19) );
  XOR U28 ( .A(n20), .B(n19), .Z(c[3]) );
  XOR U29 ( .A(a[4]), .B(b[4]), .Z(n24) );
  NAND U30 ( .A(a[3]), .B(b[3]), .Z(n22) );
  NAND U31 ( .A(n20), .B(n19), .Z(n21) );
  NAND U32 ( .A(n22), .B(n21), .Z(n23) );
  XOR U33 ( .A(n24), .B(n23), .Z(c[4]) );
  XOR U34 ( .A(a[5]), .B(b[5]), .Z(n28) );
  NAND U35 ( .A(a[4]), .B(b[4]), .Z(n26) );
  NAND U36 ( .A(n24), .B(n23), .Z(n25) );
  NAND U37 ( .A(n26), .B(n25), .Z(n27) );
  XOR U38 ( .A(n28), .B(n27), .Z(c[5]) );
  XOR U39 ( .A(a[6]), .B(b[6]), .Z(n32) );
  NAND U40 ( .A(a[5]), .B(b[5]), .Z(n30) );
  NAND U41 ( .A(n28), .B(n27), .Z(n29) );
  NAND U42 ( .A(n30), .B(n29), .Z(n31) );
  XOR U43 ( .A(n32), .B(n31), .Z(c[6]) );
  XOR U44 ( .A(a[7]), .B(b[7]), .Z(n36) );
  NAND U45 ( .A(a[6]), .B(b[6]), .Z(n34) );
  NAND U46 ( .A(n32), .B(n31), .Z(n33) );
  NAND U47 ( .A(n34), .B(n33), .Z(n35) );
  XOR U48 ( .A(n36), .B(n35), .Z(c[7]) );
  XOR U49 ( .A(b[8]), .B(a[8]), .Z(n40) );
  NAND U50 ( .A(a[7]), .B(b[7]), .Z(n38) );
  NAND U51 ( .A(n36), .B(n35), .Z(n37) );
  AND U52 ( .A(n38), .B(n37), .Z(n39) );
  XNOR U53 ( .A(n40), .B(n39), .Z(c[8]) );
  XOR U54 ( .A(b[9]), .B(a[9]), .Z(n44) );
  OR U55 ( .A(b[8]), .B(a[8]), .Z(n42) );
  NAND U56 ( .A(n40), .B(n39), .Z(n41) );
  NAND U57 ( .A(n42), .B(n41), .Z(n43) );
  XNOR U58 ( .A(n44), .B(n43), .Z(c[9]) );
  XOR U59 ( .A(a[10]), .B(b[10]), .Z(n48) );
  OR U60 ( .A(b[9]), .B(a[9]), .Z(n46) );
  NAND U61 ( .A(n44), .B(n43), .Z(n45) );
  AND U62 ( .A(n46), .B(n45), .Z(n47) );
  XOR U63 ( .A(n48), .B(n47), .Z(c[10]) );
  NAND U64 ( .A(a[10]), .B(b[10]), .Z(n50) );
  NAND U65 ( .A(n48), .B(n47), .Z(n49) );
  AND U66 ( .A(n50), .B(n49), .Z(n52) );
  XOR U67 ( .A(b[11]), .B(a[11]), .Z(n51) );
  XNOR U68 ( .A(n52), .B(n51), .Z(c[11]) );
  OR U69 ( .A(b[11]), .B(a[11]), .Z(n54) );
  NAND U70 ( .A(n52), .B(n51), .Z(n53) );
  AND U71 ( .A(n54), .B(n53), .Z(n56) );
  XOR U72 ( .A(a[12]), .B(b[12]), .Z(n55) );
  XOR U73 ( .A(n56), .B(n55), .Z(c[12]) );
  XOR U74 ( .A(a[13]), .B(b[13]), .Z(n60) );
  NAND U75 ( .A(a[12]), .B(b[12]), .Z(n58) );
  NAND U76 ( .A(n56), .B(n55), .Z(n57) );
  NAND U77 ( .A(n58), .B(n57), .Z(n59) );
  XOR U78 ( .A(n60), .B(n59), .Z(c[13]) );
  XOR U79 ( .A(a[14]), .B(b[14]), .Z(n64) );
  NAND U80 ( .A(a[13]), .B(b[13]), .Z(n62) );
  NAND U81 ( .A(n60), .B(n59), .Z(n61) );
  NAND U82 ( .A(n62), .B(n61), .Z(n63) );
  XOR U83 ( .A(n64), .B(n63), .Z(c[14]) );
  XOR U84 ( .A(a[15]), .B(b[15]), .Z(n68) );
  NAND U85 ( .A(a[14]), .B(b[14]), .Z(n66) );
  NAND U86 ( .A(n64), .B(n63), .Z(n65) );
  NAND U87 ( .A(n66), .B(n65), .Z(n67) );
  XOR U88 ( .A(n68), .B(n67), .Z(c[15]) );
  XOR U89 ( .A(a[16]), .B(b[16]), .Z(n72) );
  NAND U90 ( .A(a[15]), .B(b[15]), .Z(n70) );
  NAND U91 ( .A(n68), .B(n67), .Z(n69) );
  NAND U92 ( .A(n70), .B(n69), .Z(n71) );
  XOR U93 ( .A(n72), .B(n71), .Z(c[16]) );
  XOR U94 ( .A(a[17]), .B(b[17]), .Z(n76) );
  NAND U95 ( .A(a[16]), .B(b[16]), .Z(n74) );
  NAND U96 ( .A(n72), .B(n71), .Z(n73) );
  NAND U97 ( .A(n74), .B(n73), .Z(n75) );
  XOR U98 ( .A(n76), .B(n75), .Z(c[17]) );
  XOR U99 ( .A(a[18]), .B(b[18]), .Z(n80) );
  NAND U100 ( .A(a[17]), .B(b[17]), .Z(n78) );
  NAND U101 ( .A(n76), .B(n75), .Z(n77) );
  NAND U102 ( .A(n78), .B(n77), .Z(n79) );
  XOR U103 ( .A(n80), .B(n79), .Z(c[18]) );
  XOR U104 ( .A(a[19]), .B(b[19]), .Z(n84) );
  NAND U105 ( .A(a[18]), .B(b[18]), .Z(n82) );
  NAND U106 ( .A(n80), .B(n79), .Z(n81) );
  NAND U107 ( .A(n82), .B(n81), .Z(n83) );
  XOR U108 ( .A(n84), .B(n83), .Z(c[19]) );
  XOR U109 ( .A(a[20]), .B(b[20]), .Z(n88) );
  NAND U110 ( .A(a[19]), .B(b[19]), .Z(n86) );
  NAND U111 ( .A(n84), .B(n83), .Z(n85) );
  NAND U112 ( .A(n86), .B(n85), .Z(n87) );
  XOR U113 ( .A(n88), .B(n87), .Z(c[20]) );
  XOR U114 ( .A(a[21]), .B(b[21]), .Z(n92) );
  NAND U115 ( .A(a[20]), .B(b[20]), .Z(n90) );
  NAND U116 ( .A(n88), .B(n87), .Z(n89) );
  NAND U117 ( .A(n90), .B(n89), .Z(n91) );
  XOR U118 ( .A(n92), .B(n91), .Z(c[21]) );
  XOR U119 ( .A(a[22]), .B(b[22]), .Z(n96) );
  NAND U120 ( .A(a[21]), .B(b[21]), .Z(n94) );
  NAND U121 ( .A(n92), .B(n91), .Z(n93) );
  NAND U122 ( .A(n94), .B(n93), .Z(n95) );
  XOR U123 ( .A(n96), .B(n95), .Z(c[22]) );
  XOR U124 ( .A(a[23]), .B(b[23]), .Z(n100) );
  NAND U125 ( .A(a[22]), .B(b[22]), .Z(n98) );
  NAND U126 ( .A(n96), .B(n95), .Z(n97) );
  NAND U127 ( .A(n98), .B(n97), .Z(n99) );
  XOR U128 ( .A(n100), .B(n99), .Z(c[23]) );
  XOR U129 ( .A(a[24]), .B(b[24]), .Z(n104) );
  NAND U130 ( .A(a[23]), .B(b[23]), .Z(n102) );
  NAND U131 ( .A(n100), .B(n99), .Z(n101) );
  NAND U132 ( .A(n102), .B(n101), .Z(n103) );
  XOR U133 ( .A(n104), .B(n103), .Z(c[24]) );
  XOR U134 ( .A(a[25]), .B(b[25]), .Z(n108) );
  NAND U135 ( .A(a[24]), .B(b[24]), .Z(n106) );
  NAND U136 ( .A(n104), .B(n103), .Z(n105) );
  NAND U137 ( .A(n106), .B(n105), .Z(n107) );
  XOR U138 ( .A(n108), .B(n107), .Z(c[25]) );
  XOR U139 ( .A(a[26]), .B(b[26]), .Z(n112) );
  NAND U140 ( .A(a[25]), .B(b[25]), .Z(n110) );
  NAND U141 ( .A(n108), .B(n107), .Z(n109) );
  NAND U142 ( .A(n110), .B(n109), .Z(n111) );
  XOR U143 ( .A(n112), .B(n111), .Z(c[26]) );
  XOR U144 ( .A(a[27]), .B(b[27]), .Z(n116) );
  NAND U145 ( .A(a[26]), .B(b[26]), .Z(n114) );
  NAND U146 ( .A(n112), .B(n111), .Z(n113) );
  NAND U147 ( .A(n114), .B(n113), .Z(n115) );
  XOR U148 ( .A(n116), .B(n115), .Z(c[27]) );
  XOR U149 ( .A(a[28]), .B(b[28]), .Z(n120) );
  NAND U150 ( .A(a[27]), .B(b[27]), .Z(n118) );
  NAND U151 ( .A(n116), .B(n115), .Z(n117) );
  NAND U152 ( .A(n118), .B(n117), .Z(n119) );
  XOR U153 ( .A(n120), .B(n119), .Z(c[28]) );
  XOR U154 ( .A(a[29]), .B(b[29]), .Z(n124) );
  NAND U155 ( .A(a[28]), .B(b[28]), .Z(n122) );
  NAND U156 ( .A(n120), .B(n119), .Z(n121) );
  NAND U157 ( .A(n122), .B(n121), .Z(n123) );
  XOR U158 ( .A(n124), .B(n123), .Z(c[29]) );
  XOR U159 ( .A(a[30]), .B(b[30]), .Z(n128) );
  NAND U160 ( .A(a[29]), .B(b[29]), .Z(n126) );
  NAND U161 ( .A(n124), .B(n123), .Z(n125) );
  NAND U162 ( .A(n126), .B(n125), .Z(n127) );
  XOR U163 ( .A(n128), .B(n127), .Z(c[30]) );
  XOR U164 ( .A(a[31]), .B(b[31]), .Z(n132) );
  NAND U165 ( .A(a[30]), .B(b[30]), .Z(n130) );
  NAND U166 ( .A(n128), .B(n127), .Z(n129) );
  NAND U167 ( .A(n130), .B(n129), .Z(n131) );
  XOR U168 ( .A(n132), .B(n131), .Z(c[31]) );
  XOR U169 ( .A(a[32]), .B(b[32]), .Z(n136) );
  NAND U170 ( .A(a[31]), .B(b[31]), .Z(n134) );
  NAND U171 ( .A(n132), .B(n131), .Z(n133) );
  NAND U172 ( .A(n134), .B(n133), .Z(n135) );
  XOR U173 ( .A(n136), .B(n135), .Z(c[32]) );
  XOR U174 ( .A(a[33]), .B(b[33]), .Z(n140) );
  NAND U175 ( .A(a[32]), .B(b[32]), .Z(n138) );
  NAND U176 ( .A(n136), .B(n135), .Z(n137) );
  NAND U177 ( .A(n138), .B(n137), .Z(n139) );
  XOR U178 ( .A(n140), .B(n139), .Z(c[33]) );
  XOR U179 ( .A(a[34]), .B(b[34]), .Z(n144) );
  NAND U180 ( .A(a[33]), .B(b[33]), .Z(n142) );
  NAND U181 ( .A(n140), .B(n139), .Z(n141) );
  NAND U182 ( .A(n142), .B(n141), .Z(n143) );
  XOR U183 ( .A(n144), .B(n143), .Z(c[34]) );
  XOR U184 ( .A(a[35]), .B(b[35]), .Z(n148) );
  NAND U185 ( .A(a[34]), .B(b[34]), .Z(n146) );
  NAND U186 ( .A(n144), .B(n143), .Z(n145) );
  NAND U187 ( .A(n146), .B(n145), .Z(n147) );
  XOR U188 ( .A(n148), .B(n147), .Z(c[35]) );
  XOR U189 ( .A(a[36]), .B(b[36]), .Z(n152) );
  NAND U190 ( .A(a[35]), .B(b[35]), .Z(n150) );
  NAND U191 ( .A(n148), .B(n147), .Z(n149) );
  NAND U192 ( .A(n150), .B(n149), .Z(n151) );
  XOR U193 ( .A(n152), .B(n151), .Z(c[36]) );
  XOR U194 ( .A(a[37]), .B(b[37]), .Z(n156) );
  NAND U195 ( .A(a[36]), .B(b[36]), .Z(n154) );
  NAND U196 ( .A(n152), .B(n151), .Z(n153) );
  NAND U197 ( .A(n154), .B(n153), .Z(n155) );
  XOR U198 ( .A(n156), .B(n155), .Z(c[37]) );
  XOR U199 ( .A(a[38]), .B(b[38]), .Z(n160) );
  NAND U200 ( .A(a[37]), .B(b[37]), .Z(n158) );
  NAND U201 ( .A(n156), .B(n155), .Z(n157) );
  NAND U202 ( .A(n158), .B(n157), .Z(n159) );
  XOR U203 ( .A(n160), .B(n159), .Z(c[38]) );
  XOR U204 ( .A(a[39]), .B(b[39]), .Z(n164) );
  NAND U205 ( .A(a[38]), .B(b[38]), .Z(n162) );
  NAND U206 ( .A(n160), .B(n159), .Z(n161) );
  NAND U207 ( .A(n162), .B(n161), .Z(n163) );
  XOR U208 ( .A(n164), .B(n163), .Z(c[39]) );
  XOR U209 ( .A(a[40]), .B(b[40]), .Z(n168) );
  NAND U210 ( .A(a[39]), .B(b[39]), .Z(n166) );
  NAND U211 ( .A(n164), .B(n163), .Z(n165) );
  NAND U212 ( .A(n166), .B(n165), .Z(n167) );
  XOR U213 ( .A(n168), .B(n167), .Z(c[40]) );
  XOR U214 ( .A(a[41]), .B(b[41]), .Z(n172) );
  NAND U215 ( .A(a[40]), .B(b[40]), .Z(n170) );
  NAND U216 ( .A(n168), .B(n167), .Z(n169) );
  NAND U217 ( .A(n170), .B(n169), .Z(n171) );
  XOR U218 ( .A(n172), .B(n171), .Z(c[41]) );
  XOR U219 ( .A(a[42]), .B(b[42]), .Z(n176) );
  NAND U220 ( .A(a[41]), .B(b[41]), .Z(n174) );
  NAND U221 ( .A(n172), .B(n171), .Z(n173) );
  NAND U222 ( .A(n174), .B(n173), .Z(n175) );
  XOR U223 ( .A(n176), .B(n175), .Z(c[42]) );
  XOR U224 ( .A(a[43]), .B(b[43]), .Z(n180) );
  NAND U225 ( .A(a[42]), .B(b[42]), .Z(n178) );
  NAND U226 ( .A(n176), .B(n175), .Z(n177) );
  NAND U227 ( .A(n178), .B(n177), .Z(n179) );
  XOR U228 ( .A(n180), .B(n179), .Z(c[43]) );
  XOR U229 ( .A(a[44]), .B(b[44]), .Z(n184) );
  NAND U230 ( .A(a[43]), .B(b[43]), .Z(n182) );
  NAND U231 ( .A(n180), .B(n179), .Z(n181) );
  NAND U232 ( .A(n182), .B(n181), .Z(n183) );
  XOR U233 ( .A(n184), .B(n183), .Z(c[44]) );
  XOR U234 ( .A(a[45]), .B(b[45]), .Z(n188) );
  NAND U235 ( .A(a[44]), .B(b[44]), .Z(n186) );
  NAND U236 ( .A(n184), .B(n183), .Z(n185) );
  NAND U237 ( .A(n186), .B(n185), .Z(n187) );
  XOR U238 ( .A(n188), .B(n187), .Z(c[45]) );
  XOR U239 ( .A(a[46]), .B(b[46]), .Z(n192) );
  NAND U240 ( .A(a[45]), .B(b[45]), .Z(n190) );
  NAND U241 ( .A(n188), .B(n187), .Z(n189) );
  NAND U242 ( .A(n190), .B(n189), .Z(n191) );
  XOR U243 ( .A(n192), .B(n191), .Z(c[46]) );
  XOR U244 ( .A(a[47]), .B(b[47]), .Z(n196) );
  NAND U245 ( .A(a[46]), .B(b[46]), .Z(n194) );
  NAND U246 ( .A(n192), .B(n191), .Z(n193) );
  NAND U247 ( .A(n194), .B(n193), .Z(n195) );
  XOR U248 ( .A(n196), .B(n195), .Z(c[47]) );
  XOR U249 ( .A(a[48]), .B(b[48]), .Z(n200) );
  NAND U250 ( .A(a[47]), .B(b[47]), .Z(n198) );
  NAND U251 ( .A(n196), .B(n195), .Z(n197) );
  NAND U252 ( .A(n198), .B(n197), .Z(n199) );
  XOR U253 ( .A(n200), .B(n199), .Z(c[48]) );
  XOR U254 ( .A(a[49]), .B(b[49]), .Z(n204) );
  NAND U255 ( .A(a[48]), .B(b[48]), .Z(n202) );
  NAND U256 ( .A(n200), .B(n199), .Z(n201) );
  NAND U257 ( .A(n202), .B(n201), .Z(n203) );
  XOR U258 ( .A(n204), .B(n203), .Z(c[49]) );
  XOR U259 ( .A(a[50]), .B(b[50]), .Z(n208) );
  NAND U260 ( .A(a[49]), .B(b[49]), .Z(n206) );
  NAND U261 ( .A(n204), .B(n203), .Z(n205) );
  NAND U262 ( .A(n206), .B(n205), .Z(n207) );
  XOR U263 ( .A(n208), .B(n207), .Z(c[50]) );
  XOR U264 ( .A(a[51]), .B(b[51]), .Z(n212) );
  NAND U265 ( .A(a[50]), .B(b[50]), .Z(n210) );
  NAND U266 ( .A(n208), .B(n207), .Z(n209) );
  NAND U267 ( .A(n210), .B(n209), .Z(n211) );
  XOR U268 ( .A(n212), .B(n211), .Z(c[51]) );
  XOR U269 ( .A(a[52]), .B(b[52]), .Z(n216) );
  NAND U270 ( .A(a[51]), .B(b[51]), .Z(n214) );
  NAND U271 ( .A(n212), .B(n211), .Z(n213) );
  NAND U272 ( .A(n214), .B(n213), .Z(n215) );
  XOR U273 ( .A(n216), .B(n215), .Z(c[52]) );
  XOR U274 ( .A(a[53]), .B(b[53]), .Z(n220) );
  NAND U275 ( .A(a[52]), .B(b[52]), .Z(n218) );
  NAND U276 ( .A(n216), .B(n215), .Z(n217) );
  NAND U277 ( .A(n218), .B(n217), .Z(n219) );
  XOR U278 ( .A(n220), .B(n219), .Z(c[53]) );
  XOR U279 ( .A(a[54]), .B(b[54]), .Z(n224) );
  NAND U280 ( .A(a[53]), .B(b[53]), .Z(n222) );
  NAND U281 ( .A(n220), .B(n219), .Z(n221) );
  NAND U282 ( .A(n222), .B(n221), .Z(n223) );
  XOR U283 ( .A(n224), .B(n223), .Z(c[54]) );
  XOR U284 ( .A(a[55]), .B(b[55]), .Z(n228) );
  NAND U285 ( .A(a[54]), .B(b[54]), .Z(n226) );
  NAND U286 ( .A(n224), .B(n223), .Z(n225) );
  NAND U287 ( .A(n226), .B(n225), .Z(n227) );
  XOR U288 ( .A(n228), .B(n227), .Z(c[55]) );
  XOR U289 ( .A(a[56]), .B(b[56]), .Z(n232) );
  NAND U290 ( .A(a[55]), .B(b[55]), .Z(n230) );
  NAND U291 ( .A(n228), .B(n227), .Z(n229) );
  NAND U292 ( .A(n230), .B(n229), .Z(n231) );
  XOR U293 ( .A(n232), .B(n231), .Z(c[56]) );
  XOR U294 ( .A(a[57]), .B(b[57]), .Z(n236) );
  NAND U295 ( .A(a[56]), .B(b[56]), .Z(n234) );
  NAND U296 ( .A(n232), .B(n231), .Z(n233) );
  NAND U297 ( .A(n234), .B(n233), .Z(n235) );
  XOR U298 ( .A(n236), .B(n235), .Z(c[57]) );
  XOR U299 ( .A(a[58]), .B(b[58]), .Z(n240) );
  NAND U300 ( .A(a[57]), .B(b[57]), .Z(n238) );
  NAND U301 ( .A(n236), .B(n235), .Z(n237) );
  NAND U302 ( .A(n238), .B(n237), .Z(n239) );
  XOR U303 ( .A(n240), .B(n239), .Z(c[58]) );
  XOR U304 ( .A(a[59]), .B(b[59]), .Z(n244) );
  NAND U305 ( .A(a[58]), .B(b[58]), .Z(n242) );
  NAND U306 ( .A(n240), .B(n239), .Z(n241) );
  NAND U307 ( .A(n242), .B(n241), .Z(n243) );
  XOR U308 ( .A(n244), .B(n243), .Z(c[59]) );
  XOR U309 ( .A(a[60]), .B(b[60]), .Z(n248) );
  NAND U310 ( .A(a[59]), .B(b[59]), .Z(n246) );
  NAND U311 ( .A(n244), .B(n243), .Z(n245) );
  NAND U312 ( .A(n246), .B(n245), .Z(n247) );
  XOR U313 ( .A(n248), .B(n247), .Z(c[60]) );
  XOR U314 ( .A(a[61]), .B(b[61]), .Z(n252) );
  NAND U315 ( .A(a[60]), .B(b[60]), .Z(n250) );
  NAND U316 ( .A(n248), .B(n247), .Z(n249) );
  NAND U317 ( .A(n250), .B(n249), .Z(n251) );
  XOR U318 ( .A(n252), .B(n251), .Z(c[61]) );
  XOR U319 ( .A(a[62]), .B(b[62]), .Z(n256) );
  NAND U320 ( .A(a[61]), .B(b[61]), .Z(n254) );
  NAND U321 ( .A(n252), .B(n251), .Z(n253) );
  NAND U322 ( .A(n254), .B(n253), .Z(n255) );
  XOR U323 ( .A(n256), .B(n255), .Z(c[62]) );
  XOR U324 ( .A(a[63]), .B(b[63]), .Z(n260) );
  NAND U325 ( .A(a[62]), .B(b[62]), .Z(n258) );
  NAND U326 ( .A(n256), .B(n255), .Z(n257) );
  NAND U327 ( .A(n258), .B(n257), .Z(n259) );
  XOR U328 ( .A(n260), .B(n259), .Z(c[63]) );
  XOR U329 ( .A(b[64]), .B(a[64]), .Z(n264) );
  NAND U330 ( .A(a[63]), .B(b[63]), .Z(n262) );
  NAND U331 ( .A(n260), .B(n259), .Z(n261) );
  AND U332 ( .A(n262), .B(n261), .Z(n263) );
  XNOR U333 ( .A(n264), .B(n263), .Z(c[64]) );
  XOR U334 ( .A(b[65]), .B(a[65]), .Z(n268) );
  OR U335 ( .A(b[64]), .B(a[64]), .Z(n266) );
  NAND U336 ( .A(n264), .B(n263), .Z(n265) );
  NAND U337 ( .A(n266), .B(n265), .Z(n267) );
  XNOR U338 ( .A(n268), .B(n267), .Z(c[65]) );
  OR U339 ( .A(b[65]), .B(a[65]), .Z(n270) );
  NAND U340 ( .A(n268), .B(n267), .Z(n269) );
  AND U341 ( .A(n270), .B(n269), .Z(n272) );
  XOR U342 ( .A(a[66]), .B(b[66]), .Z(n271) );
  XOR U343 ( .A(n272), .B(n271), .Z(c[66]) );
  XOR U344 ( .A(a[67]), .B(b[67]), .Z(n276) );
  NAND U345 ( .A(a[66]), .B(b[66]), .Z(n274) );
  NAND U346 ( .A(n272), .B(n271), .Z(n273) );
  NAND U347 ( .A(n274), .B(n273), .Z(n275) );
  XOR U348 ( .A(n276), .B(n275), .Z(c[67]) );
  XOR U349 ( .A(a[68]), .B(b[68]), .Z(n280) );
  NAND U350 ( .A(a[67]), .B(b[67]), .Z(n278) );
  NAND U351 ( .A(n276), .B(n275), .Z(n277) );
  NAND U352 ( .A(n278), .B(n277), .Z(n279) );
  XOR U353 ( .A(n280), .B(n279), .Z(c[68]) );
  XOR U354 ( .A(a[69]), .B(b[69]), .Z(n284) );
  NAND U355 ( .A(a[68]), .B(b[68]), .Z(n282) );
  NAND U356 ( .A(n280), .B(n279), .Z(n281) );
  NAND U357 ( .A(n282), .B(n281), .Z(n283) );
  XOR U358 ( .A(n284), .B(n283), .Z(c[69]) );
  XOR U359 ( .A(a[70]), .B(b[70]), .Z(n288) );
  NAND U360 ( .A(a[69]), .B(b[69]), .Z(n286) );
  NAND U361 ( .A(n284), .B(n283), .Z(n285) );
  NAND U362 ( .A(n286), .B(n285), .Z(n287) );
  XOR U363 ( .A(n288), .B(n287), .Z(c[70]) );
  XOR U364 ( .A(a[71]), .B(b[71]), .Z(n292) );
  NAND U365 ( .A(a[70]), .B(b[70]), .Z(n290) );
  NAND U366 ( .A(n288), .B(n287), .Z(n289) );
  NAND U367 ( .A(n290), .B(n289), .Z(n291) );
  XOR U368 ( .A(n292), .B(n291), .Z(c[71]) );
  XOR U369 ( .A(a[72]), .B(b[72]), .Z(n296) );
  NAND U370 ( .A(a[71]), .B(b[71]), .Z(n294) );
  NAND U371 ( .A(n292), .B(n291), .Z(n293) );
  NAND U372 ( .A(n294), .B(n293), .Z(n295) );
  XOR U373 ( .A(n296), .B(n295), .Z(c[72]) );
  XOR U374 ( .A(a[73]), .B(b[73]), .Z(n300) );
  NAND U375 ( .A(a[72]), .B(b[72]), .Z(n298) );
  NAND U376 ( .A(n296), .B(n295), .Z(n297) );
  NAND U377 ( .A(n298), .B(n297), .Z(n299) );
  XOR U378 ( .A(n300), .B(n299), .Z(c[73]) );
  XOR U379 ( .A(a[74]), .B(b[74]), .Z(n304) );
  NAND U380 ( .A(a[73]), .B(b[73]), .Z(n302) );
  NAND U381 ( .A(n300), .B(n299), .Z(n301) );
  NAND U382 ( .A(n302), .B(n301), .Z(n303) );
  XOR U383 ( .A(n304), .B(n303), .Z(c[74]) );
  XOR U384 ( .A(a[75]), .B(b[75]), .Z(n308) );
  NAND U385 ( .A(a[74]), .B(b[74]), .Z(n306) );
  NAND U386 ( .A(n304), .B(n303), .Z(n305) );
  NAND U387 ( .A(n306), .B(n305), .Z(n307) );
  XOR U388 ( .A(n308), .B(n307), .Z(c[75]) );
  XOR U389 ( .A(a[76]), .B(b[76]), .Z(n312) );
  NAND U390 ( .A(a[75]), .B(b[75]), .Z(n310) );
  NAND U391 ( .A(n308), .B(n307), .Z(n309) );
  NAND U392 ( .A(n310), .B(n309), .Z(n311) );
  XOR U393 ( .A(n312), .B(n311), .Z(c[76]) );
  XOR U394 ( .A(a[77]), .B(b[77]), .Z(n316) );
  NAND U395 ( .A(a[76]), .B(b[76]), .Z(n314) );
  NAND U396 ( .A(n312), .B(n311), .Z(n313) );
  NAND U397 ( .A(n314), .B(n313), .Z(n315) );
  XOR U398 ( .A(n316), .B(n315), .Z(c[77]) );
  XOR U399 ( .A(a[78]), .B(b[78]), .Z(n320) );
  NAND U400 ( .A(a[77]), .B(b[77]), .Z(n318) );
  NAND U401 ( .A(n316), .B(n315), .Z(n317) );
  NAND U402 ( .A(n318), .B(n317), .Z(n319) );
  XOR U403 ( .A(n320), .B(n319), .Z(c[78]) );
  XOR U404 ( .A(a[79]), .B(b[79]), .Z(n324) );
  NAND U405 ( .A(a[78]), .B(b[78]), .Z(n322) );
  NAND U406 ( .A(n320), .B(n319), .Z(n321) );
  NAND U407 ( .A(n322), .B(n321), .Z(n323) );
  XOR U408 ( .A(n324), .B(n323), .Z(c[79]) );
  XOR U409 ( .A(a[80]), .B(b[80]), .Z(n328) );
  NAND U410 ( .A(a[79]), .B(b[79]), .Z(n326) );
  NAND U411 ( .A(n324), .B(n323), .Z(n325) );
  NAND U412 ( .A(n326), .B(n325), .Z(n327) );
  XOR U413 ( .A(n328), .B(n327), .Z(c[80]) );
  XOR U414 ( .A(a[81]), .B(b[81]), .Z(n332) );
  NAND U415 ( .A(a[80]), .B(b[80]), .Z(n330) );
  NAND U416 ( .A(n328), .B(n327), .Z(n329) );
  NAND U417 ( .A(n330), .B(n329), .Z(n331) );
  XOR U418 ( .A(n332), .B(n331), .Z(c[81]) );
  XOR U419 ( .A(a[82]), .B(b[82]), .Z(n336) );
  NAND U420 ( .A(a[81]), .B(b[81]), .Z(n334) );
  NAND U421 ( .A(n332), .B(n331), .Z(n333) );
  NAND U422 ( .A(n334), .B(n333), .Z(n335) );
  XOR U423 ( .A(n336), .B(n335), .Z(c[82]) );
  XOR U424 ( .A(a[83]), .B(b[83]), .Z(n340) );
  NAND U425 ( .A(a[82]), .B(b[82]), .Z(n338) );
  NAND U426 ( .A(n336), .B(n335), .Z(n337) );
  NAND U427 ( .A(n338), .B(n337), .Z(n339) );
  XOR U428 ( .A(n340), .B(n339), .Z(c[83]) );
  XOR U429 ( .A(a[84]), .B(b[84]), .Z(n344) );
  NAND U430 ( .A(a[83]), .B(b[83]), .Z(n342) );
  NAND U431 ( .A(n340), .B(n339), .Z(n341) );
  NAND U432 ( .A(n342), .B(n341), .Z(n343) );
  XOR U433 ( .A(n344), .B(n343), .Z(c[84]) );
  XOR U434 ( .A(a[85]), .B(b[85]), .Z(n348) );
  NAND U435 ( .A(a[84]), .B(b[84]), .Z(n346) );
  NAND U436 ( .A(n344), .B(n343), .Z(n345) );
  NAND U437 ( .A(n346), .B(n345), .Z(n347) );
  XOR U438 ( .A(n348), .B(n347), .Z(c[85]) );
  XOR U439 ( .A(a[86]), .B(b[86]), .Z(n352) );
  NAND U440 ( .A(a[85]), .B(b[85]), .Z(n350) );
  NAND U441 ( .A(n348), .B(n347), .Z(n349) );
  NAND U442 ( .A(n350), .B(n349), .Z(n351) );
  XOR U443 ( .A(n352), .B(n351), .Z(c[86]) );
  XOR U444 ( .A(a[87]), .B(b[87]), .Z(n356) );
  NAND U445 ( .A(a[86]), .B(b[86]), .Z(n354) );
  NAND U446 ( .A(n352), .B(n351), .Z(n353) );
  NAND U447 ( .A(n354), .B(n353), .Z(n355) );
  XOR U448 ( .A(n356), .B(n355), .Z(c[87]) );
  XOR U449 ( .A(a[88]), .B(b[88]), .Z(n360) );
  NAND U450 ( .A(a[87]), .B(b[87]), .Z(n358) );
  NAND U451 ( .A(n356), .B(n355), .Z(n357) );
  NAND U452 ( .A(n358), .B(n357), .Z(n359) );
  XOR U453 ( .A(n360), .B(n359), .Z(c[88]) );
  XOR U454 ( .A(a[89]), .B(b[89]), .Z(n364) );
  NAND U455 ( .A(a[88]), .B(b[88]), .Z(n362) );
  NAND U456 ( .A(n360), .B(n359), .Z(n361) );
  NAND U457 ( .A(n362), .B(n361), .Z(n363) );
  XOR U458 ( .A(n364), .B(n363), .Z(c[89]) );
  XOR U459 ( .A(a[90]), .B(b[90]), .Z(n368) );
  NAND U460 ( .A(a[89]), .B(b[89]), .Z(n366) );
  NAND U461 ( .A(n364), .B(n363), .Z(n365) );
  NAND U462 ( .A(n366), .B(n365), .Z(n367) );
  XOR U463 ( .A(n368), .B(n367), .Z(c[90]) );
  XOR U464 ( .A(a[91]), .B(b[91]), .Z(n372) );
  NAND U465 ( .A(a[90]), .B(b[90]), .Z(n370) );
  NAND U466 ( .A(n368), .B(n367), .Z(n369) );
  NAND U467 ( .A(n370), .B(n369), .Z(n371) );
  XOR U468 ( .A(n372), .B(n371), .Z(c[91]) );
  XOR U469 ( .A(a[92]), .B(b[92]), .Z(n376) );
  NAND U470 ( .A(a[91]), .B(b[91]), .Z(n374) );
  NAND U471 ( .A(n372), .B(n371), .Z(n373) );
  NAND U472 ( .A(n374), .B(n373), .Z(n375) );
  XOR U473 ( .A(n376), .B(n375), .Z(c[92]) );
  XOR U474 ( .A(a[93]), .B(b[93]), .Z(n380) );
  NAND U475 ( .A(a[92]), .B(b[92]), .Z(n378) );
  NAND U476 ( .A(n376), .B(n375), .Z(n377) );
  NAND U477 ( .A(n378), .B(n377), .Z(n379) );
  XOR U478 ( .A(n380), .B(n379), .Z(c[93]) );
  XOR U479 ( .A(a[94]), .B(b[94]), .Z(n384) );
  NAND U480 ( .A(a[93]), .B(b[93]), .Z(n382) );
  NAND U481 ( .A(n380), .B(n379), .Z(n381) );
  NAND U482 ( .A(n382), .B(n381), .Z(n383) );
  XOR U483 ( .A(n384), .B(n383), .Z(c[94]) );
  XOR U484 ( .A(a[95]), .B(b[95]), .Z(n388) );
  NAND U485 ( .A(a[94]), .B(b[94]), .Z(n386) );
  NAND U486 ( .A(n384), .B(n383), .Z(n385) );
  NAND U487 ( .A(n386), .B(n385), .Z(n387) );
  XOR U488 ( .A(n388), .B(n387), .Z(c[95]) );
  XOR U489 ( .A(a[96]), .B(b[96]), .Z(n392) );
  NAND U490 ( .A(a[95]), .B(b[95]), .Z(n390) );
  NAND U491 ( .A(n388), .B(n387), .Z(n389) );
  NAND U492 ( .A(n390), .B(n389), .Z(n391) );
  XOR U493 ( .A(n392), .B(n391), .Z(c[96]) );
  XOR U494 ( .A(a[97]), .B(b[97]), .Z(n396) );
  NAND U495 ( .A(a[96]), .B(b[96]), .Z(n394) );
  NAND U496 ( .A(n392), .B(n391), .Z(n393) );
  NAND U497 ( .A(n394), .B(n393), .Z(n395) );
  XOR U498 ( .A(n396), .B(n395), .Z(c[97]) );
  XOR U499 ( .A(a[98]), .B(b[98]), .Z(n400) );
  NAND U500 ( .A(a[97]), .B(b[97]), .Z(n398) );
  NAND U501 ( .A(n396), .B(n395), .Z(n397) );
  NAND U502 ( .A(n398), .B(n397), .Z(n399) );
  XOR U503 ( .A(n400), .B(n399), .Z(c[98]) );
  XOR U504 ( .A(a[99]), .B(b[99]), .Z(n404) );
  NAND U505 ( .A(a[98]), .B(b[98]), .Z(n402) );
  NAND U506 ( .A(n400), .B(n399), .Z(n401) );
  NAND U507 ( .A(n402), .B(n401), .Z(n403) );
  XOR U508 ( .A(n404), .B(n403), .Z(c[99]) );
  XOR U509 ( .A(a[100]), .B(b[100]), .Z(n408) );
  NAND U510 ( .A(a[99]), .B(b[99]), .Z(n406) );
  NAND U511 ( .A(n404), .B(n403), .Z(n405) );
  NAND U512 ( .A(n406), .B(n405), .Z(n407) );
  XOR U513 ( .A(n408), .B(n407), .Z(c[100]) );
  XOR U514 ( .A(a[101]), .B(b[101]), .Z(n412) );
  NAND U515 ( .A(a[100]), .B(b[100]), .Z(n410) );
  NAND U516 ( .A(n408), .B(n407), .Z(n409) );
  NAND U517 ( .A(n410), .B(n409), .Z(n411) );
  XOR U518 ( .A(n412), .B(n411), .Z(c[101]) );
  XOR U519 ( .A(a[102]), .B(b[102]), .Z(n416) );
  NAND U520 ( .A(a[101]), .B(b[101]), .Z(n414) );
  NAND U521 ( .A(n412), .B(n411), .Z(n413) );
  NAND U522 ( .A(n414), .B(n413), .Z(n415) );
  XOR U523 ( .A(n416), .B(n415), .Z(c[102]) );
  XOR U524 ( .A(a[103]), .B(b[103]), .Z(n420) );
  NAND U525 ( .A(a[102]), .B(b[102]), .Z(n418) );
  NAND U526 ( .A(n416), .B(n415), .Z(n417) );
  NAND U527 ( .A(n418), .B(n417), .Z(n419) );
  XOR U528 ( .A(n420), .B(n419), .Z(c[103]) );
  XOR U529 ( .A(a[104]), .B(b[104]), .Z(n424) );
  NAND U530 ( .A(a[103]), .B(b[103]), .Z(n422) );
  NAND U531 ( .A(n420), .B(n419), .Z(n421) );
  NAND U532 ( .A(n422), .B(n421), .Z(n423) );
  XOR U533 ( .A(n424), .B(n423), .Z(c[104]) );
  XOR U534 ( .A(a[105]), .B(b[105]), .Z(n428) );
  NAND U535 ( .A(a[104]), .B(b[104]), .Z(n426) );
  NAND U536 ( .A(n424), .B(n423), .Z(n425) );
  NAND U537 ( .A(n426), .B(n425), .Z(n427) );
  XOR U538 ( .A(n428), .B(n427), .Z(c[105]) );
  XOR U539 ( .A(a[106]), .B(b[106]), .Z(n432) );
  NAND U540 ( .A(a[105]), .B(b[105]), .Z(n430) );
  NAND U541 ( .A(n428), .B(n427), .Z(n429) );
  NAND U542 ( .A(n430), .B(n429), .Z(n431) );
  XOR U543 ( .A(n432), .B(n431), .Z(c[106]) );
  XOR U544 ( .A(a[107]), .B(b[107]), .Z(n436) );
  NAND U545 ( .A(a[106]), .B(b[106]), .Z(n434) );
  NAND U546 ( .A(n432), .B(n431), .Z(n433) );
  NAND U547 ( .A(n434), .B(n433), .Z(n435) );
  XOR U548 ( .A(n436), .B(n435), .Z(c[107]) );
  XOR U549 ( .A(a[108]), .B(b[108]), .Z(n440) );
  NAND U550 ( .A(a[107]), .B(b[107]), .Z(n438) );
  NAND U551 ( .A(n436), .B(n435), .Z(n437) );
  NAND U552 ( .A(n438), .B(n437), .Z(n439) );
  XOR U553 ( .A(n440), .B(n439), .Z(c[108]) );
  XOR U554 ( .A(a[109]), .B(b[109]), .Z(n444) );
  NAND U555 ( .A(a[108]), .B(b[108]), .Z(n442) );
  NAND U556 ( .A(n440), .B(n439), .Z(n441) );
  NAND U557 ( .A(n442), .B(n441), .Z(n443) );
  XOR U558 ( .A(n444), .B(n443), .Z(c[109]) );
  NAND U559 ( .A(a[109]), .B(b[109]), .Z(n446) );
  NAND U560 ( .A(n444), .B(n443), .Z(n445) );
  AND U561 ( .A(n446), .B(n445), .Z(n448) );
  XOR U562 ( .A(b[110]), .B(a[110]), .Z(n447) );
  XNOR U563 ( .A(n448), .B(n447), .Z(c[110]) );
  OR U564 ( .A(b[110]), .B(a[110]), .Z(n450) );
  NAND U565 ( .A(n448), .B(n447), .Z(n449) );
  AND U566 ( .A(n450), .B(n449), .Z(n452) );
  XOR U567 ( .A(a[111]), .B(b[111]), .Z(n451) );
  XOR U568 ( .A(n452), .B(n451), .Z(c[111]) );
  XOR U569 ( .A(b[112]), .B(a[112]), .Z(n456) );
  NAND U570 ( .A(a[111]), .B(b[111]), .Z(n454) );
  NAND U571 ( .A(n452), .B(n451), .Z(n453) );
  AND U572 ( .A(n454), .B(n453), .Z(n455) );
  XNOR U573 ( .A(n456), .B(n455), .Z(c[112]) );
  OR U574 ( .A(b[112]), .B(a[112]), .Z(n458) );
  NAND U575 ( .A(n456), .B(n455), .Z(n457) );
  AND U576 ( .A(n458), .B(n457), .Z(n460) );
  XOR U577 ( .A(a[113]), .B(b[113]), .Z(n459) );
  XOR U578 ( .A(n460), .B(n459), .Z(c[113]) );
  XOR U579 ( .A(a[114]), .B(b[114]), .Z(n464) );
  NAND U580 ( .A(a[113]), .B(b[113]), .Z(n462) );
  NAND U581 ( .A(n460), .B(n459), .Z(n461) );
  NAND U582 ( .A(n462), .B(n461), .Z(n463) );
  XOR U583 ( .A(n464), .B(n463), .Z(c[114]) );
  XOR U584 ( .A(a[115]), .B(b[115]), .Z(n468) );
  NAND U585 ( .A(a[114]), .B(b[114]), .Z(n466) );
  NAND U586 ( .A(n464), .B(n463), .Z(n465) );
  NAND U587 ( .A(n466), .B(n465), .Z(n467) );
  XOR U588 ( .A(n468), .B(n467), .Z(c[115]) );
  XOR U589 ( .A(a[116]), .B(b[116]), .Z(n472) );
  NAND U590 ( .A(a[115]), .B(b[115]), .Z(n470) );
  NAND U591 ( .A(n468), .B(n467), .Z(n469) );
  NAND U592 ( .A(n470), .B(n469), .Z(n471) );
  XOR U593 ( .A(n472), .B(n471), .Z(c[116]) );
  XOR U594 ( .A(a[117]), .B(b[117]), .Z(n476) );
  NAND U595 ( .A(a[116]), .B(b[116]), .Z(n474) );
  NAND U596 ( .A(n472), .B(n471), .Z(n473) );
  NAND U597 ( .A(n474), .B(n473), .Z(n475) );
  XOR U598 ( .A(n476), .B(n475), .Z(c[117]) );
  XOR U599 ( .A(a[118]), .B(b[118]), .Z(n480) );
  NAND U600 ( .A(a[117]), .B(b[117]), .Z(n478) );
  NAND U601 ( .A(n476), .B(n475), .Z(n477) );
  NAND U602 ( .A(n478), .B(n477), .Z(n479) );
  XOR U603 ( .A(n480), .B(n479), .Z(c[118]) );
  XOR U604 ( .A(a[119]), .B(b[119]), .Z(n484) );
  NAND U605 ( .A(a[118]), .B(b[118]), .Z(n482) );
  NAND U606 ( .A(n480), .B(n479), .Z(n481) );
  NAND U607 ( .A(n482), .B(n481), .Z(n483) );
  XOR U608 ( .A(n484), .B(n483), .Z(c[119]) );
  XOR U609 ( .A(a[120]), .B(b[120]), .Z(n488) );
  NAND U610 ( .A(a[119]), .B(b[119]), .Z(n486) );
  NAND U611 ( .A(n484), .B(n483), .Z(n485) );
  NAND U612 ( .A(n486), .B(n485), .Z(n487) );
  XOR U613 ( .A(n488), .B(n487), .Z(c[120]) );
  XOR U614 ( .A(a[121]), .B(b[121]), .Z(n492) );
  NAND U615 ( .A(a[120]), .B(b[120]), .Z(n490) );
  NAND U616 ( .A(n488), .B(n487), .Z(n489) );
  NAND U617 ( .A(n490), .B(n489), .Z(n491) );
  XOR U618 ( .A(n492), .B(n491), .Z(c[121]) );
  XOR U619 ( .A(a[122]), .B(b[122]), .Z(n496) );
  NAND U620 ( .A(a[121]), .B(b[121]), .Z(n494) );
  NAND U621 ( .A(n492), .B(n491), .Z(n493) );
  NAND U622 ( .A(n494), .B(n493), .Z(n495) );
  XOR U623 ( .A(n496), .B(n495), .Z(c[122]) );
  XOR U624 ( .A(a[123]), .B(b[123]), .Z(n500) );
  NAND U625 ( .A(a[122]), .B(b[122]), .Z(n498) );
  NAND U626 ( .A(n496), .B(n495), .Z(n497) );
  NAND U627 ( .A(n498), .B(n497), .Z(n499) );
  XOR U628 ( .A(n500), .B(n499), .Z(c[123]) );
  XOR U629 ( .A(a[124]), .B(b[124]), .Z(n504) );
  NAND U630 ( .A(a[123]), .B(b[123]), .Z(n502) );
  NAND U631 ( .A(n500), .B(n499), .Z(n501) );
  NAND U632 ( .A(n502), .B(n501), .Z(n503) );
  XOR U633 ( .A(n504), .B(n503), .Z(c[124]) );
  XOR U634 ( .A(a[125]), .B(b[125]), .Z(n508) );
  NAND U635 ( .A(a[124]), .B(b[124]), .Z(n506) );
  NAND U636 ( .A(n504), .B(n503), .Z(n505) );
  NAND U637 ( .A(n506), .B(n505), .Z(n507) );
  XOR U638 ( .A(n508), .B(n507), .Z(c[125]) );
  XOR U639 ( .A(a[126]), .B(b[126]), .Z(n512) );
  NAND U640 ( .A(a[125]), .B(b[125]), .Z(n510) );
  NAND U641 ( .A(n508), .B(n507), .Z(n509) );
  NAND U642 ( .A(n510), .B(n509), .Z(n511) );
  XOR U643 ( .A(n512), .B(n511), .Z(c[126]) );
  XOR U644 ( .A(a[127]), .B(b[127]), .Z(n516) );
  NAND U645 ( .A(a[126]), .B(b[126]), .Z(n514) );
  NAND U646 ( .A(n512), .B(n511), .Z(n513) );
  NAND U647 ( .A(n514), .B(n513), .Z(n515) );
  XOR U648 ( .A(n516), .B(n515), .Z(c[127]) );
  XOR U649 ( .A(a[128]), .B(b[128]), .Z(n520) );
  NAND U650 ( .A(a[127]), .B(b[127]), .Z(n518) );
  NAND U651 ( .A(n516), .B(n515), .Z(n517) );
  NAND U652 ( .A(n518), .B(n517), .Z(n519) );
  XOR U653 ( .A(n520), .B(n519), .Z(c[128]) );
  XOR U654 ( .A(a[129]), .B(b[129]), .Z(n524) );
  NAND U655 ( .A(a[128]), .B(b[128]), .Z(n522) );
  NAND U656 ( .A(n520), .B(n519), .Z(n521) );
  NAND U657 ( .A(n522), .B(n521), .Z(n523) );
  XOR U658 ( .A(n524), .B(n523), .Z(c[129]) );
  XOR U659 ( .A(a[130]), .B(b[130]), .Z(n528) );
  NAND U660 ( .A(a[129]), .B(b[129]), .Z(n526) );
  NAND U661 ( .A(n524), .B(n523), .Z(n525) );
  NAND U662 ( .A(n526), .B(n525), .Z(n527) );
  XOR U663 ( .A(n528), .B(n527), .Z(c[130]) );
  XOR U664 ( .A(a[131]), .B(b[131]), .Z(n532) );
  NAND U665 ( .A(a[130]), .B(b[130]), .Z(n530) );
  NAND U666 ( .A(n528), .B(n527), .Z(n529) );
  NAND U667 ( .A(n530), .B(n529), .Z(n531) );
  XOR U668 ( .A(n532), .B(n531), .Z(c[131]) );
  XOR U669 ( .A(a[132]), .B(b[132]), .Z(n536) );
  NAND U670 ( .A(a[131]), .B(b[131]), .Z(n534) );
  NAND U671 ( .A(n532), .B(n531), .Z(n533) );
  NAND U672 ( .A(n534), .B(n533), .Z(n535) );
  XOR U673 ( .A(n536), .B(n535), .Z(c[132]) );
  NAND U674 ( .A(a[132]), .B(b[132]), .Z(n538) );
  NAND U675 ( .A(n536), .B(n535), .Z(n537) );
  AND U676 ( .A(n538), .B(n537), .Z(n540) );
  XOR U677 ( .A(b[133]), .B(a[133]), .Z(n539) );
  XNOR U678 ( .A(n540), .B(n539), .Z(c[133]) );
  OR U679 ( .A(b[133]), .B(a[133]), .Z(n542) );
  NAND U680 ( .A(n540), .B(n539), .Z(n541) );
  AND U681 ( .A(n542), .B(n541), .Z(n544) );
  XOR U682 ( .A(a[134]), .B(b[134]), .Z(n543) );
  XOR U683 ( .A(n544), .B(n543), .Z(c[134]) );
  XOR U684 ( .A(a[135]), .B(b[135]), .Z(n548) );
  NAND U685 ( .A(a[134]), .B(b[134]), .Z(n546) );
  NAND U686 ( .A(n544), .B(n543), .Z(n545) );
  NAND U687 ( .A(n546), .B(n545), .Z(n547) );
  XOR U688 ( .A(n548), .B(n547), .Z(c[135]) );
  XOR U689 ( .A(a[136]), .B(b[136]), .Z(n552) );
  NAND U690 ( .A(a[135]), .B(b[135]), .Z(n550) );
  NAND U691 ( .A(n548), .B(n547), .Z(n549) );
  NAND U692 ( .A(n550), .B(n549), .Z(n551) );
  XOR U693 ( .A(n552), .B(n551), .Z(c[136]) );
  XOR U694 ( .A(a[137]), .B(b[137]), .Z(n556) );
  NAND U695 ( .A(a[136]), .B(b[136]), .Z(n554) );
  NAND U696 ( .A(n552), .B(n551), .Z(n553) );
  NAND U697 ( .A(n554), .B(n553), .Z(n555) );
  XOR U698 ( .A(n556), .B(n555), .Z(c[137]) );
  XOR U699 ( .A(a[138]), .B(b[138]), .Z(n560) );
  NAND U700 ( .A(a[137]), .B(b[137]), .Z(n558) );
  NAND U701 ( .A(n556), .B(n555), .Z(n557) );
  NAND U702 ( .A(n558), .B(n557), .Z(n559) );
  XOR U703 ( .A(n560), .B(n559), .Z(c[138]) );
  XOR U704 ( .A(a[139]), .B(b[139]), .Z(n564) );
  NAND U705 ( .A(a[138]), .B(b[138]), .Z(n562) );
  NAND U706 ( .A(n560), .B(n559), .Z(n561) );
  NAND U707 ( .A(n562), .B(n561), .Z(n563) );
  XOR U708 ( .A(n564), .B(n563), .Z(c[139]) );
  XOR U709 ( .A(a[140]), .B(b[140]), .Z(n568) );
  NAND U710 ( .A(a[139]), .B(b[139]), .Z(n566) );
  NAND U711 ( .A(n564), .B(n563), .Z(n565) );
  NAND U712 ( .A(n566), .B(n565), .Z(n567) );
  XOR U713 ( .A(n568), .B(n567), .Z(c[140]) );
  XOR U714 ( .A(a[141]), .B(b[141]), .Z(n572) );
  NAND U715 ( .A(a[140]), .B(b[140]), .Z(n570) );
  NAND U716 ( .A(n568), .B(n567), .Z(n569) );
  NAND U717 ( .A(n570), .B(n569), .Z(n571) );
  XOR U718 ( .A(n572), .B(n571), .Z(c[141]) );
  XOR U719 ( .A(a[142]), .B(b[142]), .Z(n576) );
  NAND U720 ( .A(a[141]), .B(b[141]), .Z(n574) );
  NAND U721 ( .A(n572), .B(n571), .Z(n573) );
  NAND U722 ( .A(n574), .B(n573), .Z(n575) );
  XOR U723 ( .A(n576), .B(n575), .Z(c[142]) );
  XOR U724 ( .A(a[143]), .B(b[143]), .Z(n580) );
  NAND U725 ( .A(a[142]), .B(b[142]), .Z(n578) );
  NAND U726 ( .A(n576), .B(n575), .Z(n577) );
  NAND U727 ( .A(n578), .B(n577), .Z(n579) );
  XOR U728 ( .A(n580), .B(n579), .Z(c[143]) );
  XOR U729 ( .A(a[144]), .B(b[144]), .Z(n584) );
  NAND U730 ( .A(a[143]), .B(b[143]), .Z(n582) );
  NAND U731 ( .A(n580), .B(n579), .Z(n581) );
  NAND U732 ( .A(n582), .B(n581), .Z(n583) );
  XOR U733 ( .A(n584), .B(n583), .Z(c[144]) );
  XOR U734 ( .A(a[145]), .B(b[145]), .Z(n588) );
  NAND U735 ( .A(a[144]), .B(b[144]), .Z(n586) );
  NAND U736 ( .A(n584), .B(n583), .Z(n585) );
  NAND U737 ( .A(n586), .B(n585), .Z(n587) );
  XOR U738 ( .A(n588), .B(n587), .Z(c[145]) );
  XOR U739 ( .A(a[146]), .B(b[146]), .Z(n592) );
  NAND U740 ( .A(a[145]), .B(b[145]), .Z(n590) );
  NAND U741 ( .A(n588), .B(n587), .Z(n589) );
  NAND U742 ( .A(n590), .B(n589), .Z(n591) );
  XOR U743 ( .A(n592), .B(n591), .Z(c[146]) );
  XOR U744 ( .A(a[147]), .B(b[147]), .Z(n596) );
  NAND U745 ( .A(a[146]), .B(b[146]), .Z(n594) );
  NAND U746 ( .A(n592), .B(n591), .Z(n593) );
  NAND U747 ( .A(n594), .B(n593), .Z(n595) );
  XOR U748 ( .A(n596), .B(n595), .Z(c[147]) );
  XOR U749 ( .A(a[148]), .B(b[148]), .Z(n600) );
  NAND U750 ( .A(a[147]), .B(b[147]), .Z(n598) );
  NAND U751 ( .A(n596), .B(n595), .Z(n597) );
  NAND U752 ( .A(n598), .B(n597), .Z(n599) );
  XOR U753 ( .A(n600), .B(n599), .Z(c[148]) );
  XOR U754 ( .A(a[149]), .B(b[149]), .Z(n604) );
  NAND U755 ( .A(a[148]), .B(b[148]), .Z(n602) );
  NAND U756 ( .A(n600), .B(n599), .Z(n601) );
  NAND U757 ( .A(n602), .B(n601), .Z(n603) );
  XOR U758 ( .A(n604), .B(n603), .Z(c[149]) );
  XOR U759 ( .A(a[150]), .B(b[150]), .Z(n608) );
  NAND U760 ( .A(a[149]), .B(b[149]), .Z(n606) );
  NAND U761 ( .A(n604), .B(n603), .Z(n605) );
  NAND U762 ( .A(n606), .B(n605), .Z(n607) );
  XOR U763 ( .A(n608), .B(n607), .Z(c[150]) );
  XOR U764 ( .A(a[151]), .B(b[151]), .Z(n612) );
  NAND U765 ( .A(a[150]), .B(b[150]), .Z(n610) );
  NAND U766 ( .A(n608), .B(n607), .Z(n609) );
  NAND U767 ( .A(n610), .B(n609), .Z(n611) );
  XOR U768 ( .A(n612), .B(n611), .Z(c[151]) );
  XOR U769 ( .A(a[152]), .B(b[152]), .Z(n616) );
  NAND U770 ( .A(a[151]), .B(b[151]), .Z(n614) );
  NAND U771 ( .A(n612), .B(n611), .Z(n613) );
  NAND U772 ( .A(n614), .B(n613), .Z(n615) );
  XOR U773 ( .A(n616), .B(n615), .Z(c[152]) );
  NAND U774 ( .A(a[152]), .B(b[152]), .Z(n618) );
  NAND U775 ( .A(n616), .B(n615), .Z(n617) );
  AND U776 ( .A(n618), .B(n617), .Z(n620) );
  XOR U777 ( .A(b[153]), .B(a[153]), .Z(n619) );
  XNOR U778 ( .A(n620), .B(n619), .Z(c[153]) );
  OR U779 ( .A(b[153]), .B(a[153]), .Z(n622) );
  NAND U780 ( .A(n620), .B(n619), .Z(n621) );
  AND U781 ( .A(n622), .B(n621), .Z(n624) );
  XOR U782 ( .A(a[154]), .B(b[154]), .Z(n623) );
  XOR U783 ( .A(n624), .B(n623), .Z(c[154]) );
  XOR U784 ( .A(a[155]), .B(b[155]), .Z(n628) );
  NAND U785 ( .A(a[154]), .B(b[154]), .Z(n626) );
  NAND U786 ( .A(n624), .B(n623), .Z(n625) );
  NAND U787 ( .A(n626), .B(n625), .Z(n627) );
  XOR U788 ( .A(n628), .B(n627), .Z(c[155]) );
  XOR U789 ( .A(a[156]), .B(b[156]), .Z(n632) );
  NAND U790 ( .A(a[155]), .B(b[155]), .Z(n630) );
  NAND U791 ( .A(n628), .B(n627), .Z(n629) );
  NAND U792 ( .A(n630), .B(n629), .Z(n631) );
  XOR U793 ( .A(n632), .B(n631), .Z(c[156]) );
  XOR U794 ( .A(a[157]), .B(b[157]), .Z(n636) );
  NAND U795 ( .A(a[156]), .B(b[156]), .Z(n634) );
  NAND U796 ( .A(n632), .B(n631), .Z(n633) );
  NAND U797 ( .A(n634), .B(n633), .Z(n635) );
  XOR U798 ( .A(n636), .B(n635), .Z(c[157]) );
  XOR U799 ( .A(a[158]), .B(b[158]), .Z(n640) );
  NAND U800 ( .A(a[157]), .B(b[157]), .Z(n638) );
  NAND U801 ( .A(n636), .B(n635), .Z(n637) );
  NAND U802 ( .A(n638), .B(n637), .Z(n639) );
  XOR U803 ( .A(n640), .B(n639), .Z(c[158]) );
  XOR U804 ( .A(a[159]), .B(b[159]), .Z(n644) );
  NAND U805 ( .A(a[158]), .B(b[158]), .Z(n642) );
  NAND U806 ( .A(n640), .B(n639), .Z(n641) );
  NAND U807 ( .A(n642), .B(n641), .Z(n643) );
  XOR U808 ( .A(n644), .B(n643), .Z(c[159]) );
  XOR U809 ( .A(a[160]), .B(b[160]), .Z(n648) );
  NAND U810 ( .A(a[159]), .B(b[159]), .Z(n646) );
  NAND U811 ( .A(n644), .B(n643), .Z(n645) );
  NAND U812 ( .A(n646), .B(n645), .Z(n647) );
  XOR U813 ( .A(n648), .B(n647), .Z(c[160]) );
  XOR U814 ( .A(a[161]), .B(b[161]), .Z(n652) );
  NAND U815 ( .A(a[160]), .B(b[160]), .Z(n650) );
  NAND U816 ( .A(n648), .B(n647), .Z(n649) );
  NAND U817 ( .A(n650), .B(n649), .Z(n651) );
  XOR U818 ( .A(n652), .B(n651), .Z(c[161]) );
  XOR U819 ( .A(a[162]), .B(b[162]), .Z(n656) );
  NAND U820 ( .A(a[161]), .B(b[161]), .Z(n654) );
  NAND U821 ( .A(n652), .B(n651), .Z(n653) );
  NAND U822 ( .A(n654), .B(n653), .Z(n655) );
  XOR U823 ( .A(n656), .B(n655), .Z(c[162]) );
  XOR U824 ( .A(a[163]), .B(b[163]), .Z(n660) );
  NAND U825 ( .A(a[162]), .B(b[162]), .Z(n658) );
  NAND U826 ( .A(n656), .B(n655), .Z(n657) );
  NAND U827 ( .A(n658), .B(n657), .Z(n659) );
  XOR U828 ( .A(n660), .B(n659), .Z(c[163]) );
  XOR U829 ( .A(a[164]), .B(b[164]), .Z(n664) );
  NAND U830 ( .A(a[163]), .B(b[163]), .Z(n662) );
  NAND U831 ( .A(n660), .B(n659), .Z(n661) );
  NAND U832 ( .A(n662), .B(n661), .Z(n663) );
  XOR U833 ( .A(n664), .B(n663), .Z(c[164]) );
  XOR U834 ( .A(a[165]), .B(b[165]), .Z(n668) );
  NAND U835 ( .A(a[164]), .B(b[164]), .Z(n666) );
  NAND U836 ( .A(n664), .B(n663), .Z(n665) );
  NAND U837 ( .A(n666), .B(n665), .Z(n667) );
  XOR U838 ( .A(n668), .B(n667), .Z(c[165]) );
  XOR U839 ( .A(a[166]), .B(b[166]), .Z(n672) );
  NAND U840 ( .A(a[165]), .B(b[165]), .Z(n670) );
  NAND U841 ( .A(n668), .B(n667), .Z(n669) );
  NAND U842 ( .A(n670), .B(n669), .Z(n671) );
  XOR U843 ( .A(n672), .B(n671), .Z(c[166]) );
  XOR U844 ( .A(a[167]), .B(b[167]), .Z(n676) );
  NAND U845 ( .A(a[166]), .B(b[166]), .Z(n674) );
  NAND U846 ( .A(n672), .B(n671), .Z(n673) );
  NAND U847 ( .A(n674), .B(n673), .Z(n675) );
  XOR U848 ( .A(n676), .B(n675), .Z(c[167]) );
  XOR U849 ( .A(a[168]), .B(b[168]), .Z(n680) );
  NAND U850 ( .A(a[167]), .B(b[167]), .Z(n678) );
  NAND U851 ( .A(n676), .B(n675), .Z(n677) );
  NAND U852 ( .A(n678), .B(n677), .Z(n679) );
  XOR U853 ( .A(n680), .B(n679), .Z(c[168]) );
  XOR U854 ( .A(a[169]), .B(b[169]), .Z(n684) );
  NAND U855 ( .A(a[168]), .B(b[168]), .Z(n682) );
  NAND U856 ( .A(n680), .B(n679), .Z(n681) );
  NAND U857 ( .A(n682), .B(n681), .Z(n683) );
  XOR U858 ( .A(n684), .B(n683), .Z(c[169]) );
  XOR U859 ( .A(a[170]), .B(b[170]), .Z(n688) );
  NAND U860 ( .A(a[169]), .B(b[169]), .Z(n686) );
  NAND U861 ( .A(n684), .B(n683), .Z(n685) );
  NAND U862 ( .A(n686), .B(n685), .Z(n687) );
  XOR U863 ( .A(n688), .B(n687), .Z(c[170]) );
  XOR U864 ( .A(a[171]), .B(b[171]), .Z(n692) );
  NAND U865 ( .A(a[170]), .B(b[170]), .Z(n690) );
  NAND U866 ( .A(n688), .B(n687), .Z(n689) );
  NAND U867 ( .A(n690), .B(n689), .Z(n691) );
  XOR U868 ( .A(n692), .B(n691), .Z(c[171]) );
  XOR U869 ( .A(a[172]), .B(b[172]), .Z(n696) );
  NAND U870 ( .A(a[171]), .B(b[171]), .Z(n694) );
  NAND U871 ( .A(n692), .B(n691), .Z(n693) );
  NAND U872 ( .A(n694), .B(n693), .Z(n695) );
  XOR U873 ( .A(n696), .B(n695), .Z(c[172]) );
  XOR U874 ( .A(a[173]), .B(b[173]), .Z(n700) );
  NAND U875 ( .A(a[172]), .B(b[172]), .Z(n698) );
  NAND U876 ( .A(n696), .B(n695), .Z(n697) );
  NAND U877 ( .A(n698), .B(n697), .Z(n699) );
  XOR U878 ( .A(n700), .B(n699), .Z(c[173]) );
  XOR U879 ( .A(a[174]), .B(b[174]), .Z(n704) );
  NAND U880 ( .A(a[173]), .B(b[173]), .Z(n702) );
  NAND U881 ( .A(n700), .B(n699), .Z(n701) );
  NAND U882 ( .A(n702), .B(n701), .Z(n703) );
  XOR U883 ( .A(n704), .B(n703), .Z(c[174]) );
  XOR U884 ( .A(a[175]), .B(b[175]), .Z(n708) );
  NAND U885 ( .A(a[174]), .B(b[174]), .Z(n706) );
  NAND U886 ( .A(n704), .B(n703), .Z(n705) );
  NAND U887 ( .A(n706), .B(n705), .Z(n707) );
  XOR U888 ( .A(n708), .B(n707), .Z(c[175]) );
  XOR U889 ( .A(a[176]), .B(b[176]), .Z(n712) );
  NAND U890 ( .A(a[175]), .B(b[175]), .Z(n710) );
  NAND U891 ( .A(n708), .B(n707), .Z(n709) );
  NAND U892 ( .A(n710), .B(n709), .Z(n711) );
  XOR U893 ( .A(n712), .B(n711), .Z(c[176]) );
  XOR U894 ( .A(a[177]), .B(b[177]), .Z(n716) );
  NAND U895 ( .A(a[176]), .B(b[176]), .Z(n714) );
  NAND U896 ( .A(n712), .B(n711), .Z(n713) );
  NAND U897 ( .A(n714), .B(n713), .Z(n715) );
  XOR U898 ( .A(n716), .B(n715), .Z(c[177]) );
  XOR U899 ( .A(a[178]), .B(b[178]), .Z(n720) );
  NAND U900 ( .A(a[177]), .B(b[177]), .Z(n718) );
  NAND U901 ( .A(n716), .B(n715), .Z(n717) );
  NAND U902 ( .A(n718), .B(n717), .Z(n719) );
  XOR U903 ( .A(n720), .B(n719), .Z(c[178]) );
  XOR U904 ( .A(a[179]), .B(b[179]), .Z(n724) );
  NAND U905 ( .A(a[178]), .B(b[178]), .Z(n722) );
  NAND U906 ( .A(n720), .B(n719), .Z(n721) );
  NAND U907 ( .A(n722), .B(n721), .Z(n723) );
  XOR U908 ( .A(n724), .B(n723), .Z(c[179]) );
  XOR U909 ( .A(a[180]), .B(b[180]), .Z(n728) );
  NAND U910 ( .A(a[179]), .B(b[179]), .Z(n726) );
  NAND U911 ( .A(n724), .B(n723), .Z(n725) );
  NAND U912 ( .A(n726), .B(n725), .Z(n727) );
  XOR U913 ( .A(n728), .B(n727), .Z(c[180]) );
  XOR U914 ( .A(a[181]), .B(b[181]), .Z(n732) );
  NAND U915 ( .A(a[180]), .B(b[180]), .Z(n730) );
  NAND U916 ( .A(n728), .B(n727), .Z(n729) );
  NAND U917 ( .A(n730), .B(n729), .Z(n731) );
  XOR U918 ( .A(n732), .B(n731), .Z(c[181]) );
  XOR U919 ( .A(a[182]), .B(b[182]), .Z(n736) );
  NAND U920 ( .A(a[181]), .B(b[181]), .Z(n734) );
  NAND U921 ( .A(n732), .B(n731), .Z(n733) );
  NAND U922 ( .A(n734), .B(n733), .Z(n735) );
  XOR U923 ( .A(n736), .B(n735), .Z(c[182]) );
  XOR U924 ( .A(a[183]), .B(b[183]), .Z(n740) );
  NAND U925 ( .A(a[182]), .B(b[182]), .Z(n738) );
  NAND U926 ( .A(n736), .B(n735), .Z(n737) );
  NAND U927 ( .A(n738), .B(n737), .Z(n739) );
  XOR U928 ( .A(n740), .B(n739), .Z(c[183]) );
  XOR U929 ( .A(a[184]), .B(b[184]), .Z(n744) );
  NAND U930 ( .A(a[183]), .B(b[183]), .Z(n742) );
  NAND U931 ( .A(n740), .B(n739), .Z(n741) );
  NAND U932 ( .A(n742), .B(n741), .Z(n743) );
  XOR U933 ( .A(n744), .B(n743), .Z(c[184]) );
  XOR U934 ( .A(a[185]), .B(b[185]), .Z(n748) );
  NAND U935 ( .A(a[184]), .B(b[184]), .Z(n746) );
  NAND U936 ( .A(n744), .B(n743), .Z(n745) );
  NAND U937 ( .A(n746), .B(n745), .Z(n747) );
  XOR U938 ( .A(n748), .B(n747), .Z(c[185]) );
  XOR U939 ( .A(a[186]), .B(b[186]), .Z(n752) );
  NAND U940 ( .A(a[185]), .B(b[185]), .Z(n750) );
  NAND U941 ( .A(n748), .B(n747), .Z(n749) );
  NAND U942 ( .A(n750), .B(n749), .Z(n751) );
  XOR U943 ( .A(n752), .B(n751), .Z(c[186]) );
  XOR U944 ( .A(b[187]), .B(a[187]), .Z(n756) );
  NAND U945 ( .A(a[186]), .B(b[186]), .Z(n754) );
  NAND U946 ( .A(n752), .B(n751), .Z(n753) );
  AND U947 ( .A(n754), .B(n753), .Z(n755) );
  XNOR U948 ( .A(n756), .B(n755), .Z(c[187]) );
  OR U949 ( .A(b[187]), .B(a[187]), .Z(n758) );
  NAND U950 ( .A(n756), .B(n755), .Z(n757) );
  AND U951 ( .A(n758), .B(n757), .Z(n760) );
  XOR U952 ( .A(a[188]), .B(b[188]), .Z(n759) );
  XOR U953 ( .A(n760), .B(n759), .Z(c[188]) );
  XOR U954 ( .A(a[189]), .B(b[189]), .Z(n764) );
  NAND U955 ( .A(a[188]), .B(b[188]), .Z(n762) );
  NAND U956 ( .A(n760), .B(n759), .Z(n761) );
  NAND U957 ( .A(n762), .B(n761), .Z(n763) );
  XOR U958 ( .A(n764), .B(n763), .Z(c[189]) );
  XOR U959 ( .A(a[190]), .B(b[190]), .Z(n768) );
  NAND U960 ( .A(a[189]), .B(b[189]), .Z(n766) );
  NAND U961 ( .A(n764), .B(n763), .Z(n765) );
  NAND U962 ( .A(n766), .B(n765), .Z(n767) );
  XOR U963 ( .A(n768), .B(n767), .Z(c[190]) );
  XOR U964 ( .A(a[191]), .B(b[191]), .Z(n772) );
  NAND U965 ( .A(a[190]), .B(b[190]), .Z(n770) );
  NAND U966 ( .A(n768), .B(n767), .Z(n769) );
  NAND U967 ( .A(n770), .B(n769), .Z(n771) );
  XOR U968 ( .A(n772), .B(n771), .Z(c[191]) );
  XOR U969 ( .A(b[192]), .B(a[192]), .Z(n776) );
  NAND U970 ( .A(a[191]), .B(b[191]), .Z(n774) );
  NAND U971 ( .A(n772), .B(n771), .Z(n773) );
  AND U972 ( .A(n774), .B(n773), .Z(n775) );
  XNOR U973 ( .A(n776), .B(n775), .Z(c[192]) );
  OR U974 ( .A(b[192]), .B(a[192]), .Z(n778) );
  NAND U975 ( .A(n776), .B(n775), .Z(n777) );
  AND U976 ( .A(n778), .B(n777), .Z(n780) );
  XOR U977 ( .A(a[193]), .B(b[193]), .Z(n779) );
  XOR U978 ( .A(n780), .B(n779), .Z(c[193]) );
  XOR U979 ( .A(a[194]), .B(b[194]), .Z(n784) );
  NAND U980 ( .A(a[193]), .B(b[193]), .Z(n782) );
  NAND U981 ( .A(n780), .B(n779), .Z(n781) );
  NAND U982 ( .A(n782), .B(n781), .Z(n783) );
  XOR U983 ( .A(n784), .B(n783), .Z(c[194]) );
  XOR U984 ( .A(a[195]), .B(b[195]), .Z(n788) );
  NAND U985 ( .A(a[194]), .B(b[194]), .Z(n786) );
  NAND U986 ( .A(n784), .B(n783), .Z(n785) );
  NAND U987 ( .A(n786), .B(n785), .Z(n787) );
  XOR U988 ( .A(n788), .B(n787), .Z(c[195]) );
  XOR U989 ( .A(a[196]), .B(b[196]), .Z(n792) );
  NAND U990 ( .A(a[195]), .B(b[195]), .Z(n790) );
  NAND U991 ( .A(n788), .B(n787), .Z(n789) );
  NAND U992 ( .A(n790), .B(n789), .Z(n791) );
  XOR U993 ( .A(n792), .B(n791), .Z(c[196]) );
  XOR U994 ( .A(a[197]), .B(b[197]), .Z(n796) );
  NAND U995 ( .A(a[196]), .B(b[196]), .Z(n794) );
  NAND U996 ( .A(n792), .B(n791), .Z(n793) );
  NAND U997 ( .A(n794), .B(n793), .Z(n795) );
  XOR U998 ( .A(n796), .B(n795), .Z(c[197]) );
  XOR U999 ( .A(a[198]), .B(b[198]), .Z(n800) );
  NAND U1000 ( .A(a[197]), .B(b[197]), .Z(n798) );
  NAND U1001 ( .A(n796), .B(n795), .Z(n797) );
  NAND U1002 ( .A(n798), .B(n797), .Z(n799) );
  XOR U1003 ( .A(n800), .B(n799), .Z(c[198]) );
  XOR U1004 ( .A(a[199]), .B(b[199]), .Z(n804) );
  NAND U1005 ( .A(a[198]), .B(b[198]), .Z(n802) );
  NAND U1006 ( .A(n800), .B(n799), .Z(n801) );
  NAND U1007 ( .A(n802), .B(n801), .Z(n803) );
  XOR U1008 ( .A(n804), .B(n803), .Z(c[199]) );
  XOR U1009 ( .A(a[200]), .B(b[200]), .Z(n808) );
  NAND U1010 ( .A(a[199]), .B(b[199]), .Z(n806) );
  NAND U1011 ( .A(n804), .B(n803), .Z(n805) );
  NAND U1012 ( .A(n806), .B(n805), .Z(n807) );
  XOR U1013 ( .A(n808), .B(n807), .Z(c[200]) );
  XOR U1014 ( .A(a[201]), .B(b[201]), .Z(n812) );
  NAND U1015 ( .A(a[200]), .B(b[200]), .Z(n810) );
  NAND U1016 ( .A(n808), .B(n807), .Z(n809) );
  NAND U1017 ( .A(n810), .B(n809), .Z(n811) );
  XOR U1018 ( .A(n812), .B(n811), .Z(c[201]) );
  XOR U1019 ( .A(a[202]), .B(b[202]), .Z(n816) );
  NAND U1020 ( .A(a[201]), .B(b[201]), .Z(n814) );
  NAND U1021 ( .A(n812), .B(n811), .Z(n813) );
  NAND U1022 ( .A(n814), .B(n813), .Z(n815) );
  XOR U1023 ( .A(n816), .B(n815), .Z(c[202]) );
  XOR U1024 ( .A(b[203]), .B(a[203]), .Z(n820) );
  NAND U1025 ( .A(a[202]), .B(b[202]), .Z(n818) );
  NAND U1026 ( .A(n816), .B(n815), .Z(n817) );
  AND U1027 ( .A(n818), .B(n817), .Z(n819) );
  XNOR U1028 ( .A(n820), .B(n819), .Z(c[203]) );
  XOR U1029 ( .A(b[204]), .B(a[204]), .Z(n824) );
  OR U1030 ( .A(b[203]), .B(a[203]), .Z(n822) );
  NAND U1031 ( .A(n820), .B(n819), .Z(n821) );
  NAND U1032 ( .A(n822), .B(n821), .Z(n823) );
  XNOR U1033 ( .A(n824), .B(n823), .Z(c[204]) );
  XOR U1034 ( .A(a[205]), .B(b[205]), .Z(n828) );
  OR U1035 ( .A(b[204]), .B(a[204]), .Z(n826) );
  NAND U1036 ( .A(n824), .B(n823), .Z(n825) );
  AND U1037 ( .A(n826), .B(n825), .Z(n827) );
  XOR U1038 ( .A(n828), .B(n827), .Z(c[205]) );
  NAND U1039 ( .A(a[205]), .B(b[205]), .Z(n830) );
  NAND U1040 ( .A(n828), .B(n827), .Z(n829) );
  AND U1041 ( .A(n830), .B(n829), .Z(n832) );
  XOR U1042 ( .A(b[206]), .B(a[206]), .Z(n831) );
  XNOR U1043 ( .A(n832), .B(n831), .Z(c[206]) );
  OR U1044 ( .A(b[206]), .B(a[206]), .Z(n834) );
  NAND U1045 ( .A(n832), .B(n831), .Z(n833) );
  AND U1046 ( .A(n834), .B(n833), .Z(n836) );
  XOR U1047 ( .A(a[207]), .B(b[207]), .Z(n835) );
  XOR U1048 ( .A(n836), .B(n835), .Z(c[207]) );
  XOR U1049 ( .A(a[208]), .B(b[208]), .Z(n840) );
  NAND U1050 ( .A(a[207]), .B(b[207]), .Z(n838) );
  NAND U1051 ( .A(n836), .B(n835), .Z(n837) );
  NAND U1052 ( .A(n838), .B(n837), .Z(n839) );
  XOR U1053 ( .A(n840), .B(n839), .Z(c[208]) );
  XOR U1054 ( .A(a[209]), .B(b[209]), .Z(n844) );
  NAND U1055 ( .A(a[208]), .B(b[208]), .Z(n842) );
  NAND U1056 ( .A(n840), .B(n839), .Z(n841) );
  NAND U1057 ( .A(n842), .B(n841), .Z(n843) );
  XOR U1058 ( .A(n844), .B(n843), .Z(c[209]) );
  XOR U1059 ( .A(a[210]), .B(b[210]), .Z(n848) );
  NAND U1060 ( .A(a[209]), .B(b[209]), .Z(n846) );
  NAND U1061 ( .A(n844), .B(n843), .Z(n845) );
  NAND U1062 ( .A(n846), .B(n845), .Z(n847) );
  XOR U1063 ( .A(n848), .B(n847), .Z(c[210]) );
  XOR U1064 ( .A(a[211]), .B(b[211]), .Z(n852) );
  NAND U1065 ( .A(a[210]), .B(b[210]), .Z(n850) );
  NAND U1066 ( .A(n848), .B(n847), .Z(n849) );
  NAND U1067 ( .A(n850), .B(n849), .Z(n851) );
  XOR U1068 ( .A(n852), .B(n851), .Z(c[211]) );
  XOR U1069 ( .A(a[212]), .B(b[212]), .Z(n856) );
  NAND U1070 ( .A(a[211]), .B(b[211]), .Z(n854) );
  NAND U1071 ( .A(n852), .B(n851), .Z(n853) );
  NAND U1072 ( .A(n854), .B(n853), .Z(n855) );
  XOR U1073 ( .A(n856), .B(n855), .Z(c[212]) );
  XOR U1074 ( .A(a[213]), .B(b[213]), .Z(n860) );
  NAND U1075 ( .A(a[212]), .B(b[212]), .Z(n858) );
  NAND U1076 ( .A(n856), .B(n855), .Z(n857) );
  NAND U1077 ( .A(n858), .B(n857), .Z(n859) );
  XOR U1078 ( .A(n860), .B(n859), .Z(c[213]) );
  XOR U1079 ( .A(a[214]), .B(b[214]), .Z(n864) );
  NAND U1080 ( .A(a[213]), .B(b[213]), .Z(n862) );
  NAND U1081 ( .A(n860), .B(n859), .Z(n861) );
  NAND U1082 ( .A(n862), .B(n861), .Z(n863) );
  XOR U1083 ( .A(n864), .B(n863), .Z(c[214]) );
  XOR U1084 ( .A(a[215]), .B(b[215]), .Z(n868) );
  NAND U1085 ( .A(a[214]), .B(b[214]), .Z(n866) );
  NAND U1086 ( .A(n864), .B(n863), .Z(n865) );
  NAND U1087 ( .A(n866), .B(n865), .Z(n867) );
  XOR U1088 ( .A(n868), .B(n867), .Z(c[215]) );
  XOR U1089 ( .A(a[216]), .B(b[216]), .Z(n872) );
  NAND U1090 ( .A(a[215]), .B(b[215]), .Z(n870) );
  NAND U1091 ( .A(n868), .B(n867), .Z(n869) );
  NAND U1092 ( .A(n870), .B(n869), .Z(n871) );
  XOR U1093 ( .A(n872), .B(n871), .Z(c[216]) );
  XOR U1094 ( .A(a[217]), .B(b[217]), .Z(n876) );
  NAND U1095 ( .A(a[216]), .B(b[216]), .Z(n874) );
  NAND U1096 ( .A(n872), .B(n871), .Z(n873) );
  NAND U1097 ( .A(n874), .B(n873), .Z(n875) );
  XOR U1098 ( .A(n876), .B(n875), .Z(c[217]) );
  XOR U1099 ( .A(a[218]), .B(b[218]), .Z(n880) );
  NAND U1100 ( .A(a[217]), .B(b[217]), .Z(n878) );
  NAND U1101 ( .A(n876), .B(n875), .Z(n877) );
  NAND U1102 ( .A(n878), .B(n877), .Z(n879) );
  XOR U1103 ( .A(n880), .B(n879), .Z(c[218]) );
  XOR U1104 ( .A(a[219]), .B(b[219]), .Z(n884) );
  NAND U1105 ( .A(a[218]), .B(b[218]), .Z(n882) );
  NAND U1106 ( .A(n880), .B(n879), .Z(n881) );
  NAND U1107 ( .A(n882), .B(n881), .Z(n883) );
  XOR U1108 ( .A(n884), .B(n883), .Z(c[219]) );
  XOR U1109 ( .A(a[220]), .B(b[220]), .Z(n888) );
  NAND U1110 ( .A(a[219]), .B(b[219]), .Z(n886) );
  NAND U1111 ( .A(n884), .B(n883), .Z(n885) );
  NAND U1112 ( .A(n886), .B(n885), .Z(n887) );
  XOR U1113 ( .A(n888), .B(n887), .Z(c[220]) );
  XOR U1114 ( .A(a[221]), .B(b[221]), .Z(n892) );
  NAND U1115 ( .A(a[220]), .B(b[220]), .Z(n890) );
  NAND U1116 ( .A(n888), .B(n887), .Z(n889) );
  NAND U1117 ( .A(n890), .B(n889), .Z(n891) );
  XOR U1118 ( .A(n892), .B(n891), .Z(c[221]) );
  XOR U1119 ( .A(a[222]), .B(b[222]), .Z(n896) );
  NAND U1120 ( .A(a[221]), .B(b[221]), .Z(n894) );
  NAND U1121 ( .A(n892), .B(n891), .Z(n893) );
  NAND U1122 ( .A(n894), .B(n893), .Z(n895) );
  XOR U1123 ( .A(n896), .B(n895), .Z(c[222]) );
  XOR U1124 ( .A(a[223]), .B(b[223]), .Z(n900) );
  NAND U1125 ( .A(a[222]), .B(b[222]), .Z(n898) );
  NAND U1126 ( .A(n896), .B(n895), .Z(n897) );
  NAND U1127 ( .A(n898), .B(n897), .Z(n899) );
  XOR U1128 ( .A(n900), .B(n899), .Z(c[223]) );
  XOR U1129 ( .A(a[224]), .B(b[224]), .Z(n904) );
  NAND U1130 ( .A(a[223]), .B(b[223]), .Z(n902) );
  NAND U1131 ( .A(n900), .B(n899), .Z(n901) );
  NAND U1132 ( .A(n902), .B(n901), .Z(n903) );
  XOR U1133 ( .A(n904), .B(n903), .Z(c[224]) );
  XOR U1134 ( .A(a[225]), .B(b[225]), .Z(n908) );
  NAND U1135 ( .A(a[224]), .B(b[224]), .Z(n906) );
  NAND U1136 ( .A(n904), .B(n903), .Z(n905) );
  NAND U1137 ( .A(n906), .B(n905), .Z(n907) );
  XOR U1138 ( .A(n908), .B(n907), .Z(c[225]) );
  XOR U1139 ( .A(a[226]), .B(b[226]), .Z(n912) );
  NAND U1140 ( .A(a[225]), .B(b[225]), .Z(n910) );
  NAND U1141 ( .A(n908), .B(n907), .Z(n909) );
  NAND U1142 ( .A(n910), .B(n909), .Z(n911) );
  XOR U1143 ( .A(n912), .B(n911), .Z(c[226]) );
  XOR U1144 ( .A(a[227]), .B(b[227]), .Z(n916) );
  NAND U1145 ( .A(a[226]), .B(b[226]), .Z(n914) );
  NAND U1146 ( .A(n912), .B(n911), .Z(n913) );
  NAND U1147 ( .A(n914), .B(n913), .Z(n915) );
  XOR U1148 ( .A(n916), .B(n915), .Z(c[227]) );
  XOR U1149 ( .A(a[228]), .B(b[228]), .Z(n920) );
  NAND U1150 ( .A(a[227]), .B(b[227]), .Z(n918) );
  NAND U1151 ( .A(n916), .B(n915), .Z(n917) );
  NAND U1152 ( .A(n918), .B(n917), .Z(n919) );
  XOR U1153 ( .A(n920), .B(n919), .Z(c[228]) );
  XOR U1154 ( .A(a[229]), .B(b[229]), .Z(n924) );
  NAND U1155 ( .A(a[228]), .B(b[228]), .Z(n922) );
  NAND U1156 ( .A(n920), .B(n919), .Z(n921) );
  NAND U1157 ( .A(n922), .B(n921), .Z(n923) );
  XOR U1158 ( .A(n924), .B(n923), .Z(c[229]) );
  XOR U1159 ( .A(a[230]), .B(b[230]), .Z(n928) );
  NAND U1160 ( .A(a[229]), .B(b[229]), .Z(n926) );
  NAND U1161 ( .A(n924), .B(n923), .Z(n925) );
  NAND U1162 ( .A(n926), .B(n925), .Z(n927) );
  XOR U1163 ( .A(n928), .B(n927), .Z(c[230]) );
  XOR U1164 ( .A(a[231]), .B(b[231]), .Z(n932) );
  NAND U1165 ( .A(a[230]), .B(b[230]), .Z(n930) );
  NAND U1166 ( .A(n928), .B(n927), .Z(n929) );
  NAND U1167 ( .A(n930), .B(n929), .Z(n931) );
  XOR U1168 ( .A(n932), .B(n931), .Z(c[231]) );
  XOR U1169 ( .A(a[232]), .B(b[232]), .Z(n936) );
  NAND U1170 ( .A(a[231]), .B(b[231]), .Z(n934) );
  NAND U1171 ( .A(n932), .B(n931), .Z(n933) );
  NAND U1172 ( .A(n934), .B(n933), .Z(n935) );
  XOR U1173 ( .A(n936), .B(n935), .Z(c[232]) );
  XOR U1174 ( .A(a[233]), .B(b[233]), .Z(n940) );
  NAND U1175 ( .A(a[232]), .B(b[232]), .Z(n938) );
  NAND U1176 ( .A(n936), .B(n935), .Z(n937) );
  NAND U1177 ( .A(n938), .B(n937), .Z(n939) );
  XOR U1178 ( .A(n940), .B(n939), .Z(c[233]) );
  XOR U1179 ( .A(a[234]), .B(b[234]), .Z(n944) );
  NAND U1180 ( .A(a[233]), .B(b[233]), .Z(n942) );
  NAND U1181 ( .A(n940), .B(n939), .Z(n941) );
  NAND U1182 ( .A(n942), .B(n941), .Z(n943) );
  XOR U1183 ( .A(n944), .B(n943), .Z(c[234]) );
  XOR U1184 ( .A(a[235]), .B(b[235]), .Z(n948) );
  NAND U1185 ( .A(a[234]), .B(b[234]), .Z(n946) );
  NAND U1186 ( .A(n944), .B(n943), .Z(n945) );
  NAND U1187 ( .A(n946), .B(n945), .Z(n947) );
  XOR U1188 ( .A(n948), .B(n947), .Z(c[235]) );
  XOR U1189 ( .A(a[236]), .B(b[236]), .Z(n952) );
  NAND U1190 ( .A(a[235]), .B(b[235]), .Z(n950) );
  NAND U1191 ( .A(n948), .B(n947), .Z(n949) );
  NAND U1192 ( .A(n950), .B(n949), .Z(n951) );
  XOR U1193 ( .A(n952), .B(n951), .Z(c[236]) );
  XOR U1194 ( .A(a[237]), .B(b[237]), .Z(n956) );
  NAND U1195 ( .A(a[236]), .B(b[236]), .Z(n954) );
  NAND U1196 ( .A(n952), .B(n951), .Z(n953) );
  NAND U1197 ( .A(n954), .B(n953), .Z(n955) );
  XOR U1198 ( .A(n956), .B(n955), .Z(c[237]) );
  XOR U1199 ( .A(a[238]), .B(b[238]), .Z(n960) );
  NAND U1200 ( .A(a[237]), .B(b[237]), .Z(n958) );
  NAND U1201 ( .A(n956), .B(n955), .Z(n957) );
  NAND U1202 ( .A(n958), .B(n957), .Z(n959) );
  XOR U1203 ( .A(n960), .B(n959), .Z(c[238]) );
  XOR U1204 ( .A(a[239]), .B(b[239]), .Z(n964) );
  NAND U1205 ( .A(a[238]), .B(b[238]), .Z(n962) );
  NAND U1206 ( .A(n960), .B(n959), .Z(n961) );
  NAND U1207 ( .A(n962), .B(n961), .Z(n963) );
  XOR U1208 ( .A(n964), .B(n963), .Z(c[239]) );
  XOR U1209 ( .A(a[240]), .B(b[240]), .Z(n968) );
  NAND U1210 ( .A(a[239]), .B(b[239]), .Z(n966) );
  NAND U1211 ( .A(n964), .B(n963), .Z(n965) );
  NAND U1212 ( .A(n966), .B(n965), .Z(n967) );
  XOR U1213 ( .A(n968), .B(n967), .Z(c[240]) );
  XOR U1214 ( .A(a[241]), .B(b[241]), .Z(n972) );
  NAND U1215 ( .A(a[240]), .B(b[240]), .Z(n970) );
  NAND U1216 ( .A(n968), .B(n967), .Z(n969) );
  NAND U1217 ( .A(n970), .B(n969), .Z(n971) );
  XOR U1218 ( .A(n972), .B(n971), .Z(c[241]) );
  XOR U1219 ( .A(a[242]), .B(b[242]), .Z(n976) );
  NAND U1220 ( .A(a[241]), .B(b[241]), .Z(n974) );
  NAND U1221 ( .A(n972), .B(n971), .Z(n973) );
  NAND U1222 ( .A(n974), .B(n973), .Z(n975) );
  XOR U1223 ( .A(n976), .B(n975), .Z(c[242]) );
  XOR U1224 ( .A(a[243]), .B(b[243]), .Z(n980) );
  NAND U1225 ( .A(a[242]), .B(b[242]), .Z(n978) );
  NAND U1226 ( .A(n976), .B(n975), .Z(n977) );
  NAND U1227 ( .A(n978), .B(n977), .Z(n979) );
  XOR U1228 ( .A(n980), .B(n979), .Z(c[243]) );
  XOR U1229 ( .A(a[244]), .B(b[244]), .Z(n984) );
  NAND U1230 ( .A(a[243]), .B(b[243]), .Z(n982) );
  NAND U1231 ( .A(n980), .B(n979), .Z(n981) );
  NAND U1232 ( .A(n982), .B(n981), .Z(n983) );
  XOR U1233 ( .A(n984), .B(n983), .Z(c[244]) );
  XOR U1234 ( .A(a[245]), .B(b[245]), .Z(n988) );
  NAND U1235 ( .A(a[244]), .B(b[244]), .Z(n986) );
  NAND U1236 ( .A(n984), .B(n983), .Z(n985) );
  NAND U1237 ( .A(n986), .B(n985), .Z(n987) );
  XOR U1238 ( .A(n988), .B(n987), .Z(c[245]) );
  XOR U1239 ( .A(b[246]), .B(a[246]), .Z(n992) );
  NAND U1240 ( .A(a[245]), .B(b[245]), .Z(n990) );
  NAND U1241 ( .A(n988), .B(n987), .Z(n989) );
  AND U1242 ( .A(n990), .B(n989), .Z(n991) );
  XNOR U1243 ( .A(n992), .B(n991), .Z(c[246]) );
  OR U1244 ( .A(b[246]), .B(a[246]), .Z(n994) );
  NAND U1245 ( .A(n992), .B(n991), .Z(n993) );
  AND U1246 ( .A(n994), .B(n993), .Z(n996) );
  XOR U1247 ( .A(a[247]), .B(b[247]), .Z(n995) );
  XOR U1248 ( .A(n996), .B(n995), .Z(c[247]) );
  XOR U1249 ( .A(a[248]), .B(b[248]), .Z(n1000) );
  NAND U1250 ( .A(a[247]), .B(b[247]), .Z(n998) );
  NAND U1251 ( .A(n996), .B(n995), .Z(n997) );
  NAND U1252 ( .A(n998), .B(n997), .Z(n999) );
  XOR U1253 ( .A(n1000), .B(n999), .Z(c[248]) );
  XOR U1254 ( .A(a[249]), .B(b[249]), .Z(n1004) );
  NAND U1255 ( .A(a[248]), .B(b[248]), .Z(n1002) );
  NAND U1256 ( .A(n1000), .B(n999), .Z(n1001) );
  NAND U1257 ( .A(n1002), .B(n1001), .Z(n1003) );
  XOR U1258 ( .A(n1004), .B(n1003), .Z(c[249]) );
  XOR U1259 ( .A(a[250]), .B(b[250]), .Z(n1008) );
  NAND U1260 ( .A(a[249]), .B(b[249]), .Z(n1006) );
  NAND U1261 ( .A(n1004), .B(n1003), .Z(n1005) );
  NAND U1262 ( .A(n1006), .B(n1005), .Z(n1007) );
  XOR U1263 ( .A(n1008), .B(n1007), .Z(c[250]) );
  XOR U1264 ( .A(a[251]), .B(b[251]), .Z(n1012) );
  NAND U1265 ( .A(a[250]), .B(b[250]), .Z(n1010) );
  NAND U1266 ( .A(n1008), .B(n1007), .Z(n1009) );
  NAND U1267 ( .A(n1010), .B(n1009), .Z(n1011) );
  XOR U1268 ( .A(n1012), .B(n1011), .Z(c[251]) );
  XOR U1269 ( .A(a[252]), .B(b[252]), .Z(n1016) );
  NAND U1270 ( .A(a[251]), .B(b[251]), .Z(n1014) );
  NAND U1271 ( .A(n1012), .B(n1011), .Z(n1013) );
  NAND U1272 ( .A(n1014), .B(n1013), .Z(n1015) );
  XOR U1273 ( .A(n1016), .B(n1015), .Z(c[252]) );
  XOR U1274 ( .A(a[253]), .B(b[253]), .Z(n1020) );
  NAND U1275 ( .A(a[252]), .B(b[252]), .Z(n1018) );
  NAND U1276 ( .A(n1016), .B(n1015), .Z(n1017) );
  NAND U1277 ( .A(n1018), .B(n1017), .Z(n1019) );
  XOR U1278 ( .A(n1020), .B(n1019), .Z(c[253]) );
  XOR U1279 ( .A(a[254]), .B(b[254]), .Z(n1024) );
  NAND U1280 ( .A(a[253]), .B(b[253]), .Z(n1022) );
  NAND U1281 ( .A(n1020), .B(n1019), .Z(n1021) );
  NAND U1282 ( .A(n1022), .B(n1021), .Z(n1023) );
  XOR U1283 ( .A(n1024), .B(n1023), .Z(c[254]) );
  XOR U1284 ( .A(a[255]), .B(b[255]), .Z(n1028) );
  NAND U1285 ( .A(a[254]), .B(b[254]), .Z(n1026) );
  NAND U1286 ( .A(n1024), .B(n1023), .Z(n1025) );
  NAND U1287 ( .A(n1026), .B(n1025), .Z(n1027) );
  XOR U1288 ( .A(n1028), .B(n1027), .Z(c[255]) );
  XOR U1289 ( .A(a[256]), .B(b[256]), .Z(n1032) );
  NAND U1290 ( .A(a[255]), .B(b[255]), .Z(n1030) );
  NAND U1291 ( .A(n1028), .B(n1027), .Z(n1029) );
  NAND U1292 ( .A(n1030), .B(n1029), .Z(n1031) );
  XOR U1293 ( .A(n1032), .B(n1031), .Z(c[256]) );
  XOR U1294 ( .A(a[257]), .B(b[257]), .Z(n1036) );
  NAND U1295 ( .A(a[256]), .B(b[256]), .Z(n1034) );
  NAND U1296 ( .A(n1032), .B(n1031), .Z(n1033) );
  NAND U1297 ( .A(n1034), .B(n1033), .Z(n1035) );
  XOR U1298 ( .A(n1036), .B(n1035), .Z(c[257]) );
  XOR U1299 ( .A(a[258]), .B(b[258]), .Z(n1040) );
  NAND U1300 ( .A(a[257]), .B(b[257]), .Z(n1038) );
  NAND U1301 ( .A(n1036), .B(n1035), .Z(n1037) );
  NAND U1302 ( .A(n1038), .B(n1037), .Z(n1039) );
  XOR U1303 ( .A(n1040), .B(n1039), .Z(c[258]) );
  XOR U1304 ( .A(a[259]), .B(b[259]), .Z(n1044) );
  NAND U1305 ( .A(a[258]), .B(b[258]), .Z(n1042) );
  NAND U1306 ( .A(n1040), .B(n1039), .Z(n1041) );
  NAND U1307 ( .A(n1042), .B(n1041), .Z(n1043) );
  XOR U1308 ( .A(n1044), .B(n1043), .Z(c[259]) );
  XOR U1309 ( .A(a[260]), .B(b[260]), .Z(n1048) );
  NAND U1310 ( .A(a[259]), .B(b[259]), .Z(n1046) );
  NAND U1311 ( .A(n1044), .B(n1043), .Z(n1045) );
  NAND U1312 ( .A(n1046), .B(n1045), .Z(n1047) );
  XOR U1313 ( .A(n1048), .B(n1047), .Z(c[260]) );
  XOR U1314 ( .A(a[261]), .B(b[261]), .Z(n1052) );
  NAND U1315 ( .A(a[260]), .B(b[260]), .Z(n1050) );
  NAND U1316 ( .A(n1048), .B(n1047), .Z(n1049) );
  NAND U1317 ( .A(n1050), .B(n1049), .Z(n1051) );
  XOR U1318 ( .A(n1052), .B(n1051), .Z(c[261]) );
  XOR U1319 ( .A(a[262]), .B(b[262]), .Z(n1056) );
  NAND U1320 ( .A(a[261]), .B(b[261]), .Z(n1054) );
  NAND U1321 ( .A(n1052), .B(n1051), .Z(n1053) );
  NAND U1322 ( .A(n1054), .B(n1053), .Z(n1055) );
  XOR U1323 ( .A(n1056), .B(n1055), .Z(c[262]) );
  NAND U1324 ( .A(a[262]), .B(b[262]), .Z(n1058) );
  NAND U1325 ( .A(n1056), .B(n1055), .Z(n1057) );
  AND U1326 ( .A(n1058), .B(n1057), .Z(n1060) );
  XOR U1327 ( .A(b[263]), .B(a[263]), .Z(n1059) );
  XNOR U1328 ( .A(n1060), .B(n1059), .Z(c[263]) );
  OR U1329 ( .A(b[263]), .B(a[263]), .Z(n1062) );
  NAND U1330 ( .A(n1060), .B(n1059), .Z(n1061) );
  AND U1331 ( .A(n1062), .B(n1061), .Z(n1064) );
  XOR U1332 ( .A(a[264]), .B(b[264]), .Z(n1063) );
  XOR U1333 ( .A(n1064), .B(n1063), .Z(c[264]) );
  XOR U1334 ( .A(a[265]), .B(b[265]), .Z(n1068) );
  NAND U1335 ( .A(a[264]), .B(b[264]), .Z(n1066) );
  NAND U1336 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1337 ( .A(n1066), .B(n1065), .Z(n1067) );
  XOR U1338 ( .A(n1068), .B(n1067), .Z(c[265]) );
  NAND U1339 ( .A(a[265]), .B(b[265]), .Z(n1070) );
  NAND U1340 ( .A(n1068), .B(n1067), .Z(n1069) );
  AND U1341 ( .A(n1070), .B(n1069), .Z(n1072) );
  XOR U1342 ( .A(b[266]), .B(a[266]), .Z(n1071) );
  XNOR U1343 ( .A(n1072), .B(n1071), .Z(c[266]) );
  OR U1344 ( .A(b[266]), .B(a[266]), .Z(n1074) );
  NAND U1345 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U1346 ( .A(n1074), .B(n1073), .Z(n1076) );
  XOR U1347 ( .A(a[267]), .B(b[267]), .Z(n1075) );
  XOR U1348 ( .A(n1076), .B(n1075), .Z(c[267]) );
  XOR U1349 ( .A(a[268]), .B(b[268]), .Z(n1080) );
  NAND U1350 ( .A(a[267]), .B(b[267]), .Z(n1078) );
  NAND U1351 ( .A(n1076), .B(n1075), .Z(n1077) );
  NAND U1352 ( .A(n1078), .B(n1077), .Z(n1079) );
  XOR U1353 ( .A(n1080), .B(n1079), .Z(c[268]) );
  XOR U1354 ( .A(a[269]), .B(b[269]), .Z(n1084) );
  NAND U1355 ( .A(a[268]), .B(b[268]), .Z(n1082) );
  NAND U1356 ( .A(n1080), .B(n1079), .Z(n1081) );
  NAND U1357 ( .A(n1082), .B(n1081), .Z(n1083) );
  XOR U1358 ( .A(n1084), .B(n1083), .Z(c[269]) );
  XOR U1359 ( .A(a[270]), .B(b[270]), .Z(n1088) );
  NAND U1360 ( .A(a[269]), .B(b[269]), .Z(n1086) );
  NAND U1361 ( .A(n1084), .B(n1083), .Z(n1085) );
  NAND U1362 ( .A(n1086), .B(n1085), .Z(n1087) );
  XOR U1363 ( .A(n1088), .B(n1087), .Z(c[270]) );
  XOR U1364 ( .A(a[271]), .B(b[271]), .Z(n1092) );
  NAND U1365 ( .A(a[270]), .B(b[270]), .Z(n1090) );
  NAND U1366 ( .A(n1088), .B(n1087), .Z(n1089) );
  NAND U1367 ( .A(n1090), .B(n1089), .Z(n1091) );
  XOR U1368 ( .A(n1092), .B(n1091), .Z(c[271]) );
  XOR U1369 ( .A(a[272]), .B(b[272]), .Z(n1096) );
  NAND U1370 ( .A(a[271]), .B(b[271]), .Z(n1094) );
  NAND U1371 ( .A(n1092), .B(n1091), .Z(n1093) );
  NAND U1372 ( .A(n1094), .B(n1093), .Z(n1095) );
  XOR U1373 ( .A(n1096), .B(n1095), .Z(c[272]) );
  XOR U1374 ( .A(a[273]), .B(b[273]), .Z(n1100) );
  NAND U1375 ( .A(a[272]), .B(b[272]), .Z(n1098) );
  NAND U1376 ( .A(n1096), .B(n1095), .Z(n1097) );
  NAND U1377 ( .A(n1098), .B(n1097), .Z(n1099) );
  XOR U1378 ( .A(n1100), .B(n1099), .Z(c[273]) );
  XOR U1379 ( .A(a[274]), .B(b[274]), .Z(n1104) );
  NAND U1380 ( .A(a[273]), .B(b[273]), .Z(n1102) );
  NAND U1381 ( .A(n1100), .B(n1099), .Z(n1101) );
  NAND U1382 ( .A(n1102), .B(n1101), .Z(n1103) );
  XOR U1383 ( .A(n1104), .B(n1103), .Z(c[274]) );
  XOR U1384 ( .A(a[275]), .B(b[275]), .Z(n1108) );
  NAND U1385 ( .A(a[274]), .B(b[274]), .Z(n1106) );
  NAND U1386 ( .A(n1104), .B(n1103), .Z(n1105) );
  NAND U1387 ( .A(n1106), .B(n1105), .Z(n1107) );
  XOR U1388 ( .A(n1108), .B(n1107), .Z(c[275]) );
  XOR U1389 ( .A(a[276]), .B(b[276]), .Z(n1112) );
  NAND U1390 ( .A(a[275]), .B(b[275]), .Z(n1110) );
  NAND U1391 ( .A(n1108), .B(n1107), .Z(n1109) );
  NAND U1392 ( .A(n1110), .B(n1109), .Z(n1111) );
  XOR U1393 ( .A(n1112), .B(n1111), .Z(c[276]) );
  XOR U1394 ( .A(a[277]), .B(b[277]), .Z(n1116) );
  NAND U1395 ( .A(a[276]), .B(b[276]), .Z(n1114) );
  NAND U1396 ( .A(n1112), .B(n1111), .Z(n1113) );
  NAND U1397 ( .A(n1114), .B(n1113), .Z(n1115) );
  XOR U1398 ( .A(n1116), .B(n1115), .Z(c[277]) );
  XOR U1399 ( .A(a[278]), .B(b[278]), .Z(n1120) );
  NAND U1400 ( .A(a[277]), .B(b[277]), .Z(n1118) );
  NAND U1401 ( .A(n1116), .B(n1115), .Z(n1117) );
  NAND U1402 ( .A(n1118), .B(n1117), .Z(n1119) );
  XOR U1403 ( .A(n1120), .B(n1119), .Z(c[278]) );
  XOR U1404 ( .A(a[279]), .B(b[279]), .Z(n1124) );
  NAND U1405 ( .A(a[278]), .B(b[278]), .Z(n1122) );
  NAND U1406 ( .A(n1120), .B(n1119), .Z(n1121) );
  NAND U1407 ( .A(n1122), .B(n1121), .Z(n1123) );
  XOR U1408 ( .A(n1124), .B(n1123), .Z(c[279]) );
  XOR U1409 ( .A(a[280]), .B(b[280]), .Z(n1128) );
  NAND U1410 ( .A(a[279]), .B(b[279]), .Z(n1126) );
  NAND U1411 ( .A(n1124), .B(n1123), .Z(n1125) );
  NAND U1412 ( .A(n1126), .B(n1125), .Z(n1127) );
  XOR U1413 ( .A(n1128), .B(n1127), .Z(c[280]) );
  XOR U1414 ( .A(a[281]), .B(b[281]), .Z(n1132) );
  NAND U1415 ( .A(a[280]), .B(b[280]), .Z(n1130) );
  NAND U1416 ( .A(n1128), .B(n1127), .Z(n1129) );
  NAND U1417 ( .A(n1130), .B(n1129), .Z(n1131) );
  XOR U1418 ( .A(n1132), .B(n1131), .Z(c[281]) );
  XOR U1419 ( .A(a[282]), .B(b[282]), .Z(n1136) );
  NAND U1420 ( .A(a[281]), .B(b[281]), .Z(n1134) );
  NAND U1421 ( .A(n1132), .B(n1131), .Z(n1133) );
  NAND U1422 ( .A(n1134), .B(n1133), .Z(n1135) );
  XOR U1423 ( .A(n1136), .B(n1135), .Z(c[282]) );
  XOR U1424 ( .A(a[283]), .B(b[283]), .Z(n1140) );
  NAND U1425 ( .A(a[282]), .B(b[282]), .Z(n1138) );
  NAND U1426 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U1427 ( .A(n1138), .B(n1137), .Z(n1139) );
  XOR U1428 ( .A(n1140), .B(n1139), .Z(c[283]) );
  XOR U1429 ( .A(a[284]), .B(b[284]), .Z(n1144) );
  NAND U1430 ( .A(a[283]), .B(b[283]), .Z(n1142) );
  NAND U1431 ( .A(n1140), .B(n1139), .Z(n1141) );
  NAND U1432 ( .A(n1142), .B(n1141), .Z(n1143) );
  XOR U1433 ( .A(n1144), .B(n1143), .Z(c[284]) );
  XOR U1434 ( .A(a[285]), .B(b[285]), .Z(n1148) );
  NAND U1435 ( .A(a[284]), .B(b[284]), .Z(n1146) );
  NAND U1436 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U1437 ( .A(n1146), .B(n1145), .Z(n1147) );
  XOR U1438 ( .A(n1148), .B(n1147), .Z(c[285]) );
  XOR U1439 ( .A(a[286]), .B(b[286]), .Z(n1152) );
  NAND U1440 ( .A(a[285]), .B(b[285]), .Z(n1150) );
  NAND U1441 ( .A(n1148), .B(n1147), .Z(n1149) );
  NAND U1442 ( .A(n1150), .B(n1149), .Z(n1151) );
  XOR U1443 ( .A(n1152), .B(n1151), .Z(c[286]) );
  XOR U1444 ( .A(a[287]), .B(b[287]), .Z(n1156) );
  NAND U1445 ( .A(a[286]), .B(b[286]), .Z(n1154) );
  NAND U1446 ( .A(n1152), .B(n1151), .Z(n1153) );
  NAND U1447 ( .A(n1154), .B(n1153), .Z(n1155) );
  XOR U1448 ( .A(n1156), .B(n1155), .Z(c[287]) );
  XOR U1449 ( .A(a[288]), .B(b[288]), .Z(n1160) );
  NAND U1450 ( .A(a[287]), .B(b[287]), .Z(n1158) );
  NAND U1451 ( .A(n1156), .B(n1155), .Z(n1157) );
  NAND U1452 ( .A(n1158), .B(n1157), .Z(n1159) );
  XOR U1453 ( .A(n1160), .B(n1159), .Z(c[288]) );
  XOR U1454 ( .A(a[289]), .B(b[289]), .Z(n1164) );
  NAND U1455 ( .A(a[288]), .B(b[288]), .Z(n1162) );
  NAND U1456 ( .A(n1160), .B(n1159), .Z(n1161) );
  NAND U1457 ( .A(n1162), .B(n1161), .Z(n1163) );
  XOR U1458 ( .A(n1164), .B(n1163), .Z(c[289]) );
  XOR U1459 ( .A(a[290]), .B(b[290]), .Z(n1168) );
  NAND U1460 ( .A(a[289]), .B(b[289]), .Z(n1166) );
  NAND U1461 ( .A(n1164), .B(n1163), .Z(n1165) );
  NAND U1462 ( .A(n1166), .B(n1165), .Z(n1167) );
  XOR U1463 ( .A(n1168), .B(n1167), .Z(c[290]) );
  XOR U1464 ( .A(a[291]), .B(b[291]), .Z(n1172) );
  NAND U1465 ( .A(a[290]), .B(b[290]), .Z(n1170) );
  NAND U1466 ( .A(n1168), .B(n1167), .Z(n1169) );
  NAND U1467 ( .A(n1170), .B(n1169), .Z(n1171) );
  XOR U1468 ( .A(n1172), .B(n1171), .Z(c[291]) );
  XOR U1469 ( .A(a[292]), .B(b[292]), .Z(n1176) );
  NAND U1470 ( .A(a[291]), .B(b[291]), .Z(n1174) );
  NAND U1471 ( .A(n1172), .B(n1171), .Z(n1173) );
  NAND U1472 ( .A(n1174), .B(n1173), .Z(n1175) );
  XOR U1473 ( .A(n1176), .B(n1175), .Z(c[292]) );
  XOR U1474 ( .A(a[293]), .B(b[293]), .Z(n1180) );
  NAND U1475 ( .A(a[292]), .B(b[292]), .Z(n1178) );
  NAND U1476 ( .A(n1176), .B(n1175), .Z(n1177) );
  NAND U1477 ( .A(n1178), .B(n1177), .Z(n1179) );
  XOR U1478 ( .A(n1180), .B(n1179), .Z(c[293]) );
  XOR U1479 ( .A(a[294]), .B(b[294]), .Z(n1184) );
  NAND U1480 ( .A(a[293]), .B(b[293]), .Z(n1182) );
  NAND U1481 ( .A(n1180), .B(n1179), .Z(n1181) );
  NAND U1482 ( .A(n1182), .B(n1181), .Z(n1183) );
  XOR U1483 ( .A(n1184), .B(n1183), .Z(c[294]) );
  XOR U1484 ( .A(a[295]), .B(b[295]), .Z(n1188) );
  NAND U1485 ( .A(a[294]), .B(b[294]), .Z(n1186) );
  NAND U1486 ( .A(n1184), .B(n1183), .Z(n1185) );
  NAND U1487 ( .A(n1186), .B(n1185), .Z(n1187) );
  XOR U1488 ( .A(n1188), .B(n1187), .Z(c[295]) );
  XOR U1489 ( .A(a[296]), .B(b[296]), .Z(n1192) );
  NAND U1490 ( .A(a[295]), .B(b[295]), .Z(n1190) );
  NAND U1491 ( .A(n1188), .B(n1187), .Z(n1189) );
  NAND U1492 ( .A(n1190), .B(n1189), .Z(n1191) );
  XOR U1493 ( .A(n1192), .B(n1191), .Z(c[296]) );
  XOR U1494 ( .A(a[297]), .B(b[297]), .Z(n1196) );
  NAND U1495 ( .A(a[296]), .B(b[296]), .Z(n1194) );
  NAND U1496 ( .A(n1192), .B(n1191), .Z(n1193) );
  NAND U1497 ( .A(n1194), .B(n1193), .Z(n1195) );
  XOR U1498 ( .A(n1196), .B(n1195), .Z(c[297]) );
  XOR U1499 ( .A(a[298]), .B(b[298]), .Z(n1200) );
  NAND U1500 ( .A(a[297]), .B(b[297]), .Z(n1198) );
  NAND U1501 ( .A(n1196), .B(n1195), .Z(n1197) );
  NAND U1502 ( .A(n1198), .B(n1197), .Z(n1199) );
  XOR U1503 ( .A(n1200), .B(n1199), .Z(c[298]) );
  NAND U1504 ( .A(a[298]), .B(b[298]), .Z(n1202) );
  NAND U1505 ( .A(n1200), .B(n1199), .Z(n1201) );
  AND U1506 ( .A(n1202), .B(n1201), .Z(n1204) );
  XOR U1507 ( .A(b[299]), .B(a[299]), .Z(n1203) );
  XNOR U1508 ( .A(n1204), .B(n1203), .Z(c[299]) );
  OR U1509 ( .A(b[299]), .B(a[299]), .Z(n1206) );
  NAND U1510 ( .A(n1204), .B(n1203), .Z(n1205) );
  AND U1511 ( .A(n1206), .B(n1205), .Z(n1208) );
  XOR U1512 ( .A(a[300]), .B(b[300]), .Z(n1207) );
  XOR U1513 ( .A(n1208), .B(n1207), .Z(c[300]) );
  XOR U1514 ( .A(a[301]), .B(b[301]), .Z(n1212) );
  NAND U1515 ( .A(a[300]), .B(b[300]), .Z(n1210) );
  NAND U1516 ( .A(n1208), .B(n1207), .Z(n1209) );
  NAND U1517 ( .A(n1210), .B(n1209), .Z(n1211) );
  XOR U1518 ( .A(n1212), .B(n1211), .Z(c[301]) );
  XOR U1519 ( .A(b[302]), .B(a[302]), .Z(n1216) );
  NAND U1520 ( .A(a[301]), .B(b[301]), .Z(n1214) );
  NAND U1521 ( .A(n1212), .B(n1211), .Z(n1213) );
  AND U1522 ( .A(n1214), .B(n1213), .Z(n1215) );
  XNOR U1523 ( .A(n1216), .B(n1215), .Z(c[302]) );
  XOR U1524 ( .A(a[303]), .B(b[303]), .Z(n1220) );
  OR U1525 ( .A(b[302]), .B(a[302]), .Z(n1218) );
  NAND U1526 ( .A(n1216), .B(n1215), .Z(n1217) );
  AND U1527 ( .A(n1218), .B(n1217), .Z(n1219) );
  XOR U1528 ( .A(n1220), .B(n1219), .Z(c[303]) );
  XOR U1529 ( .A(a[304]), .B(b[304]), .Z(n1224) );
  NAND U1530 ( .A(a[303]), .B(b[303]), .Z(n1222) );
  NAND U1531 ( .A(n1220), .B(n1219), .Z(n1221) );
  NAND U1532 ( .A(n1222), .B(n1221), .Z(n1223) );
  XOR U1533 ( .A(n1224), .B(n1223), .Z(c[304]) );
  XOR U1534 ( .A(a[305]), .B(b[305]), .Z(n1228) );
  NAND U1535 ( .A(a[304]), .B(b[304]), .Z(n1226) );
  NAND U1536 ( .A(n1224), .B(n1223), .Z(n1225) );
  NAND U1537 ( .A(n1226), .B(n1225), .Z(n1227) );
  XOR U1538 ( .A(n1228), .B(n1227), .Z(c[305]) );
  XOR U1539 ( .A(a[306]), .B(b[306]), .Z(n1232) );
  NAND U1540 ( .A(a[305]), .B(b[305]), .Z(n1230) );
  NAND U1541 ( .A(n1228), .B(n1227), .Z(n1229) );
  NAND U1542 ( .A(n1230), .B(n1229), .Z(n1231) );
  XOR U1543 ( .A(n1232), .B(n1231), .Z(c[306]) );
  XOR U1544 ( .A(a[307]), .B(b[307]), .Z(n1236) );
  NAND U1545 ( .A(a[306]), .B(b[306]), .Z(n1234) );
  NAND U1546 ( .A(n1232), .B(n1231), .Z(n1233) );
  NAND U1547 ( .A(n1234), .B(n1233), .Z(n1235) );
  XOR U1548 ( .A(n1236), .B(n1235), .Z(c[307]) );
  XOR U1549 ( .A(a[308]), .B(b[308]), .Z(n1240) );
  NAND U1550 ( .A(a[307]), .B(b[307]), .Z(n1238) );
  NAND U1551 ( .A(n1236), .B(n1235), .Z(n1237) );
  NAND U1552 ( .A(n1238), .B(n1237), .Z(n1239) );
  XOR U1553 ( .A(n1240), .B(n1239), .Z(c[308]) );
  XOR U1554 ( .A(a[309]), .B(b[309]), .Z(n1244) );
  NAND U1555 ( .A(a[308]), .B(b[308]), .Z(n1242) );
  NAND U1556 ( .A(n1240), .B(n1239), .Z(n1241) );
  NAND U1557 ( .A(n1242), .B(n1241), .Z(n1243) );
  XOR U1558 ( .A(n1244), .B(n1243), .Z(c[309]) );
  XOR U1559 ( .A(a[310]), .B(b[310]), .Z(n1248) );
  NAND U1560 ( .A(a[309]), .B(b[309]), .Z(n1246) );
  NAND U1561 ( .A(n1244), .B(n1243), .Z(n1245) );
  NAND U1562 ( .A(n1246), .B(n1245), .Z(n1247) );
  XOR U1563 ( .A(n1248), .B(n1247), .Z(c[310]) );
  XOR U1564 ( .A(a[311]), .B(b[311]), .Z(n1252) );
  NAND U1565 ( .A(a[310]), .B(b[310]), .Z(n1250) );
  NAND U1566 ( .A(n1248), .B(n1247), .Z(n1249) );
  NAND U1567 ( .A(n1250), .B(n1249), .Z(n1251) );
  XOR U1568 ( .A(n1252), .B(n1251), .Z(c[311]) );
  XOR U1569 ( .A(a[312]), .B(b[312]), .Z(n1256) );
  NAND U1570 ( .A(a[311]), .B(b[311]), .Z(n1254) );
  NAND U1571 ( .A(n1252), .B(n1251), .Z(n1253) );
  NAND U1572 ( .A(n1254), .B(n1253), .Z(n1255) );
  XOR U1573 ( .A(n1256), .B(n1255), .Z(c[312]) );
  XOR U1574 ( .A(a[313]), .B(b[313]), .Z(n1260) );
  NAND U1575 ( .A(a[312]), .B(b[312]), .Z(n1258) );
  NAND U1576 ( .A(n1256), .B(n1255), .Z(n1257) );
  NAND U1577 ( .A(n1258), .B(n1257), .Z(n1259) );
  XOR U1578 ( .A(n1260), .B(n1259), .Z(c[313]) );
  XOR U1579 ( .A(a[314]), .B(b[314]), .Z(n1264) );
  NAND U1580 ( .A(a[313]), .B(b[313]), .Z(n1262) );
  NAND U1581 ( .A(n1260), .B(n1259), .Z(n1261) );
  NAND U1582 ( .A(n1262), .B(n1261), .Z(n1263) );
  XOR U1583 ( .A(n1264), .B(n1263), .Z(c[314]) );
  XOR U1584 ( .A(a[315]), .B(b[315]), .Z(n1268) );
  NAND U1585 ( .A(a[314]), .B(b[314]), .Z(n1266) );
  NAND U1586 ( .A(n1264), .B(n1263), .Z(n1265) );
  NAND U1587 ( .A(n1266), .B(n1265), .Z(n1267) );
  XOR U1588 ( .A(n1268), .B(n1267), .Z(c[315]) );
  XOR U1589 ( .A(a[316]), .B(b[316]), .Z(n1272) );
  NAND U1590 ( .A(a[315]), .B(b[315]), .Z(n1270) );
  NAND U1591 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U1592 ( .A(n1270), .B(n1269), .Z(n1271) );
  XOR U1593 ( .A(n1272), .B(n1271), .Z(c[316]) );
  XOR U1594 ( .A(a[317]), .B(b[317]), .Z(n1276) );
  NAND U1595 ( .A(a[316]), .B(b[316]), .Z(n1274) );
  NAND U1596 ( .A(n1272), .B(n1271), .Z(n1273) );
  NAND U1597 ( .A(n1274), .B(n1273), .Z(n1275) );
  XOR U1598 ( .A(n1276), .B(n1275), .Z(c[317]) );
  XOR U1599 ( .A(a[318]), .B(b[318]), .Z(n1280) );
  NAND U1600 ( .A(a[317]), .B(b[317]), .Z(n1278) );
  NAND U1601 ( .A(n1276), .B(n1275), .Z(n1277) );
  NAND U1602 ( .A(n1278), .B(n1277), .Z(n1279) );
  XOR U1603 ( .A(n1280), .B(n1279), .Z(c[318]) );
  XOR U1604 ( .A(b[319]), .B(a[319]), .Z(n1284) );
  NAND U1605 ( .A(a[318]), .B(b[318]), .Z(n1282) );
  NAND U1606 ( .A(n1280), .B(n1279), .Z(n1281) );
  AND U1607 ( .A(n1282), .B(n1281), .Z(n1283) );
  XNOR U1608 ( .A(n1284), .B(n1283), .Z(c[319]) );
  OR U1609 ( .A(b[319]), .B(a[319]), .Z(n1286) );
  NAND U1610 ( .A(n1284), .B(n1283), .Z(n1285) );
  AND U1611 ( .A(n1286), .B(n1285), .Z(n1288) );
  XOR U1612 ( .A(a[320]), .B(b[320]), .Z(n1287) );
  XOR U1613 ( .A(n1288), .B(n1287), .Z(c[320]) );
  XOR U1614 ( .A(a[321]), .B(b[321]), .Z(n1292) );
  NAND U1615 ( .A(a[320]), .B(b[320]), .Z(n1290) );
  NAND U1616 ( .A(n1288), .B(n1287), .Z(n1289) );
  NAND U1617 ( .A(n1290), .B(n1289), .Z(n1291) );
  XOR U1618 ( .A(n1292), .B(n1291), .Z(c[321]) );
  XOR U1619 ( .A(a[322]), .B(b[322]), .Z(n1296) );
  NAND U1620 ( .A(a[321]), .B(b[321]), .Z(n1294) );
  NAND U1621 ( .A(n1292), .B(n1291), .Z(n1293) );
  NAND U1622 ( .A(n1294), .B(n1293), .Z(n1295) );
  XOR U1623 ( .A(n1296), .B(n1295), .Z(c[322]) );
  XOR U1624 ( .A(a[323]), .B(b[323]), .Z(n1300) );
  NAND U1625 ( .A(a[322]), .B(b[322]), .Z(n1298) );
  NAND U1626 ( .A(n1296), .B(n1295), .Z(n1297) );
  NAND U1627 ( .A(n1298), .B(n1297), .Z(n1299) );
  XOR U1628 ( .A(n1300), .B(n1299), .Z(c[323]) );
  XOR U1629 ( .A(a[324]), .B(b[324]), .Z(n1304) );
  NAND U1630 ( .A(a[323]), .B(b[323]), .Z(n1302) );
  NAND U1631 ( .A(n1300), .B(n1299), .Z(n1301) );
  NAND U1632 ( .A(n1302), .B(n1301), .Z(n1303) );
  XOR U1633 ( .A(n1304), .B(n1303), .Z(c[324]) );
  XOR U1634 ( .A(a[325]), .B(b[325]), .Z(n1308) );
  NAND U1635 ( .A(a[324]), .B(b[324]), .Z(n1306) );
  NAND U1636 ( .A(n1304), .B(n1303), .Z(n1305) );
  NAND U1637 ( .A(n1306), .B(n1305), .Z(n1307) );
  XOR U1638 ( .A(n1308), .B(n1307), .Z(c[325]) );
  XOR U1639 ( .A(a[326]), .B(b[326]), .Z(n1312) );
  NAND U1640 ( .A(a[325]), .B(b[325]), .Z(n1310) );
  NAND U1641 ( .A(n1308), .B(n1307), .Z(n1309) );
  NAND U1642 ( .A(n1310), .B(n1309), .Z(n1311) );
  XOR U1643 ( .A(n1312), .B(n1311), .Z(c[326]) );
  XOR U1644 ( .A(a[327]), .B(b[327]), .Z(n1316) );
  NAND U1645 ( .A(a[326]), .B(b[326]), .Z(n1314) );
  NAND U1646 ( .A(n1312), .B(n1311), .Z(n1313) );
  NAND U1647 ( .A(n1314), .B(n1313), .Z(n1315) );
  XOR U1648 ( .A(n1316), .B(n1315), .Z(c[327]) );
  XOR U1649 ( .A(a[328]), .B(b[328]), .Z(n1320) );
  NAND U1650 ( .A(a[327]), .B(b[327]), .Z(n1318) );
  NAND U1651 ( .A(n1316), .B(n1315), .Z(n1317) );
  NAND U1652 ( .A(n1318), .B(n1317), .Z(n1319) );
  XOR U1653 ( .A(n1320), .B(n1319), .Z(c[328]) );
  XOR U1654 ( .A(a[329]), .B(b[329]), .Z(n1324) );
  NAND U1655 ( .A(a[328]), .B(b[328]), .Z(n1322) );
  NAND U1656 ( .A(n1320), .B(n1319), .Z(n1321) );
  NAND U1657 ( .A(n1322), .B(n1321), .Z(n1323) );
  XOR U1658 ( .A(n1324), .B(n1323), .Z(c[329]) );
  XOR U1659 ( .A(a[330]), .B(b[330]), .Z(n1328) );
  NAND U1660 ( .A(a[329]), .B(b[329]), .Z(n1326) );
  NAND U1661 ( .A(n1324), .B(n1323), .Z(n1325) );
  NAND U1662 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U1663 ( .A(n1328), .B(n1327), .Z(c[330]) );
  XOR U1664 ( .A(a[331]), .B(b[331]), .Z(n1332) );
  NAND U1665 ( .A(a[330]), .B(b[330]), .Z(n1330) );
  NAND U1666 ( .A(n1328), .B(n1327), .Z(n1329) );
  NAND U1667 ( .A(n1330), .B(n1329), .Z(n1331) );
  XOR U1668 ( .A(n1332), .B(n1331), .Z(c[331]) );
  XOR U1669 ( .A(a[332]), .B(b[332]), .Z(n1336) );
  NAND U1670 ( .A(a[331]), .B(b[331]), .Z(n1334) );
  NAND U1671 ( .A(n1332), .B(n1331), .Z(n1333) );
  NAND U1672 ( .A(n1334), .B(n1333), .Z(n1335) );
  XOR U1673 ( .A(n1336), .B(n1335), .Z(c[332]) );
  XOR U1674 ( .A(b[333]), .B(a[333]), .Z(n1340) );
  NAND U1675 ( .A(a[332]), .B(b[332]), .Z(n1338) );
  NAND U1676 ( .A(n1336), .B(n1335), .Z(n1337) );
  AND U1677 ( .A(n1338), .B(n1337), .Z(n1339) );
  XNOR U1678 ( .A(n1340), .B(n1339), .Z(c[333]) );
  OR U1679 ( .A(b[333]), .B(a[333]), .Z(n1342) );
  NAND U1680 ( .A(n1340), .B(n1339), .Z(n1341) );
  AND U1681 ( .A(n1342), .B(n1341), .Z(n1344) );
  XOR U1682 ( .A(a[334]), .B(b[334]), .Z(n1343) );
  XOR U1683 ( .A(n1344), .B(n1343), .Z(c[334]) );
  XOR U1684 ( .A(a[335]), .B(b[335]), .Z(n1348) );
  NAND U1685 ( .A(a[334]), .B(b[334]), .Z(n1346) );
  NAND U1686 ( .A(n1344), .B(n1343), .Z(n1345) );
  NAND U1687 ( .A(n1346), .B(n1345), .Z(n1347) );
  XOR U1688 ( .A(n1348), .B(n1347), .Z(c[335]) );
  XOR U1689 ( .A(a[336]), .B(b[336]), .Z(n1352) );
  NAND U1690 ( .A(a[335]), .B(b[335]), .Z(n1350) );
  NAND U1691 ( .A(n1348), .B(n1347), .Z(n1349) );
  NAND U1692 ( .A(n1350), .B(n1349), .Z(n1351) );
  XOR U1693 ( .A(n1352), .B(n1351), .Z(c[336]) );
  XOR U1694 ( .A(a[337]), .B(b[337]), .Z(n1356) );
  NAND U1695 ( .A(a[336]), .B(b[336]), .Z(n1354) );
  NAND U1696 ( .A(n1352), .B(n1351), .Z(n1353) );
  NAND U1697 ( .A(n1354), .B(n1353), .Z(n1355) );
  XOR U1698 ( .A(n1356), .B(n1355), .Z(c[337]) );
  XOR U1699 ( .A(a[338]), .B(b[338]), .Z(n1360) );
  NAND U1700 ( .A(a[337]), .B(b[337]), .Z(n1358) );
  NAND U1701 ( .A(n1356), .B(n1355), .Z(n1357) );
  NAND U1702 ( .A(n1358), .B(n1357), .Z(n1359) );
  XOR U1703 ( .A(n1360), .B(n1359), .Z(c[338]) );
  XOR U1704 ( .A(a[339]), .B(b[339]), .Z(n1364) );
  NAND U1705 ( .A(a[338]), .B(b[338]), .Z(n1362) );
  NAND U1706 ( .A(n1360), .B(n1359), .Z(n1361) );
  NAND U1707 ( .A(n1362), .B(n1361), .Z(n1363) );
  XOR U1708 ( .A(n1364), .B(n1363), .Z(c[339]) );
  XOR U1709 ( .A(a[340]), .B(b[340]), .Z(n1368) );
  NAND U1710 ( .A(a[339]), .B(b[339]), .Z(n1366) );
  NAND U1711 ( .A(n1364), .B(n1363), .Z(n1365) );
  NAND U1712 ( .A(n1366), .B(n1365), .Z(n1367) );
  XOR U1713 ( .A(n1368), .B(n1367), .Z(c[340]) );
  XOR U1714 ( .A(a[341]), .B(b[341]), .Z(n1372) );
  NAND U1715 ( .A(a[340]), .B(b[340]), .Z(n1370) );
  NAND U1716 ( .A(n1368), .B(n1367), .Z(n1369) );
  NAND U1717 ( .A(n1370), .B(n1369), .Z(n1371) );
  XOR U1718 ( .A(n1372), .B(n1371), .Z(c[341]) );
  XOR U1719 ( .A(a[342]), .B(b[342]), .Z(n1376) );
  NAND U1720 ( .A(a[341]), .B(b[341]), .Z(n1374) );
  NAND U1721 ( .A(n1372), .B(n1371), .Z(n1373) );
  NAND U1722 ( .A(n1374), .B(n1373), .Z(n1375) );
  XOR U1723 ( .A(n1376), .B(n1375), .Z(c[342]) );
  XOR U1724 ( .A(a[343]), .B(b[343]), .Z(n1380) );
  NAND U1725 ( .A(a[342]), .B(b[342]), .Z(n1378) );
  NAND U1726 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U1727 ( .A(n1378), .B(n1377), .Z(n1379) );
  XOR U1728 ( .A(n1380), .B(n1379), .Z(c[343]) );
  XOR U1729 ( .A(a[344]), .B(b[344]), .Z(n1384) );
  NAND U1730 ( .A(a[343]), .B(b[343]), .Z(n1382) );
  NAND U1731 ( .A(n1380), .B(n1379), .Z(n1381) );
  NAND U1732 ( .A(n1382), .B(n1381), .Z(n1383) );
  XOR U1733 ( .A(n1384), .B(n1383), .Z(c[344]) );
  XOR U1734 ( .A(a[345]), .B(b[345]), .Z(n1388) );
  NAND U1735 ( .A(a[344]), .B(b[344]), .Z(n1386) );
  NAND U1736 ( .A(n1384), .B(n1383), .Z(n1385) );
  NAND U1737 ( .A(n1386), .B(n1385), .Z(n1387) );
  XOR U1738 ( .A(n1388), .B(n1387), .Z(c[345]) );
  XOR U1739 ( .A(a[346]), .B(b[346]), .Z(n1392) );
  NAND U1740 ( .A(a[345]), .B(b[345]), .Z(n1390) );
  NAND U1741 ( .A(n1388), .B(n1387), .Z(n1389) );
  NAND U1742 ( .A(n1390), .B(n1389), .Z(n1391) );
  XOR U1743 ( .A(n1392), .B(n1391), .Z(c[346]) );
  XOR U1744 ( .A(a[347]), .B(b[347]), .Z(n1396) );
  NAND U1745 ( .A(a[346]), .B(b[346]), .Z(n1394) );
  NAND U1746 ( .A(n1392), .B(n1391), .Z(n1393) );
  NAND U1747 ( .A(n1394), .B(n1393), .Z(n1395) );
  XOR U1748 ( .A(n1396), .B(n1395), .Z(c[347]) );
  XOR U1749 ( .A(a[348]), .B(b[348]), .Z(n1400) );
  NAND U1750 ( .A(a[347]), .B(b[347]), .Z(n1398) );
  NAND U1751 ( .A(n1396), .B(n1395), .Z(n1397) );
  NAND U1752 ( .A(n1398), .B(n1397), .Z(n1399) );
  XOR U1753 ( .A(n1400), .B(n1399), .Z(c[348]) );
  XOR U1754 ( .A(a[349]), .B(b[349]), .Z(n1404) );
  NAND U1755 ( .A(a[348]), .B(b[348]), .Z(n1402) );
  NAND U1756 ( .A(n1400), .B(n1399), .Z(n1401) );
  NAND U1757 ( .A(n1402), .B(n1401), .Z(n1403) );
  XOR U1758 ( .A(n1404), .B(n1403), .Z(c[349]) );
  XOR U1759 ( .A(a[350]), .B(b[350]), .Z(n1408) );
  NAND U1760 ( .A(a[349]), .B(b[349]), .Z(n1406) );
  NAND U1761 ( .A(n1404), .B(n1403), .Z(n1405) );
  NAND U1762 ( .A(n1406), .B(n1405), .Z(n1407) );
  XOR U1763 ( .A(n1408), .B(n1407), .Z(c[350]) );
  XOR U1764 ( .A(a[351]), .B(b[351]), .Z(n1412) );
  NAND U1765 ( .A(a[350]), .B(b[350]), .Z(n1410) );
  NAND U1766 ( .A(n1408), .B(n1407), .Z(n1409) );
  NAND U1767 ( .A(n1410), .B(n1409), .Z(n1411) );
  XOR U1768 ( .A(n1412), .B(n1411), .Z(c[351]) );
  XOR U1769 ( .A(a[352]), .B(b[352]), .Z(n1416) );
  NAND U1770 ( .A(a[351]), .B(b[351]), .Z(n1414) );
  NAND U1771 ( .A(n1412), .B(n1411), .Z(n1413) );
  NAND U1772 ( .A(n1414), .B(n1413), .Z(n1415) );
  XOR U1773 ( .A(n1416), .B(n1415), .Z(c[352]) );
  XOR U1774 ( .A(a[353]), .B(b[353]), .Z(n1420) );
  NAND U1775 ( .A(a[352]), .B(b[352]), .Z(n1418) );
  NAND U1776 ( .A(n1416), .B(n1415), .Z(n1417) );
  NAND U1777 ( .A(n1418), .B(n1417), .Z(n1419) );
  XOR U1778 ( .A(n1420), .B(n1419), .Z(c[353]) );
  XOR U1779 ( .A(a[354]), .B(b[354]), .Z(n1424) );
  NAND U1780 ( .A(a[353]), .B(b[353]), .Z(n1422) );
  NAND U1781 ( .A(n1420), .B(n1419), .Z(n1421) );
  NAND U1782 ( .A(n1422), .B(n1421), .Z(n1423) );
  XOR U1783 ( .A(n1424), .B(n1423), .Z(c[354]) );
  XOR U1784 ( .A(a[355]), .B(b[355]), .Z(n1428) );
  NAND U1785 ( .A(a[354]), .B(b[354]), .Z(n1426) );
  NAND U1786 ( .A(n1424), .B(n1423), .Z(n1425) );
  NAND U1787 ( .A(n1426), .B(n1425), .Z(n1427) );
  XOR U1788 ( .A(n1428), .B(n1427), .Z(c[355]) );
  XOR U1789 ( .A(a[356]), .B(b[356]), .Z(n1432) );
  NAND U1790 ( .A(a[355]), .B(b[355]), .Z(n1430) );
  NAND U1791 ( .A(n1428), .B(n1427), .Z(n1429) );
  NAND U1792 ( .A(n1430), .B(n1429), .Z(n1431) );
  XOR U1793 ( .A(n1432), .B(n1431), .Z(c[356]) );
  XOR U1794 ( .A(a[357]), .B(b[357]), .Z(n1436) );
  NAND U1795 ( .A(a[356]), .B(b[356]), .Z(n1434) );
  NAND U1796 ( .A(n1432), .B(n1431), .Z(n1433) );
  NAND U1797 ( .A(n1434), .B(n1433), .Z(n1435) );
  XOR U1798 ( .A(n1436), .B(n1435), .Z(c[357]) );
  XOR U1799 ( .A(a[358]), .B(b[358]), .Z(n1440) );
  NAND U1800 ( .A(a[357]), .B(b[357]), .Z(n1438) );
  NAND U1801 ( .A(n1436), .B(n1435), .Z(n1437) );
  NAND U1802 ( .A(n1438), .B(n1437), .Z(n1439) );
  XOR U1803 ( .A(n1440), .B(n1439), .Z(c[358]) );
  XOR U1804 ( .A(a[359]), .B(b[359]), .Z(n1444) );
  NAND U1805 ( .A(a[358]), .B(b[358]), .Z(n1442) );
  NAND U1806 ( .A(n1440), .B(n1439), .Z(n1441) );
  NAND U1807 ( .A(n1442), .B(n1441), .Z(n1443) );
  XOR U1808 ( .A(n1444), .B(n1443), .Z(c[359]) );
  XOR U1809 ( .A(a[360]), .B(b[360]), .Z(n1448) );
  NAND U1810 ( .A(a[359]), .B(b[359]), .Z(n1446) );
  NAND U1811 ( .A(n1444), .B(n1443), .Z(n1445) );
  NAND U1812 ( .A(n1446), .B(n1445), .Z(n1447) );
  XOR U1813 ( .A(n1448), .B(n1447), .Z(c[360]) );
  XOR U1814 ( .A(a[361]), .B(b[361]), .Z(n1452) );
  NAND U1815 ( .A(a[360]), .B(b[360]), .Z(n1450) );
  NAND U1816 ( .A(n1448), .B(n1447), .Z(n1449) );
  NAND U1817 ( .A(n1450), .B(n1449), .Z(n1451) );
  XOR U1818 ( .A(n1452), .B(n1451), .Z(c[361]) );
  XOR U1819 ( .A(a[362]), .B(b[362]), .Z(n1456) );
  NAND U1820 ( .A(a[361]), .B(b[361]), .Z(n1454) );
  NAND U1821 ( .A(n1452), .B(n1451), .Z(n1453) );
  NAND U1822 ( .A(n1454), .B(n1453), .Z(n1455) );
  XOR U1823 ( .A(n1456), .B(n1455), .Z(c[362]) );
  XOR U1824 ( .A(a[363]), .B(b[363]), .Z(n1460) );
  NAND U1825 ( .A(a[362]), .B(b[362]), .Z(n1458) );
  NAND U1826 ( .A(n1456), .B(n1455), .Z(n1457) );
  NAND U1827 ( .A(n1458), .B(n1457), .Z(n1459) );
  XOR U1828 ( .A(n1460), .B(n1459), .Z(c[363]) );
  XOR U1829 ( .A(a[364]), .B(b[364]), .Z(n1464) );
  NAND U1830 ( .A(a[363]), .B(b[363]), .Z(n1462) );
  NAND U1831 ( .A(n1460), .B(n1459), .Z(n1461) );
  NAND U1832 ( .A(n1462), .B(n1461), .Z(n1463) );
  XOR U1833 ( .A(n1464), .B(n1463), .Z(c[364]) );
  XOR U1834 ( .A(a[365]), .B(b[365]), .Z(n1468) );
  NAND U1835 ( .A(a[364]), .B(b[364]), .Z(n1466) );
  NAND U1836 ( .A(n1464), .B(n1463), .Z(n1465) );
  NAND U1837 ( .A(n1466), .B(n1465), .Z(n1467) );
  XOR U1838 ( .A(n1468), .B(n1467), .Z(c[365]) );
  XOR U1839 ( .A(a[366]), .B(b[366]), .Z(n1472) );
  NAND U1840 ( .A(a[365]), .B(b[365]), .Z(n1470) );
  NAND U1841 ( .A(n1468), .B(n1467), .Z(n1469) );
  NAND U1842 ( .A(n1470), .B(n1469), .Z(n1471) );
  XOR U1843 ( .A(n1472), .B(n1471), .Z(c[366]) );
  XOR U1844 ( .A(a[367]), .B(b[367]), .Z(n1476) );
  NAND U1845 ( .A(a[366]), .B(b[366]), .Z(n1474) );
  NAND U1846 ( .A(n1472), .B(n1471), .Z(n1473) );
  NAND U1847 ( .A(n1474), .B(n1473), .Z(n1475) );
  XOR U1848 ( .A(n1476), .B(n1475), .Z(c[367]) );
  XOR U1849 ( .A(a[368]), .B(b[368]), .Z(n1480) );
  NAND U1850 ( .A(a[367]), .B(b[367]), .Z(n1478) );
  NAND U1851 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U1852 ( .A(n1478), .B(n1477), .Z(n1479) );
  XOR U1853 ( .A(n1480), .B(n1479), .Z(c[368]) );
  XOR U1854 ( .A(a[369]), .B(b[369]), .Z(n1484) );
  NAND U1855 ( .A(a[368]), .B(b[368]), .Z(n1482) );
  NAND U1856 ( .A(n1480), .B(n1479), .Z(n1481) );
  NAND U1857 ( .A(n1482), .B(n1481), .Z(n1483) );
  XOR U1858 ( .A(n1484), .B(n1483), .Z(c[369]) );
  XOR U1859 ( .A(a[370]), .B(b[370]), .Z(n1488) );
  NAND U1860 ( .A(a[369]), .B(b[369]), .Z(n1486) );
  NAND U1861 ( .A(n1484), .B(n1483), .Z(n1485) );
  NAND U1862 ( .A(n1486), .B(n1485), .Z(n1487) );
  XOR U1863 ( .A(n1488), .B(n1487), .Z(c[370]) );
  XOR U1864 ( .A(a[371]), .B(b[371]), .Z(n1492) );
  NAND U1865 ( .A(a[370]), .B(b[370]), .Z(n1490) );
  NAND U1866 ( .A(n1488), .B(n1487), .Z(n1489) );
  NAND U1867 ( .A(n1490), .B(n1489), .Z(n1491) );
  XOR U1868 ( .A(n1492), .B(n1491), .Z(c[371]) );
  XOR U1869 ( .A(a[372]), .B(b[372]), .Z(n1496) );
  NAND U1870 ( .A(a[371]), .B(b[371]), .Z(n1494) );
  NAND U1871 ( .A(n1492), .B(n1491), .Z(n1493) );
  NAND U1872 ( .A(n1494), .B(n1493), .Z(n1495) );
  XOR U1873 ( .A(n1496), .B(n1495), .Z(c[372]) );
  XOR U1874 ( .A(a[373]), .B(b[373]), .Z(n1500) );
  NAND U1875 ( .A(a[372]), .B(b[372]), .Z(n1498) );
  NAND U1876 ( .A(n1496), .B(n1495), .Z(n1497) );
  NAND U1877 ( .A(n1498), .B(n1497), .Z(n1499) );
  XOR U1878 ( .A(n1500), .B(n1499), .Z(c[373]) );
  XOR U1879 ( .A(a[374]), .B(b[374]), .Z(n1504) );
  NAND U1880 ( .A(a[373]), .B(b[373]), .Z(n1502) );
  NAND U1881 ( .A(n1500), .B(n1499), .Z(n1501) );
  NAND U1882 ( .A(n1502), .B(n1501), .Z(n1503) );
  XOR U1883 ( .A(n1504), .B(n1503), .Z(c[374]) );
  XOR U1884 ( .A(a[375]), .B(b[375]), .Z(n1508) );
  NAND U1885 ( .A(a[374]), .B(b[374]), .Z(n1506) );
  NAND U1886 ( .A(n1504), .B(n1503), .Z(n1505) );
  NAND U1887 ( .A(n1506), .B(n1505), .Z(n1507) );
  XOR U1888 ( .A(n1508), .B(n1507), .Z(c[375]) );
  XOR U1889 ( .A(a[376]), .B(b[376]), .Z(n1512) );
  NAND U1890 ( .A(a[375]), .B(b[375]), .Z(n1510) );
  NAND U1891 ( .A(n1508), .B(n1507), .Z(n1509) );
  NAND U1892 ( .A(n1510), .B(n1509), .Z(n1511) );
  XOR U1893 ( .A(n1512), .B(n1511), .Z(c[376]) );
  XOR U1894 ( .A(a[377]), .B(b[377]), .Z(n1516) );
  NAND U1895 ( .A(a[376]), .B(b[376]), .Z(n1514) );
  NAND U1896 ( .A(n1512), .B(n1511), .Z(n1513) );
  NAND U1897 ( .A(n1514), .B(n1513), .Z(n1515) );
  XOR U1898 ( .A(n1516), .B(n1515), .Z(c[377]) );
  XOR U1899 ( .A(a[378]), .B(b[378]), .Z(n1520) );
  NAND U1900 ( .A(a[377]), .B(b[377]), .Z(n1518) );
  NAND U1901 ( .A(n1516), .B(n1515), .Z(n1517) );
  NAND U1902 ( .A(n1518), .B(n1517), .Z(n1519) );
  XOR U1903 ( .A(n1520), .B(n1519), .Z(c[378]) );
  XOR U1904 ( .A(a[379]), .B(b[379]), .Z(n1524) );
  NAND U1905 ( .A(a[378]), .B(b[378]), .Z(n1522) );
  NAND U1906 ( .A(n1520), .B(n1519), .Z(n1521) );
  NAND U1907 ( .A(n1522), .B(n1521), .Z(n1523) );
  XOR U1908 ( .A(n1524), .B(n1523), .Z(c[379]) );
  XOR U1909 ( .A(a[380]), .B(b[380]), .Z(n1528) );
  NAND U1910 ( .A(a[379]), .B(b[379]), .Z(n1526) );
  NAND U1911 ( .A(n1524), .B(n1523), .Z(n1525) );
  NAND U1912 ( .A(n1526), .B(n1525), .Z(n1527) );
  XOR U1913 ( .A(n1528), .B(n1527), .Z(c[380]) );
  XOR U1914 ( .A(a[381]), .B(b[381]), .Z(n1532) );
  NAND U1915 ( .A(a[380]), .B(b[380]), .Z(n1530) );
  NAND U1916 ( .A(n1528), .B(n1527), .Z(n1529) );
  NAND U1917 ( .A(n1530), .B(n1529), .Z(n1531) );
  XOR U1918 ( .A(n1532), .B(n1531), .Z(c[381]) );
  XOR U1919 ( .A(a[382]), .B(b[382]), .Z(n1536) );
  NAND U1920 ( .A(a[381]), .B(b[381]), .Z(n1534) );
  NAND U1921 ( .A(n1532), .B(n1531), .Z(n1533) );
  NAND U1922 ( .A(n1534), .B(n1533), .Z(n1535) );
  XOR U1923 ( .A(n1536), .B(n1535), .Z(c[382]) );
  XOR U1924 ( .A(a[383]), .B(b[383]), .Z(n1540) );
  NAND U1925 ( .A(a[382]), .B(b[382]), .Z(n1538) );
  NAND U1926 ( .A(n1536), .B(n1535), .Z(n1537) );
  NAND U1927 ( .A(n1538), .B(n1537), .Z(n1539) );
  XOR U1928 ( .A(n1540), .B(n1539), .Z(c[383]) );
  XOR U1929 ( .A(a[384]), .B(b[384]), .Z(n1544) );
  NAND U1930 ( .A(a[383]), .B(b[383]), .Z(n1542) );
  NAND U1931 ( .A(n1540), .B(n1539), .Z(n1541) );
  NAND U1932 ( .A(n1542), .B(n1541), .Z(n1543) );
  XOR U1933 ( .A(n1544), .B(n1543), .Z(c[384]) );
  XOR U1934 ( .A(a[385]), .B(b[385]), .Z(n1548) );
  NAND U1935 ( .A(a[384]), .B(b[384]), .Z(n1546) );
  NAND U1936 ( .A(n1544), .B(n1543), .Z(n1545) );
  NAND U1937 ( .A(n1546), .B(n1545), .Z(n1547) );
  XOR U1938 ( .A(n1548), .B(n1547), .Z(c[385]) );
  XOR U1939 ( .A(b[386]), .B(a[386]), .Z(n1552) );
  NAND U1940 ( .A(a[385]), .B(b[385]), .Z(n1550) );
  NAND U1941 ( .A(n1548), .B(n1547), .Z(n1549) );
  AND U1942 ( .A(n1550), .B(n1549), .Z(n1551) );
  XNOR U1943 ( .A(n1552), .B(n1551), .Z(c[386]) );
  OR U1944 ( .A(b[386]), .B(a[386]), .Z(n1554) );
  NAND U1945 ( .A(n1552), .B(n1551), .Z(n1553) );
  AND U1946 ( .A(n1554), .B(n1553), .Z(n1556) );
  XOR U1947 ( .A(a[387]), .B(b[387]), .Z(n1555) );
  XOR U1948 ( .A(n1556), .B(n1555), .Z(c[387]) );
  XOR U1949 ( .A(a[388]), .B(b[388]), .Z(n1560) );
  NAND U1950 ( .A(a[387]), .B(b[387]), .Z(n1558) );
  NAND U1951 ( .A(n1556), .B(n1555), .Z(n1557) );
  NAND U1952 ( .A(n1558), .B(n1557), .Z(n1559) );
  XOR U1953 ( .A(n1560), .B(n1559), .Z(c[388]) );
  XOR U1954 ( .A(a[389]), .B(b[389]), .Z(n1564) );
  NAND U1955 ( .A(a[388]), .B(b[388]), .Z(n1562) );
  NAND U1956 ( .A(n1560), .B(n1559), .Z(n1561) );
  NAND U1957 ( .A(n1562), .B(n1561), .Z(n1563) );
  XOR U1958 ( .A(n1564), .B(n1563), .Z(c[389]) );
  XOR U1959 ( .A(a[390]), .B(b[390]), .Z(n1568) );
  NAND U1960 ( .A(a[389]), .B(b[389]), .Z(n1566) );
  NAND U1961 ( .A(n1564), .B(n1563), .Z(n1565) );
  NAND U1962 ( .A(n1566), .B(n1565), .Z(n1567) );
  XOR U1963 ( .A(n1568), .B(n1567), .Z(c[390]) );
  XOR U1964 ( .A(a[391]), .B(b[391]), .Z(n1572) );
  NAND U1965 ( .A(a[390]), .B(b[390]), .Z(n1570) );
  NAND U1966 ( .A(n1568), .B(n1567), .Z(n1569) );
  NAND U1967 ( .A(n1570), .B(n1569), .Z(n1571) );
  XOR U1968 ( .A(n1572), .B(n1571), .Z(c[391]) );
  XOR U1969 ( .A(a[392]), .B(b[392]), .Z(n1576) );
  NAND U1970 ( .A(a[391]), .B(b[391]), .Z(n1574) );
  NAND U1971 ( .A(n1572), .B(n1571), .Z(n1573) );
  NAND U1972 ( .A(n1574), .B(n1573), .Z(n1575) );
  XOR U1973 ( .A(n1576), .B(n1575), .Z(c[392]) );
  XOR U1974 ( .A(a[393]), .B(b[393]), .Z(n1580) );
  NAND U1975 ( .A(a[392]), .B(b[392]), .Z(n1578) );
  NAND U1976 ( .A(n1576), .B(n1575), .Z(n1577) );
  NAND U1977 ( .A(n1578), .B(n1577), .Z(n1579) );
  XOR U1978 ( .A(n1580), .B(n1579), .Z(c[393]) );
  XOR U1979 ( .A(a[394]), .B(b[394]), .Z(n1584) );
  NAND U1980 ( .A(a[393]), .B(b[393]), .Z(n1582) );
  NAND U1981 ( .A(n1580), .B(n1579), .Z(n1581) );
  NAND U1982 ( .A(n1582), .B(n1581), .Z(n1583) );
  XOR U1983 ( .A(n1584), .B(n1583), .Z(c[394]) );
  XOR U1984 ( .A(a[395]), .B(b[395]), .Z(n1588) );
  NAND U1985 ( .A(a[394]), .B(b[394]), .Z(n1586) );
  NAND U1986 ( .A(n1584), .B(n1583), .Z(n1585) );
  NAND U1987 ( .A(n1586), .B(n1585), .Z(n1587) );
  XOR U1988 ( .A(n1588), .B(n1587), .Z(c[395]) );
  XOR U1989 ( .A(a[396]), .B(b[396]), .Z(n1592) );
  NAND U1990 ( .A(a[395]), .B(b[395]), .Z(n1590) );
  NAND U1991 ( .A(n1588), .B(n1587), .Z(n1589) );
  NAND U1992 ( .A(n1590), .B(n1589), .Z(n1591) );
  XOR U1993 ( .A(n1592), .B(n1591), .Z(c[396]) );
  XOR U1994 ( .A(a[397]), .B(b[397]), .Z(n1596) );
  NAND U1995 ( .A(a[396]), .B(b[396]), .Z(n1594) );
  NAND U1996 ( .A(n1592), .B(n1591), .Z(n1593) );
  NAND U1997 ( .A(n1594), .B(n1593), .Z(n1595) );
  XOR U1998 ( .A(n1596), .B(n1595), .Z(c[397]) );
  XOR U1999 ( .A(a[398]), .B(b[398]), .Z(n1600) );
  NAND U2000 ( .A(a[397]), .B(b[397]), .Z(n1598) );
  NAND U2001 ( .A(n1596), .B(n1595), .Z(n1597) );
  NAND U2002 ( .A(n1598), .B(n1597), .Z(n1599) );
  XOR U2003 ( .A(n1600), .B(n1599), .Z(c[398]) );
  XOR U2004 ( .A(a[399]), .B(b[399]), .Z(n1604) );
  NAND U2005 ( .A(a[398]), .B(b[398]), .Z(n1602) );
  NAND U2006 ( .A(n1600), .B(n1599), .Z(n1601) );
  NAND U2007 ( .A(n1602), .B(n1601), .Z(n1603) );
  XOR U2008 ( .A(n1604), .B(n1603), .Z(c[399]) );
  XOR U2009 ( .A(a[400]), .B(b[400]), .Z(n1608) );
  NAND U2010 ( .A(a[399]), .B(b[399]), .Z(n1606) );
  NAND U2011 ( .A(n1604), .B(n1603), .Z(n1605) );
  NAND U2012 ( .A(n1606), .B(n1605), .Z(n1607) );
  XOR U2013 ( .A(n1608), .B(n1607), .Z(c[400]) );
  XOR U2014 ( .A(a[401]), .B(b[401]), .Z(n1612) );
  NAND U2015 ( .A(a[400]), .B(b[400]), .Z(n1610) );
  NAND U2016 ( .A(n1608), .B(n1607), .Z(n1609) );
  NAND U2017 ( .A(n1610), .B(n1609), .Z(n1611) );
  XOR U2018 ( .A(n1612), .B(n1611), .Z(c[401]) );
  XOR U2019 ( .A(a[402]), .B(b[402]), .Z(n1616) );
  NAND U2020 ( .A(a[401]), .B(b[401]), .Z(n1614) );
  NAND U2021 ( .A(n1612), .B(n1611), .Z(n1613) );
  NAND U2022 ( .A(n1614), .B(n1613), .Z(n1615) );
  XOR U2023 ( .A(n1616), .B(n1615), .Z(c[402]) );
  XOR U2024 ( .A(a[403]), .B(b[403]), .Z(n1620) );
  NAND U2025 ( .A(a[402]), .B(b[402]), .Z(n1618) );
  NAND U2026 ( .A(n1616), .B(n1615), .Z(n1617) );
  NAND U2027 ( .A(n1618), .B(n1617), .Z(n1619) );
  XOR U2028 ( .A(n1620), .B(n1619), .Z(c[403]) );
  XOR U2029 ( .A(a[404]), .B(b[404]), .Z(n1624) );
  NAND U2030 ( .A(a[403]), .B(b[403]), .Z(n1622) );
  NAND U2031 ( .A(n1620), .B(n1619), .Z(n1621) );
  NAND U2032 ( .A(n1622), .B(n1621), .Z(n1623) );
  XOR U2033 ( .A(n1624), .B(n1623), .Z(c[404]) );
  XOR U2034 ( .A(a[405]), .B(b[405]), .Z(n1628) );
  NAND U2035 ( .A(a[404]), .B(b[404]), .Z(n1626) );
  NAND U2036 ( .A(n1624), .B(n1623), .Z(n1625) );
  NAND U2037 ( .A(n1626), .B(n1625), .Z(n1627) );
  XOR U2038 ( .A(n1628), .B(n1627), .Z(c[405]) );
  XOR U2039 ( .A(a[406]), .B(b[406]), .Z(n1632) );
  NAND U2040 ( .A(a[405]), .B(b[405]), .Z(n1630) );
  NAND U2041 ( .A(n1628), .B(n1627), .Z(n1629) );
  NAND U2042 ( .A(n1630), .B(n1629), .Z(n1631) );
  XOR U2043 ( .A(n1632), .B(n1631), .Z(c[406]) );
  XOR U2044 ( .A(a[407]), .B(b[407]), .Z(n1636) );
  NAND U2045 ( .A(a[406]), .B(b[406]), .Z(n1634) );
  NAND U2046 ( .A(n1632), .B(n1631), .Z(n1633) );
  NAND U2047 ( .A(n1634), .B(n1633), .Z(n1635) );
  XOR U2048 ( .A(n1636), .B(n1635), .Z(c[407]) );
  XOR U2049 ( .A(b[408]), .B(a[408]), .Z(n1640) );
  NAND U2050 ( .A(a[407]), .B(b[407]), .Z(n1638) );
  NAND U2051 ( .A(n1636), .B(n1635), .Z(n1637) );
  AND U2052 ( .A(n1638), .B(n1637), .Z(n1639) );
  XNOR U2053 ( .A(n1640), .B(n1639), .Z(c[408]) );
  XOR U2054 ( .A(a[409]), .B(b[409]), .Z(n1644) );
  OR U2055 ( .A(b[408]), .B(a[408]), .Z(n1642) );
  NAND U2056 ( .A(n1640), .B(n1639), .Z(n1641) );
  AND U2057 ( .A(n1642), .B(n1641), .Z(n1643) );
  XOR U2058 ( .A(n1644), .B(n1643), .Z(c[409]) );
  XOR U2059 ( .A(a[410]), .B(b[410]), .Z(n1648) );
  NAND U2060 ( .A(a[409]), .B(b[409]), .Z(n1646) );
  NAND U2061 ( .A(n1644), .B(n1643), .Z(n1645) );
  NAND U2062 ( .A(n1646), .B(n1645), .Z(n1647) );
  XOR U2063 ( .A(n1648), .B(n1647), .Z(c[410]) );
  XOR U2064 ( .A(b[411]), .B(a[411]), .Z(n1652) );
  NAND U2065 ( .A(a[410]), .B(b[410]), .Z(n1650) );
  NAND U2066 ( .A(n1648), .B(n1647), .Z(n1649) );
  AND U2067 ( .A(n1650), .B(n1649), .Z(n1651) );
  XNOR U2068 ( .A(n1652), .B(n1651), .Z(c[411]) );
  OR U2069 ( .A(b[411]), .B(a[411]), .Z(n1654) );
  NAND U2070 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U2071 ( .A(n1654), .B(n1653), .Z(n1656) );
  XOR U2072 ( .A(a[412]), .B(b[412]), .Z(n1655) );
  XOR U2073 ( .A(n1656), .B(n1655), .Z(c[412]) );
  XOR U2074 ( .A(a[413]), .B(b[413]), .Z(n1660) );
  NAND U2075 ( .A(a[412]), .B(b[412]), .Z(n1658) );
  NAND U2076 ( .A(n1656), .B(n1655), .Z(n1657) );
  NAND U2077 ( .A(n1658), .B(n1657), .Z(n1659) );
  XOR U2078 ( .A(n1660), .B(n1659), .Z(c[413]) );
  XOR U2079 ( .A(a[414]), .B(b[414]), .Z(n1664) );
  NAND U2080 ( .A(a[413]), .B(b[413]), .Z(n1662) );
  NAND U2081 ( .A(n1660), .B(n1659), .Z(n1661) );
  NAND U2082 ( .A(n1662), .B(n1661), .Z(n1663) );
  XOR U2083 ( .A(n1664), .B(n1663), .Z(c[414]) );
  XOR U2084 ( .A(a[415]), .B(b[415]), .Z(n1668) );
  NAND U2085 ( .A(a[414]), .B(b[414]), .Z(n1666) );
  NAND U2086 ( .A(n1664), .B(n1663), .Z(n1665) );
  NAND U2087 ( .A(n1666), .B(n1665), .Z(n1667) );
  XOR U2088 ( .A(n1668), .B(n1667), .Z(c[415]) );
  XOR U2089 ( .A(a[416]), .B(b[416]), .Z(n1672) );
  NAND U2090 ( .A(a[415]), .B(b[415]), .Z(n1670) );
  NAND U2091 ( .A(n1668), .B(n1667), .Z(n1669) );
  NAND U2092 ( .A(n1670), .B(n1669), .Z(n1671) );
  XOR U2093 ( .A(n1672), .B(n1671), .Z(c[416]) );
  XOR U2094 ( .A(a[417]), .B(b[417]), .Z(n1676) );
  NAND U2095 ( .A(a[416]), .B(b[416]), .Z(n1674) );
  NAND U2096 ( .A(n1672), .B(n1671), .Z(n1673) );
  NAND U2097 ( .A(n1674), .B(n1673), .Z(n1675) );
  XOR U2098 ( .A(n1676), .B(n1675), .Z(c[417]) );
  XOR U2099 ( .A(a[418]), .B(b[418]), .Z(n1680) );
  NAND U2100 ( .A(a[417]), .B(b[417]), .Z(n1678) );
  NAND U2101 ( .A(n1676), .B(n1675), .Z(n1677) );
  NAND U2102 ( .A(n1678), .B(n1677), .Z(n1679) );
  XOR U2103 ( .A(n1680), .B(n1679), .Z(c[418]) );
  XOR U2104 ( .A(a[419]), .B(b[419]), .Z(n1684) );
  NAND U2105 ( .A(a[418]), .B(b[418]), .Z(n1682) );
  NAND U2106 ( .A(n1680), .B(n1679), .Z(n1681) );
  NAND U2107 ( .A(n1682), .B(n1681), .Z(n1683) );
  XOR U2108 ( .A(n1684), .B(n1683), .Z(c[419]) );
  XOR U2109 ( .A(a[420]), .B(b[420]), .Z(n1688) );
  NAND U2110 ( .A(a[419]), .B(b[419]), .Z(n1686) );
  NAND U2111 ( .A(n1684), .B(n1683), .Z(n1685) );
  NAND U2112 ( .A(n1686), .B(n1685), .Z(n1687) );
  XOR U2113 ( .A(n1688), .B(n1687), .Z(c[420]) );
  XOR U2114 ( .A(a[421]), .B(b[421]), .Z(n1692) );
  NAND U2115 ( .A(a[420]), .B(b[420]), .Z(n1690) );
  NAND U2116 ( .A(n1688), .B(n1687), .Z(n1689) );
  NAND U2117 ( .A(n1690), .B(n1689), .Z(n1691) );
  XOR U2118 ( .A(n1692), .B(n1691), .Z(c[421]) );
  XOR U2119 ( .A(a[422]), .B(b[422]), .Z(n1696) );
  NAND U2120 ( .A(a[421]), .B(b[421]), .Z(n1694) );
  NAND U2121 ( .A(n1692), .B(n1691), .Z(n1693) );
  NAND U2122 ( .A(n1694), .B(n1693), .Z(n1695) );
  XOR U2123 ( .A(n1696), .B(n1695), .Z(c[422]) );
  XOR U2124 ( .A(a[423]), .B(b[423]), .Z(n1700) );
  NAND U2125 ( .A(a[422]), .B(b[422]), .Z(n1698) );
  NAND U2126 ( .A(n1696), .B(n1695), .Z(n1697) );
  NAND U2127 ( .A(n1698), .B(n1697), .Z(n1699) );
  XOR U2128 ( .A(n1700), .B(n1699), .Z(c[423]) );
  XOR U2129 ( .A(a[424]), .B(b[424]), .Z(n1704) );
  NAND U2130 ( .A(a[423]), .B(b[423]), .Z(n1702) );
  NAND U2131 ( .A(n1700), .B(n1699), .Z(n1701) );
  NAND U2132 ( .A(n1702), .B(n1701), .Z(n1703) );
  XOR U2133 ( .A(n1704), .B(n1703), .Z(c[424]) );
  XOR U2134 ( .A(a[425]), .B(b[425]), .Z(n1708) );
  NAND U2135 ( .A(a[424]), .B(b[424]), .Z(n1706) );
  NAND U2136 ( .A(n1704), .B(n1703), .Z(n1705) );
  NAND U2137 ( .A(n1706), .B(n1705), .Z(n1707) );
  XOR U2138 ( .A(n1708), .B(n1707), .Z(c[425]) );
  XOR U2139 ( .A(a[426]), .B(b[426]), .Z(n1712) );
  NAND U2140 ( .A(a[425]), .B(b[425]), .Z(n1710) );
  NAND U2141 ( .A(n1708), .B(n1707), .Z(n1709) );
  NAND U2142 ( .A(n1710), .B(n1709), .Z(n1711) );
  XOR U2143 ( .A(n1712), .B(n1711), .Z(c[426]) );
  XOR U2144 ( .A(a[427]), .B(b[427]), .Z(n1716) );
  NAND U2145 ( .A(a[426]), .B(b[426]), .Z(n1714) );
  NAND U2146 ( .A(n1712), .B(n1711), .Z(n1713) );
  NAND U2147 ( .A(n1714), .B(n1713), .Z(n1715) );
  XOR U2148 ( .A(n1716), .B(n1715), .Z(c[427]) );
  XOR U2149 ( .A(a[428]), .B(b[428]), .Z(n1720) );
  NAND U2150 ( .A(a[427]), .B(b[427]), .Z(n1718) );
  NAND U2151 ( .A(n1716), .B(n1715), .Z(n1717) );
  NAND U2152 ( .A(n1718), .B(n1717), .Z(n1719) );
  XOR U2153 ( .A(n1720), .B(n1719), .Z(c[428]) );
  XOR U2154 ( .A(a[429]), .B(b[429]), .Z(n1724) );
  NAND U2155 ( .A(a[428]), .B(b[428]), .Z(n1722) );
  NAND U2156 ( .A(n1720), .B(n1719), .Z(n1721) );
  NAND U2157 ( .A(n1722), .B(n1721), .Z(n1723) );
  XOR U2158 ( .A(n1724), .B(n1723), .Z(c[429]) );
  XOR U2159 ( .A(a[430]), .B(b[430]), .Z(n1728) );
  NAND U2160 ( .A(a[429]), .B(b[429]), .Z(n1726) );
  NAND U2161 ( .A(n1724), .B(n1723), .Z(n1725) );
  NAND U2162 ( .A(n1726), .B(n1725), .Z(n1727) );
  XOR U2163 ( .A(n1728), .B(n1727), .Z(c[430]) );
  XOR U2164 ( .A(a[431]), .B(b[431]), .Z(n1732) );
  NAND U2165 ( .A(a[430]), .B(b[430]), .Z(n1730) );
  NAND U2166 ( .A(n1728), .B(n1727), .Z(n1729) );
  NAND U2167 ( .A(n1730), .B(n1729), .Z(n1731) );
  XOR U2168 ( .A(n1732), .B(n1731), .Z(c[431]) );
  XOR U2169 ( .A(a[432]), .B(b[432]), .Z(n1736) );
  NAND U2170 ( .A(a[431]), .B(b[431]), .Z(n1734) );
  NAND U2171 ( .A(n1732), .B(n1731), .Z(n1733) );
  NAND U2172 ( .A(n1734), .B(n1733), .Z(n1735) );
  XOR U2173 ( .A(n1736), .B(n1735), .Z(c[432]) );
  XOR U2174 ( .A(a[433]), .B(b[433]), .Z(n1740) );
  NAND U2175 ( .A(a[432]), .B(b[432]), .Z(n1738) );
  NAND U2176 ( .A(n1736), .B(n1735), .Z(n1737) );
  NAND U2177 ( .A(n1738), .B(n1737), .Z(n1739) );
  XOR U2178 ( .A(n1740), .B(n1739), .Z(c[433]) );
  XOR U2179 ( .A(a[434]), .B(b[434]), .Z(n1744) );
  NAND U2180 ( .A(a[433]), .B(b[433]), .Z(n1742) );
  NAND U2181 ( .A(n1740), .B(n1739), .Z(n1741) );
  NAND U2182 ( .A(n1742), .B(n1741), .Z(n1743) );
  XOR U2183 ( .A(n1744), .B(n1743), .Z(c[434]) );
  XOR U2184 ( .A(a[435]), .B(b[435]), .Z(n1748) );
  NAND U2185 ( .A(a[434]), .B(b[434]), .Z(n1746) );
  NAND U2186 ( .A(n1744), .B(n1743), .Z(n1745) );
  NAND U2187 ( .A(n1746), .B(n1745), .Z(n1747) );
  XOR U2188 ( .A(n1748), .B(n1747), .Z(c[435]) );
  XOR U2189 ( .A(a[436]), .B(b[436]), .Z(n1752) );
  NAND U2190 ( .A(a[435]), .B(b[435]), .Z(n1750) );
  NAND U2191 ( .A(n1748), .B(n1747), .Z(n1749) );
  NAND U2192 ( .A(n1750), .B(n1749), .Z(n1751) );
  XOR U2193 ( .A(n1752), .B(n1751), .Z(c[436]) );
  XOR U2194 ( .A(a[437]), .B(b[437]), .Z(n1756) );
  NAND U2195 ( .A(a[436]), .B(b[436]), .Z(n1754) );
  NAND U2196 ( .A(n1752), .B(n1751), .Z(n1753) );
  NAND U2197 ( .A(n1754), .B(n1753), .Z(n1755) );
  XOR U2198 ( .A(n1756), .B(n1755), .Z(c[437]) );
  XOR U2199 ( .A(a[438]), .B(b[438]), .Z(n1760) );
  NAND U2200 ( .A(a[437]), .B(b[437]), .Z(n1758) );
  NAND U2201 ( .A(n1756), .B(n1755), .Z(n1757) );
  NAND U2202 ( .A(n1758), .B(n1757), .Z(n1759) );
  XOR U2203 ( .A(n1760), .B(n1759), .Z(c[438]) );
  XOR U2204 ( .A(a[439]), .B(b[439]), .Z(n1764) );
  NAND U2205 ( .A(a[438]), .B(b[438]), .Z(n1762) );
  NAND U2206 ( .A(n1760), .B(n1759), .Z(n1761) );
  NAND U2207 ( .A(n1762), .B(n1761), .Z(n1763) );
  XOR U2208 ( .A(n1764), .B(n1763), .Z(c[439]) );
  XOR U2209 ( .A(a[440]), .B(b[440]), .Z(n1768) );
  NAND U2210 ( .A(a[439]), .B(b[439]), .Z(n1766) );
  NAND U2211 ( .A(n1764), .B(n1763), .Z(n1765) );
  NAND U2212 ( .A(n1766), .B(n1765), .Z(n1767) );
  XOR U2213 ( .A(n1768), .B(n1767), .Z(c[440]) );
  XOR U2214 ( .A(a[441]), .B(b[441]), .Z(n1772) );
  NAND U2215 ( .A(a[440]), .B(b[440]), .Z(n1770) );
  NAND U2216 ( .A(n1768), .B(n1767), .Z(n1769) );
  NAND U2217 ( .A(n1770), .B(n1769), .Z(n1771) );
  XOR U2218 ( .A(n1772), .B(n1771), .Z(c[441]) );
  XOR U2219 ( .A(a[442]), .B(b[442]), .Z(n1776) );
  NAND U2220 ( .A(a[441]), .B(b[441]), .Z(n1774) );
  NAND U2221 ( .A(n1772), .B(n1771), .Z(n1773) );
  NAND U2222 ( .A(n1774), .B(n1773), .Z(n1775) );
  XOR U2223 ( .A(n1776), .B(n1775), .Z(c[442]) );
  NAND U2224 ( .A(a[442]), .B(b[442]), .Z(n1778) );
  NAND U2225 ( .A(n1776), .B(n1775), .Z(n1777) );
  AND U2226 ( .A(n1778), .B(n1777), .Z(n1780) );
  XOR U2227 ( .A(b[443]), .B(a[443]), .Z(n1779) );
  XNOR U2228 ( .A(n1780), .B(n1779), .Z(c[443]) );
  OR U2229 ( .A(b[443]), .B(a[443]), .Z(n1782) );
  NAND U2230 ( .A(n1780), .B(n1779), .Z(n1781) );
  AND U2231 ( .A(n1782), .B(n1781), .Z(n1784) );
  XOR U2232 ( .A(a[444]), .B(b[444]), .Z(n1783) );
  XOR U2233 ( .A(n1784), .B(n1783), .Z(c[444]) );
  XOR U2234 ( .A(a[445]), .B(b[445]), .Z(n1788) );
  NAND U2235 ( .A(a[444]), .B(b[444]), .Z(n1786) );
  NAND U2236 ( .A(n1784), .B(n1783), .Z(n1785) );
  NAND U2237 ( .A(n1786), .B(n1785), .Z(n1787) );
  XOR U2238 ( .A(n1788), .B(n1787), .Z(c[445]) );
  XOR U2239 ( .A(b[446]), .B(a[446]), .Z(n1792) );
  NAND U2240 ( .A(a[445]), .B(b[445]), .Z(n1790) );
  NAND U2241 ( .A(n1788), .B(n1787), .Z(n1789) );
  AND U2242 ( .A(n1790), .B(n1789), .Z(n1791) );
  XNOR U2243 ( .A(n1792), .B(n1791), .Z(c[446]) );
  OR U2244 ( .A(b[446]), .B(a[446]), .Z(n1794) );
  NAND U2245 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U2246 ( .A(n1794), .B(n1793), .Z(n1796) );
  XOR U2247 ( .A(a[447]), .B(b[447]), .Z(n1795) );
  XOR U2248 ( .A(n1796), .B(n1795), .Z(c[447]) );
  XOR U2249 ( .A(a[448]), .B(b[448]), .Z(n1800) );
  NAND U2250 ( .A(a[447]), .B(b[447]), .Z(n1798) );
  NAND U2251 ( .A(n1796), .B(n1795), .Z(n1797) );
  NAND U2252 ( .A(n1798), .B(n1797), .Z(n1799) );
  XOR U2253 ( .A(n1800), .B(n1799), .Z(c[448]) );
  NAND U2254 ( .A(a[448]), .B(b[448]), .Z(n1802) );
  NAND U2255 ( .A(n1800), .B(n1799), .Z(n1801) );
  AND U2256 ( .A(n1802), .B(n1801), .Z(n1804) );
  XOR U2257 ( .A(b[449]), .B(a[449]), .Z(n1803) );
  XNOR U2258 ( .A(n1804), .B(n1803), .Z(c[449]) );
  OR U2259 ( .A(b[449]), .B(a[449]), .Z(n1806) );
  NAND U2260 ( .A(n1804), .B(n1803), .Z(n1805) );
  AND U2261 ( .A(n1806), .B(n1805), .Z(n1808) );
  XOR U2262 ( .A(a[450]), .B(b[450]), .Z(n1807) );
  XOR U2263 ( .A(n1808), .B(n1807), .Z(c[450]) );
  XOR U2264 ( .A(a[451]), .B(b[451]), .Z(n1812) );
  NAND U2265 ( .A(a[450]), .B(b[450]), .Z(n1810) );
  NAND U2266 ( .A(n1808), .B(n1807), .Z(n1809) );
  NAND U2267 ( .A(n1810), .B(n1809), .Z(n1811) );
  XOR U2268 ( .A(n1812), .B(n1811), .Z(c[451]) );
  XOR U2269 ( .A(b[452]), .B(a[452]), .Z(n1816) );
  NAND U2270 ( .A(a[451]), .B(b[451]), .Z(n1814) );
  NAND U2271 ( .A(n1812), .B(n1811), .Z(n1813) );
  AND U2272 ( .A(n1814), .B(n1813), .Z(n1815) );
  XNOR U2273 ( .A(n1816), .B(n1815), .Z(c[452]) );
  OR U2274 ( .A(b[452]), .B(a[452]), .Z(n1818) );
  NAND U2275 ( .A(n1816), .B(n1815), .Z(n1817) );
  AND U2276 ( .A(n1818), .B(n1817), .Z(n1820) );
  XOR U2277 ( .A(a[453]), .B(b[453]), .Z(n1819) );
  XOR U2278 ( .A(n1820), .B(n1819), .Z(c[453]) );
  XOR U2279 ( .A(a[454]), .B(b[454]), .Z(n1824) );
  NAND U2280 ( .A(a[453]), .B(b[453]), .Z(n1822) );
  NAND U2281 ( .A(n1820), .B(n1819), .Z(n1821) );
  NAND U2282 ( .A(n1822), .B(n1821), .Z(n1823) );
  XOR U2283 ( .A(n1824), .B(n1823), .Z(c[454]) );
  XOR U2284 ( .A(a[455]), .B(b[455]), .Z(n1828) );
  NAND U2285 ( .A(a[454]), .B(b[454]), .Z(n1826) );
  NAND U2286 ( .A(n1824), .B(n1823), .Z(n1825) );
  NAND U2287 ( .A(n1826), .B(n1825), .Z(n1827) );
  XOR U2288 ( .A(n1828), .B(n1827), .Z(c[455]) );
  XOR U2289 ( .A(a[456]), .B(b[456]), .Z(n1832) );
  NAND U2290 ( .A(a[455]), .B(b[455]), .Z(n1830) );
  NAND U2291 ( .A(n1828), .B(n1827), .Z(n1829) );
  NAND U2292 ( .A(n1830), .B(n1829), .Z(n1831) );
  XOR U2293 ( .A(n1832), .B(n1831), .Z(c[456]) );
  XOR U2294 ( .A(a[457]), .B(b[457]), .Z(n1836) );
  NAND U2295 ( .A(a[456]), .B(b[456]), .Z(n1834) );
  NAND U2296 ( .A(n1832), .B(n1831), .Z(n1833) );
  NAND U2297 ( .A(n1834), .B(n1833), .Z(n1835) );
  XOR U2298 ( .A(n1836), .B(n1835), .Z(c[457]) );
  XOR U2299 ( .A(a[458]), .B(b[458]), .Z(n1840) );
  NAND U2300 ( .A(a[457]), .B(b[457]), .Z(n1838) );
  NAND U2301 ( .A(n1836), .B(n1835), .Z(n1837) );
  NAND U2302 ( .A(n1838), .B(n1837), .Z(n1839) );
  XOR U2303 ( .A(n1840), .B(n1839), .Z(c[458]) );
  XOR U2304 ( .A(a[459]), .B(b[459]), .Z(n1844) );
  NAND U2305 ( .A(a[458]), .B(b[458]), .Z(n1842) );
  NAND U2306 ( .A(n1840), .B(n1839), .Z(n1841) );
  NAND U2307 ( .A(n1842), .B(n1841), .Z(n1843) );
  XOR U2308 ( .A(n1844), .B(n1843), .Z(c[459]) );
  NAND U2309 ( .A(a[459]), .B(b[459]), .Z(n1846) );
  NAND U2310 ( .A(n1844), .B(n1843), .Z(n1845) );
  AND U2311 ( .A(n1846), .B(n1845), .Z(n1848) );
  XOR U2312 ( .A(b[460]), .B(a[460]), .Z(n1847) );
  XNOR U2313 ( .A(n1848), .B(n1847), .Z(c[460]) );
  XOR U2314 ( .A(a[461]), .B(b[461]), .Z(n1852) );
  OR U2315 ( .A(b[460]), .B(a[460]), .Z(n1850) );
  NAND U2316 ( .A(n1848), .B(n1847), .Z(n1849) );
  AND U2317 ( .A(n1850), .B(n1849), .Z(n1851) );
  XOR U2318 ( .A(n1852), .B(n1851), .Z(c[461]) );
  XOR U2319 ( .A(a[462]), .B(b[462]), .Z(n1856) );
  NAND U2320 ( .A(a[461]), .B(b[461]), .Z(n1854) );
  NAND U2321 ( .A(n1852), .B(n1851), .Z(n1853) );
  NAND U2322 ( .A(n1854), .B(n1853), .Z(n1855) );
  XOR U2323 ( .A(n1856), .B(n1855), .Z(c[462]) );
  XOR U2324 ( .A(a[463]), .B(b[463]), .Z(n1860) );
  NAND U2325 ( .A(a[462]), .B(b[462]), .Z(n1858) );
  NAND U2326 ( .A(n1856), .B(n1855), .Z(n1857) );
  NAND U2327 ( .A(n1858), .B(n1857), .Z(n1859) );
  XOR U2328 ( .A(n1860), .B(n1859), .Z(c[463]) );
  XOR U2329 ( .A(a[464]), .B(b[464]), .Z(n1864) );
  NAND U2330 ( .A(a[463]), .B(b[463]), .Z(n1862) );
  NAND U2331 ( .A(n1860), .B(n1859), .Z(n1861) );
  NAND U2332 ( .A(n1862), .B(n1861), .Z(n1863) );
  XOR U2333 ( .A(n1864), .B(n1863), .Z(c[464]) );
  XOR U2334 ( .A(a[465]), .B(b[465]), .Z(n1868) );
  NAND U2335 ( .A(a[464]), .B(b[464]), .Z(n1866) );
  NAND U2336 ( .A(n1864), .B(n1863), .Z(n1865) );
  NAND U2337 ( .A(n1866), .B(n1865), .Z(n1867) );
  XOR U2338 ( .A(n1868), .B(n1867), .Z(c[465]) );
  XOR U2339 ( .A(a[466]), .B(b[466]), .Z(n1872) );
  NAND U2340 ( .A(a[465]), .B(b[465]), .Z(n1870) );
  NAND U2341 ( .A(n1868), .B(n1867), .Z(n1869) );
  NAND U2342 ( .A(n1870), .B(n1869), .Z(n1871) );
  XOR U2343 ( .A(n1872), .B(n1871), .Z(c[466]) );
  XOR U2344 ( .A(a[467]), .B(b[467]), .Z(n1876) );
  NAND U2345 ( .A(a[466]), .B(b[466]), .Z(n1874) );
  NAND U2346 ( .A(n1872), .B(n1871), .Z(n1873) );
  NAND U2347 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U2348 ( .A(n1876), .B(n1875), .Z(c[467]) );
  XOR U2349 ( .A(a[468]), .B(b[468]), .Z(n1880) );
  NAND U2350 ( .A(a[467]), .B(b[467]), .Z(n1878) );
  NAND U2351 ( .A(n1876), .B(n1875), .Z(n1877) );
  NAND U2352 ( .A(n1878), .B(n1877), .Z(n1879) );
  XOR U2353 ( .A(n1880), .B(n1879), .Z(c[468]) );
  XOR U2354 ( .A(a[469]), .B(b[469]), .Z(n1884) );
  NAND U2355 ( .A(a[468]), .B(b[468]), .Z(n1882) );
  NAND U2356 ( .A(n1880), .B(n1879), .Z(n1881) );
  NAND U2357 ( .A(n1882), .B(n1881), .Z(n1883) );
  XOR U2358 ( .A(n1884), .B(n1883), .Z(c[469]) );
  XOR U2359 ( .A(a[470]), .B(b[470]), .Z(n1888) );
  NAND U2360 ( .A(a[469]), .B(b[469]), .Z(n1886) );
  NAND U2361 ( .A(n1884), .B(n1883), .Z(n1885) );
  NAND U2362 ( .A(n1886), .B(n1885), .Z(n1887) );
  XOR U2363 ( .A(n1888), .B(n1887), .Z(c[470]) );
  XOR U2364 ( .A(a[471]), .B(b[471]), .Z(n1892) );
  NAND U2365 ( .A(a[470]), .B(b[470]), .Z(n1890) );
  NAND U2366 ( .A(n1888), .B(n1887), .Z(n1889) );
  NAND U2367 ( .A(n1890), .B(n1889), .Z(n1891) );
  XOR U2368 ( .A(n1892), .B(n1891), .Z(c[471]) );
  XOR U2369 ( .A(a[472]), .B(b[472]), .Z(n1896) );
  NAND U2370 ( .A(a[471]), .B(b[471]), .Z(n1894) );
  NAND U2371 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U2372 ( .A(n1894), .B(n1893), .Z(n1895) );
  XOR U2373 ( .A(n1896), .B(n1895), .Z(c[472]) );
  XOR U2374 ( .A(a[473]), .B(b[473]), .Z(n1900) );
  NAND U2375 ( .A(a[472]), .B(b[472]), .Z(n1898) );
  NAND U2376 ( .A(n1896), .B(n1895), .Z(n1897) );
  NAND U2377 ( .A(n1898), .B(n1897), .Z(n1899) );
  XOR U2378 ( .A(n1900), .B(n1899), .Z(c[473]) );
  XOR U2379 ( .A(a[474]), .B(b[474]), .Z(n1904) );
  NAND U2380 ( .A(a[473]), .B(b[473]), .Z(n1902) );
  NAND U2381 ( .A(n1900), .B(n1899), .Z(n1901) );
  NAND U2382 ( .A(n1902), .B(n1901), .Z(n1903) );
  XOR U2383 ( .A(n1904), .B(n1903), .Z(c[474]) );
  XOR U2384 ( .A(a[475]), .B(b[475]), .Z(n1908) );
  NAND U2385 ( .A(a[474]), .B(b[474]), .Z(n1906) );
  NAND U2386 ( .A(n1904), .B(n1903), .Z(n1905) );
  NAND U2387 ( .A(n1906), .B(n1905), .Z(n1907) );
  XOR U2388 ( .A(n1908), .B(n1907), .Z(c[475]) );
  XOR U2389 ( .A(a[476]), .B(b[476]), .Z(n1912) );
  NAND U2390 ( .A(a[475]), .B(b[475]), .Z(n1910) );
  NAND U2391 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U2392 ( .A(n1910), .B(n1909), .Z(n1911) );
  XOR U2393 ( .A(n1912), .B(n1911), .Z(c[476]) );
  XOR U2394 ( .A(a[477]), .B(b[477]), .Z(n1916) );
  NAND U2395 ( .A(a[476]), .B(b[476]), .Z(n1914) );
  NAND U2396 ( .A(n1912), .B(n1911), .Z(n1913) );
  NAND U2397 ( .A(n1914), .B(n1913), .Z(n1915) );
  XOR U2398 ( .A(n1916), .B(n1915), .Z(c[477]) );
  XOR U2399 ( .A(a[478]), .B(b[478]), .Z(n1920) );
  NAND U2400 ( .A(a[477]), .B(b[477]), .Z(n1918) );
  NAND U2401 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U2402 ( .A(n1918), .B(n1917), .Z(n1919) );
  XOR U2403 ( .A(n1920), .B(n1919), .Z(c[478]) );
  XOR U2404 ( .A(a[479]), .B(b[479]), .Z(n1924) );
  NAND U2405 ( .A(a[478]), .B(b[478]), .Z(n1922) );
  NAND U2406 ( .A(n1920), .B(n1919), .Z(n1921) );
  NAND U2407 ( .A(n1922), .B(n1921), .Z(n1923) );
  XOR U2408 ( .A(n1924), .B(n1923), .Z(c[479]) );
  XOR U2409 ( .A(a[480]), .B(b[480]), .Z(n1928) );
  NAND U2410 ( .A(a[479]), .B(b[479]), .Z(n1926) );
  NAND U2411 ( .A(n1924), .B(n1923), .Z(n1925) );
  NAND U2412 ( .A(n1926), .B(n1925), .Z(n1927) );
  XOR U2413 ( .A(n1928), .B(n1927), .Z(c[480]) );
  XOR U2414 ( .A(a[481]), .B(b[481]), .Z(n1932) );
  NAND U2415 ( .A(a[480]), .B(b[480]), .Z(n1930) );
  NAND U2416 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U2417 ( .A(n1930), .B(n1929), .Z(n1931) );
  XOR U2418 ( .A(n1932), .B(n1931), .Z(c[481]) );
  XOR U2419 ( .A(a[482]), .B(b[482]), .Z(n1936) );
  NAND U2420 ( .A(a[481]), .B(b[481]), .Z(n1934) );
  NAND U2421 ( .A(n1932), .B(n1931), .Z(n1933) );
  NAND U2422 ( .A(n1934), .B(n1933), .Z(n1935) );
  XOR U2423 ( .A(n1936), .B(n1935), .Z(c[482]) );
  XOR U2424 ( .A(a[483]), .B(b[483]), .Z(n1940) );
  NAND U2425 ( .A(a[482]), .B(b[482]), .Z(n1938) );
  NAND U2426 ( .A(n1936), .B(n1935), .Z(n1937) );
  NAND U2427 ( .A(n1938), .B(n1937), .Z(n1939) );
  XOR U2428 ( .A(n1940), .B(n1939), .Z(c[483]) );
  XOR U2429 ( .A(a[484]), .B(b[484]), .Z(n1944) );
  NAND U2430 ( .A(a[483]), .B(b[483]), .Z(n1942) );
  NAND U2431 ( .A(n1940), .B(n1939), .Z(n1941) );
  NAND U2432 ( .A(n1942), .B(n1941), .Z(n1943) );
  XOR U2433 ( .A(n1944), .B(n1943), .Z(c[484]) );
  XOR U2434 ( .A(a[485]), .B(b[485]), .Z(n1948) );
  NAND U2435 ( .A(a[484]), .B(b[484]), .Z(n1946) );
  NAND U2436 ( .A(n1944), .B(n1943), .Z(n1945) );
  NAND U2437 ( .A(n1946), .B(n1945), .Z(n1947) );
  XOR U2438 ( .A(n1948), .B(n1947), .Z(c[485]) );
  XOR U2439 ( .A(a[486]), .B(b[486]), .Z(n1952) );
  NAND U2440 ( .A(a[485]), .B(b[485]), .Z(n1950) );
  NAND U2441 ( .A(n1948), .B(n1947), .Z(n1949) );
  NAND U2442 ( .A(n1950), .B(n1949), .Z(n1951) );
  XOR U2443 ( .A(n1952), .B(n1951), .Z(c[486]) );
  XOR U2444 ( .A(a[487]), .B(b[487]), .Z(n1956) );
  NAND U2445 ( .A(a[486]), .B(b[486]), .Z(n1954) );
  NAND U2446 ( .A(n1952), .B(n1951), .Z(n1953) );
  NAND U2447 ( .A(n1954), .B(n1953), .Z(n1955) );
  XOR U2448 ( .A(n1956), .B(n1955), .Z(c[487]) );
  XOR U2449 ( .A(a[488]), .B(b[488]), .Z(n1960) );
  NAND U2450 ( .A(a[487]), .B(b[487]), .Z(n1958) );
  NAND U2451 ( .A(n1956), .B(n1955), .Z(n1957) );
  NAND U2452 ( .A(n1958), .B(n1957), .Z(n1959) );
  XOR U2453 ( .A(n1960), .B(n1959), .Z(c[488]) );
  XOR U2454 ( .A(a[489]), .B(b[489]), .Z(n1964) );
  NAND U2455 ( .A(a[488]), .B(b[488]), .Z(n1962) );
  NAND U2456 ( .A(n1960), .B(n1959), .Z(n1961) );
  NAND U2457 ( .A(n1962), .B(n1961), .Z(n1963) );
  XOR U2458 ( .A(n1964), .B(n1963), .Z(c[489]) );
  XOR U2459 ( .A(a[490]), .B(b[490]), .Z(n1968) );
  NAND U2460 ( .A(a[489]), .B(b[489]), .Z(n1966) );
  NAND U2461 ( .A(n1964), .B(n1963), .Z(n1965) );
  NAND U2462 ( .A(n1966), .B(n1965), .Z(n1967) );
  XOR U2463 ( .A(n1968), .B(n1967), .Z(c[490]) );
  XOR U2464 ( .A(a[491]), .B(b[491]), .Z(n1972) );
  NAND U2465 ( .A(a[490]), .B(b[490]), .Z(n1970) );
  NAND U2466 ( .A(n1968), .B(n1967), .Z(n1969) );
  NAND U2467 ( .A(n1970), .B(n1969), .Z(n1971) );
  XOR U2468 ( .A(n1972), .B(n1971), .Z(c[491]) );
  XOR U2469 ( .A(a[492]), .B(b[492]), .Z(n1976) );
  NAND U2470 ( .A(a[491]), .B(b[491]), .Z(n1974) );
  NAND U2471 ( .A(n1972), .B(n1971), .Z(n1973) );
  NAND U2472 ( .A(n1974), .B(n1973), .Z(n1975) );
  XOR U2473 ( .A(n1976), .B(n1975), .Z(c[492]) );
  XOR U2474 ( .A(a[493]), .B(b[493]), .Z(n1980) );
  NAND U2475 ( .A(a[492]), .B(b[492]), .Z(n1978) );
  NAND U2476 ( .A(n1976), .B(n1975), .Z(n1977) );
  NAND U2477 ( .A(n1978), .B(n1977), .Z(n1979) );
  XOR U2478 ( .A(n1980), .B(n1979), .Z(c[493]) );
  XOR U2479 ( .A(a[494]), .B(b[494]), .Z(n1984) );
  NAND U2480 ( .A(a[493]), .B(b[493]), .Z(n1982) );
  NAND U2481 ( .A(n1980), .B(n1979), .Z(n1981) );
  NAND U2482 ( .A(n1982), .B(n1981), .Z(n1983) );
  XOR U2483 ( .A(n1984), .B(n1983), .Z(c[494]) );
  XOR U2484 ( .A(a[495]), .B(b[495]), .Z(n1988) );
  NAND U2485 ( .A(a[494]), .B(b[494]), .Z(n1986) );
  NAND U2486 ( .A(n1984), .B(n1983), .Z(n1985) );
  NAND U2487 ( .A(n1986), .B(n1985), .Z(n1987) );
  XOR U2488 ( .A(n1988), .B(n1987), .Z(c[495]) );
  XOR U2489 ( .A(a[496]), .B(b[496]), .Z(n1992) );
  NAND U2490 ( .A(a[495]), .B(b[495]), .Z(n1990) );
  NAND U2491 ( .A(n1988), .B(n1987), .Z(n1989) );
  NAND U2492 ( .A(n1990), .B(n1989), .Z(n1991) );
  XOR U2493 ( .A(n1992), .B(n1991), .Z(c[496]) );
  XOR U2494 ( .A(a[497]), .B(b[497]), .Z(n1996) );
  NAND U2495 ( .A(a[496]), .B(b[496]), .Z(n1994) );
  NAND U2496 ( .A(n1992), .B(n1991), .Z(n1993) );
  NAND U2497 ( .A(n1994), .B(n1993), .Z(n1995) );
  XOR U2498 ( .A(n1996), .B(n1995), .Z(c[497]) );
  XOR U2499 ( .A(a[498]), .B(b[498]), .Z(n2000) );
  NAND U2500 ( .A(a[497]), .B(b[497]), .Z(n1998) );
  NAND U2501 ( .A(n1996), .B(n1995), .Z(n1997) );
  NAND U2502 ( .A(n1998), .B(n1997), .Z(n1999) );
  XOR U2503 ( .A(n2000), .B(n1999), .Z(c[498]) );
  XOR U2504 ( .A(a[499]), .B(b[499]), .Z(n2004) );
  NAND U2505 ( .A(a[498]), .B(b[498]), .Z(n2002) );
  NAND U2506 ( .A(n2000), .B(n1999), .Z(n2001) );
  NAND U2507 ( .A(n2002), .B(n2001), .Z(n2003) );
  XOR U2508 ( .A(n2004), .B(n2003), .Z(c[499]) );
  XOR U2509 ( .A(a[500]), .B(b[500]), .Z(n2008) );
  NAND U2510 ( .A(a[499]), .B(b[499]), .Z(n2006) );
  NAND U2511 ( .A(n2004), .B(n2003), .Z(n2005) );
  NAND U2512 ( .A(n2006), .B(n2005), .Z(n2007) );
  XOR U2513 ( .A(n2008), .B(n2007), .Z(c[500]) );
  XOR U2514 ( .A(a[501]), .B(b[501]), .Z(n2012) );
  NAND U2515 ( .A(a[500]), .B(b[500]), .Z(n2010) );
  NAND U2516 ( .A(n2008), .B(n2007), .Z(n2009) );
  NAND U2517 ( .A(n2010), .B(n2009), .Z(n2011) );
  XOR U2518 ( .A(n2012), .B(n2011), .Z(c[501]) );
  NAND U2519 ( .A(a[501]), .B(b[501]), .Z(n2014) );
  NAND U2520 ( .A(n2012), .B(n2011), .Z(n2013) );
  NAND U2521 ( .A(n2014), .B(n2013), .Z(n2016) );
  XNOR U2522 ( .A(b[502]), .B(a[502]), .Z(n2015) );
  XNOR U2523 ( .A(n2016), .B(n2015), .Z(c[502]) );
  XOR U2524 ( .A(a[503]), .B(b[503]), .Z(n2017) );
  XOR U2525 ( .A(n2018), .B(n2017), .Z(c[503]) );
  XOR U2526 ( .A(a[504]), .B(b[504]), .Z(n2022) );
  NAND U2527 ( .A(a[503]), .B(b[503]), .Z(n2020) );
  NAND U2528 ( .A(n2018), .B(n2017), .Z(n2019) );
  NAND U2529 ( .A(n2020), .B(n2019), .Z(n2021) );
  XOR U2530 ( .A(n2022), .B(n2021), .Z(c[504]) );
  XOR U2531 ( .A(a[505]), .B(b[505]), .Z(n2026) );
  NAND U2532 ( .A(a[504]), .B(b[504]), .Z(n2024) );
  NAND U2533 ( .A(n2022), .B(n2021), .Z(n2023) );
  NAND U2534 ( .A(n2024), .B(n2023), .Z(n2025) );
  XOR U2535 ( .A(n2026), .B(n2025), .Z(c[505]) );
  XOR U2536 ( .A(a[506]), .B(b[506]), .Z(n2030) );
  NAND U2537 ( .A(a[505]), .B(b[505]), .Z(n2028) );
  NAND U2538 ( .A(n2026), .B(n2025), .Z(n2027) );
  NAND U2539 ( .A(n2028), .B(n2027), .Z(n2029) );
  XOR U2540 ( .A(n2030), .B(n2029), .Z(c[506]) );
  XOR U2541 ( .A(a[507]), .B(b[507]), .Z(n2034) );
  NAND U2542 ( .A(a[506]), .B(b[506]), .Z(n2032) );
  NAND U2543 ( .A(n2030), .B(n2029), .Z(n2031) );
  NAND U2544 ( .A(n2032), .B(n2031), .Z(n2033) );
  XOR U2545 ( .A(n2034), .B(n2033), .Z(c[507]) );
  XOR U2546 ( .A(a[508]), .B(b[508]), .Z(n2038) );
  NAND U2547 ( .A(a[507]), .B(b[507]), .Z(n2036) );
  NAND U2548 ( .A(n2034), .B(n2033), .Z(n2035) );
  NAND U2549 ( .A(n2036), .B(n2035), .Z(n2037) );
  XOR U2550 ( .A(n2038), .B(n2037), .Z(c[508]) );
  XOR U2551 ( .A(a[509]), .B(b[509]), .Z(n2042) );
  NAND U2552 ( .A(a[508]), .B(b[508]), .Z(n2040) );
  NAND U2553 ( .A(n2038), .B(n2037), .Z(n2039) );
  NAND U2554 ( .A(n2040), .B(n2039), .Z(n2041) );
  XOR U2555 ( .A(n2042), .B(n2041), .Z(c[509]) );
  XOR U2556 ( .A(a[510]), .B(b[510]), .Z(n2046) );
  NAND U2557 ( .A(a[509]), .B(b[509]), .Z(n2044) );
  NAND U2558 ( .A(n2042), .B(n2041), .Z(n2043) );
  NAND U2559 ( .A(n2044), .B(n2043), .Z(n2045) );
  XOR U2560 ( .A(n2046), .B(n2045), .Z(c[510]) );
  NAND U2561 ( .A(a[510]), .B(b[510]), .Z(n2048) );
  NAND U2562 ( .A(n2046), .B(n2045), .Z(n2047) );
  NAND U2563 ( .A(n2048), .B(n2047), .Z(n2050) );
  XNOR U2564 ( .A(a[511]), .B(b[511]), .Z(n2049) );
  XNOR U2565 ( .A(n2050), .B(n2049), .Z(c[511]) );
endmodule

