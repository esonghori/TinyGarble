
module mult_N8_CC8 ( clk, rst, a, b, c );
  input [7:0] a;
  input [0:0] b;
  output [15:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;
  wire   [15:0] sreg;

  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(sreg[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(sreg[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(sreg[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(sreg[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(sreg[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(sreg[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(sreg[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(sreg[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U4 ( .A(n40), .B(sreg[8]), .Z(n1) );
  NANDN U5 ( .A(n42), .B(n1), .Z(n2) );
  NAND U6 ( .A(n40), .B(sreg[8]), .Z(n3) );
  AND U7 ( .A(n2), .B(n3), .Z(n21) );
  XOR U8 ( .A(sreg[11]), .B(n26), .Z(n4) );
  NANDN U9 ( .A(n27), .B(n4), .Z(n5) );
  NAND U10 ( .A(sreg[11]), .B(n26), .Z(n6) );
  AND U11 ( .A(n5), .B(n6), .Z(n30) );
  XOR U12 ( .A(sreg[9]), .B(n20), .Z(n7) );
  NANDN U13 ( .A(n21), .B(n7), .Z(n8) );
  NAND U14 ( .A(sreg[9]), .B(n20), .Z(n9) );
  AND U15 ( .A(n8), .B(n9), .Z(n24) );
  XOR U16 ( .A(sreg[12]), .B(n29), .Z(n10) );
  NANDN U17 ( .A(n30), .B(n10), .Z(n11) );
  NAND U18 ( .A(sreg[12]), .B(n29), .Z(n12) );
  AND U19 ( .A(n11), .B(n12), .Z(n33) );
  XOR U20 ( .A(sreg[10]), .B(n23), .Z(n13) );
  NANDN U21 ( .A(n24), .B(n13), .Z(n14) );
  NAND U22 ( .A(sreg[10]), .B(n23), .Z(n15) );
  AND U23 ( .A(n14), .B(n15), .Z(n27) );
  XOR U24 ( .A(sreg[13]), .B(n32), .Z(n16) );
  NANDN U25 ( .A(n33), .B(n16), .Z(n17) );
  NAND U26 ( .A(sreg[13]), .B(n32), .Z(n18) );
  AND U27 ( .A(n17), .B(n18), .Z(n36) );
  AND U28 ( .A(b[0]), .B(a[2]), .Z(n20) );
  AND U29 ( .A(b[0]), .B(a[0]), .Z(n39) );
  AND U30 ( .A(n39), .B(sreg[7]), .Z(n40) );
  NAND U31 ( .A(b[0]), .B(a[1]), .Z(n42) );
  XNOR U32 ( .A(n21), .B(sreg[9]), .Z(n19) );
  XOR U33 ( .A(n20), .B(n19), .Z(c[9]) );
  AND U34 ( .A(b[0]), .B(a[3]), .Z(n23) );
  XNOR U35 ( .A(n24), .B(sreg[10]), .Z(n22) );
  XOR U36 ( .A(n23), .B(n22), .Z(c[10]) );
  AND U37 ( .A(b[0]), .B(a[4]), .Z(n26) );
  XNOR U38 ( .A(n27), .B(sreg[11]), .Z(n25) );
  XOR U39 ( .A(n26), .B(n25), .Z(c[11]) );
  AND U40 ( .A(b[0]), .B(a[5]), .Z(n29) );
  XNOR U41 ( .A(n30), .B(sreg[12]), .Z(n28) );
  XOR U42 ( .A(n29), .B(n28), .Z(c[12]) );
  AND U43 ( .A(b[0]), .B(a[6]), .Z(n32) );
  XNOR U44 ( .A(n33), .B(sreg[13]), .Z(n31) );
  XOR U45 ( .A(n32), .B(n31), .Z(c[13]) );
  NAND U46 ( .A(b[0]), .B(a[7]), .Z(n34) );
  XNOR U47 ( .A(sreg[14]), .B(n36), .Z(n35) );
  XNOR U48 ( .A(n34), .B(n35), .Z(c[14]) );
  NAND U49 ( .A(n35), .B(n34), .Z(n38) );
  NANDN U50 ( .A(sreg[14]), .B(n36), .Z(n37) );
  AND U51 ( .A(n38), .B(n37), .Z(c[15]) );
  XOR U52 ( .A(n39), .B(sreg[7]), .Z(c[7]) );
  XOR U53 ( .A(sreg[8]), .B(n40), .Z(n41) );
  XNOR U54 ( .A(n42), .B(n41), .Z(c[8]) );
endmodule

