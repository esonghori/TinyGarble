
module Inst_Mem ( inst_mem_in_wire, pc, opcode );
  input [2047:0] inst_mem_in_wire;
  input [31:2] pc;
  output [31:0] opcode;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984;

  MUX U1 ( .IN0(inst_mem_in_wire[1984]), .IN1(inst_mem_in_wire[2016]), .SEL(
        pc[2]), .F(n1) );
  MUX U2 ( .IN0(inst_mem_in_wire[1920]), .IN1(inst_mem_in_wire[1952]), .SEL(
        pc[2]), .F(n2) );
  MUX U3 ( .IN0(n2), .IN1(n1), .SEL(pc[3]), .F(n3) );
  MUX U4 ( .IN0(inst_mem_in_wire[1856]), .IN1(inst_mem_in_wire[1888]), .SEL(
        pc[2]), .F(n4) );
  MUX U5 ( .IN0(inst_mem_in_wire[1792]), .IN1(inst_mem_in_wire[1824]), .SEL(
        pc[2]), .F(n5) );
  MUX U6 ( .IN0(n5), .IN1(n4), .SEL(pc[3]), .F(n6) );
  MUX U7 ( .IN0(n6), .IN1(n3), .SEL(pc[4]), .F(n7) );
  MUX U8 ( .IN0(inst_mem_in_wire[1728]), .IN1(inst_mem_in_wire[1760]), .SEL(
        pc[2]), .F(n8) );
  MUX U9 ( .IN0(inst_mem_in_wire[1664]), .IN1(inst_mem_in_wire[1696]), .SEL(
        pc[2]), .F(n9) );
  MUX U10 ( .IN0(n9), .IN1(n8), .SEL(pc[3]), .F(n10) );
  MUX U11 ( .IN0(inst_mem_in_wire[1600]), .IN1(inst_mem_in_wire[1632]), .SEL(
        pc[2]), .F(n11) );
  MUX U12 ( .IN0(inst_mem_in_wire[1536]), .IN1(inst_mem_in_wire[1568]), .SEL(
        pc[2]), .F(n12) );
  MUX U13 ( .IN0(n12), .IN1(n11), .SEL(pc[3]), .F(n13) );
  MUX U14 ( .IN0(n13), .IN1(n10), .SEL(pc[4]), .F(n14) );
  MUX U15 ( .IN0(n14), .IN1(n7), .SEL(pc[5]), .F(n15) );
  MUX U16 ( .IN0(inst_mem_in_wire[1472]), .IN1(inst_mem_in_wire[1504]), .SEL(
        pc[2]), .F(n16) );
  MUX U17 ( .IN0(inst_mem_in_wire[1408]), .IN1(inst_mem_in_wire[1440]), .SEL(
        pc[2]), .F(n17) );
  MUX U18 ( .IN0(n17), .IN1(n16), .SEL(pc[3]), .F(n18) );
  MUX U19 ( .IN0(inst_mem_in_wire[1344]), .IN1(inst_mem_in_wire[1376]), .SEL(
        pc[2]), .F(n19) );
  MUX U20 ( .IN0(inst_mem_in_wire[1280]), .IN1(inst_mem_in_wire[1312]), .SEL(
        pc[2]), .F(n20) );
  MUX U21 ( .IN0(n20), .IN1(n19), .SEL(pc[3]), .F(n21) );
  MUX U22 ( .IN0(n21), .IN1(n18), .SEL(pc[4]), .F(n22) );
  MUX U23 ( .IN0(inst_mem_in_wire[1216]), .IN1(inst_mem_in_wire[1248]), .SEL(
        pc[2]), .F(n23) );
  MUX U24 ( .IN0(inst_mem_in_wire[1152]), .IN1(inst_mem_in_wire[1184]), .SEL(
        pc[2]), .F(n24) );
  MUX U25 ( .IN0(n24), .IN1(n23), .SEL(pc[3]), .F(n25) );
  MUX U26 ( .IN0(inst_mem_in_wire[1088]), .IN1(inst_mem_in_wire[1120]), .SEL(
        pc[2]), .F(n26) );
  MUX U27 ( .IN0(inst_mem_in_wire[1024]), .IN1(inst_mem_in_wire[1056]), .SEL(
        pc[2]), .F(n27) );
  MUX U28 ( .IN0(n27), .IN1(n26), .SEL(pc[3]), .F(n28) );
  MUX U29 ( .IN0(n28), .IN1(n25), .SEL(pc[4]), .F(n29) );
  MUX U30 ( .IN0(n29), .IN1(n22), .SEL(pc[5]), .F(n30) );
  MUX U31 ( .IN0(n30), .IN1(n15), .SEL(pc[6]), .F(n31) );
  MUX U32 ( .IN0(inst_mem_in_wire[960]), .IN1(inst_mem_in_wire[992]), .SEL(
        pc[2]), .F(n32) );
  MUX U33 ( .IN0(inst_mem_in_wire[896]), .IN1(inst_mem_in_wire[928]), .SEL(
        pc[2]), .F(n33) );
  MUX U34 ( .IN0(n33), .IN1(n32), .SEL(pc[3]), .F(n34) );
  MUX U35 ( .IN0(inst_mem_in_wire[832]), .IN1(inst_mem_in_wire[864]), .SEL(
        pc[2]), .F(n35) );
  MUX U36 ( .IN0(inst_mem_in_wire[768]), .IN1(inst_mem_in_wire[800]), .SEL(
        pc[2]), .F(n36) );
  MUX U37 ( .IN0(n36), .IN1(n35), .SEL(pc[3]), .F(n37) );
  MUX U38 ( .IN0(n37), .IN1(n34), .SEL(pc[4]), .F(n38) );
  MUX U39 ( .IN0(inst_mem_in_wire[704]), .IN1(inst_mem_in_wire[736]), .SEL(
        pc[2]), .F(n39) );
  MUX U40 ( .IN0(inst_mem_in_wire[640]), .IN1(inst_mem_in_wire[672]), .SEL(
        pc[2]), .F(n40) );
  MUX U41 ( .IN0(n40), .IN1(n39), .SEL(pc[3]), .F(n41) );
  MUX U42 ( .IN0(inst_mem_in_wire[576]), .IN1(inst_mem_in_wire[608]), .SEL(
        pc[2]), .F(n42) );
  MUX U43 ( .IN0(inst_mem_in_wire[512]), .IN1(inst_mem_in_wire[544]), .SEL(
        pc[2]), .F(n43) );
  MUX U44 ( .IN0(n43), .IN1(n42), .SEL(pc[3]), .F(n44) );
  MUX U45 ( .IN0(n44), .IN1(n41), .SEL(pc[4]), .F(n45) );
  MUX U46 ( .IN0(n45), .IN1(n38), .SEL(pc[5]), .F(n46) );
  MUX U47 ( .IN0(inst_mem_in_wire[448]), .IN1(inst_mem_in_wire[480]), .SEL(
        pc[2]), .F(n47) );
  MUX U48 ( .IN0(inst_mem_in_wire[384]), .IN1(inst_mem_in_wire[416]), .SEL(
        pc[2]), .F(n48) );
  MUX U49 ( .IN0(n48), .IN1(n47), .SEL(pc[3]), .F(n49) );
  MUX U50 ( .IN0(inst_mem_in_wire[320]), .IN1(inst_mem_in_wire[352]), .SEL(
        pc[2]), .F(n50) );
  MUX U51 ( .IN0(inst_mem_in_wire[256]), .IN1(inst_mem_in_wire[288]), .SEL(
        pc[2]), .F(n51) );
  MUX U52 ( .IN0(n51), .IN1(n50), .SEL(pc[3]), .F(n52) );
  MUX U53 ( .IN0(n52), .IN1(n49), .SEL(pc[4]), .F(n53) );
  MUX U54 ( .IN0(inst_mem_in_wire[192]), .IN1(inst_mem_in_wire[224]), .SEL(
        pc[2]), .F(n54) );
  MUX U55 ( .IN0(inst_mem_in_wire[128]), .IN1(inst_mem_in_wire[160]), .SEL(
        pc[2]), .F(n55) );
  MUX U56 ( .IN0(n55), .IN1(n54), .SEL(pc[3]), .F(n56) );
  MUX U57 ( .IN0(inst_mem_in_wire[64]), .IN1(inst_mem_in_wire[96]), .SEL(pc[2]), .F(n57) );
  MUX U58 ( .IN0(inst_mem_in_wire[0]), .IN1(inst_mem_in_wire[32]), .SEL(pc[2]), 
        .F(n58) );
  MUX U59 ( .IN0(n58), .IN1(n57), .SEL(pc[3]), .F(n59) );
  MUX U60 ( .IN0(n59), .IN1(n56), .SEL(pc[4]), .F(n60) );
  MUX U61 ( .IN0(n60), .IN1(n53), .SEL(pc[5]), .F(n61) );
  MUX U62 ( .IN0(n61), .IN1(n46), .SEL(pc[6]), .F(n62) );
  MUX U63 ( .IN0(n62), .IN1(n31), .SEL(pc[7]), .F(opcode[0]) );
  MUX U64 ( .IN0(inst_mem_in_wire[1985]), .IN1(inst_mem_in_wire[2017]), .SEL(
        pc[2]), .F(n63) );
  MUX U65 ( .IN0(inst_mem_in_wire[1921]), .IN1(inst_mem_in_wire[1953]), .SEL(
        pc[2]), .F(n64) );
  MUX U66 ( .IN0(n64), .IN1(n63), .SEL(pc[3]), .F(n65) );
  MUX U67 ( .IN0(inst_mem_in_wire[1857]), .IN1(inst_mem_in_wire[1889]), .SEL(
        pc[2]), .F(n66) );
  MUX U68 ( .IN0(inst_mem_in_wire[1793]), .IN1(inst_mem_in_wire[1825]), .SEL(
        pc[2]), .F(n67) );
  MUX U69 ( .IN0(n67), .IN1(n66), .SEL(pc[3]), .F(n68) );
  MUX U70 ( .IN0(n68), .IN1(n65), .SEL(pc[4]), .F(n69) );
  MUX U71 ( .IN0(inst_mem_in_wire[1729]), .IN1(inst_mem_in_wire[1761]), .SEL(
        pc[2]), .F(n70) );
  MUX U72 ( .IN0(inst_mem_in_wire[1665]), .IN1(inst_mem_in_wire[1697]), .SEL(
        pc[2]), .F(n71) );
  MUX U73 ( .IN0(n71), .IN1(n70), .SEL(pc[3]), .F(n72) );
  MUX U74 ( .IN0(inst_mem_in_wire[1601]), .IN1(inst_mem_in_wire[1633]), .SEL(
        pc[2]), .F(n73) );
  MUX U75 ( .IN0(inst_mem_in_wire[1537]), .IN1(inst_mem_in_wire[1569]), .SEL(
        pc[2]), .F(n74) );
  MUX U76 ( .IN0(n74), .IN1(n73), .SEL(pc[3]), .F(n75) );
  MUX U77 ( .IN0(n75), .IN1(n72), .SEL(pc[4]), .F(n76) );
  MUX U78 ( .IN0(n76), .IN1(n69), .SEL(pc[5]), .F(n77) );
  MUX U79 ( .IN0(inst_mem_in_wire[1473]), .IN1(inst_mem_in_wire[1505]), .SEL(
        pc[2]), .F(n78) );
  MUX U80 ( .IN0(inst_mem_in_wire[1409]), .IN1(inst_mem_in_wire[1441]), .SEL(
        pc[2]), .F(n79) );
  MUX U81 ( .IN0(n79), .IN1(n78), .SEL(pc[3]), .F(n80) );
  MUX U82 ( .IN0(inst_mem_in_wire[1345]), .IN1(inst_mem_in_wire[1377]), .SEL(
        pc[2]), .F(n81) );
  MUX U83 ( .IN0(inst_mem_in_wire[1281]), .IN1(inst_mem_in_wire[1313]), .SEL(
        pc[2]), .F(n82) );
  MUX U84 ( .IN0(n82), .IN1(n81), .SEL(pc[3]), .F(n83) );
  MUX U85 ( .IN0(n83), .IN1(n80), .SEL(pc[4]), .F(n84) );
  MUX U86 ( .IN0(inst_mem_in_wire[1217]), .IN1(inst_mem_in_wire[1249]), .SEL(
        pc[2]), .F(n85) );
  MUX U87 ( .IN0(inst_mem_in_wire[1153]), .IN1(inst_mem_in_wire[1185]), .SEL(
        pc[2]), .F(n86) );
  MUX U88 ( .IN0(n86), .IN1(n85), .SEL(pc[3]), .F(n87) );
  MUX U89 ( .IN0(inst_mem_in_wire[1089]), .IN1(inst_mem_in_wire[1121]), .SEL(
        pc[2]), .F(n88) );
  MUX U90 ( .IN0(inst_mem_in_wire[1025]), .IN1(inst_mem_in_wire[1057]), .SEL(
        pc[2]), .F(n89) );
  MUX U91 ( .IN0(n89), .IN1(n88), .SEL(pc[3]), .F(n90) );
  MUX U92 ( .IN0(n90), .IN1(n87), .SEL(pc[4]), .F(n91) );
  MUX U93 ( .IN0(n91), .IN1(n84), .SEL(pc[5]), .F(n92) );
  MUX U94 ( .IN0(n92), .IN1(n77), .SEL(pc[6]), .F(n93) );
  MUX U95 ( .IN0(inst_mem_in_wire[961]), .IN1(inst_mem_in_wire[993]), .SEL(
        pc[2]), .F(n94) );
  MUX U96 ( .IN0(inst_mem_in_wire[897]), .IN1(inst_mem_in_wire[929]), .SEL(
        pc[2]), .F(n95) );
  MUX U97 ( .IN0(n95), .IN1(n94), .SEL(pc[3]), .F(n96) );
  MUX U98 ( .IN0(inst_mem_in_wire[833]), .IN1(inst_mem_in_wire[865]), .SEL(
        pc[2]), .F(n97) );
  MUX U99 ( .IN0(inst_mem_in_wire[769]), .IN1(inst_mem_in_wire[801]), .SEL(
        pc[2]), .F(n98) );
  MUX U100 ( .IN0(n98), .IN1(n97), .SEL(pc[3]), .F(n99) );
  MUX U101 ( .IN0(n99), .IN1(n96), .SEL(pc[4]), .F(n100) );
  MUX U102 ( .IN0(inst_mem_in_wire[705]), .IN1(inst_mem_in_wire[737]), .SEL(
        pc[2]), .F(n101) );
  MUX U103 ( .IN0(inst_mem_in_wire[641]), .IN1(inst_mem_in_wire[673]), .SEL(
        pc[2]), .F(n102) );
  MUX U104 ( .IN0(n102), .IN1(n101), .SEL(pc[3]), .F(n103) );
  MUX U105 ( .IN0(inst_mem_in_wire[577]), .IN1(inst_mem_in_wire[609]), .SEL(
        pc[2]), .F(n104) );
  MUX U106 ( .IN0(inst_mem_in_wire[513]), .IN1(inst_mem_in_wire[545]), .SEL(
        pc[2]), .F(n105) );
  MUX U107 ( .IN0(n105), .IN1(n104), .SEL(pc[3]), .F(n106) );
  MUX U108 ( .IN0(n106), .IN1(n103), .SEL(pc[4]), .F(n107) );
  MUX U109 ( .IN0(n107), .IN1(n100), .SEL(pc[5]), .F(n108) );
  MUX U110 ( .IN0(inst_mem_in_wire[449]), .IN1(inst_mem_in_wire[481]), .SEL(
        pc[2]), .F(n109) );
  MUX U111 ( .IN0(inst_mem_in_wire[385]), .IN1(inst_mem_in_wire[417]), .SEL(
        pc[2]), .F(n110) );
  MUX U112 ( .IN0(n110), .IN1(n109), .SEL(pc[3]), .F(n111) );
  MUX U113 ( .IN0(inst_mem_in_wire[321]), .IN1(inst_mem_in_wire[353]), .SEL(
        pc[2]), .F(n112) );
  MUX U114 ( .IN0(inst_mem_in_wire[257]), .IN1(inst_mem_in_wire[289]), .SEL(
        pc[2]), .F(n113) );
  MUX U115 ( .IN0(n113), .IN1(n112), .SEL(pc[3]), .F(n114) );
  MUX U116 ( .IN0(n114), .IN1(n111), .SEL(pc[4]), .F(n115) );
  MUX U117 ( .IN0(inst_mem_in_wire[193]), .IN1(inst_mem_in_wire[225]), .SEL(
        pc[2]), .F(n116) );
  MUX U118 ( .IN0(inst_mem_in_wire[129]), .IN1(inst_mem_in_wire[161]), .SEL(
        pc[2]), .F(n117) );
  MUX U119 ( .IN0(n117), .IN1(n116), .SEL(pc[3]), .F(n118) );
  MUX U120 ( .IN0(inst_mem_in_wire[65]), .IN1(inst_mem_in_wire[97]), .SEL(
        pc[2]), .F(n119) );
  MUX U121 ( .IN0(inst_mem_in_wire[1]), .IN1(inst_mem_in_wire[33]), .SEL(pc[2]), .F(n120) );
  MUX U122 ( .IN0(n120), .IN1(n119), .SEL(pc[3]), .F(n121) );
  MUX U123 ( .IN0(n121), .IN1(n118), .SEL(pc[4]), .F(n122) );
  MUX U124 ( .IN0(n122), .IN1(n115), .SEL(pc[5]), .F(n123) );
  MUX U125 ( .IN0(n123), .IN1(n108), .SEL(pc[6]), .F(n124) );
  MUX U126 ( .IN0(n124), .IN1(n93), .SEL(pc[7]), .F(opcode[1]) );
  MUX U127 ( .IN0(inst_mem_in_wire[1986]), .IN1(inst_mem_in_wire[2018]), .SEL(
        pc[2]), .F(n125) );
  MUX U128 ( .IN0(inst_mem_in_wire[1922]), .IN1(inst_mem_in_wire[1954]), .SEL(
        pc[2]), .F(n126) );
  MUX U129 ( .IN0(n126), .IN1(n125), .SEL(pc[3]), .F(n127) );
  MUX U130 ( .IN0(inst_mem_in_wire[1858]), .IN1(inst_mem_in_wire[1890]), .SEL(
        pc[2]), .F(n128) );
  MUX U131 ( .IN0(inst_mem_in_wire[1794]), .IN1(inst_mem_in_wire[1826]), .SEL(
        pc[2]), .F(n129) );
  MUX U132 ( .IN0(n129), .IN1(n128), .SEL(pc[3]), .F(n130) );
  MUX U133 ( .IN0(n130), .IN1(n127), .SEL(pc[4]), .F(n131) );
  MUX U134 ( .IN0(inst_mem_in_wire[1730]), .IN1(inst_mem_in_wire[1762]), .SEL(
        pc[2]), .F(n132) );
  MUX U135 ( .IN0(inst_mem_in_wire[1666]), .IN1(inst_mem_in_wire[1698]), .SEL(
        pc[2]), .F(n133) );
  MUX U136 ( .IN0(n133), .IN1(n132), .SEL(pc[3]), .F(n134) );
  MUX U137 ( .IN0(inst_mem_in_wire[1602]), .IN1(inst_mem_in_wire[1634]), .SEL(
        pc[2]), .F(n135) );
  MUX U138 ( .IN0(inst_mem_in_wire[1538]), .IN1(inst_mem_in_wire[1570]), .SEL(
        pc[2]), .F(n136) );
  MUX U139 ( .IN0(n136), .IN1(n135), .SEL(pc[3]), .F(n137) );
  MUX U140 ( .IN0(n137), .IN1(n134), .SEL(pc[4]), .F(n138) );
  MUX U141 ( .IN0(n138), .IN1(n131), .SEL(pc[5]), .F(n139) );
  MUX U142 ( .IN0(inst_mem_in_wire[1474]), .IN1(inst_mem_in_wire[1506]), .SEL(
        pc[2]), .F(n140) );
  MUX U143 ( .IN0(inst_mem_in_wire[1410]), .IN1(inst_mem_in_wire[1442]), .SEL(
        pc[2]), .F(n141) );
  MUX U144 ( .IN0(n141), .IN1(n140), .SEL(pc[3]), .F(n142) );
  MUX U145 ( .IN0(inst_mem_in_wire[1346]), .IN1(inst_mem_in_wire[1378]), .SEL(
        pc[2]), .F(n143) );
  MUX U146 ( .IN0(inst_mem_in_wire[1282]), .IN1(inst_mem_in_wire[1314]), .SEL(
        pc[2]), .F(n144) );
  MUX U147 ( .IN0(n144), .IN1(n143), .SEL(pc[3]), .F(n145) );
  MUX U148 ( .IN0(n145), .IN1(n142), .SEL(pc[4]), .F(n146) );
  MUX U149 ( .IN0(inst_mem_in_wire[1218]), .IN1(inst_mem_in_wire[1250]), .SEL(
        pc[2]), .F(n147) );
  MUX U150 ( .IN0(inst_mem_in_wire[1154]), .IN1(inst_mem_in_wire[1186]), .SEL(
        pc[2]), .F(n148) );
  MUX U151 ( .IN0(n148), .IN1(n147), .SEL(pc[3]), .F(n149) );
  MUX U152 ( .IN0(inst_mem_in_wire[1090]), .IN1(inst_mem_in_wire[1122]), .SEL(
        pc[2]), .F(n150) );
  MUX U153 ( .IN0(inst_mem_in_wire[1026]), .IN1(inst_mem_in_wire[1058]), .SEL(
        pc[2]), .F(n151) );
  MUX U154 ( .IN0(n151), .IN1(n150), .SEL(pc[3]), .F(n152) );
  MUX U155 ( .IN0(n152), .IN1(n149), .SEL(pc[4]), .F(n153) );
  MUX U156 ( .IN0(n153), .IN1(n146), .SEL(pc[5]), .F(n154) );
  MUX U157 ( .IN0(n154), .IN1(n139), .SEL(pc[6]), .F(n155) );
  MUX U158 ( .IN0(inst_mem_in_wire[962]), .IN1(inst_mem_in_wire[994]), .SEL(
        pc[2]), .F(n156) );
  MUX U159 ( .IN0(inst_mem_in_wire[898]), .IN1(inst_mem_in_wire[930]), .SEL(
        pc[2]), .F(n157) );
  MUX U160 ( .IN0(n157), .IN1(n156), .SEL(pc[3]), .F(n158) );
  MUX U161 ( .IN0(inst_mem_in_wire[834]), .IN1(inst_mem_in_wire[866]), .SEL(
        pc[2]), .F(n159) );
  MUX U162 ( .IN0(inst_mem_in_wire[770]), .IN1(inst_mem_in_wire[802]), .SEL(
        pc[2]), .F(n160) );
  MUX U163 ( .IN0(n160), .IN1(n159), .SEL(pc[3]), .F(n161) );
  MUX U164 ( .IN0(n161), .IN1(n158), .SEL(pc[4]), .F(n162) );
  MUX U165 ( .IN0(inst_mem_in_wire[706]), .IN1(inst_mem_in_wire[738]), .SEL(
        pc[2]), .F(n163) );
  MUX U166 ( .IN0(inst_mem_in_wire[642]), .IN1(inst_mem_in_wire[674]), .SEL(
        pc[2]), .F(n164) );
  MUX U167 ( .IN0(n164), .IN1(n163), .SEL(pc[3]), .F(n165) );
  MUX U168 ( .IN0(inst_mem_in_wire[578]), .IN1(inst_mem_in_wire[610]), .SEL(
        pc[2]), .F(n166) );
  MUX U169 ( .IN0(inst_mem_in_wire[514]), .IN1(inst_mem_in_wire[546]), .SEL(
        pc[2]), .F(n167) );
  MUX U170 ( .IN0(n167), .IN1(n166), .SEL(pc[3]), .F(n168) );
  MUX U171 ( .IN0(n168), .IN1(n165), .SEL(pc[4]), .F(n169) );
  MUX U172 ( .IN0(n169), .IN1(n162), .SEL(pc[5]), .F(n170) );
  MUX U173 ( .IN0(inst_mem_in_wire[450]), .IN1(inst_mem_in_wire[482]), .SEL(
        pc[2]), .F(n171) );
  MUX U174 ( .IN0(inst_mem_in_wire[386]), .IN1(inst_mem_in_wire[418]), .SEL(
        pc[2]), .F(n172) );
  MUX U175 ( .IN0(n172), .IN1(n171), .SEL(pc[3]), .F(n173) );
  MUX U176 ( .IN0(inst_mem_in_wire[322]), .IN1(inst_mem_in_wire[354]), .SEL(
        pc[2]), .F(n174) );
  MUX U177 ( .IN0(inst_mem_in_wire[258]), .IN1(inst_mem_in_wire[290]), .SEL(
        pc[2]), .F(n175) );
  MUX U178 ( .IN0(n175), .IN1(n174), .SEL(pc[3]), .F(n176) );
  MUX U179 ( .IN0(n176), .IN1(n173), .SEL(pc[4]), .F(n177) );
  MUX U180 ( .IN0(inst_mem_in_wire[194]), .IN1(inst_mem_in_wire[226]), .SEL(
        pc[2]), .F(n178) );
  MUX U181 ( .IN0(inst_mem_in_wire[130]), .IN1(inst_mem_in_wire[162]), .SEL(
        pc[2]), .F(n179) );
  MUX U182 ( .IN0(n179), .IN1(n178), .SEL(pc[3]), .F(n180) );
  MUX U183 ( .IN0(inst_mem_in_wire[66]), .IN1(inst_mem_in_wire[98]), .SEL(
        pc[2]), .F(n181) );
  MUX U184 ( .IN0(inst_mem_in_wire[2]), .IN1(inst_mem_in_wire[34]), .SEL(pc[2]), .F(n182) );
  MUX U185 ( .IN0(n182), .IN1(n181), .SEL(pc[3]), .F(n183) );
  MUX U186 ( .IN0(n183), .IN1(n180), .SEL(pc[4]), .F(n184) );
  MUX U187 ( .IN0(n184), .IN1(n177), .SEL(pc[5]), .F(n185) );
  MUX U188 ( .IN0(n185), .IN1(n170), .SEL(pc[6]), .F(n186) );
  MUX U189 ( .IN0(n186), .IN1(n155), .SEL(pc[7]), .F(opcode[2]) );
  MUX U190 ( .IN0(inst_mem_in_wire[1987]), .IN1(inst_mem_in_wire[2019]), .SEL(
        pc[2]), .F(n187) );
  MUX U191 ( .IN0(inst_mem_in_wire[1923]), .IN1(inst_mem_in_wire[1955]), .SEL(
        pc[2]), .F(n188) );
  MUX U192 ( .IN0(n188), .IN1(n187), .SEL(pc[3]), .F(n189) );
  MUX U193 ( .IN0(inst_mem_in_wire[1859]), .IN1(inst_mem_in_wire[1891]), .SEL(
        pc[2]), .F(n190) );
  MUX U194 ( .IN0(inst_mem_in_wire[1795]), .IN1(inst_mem_in_wire[1827]), .SEL(
        pc[2]), .F(n191) );
  MUX U195 ( .IN0(n191), .IN1(n190), .SEL(pc[3]), .F(n192) );
  MUX U196 ( .IN0(n192), .IN1(n189), .SEL(pc[4]), .F(n193) );
  MUX U197 ( .IN0(inst_mem_in_wire[1731]), .IN1(inst_mem_in_wire[1763]), .SEL(
        pc[2]), .F(n194) );
  MUX U198 ( .IN0(inst_mem_in_wire[1667]), .IN1(inst_mem_in_wire[1699]), .SEL(
        pc[2]), .F(n195) );
  MUX U199 ( .IN0(n195), .IN1(n194), .SEL(pc[3]), .F(n196) );
  MUX U200 ( .IN0(inst_mem_in_wire[1603]), .IN1(inst_mem_in_wire[1635]), .SEL(
        pc[2]), .F(n197) );
  MUX U201 ( .IN0(inst_mem_in_wire[1539]), .IN1(inst_mem_in_wire[1571]), .SEL(
        pc[2]), .F(n198) );
  MUX U202 ( .IN0(n198), .IN1(n197), .SEL(pc[3]), .F(n199) );
  MUX U203 ( .IN0(n199), .IN1(n196), .SEL(pc[4]), .F(n200) );
  MUX U204 ( .IN0(n200), .IN1(n193), .SEL(pc[5]), .F(n201) );
  MUX U205 ( .IN0(inst_mem_in_wire[1475]), .IN1(inst_mem_in_wire[1507]), .SEL(
        pc[2]), .F(n202) );
  MUX U206 ( .IN0(inst_mem_in_wire[1411]), .IN1(inst_mem_in_wire[1443]), .SEL(
        pc[2]), .F(n203) );
  MUX U207 ( .IN0(n203), .IN1(n202), .SEL(pc[3]), .F(n204) );
  MUX U208 ( .IN0(inst_mem_in_wire[1347]), .IN1(inst_mem_in_wire[1379]), .SEL(
        pc[2]), .F(n205) );
  MUX U209 ( .IN0(inst_mem_in_wire[1283]), .IN1(inst_mem_in_wire[1315]), .SEL(
        pc[2]), .F(n206) );
  MUX U210 ( .IN0(n206), .IN1(n205), .SEL(pc[3]), .F(n207) );
  MUX U211 ( .IN0(n207), .IN1(n204), .SEL(pc[4]), .F(n208) );
  MUX U212 ( .IN0(inst_mem_in_wire[1219]), .IN1(inst_mem_in_wire[1251]), .SEL(
        pc[2]), .F(n209) );
  MUX U213 ( .IN0(inst_mem_in_wire[1155]), .IN1(inst_mem_in_wire[1187]), .SEL(
        pc[2]), .F(n210) );
  MUX U214 ( .IN0(n210), .IN1(n209), .SEL(pc[3]), .F(n211) );
  MUX U215 ( .IN0(inst_mem_in_wire[1091]), .IN1(inst_mem_in_wire[1123]), .SEL(
        pc[2]), .F(n212) );
  MUX U216 ( .IN0(inst_mem_in_wire[1027]), .IN1(inst_mem_in_wire[1059]), .SEL(
        pc[2]), .F(n213) );
  MUX U217 ( .IN0(n213), .IN1(n212), .SEL(pc[3]), .F(n214) );
  MUX U218 ( .IN0(n214), .IN1(n211), .SEL(pc[4]), .F(n215) );
  MUX U219 ( .IN0(n215), .IN1(n208), .SEL(pc[5]), .F(n216) );
  MUX U220 ( .IN0(n216), .IN1(n201), .SEL(pc[6]), .F(n217) );
  MUX U221 ( .IN0(inst_mem_in_wire[963]), .IN1(inst_mem_in_wire[995]), .SEL(
        pc[2]), .F(n218) );
  MUX U222 ( .IN0(inst_mem_in_wire[899]), .IN1(inst_mem_in_wire[931]), .SEL(
        pc[2]), .F(n219) );
  MUX U223 ( .IN0(n219), .IN1(n218), .SEL(pc[3]), .F(n220) );
  MUX U224 ( .IN0(inst_mem_in_wire[835]), .IN1(inst_mem_in_wire[867]), .SEL(
        pc[2]), .F(n221) );
  MUX U225 ( .IN0(inst_mem_in_wire[771]), .IN1(inst_mem_in_wire[803]), .SEL(
        pc[2]), .F(n222) );
  MUX U226 ( .IN0(n222), .IN1(n221), .SEL(pc[3]), .F(n223) );
  MUX U227 ( .IN0(n223), .IN1(n220), .SEL(pc[4]), .F(n224) );
  MUX U228 ( .IN0(inst_mem_in_wire[707]), .IN1(inst_mem_in_wire[739]), .SEL(
        pc[2]), .F(n225) );
  MUX U229 ( .IN0(inst_mem_in_wire[643]), .IN1(inst_mem_in_wire[675]), .SEL(
        pc[2]), .F(n226) );
  MUX U230 ( .IN0(n226), .IN1(n225), .SEL(pc[3]), .F(n227) );
  MUX U231 ( .IN0(inst_mem_in_wire[579]), .IN1(inst_mem_in_wire[611]), .SEL(
        pc[2]), .F(n228) );
  MUX U232 ( .IN0(inst_mem_in_wire[515]), .IN1(inst_mem_in_wire[547]), .SEL(
        pc[2]), .F(n229) );
  MUX U233 ( .IN0(n229), .IN1(n228), .SEL(pc[3]), .F(n230) );
  MUX U234 ( .IN0(n230), .IN1(n227), .SEL(pc[4]), .F(n231) );
  MUX U235 ( .IN0(n231), .IN1(n224), .SEL(pc[5]), .F(n232) );
  MUX U236 ( .IN0(inst_mem_in_wire[451]), .IN1(inst_mem_in_wire[483]), .SEL(
        pc[2]), .F(n233) );
  MUX U237 ( .IN0(inst_mem_in_wire[387]), .IN1(inst_mem_in_wire[419]), .SEL(
        pc[2]), .F(n234) );
  MUX U238 ( .IN0(n234), .IN1(n233), .SEL(pc[3]), .F(n235) );
  MUX U239 ( .IN0(inst_mem_in_wire[323]), .IN1(inst_mem_in_wire[355]), .SEL(
        pc[2]), .F(n236) );
  MUX U240 ( .IN0(inst_mem_in_wire[259]), .IN1(inst_mem_in_wire[291]), .SEL(
        pc[2]), .F(n237) );
  MUX U241 ( .IN0(n237), .IN1(n236), .SEL(pc[3]), .F(n238) );
  MUX U242 ( .IN0(n238), .IN1(n235), .SEL(pc[4]), .F(n239) );
  MUX U243 ( .IN0(inst_mem_in_wire[195]), .IN1(inst_mem_in_wire[227]), .SEL(
        pc[2]), .F(n240) );
  MUX U244 ( .IN0(inst_mem_in_wire[131]), .IN1(inst_mem_in_wire[163]), .SEL(
        pc[2]), .F(n241) );
  MUX U245 ( .IN0(n241), .IN1(n240), .SEL(pc[3]), .F(n242) );
  MUX U246 ( .IN0(inst_mem_in_wire[67]), .IN1(inst_mem_in_wire[99]), .SEL(
        pc[2]), .F(n243) );
  MUX U247 ( .IN0(inst_mem_in_wire[3]), .IN1(inst_mem_in_wire[35]), .SEL(pc[2]), .F(n244) );
  MUX U248 ( .IN0(n244), .IN1(n243), .SEL(pc[3]), .F(n245) );
  MUX U249 ( .IN0(n245), .IN1(n242), .SEL(pc[4]), .F(n246) );
  MUX U250 ( .IN0(n246), .IN1(n239), .SEL(pc[5]), .F(n247) );
  MUX U251 ( .IN0(n247), .IN1(n232), .SEL(pc[6]), .F(n248) );
  MUX U252 ( .IN0(n248), .IN1(n217), .SEL(pc[7]), .F(opcode[3]) );
  MUX U253 ( .IN0(inst_mem_in_wire[1988]), .IN1(inst_mem_in_wire[2020]), .SEL(
        pc[2]), .F(n249) );
  MUX U254 ( .IN0(inst_mem_in_wire[1924]), .IN1(inst_mem_in_wire[1956]), .SEL(
        pc[2]), .F(n250) );
  MUX U255 ( .IN0(n250), .IN1(n249), .SEL(pc[3]), .F(n251) );
  MUX U256 ( .IN0(inst_mem_in_wire[1860]), .IN1(inst_mem_in_wire[1892]), .SEL(
        pc[2]), .F(n252) );
  MUX U257 ( .IN0(inst_mem_in_wire[1796]), .IN1(inst_mem_in_wire[1828]), .SEL(
        pc[2]), .F(n253) );
  MUX U258 ( .IN0(n253), .IN1(n252), .SEL(pc[3]), .F(n254) );
  MUX U259 ( .IN0(n254), .IN1(n251), .SEL(pc[4]), .F(n255) );
  MUX U260 ( .IN0(inst_mem_in_wire[1732]), .IN1(inst_mem_in_wire[1764]), .SEL(
        pc[2]), .F(n256) );
  MUX U261 ( .IN0(inst_mem_in_wire[1668]), .IN1(inst_mem_in_wire[1700]), .SEL(
        pc[2]), .F(n257) );
  MUX U262 ( .IN0(n257), .IN1(n256), .SEL(pc[3]), .F(n258) );
  MUX U263 ( .IN0(inst_mem_in_wire[1604]), .IN1(inst_mem_in_wire[1636]), .SEL(
        pc[2]), .F(n259) );
  MUX U264 ( .IN0(inst_mem_in_wire[1540]), .IN1(inst_mem_in_wire[1572]), .SEL(
        pc[2]), .F(n260) );
  MUX U265 ( .IN0(n260), .IN1(n259), .SEL(pc[3]), .F(n261) );
  MUX U266 ( .IN0(n261), .IN1(n258), .SEL(pc[4]), .F(n262) );
  MUX U267 ( .IN0(n262), .IN1(n255), .SEL(pc[5]), .F(n263) );
  MUX U268 ( .IN0(inst_mem_in_wire[1476]), .IN1(inst_mem_in_wire[1508]), .SEL(
        pc[2]), .F(n264) );
  MUX U269 ( .IN0(inst_mem_in_wire[1412]), .IN1(inst_mem_in_wire[1444]), .SEL(
        pc[2]), .F(n265) );
  MUX U270 ( .IN0(n265), .IN1(n264), .SEL(pc[3]), .F(n266) );
  MUX U271 ( .IN0(inst_mem_in_wire[1348]), .IN1(inst_mem_in_wire[1380]), .SEL(
        pc[2]), .F(n267) );
  MUX U272 ( .IN0(inst_mem_in_wire[1284]), .IN1(inst_mem_in_wire[1316]), .SEL(
        pc[2]), .F(n268) );
  MUX U273 ( .IN0(n268), .IN1(n267), .SEL(pc[3]), .F(n269) );
  MUX U274 ( .IN0(n269), .IN1(n266), .SEL(pc[4]), .F(n270) );
  MUX U275 ( .IN0(inst_mem_in_wire[1220]), .IN1(inst_mem_in_wire[1252]), .SEL(
        pc[2]), .F(n271) );
  MUX U276 ( .IN0(inst_mem_in_wire[1156]), .IN1(inst_mem_in_wire[1188]), .SEL(
        pc[2]), .F(n272) );
  MUX U277 ( .IN0(n272), .IN1(n271), .SEL(pc[3]), .F(n273) );
  MUX U278 ( .IN0(inst_mem_in_wire[1092]), .IN1(inst_mem_in_wire[1124]), .SEL(
        pc[2]), .F(n274) );
  MUX U279 ( .IN0(inst_mem_in_wire[1028]), .IN1(inst_mem_in_wire[1060]), .SEL(
        pc[2]), .F(n275) );
  MUX U280 ( .IN0(n275), .IN1(n274), .SEL(pc[3]), .F(n276) );
  MUX U281 ( .IN0(n276), .IN1(n273), .SEL(pc[4]), .F(n277) );
  MUX U282 ( .IN0(n277), .IN1(n270), .SEL(pc[5]), .F(n278) );
  MUX U283 ( .IN0(n278), .IN1(n263), .SEL(pc[6]), .F(n279) );
  MUX U284 ( .IN0(inst_mem_in_wire[964]), .IN1(inst_mem_in_wire[996]), .SEL(
        pc[2]), .F(n280) );
  MUX U285 ( .IN0(inst_mem_in_wire[900]), .IN1(inst_mem_in_wire[932]), .SEL(
        pc[2]), .F(n281) );
  MUX U286 ( .IN0(n281), .IN1(n280), .SEL(pc[3]), .F(n282) );
  MUX U287 ( .IN0(inst_mem_in_wire[836]), .IN1(inst_mem_in_wire[868]), .SEL(
        pc[2]), .F(n283) );
  MUX U288 ( .IN0(inst_mem_in_wire[772]), .IN1(inst_mem_in_wire[804]), .SEL(
        pc[2]), .F(n284) );
  MUX U289 ( .IN0(n284), .IN1(n283), .SEL(pc[3]), .F(n285) );
  MUX U290 ( .IN0(n285), .IN1(n282), .SEL(pc[4]), .F(n286) );
  MUX U291 ( .IN0(inst_mem_in_wire[708]), .IN1(inst_mem_in_wire[740]), .SEL(
        pc[2]), .F(n287) );
  MUX U292 ( .IN0(inst_mem_in_wire[644]), .IN1(inst_mem_in_wire[676]), .SEL(
        pc[2]), .F(n288) );
  MUX U293 ( .IN0(n288), .IN1(n287), .SEL(pc[3]), .F(n289) );
  MUX U294 ( .IN0(inst_mem_in_wire[580]), .IN1(inst_mem_in_wire[612]), .SEL(
        pc[2]), .F(n290) );
  MUX U295 ( .IN0(inst_mem_in_wire[516]), .IN1(inst_mem_in_wire[548]), .SEL(
        pc[2]), .F(n291) );
  MUX U296 ( .IN0(n291), .IN1(n290), .SEL(pc[3]), .F(n292) );
  MUX U297 ( .IN0(n292), .IN1(n289), .SEL(pc[4]), .F(n293) );
  MUX U298 ( .IN0(n293), .IN1(n286), .SEL(pc[5]), .F(n294) );
  MUX U299 ( .IN0(inst_mem_in_wire[452]), .IN1(inst_mem_in_wire[484]), .SEL(
        pc[2]), .F(n295) );
  MUX U300 ( .IN0(inst_mem_in_wire[388]), .IN1(inst_mem_in_wire[420]), .SEL(
        pc[2]), .F(n296) );
  MUX U301 ( .IN0(n296), .IN1(n295), .SEL(pc[3]), .F(n297) );
  MUX U302 ( .IN0(inst_mem_in_wire[324]), .IN1(inst_mem_in_wire[356]), .SEL(
        pc[2]), .F(n298) );
  MUX U303 ( .IN0(inst_mem_in_wire[260]), .IN1(inst_mem_in_wire[292]), .SEL(
        pc[2]), .F(n299) );
  MUX U304 ( .IN0(n299), .IN1(n298), .SEL(pc[3]), .F(n300) );
  MUX U305 ( .IN0(n300), .IN1(n297), .SEL(pc[4]), .F(n301) );
  MUX U306 ( .IN0(inst_mem_in_wire[196]), .IN1(inst_mem_in_wire[228]), .SEL(
        pc[2]), .F(n302) );
  MUX U307 ( .IN0(inst_mem_in_wire[132]), .IN1(inst_mem_in_wire[164]), .SEL(
        pc[2]), .F(n303) );
  MUX U308 ( .IN0(n303), .IN1(n302), .SEL(pc[3]), .F(n304) );
  MUX U309 ( .IN0(inst_mem_in_wire[68]), .IN1(inst_mem_in_wire[100]), .SEL(
        pc[2]), .F(n305) );
  MUX U310 ( .IN0(inst_mem_in_wire[4]), .IN1(inst_mem_in_wire[36]), .SEL(pc[2]), .F(n306) );
  MUX U311 ( .IN0(n306), .IN1(n305), .SEL(pc[3]), .F(n307) );
  MUX U312 ( .IN0(n307), .IN1(n304), .SEL(pc[4]), .F(n308) );
  MUX U313 ( .IN0(n308), .IN1(n301), .SEL(pc[5]), .F(n309) );
  MUX U314 ( .IN0(n309), .IN1(n294), .SEL(pc[6]), .F(n310) );
  MUX U315 ( .IN0(n310), .IN1(n279), .SEL(pc[7]), .F(opcode[4]) );
  MUX U316 ( .IN0(inst_mem_in_wire[1989]), .IN1(inst_mem_in_wire[2021]), .SEL(
        pc[2]), .F(n311) );
  MUX U317 ( .IN0(inst_mem_in_wire[1925]), .IN1(inst_mem_in_wire[1957]), .SEL(
        pc[2]), .F(n312) );
  MUX U318 ( .IN0(n312), .IN1(n311), .SEL(pc[3]), .F(n313) );
  MUX U319 ( .IN0(inst_mem_in_wire[1861]), .IN1(inst_mem_in_wire[1893]), .SEL(
        pc[2]), .F(n314) );
  MUX U320 ( .IN0(inst_mem_in_wire[1797]), .IN1(inst_mem_in_wire[1829]), .SEL(
        pc[2]), .F(n315) );
  MUX U321 ( .IN0(n315), .IN1(n314), .SEL(pc[3]), .F(n316) );
  MUX U322 ( .IN0(n316), .IN1(n313), .SEL(pc[4]), .F(n317) );
  MUX U323 ( .IN0(inst_mem_in_wire[1733]), .IN1(inst_mem_in_wire[1765]), .SEL(
        pc[2]), .F(n318) );
  MUX U324 ( .IN0(inst_mem_in_wire[1669]), .IN1(inst_mem_in_wire[1701]), .SEL(
        pc[2]), .F(n319) );
  MUX U325 ( .IN0(n319), .IN1(n318), .SEL(pc[3]), .F(n320) );
  MUX U326 ( .IN0(inst_mem_in_wire[1605]), .IN1(inst_mem_in_wire[1637]), .SEL(
        pc[2]), .F(n321) );
  MUX U327 ( .IN0(inst_mem_in_wire[1541]), .IN1(inst_mem_in_wire[1573]), .SEL(
        pc[2]), .F(n322) );
  MUX U328 ( .IN0(n322), .IN1(n321), .SEL(pc[3]), .F(n323) );
  MUX U329 ( .IN0(n323), .IN1(n320), .SEL(pc[4]), .F(n324) );
  MUX U330 ( .IN0(n324), .IN1(n317), .SEL(pc[5]), .F(n325) );
  MUX U331 ( .IN0(inst_mem_in_wire[1477]), .IN1(inst_mem_in_wire[1509]), .SEL(
        pc[2]), .F(n326) );
  MUX U332 ( .IN0(inst_mem_in_wire[1413]), .IN1(inst_mem_in_wire[1445]), .SEL(
        pc[2]), .F(n327) );
  MUX U333 ( .IN0(n327), .IN1(n326), .SEL(pc[3]), .F(n328) );
  MUX U334 ( .IN0(inst_mem_in_wire[1349]), .IN1(inst_mem_in_wire[1381]), .SEL(
        pc[2]), .F(n329) );
  MUX U335 ( .IN0(inst_mem_in_wire[1285]), .IN1(inst_mem_in_wire[1317]), .SEL(
        pc[2]), .F(n330) );
  MUX U336 ( .IN0(n330), .IN1(n329), .SEL(pc[3]), .F(n331) );
  MUX U337 ( .IN0(n331), .IN1(n328), .SEL(pc[4]), .F(n332) );
  MUX U338 ( .IN0(inst_mem_in_wire[1221]), .IN1(inst_mem_in_wire[1253]), .SEL(
        pc[2]), .F(n333) );
  MUX U339 ( .IN0(inst_mem_in_wire[1157]), .IN1(inst_mem_in_wire[1189]), .SEL(
        pc[2]), .F(n334) );
  MUX U340 ( .IN0(n334), .IN1(n333), .SEL(pc[3]), .F(n335) );
  MUX U341 ( .IN0(inst_mem_in_wire[1093]), .IN1(inst_mem_in_wire[1125]), .SEL(
        pc[2]), .F(n336) );
  MUX U342 ( .IN0(inst_mem_in_wire[1029]), .IN1(inst_mem_in_wire[1061]), .SEL(
        pc[2]), .F(n337) );
  MUX U343 ( .IN0(n337), .IN1(n336), .SEL(pc[3]), .F(n338) );
  MUX U344 ( .IN0(n338), .IN1(n335), .SEL(pc[4]), .F(n339) );
  MUX U345 ( .IN0(n339), .IN1(n332), .SEL(pc[5]), .F(n340) );
  MUX U346 ( .IN0(n340), .IN1(n325), .SEL(pc[6]), .F(n341) );
  MUX U347 ( .IN0(inst_mem_in_wire[965]), .IN1(inst_mem_in_wire[997]), .SEL(
        pc[2]), .F(n342) );
  MUX U348 ( .IN0(inst_mem_in_wire[901]), .IN1(inst_mem_in_wire[933]), .SEL(
        pc[2]), .F(n343) );
  MUX U349 ( .IN0(n343), .IN1(n342), .SEL(pc[3]), .F(n344) );
  MUX U350 ( .IN0(inst_mem_in_wire[837]), .IN1(inst_mem_in_wire[869]), .SEL(
        pc[2]), .F(n345) );
  MUX U351 ( .IN0(inst_mem_in_wire[773]), .IN1(inst_mem_in_wire[805]), .SEL(
        pc[2]), .F(n346) );
  MUX U352 ( .IN0(n346), .IN1(n345), .SEL(pc[3]), .F(n347) );
  MUX U353 ( .IN0(n347), .IN1(n344), .SEL(pc[4]), .F(n348) );
  MUX U354 ( .IN0(inst_mem_in_wire[709]), .IN1(inst_mem_in_wire[741]), .SEL(
        pc[2]), .F(n349) );
  MUX U355 ( .IN0(inst_mem_in_wire[645]), .IN1(inst_mem_in_wire[677]), .SEL(
        pc[2]), .F(n350) );
  MUX U356 ( .IN0(n350), .IN1(n349), .SEL(pc[3]), .F(n351) );
  MUX U357 ( .IN0(inst_mem_in_wire[581]), .IN1(inst_mem_in_wire[613]), .SEL(
        pc[2]), .F(n352) );
  MUX U358 ( .IN0(inst_mem_in_wire[517]), .IN1(inst_mem_in_wire[549]), .SEL(
        pc[2]), .F(n353) );
  MUX U359 ( .IN0(n353), .IN1(n352), .SEL(pc[3]), .F(n354) );
  MUX U360 ( .IN0(n354), .IN1(n351), .SEL(pc[4]), .F(n355) );
  MUX U361 ( .IN0(n355), .IN1(n348), .SEL(pc[5]), .F(n356) );
  MUX U362 ( .IN0(inst_mem_in_wire[453]), .IN1(inst_mem_in_wire[485]), .SEL(
        pc[2]), .F(n357) );
  MUX U363 ( .IN0(inst_mem_in_wire[389]), .IN1(inst_mem_in_wire[421]), .SEL(
        pc[2]), .F(n358) );
  MUX U364 ( .IN0(n358), .IN1(n357), .SEL(pc[3]), .F(n359) );
  MUX U365 ( .IN0(inst_mem_in_wire[325]), .IN1(inst_mem_in_wire[357]), .SEL(
        pc[2]), .F(n360) );
  MUX U366 ( .IN0(inst_mem_in_wire[261]), .IN1(inst_mem_in_wire[293]), .SEL(
        pc[2]), .F(n361) );
  MUX U367 ( .IN0(n361), .IN1(n360), .SEL(pc[3]), .F(n362) );
  MUX U368 ( .IN0(n362), .IN1(n359), .SEL(pc[4]), .F(n363) );
  MUX U369 ( .IN0(inst_mem_in_wire[197]), .IN1(inst_mem_in_wire[229]), .SEL(
        pc[2]), .F(n364) );
  MUX U370 ( .IN0(inst_mem_in_wire[133]), .IN1(inst_mem_in_wire[165]), .SEL(
        pc[2]), .F(n365) );
  MUX U371 ( .IN0(n365), .IN1(n364), .SEL(pc[3]), .F(n366) );
  MUX U372 ( .IN0(inst_mem_in_wire[69]), .IN1(inst_mem_in_wire[101]), .SEL(
        pc[2]), .F(n367) );
  MUX U373 ( .IN0(inst_mem_in_wire[5]), .IN1(inst_mem_in_wire[37]), .SEL(pc[2]), .F(n368) );
  MUX U374 ( .IN0(n368), .IN1(n367), .SEL(pc[3]), .F(n369) );
  MUX U375 ( .IN0(n369), .IN1(n366), .SEL(pc[4]), .F(n370) );
  MUX U376 ( .IN0(n370), .IN1(n363), .SEL(pc[5]), .F(n371) );
  MUX U377 ( .IN0(n371), .IN1(n356), .SEL(pc[6]), .F(n372) );
  MUX U378 ( .IN0(n372), .IN1(n341), .SEL(pc[7]), .F(opcode[5]) );
  MUX U379 ( .IN0(inst_mem_in_wire[1990]), .IN1(inst_mem_in_wire[2022]), .SEL(
        pc[2]), .F(n373) );
  MUX U380 ( .IN0(inst_mem_in_wire[1926]), .IN1(inst_mem_in_wire[1958]), .SEL(
        pc[2]), .F(n374) );
  MUX U381 ( .IN0(n374), .IN1(n373), .SEL(pc[3]), .F(n375) );
  MUX U382 ( .IN0(inst_mem_in_wire[1862]), .IN1(inst_mem_in_wire[1894]), .SEL(
        pc[2]), .F(n376) );
  MUX U383 ( .IN0(inst_mem_in_wire[1798]), .IN1(inst_mem_in_wire[1830]), .SEL(
        pc[2]), .F(n377) );
  MUX U384 ( .IN0(n377), .IN1(n376), .SEL(pc[3]), .F(n378) );
  MUX U385 ( .IN0(n378), .IN1(n375), .SEL(pc[4]), .F(n379) );
  MUX U386 ( .IN0(inst_mem_in_wire[1734]), .IN1(inst_mem_in_wire[1766]), .SEL(
        pc[2]), .F(n380) );
  MUX U387 ( .IN0(inst_mem_in_wire[1670]), .IN1(inst_mem_in_wire[1702]), .SEL(
        pc[2]), .F(n381) );
  MUX U388 ( .IN0(n381), .IN1(n380), .SEL(pc[3]), .F(n382) );
  MUX U389 ( .IN0(inst_mem_in_wire[1606]), .IN1(inst_mem_in_wire[1638]), .SEL(
        pc[2]), .F(n383) );
  MUX U390 ( .IN0(inst_mem_in_wire[1542]), .IN1(inst_mem_in_wire[1574]), .SEL(
        pc[2]), .F(n384) );
  MUX U391 ( .IN0(n384), .IN1(n383), .SEL(pc[3]), .F(n385) );
  MUX U392 ( .IN0(n385), .IN1(n382), .SEL(pc[4]), .F(n386) );
  MUX U393 ( .IN0(n386), .IN1(n379), .SEL(pc[5]), .F(n387) );
  MUX U394 ( .IN0(inst_mem_in_wire[1478]), .IN1(inst_mem_in_wire[1510]), .SEL(
        pc[2]), .F(n388) );
  MUX U395 ( .IN0(inst_mem_in_wire[1414]), .IN1(inst_mem_in_wire[1446]), .SEL(
        pc[2]), .F(n389) );
  MUX U396 ( .IN0(n389), .IN1(n388), .SEL(pc[3]), .F(n390) );
  MUX U397 ( .IN0(inst_mem_in_wire[1350]), .IN1(inst_mem_in_wire[1382]), .SEL(
        pc[2]), .F(n391) );
  MUX U398 ( .IN0(inst_mem_in_wire[1286]), .IN1(inst_mem_in_wire[1318]), .SEL(
        pc[2]), .F(n392) );
  MUX U399 ( .IN0(n392), .IN1(n391), .SEL(pc[3]), .F(n393) );
  MUX U400 ( .IN0(n393), .IN1(n390), .SEL(pc[4]), .F(n394) );
  MUX U401 ( .IN0(inst_mem_in_wire[1222]), .IN1(inst_mem_in_wire[1254]), .SEL(
        pc[2]), .F(n395) );
  MUX U402 ( .IN0(inst_mem_in_wire[1158]), .IN1(inst_mem_in_wire[1190]), .SEL(
        pc[2]), .F(n396) );
  MUX U403 ( .IN0(n396), .IN1(n395), .SEL(pc[3]), .F(n397) );
  MUX U404 ( .IN0(inst_mem_in_wire[1094]), .IN1(inst_mem_in_wire[1126]), .SEL(
        pc[2]), .F(n398) );
  MUX U405 ( .IN0(inst_mem_in_wire[1030]), .IN1(inst_mem_in_wire[1062]), .SEL(
        pc[2]), .F(n399) );
  MUX U406 ( .IN0(n399), .IN1(n398), .SEL(pc[3]), .F(n400) );
  MUX U407 ( .IN0(n400), .IN1(n397), .SEL(pc[4]), .F(n401) );
  MUX U408 ( .IN0(n401), .IN1(n394), .SEL(pc[5]), .F(n402) );
  MUX U409 ( .IN0(n402), .IN1(n387), .SEL(pc[6]), .F(n403) );
  MUX U410 ( .IN0(inst_mem_in_wire[966]), .IN1(inst_mem_in_wire[998]), .SEL(
        pc[2]), .F(n404) );
  MUX U411 ( .IN0(inst_mem_in_wire[902]), .IN1(inst_mem_in_wire[934]), .SEL(
        pc[2]), .F(n405) );
  MUX U412 ( .IN0(n405), .IN1(n404), .SEL(pc[3]), .F(n406) );
  MUX U413 ( .IN0(inst_mem_in_wire[838]), .IN1(inst_mem_in_wire[870]), .SEL(
        pc[2]), .F(n407) );
  MUX U414 ( .IN0(inst_mem_in_wire[774]), .IN1(inst_mem_in_wire[806]), .SEL(
        pc[2]), .F(n408) );
  MUX U415 ( .IN0(n408), .IN1(n407), .SEL(pc[3]), .F(n409) );
  MUX U416 ( .IN0(n409), .IN1(n406), .SEL(pc[4]), .F(n410) );
  MUX U417 ( .IN0(inst_mem_in_wire[710]), .IN1(inst_mem_in_wire[742]), .SEL(
        pc[2]), .F(n411) );
  MUX U418 ( .IN0(inst_mem_in_wire[646]), .IN1(inst_mem_in_wire[678]), .SEL(
        pc[2]), .F(n412) );
  MUX U419 ( .IN0(n412), .IN1(n411), .SEL(pc[3]), .F(n413) );
  MUX U420 ( .IN0(inst_mem_in_wire[582]), .IN1(inst_mem_in_wire[614]), .SEL(
        pc[2]), .F(n414) );
  MUX U421 ( .IN0(inst_mem_in_wire[518]), .IN1(inst_mem_in_wire[550]), .SEL(
        pc[2]), .F(n415) );
  MUX U422 ( .IN0(n415), .IN1(n414), .SEL(pc[3]), .F(n416) );
  MUX U423 ( .IN0(n416), .IN1(n413), .SEL(pc[4]), .F(n417) );
  MUX U424 ( .IN0(n417), .IN1(n410), .SEL(pc[5]), .F(n418) );
  MUX U425 ( .IN0(inst_mem_in_wire[454]), .IN1(inst_mem_in_wire[486]), .SEL(
        pc[2]), .F(n419) );
  MUX U426 ( .IN0(inst_mem_in_wire[390]), .IN1(inst_mem_in_wire[422]), .SEL(
        pc[2]), .F(n420) );
  MUX U427 ( .IN0(n420), .IN1(n419), .SEL(pc[3]), .F(n421) );
  MUX U428 ( .IN0(inst_mem_in_wire[326]), .IN1(inst_mem_in_wire[358]), .SEL(
        pc[2]), .F(n422) );
  MUX U429 ( .IN0(inst_mem_in_wire[262]), .IN1(inst_mem_in_wire[294]), .SEL(
        pc[2]), .F(n423) );
  MUX U430 ( .IN0(n423), .IN1(n422), .SEL(pc[3]), .F(n424) );
  MUX U431 ( .IN0(n424), .IN1(n421), .SEL(pc[4]), .F(n425) );
  MUX U432 ( .IN0(inst_mem_in_wire[198]), .IN1(inst_mem_in_wire[230]), .SEL(
        pc[2]), .F(n426) );
  MUX U433 ( .IN0(inst_mem_in_wire[134]), .IN1(inst_mem_in_wire[166]), .SEL(
        pc[2]), .F(n427) );
  MUX U434 ( .IN0(n427), .IN1(n426), .SEL(pc[3]), .F(n428) );
  MUX U435 ( .IN0(inst_mem_in_wire[70]), .IN1(inst_mem_in_wire[102]), .SEL(
        pc[2]), .F(n429) );
  MUX U436 ( .IN0(inst_mem_in_wire[6]), .IN1(inst_mem_in_wire[38]), .SEL(pc[2]), .F(n430) );
  MUX U437 ( .IN0(n430), .IN1(n429), .SEL(pc[3]), .F(n431) );
  MUX U438 ( .IN0(n431), .IN1(n428), .SEL(pc[4]), .F(n432) );
  MUX U439 ( .IN0(n432), .IN1(n425), .SEL(pc[5]), .F(n433) );
  MUX U440 ( .IN0(n433), .IN1(n418), .SEL(pc[6]), .F(n434) );
  MUX U441 ( .IN0(n434), .IN1(n403), .SEL(pc[7]), .F(opcode[6]) );
  MUX U442 ( .IN0(inst_mem_in_wire[1991]), .IN1(inst_mem_in_wire[2023]), .SEL(
        pc[2]), .F(n435) );
  MUX U443 ( .IN0(inst_mem_in_wire[1927]), .IN1(inst_mem_in_wire[1959]), .SEL(
        pc[2]), .F(n436) );
  MUX U444 ( .IN0(n436), .IN1(n435), .SEL(pc[3]), .F(n437) );
  MUX U445 ( .IN0(inst_mem_in_wire[1863]), .IN1(inst_mem_in_wire[1895]), .SEL(
        pc[2]), .F(n438) );
  MUX U446 ( .IN0(inst_mem_in_wire[1799]), .IN1(inst_mem_in_wire[1831]), .SEL(
        pc[2]), .F(n439) );
  MUX U447 ( .IN0(n439), .IN1(n438), .SEL(pc[3]), .F(n440) );
  MUX U448 ( .IN0(n440), .IN1(n437), .SEL(pc[4]), .F(n441) );
  MUX U449 ( .IN0(inst_mem_in_wire[1735]), .IN1(inst_mem_in_wire[1767]), .SEL(
        pc[2]), .F(n442) );
  MUX U450 ( .IN0(inst_mem_in_wire[1671]), .IN1(inst_mem_in_wire[1703]), .SEL(
        pc[2]), .F(n443) );
  MUX U451 ( .IN0(n443), .IN1(n442), .SEL(pc[3]), .F(n444) );
  MUX U452 ( .IN0(inst_mem_in_wire[1607]), .IN1(inst_mem_in_wire[1639]), .SEL(
        pc[2]), .F(n445) );
  MUX U453 ( .IN0(inst_mem_in_wire[1543]), .IN1(inst_mem_in_wire[1575]), .SEL(
        pc[2]), .F(n446) );
  MUX U454 ( .IN0(n446), .IN1(n445), .SEL(pc[3]), .F(n447) );
  MUX U455 ( .IN0(n447), .IN1(n444), .SEL(pc[4]), .F(n448) );
  MUX U456 ( .IN0(n448), .IN1(n441), .SEL(pc[5]), .F(n449) );
  MUX U457 ( .IN0(inst_mem_in_wire[1479]), .IN1(inst_mem_in_wire[1511]), .SEL(
        pc[2]), .F(n450) );
  MUX U458 ( .IN0(inst_mem_in_wire[1415]), .IN1(inst_mem_in_wire[1447]), .SEL(
        pc[2]), .F(n451) );
  MUX U459 ( .IN0(n451), .IN1(n450), .SEL(pc[3]), .F(n452) );
  MUX U460 ( .IN0(inst_mem_in_wire[1351]), .IN1(inst_mem_in_wire[1383]), .SEL(
        pc[2]), .F(n453) );
  MUX U461 ( .IN0(inst_mem_in_wire[1287]), .IN1(inst_mem_in_wire[1319]), .SEL(
        pc[2]), .F(n454) );
  MUX U462 ( .IN0(n454), .IN1(n453), .SEL(pc[3]), .F(n455) );
  MUX U463 ( .IN0(n455), .IN1(n452), .SEL(pc[4]), .F(n456) );
  MUX U464 ( .IN0(inst_mem_in_wire[1223]), .IN1(inst_mem_in_wire[1255]), .SEL(
        pc[2]), .F(n457) );
  MUX U465 ( .IN0(inst_mem_in_wire[1159]), .IN1(inst_mem_in_wire[1191]), .SEL(
        pc[2]), .F(n458) );
  MUX U466 ( .IN0(n458), .IN1(n457), .SEL(pc[3]), .F(n459) );
  MUX U467 ( .IN0(inst_mem_in_wire[1095]), .IN1(inst_mem_in_wire[1127]), .SEL(
        pc[2]), .F(n460) );
  MUX U468 ( .IN0(inst_mem_in_wire[1031]), .IN1(inst_mem_in_wire[1063]), .SEL(
        pc[2]), .F(n461) );
  MUX U469 ( .IN0(n461), .IN1(n460), .SEL(pc[3]), .F(n462) );
  MUX U470 ( .IN0(n462), .IN1(n459), .SEL(pc[4]), .F(n463) );
  MUX U471 ( .IN0(n463), .IN1(n456), .SEL(pc[5]), .F(n464) );
  MUX U472 ( .IN0(n464), .IN1(n449), .SEL(pc[6]), .F(n465) );
  MUX U473 ( .IN0(inst_mem_in_wire[967]), .IN1(inst_mem_in_wire[999]), .SEL(
        pc[2]), .F(n466) );
  MUX U474 ( .IN0(inst_mem_in_wire[903]), .IN1(inst_mem_in_wire[935]), .SEL(
        pc[2]), .F(n467) );
  MUX U475 ( .IN0(n467), .IN1(n466), .SEL(pc[3]), .F(n468) );
  MUX U476 ( .IN0(inst_mem_in_wire[839]), .IN1(inst_mem_in_wire[871]), .SEL(
        pc[2]), .F(n469) );
  MUX U477 ( .IN0(inst_mem_in_wire[775]), .IN1(inst_mem_in_wire[807]), .SEL(
        pc[2]), .F(n470) );
  MUX U478 ( .IN0(n470), .IN1(n469), .SEL(pc[3]), .F(n471) );
  MUX U479 ( .IN0(n471), .IN1(n468), .SEL(pc[4]), .F(n472) );
  MUX U480 ( .IN0(inst_mem_in_wire[711]), .IN1(inst_mem_in_wire[743]), .SEL(
        pc[2]), .F(n473) );
  MUX U481 ( .IN0(inst_mem_in_wire[647]), .IN1(inst_mem_in_wire[679]), .SEL(
        pc[2]), .F(n474) );
  MUX U482 ( .IN0(n474), .IN1(n473), .SEL(pc[3]), .F(n475) );
  MUX U483 ( .IN0(inst_mem_in_wire[583]), .IN1(inst_mem_in_wire[615]), .SEL(
        pc[2]), .F(n476) );
  MUX U484 ( .IN0(inst_mem_in_wire[519]), .IN1(inst_mem_in_wire[551]), .SEL(
        pc[2]), .F(n477) );
  MUX U485 ( .IN0(n477), .IN1(n476), .SEL(pc[3]), .F(n478) );
  MUX U486 ( .IN0(n478), .IN1(n475), .SEL(pc[4]), .F(n479) );
  MUX U487 ( .IN0(n479), .IN1(n472), .SEL(pc[5]), .F(n480) );
  MUX U488 ( .IN0(inst_mem_in_wire[455]), .IN1(inst_mem_in_wire[487]), .SEL(
        pc[2]), .F(n481) );
  MUX U489 ( .IN0(inst_mem_in_wire[391]), .IN1(inst_mem_in_wire[423]), .SEL(
        pc[2]), .F(n482) );
  MUX U490 ( .IN0(n482), .IN1(n481), .SEL(pc[3]), .F(n483) );
  MUX U491 ( .IN0(inst_mem_in_wire[327]), .IN1(inst_mem_in_wire[359]), .SEL(
        pc[2]), .F(n484) );
  MUX U492 ( .IN0(inst_mem_in_wire[263]), .IN1(inst_mem_in_wire[295]), .SEL(
        pc[2]), .F(n485) );
  MUX U493 ( .IN0(n485), .IN1(n484), .SEL(pc[3]), .F(n486) );
  MUX U494 ( .IN0(n486), .IN1(n483), .SEL(pc[4]), .F(n487) );
  MUX U495 ( .IN0(inst_mem_in_wire[199]), .IN1(inst_mem_in_wire[231]), .SEL(
        pc[2]), .F(n488) );
  MUX U496 ( .IN0(inst_mem_in_wire[135]), .IN1(inst_mem_in_wire[167]), .SEL(
        pc[2]), .F(n489) );
  MUX U497 ( .IN0(n489), .IN1(n488), .SEL(pc[3]), .F(n490) );
  MUX U498 ( .IN0(inst_mem_in_wire[71]), .IN1(inst_mem_in_wire[103]), .SEL(
        pc[2]), .F(n491) );
  MUX U499 ( .IN0(inst_mem_in_wire[7]), .IN1(inst_mem_in_wire[39]), .SEL(pc[2]), .F(n492) );
  MUX U500 ( .IN0(n492), .IN1(n491), .SEL(pc[3]), .F(n493) );
  MUX U501 ( .IN0(n493), .IN1(n490), .SEL(pc[4]), .F(n494) );
  MUX U502 ( .IN0(n494), .IN1(n487), .SEL(pc[5]), .F(n495) );
  MUX U503 ( .IN0(n495), .IN1(n480), .SEL(pc[6]), .F(n496) );
  MUX U504 ( .IN0(n496), .IN1(n465), .SEL(pc[7]), .F(opcode[7]) );
  MUX U505 ( .IN0(inst_mem_in_wire[1992]), .IN1(inst_mem_in_wire[2024]), .SEL(
        pc[2]), .F(n497) );
  MUX U506 ( .IN0(inst_mem_in_wire[1928]), .IN1(inst_mem_in_wire[1960]), .SEL(
        pc[2]), .F(n498) );
  MUX U507 ( .IN0(n498), .IN1(n497), .SEL(pc[3]), .F(n499) );
  MUX U508 ( .IN0(inst_mem_in_wire[1864]), .IN1(inst_mem_in_wire[1896]), .SEL(
        pc[2]), .F(n500) );
  MUX U509 ( .IN0(inst_mem_in_wire[1800]), .IN1(inst_mem_in_wire[1832]), .SEL(
        pc[2]), .F(n501) );
  MUX U510 ( .IN0(n501), .IN1(n500), .SEL(pc[3]), .F(n502) );
  MUX U511 ( .IN0(n502), .IN1(n499), .SEL(pc[4]), .F(n503) );
  MUX U512 ( .IN0(inst_mem_in_wire[1736]), .IN1(inst_mem_in_wire[1768]), .SEL(
        pc[2]), .F(n504) );
  MUX U513 ( .IN0(inst_mem_in_wire[1672]), .IN1(inst_mem_in_wire[1704]), .SEL(
        pc[2]), .F(n505) );
  MUX U514 ( .IN0(n505), .IN1(n504), .SEL(pc[3]), .F(n506) );
  MUX U515 ( .IN0(inst_mem_in_wire[1608]), .IN1(inst_mem_in_wire[1640]), .SEL(
        pc[2]), .F(n507) );
  MUX U516 ( .IN0(inst_mem_in_wire[1544]), .IN1(inst_mem_in_wire[1576]), .SEL(
        pc[2]), .F(n508) );
  MUX U517 ( .IN0(n508), .IN1(n507), .SEL(pc[3]), .F(n509) );
  MUX U518 ( .IN0(n509), .IN1(n506), .SEL(pc[4]), .F(n510) );
  MUX U519 ( .IN0(n510), .IN1(n503), .SEL(pc[5]), .F(n511) );
  MUX U520 ( .IN0(inst_mem_in_wire[1480]), .IN1(inst_mem_in_wire[1512]), .SEL(
        pc[2]), .F(n512) );
  MUX U521 ( .IN0(inst_mem_in_wire[1416]), .IN1(inst_mem_in_wire[1448]), .SEL(
        pc[2]), .F(n513) );
  MUX U522 ( .IN0(n513), .IN1(n512), .SEL(pc[3]), .F(n514) );
  MUX U523 ( .IN0(inst_mem_in_wire[1352]), .IN1(inst_mem_in_wire[1384]), .SEL(
        pc[2]), .F(n515) );
  MUX U524 ( .IN0(inst_mem_in_wire[1288]), .IN1(inst_mem_in_wire[1320]), .SEL(
        pc[2]), .F(n516) );
  MUX U525 ( .IN0(n516), .IN1(n515), .SEL(pc[3]), .F(n517) );
  MUX U526 ( .IN0(n517), .IN1(n514), .SEL(pc[4]), .F(n518) );
  MUX U527 ( .IN0(inst_mem_in_wire[1224]), .IN1(inst_mem_in_wire[1256]), .SEL(
        pc[2]), .F(n519) );
  MUX U528 ( .IN0(inst_mem_in_wire[1160]), .IN1(inst_mem_in_wire[1192]), .SEL(
        pc[2]), .F(n520) );
  MUX U529 ( .IN0(n520), .IN1(n519), .SEL(pc[3]), .F(n521) );
  MUX U530 ( .IN0(inst_mem_in_wire[1096]), .IN1(inst_mem_in_wire[1128]), .SEL(
        pc[2]), .F(n522) );
  MUX U531 ( .IN0(inst_mem_in_wire[1032]), .IN1(inst_mem_in_wire[1064]), .SEL(
        pc[2]), .F(n523) );
  MUX U532 ( .IN0(n523), .IN1(n522), .SEL(pc[3]), .F(n524) );
  MUX U533 ( .IN0(n524), .IN1(n521), .SEL(pc[4]), .F(n525) );
  MUX U534 ( .IN0(n525), .IN1(n518), .SEL(pc[5]), .F(n526) );
  MUX U535 ( .IN0(n526), .IN1(n511), .SEL(pc[6]), .F(n527) );
  MUX U536 ( .IN0(inst_mem_in_wire[968]), .IN1(inst_mem_in_wire[1000]), .SEL(
        pc[2]), .F(n528) );
  MUX U537 ( .IN0(inst_mem_in_wire[904]), .IN1(inst_mem_in_wire[936]), .SEL(
        pc[2]), .F(n529) );
  MUX U538 ( .IN0(n529), .IN1(n528), .SEL(pc[3]), .F(n530) );
  MUX U539 ( .IN0(inst_mem_in_wire[840]), .IN1(inst_mem_in_wire[872]), .SEL(
        pc[2]), .F(n531) );
  MUX U540 ( .IN0(inst_mem_in_wire[776]), .IN1(inst_mem_in_wire[808]), .SEL(
        pc[2]), .F(n532) );
  MUX U541 ( .IN0(n532), .IN1(n531), .SEL(pc[3]), .F(n533) );
  MUX U542 ( .IN0(n533), .IN1(n530), .SEL(pc[4]), .F(n534) );
  MUX U543 ( .IN0(inst_mem_in_wire[712]), .IN1(inst_mem_in_wire[744]), .SEL(
        pc[2]), .F(n535) );
  MUX U544 ( .IN0(inst_mem_in_wire[648]), .IN1(inst_mem_in_wire[680]), .SEL(
        pc[2]), .F(n536) );
  MUX U545 ( .IN0(n536), .IN1(n535), .SEL(pc[3]), .F(n537) );
  MUX U546 ( .IN0(inst_mem_in_wire[584]), .IN1(inst_mem_in_wire[616]), .SEL(
        pc[2]), .F(n538) );
  MUX U547 ( .IN0(inst_mem_in_wire[520]), .IN1(inst_mem_in_wire[552]), .SEL(
        pc[2]), .F(n539) );
  MUX U548 ( .IN0(n539), .IN1(n538), .SEL(pc[3]), .F(n540) );
  MUX U549 ( .IN0(n540), .IN1(n537), .SEL(pc[4]), .F(n541) );
  MUX U550 ( .IN0(n541), .IN1(n534), .SEL(pc[5]), .F(n542) );
  MUX U551 ( .IN0(inst_mem_in_wire[456]), .IN1(inst_mem_in_wire[488]), .SEL(
        pc[2]), .F(n543) );
  MUX U552 ( .IN0(inst_mem_in_wire[392]), .IN1(inst_mem_in_wire[424]), .SEL(
        pc[2]), .F(n544) );
  MUX U553 ( .IN0(n544), .IN1(n543), .SEL(pc[3]), .F(n545) );
  MUX U554 ( .IN0(inst_mem_in_wire[328]), .IN1(inst_mem_in_wire[360]), .SEL(
        pc[2]), .F(n546) );
  MUX U555 ( .IN0(inst_mem_in_wire[264]), .IN1(inst_mem_in_wire[296]), .SEL(
        pc[2]), .F(n547) );
  MUX U556 ( .IN0(n547), .IN1(n546), .SEL(pc[3]), .F(n548) );
  MUX U557 ( .IN0(n548), .IN1(n545), .SEL(pc[4]), .F(n549) );
  MUX U558 ( .IN0(inst_mem_in_wire[200]), .IN1(inst_mem_in_wire[232]), .SEL(
        pc[2]), .F(n550) );
  MUX U559 ( .IN0(inst_mem_in_wire[136]), .IN1(inst_mem_in_wire[168]), .SEL(
        pc[2]), .F(n551) );
  MUX U560 ( .IN0(n551), .IN1(n550), .SEL(pc[3]), .F(n552) );
  MUX U561 ( .IN0(inst_mem_in_wire[72]), .IN1(inst_mem_in_wire[104]), .SEL(
        pc[2]), .F(n553) );
  MUX U562 ( .IN0(inst_mem_in_wire[8]), .IN1(inst_mem_in_wire[40]), .SEL(pc[2]), .F(n554) );
  MUX U563 ( .IN0(n554), .IN1(n553), .SEL(pc[3]), .F(n555) );
  MUX U564 ( .IN0(n555), .IN1(n552), .SEL(pc[4]), .F(n556) );
  MUX U565 ( .IN0(n556), .IN1(n549), .SEL(pc[5]), .F(n557) );
  MUX U566 ( .IN0(n557), .IN1(n542), .SEL(pc[6]), .F(n558) );
  MUX U567 ( .IN0(n558), .IN1(n527), .SEL(pc[7]), .F(opcode[8]) );
  MUX U568 ( .IN0(inst_mem_in_wire[1993]), .IN1(inst_mem_in_wire[2025]), .SEL(
        pc[2]), .F(n559) );
  MUX U569 ( .IN0(inst_mem_in_wire[1929]), .IN1(inst_mem_in_wire[1961]), .SEL(
        pc[2]), .F(n560) );
  MUX U570 ( .IN0(n560), .IN1(n559), .SEL(pc[3]), .F(n561) );
  MUX U571 ( .IN0(inst_mem_in_wire[1865]), .IN1(inst_mem_in_wire[1897]), .SEL(
        pc[2]), .F(n562) );
  MUX U572 ( .IN0(inst_mem_in_wire[1801]), .IN1(inst_mem_in_wire[1833]), .SEL(
        pc[2]), .F(n563) );
  MUX U573 ( .IN0(n563), .IN1(n562), .SEL(pc[3]), .F(n564) );
  MUX U574 ( .IN0(n564), .IN1(n561), .SEL(pc[4]), .F(n565) );
  MUX U575 ( .IN0(inst_mem_in_wire[1737]), .IN1(inst_mem_in_wire[1769]), .SEL(
        pc[2]), .F(n566) );
  MUX U576 ( .IN0(inst_mem_in_wire[1673]), .IN1(inst_mem_in_wire[1705]), .SEL(
        pc[2]), .F(n567) );
  MUX U577 ( .IN0(n567), .IN1(n566), .SEL(pc[3]), .F(n568) );
  MUX U578 ( .IN0(inst_mem_in_wire[1609]), .IN1(inst_mem_in_wire[1641]), .SEL(
        pc[2]), .F(n569) );
  MUX U579 ( .IN0(inst_mem_in_wire[1545]), .IN1(inst_mem_in_wire[1577]), .SEL(
        pc[2]), .F(n570) );
  MUX U580 ( .IN0(n570), .IN1(n569), .SEL(pc[3]), .F(n571) );
  MUX U581 ( .IN0(n571), .IN1(n568), .SEL(pc[4]), .F(n572) );
  MUX U582 ( .IN0(n572), .IN1(n565), .SEL(pc[5]), .F(n573) );
  MUX U583 ( .IN0(inst_mem_in_wire[1481]), .IN1(inst_mem_in_wire[1513]), .SEL(
        pc[2]), .F(n574) );
  MUX U584 ( .IN0(inst_mem_in_wire[1417]), .IN1(inst_mem_in_wire[1449]), .SEL(
        pc[2]), .F(n575) );
  MUX U585 ( .IN0(n575), .IN1(n574), .SEL(pc[3]), .F(n576) );
  MUX U586 ( .IN0(inst_mem_in_wire[1353]), .IN1(inst_mem_in_wire[1385]), .SEL(
        pc[2]), .F(n577) );
  MUX U587 ( .IN0(inst_mem_in_wire[1289]), .IN1(inst_mem_in_wire[1321]), .SEL(
        pc[2]), .F(n578) );
  MUX U588 ( .IN0(n578), .IN1(n577), .SEL(pc[3]), .F(n579) );
  MUX U589 ( .IN0(n579), .IN1(n576), .SEL(pc[4]), .F(n580) );
  MUX U590 ( .IN0(inst_mem_in_wire[1225]), .IN1(inst_mem_in_wire[1257]), .SEL(
        pc[2]), .F(n581) );
  MUX U591 ( .IN0(inst_mem_in_wire[1161]), .IN1(inst_mem_in_wire[1193]), .SEL(
        pc[2]), .F(n582) );
  MUX U592 ( .IN0(n582), .IN1(n581), .SEL(pc[3]), .F(n583) );
  MUX U593 ( .IN0(inst_mem_in_wire[1097]), .IN1(inst_mem_in_wire[1129]), .SEL(
        pc[2]), .F(n584) );
  MUX U594 ( .IN0(inst_mem_in_wire[1033]), .IN1(inst_mem_in_wire[1065]), .SEL(
        pc[2]), .F(n585) );
  MUX U595 ( .IN0(n585), .IN1(n584), .SEL(pc[3]), .F(n586) );
  MUX U596 ( .IN0(n586), .IN1(n583), .SEL(pc[4]), .F(n587) );
  MUX U597 ( .IN0(n587), .IN1(n580), .SEL(pc[5]), .F(n588) );
  MUX U598 ( .IN0(n588), .IN1(n573), .SEL(pc[6]), .F(n589) );
  MUX U599 ( .IN0(inst_mem_in_wire[969]), .IN1(inst_mem_in_wire[1001]), .SEL(
        pc[2]), .F(n590) );
  MUX U600 ( .IN0(inst_mem_in_wire[905]), .IN1(inst_mem_in_wire[937]), .SEL(
        pc[2]), .F(n591) );
  MUX U601 ( .IN0(n591), .IN1(n590), .SEL(pc[3]), .F(n592) );
  MUX U602 ( .IN0(inst_mem_in_wire[841]), .IN1(inst_mem_in_wire[873]), .SEL(
        pc[2]), .F(n593) );
  MUX U603 ( .IN0(inst_mem_in_wire[777]), .IN1(inst_mem_in_wire[809]), .SEL(
        pc[2]), .F(n594) );
  MUX U604 ( .IN0(n594), .IN1(n593), .SEL(pc[3]), .F(n595) );
  MUX U605 ( .IN0(n595), .IN1(n592), .SEL(pc[4]), .F(n596) );
  MUX U606 ( .IN0(inst_mem_in_wire[713]), .IN1(inst_mem_in_wire[745]), .SEL(
        pc[2]), .F(n597) );
  MUX U607 ( .IN0(inst_mem_in_wire[649]), .IN1(inst_mem_in_wire[681]), .SEL(
        pc[2]), .F(n598) );
  MUX U608 ( .IN0(n598), .IN1(n597), .SEL(pc[3]), .F(n599) );
  MUX U609 ( .IN0(inst_mem_in_wire[585]), .IN1(inst_mem_in_wire[617]), .SEL(
        pc[2]), .F(n600) );
  MUX U610 ( .IN0(inst_mem_in_wire[521]), .IN1(inst_mem_in_wire[553]), .SEL(
        pc[2]), .F(n601) );
  MUX U611 ( .IN0(n601), .IN1(n600), .SEL(pc[3]), .F(n602) );
  MUX U612 ( .IN0(n602), .IN1(n599), .SEL(pc[4]), .F(n603) );
  MUX U613 ( .IN0(n603), .IN1(n596), .SEL(pc[5]), .F(n604) );
  MUX U614 ( .IN0(inst_mem_in_wire[457]), .IN1(inst_mem_in_wire[489]), .SEL(
        pc[2]), .F(n605) );
  MUX U615 ( .IN0(inst_mem_in_wire[393]), .IN1(inst_mem_in_wire[425]), .SEL(
        pc[2]), .F(n606) );
  MUX U616 ( .IN0(n606), .IN1(n605), .SEL(pc[3]), .F(n607) );
  MUX U617 ( .IN0(inst_mem_in_wire[329]), .IN1(inst_mem_in_wire[361]), .SEL(
        pc[2]), .F(n608) );
  MUX U618 ( .IN0(inst_mem_in_wire[265]), .IN1(inst_mem_in_wire[297]), .SEL(
        pc[2]), .F(n609) );
  MUX U619 ( .IN0(n609), .IN1(n608), .SEL(pc[3]), .F(n610) );
  MUX U620 ( .IN0(n610), .IN1(n607), .SEL(pc[4]), .F(n611) );
  MUX U621 ( .IN0(inst_mem_in_wire[201]), .IN1(inst_mem_in_wire[233]), .SEL(
        pc[2]), .F(n612) );
  MUX U622 ( .IN0(inst_mem_in_wire[137]), .IN1(inst_mem_in_wire[169]), .SEL(
        pc[2]), .F(n613) );
  MUX U623 ( .IN0(n613), .IN1(n612), .SEL(pc[3]), .F(n614) );
  MUX U624 ( .IN0(inst_mem_in_wire[73]), .IN1(inst_mem_in_wire[105]), .SEL(
        pc[2]), .F(n615) );
  MUX U625 ( .IN0(inst_mem_in_wire[9]), .IN1(inst_mem_in_wire[41]), .SEL(pc[2]), .F(n616) );
  MUX U626 ( .IN0(n616), .IN1(n615), .SEL(pc[3]), .F(n617) );
  MUX U627 ( .IN0(n617), .IN1(n614), .SEL(pc[4]), .F(n618) );
  MUX U628 ( .IN0(n618), .IN1(n611), .SEL(pc[5]), .F(n619) );
  MUX U629 ( .IN0(n619), .IN1(n604), .SEL(pc[6]), .F(n620) );
  MUX U630 ( .IN0(n620), .IN1(n589), .SEL(pc[7]), .F(opcode[9]) );
  MUX U631 ( .IN0(inst_mem_in_wire[1994]), .IN1(inst_mem_in_wire[2026]), .SEL(
        pc[2]), .F(n621) );
  MUX U632 ( .IN0(inst_mem_in_wire[1930]), .IN1(inst_mem_in_wire[1962]), .SEL(
        pc[2]), .F(n622) );
  MUX U633 ( .IN0(n622), .IN1(n621), .SEL(pc[3]), .F(n623) );
  MUX U634 ( .IN0(inst_mem_in_wire[1866]), .IN1(inst_mem_in_wire[1898]), .SEL(
        pc[2]), .F(n624) );
  MUX U635 ( .IN0(inst_mem_in_wire[1802]), .IN1(inst_mem_in_wire[1834]), .SEL(
        pc[2]), .F(n625) );
  MUX U636 ( .IN0(n625), .IN1(n624), .SEL(pc[3]), .F(n626) );
  MUX U637 ( .IN0(n626), .IN1(n623), .SEL(pc[4]), .F(n627) );
  MUX U638 ( .IN0(inst_mem_in_wire[1738]), .IN1(inst_mem_in_wire[1770]), .SEL(
        pc[2]), .F(n628) );
  MUX U639 ( .IN0(inst_mem_in_wire[1674]), .IN1(inst_mem_in_wire[1706]), .SEL(
        pc[2]), .F(n629) );
  MUX U640 ( .IN0(n629), .IN1(n628), .SEL(pc[3]), .F(n630) );
  MUX U641 ( .IN0(inst_mem_in_wire[1610]), .IN1(inst_mem_in_wire[1642]), .SEL(
        pc[2]), .F(n631) );
  MUX U642 ( .IN0(inst_mem_in_wire[1546]), .IN1(inst_mem_in_wire[1578]), .SEL(
        pc[2]), .F(n632) );
  MUX U643 ( .IN0(n632), .IN1(n631), .SEL(pc[3]), .F(n633) );
  MUX U644 ( .IN0(n633), .IN1(n630), .SEL(pc[4]), .F(n634) );
  MUX U645 ( .IN0(n634), .IN1(n627), .SEL(pc[5]), .F(n635) );
  MUX U646 ( .IN0(inst_mem_in_wire[1482]), .IN1(inst_mem_in_wire[1514]), .SEL(
        pc[2]), .F(n636) );
  MUX U647 ( .IN0(inst_mem_in_wire[1418]), .IN1(inst_mem_in_wire[1450]), .SEL(
        pc[2]), .F(n637) );
  MUX U648 ( .IN0(n637), .IN1(n636), .SEL(pc[3]), .F(n638) );
  MUX U649 ( .IN0(inst_mem_in_wire[1354]), .IN1(inst_mem_in_wire[1386]), .SEL(
        pc[2]), .F(n639) );
  MUX U650 ( .IN0(inst_mem_in_wire[1290]), .IN1(inst_mem_in_wire[1322]), .SEL(
        pc[2]), .F(n640) );
  MUX U651 ( .IN0(n640), .IN1(n639), .SEL(pc[3]), .F(n641) );
  MUX U652 ( .IN0(n641), .IN1(n638), .SEL(pc[4]), .F(n642) );
  MUX U653 ( .IN0(inst_mem_in_wire[1226]), .IN1(inst_mem_in_wire[1258]), .SEL(
        pc[2]), .F(n643) );
  MUX U654 ( .IN0(inst_mem_in_wire[1162]), .IN1(inst_mem_in_wire[1194]), .SEL(
        pc[2]), .F(n644) );
  MUX U655 ( .IN0(n644), .IN1(n643), .SEL(pc[3]), .F(n645) );
  MUX U656 ( .IN0(inst_mem_in_wire[1098]), .IN1(inst_mem_in_wire[1130]), .SEL(
        pc[2]), .F(n646) );
  MUX U657 ( .IN0(inst_mem_in_wire[1034]), .IN1(inst_mem_in_wire[1066]), .SEL(
        pc[2]), .F(n647) );
  MUX U658 ( .IN0(n647), .IN1(n646), .SEL(pc[3]), .F(n648) );
  MUX U659 ( .IN0(n648), .IN1(n645), .SEL(pc[4]), .F(n649) );
  MUX U660 ( .IN0(n649), .IN1(n642), .SEL(pc[5]), .F(n650) );
  MUX U661 ( .IN0(n650), .IN1(n635), .SEL(pc[6]), .F(n651) );
  MUX U662 ( .IN0(inst_mem_in_wire[970]), .IN1(inst_mem_in_wire[1002]), .SEL(
        pc[2]), .F(n652) );
  MUX U663 ( .IN0(inst_mem_in_wire[906]), .IN1(inst_mem_in_wire[938]), .SEL(
        pc[2]), .F(n653) );
  MUX U664 ( .IN0(n653), .IN1(n652), .SEL(pc[3]), .F(n654) );
  MUX U665 ( .IN0(inst_mem_in_wire[842]), .IN1(inst_mem_in_wire[874]), .SEL(
        pc[2]), .F(n655) );
  MUX U666 ( .IN0(inst_mem_in_wire[778]), .IN1(inst_mem_in_wire[810]), .SEL(
        pc[2]), .F(n656) );
  MUX U667 ( .IN0(n656), .IN1(n655), .SEL(pc[3]), .F(n657) );
  MUX U668 ( .IN0(n657), .IN1(n654), .SEL(pc[4]), .F(n658) );
  MUX U669 ( .IN0(inst_mem_in_wire[714]), .IN1(inst_mem_in_wire[746]), .SEL(
        pc[2]), .F(n659) );
  MUX U670 ( .IN0(inst_mem_in_wire[650]), .IN1(inst_mem_in_wire[682]), .SEL(
        pc[2]), .F(n660) );
  MUX U671 ( .IN0(n660), .IN1(n659), .SEL(pc[3]), .F(n661) );
  MUX U672 ( .IN0(inst_mem_in_wire[586]), .IN1(inst_mem_in_wire[618]), .SEL(
        pc[2]), .F(n662) );
  MUX U673 ( .IN0(inst_mem_in_wire[522]), .IN1(inst_mem_in_wire[554]), .SEL(
        pc[2]), .F(n663) );
  MUX U674 ( .IN0(n663), .IN1(n662), .SEL(pc[3]), .F(n664) );
  MUX U675 ( .IN0(n664), .IN1(n661), .SEL(pc[4]), .F(n665) );
  MUX U676 ( .IN0(n665), .IN1(n658), .SEL(pc[5]), .F(n666) );
  MUX U677 ( .IN0(inst_mem_in_wire[458]), .IN1(inst_mem_in_wire[490]), .SEL(
        pc[2]), .F(n667) );
  MUX U678 ( .IN0(inst_mem_in_wire[394]), .IN1(inst_mem_in_wire[426]), .SEL(
        pc[2]), .F(n668) );
  MUX U679 ( .IN0(n668), .IN1(n667), .SEL(pc[3]), .F(n669) );
  MUX U680 ( .IN0(inst_mem_in_wire[330]), .IN1(inst_mem_in_wire[362]), .SEL(
        pc[2]), .F(n670) );
  MUX U681 ( .IN0(inst_mem_in_wire[266]), .IN1(inst_mem_in_wire[298]), .SEL(
        pc[2]), .F(n671) );
  MUX U682 ( .IN0(n671), .IN1(n670), .SEL(pc[3]), .F(n672) );
  MUX U683 ( .IN0(n672), .IN1(n669), .SEL(pc[4]), .F(n673) );
  MUX U684 ( .IN0(inst_mem_in_wire[202]), .IN1(inst_mem_in_wire[234]), .SEL(
        pc[2]), .F(n674) );
  MUX U685 ( .IN0(inst_mem_in_wire[138]), .IN1(inst_mem_in_wire[170]), .SEL(
        pc[2]), .F(n675) );
  MUX U686 ( .IN0(n675), .IN1(n674), .SEL(pc[3]), .F(n676) );
  MUX U687 ( .IN0(inst_mem_in_wire[74]), .IN1(inst_mem_in_wire[106]), .SEL(
        pc[2]), .F(n677) );
  MUX U688 ( .IN0(inst_mem_in_wire[10]), .IN1(inst_mem_in_wire[42]), .SEL(
        pc[2]), .F(n678) );
  MUX U689 ( .IN0(n678), .IN1(n677), .SEL(pc[3]), .F(n679) );
  MUX U690 ( .IN0(n679), .IN1(n676), .SEL(pc[4]), .F(n680) );
  MUX U691 ( .IN0(n680), .IN1(n673), .SEL(pc[5]), .F(n681) );
  MUX U692 ( .IN0(n681), .IN1(n666), .SEL(pc[6]), .F(n682) );
  MUX U693 ( .IN0(n682), .IN1(n651), .SEL(pc[7]), .F(opcode[10]) );
  MUX U694 ( .IN0(inst_mem_in_wire[1995]), .IN1(inst_mem_in_wire[2027]), .SEL(
        pc[2]), .F(n683) );
  MUX U695 ( .IN0(inst_mem_in_wire[1931]), .IN1(inst_mem_in_wire[1963]), .SEL(
        pc[2]), .F(n684) );
  MUX U696 ( .IN0(n684), .IN1(n683), .SEL(pc[3]), .F(n685) );
  MUX U697 ( .IN0(inst_mem_in_wire[1867]), .IN1(inst_mem_in_wire[1899]), .SEL(
        pc[2]), .F(n686) );
  MUX U698 ( .IN0(inst_mem_in_wire[1803]), .IN1(inst_mem_in_wire[1835]), .SEL(
        pc[2]), .F(n687) );
  MUX U699 ( .IN0(n687), .IN1(n686), .SEL(pc[3]), .F(n688) );
  MUX U700 ( .IN0(n688), .IN1(n685), .SEL(pc[4]), .F(n689) );
  MUX U701 ( .IN0(inst_mem_in_wire[1739]), .IN1(inst_mem_in_wire[1771]), .SEL(
        pc[2]), .F(n690) );
  MUX U702 ( .IN0(inst_mem_in_wire[1675]), .IN1(inst_mem_in_wire[1707]), .SEL(
        pc[2]), .F(n691) );
  MUX U703 ( .IN0(n691), .IN1(n690), .SEL(pc[3]), .F(n692) );
  MUX U704 ( .IN0(inst_mem_in_wire[1611]), .IN1(inst_mem_in_wire[1643]), .SEL(
        pc[2]), .F(n693) );
  MUX U705 ( .IN0(inst_mem_in_wire[1547]), .IN1(inst_mem_in_wire[1579]), .SEL(
        pc[2]), .F(n694) );
  MUX U706 ( .IN0(n694), .IN1(n693), .SEL(pc[3]), .F(n695) );
  MUX U707 ( .IN0(n695), .IN1(n692), .SEL(pc[4]), .F(n696) );
  MUX U708 ( .IN0(n696), .IN1(n689), .SEL(pc[5]), .F(n697) );
  MUX U709 ( .IN0(inst_mem_in_wire[1483]), .IN1(inst_mem_in_wire[1515]), .SEL(
        pc[2]), .F(n698) );
  MUX U710 ( .IN0(inst_mem_in_wire[1419]), .IN1(inst_mem_in_wire[1451]), .SEL(
        pc[2]), .F(n699) );
  MUX U711 ( .IN0(n699), .IN1(n698), .SEL(pc[3]), .F(n700) );
  MUX U712 ( .IN0(inst_mem_in_wire[1355]), .IN1(inst_mem_in_wire[1387]), .SEL(
        pc[2]), .F(n701) );
  MUX U713 ( .IN0(inst_mem_in_wire[1291]), .IN1(inst_mem_in_wire[1323]), .SEL(
        pc[2]), .F(n702) );
  MUX U714 ( .IN0(n702), .IN1(n701), .SEL(pc[3]), .F(n703) );
  MUX U715 ( .IN0(n703), .IN1(n700), .SEL(pc[4]), .F(n704) );
  MUX U716 ( .IN0(inst_mem_in_wire[1227]), .IN1(inst_mem_in_wire[1259]), .SEL(
        pc[2]), .F(n705) );
  MUX U717 ( .IN0(inst_mem_in_wire[1163]), .IN1(inst_mem_in_wire[1195]), .SEL(
        pc[2]), .F(n706) );
  MUX U718 ( .IN0(n706), .IN1(n705), .SEL(pc[3]), .F(n707) );
  MUX U719 ( .IN0(inst_mem_in_wire[1099]), .IN1(inst_mem_in_wire[1131]), .SEL(
        pc[2]), .F(n708) );
  MUX U720 ( .IN0(inst_mem_in_wire[1035]), .IN1(inst_mem_in_wire[1067]), .SEL(
        pc[2]), .F(n709) );
  MUX U721 ( .IN0(n709), .IN1(n708), .SEL(pc[3]), .F(n710) );
  MUX U722 ( .IN0(n710), .IN1(n707), .SEL(pc[4]), .F(n711) );
  MUX U723 ( .IN0(n711), .IN1(n704), .SEL(pc[5]), .F(n712) );
  MUX U724 ( .IN0(n712), .IN1(n697), .SEL(pc[6]), .F(n713) );
  MUX U725 ( .IN0(inst_mem_in_wire[971]), .IN1(inst_mem_in_wire[1003]), .SEL(
        pc[2]), .F(n714) );
  MUX U726 ( .IN0(inst_mem_in_wire[907]), .IN1(inst_mem_in_wire[939]), .SEL(
        pc[2]), .F(n715) );
  MUX U727 ( .IN0(n715), .IN1(n714), .SEL(pc[3]), .F(n716) );
  MUX U728 ( .IN0(inst_mem_in_wire[843]), .IN1(inst_mem_in_wire[875]), .SEL(
        pc[2]), .F(n717) );
  MUX U729 ( .IN0(inst_mem_in_wire[779]), .IN1(inst_mem_in_wire[811]), .SEL(
        pc[2]), .F(n718) );
  MUX U730 ( .IN0(n718), .IN1(n717), .SEL(pc[3]), .F(n719) );
  MUX U731 ( .IN0(n719), .IN1(n716), .SEL(pc[4]), .F(n720) );
  MUX U732 ( .IN0(inst_mem_in_wire[715]), .IN1(inst_mem_in_wire[747]), .SEL(
        pc[2]), .F(n721) );
  MUX U733 ( .IN0(inst_mem_in_wire[651]), .IN1(inst_mem_in_wire[683]), .SEL(
        pc[2]), .F(n722) );
  MUX U734 ( .IN0(n722), .IN1(n721), .SEL(pc[3]), .F(n723) );
  MUX U735 ( .IN0(inst_mem_in_wire[587]), .IN1(inst_mem_in_wire[619]), .SEL(
        pc[2]), .F(n724) );
  MUX U736 ( .IN0(inst_mem_in_wire[523]), .IN1(inst_mem_in_wire[555]), .SEL(
        pc[2]), .F(n725) );
  MUX U737 ( .IN0(n725), .IN1(n724), .SEL(pc[3]), .F(n726) );
  MUX U738 ( .IN0(n726), .IN1(n723), .SEL(pc[4]), .F(n727) );
  MUX U739 ( .IN0(n727), .IN1(n720), .SEL(pc[5]), .F(n728) );
  MUX U740 ( .IN0(inst_mem_in_wire[459]), .IN1(inst_mem_in_wire[491]), .SEL(
        pc[2]), .F(n729) );
  MUX U741 ( .IN0(inst_mem_in_wire[395]), .IN1(inst_mem_in_wire[427]), .SEL(
        pc[2]), .F(n730) );
  MUX U742 ( .IN0(n730), .IN1(n729), .SEL(pc[3]), .F(n731) );
  MUX U743 ( .IN0(inst_mem_in_wire[331]), .IN1(inst_mem_in_wire[363]), .SEL(
        pc[2]), .F(n732) );
  MUX U744 ( .IN0(inst_mem_in_wire[267]), .IN1(inst_mem_in_wire[299]), .SEL(
        pc[2]), .F(n733) );
  MUX U745 ( .IN0(n733), .IN1(n732), .SEL(pc[3]), .F(n734) );
  MUX U746 ( .IN0(n734), .IN1(n731), .SEL(pc[4]), .F(n735) );
  MUX U747 ( .IN0(inst_mem_in_wire[203]), .IN1(inst_mem_in_wire[235]), .SEL(
        pc[2]), .F(n736) );
  MUX U748 ( .IN0(inst_mem_in_wire[139]), .IN1(inst_mem_in_wire[171]), .SEL(
        pc[2]), .F(n737) );
  MUX U749 ( .IN0(n737), .IN1(n736), .SEL(pc[3]), .F(n738) );
  MUX U750 ( .IN0(inst_mem_in_wire[75]), .IN1(inst_mem_in_wire[107]), .SEL(
        pc[2]), .F(n739) );
  MUX U751 ( .IN0(inst_mem_in_wire[11]), .IN1(inst_mem_in_wire[43]), .SEL(
        pc[2]), .F(n740) );
  MUX U752 ( .IN0(n740), .IN1(n739), .SEL(pc[3]), .F(n741) );
  MUX U753 ( .IN0(n741), .IN1(n738), .SEL(pc[4]), .F(n742) );
  MUX U754 ( .IN0(n742), .IN1(n735), .SEL(pc[5]), .F(n743) );
  MUX U755 ( .IN0(n743), .IN1(n728), .SEL(pc[6]), .F(n744) );
  MUX U756 ( .IN0(n744), .IN1(n713), .SEL(pc[7]), .F(opcode[11]) );
  MUX U757 ( .IN0(inst_mem_in_wire[1996]), .IN1(inst_mem_in_wire[2028]), .SEL(
        pc[2]), .F(n745) );
  MUX U758 ( .IN0(inst_mem_in_wire[1932]), .IN1(inst_mem_in_wire[1964]), .SEL(
        pc[2]), .F(n746) );
  MUX U759 ( .IN0(n746), .IN1(n745), .SEL(pc[3]), .F(n747) );
  MUX U760 ( .IN0(inst_mem_in_wire[1868]), .IN1(inst_mem_in_wire[1900]), .SEL(
        pc[2]), .F(n748) );
  MUX U761 ( .IN0(inst_mem_in_wire[1804]), .IN1(inst_mem_in_wire[1836]), .SEL(
        pc[2]), .F(n749) );
  MUX U762 ( .IN0(n749), .IN1(n748), .SEL(pc[3]), .F(n750) );
  MUX U763 ( .IN0(n750), .IN1(n747), .SEL(pc[4]), .F(n751) );
  MUX U764 ( .IN0(inst_mem_in_wire[1740]), .IN1(inst_mem_in_wire[1772]), .SEL(
        pc[2]), .F(n752) );
  MUX U765 ( .IN0(inst_mem_in_wire[1676]), .IN1(inst_mem_in_wire[1708]), .SEL(
        pc[2]), .F(n753) );
  MUX U766 ( .IN0(n753), .IN1(n752), .SEL(pc[3]), .F(n754) );
  MUX U767 ( .IN0(inst_mem_in_wire[1612]), .IN1(inst_mem_in_wire[1644]), .SEL(
        pc[2]), .F(n755) );
  MUX U768 ( .IN0(inst_mem_in_wire[1548]), .IN1(inst_mem_in_wire[1580]), .SEL(
        pc[2]), .F(n756) );
  MUX U769 ( .IN0(n756), .IN1(n755), .SEL(pc[3]), .F(n757) );
  MUX U770 ( .IN0(n757), .IN1(n754), .SEL(pc[4]), .F(n758) );
  MUX U771 ( .IN0(n758), .IN1(n751), .SEL(pc[5]), .F(n759) );
  MUX U772 ( .IN0(inst_mem_in_wire[1484]), .IN1(inst_mem_in_wire[1516]), .SEL(
        pc[2]), .F(n760) );
  MUX U773 ( .IN0(inst_mem_in_wire[1420]), .IN1(inst_mem_in_wire[1452]), .SEL(
        pc[2]), .F(n761) );
  MUX U774 ( .IN0(n761), .IN1(n760), .SEL(pc[3]), .F(n762) );
  MUX U775 ( .IN0(inst_mem_in_wire[1356]), .IN1(inst_mem_in_wire[1388]), .SEL(
        pc[2]), .F(n763) );
  MUX U776 ( .IN0(inst_mem_in_wire[1292]), .IN1(inst_mem_in_wire[1324]), .SEL(
        pc[2]), .F(n764) );
  MUX U777 ( .IN0(n764), .IN1(n763), .SEL(pc[3]), .F(n765) );
  MUX U778 ( .IN0(n765), .IN1(n762), .SEL(pc[4]), .F(n766) );
  MUX U779 ( .IN0(inst_mem_in_wire[1228]), .IN1(inst_mem_in_wire[1260]), .SEL(
        pc[2]), .F(n767) );
  MUX U780 ( .IN0(inst_mem_in_wire[1164]), .IN1(inst_mem_in_wire[1196]), .SEL(
        pc[2]), .F(n768) );
  MUX U781 ( .IN0(n768), .IN1(n767), .SEL(pc[3]), .F(n769) );
  MUX U782 ( .IN0(inst_mem_in_wire[1100]), .IN1(inst_mem_in_wire[1132]), .SEL(
        pc[2]), .F(n770) );
  MUX U783 ( .IN0(inst_mem_in_wire[1036]), .IN1(inst_mem_in_wire[1068]), .SEL(
        pc[2]), .F(n771) );
  MUX U784 ( .IN0(n771), .IN1(n770), .SEL(pc[3]), .F(n772) );
  MUX U785 ( .IN0(n772), .IN1(n769), .SEL(pc[4]), .F(n773) );
  MUX U786 ( .IN0(n773), .IN1(n766), .SEL(pc[5]), .F(n774) );
  MUX U787 ( .IN0(n774), .IN1(n759), .SEL(pc[6]), .F(n775) );
  MUX U788 ( .IN0(inst_mem_in_wire[972]), .IN1(inst_mem_in_wire[1004]), .SEL(
        pc[2]), .F(n776) );
  MUX U789 ( .IN0(inst_mem_in_wire[908]), .IN1(inst_mem_in_wire[940]), .SEL(
        pc[2]), .F(n777) );
  MUX U790 ( .IN0(n777), .IN1(n776), .SEL(pc[3]), .F(n778) );
  MUX U791 ( .IN0(inst_mem_in_wire[844]), .IN1(inst_mem_in_wire[876]), .SEL(
        pc[2]), .F(n779) );
  MUX U792 ( .IN0(inst_mem_in_wire[780]), .IN1(inst_mem_in_wire[812]), .SEL(
        pc[2]), .F(n780) );
  MUX U793 ( .IN0(n780), .IN1(n779), .SEL(pc[3]), .F(n781) );
  MUX U794 ( .IN0(n781), .IN1(n778), .SEL(pc[4]), .F(n782) );
  MUX U795 ( .IN0(inst_mem_in_wire[716]), .IN1(inst_mem_in_wire[748]), .SEL(
        pc[2]), .F(n783) );
  MUX U796 ( .IN0(inst_mem_in_wire[652]), .IN1(inst_mem_in_wire[684]), .SEL(
        pc[2]), .F(n784) );
  MUX U797 ( .IN0(n784), .IN1(n783), .SEL(pc[3]), .F(n785) );
  MUX U798 ( .IN0(inst_mem_in_wire[588]), .IN1(inst_mem_in_wire[620]), .SEL(
        pc[2]), .F(n786) );
  MUX U799 ( .IN0(inst_mem_in_wire[524]), .IN1(inst_mem_in_wire[556]), .SEL(
        pc[2]), .F(n787) );
  MUX U800 ( .IN0(n787), .IN1(n786), .SEL(pc[3]), .F(n788) );
  MUX U801 ( .IN0(n788), .IN1(n785), .SEL(pc[4]), .F(n789) );
  MUX U802 ( .IN0(n789), .IN1(n782), .SEL(pc[5]), .F(n790) );
  MUX U803 ( .IN0(inst_mem_in_wire[460]), .IN1(inst_mem_in_wire[492]), .SEL(
        pc[2]), .F(n791) );
  MUX U804 ( .IN0(inst_mem_in_wire[396]), .IN1(inst_mem_in_wire[428]), .SEL(
        pc[2]), .F(n792) );
  MUX U805 ( .IN0(n792), .IN1(n791), .SEL(pc[3]), .F(n793) );
  MUX U806 ( .IN0(inst_mem_in_wire[332]), .IN1(inst_mem_in_wire[364]), .SEL(
        pc[2]), .F(n794) );
  MUX U807 ( .IN0(inst_mem_in_wire[268]), .IN1(inst_mem_in_wire[300]), .SEL(
        pc[2]), .F(n795) );
  MUX U808 ( .IN0(n795), .IN1(n794), .SEL(pc[3]), .F(n796) );
  MUX U809 ( .IN0(n796), .IN1(n793), .SEL(pc[4]), .F(n797) );
  MUX U810 ( .IN0(inst_mem_in_wire[204]), .IN1(inst_mem_in_wire[236]), .SEL(
        pc[2]), .F(n798) );
  MUX U811 ( .IN0(inst_mem_in_wire[140]), .IN1(inst_mem_in_wire[172]), .SEL(
        pc[2]), .F(n799) );
  MUX U812 ( .IN0(n799), .IN1(n798), .SEL(pc[3]), .F(n800) );
  MUX U813 ( .IN0(inst_mem_in_wire[76]), .IN1(inst_mem_in_wire[108]), .SEL(
        pc[2]), .F(n801) );
  MUX U814 ( .IN0(inst_mem_in_wire[12]), .IN1(inst_mem_in_wire[44]), .SEL(
        pc[2]), .F(n802) );
  MUX U815 ( .IN0(n802), .IN1(n801), .SEL(pc[3]), .F(n803) );
  MUX U816 ( .IN0(n803), .IN1(n800), .SEL(pc[4]), .F(n804) );
  MUX U817 ( .IN0(n804), .IN1(n797), .SEL(pc[5]), .F(n805) );
  MUX U818 ( .IN0(n805), .IN1(n790), .SEL(pc[6]), .F(n806) );
  MUX U819 ( .IN0(n806), .IN1(n775), .SEL(pc[7]), .F(opcode[12]) );
  MUX U820 ( .IN0(inst_mem_in_wire[1997]), .IN1(inst_mem_in_wire[2029]), .SEL(
        pc[2]), .F(n807) );
  MUX U821 ( .IN0(inst_mem_in_wire[1933]), .IN1(inst_mem_in_wire[1965]), .SEL(
        pc[2]), .F(n808) );
  MUX U822 ( .IN0(n808), .IN1(n807), .SEL(pc[3]), .F(n809) );
  MUX U823 ( .IN0(inst_mem_in_wire[1869]), .IN1(inst_mem_in_wire[1901]), .SEL(
        pc[2]), .F(n810) );
  MUX U824 ( .IN0(inst_mem_in_wire[1805]), .IN1(inst_mem_in_wire[1837]), .SEL(
        pc[2]), .F(n811) );
  MUX U825 ( .IN0(n811), .IN1(n810), .SEL(pc[3]), .F(n812) );
  MUX U826 ( .IN0(n812), .IN1(n809), .SEL(pc[4]), .F(n813) );
  MUX U827 ( .IN0(inst_mem_in_wire[1741]), .IN1(inst_mem_in_wire[1773]), .SEL(
        pc[2]), .F(n814) );
  MUX U828 ( .IN0(inst_mem_in_wire[1677]), .IN1(inst_mem_in_wire[1709]), .SEL(
        pc[2]), .F(n815) );
  MUX U829 ( .IN0(n815), .IN1(n814), .SEL(pc[3]), .F(n816) );
  MUX U830 ( .IN0(inst_mem_in_wire[1613]), .IN1(inst_mem_in_wire[1645]), .SEL(
        pc[2]), .F(n817) );
  MUX U831 ( .IN0(inst_mem_in_wire[1549]), .IN1(inst_mem_in_wire[1581]), .SEL(
        pc[2]), .F(n818) );
  MUX U832 ( .IN0(n818), .IN1(n817), .SEL(pc[3]), .F(n819) );
  MUX U833 ( .IN0(n819), .IN1(n816), .SEL(pc[4]), .F(n820) );
  MUX U834 ( .IN0(n820), .IN1(n813), .SEL(pc[5]), .F(n821) );
  MUX U835 ( .IN0(inst_mem_in_wire[1485]), .IN1(inst_mem_in_wire[1517]), .SEL(
        pc[2]), .F(n822) );
  MUX U836 ( .IN0(inst_mem_in_wire[1421]), .IN1(inst_mem_in_wire[1453]), .SEL(
        pc[2]), .F(n823) );
  MUX U837 ( .IN0(n823), .IN1(n822), .SEL(pc[3]), .F(n824) );
  MUX U838 ( .IN0(inst_mem_in_wire[1357]), .IN1(inst_mem_in_wire[1389]), .SEL(
        pc[2]), .F(n825) );
  MUX U839 ( .IN0(inst_mem_in_wire[1293]), .IN1(inst_mem_in_wire[1325]), .SEL(
        pc[2]), .F(n826) );
  MUX U840 ( .IN0(n826), .IN1(n825), .SEL(pc[3]), .F(n827) );
  MUX U841 ( .IN0(n827), .IN1(n824), .SEL(pc[4]), .F(n828) );
  MUX U842 ( .IN0(inst_mem_in_wire[1229]), .IN1(inst_mem_in_wire[1261]), .SEL(
        pc[2]), .F(n829) );
  MUX U843 ( .IN0(inst_mem_in_wire[1165]), .IN1(inst_mem_in_wire[1197]), .SEL(
        pc[2]), .F(n830) );
  MUX U844 ( .IN0(n830), .IN1(n829), .SEL(pc[3]), .F(n831) );
  MUX U845 ( .IN0(inst_mem_in_wire[1101]), .IN1(inst_mem_in_wire[1133]), .SEL(
        pc[2]), .F(n832) );
  MUX U846 ( .IN0(inst_mem_in_wire[1037]), .IN1(inst_mem_in_wire[1069]), .SEL(
        pc[2]), .F(n833) );
  MUX U847 ( .IN0(n833), .IN1(n832), .SEL(pc[3]), .F(n834) );
  MUX U848 ( .IN0(n834), .IN1(n831), .SEL(pc[4]), .F(n835) );
  MUX U849 ( .IN0(n835), .IN1(n828), .SEL(pc[5]), .F(n836) );
  MUX U850 ( .IN0(n836), .IN1(n821), .SEL(pc[6]), .F(n837) );
  MUX U851 ( .IN0(inst_mem_in_wire[973]), .IN1(inst_mem_in_wire[1005]), .SEL(
        pc[2]), .F(n838) );
  MUX U852 ( .IN0(inst_mem_in_wire[909]), .IN1(inst_mem_in_wire[941]), .SEL(
        pc[2]), .F(n839) );
  MUX U853 ( .IN0(n839), .IN1(n838), .SEL(pc[3]), .F(n840) );
  MUX U854 ( .IN0(inst_mem_in_wire[845]), .IN1(inst_mem_in_wire[877]), .SEL(
        pc[2]), .F(n841) );
  MUX U855 ( .IN0(inst_mem_in_wire[781]), .IN1(inst_mem_in_wire[813]), .SEL(
        pc[2]), .F(n842) );
  MUX U856 ( .IN0(n842), .IN1(n841), .SEL(pc[3]), .F(n843) );
  MUX U857 ( .IN0(n843), .IN1(n840), .SEL(pc[4]), .F(n844) );
  MUX U858 ( .IN0(inst_mem_in_wire[717]), .IN1(inst_mem_in_wire[749]), .SEL(
        pc[2]), .F(n845) );
  MUX U859 ( .IN0(inst_mem_in_wire[653]), .IN1(inst_mem_in_wire[685]), .SEL(
        pc[2]), .F(n846) );
  MUX U860 ( .IN0(n846), .IN1(n845), .SEL(pc[3]), .F(n847) );
  MUX U861 ( .IN0(inst_mem_in_wire[589]), .IN1(inst_mem_in_wire[621]), .SEL(
        pc[2]), .F(n848) );
  MUX U862 ( .IN0(inst_mem_in_wire[525]), .IN1(inst_mem_in_wire[557]), .SEL(
        pc[2]), .F(n849) );
  MUX U863 ( .IN0(n849), .IN1(n848), .SEL(pc[3]), .F(n850) );
  MUX U864 ( .IN0(n850), .IN1(n847), .SEL(pc[4]), .F(n851) );
  MUX U865 ( .IN0(n851), .IN1(n844), .SEL(pc[5]), .F(n852) );
  MUX U866 ( .IN0(inst_mem_in_wire[461]), .IN1(inst_mem_in_wire[493]), .SEL(
        pc[2]), .F(n853) );
  MUX U867 ( .IN0(inst_mem_in_wire[397]), .IN1(inst_mem_in_wire[429]), .SEL(
        pc[2]), .F(n854) );
  MUX U868 ( .IN0(n854), .IN1(n853), .SEL(pc[3]), .F(n855) );
  MUX U869 ( .IN0(inst_mem_in_wire[333]), .IN1(inst_mem_in_wire[365]), .SEL(
        pc[2]), .F(n856) );
  MUX U870 ( .IN0(inst_mem_in_wire[269]), .IN1(inst_mem_in_wire[301]), .SEL(
        pc[2]), .F(n857) );
  MUX U871 ( .IN0(n857), .IN1(n856), .SEL(pc[3]), .F(n858) );
  MUX U872 ( .IN0(n858), .IN1(n855), .SEL(pc[4]), .F(n859) );
  MUX U873 ( .IN0(inst_mem_in_wire[205]), .IN1(inst_mem_in_wire[237]), .SEL(
        pc[2]), .F(n860) );
  MUX U874 ( .IN0(inst_mem_in_wire[141]), .IN1(inst_mem_in_wire[173]), .SEL(
        pc[2]), .F(n861) );
  MUX U875 ( .IN0(n861), .IN1(n860), .SEL(pc[3]), .F(n862) );
  MUX U876 ( .IN0(inst_mem_in_wire[77]), .IN1(inst_mem_in_wire[109]), .SEL(
        pc[2]), .F(n863) );
  MUX U877 ( .IN0(inst_mem_in_wire[13]), .IN1(inst_mem_in_wire[45]), .SEL(
        pc[2]), .F(n864) );
  MUX U878 ( .IN0(n864), .IN1(n863), .SEL(pc[3]), .F(n865) );
  MUX U879 ( .IN0(n865), .IN1(n862), .SEL(pc[4]), .F(n866) );
  MUX U880 ( .IN0(n866), .IN1(n859), .SEL(pc[5]), .F(n867) );
  MUX U881 ( .IN0(n867), .IN1(n852), .SEL(pc[6]), .F(n868) );
  MUX U882 ( .IN0(n868), .IN1(n837), .SEL(pc[7]), .F(opcode[13]) );
  MUX U883 ( .IN0(inst_mem_in_wire[1998]), .IN1(inst_mem_in_wire[2030]), .SEL(
        pc[2]), .F(n869) );
  MUX U884 ( .IN0(inst_mem_in_wire[1934]), .IN1(inst_mem_in_wire[1966]), .SEL(
        pc[2]), .F(n870) );
  MUX U885 ( .IN0(n870), .IN1(n869), .SEL(pc[3]), .F(n871) );
  MUX U886 ( .IN0(inst_mem_in_wire[1870]), .IN1(inst_mem_in_wire[1902]), .SEL(
        pc[2]), .F(n872) );
  MUX U887 ( .IN0(inst_mem_in_wire[1806]), .IN1(inst_mem_in_wire[1838]), .SEL(
        pc[2]), .F(n873) );
  MUX U888 ( .IN0(n873), .IN1(n872), .SEL(pc[3]), .F(n874) );
  MUX U889 ( .IN0(n874), .IN1(n871), .SEL(pc[4]), .F(n875) );
  MUX U890 ( .IN0(inst_mem_in_wire[1742]), .IN1(inst_mem_in_wire[1774]), .SEL(
        pc[2]), .F(n876) );
  MUX U891 ( .IN0(inst_mem_in_wire[1678]), .IN1(inst_mem_in_wire[1710]), .SEL(
        pc[2]), .F(n877) );
  MUX U892 ( .IN0(n877), .IN1(n876), .SEL(pc[3]), .F(n878) );
  MUX U893 ( .IN0(inst_mem_in_wire[1614]), .IN1(inst_mem_in_wire[1646]), .SEL(
        pc[2]), .F(n879) );
  MUX U894 ( .IN0(inst_mem_in_wire[1550]), .IN1(inst_mem_in_wire[1582]), .SEL(
        pc[2]), .F(n880) );
  MUX U895 ( .IN0(n880), .IN1(n879), .SEL(pc[3]), .F(n881) );
  MUX U896 ( .IN0(n881), .IN1(n878), .SEL(pc[4]), .F(n882) );
  MUX U897 ( .IN0(n882), .IN1(n875), .SEL(pc[5]), .F(n883) );
  MUX U898 ( .IN0(inst_mem_in_wire[1486]), .IN1(inst_mem_in_wire[1518]), .SEL(
        pc[2]), .F(n884) );
  MUX U899 ( .IN0(inst_mem_in_wire[1422]), .IN1(inst_mem_in_wire[1454]), .SEL(
        pc[2]), .F(n885) );
  MUX U900 ( .IN0(n885), .IN1(n884), .SEL(pc[3]), .F(n886) );
  MUX U901 ( .IN0(inst_mem_in_wire[1358]), .IN1(inst_mem_in_wire[1390]), .SEL(
        pc[2]), .F(n887) );
  MUX U902 ( .IN0(inst_mem_in_wire[1294]), .IN1(inst_mem_in_wire[1326]), .SEL(
        pc[2]), .F(n888) );
  MUX U903 ( .IN0(n888), .IN1(n887), .SEL(pc[3]), .F(n889) );
  MUX U904 ( .IN0(n889), .IN1(n886), .SEL(pc[4]), .F(n890) );
  MUX U905 ( .IN0(inst_mem_in_wire[1230]), .IN1(inst_mem_in_wire[1262]), .SEL(
        pc[2]), .F(n891) );
  MUX U906 ( .IN0(inst_mem_in_wire[1166]), .IN1(inst_mem_in_wire[1198]), .SEL(
        pc[2]), .F(n892) );
  MUX U907 ( .IN0(n892), .IN1(n891), .SEL(pc[3]), .F(n893) );
  MUX U908 ( .IN0(inst_mem_in_wire[1102]), .IN1(inst_mem_in_wire[1134]), .SEL(
        pc[2]), .F(n894) );
  MUX U909 ( .IN0(inst_mem_in_wire[1038]), .IN1(inst_mem_in_wire[1070]), .SEL(
        pc[2]), .F(n895) );
  MUX U910 ( .IN0(n895), .IN1(n894), .SEL(pc[3]), .F(n896) );
  MUX U911 ( .IN0(n896), .IN1(n893), .SEL(pc[4]), .F(n897) );
  MUX U912 ( .IN0(n897), .IN1(n890), .SEL(pc[5]), .F(n898) );
  MUX U913 ( .IN0(n898), .IN1(n883), .SEL(pc[6]), .F(n899) );
  MUX U914 ( .IN0(inst_mem_in_wire[974]), .IN1(inst_mem_in_wire[1006]), .SEL(
        pc[2]), .F(n900) );
  MUX U915 ( .IN0(inst_mem_in_wire[910]), .IN1(inst_mem_in_wire[942]), .SEL(
        pc[2]), .F(n901) );
  MUX U916 ( .IN0(n901), .IN1(n900), .SEL(pc[3]), .F(n902) );
  MUX U917 ( .IN0(inst_mem_in_wire[846]), .IN1(inst_mem_in_wire[878]), .SEL(
        pc[2]), .F(n903) );
  MUX U918 ( .IN0(inst_mem_in_wire[782]), .IN1(inst_mem_in_wire[814]), .SEL(
        pc[2]), .F(n904) );
  MUX U919 ( .IN0(n904), .IN1(n903), .SEL(pc[3]), .F(n905) );
  MUX U920 ( .IN0(n905), .IN1(n902), .SEL(pc[4]), .F(n906) );
  MUX U921 ( .IN0(inst_mem_in_wire[718]), .IN1(inst_mem_in_wire[750]), .SEL(
        pc[2]), .F(n907) );
  MUX U922 ( .IN0(inst_mem_in_wire[654]), .IN1(inst_mem_in_wire[686]), .SEL(
        pc[2]), .F(n908) );
  MUX U923 ( .IN0(n908), .IN1(n907), .SEL(pc[3]), .F(n909) );
  MUX U924 ( .IN0(inst_mem_in_wire[590]), .IN1(inst_mem_in_wire[622]), .SEL(
        pc[2]), .F(n910) );
  MUX U925 ( .IN0(inst_mem_in_wire[526]), .IN1(inst_mem_in_wire[558]), .SEL(
        pc[2]), .F(n911) );
  MUX U926 ( .IN0(n911), .IN1(n910), .SEL(pc[3]), .F(n912) );
  MUX U927 ( .IN0(n912), .IN1(n909), .SEL(pc[4]), .F(n913) );
  MUX U928 ( .IN0(n913), .IN1(n906), .SEL(pc[5]), .F(n914) );
  MUX U929 ( .IN0(inst_mem_in_wire[462]), .IN1(inst_mem_in_wire[494]), .SEL(
        pc[2]), .F(n915) );
  MUX U930 ( .IN0(inst_mem_in_wire[398]), .IN1(inst_mem_in_wire[430]), .SEL(
        pc[2]), .F(n916) );
  MUX U931 ( .IN0(n916), .IN1(n915), .SEL(pc[3]), .F(n917) );
  MUX U932 ( .IN0(inst_mem_in_wire[334]), .IN1(inst_mem_in_wire[366]), .SEL(
        pc[2]), .F(n918) );
  MUX U933 ( .IN0(inst_mem_in_wire[270]), .IN1(inst_mem_in_wire[302]), .SEL(
        pc[2]), .F(n919) );
  MUX U934 ( .IN0(n919), .IN1(n918), .SEL(pc[3]), .F(n920) );
  MUX U935 ( .IN0(n920), .IN1(n917), .SEL(pc[4]), .F(n921) );
  MUX U936 ( .IN0(inst_mem_in_wire[206]), .IN1(inst_mem_in_wire[238]), .SEL(
        pc[2]), .F(n922) );
  MUX U937 ( .IN0(inst_mem_in_wire[142]), .IN1(inst_mem_in_wire[174]), .SEL(
        pc[2]), .F(n923) );
  MUX U938 ( .IN0(n923), .IN1(n922), .SEL(pc[3]), .F(n924) );
  MUX U939 ( .IN0(inst_mem_in_wire[78]), .IN1(inst_mem_in_wire[110]), .SEL(
        pc[2]), .F(n925) );
  MUX U940 ( .IN0(inst_mem_in_wire[14]), .IN1(inst_mem_in_wire[46]), .SEL(
        pc[2]), .F(n926) );
  MUX U941 ( .IN0(n926), .IN1(n925), .SEL(pc[3]), .F(n927) );
  MUX U942 ( .IN0(n927), .IN1(n924), .SEL(pc[4]), .F(n928) );
  MUX U943 ( .IN0(n928), .IN1(n921), .SEL(pc[5]), .F(n929) );
  MUX U944 ( .IN0(n929), .IN1(n914), .SEL(pc[6]), .F(n930) );
  MUX U945 ( .IN0(n930), .IN1(n899), .SEL(pc[7]), .F(opcode[14]) );
  MUX U946 ( .IN0(inst_mem_in_wire[1999]), .IN1(inst_mem_in_wire[2031]), .SEL(
        pc[2]), .F(n931) );
  MUX U947 ( .IN0(inst_mem_in_wire[1935]), .IN1(inst_mem_in_wire[1967]), .SEL(
        pc[2]), .F(n932) );
  MUX U948 ( .IN0(n932), .IN1(n931), .SEL(pc[3]), .F(n933) );
  MUX U949 ( .IN0(inst_mem_in_wire[1871]), .IN1(inst_mem_in_wire[1903]), .SEL(
        pc[2]), .F(n934) );
  MUX U950 ( .IN0(inst_mem_in_wire[1807]), .IN1(inst_mem_in_wire[1839]), .SEL(
        pc[2]), .F(n935) );
  MUX U951 ( .IN0(n935), .IN1(n934), .SEL(pc[3]), .F(n936) );
  MUX U952 ( .IN0(n936), .IN1(n933), .SEL(pc[4]), .F(n937) );
  MUX U953 ( .IN0(inst_mem_in_wire[1743]), .IN1(inst_mem_in_wire[1775]), .SEL(
        pc[2]), .F(n938) );
  MUX U954 ( .IN0(inst_mem_in_wire[1679]), .IN1(inst_mem_in_wire[1711]), .SEL(
        pc[2]), .F(n939) );
  MUX U955 ( .IN0(n939), .IN1(n938), .SEL(pc[3]), .F(n940) );
  MUX U956 ( .IN0(inst_mem_in_wire[1615]), .IN1(inst_mem_in_wire[1647]), .SEL(
        pc[2]), .F(n941) );
  MUX U957 ( .IN0(inst_mem_in_wire[1551]), .IN1(inst_mem_in_wire[1583]), .SEL(
        pc[2]), .F(n942) );
  MUX U958 ( .IN0(n942), .IN1(n941), .SEL(pc[3]), .F(n943) );
  MUX U959 ( .IN0(n943), .IN1(n940), .SEL(pc[4]), .F(n944) );
  MUX U960 ( .IN0(n944), .IN1(n937), .SEL(pc[5]), .F(n945) );
  MUX U961 ( .IN0(inst_mem_in_wire[1487]), .IN1(inst_mem_in_wire[1519]), .SEL(
        pc[2]), .F(n946) );
  MUX U962 ( .IN0(inst_mem_in_wire[1423]), .IN1(inst_mem_in_wire[1455]), .SEL(
        pc[2]), .F(n947) );
  MUX U963 ( .IN0(n947), .IN1(n946), .SEL(pc[3]), .F(n948) );
  MUX U964 ( .IN0(inst_mem_in_wire[1359]), .IN1(inst_mem_in_wire[1391]), .SEL(
        pc[2]), .F(n949) );
  MUX U965 ( .IN0(inst_mem_in_wire[1295]), .IN1(inst_mem_in_wire[1327]), .SEL(
        pc[2]), .F(n950) );
  MUX U966 ( .IN0(n950), .IN1(n949), .SEL(pc[3]), .F(n951) );
  MUX U967 ( .IN0(n951), .IN1(n948), .SEL(pc[4]), .F(n952) );
  MUX U968 ( .IN0(inst_mem_in_wire[1231]), .IN1(inst_mem_in_wire[1263]), .SEL(
        pc[2]), .F(n953) );
  MUX U969 ( .IN0(inst_mem_in_wire[1167]), .IN1(inst_mem_in_wire[1199]), .SEL(
        pc[2]), .F(n954) );
  MUX U970 ( .IN0(n954), .IN1(n953), .SEL(pc[3]), .F(n955) );
  MUX U971 ( .IN0(inst_mem_in_wire[1103]), .IN1(inst_mem_in_wire[1135]), .SEL(
        pc[2]), .F(n956) );
  MUX U972 ( .IN0(inst_mem_in_wire[1039]), .IN1(inst_mem_in_wire[1071]), .SEL(
        pc[2]), .F(n957) );
  MUX U973 ( .IN0(n957), .IN1(n956), .SEL(pc[3]), .F(n958) );
  MUX U974 ( .IN0(n958), .IN1(n955), .SEL(pc[4]), .F(n959) );
  MUX U975 ( .IN0(n959), .IN1(n952), .SEL(pc[5]), .F(n960) );
  MUX U976 ( .IN0(n960), .IN1(n945), .SEL(pc[6]), .F(n961) );
  MUX U977 ( .IN0(inst_mem_in_wire[975]), .IN1(inst_mem_in_wire[1007]), .SEL(
        pc[2]), .F(n962) );
  MUX U978 ( .IN0(inst_mem_in_wire[911]), .IN1(inst_mem_in_wire[943]), .SEL(
        pc[2]), .F(n963) );
  MUX U979 ( .IN0(n963), .IN1(n962), .SEL(pc[3]), .F(n964) );
  MUX U980 ( .IN0(inst_mem_in_wire[847]), .IN1(inst_mem_in_wire[879]), .SEL(
        pc[2]), .F(n965) );
  MUX U981 ( .IN0(inst_mem_in_wire[783]), .IN1(inst_mem_in_wire[815]), .SEL(
        pc[2]), .F(n966) );
  MUX U982 ( .IN0(n966), .IN1(n965), .SEL(pc[3]), .F(n967) );
  MUX U983 ( .IN0(n967), .IN1(n964), .SEL(pc[4]), .F(n968) );
  MUX U984 ( .IN0(inst_mem_in_wire[719]), .IN1(inst_mem_in_wire[751]), .SEL(
        pc[2]), .F(n969) );
  MUX U985 ( .IN0(inst_mem_in_wire[655]), .IN1(inst_mem_in_wire[687]), .SEL(
        pc[2]), .F(n970) );
  MUX U986 ( .IN0(n970), .IN1(n969), .SEL(pc[3]), .F(n971) );
  MUX U987 ( .IN0(inst_mem_in_wire[591]), .IN1(inst_mem_in_wire[623]), .SEL(
        pc[2]), .F(n972) );
  MUX U988 ( .IN0(inst_mem_in_wire[527]), .IN1(inst_mem_in_wire[559]), .SEL(
        pc[2]), .F(n973) );
  MUX U989 ( .IN0(n973), .IN1(n972), .SEL(pc[3]), .F(n974) );
  MUX U990 ( .IN0(n974), .IN1(n971), .SEL(pc[4]), .F(n975) );
  MUX U991 ( .IN0(n975), .IN1(n968), .SEL(pc[5]), .F(n976) );
  MUX U992 ( .IN0(inst_mem_in_wire[463]), .IN1(inst_mem_in_wire[495]), .SEL(
        pc[2]), .F(n977) );
  MUX U993 ( .IN0(inst_mem_in_wire[399]), .IN1(inst_mem_in_wire[431]), .SEL(
        pc[2]), .F(n978) );
  MUX U994 ( .IN0(n978), .IN1(n977), .SEL(pc[3]), .F(n979) );
  MUX U995 ( .IN0(inst_mem_in_wire[335]), .IN1(inst_mem_in_wire[367]), .SEL(
        pc[2]), .F(n980) );
  MUX U996 ( .IN0(inst_mem_in_wire[271]), .IN1(inst_mem_in_wire[303]), .SEL(
        pc[2]), .F(n981) );
  MUX U997 ( .IN0(n981), .IN1(n980), .SEL(pc[3]), .F(n982) );
  MUX U998 ( .IN0(n982), .IN1(n979), .SEL(pc[4]), .F(n983) );
  MUX U999 ( .IN0(inst_mem_in_wire[207]), .IN1(inst_mem_in_wire[239]), .SEL(
        pc[2]), .F(n984) );
  MUX U1000 ( .IN0(inst_mem_in_wire[143]), .IN1(inst_mem_in_wire[175]), .SEL(
        pc[2]), .F(n985) );
  MUX U1001 ( .IN0(n985), .IN1(n984), .SEL(pc[3]), .F(n986) );
  MUX U1002 ( .IN0(inst_mem_in_wire[79]), .IN1(inst_mem_in_wire[111]), .SEL(
        pc[2]), .F(n987) );
  MUX U1003 ( .IN0(inst_mem_in_wire[15]), .IN1(inst_mem_in_wire[47]), .SEL(
        pc[2]), .F(n988) );
  MUX U1004 ( .IN0(n988), .IN1(n987), .SEL(pc[3]), .F(n989) );
  MUX U1005 ( .IN0(n989), .IN1(n986), .SEL(pc[4]), .F(n990) );
  MUX U1006 ( .IN0(n990), .IN1(n983), .SEL(pc[5]), .F(n991) );
  MUX U1007 ( .IN0(n991), .IN1(n976), .SEL(pc[6]), .F(n992) );
  MUX U1008 ( .IN0(n992), .IN1(n961), .SEL(pc[7]), .F(opcode[15]) );
  MUX U1009 ( .IN0(inst_mem_in_wire[2000]), .IN1(inst_mem_in_wire[2032]), 
        .SEL(pc[2]), .F(n993) );
  MUX U1010 ( .IN0(inst_mem_in_wire[1936]), .IN1(inst_mem_in_wire[1968]), 
        .SEL(pc[2]), .F(n994) );
  MUX U1011 ( .IN0(n994), .IN1(n993), .SEL(pc[3]), .F(n995) );
  MUX U1012 ( .IN0(inst_mem_in_wire[1872]), .IN1(inst_mem_in_wire[1904]), 
        .SEL(pc[2]), .F(n996) );
  MUX U1013 ( .IN0(inst_mem_in_wire[1808]), .IN1(inst_mem_in_wire[1840]), 
        .SEL(pc[2]), .F(n997) );
  MUX U1014 ( .IN0(n997), .IN1(n996), .SEL(pc[3]), .F(n998) );
  MUX U1015 ( .IN0(n998), .IN1(n995), .SEL(pc[4]), .F(n999) );
  MUX U1016 ( .IN0(inst_mem_in_wire[1744]), .IN1(inst_mem_in_wire[1776]), 
        .SEL(pc[2]), .F(n1000) );
  MUX U1017 ( .IN0(inst_mem_in_wire[1680]), .IN1(inst_mem_in_wire[1712]), 
        .SEL(pc[2]), .F(n1001) );
  MUX U1018 ( .IN0(n1001), .IN1(n1000), .SEL(pc[3]), .F(n1002) );
  MUX U1019 ( .IN0(inst_mem_in_wire[1616]), .IN1(inst_mem_in_wire[1648]), 
        .SEL(pc[2]), .F(n1003) );
  MUX U1020 ( .IN0(inst_mem_in_wire[1552]), .IN1(inst_mem_in_wire[1584]), 
        .SEL(pc[2]), .F(n1004) );
  MUX U1021 ( .IN0(n1004), .IN1(n1003), .SEL(pc[3]), .F(n1005) );
  MUX U1022 ( .IN0(n1005), .IN1(n1002), .SEL(pc[4]), .F(n1006) );
  MUX U1023 ( .IN0(n1006), .IN1(n999), .SEL(pc[5]), .F(n1007) );
  MUX U1024 ( .IN0(inst_mem_in_wire[1488]), .IN1(inst_mem_in_wire[1520]), 
        .SEL(pc[2]), .F(n1008) );
  MUX U1025 ( .IN0(inst_mem_in_wire[1424]), .IN1(inst_mem_in_wire[1456]), 
        .SEL(pc[2]), .F(n1009) );
  MUX U1026 ( .IN0(n1009), .IN1(n1008), .SEL(pc[3]), .F(n1010) );
  MUX U1027 ( .IN0(inst_mem_in_wire[1360]), .IN1(inst_mem_in_wire[1392]), 
        .SEL(pc[2]), .F(n1011) );
  MUX U1028 ( .IN0(inst_mem_in_wire[1296]), .IN1(inst_mem_in_wire[1328]), 
        .SEL(pc[2]), .F(n1012) );
  MUX U1029 ( .IN0(n1012), .IN1(n1011), .SEL(pc[3]), .F(n1013) );
  MUX U1030 ( .IN0(n1013), .IN1(n1010), .SEL(pc[4]), .F(n1014) );
  MUX U1031 ( .IN0(inst_mem_in_wire[1232]), .IN1(inst_mem_in_wire[1264]), 
        .SEL(pc[2]), .F(n1015) );
  MUX U1032 ( .IN0(inst_mem_in_wire[1168]), .IN1(inst_mem_in_wire[1200]), 
        .SEL(pc[2]), .F(n1016) );
  MUX U1033 ( .IN0(n1016), .IN1(n1015), .SEL(pc[3]), .F(n1017) );
  MUX U1034 ( .IN0(inst_mem_in_wire[1104]), .IN1(inst_mem_in_wire[1136]), 
        .SEL(pc[2]), .F(n1018) );
  MUX U1035 ( .IN0(inst_mem_in_wire[1040]), .IN1(inst_mem_in_wire[1072]), 
        .SEL(pc[2]), .F(n1019) );
  MUX U1036 ( .IN0(n1019), .IN1(n1018), .SEL(pc[3]), .F(n1020) );
  MUX U1037 ( .IN0(n1020), .IN1(n1017), .SEL(pc[4]), .F(n1021) );
  MUX U1038 ( .IN0(n1021), .IN1(n1014), .SEL(pc[5]), .F(n1022) );
  MUX U1039 ( .IN0(n1022), .IN1(n1007), .SEL(pc[6]), .F(n1023) );
  MUX U1040 ( .IN0(inst_mem_in_wire[976]), .IN1(inst_mem_in_wire[1008]), .SEL(
        pc[2]), .F(n1024) );
  MUX U1041 ( .IN0(inst_mem_in_wire[912]), .IN1(inst_mem_in_wire[944]), .SEL(
        pc[2]), .F(n1025) );
  MUX U1042 ( .IN0(n1025), .IN1(n1024), .SEL(pc[3]), .F(n1026) );
  MUX U1043 ( .IN0(inst_mem_in_wire[848]), .IN1(inst_mem_in_wire[880]), .SEL(
        pc[2]), .F(n1027) );
  MUX U1044 ( .IN0(inst_mem_in_wire[784]), .IN1(inst_mem_in_wire[816]), .SEL(
        pc[2]), .F(n1028) );
  MUX U1045 ( .IN0(n1028), .IN1(n1027), .SEL(pc[3]), .F(n1029) );
  MUX U1046 ( .IN0(n1029), .IN1(n1026), .SEL(pc[4]), .F(n1030) );
  MUX U1047 ( .IN0(inst_mem_in_wire[720]), .IN1(inst_mem_in_wire[752]), .SEL(
        pc[2]), .F(n1031) );
  MUX U1048 ( .IN0(inst_mem_in_wire[656]), .IN1(inst_mem_in_wire[688]), .SEL(
        pc[2]), .F(n1032) );
  MUX U1049 ( .IN0(n1032), .IN1(n1031), .SEL(pc[3]), .F(n1033) );
  MUX U1050 ( .IN0(inst_mem_in_wire[592]), .IN1(inst_mem_in_wire[624]), .SEL(
        pc[2]), .F(n1034) );
  MUX U1051 ( .IN0(inst_mem_in_wire[528]), .IN1(inst_mem_in_wire[560]), .SEL(
        pc[2]), .F(n1035) );
  MUX U1052 ( .IN0(n1035), .IN1(n1034), .SEL(pc[3]), .F(n1036) );
  MUX U1053 ( .IN0(n1036), .IN1(n1033), .SEL(pc[4]), .F(n1037) );
  MUX U1054 ( .IN0(n1037), .IN1(n1030), .SEL(pc[5]), .F(n1038) );
  MUX U1055 ( .IN0(inst_mem_in_wire[464]), .IN1(inst_mem_in_wire[496]), .SEL(
        pc[2]), .F(n1039) );
  MUX U1056 ( .IN0(inst_mem_in_wire[400]), .IN1(inst_mem_in_wire[432]), .SEL(
        pc[2]), .F(n1040) );
  MUX U1057 ( .IN0(n1040), .IN1(n1039), .SEL(pc[3]), .F(n1041) );
  MUX U1058 ( .IN0(inst_mem_in_wire[336]), .IN1(inst_mem_in_wire[368]), .SEL(
        pc[2]), .F(n1042) );
  MUX U1059 ( .IN0(inst_mem_in_wire[272]), .IN1(inst_mem_in_wire[304]), .SEL(
        pc[2]), .F(n1043) );
  MUX U1060 ( .IN0(n1043), .IN1(n1042), .SEL(pc[3]), .F(n1044) );
  MUX U1061 ( .IN0(n1044), .IN1(n1041), .SEL(pc[4]), .F(n1045) );
  MUX U1062 ( .IN0(inst_mem_in_wire[208]), .IN1(inst_mem_in_wire[240]), .SEL(
        pc[2]), .F(n1046) );
  MUX U1063 ( .IN0(inst_mem_in_wire[144]), .IN1(inst_mem_in_wire[176]), .SEL(
        pc[2]), .F(n1047) );
  MUX U1064 ( .IN0(n1047), .IN1(n1046), .SEL(pc[3]), .F(n1048) );
  MUX U1065 ( .IN0(inst_mem_in_wire[80]), .IN1(inst_mem_in_wire[112]), .SEL(
        pc[2]), .F(n1049) );
  MUX U1066 ( .IN0(inst_mem_in_wire[16]), .IN1(inst_mem_in_wire[48]), .SEL(
        pc[2]), .F(n1050) );
  MUX U1067 ( .IN0(n1050), .IN1(n1049), .SEL(pc[3]), .F(n1051) );
  MUX U1068 ( .IN0(n1051), .IN1(n1048), .SEL(pc[4]), .F(n1052) );
  MUX U1069 ( .IN0(n1052), .IN1(n1045), .SEL(pc[5]), .F(n1053) );
  MUX U1070 ( .IN0(n1053), .IN1(n1038), .SEL(pc[6]), .F(n1054) );
  MUX U1071 ( .IN0(n1054), .IN1(n1023), .SEL(pc[7]), .F(opcode[16]) );
  MUX U1072 ( .IN0(inst_mem_in_wire[2001]), .IN1(inst_mem_in_wire[2033]), 
        .SEL(pc[2]), .F(n1055) );
  MUX U1073 ( .IN0(inst_mem_in_wire[1937]), .IN1(inst_mem_in_wire[1969]), 
        .SEL(pc[2]), .F(n1056) );
  MUX U1074 ( .IN0(n1056), .IN1(n1055), .SEL(pc[3]), .F(n1057) );
  MUX U1075 ( .IN0(inst_mem_in_wire[1873]), .IN1(inst_mem_in_wire[1905]), 
        .SEL(pc[2]), .F(n1058) );
  MUX U1076 ( .IN0(inst_mem_in_wire[1809]), .IN1(inst_mem_in_wire[1841]), 
        .SEL(pc[2]), .F(n1059) );
  MUX U1077 ( .IN0(n1059), .IN1(n1058), .SEL(pc[3]), .F(n1060) );
  MUX U1078 ( .IN0(n1060), .IN1(n1057), .SEL(pc[4]), .F(n1061) );
  MUX U1079 ( .IN0(inst_mem_in_wire[1745]), .IN1(inst_mem_in_wire[1777]), 
        .SEL(pc[2]), .F(n1062) );
  MUX U1080 ( .IN0(inst_mem_in_wire[1681]), .IN1(inst_mem_in_wire[1713]), 
        .SEL(pc[2]), .F(n1063) );
  MUX U1081 ( .IN0(n1063), .IN1(n1062), .SEL(pc[3]), .F(n1064) );
  MUX U1082 ( .IN0(inst_mem_in_wire[1617]), .IN1(inst_mem_in_wire[1649]), 
        .SEL(pc[2]), .F(n1065) );
  MUX U1083 ( .IN0(inst_mem_in_wire[1553]), .IN1(inst_mem_in_wire[1585]), 
        .SEL(pc[2]), .F(n1066) );
  MUX U1084 ( .IN0(n1066), .IN1(n1065), .SEL(pc[3]), .F(n1067) );
  MUX U1085 ( .IN0(n1067), .IN1(n1064), .SEL(pc[4]), .F(n1068) );
  MUX U1086 ( .IN0(n1068), .IN1(n1061), .SEL(pc[5]), .F(n1069) );
  MUX U1087 ( .IN0(inst_mem_in_wire[1489]), .IN1(inst_mem_in_wire[1521]), 
        .SEL(pc[2]), .F(n1070) );
  MUX U1088 ( .IN0(inst_mem_in_wire[1425]), .IN1(inst_mem_in_wire[1457]), 
        .SEL(pc[2]), .F(n1071) );
  MUX U1089 ( .IN0(n1071), .IN1(n1070), .SEL(pc[3]), .F(n1072) );
  MUX U1090 ( .IN0(inst_mem_in_wire[1361]), .IN1(inst_mem_in_wire[1393]), 
        .SEL(pc[2]), .F(n1073) );
  MUX U1091 ( .IN0(inst_mem_in_wire[1297]), .IN1(inst_mem_in_wire[1329]), 
        .SEL(pc[2]), .F(n1074) );
  MUX U1092 ( .IN0(n1074), .IN1(n1073), .SEL(pc[3]), .F(n1075) );
  MUX U1093 ( .IN0(n1075), .IN1(n1072), .SEL(pc[4]), .F(n1076) );
  MUX U1094 ( .IN0(inst_mem_in_wire[1233]), .IN1(inst_mem_in_wire[1265]), 
        .SEL(pc[2]), .F(n1077) );
  MUX U1095 ( .IN0(inst_mem_in_wire[1169]), .IN1(inst_mem_in_wire[1201]), 
        .SEL(pc[2]), .F(n1078) );
  MUX U1096 ( .IN0(n1078), .IN1(n1077), .SEL(pc[3]), .F(n1079) );
  MUX U1097 ( .IN0(inst_mem_in_wire[1105]), .IN1(inst_mem_in_wire[1137]), 
        .SEL(pc[2]), .F(n1080) );
  MUX U1098 ( .IN0(inst_mem_in_wire[1041]), .IN1(inst_mem_in_wire[1073]), 
        .SEL(pc[2]), .F(n1081) );
  MUX U1099 ( .IN0(n1081), .IN1(n1080), .SEL(pc[3]), .F(n1082) );
  MUX U1100 ( .IN0(n1082), .IN1(n1079), .SEL(pc[4]), .F(n1083) );
  MUX U1101 ( .IN0(n1083), .IN1(n1076), .SEL(pc[5]), .F(n1084) );
  MUX U1102 ( .IN0(n1084), .IN1(n1069), .SEL(pc[6]), .F(n1085) );
  MUX U1103 ( .IN0(inst_mem_in_wire[977]), .IN1(inst_mem_in_wire[1009]), .SEL(
        pc[2]), .F(n1086) );
  MUX U1104 ( .IN0(inst_mem_in_wire[913]), .IN1(inst_mem_in_wire[945]), .SEL(
        pc[2]), .F(n1087) );
  MUX U1105 ( .IN0(n1087), .IN1(n1086), .SEL(pc[3]), .F(n1088) );
  MUX U1106 ( .IN0(inst_mem_in_wire[849]), .IN1(inst_mem_in_wire[881]), .SEL(
        pc[2]), .F(n1089) );
  MUX U1107 ( .IN0(inst_mem_in_wire[785]), .IN1(inst_mem_in_wire[817]), .SEL(
        pc[2]), .F(n1090) );
  MUX U1108 ( .IN0(n1090), .IN1(n1089), .SEL(pc[3]), .F(n1091) );
  MUX U1109 ( .IN0(n1091), .IN1(n1088), .SEL(pc[4]), .F(n1092) );
  MUX U1110 ( .IN0(inst_mem_in_wire[721]), .IN1(inst_mem_in_wire[753]), .SEL(
        pc[2]), .F(n1093) );
  MUX U1111 ( .IN0(inst_mem_in_wire[657]), .IN1(inst_mem_in_wire[689]), .SEL(
        pc[2]), .F(n1094) );
  MUX U1112 ( .IN0(n1094), .IN1(n1093), .SEL(pc[3]), .F(n1095) );
  MUX U1113 ( .IN0(inst_mem_in_wire[593]), .IN1(inst_mem_in_wire[625]), .SEL(
        pc[2]), .F(n1096) );
  MUX U1114 ( .IN0(inst_mem_in_wire[529]), .IN1(inst_mem_in_wire[561]), .SEL(
        pc[2]), .F(n1097) );
  MUX U1115 ( .IN0(n1097), .IN1(n1096), .SEL(pc[3]), .F(n1098) );
  MUX U1116 ( .IN0(n1098), .IN1(n1095), .SEL(pc[4]), .F(n1099) );
  MUX U1117 ( .IN0(n1099), .IN1(n1092), .SEL(pc[5]), .F(n1100) );
  MUX U1118 ( .IN0(inst_mem_in_wire[465]), .IN1(inst_mem_in_wire[497]), .SEL(
        pc[2]), .F(n1101) );
  MUX U1119 ( .IN0(inst_mem_in_wire[401]), .IN1(inst_mem_in_wire[433]), .SEL(
        pc[2]), .F(n1102) );
  MUX U1120 ( .IN0(n1102), .IN1(n1101), .SEL(pc[3]), .F(n1103) );
  MUX U1121 ( .IN0(inst_mem_in_wire[337]), .IN1(inst_mem_in_wire[369]), .SEL(
        pc[2]), .F(n1104) );
  MUX U1122 ( .IN0(inst_mem_in_wire[273]), .IN1(inst_mem_in_wire[305]), .SEL(
        pc[2]), .F(n1105) );
  MUX U1123 ( .IN0(n1105), .IN1(n1104), .SEL(pc[3]), .F(n1106) );
  MUX U1124 ( .IN0(n1106), .IN1(n1103), .SEL(pc[4]), .F(n1107) );
  MUX U1125 ( .IN0(inst_mem_in_wire[209]), .IN1(inst_mem_in_wire[241]), .SEL(
        pc[2]), .F(n1108) );
  MUX U1126 ( .IN0(inst_mem_in_wire[145]), .IN1(inst_mem_in_wire[177]), .SEL(
        pc[2]), .F(n1109) );
  MUX U1127 ( .IN0(n1109), .IN1(n1108), .SEL(pc[3]), .F(n1110) );
  MUX U1128 ( .IN0(inst_mem_in_wire[81]), .IN1(inst_mem_in_wire[113]), .SEL(
        pc[2]), .F(n1111) );
  MUX U1129 ( .IN0(inst_mem_in_wire[17]), .IN1(inst_mem_in_wire[49]), .SEL(
        pc[2]), .F(n1112) );
  MUX U1130 ( .IN0(n1112), .IN1(n1111), .SEL(pc[3]), .F(n1113) );
  MUX U1131 ( .IN0(n1113), .IN1(n1110), .SEL(pc[4]), .F(n1114) );
  MUX U1132 ( .IN0(n1114), .IN1(n1107), .SEL(pc[5]), .F(n1115) );
  MUX U1133 ( .IN0(n1115), .IN1(n1100), .SEL(pc[6]), .F(n1116) );
  MUX U1134 ( .IN0(n1116), .IN1(n1085), .SEL(pc[7]), .F(opcode[17]) );
  MUX U1135 ( .IN0(inst_mem_in_wire[2002]), .IN1(inst_mem_in_wire[2034]), 
        .SEL(pc[2]), .F(n1117) );
  MUX U1136 ( .IN0(inst_mem_in_wire[1938]), .IN1(inst_mem_in_wire[1970]), 
        .SEL(pc[2]), .F(n1118) );
  MUX U1137 ( .IN0(n1118), .IN1(n1117), .SEL(pc[3]), .F(n1119) );
  MUX U1138 ( .IN0(inst_mem_in_wire[1874]), .IN1(inst_mem_in_wire[1906]), 
        .SEL(pc[2]), .F(n1120) );
  MUX U1139 ( .IN0(inst_mem_in_wire[1810]), .IN1(inst_mem_in_wire[1842]), 
        .SEL(pc[2]), .F(n1121) );
  MUX U1140 ( .IN0(n1121), .IN1(n1120), .SEL(pc[3]), .F(n1122) );
  MUX U1141 ( .IN0(n1122), .IN1(n1119), .SEL(pc[4]), .F(n1123) );
  MUX U1142 ( .IN0(inst_mem_in_wire[1746]), .IN1(inst_mem_in_wire[1778]), 
        .SEL(pc[2]), .F(n1124) );
  MUX U1143 ( .IN0(inst_mem_in_wire[1682]), .IN1(inst_mem_in_wire[1714]), 
        .SEL(pc[2]), .F(n1125) );
  MUX U1144 ( .IN0(n1125), .IN1(n1124), .SEL(pc[3]), .F(n1126) );
  MUX U1145 ( .IN0(inst_mem_in_wire[1618]), .IN1(inst_mem_in_wire[1650]), 
        .SEL(pc[2]), .F(n1127) );
  MUX U1146 ( .IN0(inst_mem_in_wire[1554]), .IN1(inst_mem_in_wire[1586]), 
        .SEL(pc[2]), .F(n1128) );
  MUX U1147 ( .IN0(n1128), .IN1(n1127), .SEL(pc[3]), .F(n1129) );
  MUX U1148 ( .IN0(n1129), .IN1(n1126), .SEL(pc[4]), .F(n1130) );
  MUX U1149 ( .IN0(n1130), .IN1(n1123), .SEL(pc[5]), .F(n1131) );
  MUX U1150 ( .IN0(inst_mem_in_wire[1490]), .IN1(inst_mem_in_wire[1522]), 
        .SEL(pc[2]), .F(n1132) );
  MUX U1151 ( .IN0(inst_mem_in_wire[1426]), .IN1(inst_mem_in_wire[1458]), 
        .SEL(pc[2]), .F(n1133) );
  MUX U1152 ( .IN0(n1133), .IN1(n1132), .SEL(pc[3]), .F(n1134) );
  MUX U1153 ( .IN0(inst_mem_in_wire[1362]), .IN1(inst_mem_in_wire[1394]), 
        .SEL(pc[2]), .F(n1135) );
  MUX U1154 ( .IN0(inst_mem_in_wire[1298]), .IN1(inst_mem_in_wire[1330]), 
        .SEL(pc[2]), .F(n1136) );
  MUX U1155 ( .IN0(n1136), .IN1(n1135), .SEL(pc[3]), .F(n1137) );
  MUX U1156 ( .IN0(n1137), .IN1(n1134), .SEL(pc[4]), .F(n1138) );
  MUX U1157 ( .IN0(inst_mem_in_wire[1234]), .IN1(inst_mem_in_wire[1266]), 
        .SEL(pc[2]), .F(n1139) );
  MUX U1158 ( .IN0(inst_mem_in_wire[1170]), .IN1(inst_mem_in_wire[1202]), 
        .SEL(pc[2]), .F(n1140) );
  MUX U1159 ( .IN0(n1140), .IN1(n1139), .SEL(pc[3]), .F(n1141) );
  MUX U1160 ( .IN0(inst_mem_in_wire[1106]), .IN1(inst_mem_in_wire[1138]), 
        .SEL(pc[2]), .F(n1142) );
  MUX U1161 ( .IN0(inst_mem_in_wire[1042]), .IN1(inst_mem_in_wire[1074]), 
        .SEL(pc[2]), .F(n1143) );
  MUX U1162 ( .IN0(n1143), .IN1(n1142), .SEL(pc[3]), .F(n1144) );
  MUX U1163 ( .IN0(n1144), .IN1(n1141), .SEL(pc[4]), .F(n1145) );
  MUX U1164 ( .IN0(n1145), .IN1(n1138), .SEL(pc[5]), .F(n1146) );
  MUX U1165 ( .IN0(n1146), .IN1(n1131), .SEL(pc[6]), .F(n1147) );
  MUX U1166 ( .IN0(inst_mem_in_wire[978]), .IN1(inst_mem_in_wire[1010]), .SEL(
        pc[2]), .F(n1148) );
  MUX U1167 ( .IN0(inst_mem_in_wire[914]), .IN1(inst_mem_in_wire[946]), .SEL(
        pc[2]), .F(n1149) );
  MUX U1168 ( .IN0(n1149), .IN1(n1148), .SEL(pc[3]), .F(n1150) );
  MUX U1169 ( .IN0(inst_mem_in_wire[850]), .IN1(inst_mem_in_wire[882]), .SEL(
        pc[2]), .F(n1151) );
  MUX U1170 ( .IN0(inst_mem_in_wire[786]), .IN1(inst_mem_in_wire[818]), .SEL(
        pc[2]), .F(n1152) );
  MUX U1171 ( .IN0(n1152), .IN1(n1151), .SEL(pc[3]), .F(n1153) );
  MUX U1172 ( .IN0(n1153), .IN1(n1150), .SEL(pc[4]), .F(n1154) );
  MUX U1173 ( .IN0(inst_mem_in_wire[722]), .IN1(inst_mem_in_wire[754]), .SEL(
        pc[2]), .F(n1155) );
  MUX U1174 ( .IN0(inst_mem_in_wire[658]), .IN1(inst_mem_in_wire[690]), .SEL(
        pc[2]), .F(n1156) );
  MUX U1175 ( .IN0(n1156), .IN1(n1155), .SEL(pc[3]), .F(n1157) );
  MUX U1176 ( .IN0(inst_mem_in_wire[594]), .IN1(inst_mem_in_wire[626]), .SEL(
        pc[2]), .F(n1158) );
  MUX U1177 ( .IN0(inst_mem_in_wire[530]), .IN1(inst_mem_in_wire[562]), .SEL(
        pc[2]), .F(n1159) );
  MUX U1178 ( .IN0(n1159), .IN1(n1158), .SEL(pc[3]), .F(n1160) );
  MUX U1179 ( .IN0(n1160), .IN1(n1157), .SEL(pc[4]), .F(n1161) );
  MUX U1180 ( .IN0(n1161), .IN1(n1154), .SEL(pc[5]), .F(n1162) );
  MUX U1181 ( .IN0(inst_mem_in_wire[466]), .IN1(inst_mem_in_wire[498]), .SEL(
        pc[2]), .F(n1163) );
  MUX U1182 ( .IN0(inst_mem_in_wire[402]), .IN1(inst_mem_in_wire[434]), .SEL(
        pc[2]), .F(n1164) );
  MUX U1183 ( .IN0(n1164), .IN1(n1163), .SEL(pc[3]), .F(n1165) );
  MUX U1184 ( .IN0(inst_mem_in_wire[338]), .IN1(inst_mem_in_wire[370]), .SEL(
        pc[2]), .F(n1166) );
  MUX U1185 ( .IN0(inst_mem_in_wire[274]), .IN1(inst_mem_in_wire[306]), .SEL(
        pc[2]), .F(n1167) );
  MUX U1186 ( .IN0(n1167), .IN1(n1166), .SEL(pc[3]), .F(n1168) );
  MUX U1187 ( .IN0(n1168), .IN1(n1165), .SEL(pc[4]), .F(n1169) );
  MUX U1188 ( .IN0(inst_mem_in_wire[210]), .IN1(inst_mem_in_wire[242]), .SEL(
        pc[2]), .F(n1170) );
  MUX U1189 ( .IN0(inst_mem_in_wire[146]), .IN1(inst_mem_in_wire[178]), .SEL(
        pc[2]), .F(n1171) );
  MUX U1190 ( .IN0(n1171), .IN1(n1170), .SEL(pc[3]), .F(n1172) );
  MUX U1191 ( .IN0(inst_mem_in_wire[82]), .IN1(inst_mem_in_wire[114]), .SEL(
        pc[2]), .F(n1173) );
  MUX U1192 ( .IN0(inst_mem_in_wire[18]), .IN1(inst_mem_in_wire[50]), .SEL(
        pc[2]), .F(n1174) );
  MUX U1193 ( .IN0(n1174), .IN1(n1173), .SEL(pc[3]), .F(n1175) );
  MUX U1194 ( .IN0(n1175), .IN1(n1172), .SEL(pc[4]), .F(n1176) );
  MUX U1195 ( .IN0(n1176), .IN1(n1169), .SEL(pc[5]), .F(n1177) );
  MUX U1196 ( .IN0(n1177), .IN1(n1162), .SEL(pc[6]), .F(n1178) );
  MUX U1197 ( .IN0(n1178), .IN1(n1147), .SEL(pc[7]), .F(opcode[18]) );
  MUX U1198 ( .IN0(inst_mem_in_wire[2003]), .IN1(inst_mem_in_wire[2035]), 
        .SEL(pc[2]), .F(n1179) );
  MUX U1199 ( .IN0(inst_mem_in_wire[1939]), .IN1(inst_mem_in_wire[1971]), 
        .SEL(pc[2]), .F(n1180) );
  MUX U1200 ( .IN0(n1180), .IN1(n1179), .SEL(pc[3]), .F(n1181) );
  MUX U1201 ( .IN0(inst_mem_in_wire[1875]), .IN1(inst_mem_in_wire[1907]), 
        .SEL(pc[2]), .F(n1182) );
  MUX U1202 ( .IN0(inst_mem_in_wire[1811]), .IN1(inst_mem_in_wire[1843]), 
        .SEL(pc[2]), .F(n1183) );
  MUX U1203 ( .IN0(n1183), .IN1(n1182), .SEL(pc[3]), .F(n1184) );
  MUX U1204 ( .IN0(n1184), .IN1(n1181), .SEL(pc[4]), .F(n1185) );
  MUX U1205 ( .IN0(inst_mem_in_wire[1747]), .IN1(inst_mem_in_wire[1779]), 
        .SEL(pc[2]), .F(n1186) );
  MUX U1206 ( .IN0(inst_mem_in_wire[1683]), .IN1(inst_mem_in_wire[1715]), 
        .SEL(pc[2]), .F(n1187) );
  MUX U1207 ( .IN0(n1187), .IN1(n1186), .SEL(pc[3]), .F(n1188) );
  MUX U1208 ( .IN0(inst_mem_in_wire[1619]), .IN1(inst_mem_in_wire[1651]), 
        .SEL(pc[2]), .F(n1189) );
  MUX U1209 ( .IN0(inst_mem_in_wire[1555]), .IN1(inst_mem_in_wire[1587]), 
        .SEL(pc[2]), .F(n1190) );
  MUX U1210 ( .IN0(n1190), .IN1(n1189), .SEL(pc[3]), .F(n1191) );
  MUX U1211 ( .IN0(n1191), .IN1(n1188), .SEL(pc[4]), .F(n1192) );
  MUX U1212 ( .IN0(n1192), .IN1(n1185), .SEL(pc[5]), .F(n1193) );
  MUX U1213 ( .IN0(inst_mem_in_wire[1491]), .IN1(inst_mem_in_wire[1523]), 
        .SEL(pc[2]), .F(n1194) );
  MUX U1214 ( .IN0(inst_mem_in_wire[1427]), .IN1(inst_mem_in_wire[1459]), 
        .SEL(pc[2]), .F(n1195) );
  MUX U1215 ( .IN0(n1195), .IN1(n1194), .SEL(pc[3]), .F(n1196) );
  MUX U1216 ( .IN0(inst_mem_in_wire[1363]), .IN1(inst_mem_in_wire[1395]), 
        .SEL(pc[2]), .F(n1197) );
  MUX U1217 ( .IN0(inst_mem_in_wire[1299]), .IN1(inst_mem_in_wire[1331]), 
        .SEL(pc[2]), .F(n1198) );
  MUX U1218 ( .IN0(n1198), .IN1(n1197), .SEL(pc[3]), .F(n1199) );
  MUX U1219 ( .IN0(n1199), .IN1(n1196), .SEL(pc[4]), .F(n1200) );
  MUX U1220 ( .IN0(inst_mem_in_wire[1235]), .IN1(inst_mem_in_wire[1267]), 
        .SEL(pc[2]), .F(n1201) );
  MUX U1221 ( .IN0(inst_mem_in_wire[1171]), .IN1(inst_mem_in_wire[1203]), 
        .SEL(pc[2]), .F(n1202) );
  MUX U1222 ( .IN0(n1202), .IN1(n1201), .SEL(pc[3]), .F(n1203) );
  MUX U1223 ( .IN0(inst_mem_in_wire[1107]), .IN1(inst_mem_in_wire[1139]), 
        .SEL(pc[2]), .F(n1204) );
  MUX U1224 ( .IN0(inst_mem_in_wire[1043]), .IN1(inst_mem_in_wire[1075]), 
        .SEL(pc[2]), .F(n1205) );
  MUX U1225 ( .IN0(n1205), .IN1(n1204), .SEL(pc[3]), .F(n1206) );
  MUX U1226 ( .IN0(n1206), .IN1(n1203), .SEL(pc[4]), .F(n1207) );
  MUX U1227 ( .IN0(n1207), .IN1(n1200), .SEL(pc[5]), .F(n1208) );
  MUX U1228 ( .IN0(n1208), .IN1(n1193), .SEL(pc[6]), .F(n1209) );
  MUX U1229 ( .IN0(inst_mem_in_wire[979]), .IN1(inst_mem_in_wire[1011]), .SEL(
        pc[2]), .F(n1210) );
  MUX U1230 ( .IN0(inst_mem_in_wire[915]), .IN1(inst_mem_in_wire[947]), .SEL(
        pc[2]), .F(n1211) );
  MUX U1231 ( .IN0(n1211), .IN1(n1210), .SEL(pc[3]), .F(n1212) );
  MUX U1232 ( .IN0(inst_mem_in_wire[851]), .IN1(inst_mem_in_wire[883]), .SEL(
        pc[2]), .F(n1213) );
  MUX U1233 ( .IN0(inst_mem_in_wire[787]), .IN1(inst_mem_in_wire[819]), .SEL(
        pc[2]), .F(n1214) );
  MUX U1234 ( .IN0(n1214), .IN1(n1213), .SEL(pc[3]), .F(n1215) );
  MUX U1235 ( .IN0(n1215), .IN1(n1212), .SEL(pc[4]), .F(n1216) );
  MUX U1236 ( .IN0(inst_mem_in_wire[723]), .IN1(inst_mem_in_wire[755]), .SEL(
        pc[2]), .F(n1217) );
  MUX U1237 ( .IN0(inst_mem_in_wire[659]), .IN1(inst_mem_in_wire[691]), .SEL(
        pc[2]), .F(n1218) );
  MUX U1238 ( .IN0(n1218), .IN1(n1217), .SEL(pc[3]), .F(n1219) );
  MUX U1239 ( .IN0(inst_mem_in_wire[595]), .IN1(inst_mem_in_wire[627]), .SEL(
        pc[2]), .F(n1220) );
  MUX U1240 ( .IN0(inst_mem_in_wire[531]), .IN1(inst_mem_in_wire[563]), .SEL(
        pc[2]), .F(n1221) );
  MUX U1241 ( .IN0(n1221), .IN1(n1220), .SEL(pc[3]), .F(n1222) );
  MUX U1242 ( .IN0(n1222), .IN1(n1219), .SEL(pc[4]), .F(n1223) );
  MUX U1243 ( .IN0(n1223), .IN1(n1216), .SEL(pc[5]), .F(n1224) );
  MUX U1244 ( .IN0(inst_mem_in_wire[467]), .IN1(inst_mem_in_wire[499]), .SEL(
        pc[2]), .F(n1225) );
  MUX U1245 ( .IN0(inst_mem_in_wire[403]), .IN1(inst_mem_in_wire[435]), .SEL(
        pc[2]), .F(n1226) );
  MUX U1246 ( .IN0(n1226), .IN1(n1225), .SEL(pc[3]), .F(n1227) );
  MUX U1247 ( .IN0(inst_mem_in_wire[339]), .IN1(inst_mem_in_wire[371]), .SEL(
        pc[2]), .F(n1228) );
  MUX U1248 ( .IN0(inst_mem_in_wire[275]), .IN1(inst_mem_in_wire[307]), .SEL(
        pc[2]), .F(n1229) );
  MUX U1249 ( .IN0(n1229), .IN1(n1228), .SEL(pc[3]), .F(n1230) );
  MUX U1250 ( .IN0(n1230), .IN1(n1227), .SEL(pc[4]), .F(n1231) );
  MUX U1251 ( .IN0(inst_mem_in_wire[211]), .IN1(inst_mem_in_wire[243]), .SEL(
        pc[2]), .F(n1232) );
  MUX U1252 ( .IN0(inst_mem_in_wire[147]), .IN1(inst_mem_in_wire[179]), .SEL(
        pc[2]), .F(n1233) );
  MUX U1253 ( .IN0(n1233), .IN1(n1232), .SEL(pc[3]), .F(n1234) );
  MUX U1254 ( .IN0(inst_mem_in_wire[83]), .IN1(inst_mem_in_wire[115]), .SEL(
        pc[2]), .F(n1235) );
  MUX U1255 ( .IN0(inst_mem_in_wire[19]), .IN1(inst_mem_in_wire[51]), .SEL(
        pc[2]), .F(n1236) );
  MUX U1256 ( .IN0(n1236), .IN1(n1235), .SEL(pc[3]), .F(n1237) );
  MUX U1257 ( .IN0(n1237), .IN1(n1234), .SEL(pc[4]), .F(n1238) );
  MUX U1258 ( .IN0(n1238), .IN1(n1231), .SEL(pc[5]), .F(n1239) );
  MUX U1259 ( .IN0(n1239), .IN1(n1224), .SEL(pc[6]), .F(n1240) );
  MUX U1260 ( .IN0(n1240), .IN1(n1209), .SEL(pc[7]), .F(opcode[19]) );
  MUX U1261 ( .IN0(inst_mem_in_wire[2004]), .IN1(inst_mem_in_wire[2036]), 
        .SEL(pc[2]), .F(n1241) );
  MUX U1262 ( .IN0(inst_mem_in_wire[1940]), .IN1(inst_mem_in_wire[1972]), 
        .SEL(pc[2]), .F(n1242) );
  MUX U1263 ( .IN0(n1242), .IN1(n1241), .SEL(pc[3]), .F(n1243) );
  MUX U1264 ( .IN0(inst_mem_in_wire[1876]), .IN1(inst_mem_in_wire[1908]), 
        .SEL(pc[2]), .F(n1244) );
  MUX U1265 ( .IN0(inst_mem_in_wire[1812]), .IN1(inst_mem_in_wire[1844]), 
        .SEL(pc[2]), .F(n1245) );
  MUX U1266 ( .IN0(n1245), .IN1(n1244), .SEL(pc[3]), .F(n1246) );
  MUX U1267 ( .IN0(n1246), .IN1(n1243), .SEL(pc[4]), .F(n1247) );
  MUX U1268 ( .IN0(inst_mem_in_wire[1748]), .IN1(inst_mem_in_wire[1780]), 
        .SEL(pc[2]), .F(n1248) );
  MUX U1269 ( .IN0(inst_mem_in_wire[1684]), .IN1(inst_mem_in_wire[1716]), 
        .SEL(pc[2]), .F(n1249) );
  MUX U1270 ( .IN0(n1249), .IN1(n1248), .SEL(pc[3]), .F(n1250) );
  MUX U1271 ( .IN0(inst_mem_in_wire[1620]), .IN1(inst_mem_in_wire[1652]), 
        .SEL(pc[2]), .F(n1251) );
  MUX U1272 ( .IN0(inst_mem_in_wire[1556]), .IN1(inst_mem_in_wire[1588]), 
        .SEL(pc[2]), .F(n1252) );
  MUX U1273 ( .IN0(n1252), .IN1(n1251), .SEL(pc[3]), .F(n1253) );
  MUX U1274 ( .IN0(n1253), .IN1(n1250), .SEL(pc[4]), .F(n1254) );
  MUX U1275 ( .IN0(n1254), .IN1(n1247), .SEL(pc[5]), .F(n1255) );
  MUX U1276 ( .IN0(inst_mem_in_wire[1492]), .IN1(inst_mem_in_wire[1524]), 
        .SEL(pc[2]), .F(n1256) );
  MUX U1277 ( .IN0(inst_mem_in_wire[1428]), .IN1(inst_mem_in_wire[1460]), 
        .SEL(pc[2]), .F(n1257) );
  MUX U1278 ( .IN0(n1257), .IN1(n1256), .SEL(pc[3]), .F(n1258) );
  MUX U1279 ( .IN0(inst_mem_in_wire[1364]), .IN1(inst_mem_in_wire[1396]), 
        .SEL(pc[2]), .F(n1259) );
  MUX U1280 ( .IN0(inst_mem_in_wire[1300]), .IN1(inst_mem_in_wire[1332]), 
        .SEL(pc[2]), .F(n1260) );
  MUX U1281 ( .IN0(n1260), .IN1(n1259), .SEL(pc[3]), .F(n1261) );
  MUX U1282 ( .IN0(n1261), .IN1(n1258), .SEL(pc[4]), .F(n1262) );
  MUX U1283 ( .IN0(inst_mem_in_wire[1236]), .IN1(inst_mem_in_wire[1268]), 
        .SEL(pc[2]), .F(n1263) );
  MUX U1284 ( .IN0(inst_mem_in_wire[1172]), .IN1(inst_mem_in_wire[1204]), 
        .SEL(pc[2]), .F(n1264) );
  MUX U1285 ( .IN0(n1264), .IN1(n1263), .SEL(pc[3]), .F(n1265) );
  MUX U1286 ( .IN0(inst_mem_in_wire[1108]), .IN1(inst_mem_in_wire[1140]), 
        .SEL(pc[2]), .F(n1266) );
  MUX U1287 ( .IN0(inst_mem_in_wire[1044]), .IN1(inst_mem_in_wire[1076]), 
        .SEL(pc[2]), .F(n1267) );
  MUX U1288 ( .IN0(n1267), .IN1(n1266), .SEL(pc[3]), .F(n1268) );
  MUX U1289 ( .IN0(n1268), .IN1(n1265), .SEL(pc[4]), .F(n1269) );
  MUX U1290 ( .IN0(n1269), .IN1(n1262), .SEL(pc[5]), .F(n1270) );
  MUX U1291 ( .IN0(n1270), .IN1(n1255), .SEL(pc[6]), .F(n1271) );
  MUX U1292 ( .IN0(inst_mem_in_wire[980]), .IN1(inst_mem_in_wire[1012]), .SEL(
        pc[2]), .F(n1272) );
  MUX U1293 ( .IN0(inst_mem_in_wire[916]), .IN1(inst_mem_in_wire[948]), .SEL(
        pc[2]), .F(n1273) );
  MUX U1294 ( .IN0(n1273), .IN1(n1272), .SEL(pc[3]), .F(n1274) );
  MUX U1295 ( .IN0(inst_mem_in_wire[852]), .IN1(inst_mem_in_wire[884]), .SEL(
        pc[2]), .F(n1275) );
  MUX U1296 ( .IN0(inst_mem_in_wire[788]), .IN1(inst_mem_in_wire[820]), .SEL(
        pc[2]), .F(n1276) );
  MUX U1297 ( .IN0(n1276), .IN1(n1275), .SEL(pc[3]), .F(n1277) );
  MUX U1298 ( .IN0(n1277), .IN1(n1274), .SEL(pc[4]), .F(n1278) );
  MUX U1299 ( .IN0(inst_mem_in_wire[724]), .IN1(inst_mem_in_wire[756]), .SEL(
        pc[2]), .F(n1279) );
  MUX U1300 ( .IN0(inst_mem_in_wire[660]), .IN1(inst_mem_in_wire[692]), .SEL(
        pc[2]), .F(n1280) );
  MUX U1301 ( .IN0(n1280), .IN1(n1279), .SEL(pc[3]), .F(n1281) );
  MUX U1302 ( .IN0(inst_mem_in_wire[596]), .IN1(inst_mem_in_wire[628]), .SEL(
        pc[2]), .F(n1282) );
  MUX U1303 ( .IN0(inst_mem_in_wire[532]), .IN1(inst_mem_in_wire[564]), .SEL(
        pc[2]), .F(n1283) );
  MUX U1304 ( .IN0(n1283), .IN1(n1282), .SEL(pc[3]), .F(n1284) );
  MUX U1305 ( .IN0(n1284), .IN1(n1281), .SEL(pc[4]), .F(n1285) );
  MUX U1306 ( .IN0(n1285), .IN1(n1278), .SEL(pc[5]), .F(n1286) );
  MUX U1307 ( .IN0(inst_mem_in_wire[468]), .IN1(inst_mem_in_wire[500]), .SEL(
        pc[2]), .F(n1287) );
  MUX U1308 ( .IN0(inst_mem_in_wire[404]), .IN1(inst_mem_in_wire[436]), .SEL(
        pc[2]), .F(n1288) );
  MUX U1309 ( .IN0(n1288), .IN1(n1287), .SEL(pc[3]), .F(n1289) );
  MUX U1310 ( .IN0(inst_mem_in_wire[340]), .IN1(inst_mem_in_wire[372]), .SEL(
        pc[2]), .F(n1290) );
  MUX U1311 ( .IN0(inst_mem_in_wire[276]), .IN1(inst_mem_in_wire[308]), .SEL(
        pc[2]), .F(n1291) );
  MUX U1312 ( .IN0(n1291), .IN1(n1290), .SEL(pc[3]), .F(n1292) );
  MUX U1313 ( .IN0(n1292), .IN1(n1289), .SEL(pc[4]), .F(n1293) );
  MUX U1314 ( .IN0(inst_mem_in_wire[212]), .IN1(inst_mem_in_wire[244]), .SEL(
        pc[2]), .F(n1294) );
  MUX U1315 ( .IN0(inst_mem_in_wire[148]), .IN1(inst_mem_in_wire[180]), .SEL(
        pc[2]), .F(n1295) );
  MUX U1316 ( .IN0(n1295), .IN1(n1294), .SEL(pc[3]), .F(n1296) );
  MUX U1317 ( .IN0(inst_mem_in_wire[84]), .IN1(inst_mem_in_wire[116]), .SEL(
        pc[2]), .F(n1297) );
  MUX U1318 ( .IN0(inst_mem_in_wire[20]), .IN1(inst_mem_in_wire[52]), .SEL(
        pc[2]), .F(n1298) );
  MUX U1319 ( .IN0(n1298), .IN1(n1297), .SEL(pc[3]), .F(n1299) );
  MUX U1320 ( .IN0(n1299), .IN1(n1296), .SEL(pc[4]), .F(n1300) );
  MUX U1321 ( .IN0(n1300), .IN1(n1293), .SEL(pc[5]), .F(n1301) );
  MUX U1322 ( .IN0(n1301), .IN1(n1286), .SEL(pc[6]), .F(n1302) );
  MUX U1323 ( .IN0(n1302), .IN1(n1271), .SEL(pc[7]), .F(opcode[20]) );
  MUX U1324 ( .IN0(inst_mem_in_wire[2005]), .IN1(inst_mem_in_wire[2037]), 
        .SEL(pc[2]), .F(n1303) );
  MUX U1325 ( .IN0(inst_mem_in_wire[1941]), .IN1(inst_mem_in_wire[1973]), 
        .SEL(pc[2]), .F(n1304) );
  MUX U1326 ( .IN0(n1304), .IN1(n1303), .SEL(pc[3]), .F(n1305) );
  MUX U1327 ( .IN0(inst_mem_in_wire[1877]), .IN1(inst_mem_in_wire[1909]), 
        .SEL(pc[2]), .F(n1306) );
  MUX U1328 ( .IN0(inst_mem_in_wire[1813]), .IN1(inst_mem_in_wire[1845]), 
        .SEL(pc[2]), .F(n1307) );
  MUX U1329 ( .IN0(n1307), .IN1(n1306), .SEL(pc[3]), .F(n1308) );
  MUX U1330 ( .IN0(n1308), .IN1(n1305), .SEL(pc[4]), .F(n1309) );
  MUX U1331 ( .IN0(inst_mem_in_wire[1749]), .IN1(inst_mem_in_wire[1781]), 
        .SEL(pc[2]), .F(n1310) );
  MUX U1332 ( .IN0(inst_mem_in_wire[1685]), .IN1(inst_mem_in_wire[1717]), 
        .SEL(pc[2]), .F(n1311) );
  MUX U1333 ( .IN0(n1311), .IN1(n1310), .SEL(pc[3]), .F(n1312) );
  MUX U1334 ( .IN0(inst_mem_in_wire[1621]), .IN1(inst_mem_in_wire[1653]), 
        .SEL(pc[2]), .F(n1313) );
  MUX U1335 ( .IN0(inst_mem_in_wire[1557]), .IN1(inst_mem_in_wire[1589]), 
        .SEL(pc[2]), .F(n1314) );
  MUX U1336 ( .IN0(n1314), .IN1(n1313), .SEL(pc[3]), .F(n1315) );
  MUX U1337 ( .IN0(n1315), .IN1(n1312), .SEL(pc[4]), .F(n1316) );
  MUX U1338 ( .IN0(n1316), .IN1(n1309), .SEL(pc[5]), .F(n1317) );
  MUX U1339 ( .IN0(inst_mem_in_wire[1493]), .IN1(inst_mem_in_wire[1525]), 
        .SEL(pc[2]), .F(n1318) );
  MUX U1340 ( .IN0(inst_mem_in_wire[1429]), .IN1(inst_mem_in_wire[1461]), 
        .SEL(pc[2]), .F(n1319) );
  MUX U1341 ( .IN0(n1319), .IN1(n1318), .SEL(pc[3]), .F(n1320) );
  MUX U1342 ( .IN0(inst_mem_in_wire[1365]), .IN1(inst_mem_in_wire[1397]), 
        .SEL(pc[2]), .F(n1321) );
  MUX U1343 ( .IN0(inst_mem_in_wire[1301]), .IN1(inst_mem_in_wire[1333]), 
        .SEL(pc[2]), .F(n1322) );
  MUX U1344 ( .IN0(n1322), .IN1(n1321), .SEL(pc[3]), .F(n1323) );
  MUX U1345 ( .IN0(n1323), .IN1(n1320), .SEL(pc[4]), .F(n1324) );
  MUX U1346 ( .IN0(inst_mem_in_wire[1237]), .IN1(inst_mem_in_wire[1269]), 
        .SEL(pc[2]), .F(n1325) );
  MUX U1347 ( .IN0(inst_mem_in_wire[1173]), .IN1(inst_mem_in_wire[1205]), 
        .SEL(pc[2]), .F(n1326) );
  MUX U1348 ( .IN0(n1326), .IN1(n1325), .SEL(pc[3]), .F(n1327) );
  MUX U1349 ( .IN0(inst_mem_in_wire[1109]), .IN1(inst_mem_in_wire[1141]), 
        .SEL(pc[2]), .F(n1328) );
  MUX U1350 ( .IN0(inst_mem_in_wire[1045]), .IN1(inst_mem_in_wire[1077]), 
        .SEL(pc[2]), .F(n1329) );
  MUX U1351 ( .IN0(n1329), .IN1(n1328), .SEL(pc[3]), .F(n1330) );
  MUX U1352 ( .IN0(n1330), .IN1(n1327), .SEL(pc[4]), .F(n1331) );
  MUX U1353 ( .IN0(n1331), .IN1(n1324), .SEL(pc[5]), .F(n1332) );
  MUX U1354 ( .IN0(n1332), .IN1(n1317), .SEL(pc[6]), .F(n1333) );
  MUX U1355 ( .IN0(inst_mem_in_wire[981]), .IN1(inst_mem_in_wire[1013]), .SEL(
        pc[2]), .F(n1334) );
  MUX U1356 ( .IN0(inst_mem_in_wire[917]), .IN1(inst_mem_in_wire[949]), .SEL(
        pc[2]), .F(n1335) );
  MUX U1357 ( .IN0(n1335), .IN1(n1334), .SEL(pc[3]), .F(n1336) );
  MUX U1358 ( .IN0(inst_mem_in_wire[853]), .IN1(inst_mem_in_wire[885]), .SEL(
        pc[2]), .F(n1337) );
  MUX U1359 ( .IN0(inst_mem_in_wire[789]), .IN1(inst_mem_in_wire[821]), .SEL(
        pc[2]), .F(n1338) );
  MUX U1360 ( .IN0(n1338), .IN1(n1337), .SEL(pc[3]), .F(n1339) );
  MUX U1361 ( .IN0(n1339), .IN1(n1336), .SEL(pc[4]), .F(n1340) );
  MUX U1362 ( .IN0(inst_mem_in_wire[725]), .IN1(inst_mem_in_wire[757]), .SEL(
        pc[2]), .F(n1341) );
  MUX U1363 ( .IN0(inst_mem_in_wire[661]), .IN1(inst_mem_in_wire[693]), .SEL(
        pc[2]), .F(n1342) );
  MUX U1364 ( .IN0(n1342), .IN1(n1341), .SEL(pc[3]), .F(n1343) );
  MUX U1365 ( .IN0(inst_mem_in_wire[597]), .IN1(inst_mem_in_wire[629]), .SEL(
        pc[2]), .F(n1344) );
  MUX U1366 ( .IN0(inst_mem_in_wire[533]), .IN1(inst_mem_in_wire[565]), .SEL(
        pc[2]), .F(n1345) );
  MUX U1367 ( .IN0(n1345), .IN1(n1344), .SEL(pc[3]), .F(n1346) );
  MUX U1368 ( .IN0(n1346), .IN1(n1343), .SEL(pc[4]), .F(n1347) );
  MUX U1369 ( .IN0(n1347), .IN1(n1340), .SEL(pc[5]), .F(n1348) );
  MUX U1370 ( .IN0(inst_mem_in_wire[469]), .IN1(inst_mem_in_wire[501]), .SEL(
        pc[2]), .F(n1349) );
  MUX U1371 ( .IN0(inst_mem_in_wire[405]), .IN1(inst_mem_in_wire[437]), .SEL(
        pc[2]), .F(n1350) );
  MUX U1372 ( .IN0(n1350), .IN1(n1349), .SEL(pc[3]), .F(n1351) );
  MUX U1373 ( .IN0(inst_mem_in_wire[341]), .IN1(inst_mem_in_wire[373]), .SEL(
        pc[2]), .F(n1352) );
  MUX U1374 ( .IN0(inst_mem_in_wire[277]), .IN1(inst_mem_in_wire[309]), .SEL(
        pc[2]), .F(n1353) );
  MUX U1375 ( .IN0(n1353), .IN1(n1352), .SEL(pc[3]), .F(n1354) );
  MUX U1376 ( .IN0(n1354), .IN1(n1351), .SEL(pc[4]), .F(n1355) );
  MUX U1377 ( .IN0(inst_mem_in_wire[213]), .IN1(inst_mem_in_wire[245]), .SEL(
        pc[2]), .F(n1356) );
  MUX U1378 ( .IN0(inst_mem_in_wire[149]), .IN1(inst_mem_in_wire[181]), .SEL(
        pc[2]), .F(n1357) );
  MUX U1379 ( .IN0(n1357), .IN1(n1356), .SEL(pc[3]), .F(n1358) );
  MUX U1380 ( .IN0(inst_mem_in_wire[85]), .IN1(inst_mem_in_wire[117]), .SEL(
        pc[2]), .F(n1359) );
  MUX U1381 ( .IN0(inst_mem_in_wire[21]), .IN1(inst_mem_in_wire[53]), .SEL(
        pc[2]), .F(n1360) );
  MUX U1382 ( .IN0(n1360), .IN1(n1359), .SEL(pc[3]), .F(n1361) );
  MUX U1383 ( .IN0(n1361), .IN1(n1358), .SEL(pc[4]), .F(n1362) );
  MUX U1384 ( .IN0(n1362), .IN1(n1355), .SEL(pc[5]), .F(n1363) );
  MUX U1385 ( .IN0(n1363), .IN1(n1348), .SEL(pc[6]), .F(n1364) );
  MUX U1386 ( .IN0(n1364), .IN1(n1333), .SEL(pc[7]), .F(opcode[21]) );
  MUX U1387 ( .IN0(inst_mem_in_wire[2006]), .IN1(inst_mem_in_wire[2038]), 
        .SEL(pc[2]), .F(n1365) );
  MUX U1388 ( .IN0(inst_mem_in_wire[1942]), .IN1(inst_mem_in_wire[1974]), 
        .SEL(pc[2]), .F(n1366) );
  MUX U1389 ( .IN0(n1366), .IN1(n1365), .SEL(pc[3]), .F(n1367) );
  MUX U1390 ( .IN0(inst_mem_in_wire[1878]), .IN1(inst_mem_in_wire[1910]), 
        .SEL(pc[2]), .F(n1368) );
  MUX U1391 ( .IN0(inst_mem_in_wire[1814]), .IN1(inst_mem_in_wire[1846]), 
        .SEL(pc[2]), .F(n1369) );
  MUX U1392 ( .IN0(n1369), .IN1(n1368), .SEL(pc[3]), .F(n1370) );
  MUX U1393 ( .IN0(n1370), .IN1(n1367), .SEL(pc[4]), .F(n1371) );
  MUX U1394 ( .IN0(inst_mem_in_wire[1750]), .IN1(inst_mem_in_wire[1782]), 
        .SEL(pc[2]), .F(n1372) );
  MUX U1395 ( .IN0(inst_mem_in_wire[1686]), .IN1(inst_mem_in_wire[1718]), 
        .SEL(pc[2]), .F(n1373) );
  MUX U1396 ( .IN0(n1373), .IN1(n1372), .SEL(pc[3]), .F(n1374) );
  MUX U1397 ( .IN0(inst_mem_in_wire[1622]), .IN1(inst_mem_in_wire[1654]), 
        .SEL(pc[2]), .F(n1375) );
  MUX U1398 ( .IN0(inst_mem_in_wire[1558]), .IN1(inst_mem_in_wire[1590]), 
        .SEL(pc[2]), .F(n1376) );
  MUX U1399 ( .IN0(n1376), .IN1(n1375), .SEL(pc[3]), .F(n1377) );
  MUX U1400 ( .IN0(n1377), .IN1(n1374), .SEL(pc[4]), .F(n1378) );
  MUX U1401 ( .IN0(n1378), .IN1(n1371), .SEL(pc[5]), .F(n1379) );
  MUX U1402 ( .IN0(inst_mem_in_wire[1494]), .IN1(inst_mem_in_wire[1526]), 
        .SEL(pc[2]), .F(n1380) );
  MUX U1403 ( .IN0(inst_mem_in_wire[1430]), .IN1(inst_mem_in_wire[1462]), 
        .SEL(pc[2]), .F(n1381) );
  MUX U1404 ( .IN0(n1381), .IN1(n1380), .SEL(pc[3]), .F(n1382) );
  MUX U1405 ( .IN0(inst_mem_in_wire[1366]), .IN1(inst_mem_in_wire[1398]), 
        .SEL(pc[2]), .F(n1383) );
  MUX U1406 ( .IN0(inst_mem_in_wire[1302]), .IN1(inst_mem_in_wire[1334]), 
        .SEL(pc[2]), .F(n1384) );
  MUX U1407 ( .IN0(n1384), .IN1(n1383), .SEL(pc[3]), .F(n1385) );
  MUX U1408 ( .IN0(n1385), .IN1(n1382), .SEL(pc[4]), .F(n1386) );
  MUX U1409 ( .IN0(inst_mem_in_wire[1238]), .IN1(inst_mem_in_wire[1270]), 
        .SEL(pc[2]), .F(n1387) );
  MUX U1410 ( .IN0(inst_mem_in_wire[1174]), .IN1(inst_mem_in_wire[1206]), 
        .SEL(pc[2]), .F(n1388) );
  MUX U1411 ( .IN0(n1388), .IN1(n1387), .SEL(pc[3]), .F(n1389) );
  MUX U1412 ( .IN0(inst_mem_in_wire[1110]), .IN1(inst_mem_in_wire[1142]), 
        .SEL(pc[2]), .F(n1390) );
  MUX U1413 ( .IN0(inst_mem_in_wire[1046]), .IN1(inst_mem_in_wire[1078]), 
        .SEL(pc[2]), .F(n1391) );
  MUX U1414 ( .IN0(n1391), .IN1(n1390), .SEL(pc[3]), .F(n1392) );
  MUX U1415 ( .IN0(n1392), .IN1(n1389), .SEL(pc[4]), .F(n1393) );
  MUX U1416 ( .IN0(n1393), .IN1(n1386), .SEL(pc[5]), .F(n1394) );
  MUX U1417 ( .IN0(n1394), .IN1(n1379), .SEL(pc[6]), .F(n1395) );
  MUX U1418 ( .IN0(inst_mem_in_wire[982]), .IN1(inst_mem_in_wire[1014]), .SEL(
        pc[2]), .F(n1396) );
  MUX U1419 ( .IN0(inst_mem_in_wire[918]), .IN1(inst_mem_in_wire[950]), .SEL(
        pc[2]), .F(n1397) );
  MUX U1420 ( .IN0(n1397), .IN1(n1396), .SEL(pc[3]), .F(n1398) );
  MUX U1421 ( .IN0(inst_mem_in_wire[854]), .IN1(inst_mem_in_wire[886]), .SEL(
        pc[2]), .F(n1399) );
  MUX U1422 ( .IN0(inst_mem_in_wire[790]), .IN1(inst_mem_in_wire[822]), .SEL(
        pc[2]), .F(n1400) );
  MUX U1423 ( .IN0(n1400), .IN1(n1399), .SEL(pc[3]), .F(n1401) );
  MUX U1424 ( .IN0(n1401), .IN1(n1398), .SEL(pc[4]), .F(n1402) );
  MUX U1425 ( .IN0(inst_mem_in_wire[726]), .IN1(inst_mem_in_wire[758]), .SEL(
        pc[2]), .F(n1403) );
  MUX U1426 ( .IN0(inst_mem_in_wire[662]), .IN1(inst_mem_in_wire[694]), .SEL(
        pc[2]), .F(n1404) );
  MUX U1427 ( .IN0(n1404), .IN1(n1403), .SEL(pc[3]), .F(n1405) );
  MUX U1428 ( .IN0(inst_mem_in_wire[598]), .IN1(inst_mem_in_wire[630]), .SEL(
        pc[2]), .F(n1406) );
  MUX U1429 ( .IN0(inst_mem_in_wire[534]), .IN1(inst_mem_in_wire[566]), .SEL(
        pc[2]), .F(n1407) );
  MUX U1430 ( .IN0(n1407), .IN1(n1406), .SEL(pc[3]), .F(n1408) );
  MUX U1431 ( .IN0(n1408), .IN1(n1405), .SEL(pc[4]), .F(n1409) );
  MUX U1432 ( .IN0(n1409), .IN1(n1402), .SEL(pc[5]), .F(n1410) );
  MUX U1433 ( .IN0(inst_mem_in_wire[470]), .IN1(inst_mem_in_wire[502]), .SEL(
        pc[2]), .F(n1411) );
  MUX U1434 ( .IN0(inst_mem_in_wire[406]), .IN1(inst_mem_in_wire[438]), .SEL(
        pc[2]), .F(n1412) );
  MUX U1435 ( .IN0(n1412), .IN1(n1411), .SEL(pc[3]), .F(n1413) );
  MUX U1436 ( .IN0(inst_mem_in_wire[342]), .IN1(inst_mem_in_wire[374]), .SEL(
        pc[2]), .F(n1414) );
  MUX U1437 ( .IN0(inst_mem_in_wire[278]), .IN1(inst_mem_in_wire[310]), .SEL(
        pc[2]), .F(n1415) );
  MUX U1438 ( .IN0(n1415), .IN1(n1414), .SEL(pc[3]), .F(n1416) );
  MUX U1439 ( .IN0(n1416), .IN1(n1413), .SEL(pc[4]), .F(n1417) );
  MUX U1440 ( .IN0(inst_mem_in_wire[214]), .IN1(inst_mem_in_wire[246]), .SEL(
        pc[2]), .F(n1418) );
  MUX U1441 ( .IN0(inst_mem_in_wire[150]), .IN1(inst_mem_in_wire[182]), .SEL(
        pc[2]), .F(n1419) );
  MUX U1442 ( .IN0(n1419), .IN1(n1418), .SEL(pc[3]), .F(n1420) );
  MUX U1443 ( .IN0(inst_mem_in_wire[86]), .IN1(inst_mem_in_wire[118]), .SEL(
        pc[2]), .F(n1421) );
  MUX U1444 ( .IN0(inst_mem_in_wire[22]), .IN1(inst_mem_in_wire[54]), .SEL(
        pc[2]), .F(n1422) );
  MUX U1445 ( .IN0(n1422), .IN1(n1421), .SEL(pc[3]), .F(n1423) );
  MUX U1446 ( .IN0(n1423), .IN1(n1420), .SEL(pc[4]), .F(n1424) );
  MUX U1447 ( .IN0(n1424), .IN1(n1417), .SEL(pc[5]), .F(n1425) );
  MUX U1448 ( .IN0(n1425), .IN1(n1410), .SEL(pc[6]), .F(n1426) );
  MUX U1449 ( .IN0(n1426), .IN1(n1395), .SEL(pc[7]), .F(opcode[22]) );
  MUX U1450 ( .IN0(inst_mem_in_wire[2007]), .IN1(inst_mem_in_wire[2039]), 
        .SEL(pc[2]), .F(n1427) );
  MUX U1451 ( .IN0(inst_mem_in_wire[1943]), .IN1(inst_mem_in_wire[1975]), 
        .SEL(pc[2]), .F(n1428) );
  MUX U1452 ( .IN0(n1428), .IN1(n1427), .SEL(pc[3]), .F(n1429) );
  MUX U1453 ( .IN0(inst_mem_in_wire[1879]), .IN1(inst_mem_in_wire[1911]), 
        .SEL(pc[2]), .F(n1430) );
  MUX U1454 ( .IN0(inst_mem_in_wire[1815]), .IN1(inst_mem_in_wire[1847]), 
        .SEL(pc[2]), .F(n1431) );
  MUX U1455 ( .IN0(n1431), .IN1(n1430), .SEL(pc[3]), .F(n1432) );
  MUX U1456 ( .IN0(n1432), .IN1(n1429), .SEL(pc[4]), .F(n1433) );
  MUX U1457 ( .IN0(inst_mem_in_wire[1751]), .IN1(inst_mem_in_wire[1783]), 
        .SEL(pc[2]), .F(n1434) );
  MUX U1458 ( .IN0(inst_mem_in_wire[1687]), .IN1(inst_mem_in_wire[1719]), 
        .SEL(pc[2]), .F(n1435) );
  MUX U1459 ( .IN0(n1435), .IN1(n1434), .SEL(pc[3]), .F(n1436) );
  MUX U1460 ( .IN0(inst_mem_in_wire[1623]), .IN1(inst_mem_in_wire[1655]), 
        .SEL(pc[2]), .F(n1437) );
  MUX U1461 ( .IN0(inst_mem_in_wire[1559]), .IN1(inst_mem_in_wire[1591]), 
        .SEL(pc[2]), .F(n1438) );
  MUX U1462 ( .IN0(n1438), .IN1(n1437), .SEL(pc[3]), .F(n1439) );
  MUX U1463 ( .IN0(n1439), .IN1(n1436), .SEL(pc[4]), .F(n1440) );
  MUX U1464 ( .IN0(n1440), .IN1(n1433), .SEL(pc[5]), .F(n1441) );
  MUX U1465 ( .IN0(inst_mem_in_wire[1495]), .IN1(inst_mem_in_wire[1527]), 
        .SEL(pc[2]), .F(n1442) );
  MUX U1466 ( .IN0(inst_mem_in_wire[1431]), .IN1(inst_mem_in_wire[1463]), 
        .SEL(pc[2]), .F(n1443) );
  MUX U1467 ( .IN0(n1443), .IN1(n1442), .SEL(pc[3]), .F(n1444) );
  MUX U1468 ( .IN0(inst_mem_in_wire[1367]), .IN1(inst_mem_in_wire[1399]), 
        .SEL(pc[2]), .F(n1445) );
  MUX U1469 ( .IN0(inst_mem_in_wire[1303]), .IN1(inst_mem_in_wire[1335]), 
        .SEL(pc[2]), .F(n1446) );
  MUX U1470 ( .IN0(n1446), .IN1(n1445), .SEL(pc[3]), .F(n1447) );
  MUX U1471 ( .IN0(n1447), .IN1(n1444), .SEL(pc[4]), .F(n1448) );
  MUX U1472 ( .IN0(inst_mem_in_wire[1239]), .IN1(inst_mem_in_wire[1271]), 
        .SEL(pc[2]), .F(n1449) );
  MUX U1473 ( .IN0(inst_mem_in_wire[1175]), .IN1(inst_mem_in_wire[1207]), 
        .SEL(pc[2]), .F(n1450) );
  MUX U1474 ( .IN0(n1450), .IN1(n1449), .SEL(pc[3]), .F(n1451) );
  MUX U1475 ( .IN0(inst_mem_in_wire[1111]), .IN1(inst_mem_in_wire[1143]), 
        .SEL(pc[2]), .F(n1452) );
  MUX U1476 ( .IN0(inst_mem_in_wire[1047]), .IN1(inst_mem_in_wire[1079]), 
        .SEL(pc[2]), .F(n1453) );
  MUX U1477 ( .IN0(n1453), .IN1(n1452), .SEL(pc[3]), .F(n1454) );
  MUX U1478 ( .IN0(n1454), .IN1(n1451), .SEL(pc[4]), .F(n1455) );
  MUX U1479 ( .IN0(n1455), .IN1(n1448), .SEL(pc[5]), .F(n1456) );
  MUX U1480 ( .IN0(n1456), .IN1(n1441), .SEL(pc[6]), .F(n1457) );
  MUX U1481 ( .IN0(inst_mem_in_wire[983]), .IN1(inst_mem_in_wire[1015]), .SEL(
        pc[2]), .F(n1458) );
  MUX U1482 ( .IN0(inst_mem_in_wire[919]), .IN1(inst_mem_in_wire[951]), .SEL(
        pc[2]), .F(n1459) );
  MUX U1483 ( .IN0(n1459), .IN1(n1458), .SEL(pc[3]), .F(n1460) );
  MUX U1484 ( .IN0(inst_mem_in_wire[855]), .IN1(inst_mem_in_wire[887]), .SEL(
        pc[2]), .F(n1461) );
  MUX U1485 ( .IN0(inst_mem_in_wire[791]), .IN1(inst_mem_in_wire[823]), .SEL(
        pc[2]), .F(n1462) );
  MUX U1486 ( .IN0(n1462), .IN1(n1461), .SEL(pc[3]), .F(n1463) );
  MUX U1487 ( .IN0(n1463), .IN1(n1460), .SEL(pc[4]), .F(n1464) );
  MUX U1488 ( .IN0(inst_mem_in_wire[727]), .IN1(inst_mem_in_wire[759]), .SEL(
        pc[2]), .F(n1465) );
  MUX U1489 ( .IN0(inst_mem_in_wire[663]), .IN1(inst_mem_in_wire[695]), .SEL(
        pc[2]), .F(n1466) );
  MUX U1490 ( .IN0(n1466), .IN1(n1465), .SEL(pc[3]), .F(n1467) );
  MUX U1491 ( .IN0(inst_mem_in_wire[599]), .IN1(inst_mem_in_wire[631]), .SEL(
        pc[2]), .F(n1468) );
  MUX U1492 ( .IN0(inst_mem_in_wire[535]), .IN1(inst_mem_in_wire[567]), .SEL(
        pc[2]), .F(n1469) );
  MUX U1493 ( .IN0(n1469), .IN1(n1468), .SEL(pc[3]), .F(n1470) );
  MUX U1494 ( .IN0(n1470), .IN1(n1467), .SEL(pc[4]), .F(n1471) );
  MUX U1495 ( .IN0(n1471), .IN1(n1464), .SEL(pc[5]), .F(n1472) );
  MUX U1496 ( .IN0(inst_mem_in_wire[471]), .IN1(inst_mem_in_wire[503]), .SEL(
        pc[2]), .F(n1473) );
  MUX U1497 ( .IN0(inst_mem_in_wire[407]), .IN1(inst_mem_in_wire[439]), .SEL(
        pc[2]), .F(n1474) );
  MUX U1498 ( .IN0(n1474), .IN1(n1473), .SEL(pc[3]), .F(n1475) );
  MUX U1499 ( .IN0(inst_mem_in_wire[343]), .IN1(inst_mem_in_wire[375]), .SEL(
        pc[2]), .F(n1476) );
  MUX U1500 ( .IN0(inst_mem_in_wire[279]), .IN1(inst_mem_in_wire[311]), .SEL(
        pc[2]), .F(n1477) );
  MUX U1501 ( .IN0(n1477), .IN1(n1476), .SEL(pc[3]), .F(n1478) );
  MUX U1502 ( .IN0(n1478), .IN1(n1475), .SEL(pc[4]), .F(n1479) );
  MUX U1503 ( .IN0(inst_mem_in_wire[215]), .IN1(inst_mem_in_wire[247]), .SEL(
        pc[2]), .F(n1480) );
  MUX U1504 ( .IN0(inst_mem_in_wire[151]), .IN1(inst_mem_in_wire[183]), .SEL(
        pc[2]), .F(n1481) );
  MUX U1505 ( .IN0(n1481), .IN1(n1480), .SEL(pc[3]), .F(n1482) );
  MUX U1506 ( .IN0(inst_mem_in_wire[87]), .IN1(inst_mem_in_wire[119]), .SEL(
        pc[2]), .F(n1483) );
  MUX U1507 ( .IN0(inst_mem_in_wire[23]), .IN1(inst_mem_in_wire[55]), .SEL(
        pc[2]), .F(n1484) );
  MUX U1508 ( .IN0(n1484), .IN1(n1483), .SEL(pc[3]), .F(n1485) );
  MUX U1509 ( .IN0(n1485), .IN1(n1482), .SEL(pc[4]), .F(n1486) );
  MUX U1510 ( .IN0(n1486), .IN1(n1479), .SEL(pc[5]), .F(n1487) );
  MUX U1511 ( .IN0(n1487), .IN1(n1472), .SEL(pc[6]), .F(n1488) );
  MUX U1512 ( .IN0(n1488), .IN1(n1457), .SEL(pc[7]), .F(opcode[23]) );
  MUX U1513 ( .IN0(inst_mem_in_wire[2008]), .IN1(inst_mem_in_wire[2040]), 
        .SEL(pc[2]), .F(n1489) );
  MUX U1514 ( .IN0(inst_mem_in_wire[1944]), .IN1(inst_mem_in_wire[1976]), 
        .SEL(pc[2]), .F(n1490) );
  MUX U1515 ( .IN0(n1490), .IN1(n1489), .SEL(pc[3]), .F(n1491) );
  MUX U1516 ( .IN0(inst_mem_in_wire[1880]), .IN1(inst_mem_in_wire[1912]), 
        .SEL(pc[2]), .F(n1492) );
  MUX U1517 ( .IN0(inst_mem_in_wire[1816]), .IN1(inst_mem_in_wire[1848]), 
        .SEL(pc[2]), .F(n1493) );
  MUX U1518 ( .IN0(n1493), .IN1(n1492), .SEL(pc[3]), .F(n1494) );
  MUX U1519 ( .IN0(n1494), .IN1(n1491), .SEL(pc[4]), .F(n1495) );
  MUX U1520 ( .IN0(inst_mem_in_wire[1752]), .IN1(inst_mem_in_wire[1784]), 
        .SEL(pc[2]), .F(n1496) );
  MUX U1521 ( .IN0(inst_mem_in_wire[1688]), .IN1(inst_mem_in_wire[1720]), 
        .SEL(pc[2]), .F(n1497) );
  MUX U1522 ( .IN0(n1497), .IN1(n1496), .SEL(pc[3]), .F(n1498) );
  MUX U1523 ( .IN0(inst_mem_in_wire[1624]), .IN1(inst_mem_in_wire[1656]), 
        .SEL(pc[2]), .F(n1499) );
  MUX U1524 ( .IN0(inst_mem_in_wire[1560]), .IN1(inst_mem_in_wire[1592]), 
        .SEL(pc[2]), .F(n1500) );
  MUX U1525 ( .IN0(n1500), .IN1(n1499), .SEL(pc[3]), .F(n1501) );
  MUX U1526 ( .IN0(n1501), .IN1(n1498), .SEL(pc[4]), .F(n1502) );
  MUX U1527 ( .IN0(n1502), .IN1(n1495), .SEL(pc[5]), .F(n1503) );
  MUX U1528 ( .IN0(inst_mem_in_wire[1496]), .IN1(inst_mem_in_wire[1528]), 
        .SEL(pc[2]), .F(n1504) );
  MUX U1529 ( .IN0(inst_mem_in_wire[1432]), .IN1(inst_mem_in_wire[1464]), 
        .SEL(pc[2]), .F(n1505) );
  MUX U1530 ( .IN0(n1505), .IN1(n1504), .SEL(pc[3]), .F(n1506) );
  MUX U1531 ( .IN0(inst_mem_in_wire[1368]), .IN1(inst_mem_in_wire[1400]), 
        .SEL(pc[2]), .F(n1507) );
  MUX U1532 ( .IN0(inst_mem_in_wire[1304]), .IN1(inst_mem_in_wire[1336]), 
        .SEL(pc[2]), .F(n1508) );
  MUX U1533 ( .IN0(n1508), .IN1(n1507), .SEL(pc[3]), .F(n1509) );
  MUX U1534 ( .IN0(n1509), .IN1(n1506), .SEL(pc[4]), .F(n1510) );
  MUX U1535 ( .IN0(inst_mem_in_wire[1240]), .IN1(inst_mem_in_wire[1272]), 
        .SEL(pc[2]), .F(n1511) );
  MUX U1536 ( .IN0(inst_mem_in_wire[1176]), .IN1(inst_mem_in_wire[1208]), 
        .SEL(pc[2]), .F(n1512) );
  MUX U1537 ( .IN0(n1512), .IN1(n1511), .SEL(pc[3]), .F(n1513) );
  MUX U1538 ( .IN0(inst_mem_in_wire[1112]), .IN1(inst_mem_in_wire[1144]), 
        .SEL(pc[2]), .F(n1514) );
  MUX U1539 ( .IN0(inst_mem_in_wire[1048]), .IN1(inst_mem_in_wire[1080]), 
        .SEL(pc[2]), .F(n1515) );
  MUX U1540 ( .IN0(n1515), .IN1(n1514), .SEL(pc[3]), .F(n1516) );
  MUX U1541 ( .IN0(n1516), .IN1(n1513), .SEL(pc[4]), .F(n1517) );
  MUX U1542 ( .IN0(n1517), .IN1(n1510), .SEL(pc[5]), .F(n1518) );
  MUX U1543 ( .IN0(n1518), .IN1(n1503), .SEL(pc[6]), .F(n1519) );
  MUX U1544 ( .IN0(inst_mem_in_wire[984]), .IN1(inst_mem_in_wire[1016]), .SEL(
        pc[2]), .F(n1520) );
  MUX U1545 ( .IN0(inst_mem_in_wire[920]), .IN1(inst_mem_in_wire[952]), .SEL(
        pc[2]), .F(n1521) );
  MUX U1546 ( .IN0(n1521), .IN1(n1520), .SEL(pc[3]), .F(n1522) );
  MUX U1547 ( .IN0(inst_mem_in_wire[856]), .IN1(inst_mem_in_wire[888]), .SEL(
        pc[2]), .F(n1523) );
  MUX U1548 ( .IN0(inst_mem_in_wire[792]), .IN1(inst_mem_in_wire[824]), .SEL(
        pc[2]), .F(n1524) );
  MUX U1549 ( .IN0(n1524), .IN1(n1523), .SEL(pc[3]), .F(n1525) );
  MUX U1550 ( .IN0(n1525), .IN1(n1522), .SEL(pc[4]), .F(n1526) );
  MUX U1551 ( .IN0(inst_mem_in_wire[728]), .IN1(inst_mem_in_wire[760]), .SEL(
        pc[2]), .F(n1527) );
  MUX U1552 ( .IN0(inst_mem_in_wire[664]), .IN1(inst_mem_in_wire[696]), .SEL(
        pc[2]), .F(n1528) );
  MUX U1553 ( .IN0(n1528), .IN1(n1527), .SEL(pc[3]), .F(n1529) );
  MUX U1554 ( .IN0(inst_mem_in_wire[600]), .IN1(inst_mem_in_wire[632]), .SEL(
        pc[2]), .F(n1530) );
  MUX U1555 ( .IN0(inst_mem_in_wire[536]), .IN1(inst_mem_in_wire[568]), .SEL(
        pc[2]), .F(n1531) );
  MUX U1556 ( .IN0(n1531), .IN1(n1530), .SEL(pc[3]), .F(n1532) );
  MUX U1557 ( .IN0(n1532), .IN1(n1529), .SEL(pc[4]), .F(n1533) );
  MUX U1558 ( .IN0(n1533), .IN1(n1526), .SEL(pc[5]), .F(n1534) );
  MUX U1559 ( .IN0(inst_mem_in_wire[472]), .IN1(inst_mem_in_wire[504]), .SEL(
        pc[2]), .F(n1535) );
  MUX U1560 ( .IN0(inst_mem_in_wire[408]), .IN1(inst_mem_in_wire[440]), .SEL(
        pc[2]), .F(n1536) );
  MUX U1561 ( .IN0(n1536), .IN1(n1535), .SEL(pc[3]), .F(n1537) );
  MUX U1562 ( .IN0(inst_mem_in_wire[344]), .IN1(inst_mem_in_wire[376]), .SEL(
        pc[2]), .F(n1538) );
  MUX U1563 ( .IN0(inst_mem_in_wire[280]), .IN1(inst_mem_in_wire[312]), .SEL(
        pc[2]), .F(n1539) );
  MUX U1564 ( .IN0(n1539), .IN1(n1538), .SEL(pc[3]), .F(n1540) );
  MUX U1565 ( .IN0(n1540), .IN1(n1537), .SEL(pc[4]), .F(n1541) );
  MUX U1566 ( .IN0(inst_mem_in_wire[216]), .IN1(inst_mem_in_wire[248]), .SEL(
        pc[2]), .F(n1542) );
  MUX U1567 ( .IN0(inst_mem_in_wire[152]), .IN1(inst_mem_in_wire[184]), .SEL(
        pc[2]), .F(n1543) );
  MUX U1568 ( .IN0(n1543), .IN1(n1542), .SEL(pc[3]), .F(n1544) );
  MUX U1569 ( .IN0(inst_mem_in_wire[88]), .IN1(inst_mem_in_wire[120]), .SEL(
        pc[2]), .F(n1545) );
  MUX U1570 ( .IN0(inst_mem_in_wire[24]), .IN1(inst_mem_in_wire[56]), .SEL(
        pc[2]), .F(n1546) );
  MUX U1571 ( .IN0(n1546), .IN1(n1545), .SEL(pc[3]), .F(n1547) );
  MUX U1572 ( .IN0(n1547), .IN1(n1544), .SEL(pc[4]), .F(n1548) );
  MUX U1573 ( .IN0(n1548), .IN1(n1541), .SEL(pc[5]), .F(n1549) );
  MUX U1574 ( .IN0(n1549), .IN1(n1534), .SEL(pc[6]), .F(n1550) );
  MUX U1575 ( .IN0(n1550), .IN1(n1519), .SEL(pc[7]), .F(opcode[24]) );
  MUX U1576 ( .IN0(inst_mem_in_wire[2009]), .IN1(inst_mem_in_wire[2041]), 
        .SEL(pc[2]), .F(n1551) );
  MUX U1577 ( .IN0(inst_mem_in_wire[1945]), .IN1(inst_mem_in_wire[1977]), 
        .SEL(pc[2]), .F(n1552) );
  MUX U1578 ( .IN0(n1552), .IN1(n1551), .SEL(pc[3]), .F(n1553) );
  MUX U1579 ( .IN0(inst_mem_in_wire[1881]), .IN1(inst_mem_in_wire[1913]), 
        .SEL(pc[2]), .F(n1554) );
  MUX U1580 ( .IN0(inst_mem_in_wire[1817]), .IN1(inst_mem_in_wire[1849]), 
        .SEL(pc[2]), .F(n1555) );
  MUX U1581 ( .IN0(n1555), .IN1(n1554), .SEL(pc[3]), .F(n1556) );
  MUX U1582 ( .IN0(n1556), .IN1(n1553), .SEL(pc[4]), .F(n1557) );
  MUX U1583 ( .IN0(inst_mem_in_wire[1753]), .IN1(inst_mem_in_wire[1785]), 
        .SEL(pc[2]), .F(n1558) );
  MUX U1584 ( .IN0(inst_mem_in_wire[1689]), .IN1(inst_mem_in_wire[1721]), 
        .SEL(pc[2]), .F(n1559) );
  MUX U1585 ( .IN0(n1559), .IN1(n1558), .SEL(pc[3]), .F(n1560) );
  MUX U1586 ( .IN0(inst_mem_in_wire[1625]), .IN1(inst_mem_in_wire[1657]), 
        .SEL(pc[2]), .F(n1561) );
  MUX U1587 ( .IN0(inst_mem_in_wire[1561]), .IN1(inst_mem_in_wire[1593]), 
        .SEL(pc[2]), .F(n1562) );
  MUX U1588 ( .IN0(n1562), .IN1(n1561), .SEL(pc[3]), .F(n1563) );
  MUX U1589 ( .IN0(n1563), .IN1(n1560), .SEL(pc[4]), .F(n1564) );
  MUX U1590 ( .IN0(n1564), .IN1(n1557), .SEL(pc[5]), .F(n1565) );
  MUX U1591 ( .IN0(inst_mem_in_wire[1497]), .IN1(inst_mem_in_wire[1529]), 
        .SEL(pc[2]), .F(n1566) );
  MUX U1592 ( .IN0(inst_mem_in_wire[1433]), .IN1(inst_mem_in_wire[1465]), 
        .SEL(pc[2]), .F(n1567) );
  MUX U1593 ( .IN0(n1567), .IN1(n1566), .SEL(pc[3]), .F(n1568) );
  MUX U1594 ( .IN0(inst_mem_in_wire[1369]), .IN1(inst_mem_in_wire[1401]), 
        .SEL(pc[2]), .F(n1569) );
  MUX U1595 ( .IN0(inst_mem_in_wire[1305]), .IN1(inst_mem_in_wire[1337]), 
        .SEL(pc[2]), .F(n1570) );
  MUX U1596 ( .IN0(n1570), .IN1(n1569), .SEL(pc[3]), .F(n1571) );
  MUX U1597 ( .IN0(n1571), .IN1(n1568), .SEL(pc[4]), .F(n1572) );
  MUX U1598 ( .IN0(inst_mem_in_wire[1241]), .IN1(inst_mem_in_wire[1273]), 
        .SEL(pc[2]), .F(n1573) );
  MUX U1599 ( .IN0(inst_mem_in_wire[1177]), .IN1(inst_mem_in_wire[1209]), 
        .SEL(pc[2]), .F(n1574) );
  MUX U1600 ( .IN0(n1574), .IN1(n1573), .SEL(pc[3]), .F(n1575) );
  MUX U1601 ( .IN0(inst_mem_in_wire[1113]), .IN1(inst_mem_in_wire[1145]), 
        .SEL(pc[2]), .F(n1576) );
  MUX U1602 ( .IN0(inst_mem_in_wire[1049]), .IN1(inst_mem_in_wire[1081]), 
        .SEL(pc[2]), .F(n1577) );
  MUX U1603 ( .IN0(n1577), .IN1(n1576), .SEL(pc[3]), .F(n1578) );
  MUX U1604 ( .IN0(n1578), .IN1(n1575), .SEL(pc[4]), .F(n1579) );
  MUX U1605 ( .IN0(n1579), .IN1(n1572), .SEL(pc[5]), .F(n1580) );
  MUX U1606 ( .IN0(n1580), .IN1(n1565), .SEL(pc[6]), .F(n1581) );
  MUX U1607 ( .IN0(inst_mem_in_wire[985]), .IN1(inst_mem_in_wire[1017]), .SEL(
        pc[2]), .F(n1582) );
  MUX U1608 ( .IN0(inst_mem_in_wire[921]), .IN1(inst_mem_in_wire[953]), .SEL(
        pc[2]), .F(n1583) );
  MUX U1609 ( .IN0(n1583), .IN1(n1582), .SEL(pc[3]), .F(n1584) );
  MUX U1610 ( .IN0(inst_mem_in_wire[857]), .IN1(inst_mem_in_wire[889]), .SEL(
        pc[2]), .F(n1585) );
  MUX U1611 ( .IN0(inst_mem_in_wire[793]), .IN1(inst_mem_in_wire[825]), .SEL(
        pc[2]), .F(n1586) );
  MUX U1612 ( .IN0(n1586), .IN1(n1585), .SEL(pc[3]), .F(n1587) );
  MUX U1613 ( .IN0(n1587), .IN1(n1584), .SEL(pc[4]), .F(n1588) );
  MUX U1614 ( .IN0(inst_mem_in_wire[729]), .IN1(inst_mem_in_wire[761]), .SEL(
        pc[2]), .F(n1589) );
  MUX U1615 ( .IN0(inst_mem_in_wire[665]), .IN1(inst_mem_in_wire[697]), .SEL(
        pc[2]), .F(n1590) );
  MUX U1616 ( .IN0(n1590), .IN1(n1589), .SEL(pc[3]), .F(n1591) );
  MUX U1617 ( .IN0(inst_mem_in_wire[601]), .IN1(inst_mem_in_wire[633]), .SEL(
        pc[2]), .F(n1592) );
  MUX U1618 ( .IN0(inst_mem_in_wire[537]), .IN1(inst_mem_in_wire[569]), .SEL(
        pc[2]), .F(n1593) );
  MUX U1619 ( .IN0(n1593), .IN1(n1592), .SEL(pc[3]), .F(n1594) );
  MUX U1620 ( .IN0(n1594), .IN1(n1591), .SEL(pc[4]), .F(n1595) );
  MUX U1621 ( .IN0(n1595), .IN1(n1588), .SEL(pc[5]), .F(n1596) );
  MUX U1622 ( .IN0(inst_mem_in_wire[473]), .IN1(inst_mem_in_wire[505]), .SEL(
        pc[2]), .F(n1597) );
  MUX U1623 ( .IN0(inst_mem_in_wire[409]), .IN1(inst_mem_in_wire[441]), .SEL(
        pc[2]), .F(n1598) );
  MUX U1624 ( .IN0(n1598), .IN1(n1597), .SEL(pc[3]), .F(n1599) );
  MUX U1625 ( .IN0(inst_mem_in_wire[345]), .IN1(inst_mem_in_wire[377]), .SEL(
        pc[2]), .F(n1600) );
  MUX U1626 ( .IN0(inst_mem_in_wire[281]), .IN1(inst_mem_in_wire[313]), .SEL(
        pc[2]), .F(n1601) );
  MUX U1627 ( .IN0(n1601), .IN1(n1600), .SEL(pc[3]), .F(n1602) );
  MUX U1628 ( .IN0(n1602), .IN1(n1599), .SEL(pc[4]), .F(n1603) );
  MUX U1629 ( .IN0(inst_mem_in_wire[217]), .IN1(inst_mem_in_wire[249]), .SEL(
        pc[2]), .F(n1604) );
  MUX U1630 ( .IN0(inst_mem_in_wire[153]), .IN1(inst_mem_in_wire[185]), .SEL(
        pc[2]), .F(n1605) );
  MUX U1631 ( .IN0(n1605), .IN1(n1604), .SEL(pc[3]), .F(n1606) );
  MUX U1632 ( .IN0(inst_mem_in_wire[89]), .IN1(inst_mem_in_wire[121]), .SEL(
        pc[2]), .F(n1607) );
  MUX U1633 ( .IN0(inst_mem_in_wire[25]), .IN1(inst_mem_in_wire[57]), .SEL(
        pc[2]), .F(n1608) );
  MUX U1634 ( .IN0(n1608), .IN1(n1607), .SEL(pc[3]), .F(n1609) );
  MUX U1635 ( .IN0(n1609), .IN1(n1606), .SEL(pc[4]), .F(n1610) );
  MUX U1636 ( .IN0(n1610), .IN1(n1603), .SEL(pc[5]), .F(n1611) );
  MUX U1637 ( .IN0(n1611), .IN1(n1596), .SEL(pc[6]), .F(n1612) );
  MUX U1638 ( .IN0(n1612), .IN1(n1581), .SEL(pc[7]), .F(opcode[25]) );
  MUX U1639 ( .IN0(inst_mem_in_wire[2010]), .IN1(inst_mem_in_wire[2042]), 
        .SEL(pc[2]), .F(n1613) );
  MUX U1640 ( .IN0(inst_mem_in_wire[1946]), .IN1(inst_mem_in_wire[1978]), 
        .SEL(pc[2]), .F(n1614) );
  MUX U1641 ( .IN0(n1614), .IN1(n1613), .SEL(pc[3]), .F(n1615) );
  MUX U1642 ( .IN0(inst_mem_in_wire[1882]), .IN1(inst_mem_in_wire[1914]), 
        .SEL(pc[2]), .F(n1616) );
  MUX U1643 ( .IN0(inst_mem_in_wire[1818]), .IN1(inst_mem_in_wire[1850]), 
        .SEL(pc[2]), .F(n1617) );
  MUX U1644 ( .IN0(n1617), .IN1(n1616), .SEL(pc[3]), .F(n1618) );
  MUX U1645 ( .IN0(n1618), .IN1(n1615), .SEL(pc[4]), .F(n1619) );
  MUX U1646 ( .IN0(inst_mem_in_wire[1754]), .IN1(inst_mem_in_wire[1786]), 
        .SEL(pc[2]), .F(n1620) );
  MUX U1647 ( .IN0(inst_mem_in_wire[1690]), .IN1(inst_mem_in_wire[1722]), 
        .SEL(pc[2]), .F(n1621) );
  MUX U1648 ( .IN0(n1621), .IN1(n1620), .SEL(pc[3]), .F(n1622) );
  MUX U1649 ( .IN0(inst_mem_in_wire[1626]), .IN1(inst_mem_in_wire[1658]), 
        .SEL(pc[2]), .F(n1623) );
  MUX U1650 ( .IN0(inst_mem_in_wire[1562]), .IN1(inst_mem_in_wire[1594]), 
        .SEL(pc[2]), .F(n1624) );
  MUX U1651 ( .IN0(n1624), .IN1(n1623), .SEL(pc[3]), .F(n1625) );
  MUX U1652 ( .IN0(n1625), .IN1(n1622), .SEL(pc[4]), .F(n1626) );
  MUX U1653 ( .IN0(n1626), .IN1(n1619), .SEL(pc[5]), .F(n1627) );
  MUX U1654 ( .IN0(inst_mem_in_wire[1498]), .IN1(inst_mem_in_wire[1530]), 
        .SEL(pc[2]), .F(n1628) );
  MUX U1655 ( .IN0(inst_mem_in_wire[1434]), .IN1(inst_mem_in_wire[1466]), 
        .SEL(pc[2]), .F(n1629) );
  MUX U1656 ( .IN0(n1629), .IN1(n1628), .SEL(pc[3]), .F(n1630) );
  MUX U1657 ( .IN0(inst_mem_in_wire[1370]), .IN1(inst_mem_in_wire[1402]), 
        .SEL(pc[2]), .F(n1631) );
  MUX U1658 ( .IN0(inst_mem_in_wire[1306]), .IN1(inst_mem_in_wire[1338]), 
        .SEL(pc[2]), .F(n1632) );
  MUX U1659 ( .IN0(n1632), .IN1(n1631), .SEL(pc[3]), .F(n1633) );
  MUX U1660 ( .IN0(n1633), .IN1(n1630), .SEL(pc[4]), .F(n1634) );
  MUX U1661 ( .IN0(inst_mem_in_wire[1242]), .IN1(inst_mem_in_wire[1274]), 
        .SEL(pc[2]), .F(n1635) );
  MUX U1662 ( .IN0(inst_mem_in_wire[1178]), .IN1(inst_mem_in_wire[1210]), 
        .SEL(pc[2]), .F(n1636) );
  MUX U1663 ( .IN0(n1636), .IN1(n1635), .SEL(pc[3]), .F(n1637) );
  MUX U1664 ( .IN0(inst_mem_in_wire[1114]), .IN1(inst_mem_in_wire[1146]), 
        .SEL(pc[2]), .F(n1638) );
  MUX U1665 ( .IN0(inst_mem_in_wire[1050]), .IN1(inst_mem_in_wire[1082]), 
        .SEL(pc[2]), .F(n1639) );
  MUX U1666 ( .IN0(n1639), .IN1(n1638), .SEL(pc[3]), .F(n1640) );
  MUX U1667 ( .IN0(n1640), .IN1(n1637), .SEL(pc[4]), .F(n1641) );
  MUX U1668 ( .IN0(n1641), .IN1(n1634), .SEL(pc[5]), .F(n1642) );
  MUX U1669 ( .IN0(n1642), .IN1(n1627), .SEL(pc[6]), .F(n1643) );
  MUX U1670 ( .IN0(inst_mem_in_wire[986]), .IN1(inst_mem_in_wire[1018]), .SEL(
        pc[2]), .F(n1644) );
  MUX U1671 ( .IN0(inst_mem_in_wire[922]), .IN1(inst_mem_in_wire[954]), .SEL(
        pc[2]), .F(n1645) );
  MUX U1672 ( .IN0(n1645), .IN1(n1644), .SEL(pc[3]), .F(n1646) );
  MUX U1673 ( .IN0(inst_mem_in_wire[858]), .IN1(inst_mem_in_wire[890]), .SEL(
        pc[2]), .F(n1647) );
  MUX U1674 ( .IN0(inst_mem_in_wire[794]), .IN1(inst_mem_in_wire[826]), .SEL(
        pc[2]), .F(n1648) );
  MUX U1675 ( .IN0(n1648), .IN1(n1647), .SEL(pc[3]), .F(n1649) );
  MUX U1676 ( .IN0(n1649), .IN1(n1646), .SEL(pc[4]), .F(n1650) );
  MUX U1677 ( .IN0(inst_mem_in_wire[730]), .IN1(inst_mem_in_wire[762]), .SEL(
        pc[2]), .F(n1651) );
  MUX U1678 ( .IN0(inst_mem_in_wire[666]), .IN1(inst_mem_in_wire[698]), .SEL(
        pc[2]), .F(n1652) );
  MUX U1679 ( .IN0(n1652), .IN1(n1651), .SEL(pc[3]), .F(n1653) );
  MUX U1680 ( .IN0(inst_mem_in_wire[602]), .IN1(inst_mem_in_wire[634]), .SEL(
        pc[2]), .F(n1654) );
  MUX U1681 ( .IN0(inst_mem_in_wire[538]), .IN1(inst_mem_in_wire[570]), .SEL(
        pc[2]), .F(n1655) );
  MUX U1682 ( .IN0(n1655), .IN1(n1654), .SEL(pc[3]), .F(n1656) );
  MUX U1683 ( .IN0(n1656), .IN1(n1653), .SEL(pc[4]), .F(n1657) );
  MUX U1684 ( .IN0(n1657), .IN1(n1650), .SEL(pc[5]), .F(n1658) );
  MUX U1685 ( .IN0(inst_mem_in_wire[474]), .IN1(inst_mem_in_wire[506]), .SEL(
        pc[2]), .F(n1659) );
  MUX U1686 ( .IN0(inst_mem_in_wire[410]), .IN1(inst_mem_in_wire[442]), .SEL(
        pc[2]), .F(n1660) );
  MUX U1687 ( .IN0(n1660), .IN1(n1659), .SEL(pc[3]), .F(n1661) );
  MUX U1688 ( .IN0(inst_mem_in_wire[346]), .IN1(inst_mem_in_wire[378]), .SEL(
        pc[2]), .F(n1662) );
  MUX U1689 ( .IN0(inst_mem_in_wire[282]), .IN1(inst_mem_in_wire[314]), .SEL(
        pc[2]), .F(n1663) );
  MUX U1690 ( .IN0(n1663), .IN1(n1662), .SEL(pc[3]), .F(n1664) );
  MUX U1691 ( .IN0(n1664), .IN1(n1661), .SEL(pc[4]), .F(n1665) );
  MUX U1692 ( .IN0(inst_mem_in_wire[218]), .IN1(inst_mem_in_wire[250]), .SEL(
        pc[2]), .F(n1666) );
  MUX U1693 ( .IN0(inst_mem_in_wire[154]), .IN1(inst_mem_in_wire[186]), .SEL(
        pc[2]), .F(n1667) );
  MUX U1694 ( .IN0(n1667), .IN1(n1666), .SEL(pc[3]), .F(n1668) );
  MUX U1695 ( .IN0(inst_mem_in_wire[90]), .IN1(inst_mem_in_wire[122]), .SEL(
        pc[2]), .F(n1669) );
  MUX U1696 ( .IN0(inst_mem_in_wire[26]), .IN1(inst_mem_in_wire[58]), .SEL(
        pc[2]), .F(n1670) );
  MUX U1697 ( .IN0(n1670), .IN1(n1669), .SEL(pc[3]), .F(n1671) );
  MUX U1698 ( .IN0(n1671), .IN1(n1668), .SEL(pc[4]), .F(n1672) );
  MUX U1699 ( .IN0(n1672), .IN1(n1665), .SEL(pc[5]), .F(n1673) );
  MUX U1700 ( .IN0(n1673), .IN1(n1658), .SEL(pc[6]), .F(n1674) );
  MUX U1701 ( .IN0(n1674), .IN1(n1643), .SEL(pc[7]), .F(opcode[26]) );
  MUX U1702 ( .IN0(inst_mem_in_wire[2011]), .IN1(inst_mem_in_wire[2043]), 
        .SEL(pc[2]), .F(n1675) );
  MUX U1703 ( .IN0(inst_mem_in_wire[1947]), .IN1(inst_mem_in_wire[1979]), 
        .SEL(pc[2]), .F(n1676) );
  MUX U1704 ( .IN0(n1676), .IN1(n1675), .SEL(pc[3]), .F(n1677) );
  MUX U1705 ( .IN0(inst_mem_in_wire[1883]), .IN1(inst_mem_in_wire[1915]), 
        .SEL(pc[2]), .F(n1678) );
  MUX U1706 ( .IN0(inst_mem_in_wire[1819]), .IN1(inst_mem_in_wire[1851]), 
        .SEL(pc[2]), .F(n1679) );
  MUX U1707 ( .IN0(n1679), .IN1(n1678), .SEL(pc[3]), .F(n1680) );
  MUX U1708 ( .IN0(n1680), .IN1(n1677), .SEL(pc[4]), .F(n1681) );
  MUX U1709 ( .IN0(inst_mem_in_wire[1755]), .IN1(inst_mem_in_wire[1787]), 
        .SEL(pc[2]), .F(n1682) );
  MUX U1710 ( .IN0(inst_mem_in_wire[1691]), .IN1(inst_mem_in_wire[1723]), 
        .SEL(pc[2]), .F(n1683) );
  MUX U1711 ( .IN0(n1683), .IN1(n1682), .SEL(pc[3]), .F(n1684) );
  MUX U1712 ( .IN0(inst_mem_in_wire[1627]), .IN1(inst_mem_in_wire[1659]), 
        .SEL(pc[2]), .F(n1685) );
  MUX U1713 ( .IN0(inst_mem_in_wire[1563]), .IN1(inst_mem_in_wire[1595]), 
        .SEL(pc[2]), .F(n1686) );
  MUX U1714 ( .IN0(n1686), .IN1(n1685), .SEL(pc[3]), .F(n1687) );
  MUX U1715 ( .IN0(n1687), .IN1(n1684), .SEL(pc[4]), .F(n1688) );
  MUX U1716 ( .IN0(n1688), .IN1(n1681), .SEL(pc[5]), .F(n1689) );
  MUX U1717 ( .IN0(inst_mem_in_wire[1499]), .IN1(inst_mem_in_wire[1531]), 
        .SEL(pc[2]), .F(n1690) );
  MUX U1718 ( .IN0(inst_mem_in_wire[1435]), .IN1(inst_mem_in_wire[1467]), 
        .SEL(pc[2]), .F(n1691) );
  MUX U1719 ( .IN0(n1691), .IN1(n1690), .SEL(pc[3]), .F(n1692) );
  MUX U1720 ( .IN0(inst_mem_in_wire[1371]), .IN1(inst_mem_in_wire[1403]), 
        .SEL(pc[2]), .F(n1693) );
  MUX U1721 ( .IN0(inst_mem_in_wire[1307]), .IN1(inst_mem_in_wire[1339]), 
        .SEL(pc[2]), .F(n1694) );
  MUX U1722 ( .IN0(n1694), .IN1(n1693), .SEL(pc[3]), .F(n1695) );
  MUX U1723 ( .IN0(n1695), .IN1(n1692), .SEL(pc[4]), .F(n1696) );
  MUX U1724 ( .IN0(inst_mem_in_wire[1243]), .IN1(inst_mem_in_wire[1275]), 
        .SEL(pc[2]), .F(n1697) );
  MUX U1725 ( .IN0(inst_mem_in_wire[1179]), .IN1(inst_mem_in_wire[1211]), 
        .SEL(pc[2]), .F(n1698) );
  MUX U1726 ( .IN0(n1698), .IN1(n1697), .SEL(pc[3]), .F(n1699) );
  MUX U1727 ( .IN0(inst_mem_in_wire[1115]), .IN1(inst_mem_in_wire[1147]), 
        .SEL(pc[2]), .F(n1700) );
  MUX U1728 ( .IN0(inst_mem_in_wire[1051]), .IN1(inst_mem_in_wire[1083]), 
        .SEL(pc[2]), .F(n1701) );
  MUX U1729 ( .IN0(n1701), .IN1(n1700), .SEL(pc[3]), .F(n1702) );
  MUX U1730 ( .IN0(n1702), .IN1(n1699), .SEL(pc[4]), .F(n1703) );
  MUX U1731 ( .IN0(n1703), .IN1(n1696), .SEL(pc[5]), .F(n1704) );
  MUX U1732 ( .IN0(n1704), .IN1(n1689), .SEL(pc[6]), .F(n1705) );
  MUX U1733 ( .IN0(inst_mem_in_wire[987]), .IN1(inst_mem_in_wire[1019]), .SEL(
        pc[2]), .F(n1706) );
  MUX U1734 ( .IN0(inst_mem_in_wire[923]), .IN1(inst_mem_in_wire[955]), .SEL(
        pc[2]), .F(n1707) );
  MUX U1735 ( .IN0(n1707), .IN1(n1706), .SEL(pc[3]), .F(n1708) );
  MUX U1736 ( .IN0(inst_mem_in_wire[859]), .IN1(inst_mem_in_wire[891]), .SEL(
        pc[2]), .F(n1709) );
  MUX U1737 ( .IN0(inst_mem_in_wire[795]), .IN1(inst_mem_in_wire[827]), .SEL(
        pc[2]), .F(n1710) );
  MUX U1738 ( .IN0(n1710), .IN1(n1709), .SEL(pc[3]), .F(n1711) );
  MUX U1739 ( .IN0(n1711), .IN1(n1708), .SEL(pc[4]), .F(n1712) );
  MUX U1740 ( .IN0(inst_mem_in_wire[731]), .IN1(inst_mem_in_wire[763]), .SEL(
        pc[2]), .F(n1713) );
  MUX U1741 ( .IN0(inst_mem_in_wire[667]), .IN1(inst_mem_in_wire[699]), .SEL(
        pc[2]), .F(n1714) );
  MUX U1742 ( .IN0(n1714), .IN1(n1713), .SEL(pc[3]), .F(n1715) );
  MUX U1743 ( .IN0(inst_mem_in_wire[603]), .IN1(inst_mem_in_wire[635]), .SEL(
        pc[2]), .F(n1716) );
  MUX U1744 ( .IN0(inst_mem_in_wire[539]), .IN1(inst_mem_in_wire[571]), .SEL(
        pc[2]), .F(n1717) );
  MUX U1745 ( .IN0(n1717), .IN1(n1716), .SEL(pc[3]), .F(n1718) );
  MUX U1746 ( .IN0(n1718), .IN1(n1715), .SEL(pc[4]), .F(n1719) );
  MUX U1747 ( .IN0(n1719), .IN1(n1712), .SEL(pc[5]), .F(n1720) );
  MUX U1748 ( .IN0(inst_mem_in_wire[475]), .IN1(inst_mem_in_wire[507]), .SEL(
        pc[2]), .F(n1721) );
  MUX U1749 ( .IN0(inst_mem_in_wire[411]), .IN1(inst_mem_in_wire[443]), .SEL(
        pc[2]), .F(n1722) );
  MUX U1750 ( .IN0(n1722), .IN1(n1721), .SEL(pc[3]), .F(n1723) );
  MUX U1751 ( .IN0(inst_mem_in_wire[347]), .IN1(inst_mem_in_wire[379]), .SEL(
        pc[2]), .F(n1724) );
  MUX U1752 ( .IN0(inst_mem_in_wire[283]), .IN1(inst_mem_in_wire[315]), .SEL(
        pc[2]), .F(n1725) );
  MUX U1753 ( .IN0(n1725), .IN1(n1724), .SEL(pc[3]), .F(n1726) );
  MUX U1754 ( .IN0(n1726), .IN1(n1723), .SEL(pc[4]), .F(n1727) );
  MUX U1755 ( .IN0(inst_mem_in_wire[219]), .IN1(inst_mem_in_wire[251]), .SEL(
        pc[2]), .F(n1728) );
  MUX U1756 ( .IN0(inst_mem_in_wire[155]), .IN1(inst_mem_in_wire[187]), .SEL(
        pc[2]), .F(n1729) );
  MUX U1757 ( .IN0(n1729), .IN1(n1728), .SEL(pc[3]), .F(n1730) );
  MUX U1758 ( .IN0(inst_mem_in_wire[91]), .IN1(inst_mem_in_wire[123]), .SEL(
        pc[2]), .F(n1731) );
  MUX U1759 ( .IN0(inst_mem_in_wire[27]), .IN1(inst_mem_in_wire[59]), .SEL(
        pc[2]), .F(n1732) );
  MUX U1760 ( .IN0(n1732), .IN1(n1731), .SEL(pc[3]), .F(n1733) );
  MUX U1761 ( .IN0(n1733), .IN1(n1730), .SEL(pc[4]), .F(n1734) );
  MUX U1762 ( .IN0(n1734), .IN1(n1727), .SEL(pc[5]), .F(n1735) );
  MUX U1763 ( .IN0(n1735), .IN1(n1720), .SEL(pc[6]), .F(n1736) );
  MUX U1764 ( .IN0(n1736), .IN1(n1705), .SEL(pc[7]), .F(opcode[27]) );
  MUX U1765 ( .IN0(inst_mem_in_wire[2012]), .IN1(inst_mem_in_wire[2044]), 
        .SEL(pc[2]), .F(n1737) );
  MUX U1766 ( .IN0(inst_mem_in_wire[1948]), .IN1(inst_mem_in_wire[1980]), 
        .SEL(pc[2]), .F(n1738) );
  MUX U1767 ( .IN0(n1738), .IN1(n1737), .SEL(pc[3]), .F(n1739) );
  MUX U1768 ( .IN0(inst_mem_in_wire[1884]), .IN1(inst_mem_in_wire[1916]), 
        .SEL(pc[2]), .F(n1740) );
  MUX U1769 ( .IN0(inst_mem_in_wire[1820]), .IN1(inst_mem_in_wire[1852]), 
        .SEL(pc[2]), .F(n1741) );
  MUX U1770 ( .IN0(n1741), .IN1(n1740), .SEL(pc[3]), .F(n1742) );
  MUX U1771 ( .IN0(n1742), .IN1(n1739), .SEL(pc[4]), .F(n1743) );
  MUX U1772 ( .IN0(inst_mem_in_wire[1756]), .IN1(inst_mem_in_wire[1788]), 
        .SEL(pc[2]), .F(n1744) );
  MUX U1773 ( .IN0(inst_mem_in_wire[1692]), .IN1(inst_mem_in_wire[1724]), 
        .SEL(pc[2]), .F(n1745) );
  MUX U1774 ( .IN0(n1745), .IN1(n1744), .SEL(pc[3]), .F(n1746) );
  MUX U1775 ( .IN0(inst_mem_in_wire[1628]), .IN1(inst_mem_in_wire[1660]), 
        .SEL(pc[2]), .F(n1747) );
  MUX U1776 ( .IN0(inst_mem_in_wire[1564]), .IN1(inst_mem_in_wire[1596]), 
        .SEL(pc[2]), .F(n1748) );
  MUX U1777 ( .IN0(n1748), .IN1(n1747), .SEL(pc[3]), .F(n1749) );
  MUX U1778 ( .IN0(n1749), .IN1(n1746), .SEL(pc[4]), .F(n1750) );
  MUX U1779 ( .IN0(n1750), .IN1(n1743), .SEL(pc[5]), .F(n1751) );
  MUX U1780 ( .IN0(inst_mem_in_wire[1500]), .IN1(inst_mem_in_wire[1532]), 
        .SEL(pc[2]), .F(n1752) );
  MUX U1781 ( .IN0(inst_mem_in_wire[1436]), .IN1(inst_mem_in_wire[1468]), 
        .SEL(pc[2]), .F(n1753) );
  MUX U1782 ( .IN0(n1753), .IN1(n1752), .SEL(pc[3]), .F(n1754) );
  MUX U1783 ( .IN0(inst_mem_in_wire[1372]), .IN1(inst_mem_in_wire[1404]), 
        .SEL(pc[2]), .F(n1755) );
  MUX U1784 ( .IN0(inst_mem_in_wire[1308]), .IN1(inst_mem_in_wire[1340]), 
        .SEL(pc[2]), .F(n1756) );
  MUX U1785 ( .IN0(n1756), .IN1(n1755), .SEL(pc[3]), .F(n1757) );
  MUX U1786 ( .IN0(n1757), .IN1(n1754), .SEL(pc[4]), .F(n1758) );
  MUX U1787 ( .IN0(inst_mem_in_wire[1244]), .IN1(inst_mem_in_wire[1276]), 
        .SEL(pc[2]), .F(n1759) );
  MUX U1788 ( .IN0(inst_mem_in_wire[1180]), .IN1(inst_mem_in_wire[1212]), 
        .SEL(pc[2]), .F(n1760) );
  MUX U1789 ( .IN0(n1760), .IN1(n1759), .SEL(pc[3]), .F(n1761) );
  MUX U1790 ( .IN0(inst_mem_in_wire[1116]), .IN1(inst_mem_in_wire[1148]), 
        .SEL(pc[2]), .F(n1762) );
  MUX U1791 ( .IN0(inst_mem_in_wire[1052]), .IN1(inst_mem_in_wire[1084]), 
        .SEL(pc[2]), .F(n1763) );
  MUX U1792 ( .IN0(n1763), .IN1(n1762), .SEL(pc[3]), .F(n1764) );
  MUX U1793 ( .IN0(n1764), .IN1(n1761), .SEL(pc[4]), .F(n1765) );
  MUX U1794 ( .IN0(n1765), .IN1(n1758), .SEL(pc[5]), .F(n1766) );
  MUX U1795 ( .IN0(n1766), .IN1(n1751), .SEL(pc[6]), .F(n1767) );
  MUX U1796 ( .IN0(inst_mem_in_wire[988]), .IN1(inst_mem_in_wire[1020]), .SEL(
        pc[2]), .F(n1768) );
  MUX U1797 ( .IN0(inst_mem_in_wire[924]), .IN1(inst_mem_in_wire[956]), .SEL(
        pc[2]), .F(n1769) );
  MUX U1798 ( .IN0(n1769), .IN1(n1768), .SEL(pc[3]), .F(n1770) );
  MUX U1799 ( .IN0(inst_mem_in_wire[860]), .IN1(inst_mem_in_wire[892]), .SEL(
        pc[2]), .F(n1771) );
  MUX U1800 ( .IN0(inst_mem_in_wire[796]), .IN1(inst_mem_in_wire[828]), .SEL(
        pc[2]), .F(n1772) );
  MUX U1801 ( .IN0(n1772), .IN1(n1771), .SEL(pc[3]), .F(n1773) );
  MUX U1802 ( .IN0(n1773), .IN1(n1770), .SEL(pc[4]), .F(n1774) );
  MUX U1803 ( .IN0(inst_mem_in_wire[732]), .IN1(inst_mem_in_wire[764]), .SEL(
        pc[2]), .F(n1775) );
  MUX U1804 ( .IN0(inst_mem_in_wire[668]), .IN1(inst_mem_in_wire[700]), .SEL(
        pc[2]), .F(n1776) );
  MUX U1805 ( .IN0(n1776), .IN1(n1775), .SEL(pc[3]), .F(n1777) );
  MUX U1806 ( .IN0(inst_mem_in_wire[604]), .IN1(inst_mem_in_wire[636]), .SEL(
        pc[2]), .F(n1778) );
  MUX U1807 ( .IN0(inst_mem_in_wire[540]), .IN1(inst_mem_in_wire[572]), .SEL(
        pc[2]), .F(n1779) );
  MUX U1808 ( .IN0(n1779), .IN1(n1778), .SEL(pc[3]), .F(n1780) );
  MUX U1809 ( .IN0(n1780), .IN1(n1777), .SEL(pc[4]), .F(n1781) );
  MUX U1810 ( .IN0(n1781), .IN1(n1774), .SEL(pc[5]), .F(n1782) );
  MUX U1811 ( .IN0(inst_mem_in_wire[476]), .IN1(inst_mem_in_wire[508]), .SEL(
        pc[2]), .F(n1783) );
  MUX U1812 ( .IN0(inst_mem_in_wire[412]), .IN1(inst_mem_in_wire[444]), .SEL(
        pc[2]), .F(n1784) );
  MUX U1813 ( .IN0(n1784), .IN1(n1783), .SEL(pc[3]), .F(n1785) );
  MUX U1814 ( .IN0(inst_mem_in_wire[348]), .IN1(inst_mem_in_wire[380]), .SEL(
        pc[2]), .F(n1786) );
  MUX U1815 ( .IN0(inst_mem_in_wire[284]), .IN1(inst_mem_in_wire[316]), .SEL(
        pc[2]), .F(n1787) );
  MUX U1816 ( .IN0(n1787), .IN1(n1786), .SEL(pc[3]), .F(n1788) );
  MUX U1817 ( .IN0(n1788), .IN1(n1785), .SEL(pc[4]), .F(n1789) );
  MUX U1818 ( .IN0(inst_mem_in_wire[220]), .IN1(inst_mem_in_wire[252]), .SEL(
        pc[2]), .F(n1790) );
  MUX U1819 ( .IN0(inst_mem_in_wire[156]), .IN1(inst_mem_in_wire[188]), .SEL(
        pc[2]), .F(n1791) );
  MUX U1820 ( .IN0(n1791), .IN1(n1790), .SEL(pc[3]), .F(n1792) );
  MUX U1821 ( .IN0(inst_mem_in_wire[92]), .IN1(inst_mem_in_wire[124]), .SEL(
        pc[2]), .F(n1793) );
  MUX U1822 ( .IN0(inst_mem_in_wire[28]), .IN1(inst_mem_in_wire[60]), .SEL(
        pc[2]), .F(n1794) );
  MUX U1823 ( .IN0(n1794), .IN1(n1793), .SEL(pc[3]), .F(n1795) );
  MUX U1824 ( .IN0(n1795), .IN1(n1792), .SEL(pc[4]), .F(n1796) );
  MUX U1825 ( .IN0(n1796), .IN1(n1789), .SEL(pc[5]), .F(n1797) );
  MUX U1826 ( .IN0(n1797), .IN1(n1782), .SEL(pc[6]), .F(n1798) );
  MUX U1827 ( .IN0(n1798), .IN1(n1767), .SEL(pc[7]), .F(opcode[28]) );
  MUX U1828 ( .IN0(inst_mem_in_wire[2013]), .IN1(inst_mem_in_wire[2045]), 
        .SEL(pc[2]), .F(n1799) );
  MUX U1829 ( .IN0(inst_mem_in_wire[1949]), .IN1(inst_mem_in_wire[1981]), 
        .SEL(pc[2]), .F(n1800) );
  MUX U1830 ( .IN0(n1800), .IN1(n1799), .SEL(pc[3]), .F(n1801) );
  MUX U1831 ( .IN0(inst_mem_in_wire[1885]), .IN1(inst_mem_in_wire[1917]), 
        .SEL(pc[2]), .F(n1802) );
  MUX U1832 ( .IN0(inst_mem_in_wire[1821]), .IN1(inst_mem_in_wire[1853]), 
        .SEL(pc[2]), .F(n1803) );
  MUX U1833 ( .IN0(n1803), .IN1(n1802), .SEL(pc[3]), .F(n1804) );
  MUX U1834 ( .IN0(n1804), .IN1(n1801), .SEL(pc[4]), .F(n1805) );
  MUX U1835 ( .IN0(inst_mem_in_wire[1757]), .IN1(inst_mem_in_wire[1789]), 
        .SEL(pc[2]), .F(n1806) );
  MUX U1836 ( .IN0(inst_mem_in_wire[1693]), .IN1(inst_mem_in_wire[1725]), 
        .SEL(pc[2]), .F(n1807) );
  MUX U1837 ( .IN0(n1807), .IN1(n1806), .SEL(pc[3]), .F(n1808) );
  MUX U1838 ( .IN0(inst_mem_in_wire[1629]), .IN1(inst_mem_in_wire[1661]), 
        .SEL(pc[2]), .F(n1809) );
  MUX U1839 ( .IN0(inst_mem_in_wire[1565]), .IN1(inst_mem_in_wire[1597]), 
        .SEL(pc[2]), .F(n1810) );
  MUX U1840 ( .IN0(n1810), .IN1(n1809), .SEL(pc[3]), .F(n1811) );
  MUX U1841 ( .IN0(n1811), .IN1(n1808), .SEL(pc[4]), .F(n1812) );
  MUX U1842 ( .IN0(n1812), .IN1(n1805), .SEL(pc[5]), .F(n1813) );
  MUX U1843 ( .IN0(inst_mem_in_wire[1501]), .IN1(inst_mem_in_wire[1533]), 
        .SEL(pc[2]), .F(n1814) );
  MUX U1844 ( .IN0(inst_mem_in_wire[1437]), .IN1(inst_mem_in_wire[1469]), 
        .SEL(pc[2]), .F(n1815) );
  MUX U1845 ( .IN0(n1815), .IN1(n1814), .SEL(pc[3]), .F(n1816) );
  MUX U1846 ( .IN0(inst_mem_in_wire[1373]), .IN1(inst_mem_in_wire[1405]), 
        .SEL(pc[2]), .F(n1817) );
  MUX U1847 ( .IN0(inst_mem_in_wire[1309]), .IN1(inst_mem_in_wire[1341]), 
        .SEL(pc[2]), .F(n1818) );
  MUX U1848 ( .IN0(n1818), .IN1(n1817), .SEL(pc[3]), .F(n1819) );
  MUX U1849 ( .IN0(n1819), .IN1(n1816), .SEL(pc[4]), .F(n1820) );
  MUX U1850 ( .IN0(inst_mem_in_wire[1245]), .IN1(inst_mem_in_wire[1277]), 
        .SEL(pc[2]), .F(n1821) );
  MUX U1851 ( .IN0(inst_mem_in_wire[1181]), .IN1(inst_mem_in_wire[1213]), 
        .SEL(pc[2]), .F(n1822) );
  MUX U1852 ( .IN0(n1822), .IN1(n1821), .SEL(pc[3]), .F(n1823) );
  MUX U1853 ( .IN0(inst_mem_in_wire[1117]), .IN1(inst_mem_in_wire[1149]), 
        .SEL(pc[2]), .F(n1824) );
  MUX U1854 ( .IN0(inst_mem_in_wire[1053]), .IN1(inst_mem_in_wire[1085]), 
        .SEL(pc[2]), .F(n1825) );
  MUX U1855 ( .IN0(n1825), .IN1(n1824), .SEL(pc[3]), .F(n1826) );
  MUX U1856 ( .IN0(n1826), .IN1(n1823), .SEL(pc[4]), .F(n1827) );
  MUX U1857 ( .IN0(n1827), .IN1(n1820), .SEL(pc[5]), .F(n1828) );
  MUX U1858 ( .IN0(n1828), .IN1(n1813), .SEL(pc[6]), .F(n1829) );
  MUX U1859 ( .IN0(inst_mem_in_wire[989]), .IN1(inst_mem_in_wire[1021]), .SEL(
        pc[2]), .F(n1830) );
  MUX U1860 ( .IN0(inst_mem_in_wire[925]), .IN1(inst_mem_in_wire[957]), .SEL(
        pc[2]), .F(n1831) );
  MUX U1861 ( .IN0(n1831), .IN1(n1830), .SEL(pc[3]), .F(n1832) );
  MUX U1862 ( .IN0(inst_mem_in_wire[861]), .IN1(inst_mem_in_wire[893]), .SEL(
        pc[2]), .F(n1833) );
  MUX U1863 ( .IN0(inst_mem_in_wire[797]), .IN1(inst_mem_in_wire[829]), .SEL(
        pc[2]), .F(n1834) );
  MUX U1864 ( .IN0(n1834), .IN1(n1833), .SEL(pc[3]), .F(n1835) );
  MUX U1865 ( .IN0(n1835), .IN1(n1832), .SEL(pc[4]), .F(n1836) );
  MUX U1866 ( .IN0(inst_mem_in_wire[733]), .IN1(inst_mem_in_wire[765]), .SEL(
        pc[2]), .F(n1837) );
  MUX U1867 ( .IN0(inst_mem_in_wire[669]), .IN1(inst_mem_in_wire[701]), .SEL(
        pc[2]), .F(n1838) );
  MUX U1868 ( .IN0(n1838), .IN1(n1837), .SEL(pc[3]), .F(n1839) );
  MUX U1869 ( .IN0(inst_mem_in_wire[605]), .IN1(inst_mem_in_wire[637]), .SEL(
        pc[2]), .F(n1840) );
  MUX U1870 ( .IN0(inst_mem_in_wire[541]), .IN1(inst_mem_in_wire[573]), .SEL(
        pc[2]), .F(n1841) );
  MUX U1871 ( .IN0(n1841), .IN1(n1840), .SEL(pc[3]), .F(n1842) );
  MUX U1872 ( .IN0(n1842), .IN1(n1839), .SEL(pc[4]), .F(n1843) );
  MUX U1873 ( .IN0(n1843), .IN1(n1836), .SEL(pc[5]), .F(n1844) );
  MUX U1874 ( .IN0(inst_mem_in_wire[477]), .IN1(inst_mem_in_wire[509]), .SEL(
        pc[2]), .F(n1845) );
  MUX U1875 ( .IN0(inst_mem_in_wire[413]), .IN1(inst_mem_in_wire[445]), .SEL(
        pc[2]), .F(n1846) );
  MUX U1876 ( .IN0(n1846), .IN1(n1845), .SEL(pc[3]), .F(n1847) );
  MUX U1877 ( .IN0(inst_mem_in_wire[349]), .IN1(inst_mem_in_wire[381]), .SEL(
        pc[2]), .F(n1848) );
  MUX U1878 ( .IN0(inst_mem_in_wire[285]), .IN1(inst_mem_in_wire[317]), .SEL(
        pc[2]), .F(n1849) );
  MUX U1879 ( .IN0(n1849), .IN1(n1848), .SEL(pc[3]), .F(n1850) );
  MUX U1880 ( .IN0(n1850), .IN1(n1847), .SEL(pc[4]), .F(n1851) );
  MUX U1881 ( .IN0(inst_mem_in_wire[221]), .IN1(inst_mem_in_wire[253]), .SEL(
        pc[2]), .F(n1852) );
  MUX U1882 ( .IN0(inst_mem_in_wire[157]), .IN1(inst_mem_in_wire[189]), .SEL(
        pc[2]), .F(n1853) );
  MUX U1883 ( .IN0(n1853), .IN1(n1852), .SEL(pc[3]), .F(n1854) );
  MUX U1884 ( .IN0(inst_mem_in_wire[93]), .IN1(inst_mem_in_wire[125]), .SEL(
        pc[2]), .F(n1855) );
  MUX U1885 ( .IN0(inst_mem_in_wire[29]), .IN1(inst_mem_in_wire[61]), .SEL(
        pc[2]), .F(n1856) );
  MUX U1886 ( .IN0(n1856), .IN1(n1855), .SEL(pc[3]), .F(n1857) );
  MUX U1887 ( .IN0(n1857), .IN1(n1854), .SEL(pc[4]), .F(n1858) );
  MUX U1888 ( .IN0(n1858), .IN1(n1851), .SEL(pc[5]), .F(n1859) );
  MUX U1889 ( .IN0(n1859), .IN1(n1844), .SEL(pc[6]), .F(n1860) );
  MUX U1890 ( .IN0(n1860), .IN1(n1829), .SEL(pc[7]), .F(opcode[29]) );
  MUX U1891 ( .IN0(inst_mem_in_wire[2014]), .IN1(inst_mem_in_wire[2046]), 
        .SEL(pc[2]), .F(n1861) );
  MUX U1892 ( .IN0(inst_mem_in_wire[1950]), .IN1(inst_mem_in_wire[1982]), 
        .SEL(pc[2]), .F(n1862) );
  MUX U1893 ( .IN0(n1862), .IN1(n1861), .SEL(pc[3]), .F(n1863) );
  MUX U1894 ( .IN0(inst_mem_in_wire[1886]), .IN1(inst_mem_in_wire[1918]), 
        .SEL(pc[2]), .F(n1864) );
  MUX U1895 ( .IN0(inst_mem_in_wire[1822]), .IN1(inst_mem_in_wire[1854]), 
        .SEL(pc[2]), .F(n1865) );
  MUX U1896 ( .IN0(n1865), .IN1(n1864), .SEL(pc[3]), .F(n1866) );
  MUX U1897 ( .IN0(n1866), .IN1(n1863), .SEL(pc[4]), .F(n1867) );
  MUX U1898 ( .IN0(inst_mem_in_wire[1758]), .IN1(inst_mem_in_wire[1790]), 
        .SEL(pc[2]), .F(n1868) );
  MUX U1899 ( .IN0(inst_mem_in_wire[1694]), .IN1(inst_mem_in_wire[1726]), 
        .SEL(pc[2]), .F(n1869) );
  MUX U1900 ( .IN0(n1869), .IN1(n1868), .SEL(pc[3]), .F(n1870) );
  MUX U1901 ( .IN0(inst_mem_in_wire[1630]), .IN1(inst_mem_in_wire[1662]), 
        .SEL(pc[2]), .F(n1871) );
  MUX U1902 ( .IN0(inst_mem_in_wire[1566]), .IN1(inst_mem_in_wire[1598]), 
        .SEL(pc[2]), .F(n1872) );
  MUX U1903 ( .IN0(n1872), .IN1(n1871), .SEL(pc[3]), .F(n1873) );
  MUX U1904 ( .IN0(n1873), .IN1(n1870), .SEL(pc[4]), .F(n1874) );
  MUX U1905 ( .IN0(n1874), .IN1(n1867), .SEL(pc[5]), .F(n1875) );
  MUX U1906 ( .IN0(inst_mem_in_wire[1502]), .IN1(inst_mem_in_wire[1534]), 
        .SEL(pc[2]), .F(n1876) );
  MUX U1907 ( .IN0(inst_mem_in_wire[1438]), .IN1(inst_mem_in_wire[1470]), 
        .SEL(pc[2]), .F(n1877) );
  MUX U1908 ( .IN0(n1877), .IN1(n1876), .SEL(pc[3]), .F(n1878) );
  MUX U1909 ( .IN0(inst_mem_in_wire[1374]), .IN1(inst_mem_in_wire[1406]), 
        .SEL(pc[2]), .F(n1879) );
  MUX U1910 ( .IN0(inst_mem_in_wire[1310]), .IN1(inst_mem_in_wire[1342]), 
        .SEL(pc[2]), .F(n1880) );
  MUX U1911 ( .IN0(n1880), .IN1(n1879), .SEL(pc[3]), .F(n1881) );
  MUX U1912 ( .IN0(n1881), .IN1(n1878), .SEL(pc[4]), .F(n1882) );
  MUX U1913 ( .IN0(inst_mem_in_wire[1246]), .IN1(inst_mem_in_wire[1278]), 
        .SEL(pc[2]), .F(n1883) );
  MUX U1914 ( .IN0(inst_mem_in_wire[1182]), .IN1(inst_mem_in_wire[1214]), 
        .SEL(pc[2]), .F(n1884) );
  MUX U1915 ( .IN0(n1884), .IN1(n1883), .SEL(pc[3]), .F(n1885) );
  MUX U1916 ( .IN0(inst_mem_in_wire[1118]), .IN1(inst_mem_in_wire[1150]), 
        .SEL(pc[2]), .F(n1886) );
  MUX U1917 ( .IN0(inst_mem_in_wire[1054]), .IN1(inst_mem_in_wire[1086]), 
        .SEL(pc[2]), .F(n1887) );
  MUX U1918 ( .IN0(n1887), .IN1(n1886), .SEL(pc[3]), .F(n1888) );
  MUX U1919 ( .IN0(n1888), .IN1(n1885), .SEL(pc[4]), .F(n1889) );
  MUX U1920 ( .IN0(n1889), .IN1(n1882), .SEL(pc[5]), .F(n1890) );
  MUX U1921 ( .IN0(n1890), .IN1(n1875), .SEL(pc[6]), .F(n1891) );
  MUX U1922 ( .IN0(inst_mem_in_wire[990]), .IN1(inst_mem_in_wire[1022]), .SEL(
        pc[2]), .F(n1892) );
  MUX U1923 ( .IN0(inst_mem_in_wire[926]), .IN1(inst_mem_in_wire[958]), .SEL(
        pc[2]), .F(n1893) );
  MUX U1924 ( .IN0(n1893), .IN1(n1892), .SEL(pc[3]), .F(n1894) );
  MUX U1925 ( .IN0(inst_mem_in_wire[862]), .IN1(inst_mem_in_wire[894]), .SEL(
        pc[2]), .F(n1895) );
  MUX U1926 ( .IN0(inst_mem_in_wire[798]), .IN1(inst_mem_in_wire[830]), .SEL(
        pc[2]), .F(n1896) );
  MUX U1927 ( .IN0(n1896), .IN1(n1895), .SEL(pc[3]), .F(n1897) );
  MUX U1928 ( .IN0(n1897), .IN1(n1894), .SEL(pc[4]), .F(n1898) );
  MUX U1929 ( .IN0(inst_mem_in_wire[734]), .IN1(inst_mem_in_wire[766]), .SEL(
        pc[2]), .F(n1899) );
  MUX U1930 ( .IN0(inst_mem_in_wire[670]), .IN1(inst_mem_in_wire[702]), .SEL(
        pc[2]), .F(n1900) );
  MUX U1931 ( .IN0(n1900), .IN1(n1899), .SEL(pc[3]), .F(n1901) );
  MUX U1932 ( .IN0(inst_mem_in_wire[606]), .IN1(inst_mem_in_wire[638]), .SEL(
        pc[2]), .F(n1902) );
  MUX U1933 ( .IN0(inst_mem_in_wire[542]), .IN1(inst_mem_in_wire[574]), .SEL(
        pc[2]), .F(n1903) );
  MUX U1934 ( .IN0(n1903), .IN1(n1902), .SEL(pc[3]), .F(n1904) );
  MUX U1935 ( .IN0(n1904), .IN1(n1901), .SEL(pc[4]), .F(n1905) );
  MUX U1936 ( .IN0(n1905), .IN1(n1898), .SEL(pc[5]), .F(n1906) );
  MUX U1937 ( .IN0(inst_mem_in_wire[478]), .IN1(inst_mem_in_wire[510]), .SEL(
        pc[2]), .F(n1907) );
  MUX U1938 ( .IN0(inst_mem_in_wire[414]), .IN1(inst_mem_in_wire[446]), .SEL(
        pc[2]), .F(n1908) );
  MUX U1939 ( .IN0(n1908), .IN1(n1907), .SEL(pc[3]), .F(n1909) );
  MUX U1940 ( .IN0(inst_mem_in_wire[350]), .IN1(inst_mem_in_wire[382]), .SEL(
        pc[2]), .F(n1910) );
  MUX U1941 ( .IN0(inst_mem_in_wire[286]), .IN1(inst_mem_in_wire[318]), .SEL(
        pc[2]), .F(n1911) );
  MUX U1942 ( .IN0(n1911), .IN1(n1910), .SEL(pc[3]), .F(n1912) );
  MUX U1943 ( .IN0(n1912), .IN1(n1909), .SEL(pc[4]), .F(n1913) );
  MUX U1944 ( .IN0(inst_mem_in_wire[222]), .IN1(inst_mem_in_wire[254]), .SEL(
        pc[2]), .F(n1914) );
  MUX U1945 ( .IN0(inst_mem_in_wire[158]), .IN1(inst_mem_in_wire[190]), .SEL(
        pc[2]), .F(n1915) );
  MUX U1946 ( .IN0(n1915), .IN1(n1914), .SEL(pc[3]), .F(n1916) );
  MUX U1947 ( .IN0(inst_mem_in_wire[94]), .IN1(inst_mem_in_wire[126]), .SEL(
        pc[2]), .F(n1917) );
  MUX U1948 ( .IN0(inst_mem_in_wire[30]), .IN1(inst_mem_in_wire[62]), .SEL(
        pc[2]), .F(n1918) );
  MUX U1949 ( .IN0(n1918), .IN1(n1917), .SEL(pc[3]), .F(n1919) );
  MUX U1950 ( .IN0(n1919), .IN1(n1916), .SEL(pc[4]), .F(n1920) );
  MUX U1951 ( .IN0(n1920), .IN1(n1913), .SEL(pc[5]), .F(n1921) );
  MUX U1952 ( .IN0(n1921), .IN1(n1906), .SEL(pc[6]), .F(n1922) );
  MUX U1953 ( .IN0(n1922), .IN1(n1891), .SEL(pc[7]), .F(opcode[30]) );
  MUX U1954 ( .IN0(inst_mem_in_wire[2015]), .IN1(inst_mem_in_wire[2047]), 
        .SEL(pc[2]), .F(n1923) );
  MUX U1955 ( .IN0(inst_mem_in_wire[1951]), .IN1(inst_mem_in_wire[1983]), 
        .SEL(pc[2]), .F(n1924) );
  MUX U1956 ( .IN0(n1924), .IN1(n1923), .SEL(pc[3]), .F(n1925) );
  MUX U1957 ( .IN0(inst_mem_in_wire[1887]), .IN1(inst_mem_in_wire[1919]), 
        .SEL(pc[2]), .F(n1926) );
  MUX U1958 ( .IN0(inst_mem_in_wire[1823]), .IN1(inst_mem_in_wire[1855]), 
        .SEL(pc[2]), .F(n1927) );
  MUX U1959 ( .IN0(n1927), .IN1(n1926), .SEL(pc[3]), .F(n1928) );
  MUX U1960 ( .IN0(n1928), .IN1(n1925), .SEL(pc[4]), .F(n1929) );
  MUX U1961 ( .IN0(inst_mem_in_wire[1759]), .IN1(inst_mem_in_wire[1791]), 
        .SEL(pc[2]), .F(n1930) );
  MUX U1962 ( .IN0(inst_mem_in_wire[1695]), .IN1(inst_mem_in_wire[1727]), 
        .SEL(pc[2]), .F(n1931) );
  MUX U1963 ( .IN0(n1931), .IN1(n1930), .SEL(pc[3]), .F(n1932) );
  MUX U1964 ( .IN0(inst_mem_in_wire[1631]), .IN1(inst_mem_in_wire[1663]), 
        .SEL(pc[2]), .F(n1933) );
  MUX U1965 ( .IN0(inst_mem_in_wire[1567]), .IN1(inst_mem_in_wire[1599]), 
        .SEL(pc[2]), .F(n1934) );
  MUX U1966 ( .IN0(n1934), .IN1(n1933), .SEL(pc[3]), .F(n1935) );
  MUX U1967 ( .IN0(n1935), .IN1(n1932), .SEL(pc[4]), .F(n1936) );
  MUX U1968 ( .IN0(n1936), .IN1(n1929), .SEL(pc[5]), .F(n1937) );
  MUX U1969 ( .IN0(inst_mem_in_wire[1503]), .IN1(inst_mem_in_wire[1535]), 
        .SEL(pc[2]), .F(n1938) );
  MUX U1970 ( .IN0(inst_mem_in_wire[1439]), .IN1(inst_mem_in_wire[1471]), 
        .SEL(pc[2]), .F(n1939) );
  MUX U1971 ( .IN0(n1939), .IN1(n1938), .SEL(pc[3]), .F(n1940) );
  MUX U1972 ( .IN0(inst_mem_in_wire[1375]), .IN1(inst_mem_in_wire[1407]), 
        .SEL(pc[2]), .F(n1941) );
  MUX U1973 ( .IN0(inst_mem_in_wire[1311]), .IN1(inst_mem_in_wire[1343]), 
        .SEL(pc[2]), .F(n1942) );
  MUX U1974 ( .IN0(n1942), .IN1(n1941), .SEL(pc[3]), .F(n1943) );
  MUX U1975 ( .IN0(n1943), .IN1(n1940), .SEL(pc[4]), .F(n1944) );
  MUX U1976 ( .IN0(inst_mem_in_wire[1247]), .IN1(inst_mem_in_wire[1279]), 
        .SEL(pc[2]), .F(n1945) );
  MUX U1977 ( .IN0(inst_mem_in_wire[1183]), .IN1(inst_mem_in_wire[1215]), 
        .SEL(pc[2]), .F(n1946) );
  MUX U1978 ( .IN0(n1946), .IN1(n1945), .SEL(pc[3]), .F(n1947) );
  MUX U1979 ( .IN0(inst_mem_in_wire[1119]), .IN1(inst_mem_in_wire[1151]), 
        .SEL(pc[2]), .F(n1948) );
  MUX U1980 ( .IN0(inst_mem_in_wire[1055]), .IN1(inst_mem_in_wire[1087]), 
        .SEL(pc[2]), .F(n1949) );
  MUX U1981 ( .IN0(n1949), .IN1(n1948), .SEL(pc[3]), .F(n1950) );
  MUX U1982 ( .IN0(n1950), .IN1(n1947), .SEL(pc[4]), .F(n1951) );
  MUX U1983 ( .IN0(n1951), .IN1(n1944), .SEL(pc[5]), .F(n1952) );
  MUX U1984 ( .IN0(n1952), .IN1(n1937), .SEL(pc[6]), .F(n1953) );
  MUX U1985 ( .IN0(inst_mem_in_wire[991]), .IN1(inst_mem_in_wire[1023]), .SEL(
        pc[2]), .F(n1954) );
  MUX U1986 ( .IN0(inst_mem_in_wire[927]), .IN1(inst_mem_in_wire[959]), .SEL(
        pc[2]), .F(n1955) );
  MUX U1987 ( .IN0(n1955), .IN1(n1954), .SEL(pc[3]), .F(n1956) );
  MUX U1988 ( .IN0(inst_mem_in_wire[863]), .IN1(inst_mem_in_wire[895]), .SEL(
        pc[2]), .F(n1957) );
  MUX U1989 ( .IN0(inst_mem_in_wire[799]), .IN1(inst_mem_in_wire[831]), .SEL(
        pc[2]), .F(n1958) );
  MUX U1990 ( .IN0(n1958), .IN1(n1957), .SEL(pc[3]), .F(n1959) );
  MUX U1991 ( .IN0(n1959), .IN1(n1956), .SEL(pc[4]), .F(n1960) );
  MUX U1992 ( .IN0(inst_mem_in_wire[735]), .IN1(inst_mem_in_wire[767]), .SEL(
        pc[2]), .F(n1961) );
  MUX U1993 ( .IN0(inst_mem_in_wire[671]), .IN1(inst_mem_in_wire[703]), .SEL(
        pc[2]), .F(n1962) );
  MUX U1994 ( .IN0(n1962), .IN1(n1961), .SEL(pc[3]), .F(n1963) );
  MUX U1995 ( .IN0(inst_mem_in_wire[607]), .IN1(inst_mem_in_wire[639]), .SEL(
        pc[2]), .F(n1964) );
  MUX U1996 ( .IN0(inst_mem_in_wire[543]), .IN1(inst_mem_in_wire[575]), .SEL(
        pc[2]), .F(n1965) );
  MUX U1997 ( .IN0(n1965), .IN1(n1964), .SEL(pc[3]), .F(n1966) );
  MUX U1998 ( .IN0(n1966), .IN1(n1963), .SEL(pc[4]), .F(n1967) );
  MUX U1999 ( .IN0(n1967), .IN1(n1960), .SEL(pc[5]), .F(n1968) );
  MUX U2000 ( .IN0(inst_mem_in_wire[479]), .IN1(inst_mem_in_wire[511]), .SEL(
        pc[2]), .F(n1969) );
  MUX U2001 ( .IN0(inst_mem_in_wire[415]), .IN1(inst_mem_in_wire[447]), .SEL(
        pc[2]), .F(n1970) );
  MUX U2002 ( .IN0(n1970), .IN1(n1969), .SEL(pc[3]), .F(n1971) );
  MUX U2003 ( .IN0(inst_mem_in_wire[351]), .IN1(inst_mem_in_wire[383]), .SEL(
        pc[2]), .F(n1972) );
  MUX U2004 ( .IN0(inst_mem_in_wire[287]), .IN1(inst_mem_in_wire[319]), .SEL(
        pc[2]), .F(n1973) );
  MUX U2005 ( .IN0(n1973), .IN1(n1972), .SEL(pc[3]), .F(n1974) );
  MUX U2006 ( .IN0(n1974), .IN1(n1971), .SEL(pc[4]), .F(n1975) );
  MUX U2007 ( .IN0(inst_mem_in_wire[223]), .IN1(inst_mem_in_wire[255]), .SEL(
        pc[2]), .F(n1976) );
  MUX U2008 ( .IN0(inst_mem_in_wire[159]), .IN1(inst_mem_in_wire[191]), .SEL(
        pc[2]), .F(n1977) );
  MUX U2009 ( .IN0(n1977), .IN1(n1976), .SEL(pc[3]), .F(n1978) );
  MUX U2010 ( .IN0(inst_mem_in_wire[95]), .IN1(inst_mem_in_wire[127]), .SEL(
        pc[2]), .F(n1979) );
  MUX U2011 ( .IN0(inst_mem_in_wire[31]), .IN1(inst_mem_in_wire[63]), .SEL(
        pc[2]), .F(n1980) );
  MUX U2012 ( .IN0(n1980), .IN1(n1979), .SEL(pc[3]), .F(n1981) );
  MUX U2013 ( .IN0(n1981), .IN1(n1978), .SEL(pc[4]), .F(n1982) );
  MUX U2014 ( .IN0(n1982), .IN1(n1975), .SEL(pc[5]), .F(n1983) );
  MUX U2015 ( .IN0(n1983), .IN1(n1968), .SEL(pc[6]), .F(n1984) );
  MUX U2016 ( .IN0(n1984), .IN1(n1953), .SEL(pc[7]), .F(opcode[31]) );
endmodule

