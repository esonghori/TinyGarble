
module Reg_Bank ( clk, rst, rs_index, rt_index, rd_index, reg_source_out, 
        reg_target_out, reg_dest_new );
  input [4:0] rs_index;
  input [4:0] rt_index;
  input [4:0] rd_index;
  output [31:0] reg_source_out;
  output [31:0] reg_target_out;
  input [31:0] reg_dest_new;
  input clk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, \registers[31][31] ,
         \registers[31][30] , \registers[31][29] , \registers[31][28] ,
         \registers[31][27] , \registers[31][26] , \registers[31][25] ,
         \registers[31][24] , \registers[31][23] , \registers[31][22] ,
         \registers[31][21] , \registers[31][20] , \registers[31][19] ,
         \registers[31][18] , \registers[31][17] , \registers[31][16] ,
         \registers[31][15] , \registers[31][14] , \registers[31][13] ,
         \registers[31][12] , \registers[31][11] , \registers[31][10] ,
         \registers[31][9] , \registers[31][8] , \registers[31][7] ,
         \registers[31][6] , \registers[31][5] , \registers[31][4] ,
         \registers[31][3] , \registers[31][2] , \registers[31][1] ,
         \registers[31][0] , \registers[30][31] , \registers[30][30] ,
         \registers[30][29] , \registers[30][28] , \registers[30][27] ,
         \registers[30][26] , \registers[30][25] , \registers[30][24] ,
         \registers[30][23] , \registers[30][22] , \registers[30][21] ,
         \registers[30][20] , \registers[30][19] , \registers[30][18] ,
         \registers[30][17] , \registers[30][16] , \registers[30][15] ,
         \registers[30][14] , \registers[30][13] , \registers[30][12] ,
         \registers[30][11] , \registers[30][10] , \registers[30][9] ,
         \registers[30][8] , \registers[30][7] , \registers[30][6] ,
         \registers[30][5] , \registers[30][4] , \registers[30][3] ,
         \registers[30][2] , \registers[30][1] , \registers[30][0] ,
         \registers[29][31] , \registers[29][30] , \registers[29][29] ,
         \registers[29][28] , \registers[29][27] , \registers[29][26] ,
         \registers[29][25] , \registers[29][24] , \registers[29][23] ,
         \registers[29][22] , \registers[29][21] , \registers[29][20] ,
         \registers[29][19] , \registers[29][18] , \registers[29][17] ,
         \registers[29][16] , \registers[29][15] , \registers[29][14] ,
         \registers[29][13] , \registers[29][12] , \registers[29][11] ,
         \registers[29][10] , \registers[29][9] , \registers[29][8] ,
         \registers[29][7] , \registers[29][6] , \registers[29][5] ,
         \registers[29][4] , \registers[29][3] , \registers[29][2] ,
         \registers[29][1] , \registers[29][0] , \registers[28][31] ,
         \registers[28][30] , \registers[28][29] , \registers[28][28] ,
         \registers[28][27] , \registers[28][26] , \registers[28][25] ,
         \registers[28][24] , \registers[28][23] , \registers[28][22] ,
         \registers[28][21] , \registers[28][20] , \registers[28][19] ,
         \registers[28][18] , \registers[28][17] , \registers[28][16] ,
         \registers[28][15] , \registers[28][14] , \registers[28][13] ,
         \registers[28][12] , \registers[28][11] , \registers[28][10] ,
         \registers[28][9] , \registers[28][8] , \registers[28][7] ,
         \registers[28][6] , \registers[28][5] , \registers[28][4] ,
         \registers[28][3] , \registers[28][2] , \registers[28][1] ,
         \registers[28][0] , \registers[27][31] , \registers[27][30] ,
         \registers[27][29] , \registers[27][28] , \registers[27][27] ,
         \registers[27][26] , \registers[27][25] , \registers[27][24] ,
         \registers[27][23] , \registers[27][22] , \registers[27][21] ,
         \registers[27][20] , \registers[27][19] , \registers[27][18] ,
         \registers[27][17] , \registers[27][16] , \registers[27][15] ,
         \registers[27][14] , \registers[27][13] , \registers[27][12] ,
         \registers[27][11] , \registers[27][10] , \registers[27][9] ,
         \registers[27][8] , \registers[27][7] , \registers[27][6] ,
         \registers[27][5] , \registers[27][4] , \registers[27][3] ,
         \registers[27][2] , \registers[27][1] , \registers[27][0] ,
         \registers[26][31] , \registers[26][30] , \registers[26][29] ,
         \registers[26][28] , \registers[26][27] , \registers[26][26] ,
         \registers[26][25] , \registers[26][24] , \registers[26][23] ,
         \registers[26][22] , \registers[26][21] , \registers[26][20] ,
         \registers[26][19] , \registers[26][18] , \registers[26][17] ,
         \registers[26][16] , \registers[26][15] , \registers[26][14] ,
         \registers[26][13] , \registers[26][12] , \registers[26][11] ,
         \registers[26][10] , \registers[26][9] , \registers[26][8] ,
         \registers[26][7] , \registers[26][6] , \registers[26][5] ,
         \registers[26][4] , \registers[26][3] , \registers[26][2] ,
         \registers[26][1] , \registers[26][0] , \registers[25][31] ,
         \registers[25][30] , \registers[25][29] , \registers[25][28] ,
         \registers[25][27] , \registers[25][26] , \registers[25][25] ,
         \registers[25][24] , \registers[25][23] , \registers[25][22] ,
         \registers[25][21] , \registers[25][20] , \registers[25][19] ,
         \registers[25][18] , \registers[25][17] , \registers[25][16] ,
         \registers[25][15] , \registers[25][14] , \registers[25][13] ,
         \registers[25][12] , \registers[25][11] , \registers[25][10] ,
         \registers[25][9] , \registers[25][8] , \registers[25][7] ,
         \registers[25][6] , \registers[25][5] , \registers[25][4] ,
         \registers[25][3] , \registers[25][2] , \registers[25][1] ,
         \registers[25][0] , \registers[24][31] , \registers[24][30] ,
         \registers[24][29] , \registers[24][28] , \registers[24][27] ,
         \registers[24][26] , \registers[24][25] , \registers[24][24] ,
         \registers[24][23] , \registers[24][22] , \registers[24][21] ,
         \registers[24][20] , \registers[24][19] , \registers[24][18] ,
         \registers[24][17] , \registers[24][16] , \registers[24][15] ,
         \registers[24][14] , \registers[24][13] , \registers[24][12] ,
         \registers[24][11] , \registers[24][10] , \registers[24][9] ,
         \registers[24][8] , \registers[24][7] , \registers[24][6] ,
         \registers[24][5] , \registers[24][4] , \registers[24][3] ,
         \registers[24][2] , \registers[24][1] , \registers[24][0] ,
         \registers[23][31] , \registers[23][30] , \registers[23][29] ,
         \registers[23][28] , \registers[23][27] , \registers[23][26] ,
         \registers[23][25] , \registers[23][24] , \registers[23][23] ,
         \registers[23][22] , \registers[23][21] , \registers[23][20] ,
         \registers[23][19] , \registers[23][18] , \registers[23][17] ,
         \registers[23][16] , \registers[23][15] , \registers[23][14] ,
         \registers[23][13] , \registers[23][12] , \registers[23][11] ,
         \registers[23][10] , \registers[23][9] , \registers[23][8] ,
         \registers[23][7] , \registers[23][6] , \registers[23][5] ,
         \registers[23][4] , \registers[23][3] , \registers[23][2] ,
         \registers[23][1] , \registers[23][0] , \registers[22][31] ,
         \registers[22][30] , \registers[22][29] , \registers[22][28] ,
         \registers[22][27] , \registers[22][26] , \registers[22][25] ,
         \registers[22][24] , \registers[22][23] , \registers[22][22] ,
         \registers[22][21] , \registers[22][20] , \registers[22][19] ,
         \registers[22][18] , \registers[22][17] , \registers[22][16] ,
         \registers[22][15] , \registers[22][14] , \registers[22][13] ,
         \registers[22][12] , \registers[22][11] , \registers[22][10] ,
         \registers[22][9] , \registers[22][8] , \registers[22][7] ,
         \registers[22][6] , \registers[22][5] , \registers[22][4] ,
         \registers[22][3] , \registers[22][2] , \registers[22][1] ,
         \registers[22][0] , \registers[21][31] , \registers[21][30] ,
         \registers[21][29] , \registers[21][28] , \registers[21][27] ,
         \registers[21][26] , \registers[21][25] , \registers[21][24] ,
         \registers[21][23] , \registers[21][22] , \registers[21][21] ,
         \registers[21][20] , \registers[21][19] , \registers[21][18] ,
         \registers[21][17] , \registers[21][16] , \registers[21][15] ,
         \registers[21][14] , \registers[21][13] , \registers[21][12] ,
         \registers[21][11] , \registers[21][10] , \registers[21][9] ,
         \registers[21][8] , \registers[21][7] , \registers[21][6] ,
         \registers[21][5] , \registers[21][4] , \registers[21][3] ,
         \registers[21][2] , \registers[21][1] , \registers[21][0] ,
         \registers[20][31] , \registers[20][30] , \registers[20][29] ,
         \registers[20][28] , \registers[20][27] , \registers[20][26] ,
         \registers[20][25] , \registers[20][24] , \registers[20][23] ,
         \registers[20][22] , \registers[20][21] , \registers[20][20] ,
         \registers[20][19] , \registers[20][18] , \registers[20][17] ,
         \registers[20][16] , \registers[20][15] , \registers[20][14] ,
         \registers[20][13] , \registers[20][12] , \registers[20][11] ,
         \registers[20][10] , \registers[20][9] , \registers[20][8] ,
         \registers[20][7] , \registers[20][6] , \registers[20][5] ,
         \registers[20][4] , \registers[20][3] , \registers[20][2] ,
         \registers[20][1] , \registers[20][0] , \registers[19][31] ,
         \registers[19][30] , \registers[19][29] , \registers[19][28] ,
         \registers[19][27] , \registers[19][26] , \registers[19][25] ,
         \registers[19][24] , \registers[19][23] , \registers[19][22] ,
         \registers[19][21] , \registers[19][20] , \registers[19][19] ,
         \registers[19][18] , \registers[19][17] , \registers[19][16] ,
         \registers[19][15] , \registers[19][14] , \registers[19][13] ,
         \registers[19][12] , \registers[19][11] , \registers[19][10] ,
         \registers[19][9] , \registers[19][8] , \registers[19][7] ,
         \registers[19][6] , \registers[19][5] , \registers[19][4] ,
         \registers[19][3] , \registers[19][2] , \registers[19][1] ,
         \registers[19][0] , \registers[18][31] , \registers[18][30] ,
         \registers[18][29] , \registers[18][28] , \registers[18][27] ,
         \registers[18][26] , \registers[18][25] , \registers[18][24] ,
         \registers[18][23] , \registers[18][22] , \registers[18][21] ,
         \registers[18][20] , \registers[18][19] , \registers[18][18] ,
         \registers[18][17] , \registers[18][16] , \registers[18][15] ,
         \registers[18][14] , \registers[18][13] , \registers[18][12] ,
         \registers[18][11] , \registers[18][10] , \registers[18][9] ,
         \registers[18][8] , \registers[18][7] , \registers[18][6] ,
         \registers[18][5] , \registers[18][4] , \registers[18][3] ,
         \registers[18][2] , \registers[18][1] , \registers[18][0] ,
         \registers[17][31] , \registers[17][30] , \registers[17][29] ,
         \registers[17][28] , \registers[17][27] , \registers[17][26] ,
         \registers[17][25] , \registers[17][24] , \registers[17][23] ,
         \registers[17][22] , \registers[17][21] , \registers[17][20] ,
         \registers[17][19] , \registers[17][18] , \registers[17][17] ,
         \registers[17][16] , \registers[17][15] , \registers[17][14] ,
         \registers[17][13] , \registers[17][12] , \registers[17][11] ,
         \registers[17][10] , \registers[17][9] , \registers[17][8] ,
         \registers[17][7] , \registers[17][6] , \registers[17][5] ,
         \registers[17][4] , \registers[17][3] , \registers[17][2] ,
         \registers[17][1] , \registers[17][0] , \registers[16][31] ,
         \registers[16][30] , \registers[16][29] , \registers[16][28] ,
         \registers[16][27] , \registers[16][26] , \registers[16][25] ,
         \registers[16][24] , \registers[16][23] , \registers[16][22] ,
         \registers[16][21] , \registers[16][20] , \registers[16][19] ,
         \registers[16][18] , \registers[16][17] , \registers[16][16] ,
         \registers[16][15] , \registers[16][14] , \registers[16][13] ,
         \registers[16][12] , \registers[16][11] , \registers[16][10] ,
         \registers[16][9] , \registers[16][8] , \registers[16][7] ,
         \registers[16][6] , \registers[16][5] , \registers[16][4] ,
         \registers[16][3] , \registers[16][2] , \registers[16][1] ,
         \registers[16][0] , \registers[15][31] , \registers[15][30] ,
         \registers[15][29] , \registers[15][28] , \registers[15][27] ,
         \registers[15][26] , \registers[15][25] , \registers[15][24] ,
         \registers[15][23] , \registers[15][22] , \registers[15][21] ,
         \registers[15][20] , \registers[15][19] , \registers[15][18] ,
         \registers[15][17] , \registers[15][16] , \registers[15][15] ,
         \registers[15][14] , \registers[15][13] , \registers[15][12] ,
         \registers[15][11] , \registers[15][10] , \registers[15][9] ,
         \registers[15][8] , \registers[15][7] , \registers[15][6] ,
         \registers[15][5] , \registers[15][4] , \registers[15][3] ,
         \registers[15][2] , \registers[15][1] , \registers[15][0] ,
         \registers[14][31] , \registers[14][30] , \registers[14][29] ,
         \registers[14][28] , \registers[14][27] , \registers[14][26] ,
         \registers[14][25] , \registers[14][24] , \registers[14][23] ,
         \registers[14][22] , \registers[14][21] , \registers[14][20] ,
         \registers[14][19] , \registers[14][18] , \registers[14][17] ,
         \registers[14][16] , \registers[14][15] , \registers[14][14] ,
         \registers[14][13] , \registers[14][12] , \registers[14][11] ,
         \registers[14][10] , \registers[14][9] , \registers[14][8] ,
         \registers[14][7] , \registers[14][6] , \registers[14][5] ,
         \registers[14][4] , \registers[14][3] , \registers[14][2] ,
         \registers[14][1] , \registers[14][0] , \registers[13][31] ,
         \registers[13][30] , \registers[13][29] , \registers[13][28] ,
         \registers[13][27] , \registers[13][26] , \registers[13][25] ,
         \registers[13][24] , \registers[13][23] , \registers[13][22] ,
         \registers[13][21] , \registers[13][20] , \registers[13][19] ,
         \registers[13][18] , \registers[13][17] , \registers[13][16] ,
         \registers[13][15] , \registers[13][14] , \registers[13][13] ,
         \registers[13][12] , \registers[13][11] , \registers[13][10] ,
         \registers[13][9] , \registers[13][8] , \registers[13][7] ,
         \registers[13][6] , \registers[13][5] , \registers[13][4] ,
         \registers[13][3] , \registers[13][2] , \registers[13][1] ,
         \registers[13][0] , \registers[12][31] , \registers[12][30] ,
         \registers[12][29] , \registers[12][28] , \registers[12][27] ,
         \registers[12][26] , \registers[12][25] , \registers[12][24] ,
         \registers[12][23] , \registers[12][22] , \registers[12][21] ,
         \registers[12][20] , \registers[12][19] , \registers[12][18] ,
         \registers[12][17] , \registers[12][16] , \registers[12][15] ,
         \registers[12][14] , \registers[12][13] , \registers[12][12] ,
         \registers[12][11] , \registers[12][10] , \registers[12][9] ,
         \registers[12][8] , \registers[12][7] , \registers[12][6] ,
         \registers[12][5] , \registers[12][4] , \registers[12][3] ,
         \registers[12][2] , \registers[12][1] , \registers[12][0] ,
         \registers[11][31] , \registers[11][30] , \registers[11][29] ,
         \registers[11][28] , \registers[11][27] , \registers[11][26] ,
         \registers[11][25] , \registers[11][24] , \registers[11][23] ,
         \registers[11][22] , \registers[11][21] , \registers[11][20] ,
         \registers[11][19] , \registers[11][18] , \registers[11][17] ,
         \registers[11][16] , \registers[11][15] , \registers[11][14] ,
         \registers[11][13] , \registers[11][12] , \registers[11][11] ,
         \registers[11][10] , \registers[11][9] , \registers[11][8] ,
         \registers[11][7] , \registers[11][6] , \registers[11][5] ,
         \registers[11][4] , \registers[11][3] , \registers[11][2] ,
         \registers[11][1] , \registers[11][0] , \registers[10][31] ,
         \registers[10][30] , \registers[10][29] , \registers[10][28] ,
         \registers[10][27] , \registers[10][26] , \registers[10][25] ,
         \registers[10][24] , \registers[10][23] , \registers[10][22] ,
         \registers[10][21] , \registers[10][20] , \registers[10][19] ,
         \registers[10][18] , \registers[10][17] , \registers[10][16] ,
         \registers[10][15] , \registers[10][14] , \registers[10][13] ,
         \registers[10][12] , \registers[10][11] , \registers[10][10] ,
         \registers[10][9] , \registers[10][8] , \registers[10][7] ,
         \registers[10][6] , \registers[10][5] , \registers[10][4] ,
         \registers[10][3] , \registers[10][2] , \registers[10][1] ,
         \registers[10][0] , \registers[9][31] , \registers[9][30] ,
         \registers[9][29] , \registers[9][28] , \registers[9][27] ,
         \registers[9][26] , \registers[9][25] , \registers[9][24] ,
         \registers[9][23] , \registers[9][22] , \registers[9][21] ,
         \registers[9][20] , \registers[9][19] , \registers[9][18] ,
         \registers[9][17] , \registers[9][16] , \registers[9][15] ,
         \registers[9][14] , \registers[9][13] , \registers[9][12] ,
         \registers[9][11] , \registers[9][10] , \registers[9][9] ,
         \registers[9][8] , \registers[9][7] , \registers[9][6] ,
         \registers[9][5] , \registers[9][4] , \registers[9][3] ,
         \registers[9][2] , \registers[9][1] , \registers[9][0] ,
         \registers[8][31] , \registers[8][30] , \registers[8][29] ,
         \registers[8][28] , \registers[8][27] , \registers[8][26] ,
         \registers[8][25] , \registers[8][24] , \registers[8][23] ,
         \registers[8][22] , \registers[8][21] , \registers[8][20] ,
         \registers[8][19] , \registers[8][18] , \registers[8][17] ,
         \registers[8][16] , \registers[8][15] , \registers[8][14] ,
         \registers[8][13] , \registers[8][12] , \registers[8][11] ,
         \registers[8][10] , \registers[8][9] , \registers[8][8] ,
         \registers[8][7] , \registers[8][6] , \registers[8][5] ,
         \registers[8][4] , \registers[8][3] , \registers[8][2] ,
         \registers[8][1] , \registers[8][0] , \registers[7][31] ,
         \registers[7][30] , \registers[7][29] , \registers[7][28] ,
         \registers[7][27] , \registers[7][26] , \registers[7][25] ,
         \registers[7][24] , \registers[7][23] , \registers[7][22] ,
         \registers[7][21] , \registers[7][20] , \registers[7][19] ,
         \registers[7][18] , \registers[7][17] , \registers[7][16] ,
         \registers[7][15] , \registers[7][14] , \registers[7][13] ,
         \registers[7][12] , \registers[7][11] , \registers[7][10] ,
         \registers[7][9] , \registers[7][8] , \registers[7][7] ,
         \registers[7][6] , \registers[7][5] , \registers[7][4] ,
         \registers[7][3] , \registers[7][2] , \registers[7][1] ,
         \registers[7][0] , \registers[6][31] , \registers[6][30] ,
         \registers[6][29] , \registers[6][28] , \registers[6][27] ,
         \registers[6][26] , \registers[6][25] , \registers[6][24] ,
         \registers[6][23] , \registers[6][22] , \registers[6][21] ,
         \registers[6][20] , \registers[6][19] , \registers[6][18] ,
         \registers[6][17] , \registers[6][16] , \registers[6][15] ,
         \registers[6][14] , \registers[6][13] , \registers[6][12] ,
         \registers[6][11] , \registers[6][10] , \registers[6][9] ,
         \registers[6][8] , \registers[6][7] , \registers[6][6] ,
         \registers[6][5] , \registers[6][4] , \registers[6][3] ,
         \registers[6][2] , \registers[6][1] , \registers[6][0] ,
         \registers[5][31] , \registers[5][30] , \registers[5][29] ,
         \registers[5][28] , \registers[5][27] , \registers[5][26] ,
         \registers[5][25] , \registers[5][24] , \registers[5][23] ,
         \registers[5][22] , \registers[5][21] , \registers[5][20] ,
         \registers[5][19] , \registers[5][18] , \registers[5][17] ,
         \registers[5][16] , \registers[5][15] , \registers[5][14] ,
         \registers[5][13] , \registers[5][12] , \registers[5][11] ,
         \registers[5][10] , \registers[5][9] , \registers[5][8] ,
         \registers[5][7] , \registers[5][6] , \registers[5][5] ,
         \registers[5][4] , \registers[5][3] , \registers[5][2] ,
         \registers[5][1] , \registers[5][0] , \registers[4][31] ,
         \registers[4][30] , \registers[4][29] , \registers[4][28] ,
         \registers[4][27] , \registers[4][26] , \registers[4][25] ,
         \registers[4][24] , \registers[4][23] , \registers[4][22] ,
         \registers[4][21] , \registers[4][20] , \registers[4][19] ,
         \registers[4][18] , \registers[4][17] , \registers[4][16] ,
         \registers[4][15] , \registers[4][14] , \registers[4][13] ,
         \registers[4][12] , \registers[4][11] , \registers[4][10] ,
         \registers[4][9] , \registers[4][8] , \registers[4][7] ,
         \registers[4][6] , \registers[4][5] , \registers[4][4] ,
         \registers[4][3] , \registers[4][2] , \registers[4][1] ,
         \registers[4][0] , \registers[3][31] , \registers[3][30] ,
         \registers[3][29] , \registers[3][28] , \registers[3][27] ,
         \registers[3][26] , \registers[3][25] , \registers[3][24] ,
         \registers[3][23] , \registers[3][22] , \registers[3][21] ,
         \registers[3][20] , \registers[3][19] , \registers[3][18] ,
         \registers[3][17] , \registers[3][16] , \registers[3][15] ,
         \registers[3][14] , \registers[3][13] , \registers[3][12] ,
         \registers[3][11] , \registers[3][10] , \registers[3][9] ,
         \registers[3][8] , \registers[3][7] , \registers[3][6] ,
         \registers[3][5] , \registers[3][4] , \registers[3][3] ,
         \registers[3][2] , \registers[3][1] , \registers[3][0] ,
         \registers[2][31] , \registers[2][30] , \registers[2][29] ,
         \registers[2][28] , \registers[2][27] , \registers[2][26] ,
         \registers[2][25] , \registers[2][24] , \registers[2][23] ,
         \registers[2][22] , \registers[2][21] , \registers[2][20] ,
         \registers[2][19] , \registers[2][18] , \registers[2][17] ,
         \registers[2][16] , \registers[2][15] , \registers[2][14] ,
         \registers[2][13] , \registers[2][12] , \registers[2][11] ,
         \registers[2][10] , \registers[2][9] , \registers[2][8] ,
         \registers[2][7] , \registers[2][6] , \registers[2][5] ,
         \registers[2][4] , \registers[2][3] , \registers[2][2] ,
         \registers[2][1] , \registers[2][0] , \registers[1][31] ,
         \registers[1][30] , \registers[1][29] , \registers[1][28] ,
         \registers[1][27] , \registers[1][26] , \registers[1][25] ,
         \registers[1][24] , \registers[1][23] , \registers[1][22] ,
         \registers[1][21] , \registers[1][20] , \registers[1][19] ,
         \registers[1][18] , \registers[1][17] , \registers[1][16] ,
         \registers[1][15] , \registers[1][14] , \registers[1][13] ,
         \registers[1][12] , \registers[1][11] , \registers[1][10] ,
         \registers[1][9] , \registers[1][8] , \registers[1][7] ,
         \registers[1][6] , \registers[1][5] , \registers[1][4] ,
         \registers[1][3] , \registers[1][2] , \registers[1][1] ,
         \registers[1][0] , n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017;
  assign N9 = rs_index[0];
  assign N10 = rs_index[1];
  assign N11 = rs_index[2];
  assign N12 = rs_index[3];
  assign N13 = rs_index[4];
  assign N14 = rt_index[0];
  assign N15 = rt_index[1];
  assign N16 = rt_index[2];
  assign N17 = rt_index[3];
  assign N18 = rt_index[4];

  DFF \registers_reg[31][31]  ( .D(n4017), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][31] ) );
  DFF \registers_reg[31][30]  ( .D(n4016), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][30] ) );
  DFF \registers_reg[31][29]  ( .D(n4015), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][29] ) );
  DFF \registers_reg[31][28]  ( .D(n4014), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][28] ) );
  DFF \registers_reg[31][27]  ( .D(n4013), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][27] ) );
  DFF \registers_reg[31][26]  ( .D(n4012), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][26] ) );
  DFF \registers_reg[31][25]  ( .D(n4011), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][25] ) );
  DFF \registers_reg[31][24]  ( .D(n4010), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][24] ) );
  DFF \registers_reg[31][23]  ( .D(n4009), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][23] ) );
  DFF \registers_reg[31][22]  ( .D(n4008), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][22] ) );
  DFF \registers_reg[31][21]  ( .D(n4007), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][21] ) );
  DFF \registers_reg[31][20]  ( .D(n4006), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][20] ) );
  DFF \registers_reg[31][19]  ( .D(n4005), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][19] ) );
  DFF \registers_reg[31][18]  ( .D(n4004), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][18] ) );
  DFF \registers_reg[31][17]  ( .D(n4003), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][17] ) );
  DFF \registers_reg[31][16]  ( .D(n4002), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][16] ) );
  DFF \registers_reg[31][15]  ( .D(n4001), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][15] ) );
  DFF \registers_reg[31][14]  ( .D(n4000), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][14] ) );
  DFF \registers_reg[31][13]  ( .D(n3999), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][13] ) );
  DFF \registers_reg[31][12]  ( .D(n3998), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][12] ) );
  DFF \registers_reg[31][11]  ( .D(n3997), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][11] ) );
  DFF \registers_reg[31][10]  ( .D(n3996), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][10] ) );
  DFF \registers_reg[31][9]  ( .D(n3995), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][9] ) );
  DFF \registers_reg[31][8]  ( .D(n3994), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][8] ) );
  DFF \registers_reg[31][7]  ( .D(n3993), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][7] ) );
  DFF \registers_reg[31][6]  ( .D(n3992), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][6] ) );
  DFF \registers_reg[31][5]  ( .D(n3991), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][5] ) );
  DFF \registers_reg[31][4]  ( .D(n3990), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][4] ) );
  DFF \registers_reg[31][3]  ( .D(n3989), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][3] ) );
  DFF \registers_reg[31][2]  ( .D(n3988), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][2] ) );
  DFF \registers_reg[31][1]  ( .D(n3987), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][1] ) );
  DFF \registers_reg[31][0]  ( .D(n3986), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[31][0] ) );
  DFF \registers_reg[30][31]  ( .D(n3985), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][31] ) );
  DFF \registers_reg[30][30]  ( .D(n3984), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][30] ) );
  DFF \registers_reg[30][29]  ( .D(n3983), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][29] ) );
  DFF \registers_reg[30][28]  ( .D(n3982), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][28] ) );
  DFF \registers_reg[30][27]  ( .D(n3981), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][27] ) );
  DFF \registers_reg[30][26]  ( .D(n3980), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][26] ) );
  DFF \registers_reg[30][25]  ( .D(n3979), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][25] ) );
  DFF \registers_reg[30][24]  ( .D(n3978), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][24] ) );
  DFF \registers_reg[30][23]  ( .D(n3977), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][23] ) );
  DFF \registers_reg[30][22]  ( .D(n3976), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][22] ) );
  DFF \registers_reg[30][21]  ( .D(n3975), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][21] ) );
  DFF \registers_reg[30][20]  ( .D(n3974), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][20] ) );
  DFF \registers_reg[30][19]  ( .D(n3973), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][19] ) );
  DFF \registers_reg[30][18]  ( .D(n3972), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][18] ) );
  DFF \registers_reg[30][17]  ( .D(n3971), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][17] ) );
  DFF \registers_reg[30][16]  ( .D(n3970), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][16] ) );
  DFF \registers_reg[30][15]  ( .D(n3969), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][15] ) );
  DFF \registers_reg[30][14]  ( .D(n3968), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][14] ) );
  DFF \registers_reg[30][13]  ( .D(n3967), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][13] ) );
  DFF \registers_reg[30][12]  ( .D(n3966), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][12] ) );
  DFF \registers_reg[30][11]  ( .D(n3965), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][11] ) );
  DFF \registers_reg[30][10]  ( .D(n3964), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][10] ) );
  DFF \registers_reg[30][9]  ( .D(n3963), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][9] ) );
  DFF \registers_reg[30][8]  ( .D(n3962), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][8] ) );
  DFF \registers_reg[30][7]  ( .D(n3961), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][7] ) );
  DFF \registers_reg[30][6]  ( .D(n3960), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][6] ) );
  DFF \registers_reg[30][5]  ( .D(n3959), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][5] ) );
  DFF \registers_reg[30][4]  ( .D(n3958), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][4] ) );
  DFF \registers_reg[30][3]  ( .D(n3957), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][3] ) );
  DFF \registers_reg[30][2]  ( .D(n3956), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][2] ) );
  DFF \registers_reg[30][1]  ( .D(n3955), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][1] ) );
  DFF \registers_reg[30][0]  ( .D(n3954), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[30][0] ) );
  DFF \registers_reg[29][31]  ( .D(n3953), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][31] ) );
  DFF \registers_reg[29][30]  ( .D(n3952), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][30] ) );
  DFF \registers_reg[29][29]  ( .D(n3951), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][29] ) );
  DFF \registers_reg[29][28]  ( .D(n3950), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][28] ) );
  DFF \registers_reg[29][27]  ( .D(n3949), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][27] ) );
  DFF \registers_reg[29][26]  ( .D(n3948), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][26] ) );
  DFF \registers_reg[29][25]  ( .D(n3947), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][25] ) );
  DFF \registers_reg[29][24]  ( .D(n3946), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][24] ) );
  DFF \registers_reg[29][23]  ( .D(n3945), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][23] ) );
  DFF \registers_reg[29][22]  ( .D(n3944), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][22] ) );
  DFF \registers_reg[29][21]  ( .D(n3943), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][21] ) );
  DFF \registers_reg[29][20]  ( .D(n3942), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][20] ) );
  DFF \registers_reg[29][19]  ( .D(n3941), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][19] ) );
  DFF \registers_reg[29][18]  ( .D(n3940), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][18] ) );
  DFF \registers_reg[29][17]  ( .D(n3939), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][17] ) );
  DFF \registers_reg[29][16]  ( .D(n3938), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][16] ) );
  DFF \registers_reg[29][15]  ( .D(n3937), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][15] ) );
  DFF \registers_reg[29][14]  ( .D(n3936), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][14] ) );
  DFF \registers_reg[29][13]  ( .D(n3935), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][13] ) );
  DFF \registers_reg[29][12]  ( .D(n3934), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][12] ) );
  DFF \registers_reg[29][11]  ( .D(n3933), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][11] ) );
  DFF \registers_reg[29][10]  ( .D(n3932), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][10] ) );
  DFF \registers_reg[29][9]  ( .D(n3931), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][9] ) );
  DFF \registers_reg[29][8]  ( .D(n3930), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][8] ) );
  DFF \registers_reg[29][7]  ( .D(n3929), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][7] ) );
  DFF \registers_reg[29][6]  ( .D(n3928), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][6] ) );
  DFF \registers_reg[29][5]  ( .D(n3927), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][5] ) );
  DFF \registers_reg[29][4]  ( .D(n3926), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][4] ) );
  DFF \registers_reg[29][3]  ( .D(n3925), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][3] ) );
  DFF \registers_reg[29][2]  ( .D(n3924), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][2] ) );
  DFF \registers_reg[29][1]  ( .D(n3923), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][1] ) );
  DFF \registers_reg[29][0]  ( .D(n3922), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[29][0] ) );
  DFF \registers_reg[28][31]  ( .D(n3921), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][31] ) );
  DFF \registers_reg[28][30]  ( .D(n3920), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][30] ) );
  DFF \registers_reg[28][29]  ( .D(n3919), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][29] ) );
  DFF \registers_reg[28][28]  ( .D(n3918), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][28] ) );
  DFF \registers_reg[28][27]  ( .D(n3917), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][27] ) );
  DFF \registers_reg[28][26]  ( .D(n3916), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][26] ) );
  DFF \registers_reg[28][25]  ( .D(n3915), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][25] ) );
  DFF \registers_reg[28][24]  ( .D(n3914), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][24] ) );
  DFF \registers_reg[28][23]  ( .D(n3913), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][23] ) );
  DFF \registers_reg[28][22]  ( .D(n3912), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][22] ) );
  DFF \registers_reg[28][21]  ( .D(n3911), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][21] ) );
  DFF \registers_reg[28][20]  ( .D(n3910), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][20] ) );
  DFF \registers_reg[28][19]  ( .D(n3909), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][19] ) );
  DFF \registers_reg[28][18]  ( .D(n3908), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][18] ) );
  DFF \registers_reg[28][17]  ( .D(n3907), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][17] ) );
  DFF \registers_reg[28][16]  ( .D(n3906), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][16] ) );
  DFF \registers_reg[28][15]  ( .D(n3905), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][15] ) );
  DFF \registers_reg[28][14]  ( .D(n3904), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][14] ) );
  DFF \registers_reg[28][13]  ( .D(n3903), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][13] ) );
  DFF \registers_reg[28][12]  ( .D(n3902), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][12] ) );
  DFF \registers_reg[28][11]  ( .D(n3901), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][11] ) );
  DFF \registers_reg[28][10]  ( .D(n3900), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][10] ) );
  DFF \registers_reg[28][9]  ( .D(n3899), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][9] ) );
  DFF \registers_reg[28][8]  ( .D(n3898), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][8] ) );
  DFF \registers_reg[28][7]  ( .D(n3897), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][7] ) );
  DFF \registers_reg[28][6]  ( .D(n3896), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][6] ) );
  DFF \registers_reg[28][5]  ( .D(n3895), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][5] ) );
  DFF \registers_reg[28][4]  ( .D(n3894), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][4] ) );
  DFF \registers_reg[28][3]  ( .D(n3893), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][3] ) );
  DFF \registers_reg[28][2]  ( .D(n3892), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][2] ) );
  DFF \registers_reg[28][1]  ( .D(n3891), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][1] ) );
  DFF \registers_reg[28][0]  ( .D(n3890), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[28][0] ) );
  DFF \registers_reg[27][31]  ( .D(n3889), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][31] ) );
  DFF \registers_reg[27][30]  ( .D(n3888), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][30] ) );
  DFF \registers_reg[27][29]  ( .D(n3887), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][29] ) );
  DFF \registers_reg[27][28]  ( .D(n3886), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][28] ) );
  DFF \registers_reg[27][27]  ( .D(n3885), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][27] ) );
  DFF \registers_reg[27][26]  ( .D(n3884), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][26] ) );
  DFF \registers_reg[27][25]  ( .D(n3883), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][25] ) );
  DFF \registers_reg[27][24]  ( .D(n3882), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][24] ) );
  DFF \registers_reg[27][23]  ( .D(n3881), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][23] ) );
  DFF \registers_reg[27][22]  ( .D(n3880), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][22] ) );
  DFF \registers_reg[27][21]  ( .D(n3879), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][21] ) );
  DFF \registers_reg[27][20]  ( .D(n3878), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][20] ) );
  DFF \registers_reg[27][19]  ( .D(n3877), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][19] ) );
  DFF \registers_reg[27][18]  ( .D(n3876), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][18] ) );
  DFF \registers_reg[27][17]  ( .D(n3875), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][17] ) );
  DFF \registers_reg[27][16]  ( .D(n3874), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][16] ) );
  DFF \registers_reg[27][15]  ( .D(n3873), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][15] ) );
  DFF \registers_reg[27][14]  ( .D(n3872), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][14] ) );
  DFF \registers_reg[27][13]  ( .D(n3871), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][13] ) );
  DFF \registers_reg[27][12]  ( .D(n3870), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][12] ) );
  DFF \registers_reg[27][11]  ( .D(n3869), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][11] ) );
  DFF \registers_reg[27][10]  ( .D(n3868), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][10] ) );
  DFF \registers_reg[27][9]  ( .D(n3867), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][9] ) );
  DFF \registers_reg[27][8]  ( .D(n3866), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][8] ) );
  DFF \registers_reg[27][7]  ( .D(n3865), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][7] ) );
  DFF \registers_reg[27][6]  ( .D(n3864), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][6] ) );
  DFF \registers_reg[27][5]  ( .D(n3863), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][5] ) );
  DFF \registers_reg[27][4]  ( .D(n3862), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][4] ) );
  DFF \registers_reg[27][3]  ( .D(n3861), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][3] ) );
  DFF \registers_reg[27][2]  ( .D(n3860), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][2] ) );
  DFF \registers_reg[27][1]  ( .D(n3859), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][1] ) );
  DFF \registers_reg[27][0]  ( .D(n3858), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[27][0] ) );
  DFF \registers_reg[26][31]  ( .D(n3857), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][31] ) );
  DFF \registers_reg[26][30]  ( .D(n3856), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][30] ) );
  DFF \registers_reg[26][29]  ( .D(n3855), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][29] ) );
  DFF \registers_reg[26][28]  ( .D(n3854), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][28] ) );
  DFF \registers_reg[26][27]  ( .D(n3853), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][27] ) );
  DFF \registers_reg[26][26]  ( .D(n3852), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][26] ) );
  DFF \registers_reg[26][25]  ( .D(n3851), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][25] ) );
  DFF \registers_reg[26][24]  ( .D(n3850), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][24] ) );
  DFF \registers_reg[26][23]  ( .D(n3849), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][23] ) );
  DFF \registers_reg[26][22]  ( .D(n3848), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][22] ) );
  DFF \registers_reg[26][21]  ( .D(n3847), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][21] ) );
  DFF \registers_reg[26][20]  ( .D(n3846), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][20] ) );
  DFF \registers_reg[26][19]  ( .D(n3845), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][19] ) );
  DFF \registers_reg[26][18]  ( .D(n3844), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][18] ) );
  DFF \registers_reg[26][17]  ( .D(n3843), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][17] ) );
  DFF \registers_reg[26][16]  ( .D(n3842), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][16] ) );
  DFF \registers_reg[26][15]  ( .D(n3841), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][15] ) );
  DFF \registers_reg[26][14]  ( .D(n3840), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][14] ) );
  DFF \registers_reg[26][13]  ( .D(n3839), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][13] ) );
  DFF \registers_reg[26][12]  ( .D(n3838), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][12] ) );
  DFF \registers_reg[26][11]  ( .D(n3837), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][11] ) );
  DFF \registers_reg[26][10]  ( .D(n3836), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][10] ) );
  DFF \registers_reg[26][9]  ( .D(n3835), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][9] ) );
  DFF \registers_reg[26][8]  ( .D(n3834), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][8] ) );
  DFF \registers_reg[26][7]  ( .D(n3833), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][7] ) );
  DFF \registers_reg[26][6]  ( .D(n3832), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][6] ) );
  DFF \registers_reg[26][5]  ( .D(n3831), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][5] ) );
  DFF \registers_reg[26][4]  ( .D(n3830), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][4] ) );
  DFF \registers_reg[26][3]  ( .D(n3829), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][3] ) );
  DFF \registers_reg[26][2]  ( .D(n3828), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][2] ) );
  DFF \registers_reg[26][1]  ( .D(n3827), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][1] ) );
  DFF \registers_reg[26][0]  ( .D(n3826), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[26][0] ) );
  DFF \registers_reg[25][31]  ( .D(n3825), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][31] ) );
  DFF \registers_reg[25][30]  ( .D(n3824), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][30] ) );
  DFF \registers_reg[25][29]  ( .D(n3823), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][29] ) );
  DFF \registers_reg[25][28]  ( .D(n3822), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][28] ) );
  DFF \registers_reg[25][27]  ( .D(n3821), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][27] ) );
  DFF \registers_reg[25][26]  ( .D(n3820), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][26] ) );
  DFF \registers_reg[25][25]  ( .D(n3819), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][25] ) );
  DFF \registers_reg[25][24]  ( .D(n3818), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][24] ) );
  DFF \registers_reg[25][23]  ( .D(n3817), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][23] ) );
  DFF \registers_reg[25][22]  ( .D(n3816), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][22] ) );
  DFF \registers_reg[25][21]  ( .D(n3815), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][21] ) );
  DFF \registers_reg[25][20]  ( .D(n3814), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][20] ) );
  DFF \registers_reg[25][19]  ( .D(n3813), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][19] ) );
  DFF \registers_reg[25][18]  ( .D(n3812), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][18] ) );
  DFF \registers_reg[25][17]  ( .D(n3811), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][17] ) );
  DFF \registers_reg[25][16]  ( .D(n3810), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][16] ) );
  DFF \registers_reg[25][15]  ( .D(n3809), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][15] ) );
  DFF \registers_reg[25][14]  ( .D(n3808), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][14] ) );
  DFF \registers_reg[25][13]  ( .D(n3807), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][13] ) );
  DFF \registers_reg[25][12]  ( .D(n3806), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][12] ) );
  DFF \registers_reg[25][11]  ( .D(n3805), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][11] ) );
  DFF \registers_reg[25][10]  ( .D(n3804), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][10] ) );
  DFF \registers_reg[25][9]  ( .D(n3803), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][9] ) );
  DFF \registers_reg[25][8]  ( .D(n3802), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][8] ) );
  DFF \registers_reg[25][7]  ( .D(n3801), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][7] ) );
  DFF \registers_reg[25][6]  ( .D(n3800), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][6] ) );
  DFF \registers_reg[25][5]  ( .D(n3799), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][5] ) );
  DFF \registers_reg[25][4]  ( .D(n3798), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][4] ) );
  DFF \registers_reg[25][3]  ( .D(n3797), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][3] ) );
  DFF \registers_reg[25][2]  ( .D(n3796), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][2] ) );
  DFF \registers_reg[25][1]  ( .D(n3795), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][1] ) );
  DFF \registers_reg[25][0]  ( .D(n3794), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[25][0] ) );
  DFF \registers_reg[24][31]  ( .D(n3793), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][31] ) );
  DFF \registers_reg[24][30]  ( .D(n3792), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][30] ) );
  DFF \registers_reg[24][29]  ( .D(n3791), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][29] ) );
  DFF \registers_reg[24][28]  ( .D(n3790), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][28] ) );
  DFF \registers_reg[24][27]  ( .D(n3789), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][27] ) );
  DFF \registers_reg[24][26]  ( .D(n3788), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][26] ) );
  DFF \registers_reg[24][25]  ( .D(n3787), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][25] ) );
  DFF \registers_reg[24][24]  ( .D(n3786), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][24] ) );
  DFF \registers_reg[24][23]  ( .D(n3785), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][23] ) );
  DFF \registers_reg[24][22]  ( .D(n3784), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][22] ) );
  DFF \registers_reg[24][21]  ( .D(n3783), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][21] ) );
  DFF \registers_reg[24][20]  ( .D(n3782), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][20] ) );
  DFF \registers_reg[24][19]  ( .D(n3781), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][19] ) );
  DFF \registers_reg[24][18]  ( .D(n3780), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][18] ) );
  DFF \registers_reg[24][17]  ( .D(n3779), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][17] ) );
  DFF \registers_reg[24][16]  ( .D(n3778), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][16] ) );
  DFF \registers_reg[24][15]  ( .D(n3777), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][15] ) );
  DFF \registers_reg[24][14]  ( .D(n3776), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][14] ) );
  DFF \registers_reg[24][13]  ( .D(n3775), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][13] ) );
  DFF \registers_reg[24][12]  ( .D(n3774), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][12] ) );
  DFF \registers_reg[24][11]  ( .D(n3773), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][11] ) );
  DFF \registers_reg[24][10]  ( .D(n3772), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][10] ) );
  DFF \registers_reg[24][9]  ( .D(n3771), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][9] ) );
  DFF \registers_reg[24][8]  ( .D(n3770), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][8] ) );
  DFF \registers_reg[24][7]  ( .D(n3769), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][7] ) );
  DFF \registers_reg[24][6]  ( .D(n3768), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][6] ) );
  DFF \registers_reg[24][5]  ( .D(n3767), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][5] ) );
  DFF \registers_reg[24][4]  ( .D(n3766), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][4] ) );
  DFF \registers_reg[24][3]  ( .D(n3765), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][3] ) );
  DFF \registers_reg[24][2]  ( .D(n3764), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][2] ) );
  DFF \registers_reg[24][1]  ( .D(n3763), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][1] ) );
  DFF \registers_reg[24][0]  ( .D(n3762), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[24][0] ) );
  DFF \registers_reg[23][31]  ( .D(n3761), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][31] ) );
  DFF \registers_reg[23][30]  ( .D(n3760), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][30] ) );
  DFF \registers_reg[23][29]  ( .D(n3759), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][29] ) );
  DFF \registers_reg[23][28]  ( .D(n3758), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][28] ) );
  DFF \registers_reg[23][27]  ( .D(n3757), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][27] ) );
  DFF \registers_reg[23][26]  ( .D(n3756), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][26] ) );
  DFF \registers_reg[23][25]  ( .D(n3755), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][25] ) );
  DFF \registers_reg[23][24]  ( .D(n3754), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][24] ) );
  DFF \registers_reg[23][23]  ( .D(n3753), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][23] ) );
  DFF \registers_reg[23][22]  ( .D(n3752), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][22] ) );
  DFF \registers_reg[23][21]  ( .D(n3751), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][21] ) );
  DFF \registers_reg[23][20]  ( .D(n3750), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][20] ) );
  DFF \registers_reg[23][19]  ( .D(n3749), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][19] ) );
  DFF \registers_reg[23][18]  ( .D(n3748), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][18] ) );
  DFF \registers_reg[23][17]  ( .D(n3747), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][17] ) );
  DFF \registers_reg[23][16]  ( .D(n3746), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][16] ) );
  DFF \registers_reg[23][15]  ( .D(n3745), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][15] ) );
  DFF \registers_reg[23][14]  ( .D(n3744), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][14] ) );
  DFF \registers_reg[23][13]  ( .D(n3743), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][13] ) );
  DFF \registers_reg[23][12]  ( .D(n3742), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][12] ) );
  DFF \registers_reg[23][11]  ( .D(n3741), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][11] ) );
  DFF \registers_reg[23][10]  ( .D(n3740), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][10] ) );
  DFF \registers_reg[23][9]  ( .D(n3739), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][9] ) );
  DFF \registers_reg[23][8]  ( .D(n3738), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][8] ) );
  DFF \registers_reg[23][7]  ( .D(n3737), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][7] ) );
  DFF \registers_reg[23][6]  ( .D(n3736), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][6] ) );
  DFF \registers_reg[23][5]  ( .D(n3735), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][5] ) );
  DFF \registers_reg[23][4]  ( .D(n3734), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][4] ) );
  DFF \registers_reg[23][3]  ( .D(n3733), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][3] ) );
  DFF \registers_reg[23][2]  ( .D(n3732), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][2] ) );
  DFF \registers_reg[23][1]  ( .D(n3731), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][1] ) );
  DFF \registers_reg[23][0]  ( .D(n3730), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[23][0] ) );
  DFF \registers_reg[22][31]  ( .D(n3729), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][31] ) );
  DFF \registers_reg[22][30]  ( .D(n3728), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][30] ) );
  DFF \registers_reg[22][29]  ( .D(n3727), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][29] ) );
  DFF \registers_reg[22][28]  ( .D(n3726), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][28] ) );
  DFF \registers_reg[22][27]  ( .D(n3725), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][27] ) );
  DFF \registers_reg[22][26]  ( .D(n3724), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][26] ) );
  DFF \registers_reg[22][25]  ( .D(n3723), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][25] ) );
  DFF \registers_reg[22][24]  ( .D(n3722), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][24] ) );
  DFF \registers_reg[22][23]  ( .D(n3721), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][23] ) );
  DFF \registers_reg[22][22]  ( .D(n3720), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][22] ) );
  DFF \registers_reg[22][21]  ( .D(n3719), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][21] ) );
  DFF \registers_reg[22][20]  ( .D(n3718), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][20] ) );
  DFF \registers_reg[22][19]  ( .D(n3717), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][19] ) );
  DFF \registers_reg[22][18]  ( .D(n3716), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][18] ) );
  DFF \registers_reg[22][17]  ( .D(n3715), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][17] ) );
  DFF \registers_reg[22][16]  ( .D(n3714), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][16] ) );
  DFF \registers_reg[22][15]  ( .D(n3713), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][15] ) );
  DFF \registers_reg[22][14]  ( .D(n3712), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][14] ) );
  DFF \registers_reg[22][13]  ( .D(n3711), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][13] ) );
  DFF \registers_reg[22][12]  ( .D(n3710), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][12] ) );
  DFF \registers_reg[22][11]  ( .D(n3709), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][11] ) );
  DFF \registers_reg[22][10]  ( .D(n3708), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][10] ) );
  DFF \registers_reg[22][9]  ( .D(n3707), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][9] ) );
  DFF \registers_reg[22][8]  ( .D(n3706), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][8] ) );
  DFF \registers_reg[22][7]  ( .D(n3705), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][7] ) );
  DFF \registers_reg[22][6]  ( .D(n3704), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][6] ) );
  DFF \registers_reg[22][5]  ( .D(n3703), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][5] ) );
  DFF \registers_reg[22][4]  ( .D(n3702), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][4] ) );
  DFF \registers_reg[22][3]  ( .D(n3701), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][3] ) );
  DFF \registers_reg[22][2]  ( .D(n3700), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][2] ) );
  DFF \registers_reg[22][1]  ( .D(n3699), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][1] ) );
  DFF \registers_reg[22][0]  ( .D(n3698), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[22][0] ) );
  DFF \registers_reg[21][31]  ( .D(n3697), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][31] ) );
  DFF \registers_reg[21][30]  ( .D(n3696), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][30] ) );
  DFF \registers_reg[21][29]  ( .D(n3695), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][29] ) );
  DFF \registers_reg[21][28]  ( .D(n3694), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][28] ) );
  DFF \registers_reg[21][27]  ( .D(n3693), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][27] ) );
  DFF \registers_reg[21][26]  ( .D(n3692), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][26] ) );
  DFF \registers_reg[21][25]  ( .D(n3691), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][25] ) );
  DFF \registers_reg[21][24]  ( .D(n3690), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][24] ) );
  DFF \registers_reg[21][23]  ( .D(n3689), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][23] ) );
  DFF \registers_reg[21][22]  ( .D(n3688), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][22] ) );
  DFF \registers_reg[21][21]  ( .D(n3687), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][21] ) );
  DFF \registers_reg[21][20]  ( .D(n3686), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][20] ) );
  DFF \registers_reg[21][19]  ( .D(n3685), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][19] ) );
  DFF \registers_reg[21][18]  ( .D(n3684), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][18] ) );
  DFF \registers_reg[21][17]  ( .D(n3683), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][17] ) );
  DFF \registers_reg[21][16]  ( .D(n3682), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][16] ) );
  DFF \registers_reg[21][15]  ( .D(n3681), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][15] ) );
  DFF \registers_reg[21][14]  ( .D(n3680), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][14] ) );
  DFF \registers_reg[21][13]  ( .D(n3679), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][13] ) );
  DFF \registers_reg[21][12]  ( .D(n3678), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][12] ) );
  DFF \registers_reg[21][11]  ( .D(n3677), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][11] ) );
  DFF \registers_reg[21][10]  ( .D(n3676), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][10] ) );
  DFF \registers_reg[21][9]  ( .D(n3675), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][9] ) );
  DFF \registers_reg[21][8]  ( .D(n3674), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][8] ) );
  DFF \registers_reg[21][7]  ( .D(n3673), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][7] ) );
  DFF \registers_reg[21][6]  ( .D(n3672), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][6] ) );
  DFF \registers_reg[21][5]  ( .D(n3671), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][5] ) );
  DFF \registers_reg[21][4]  ( .D(n3670), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][4] ) );
  DFF \registers_reg[21][3]  ( .D(n3669), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][3] ) );
  DFF \registers_reg[21][2]  ( .D(n3668), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][2] ) );
  DFF \registers_reg[21][1]  ( .D(n3667), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][1] ) );
  DFF \registers_reg[21][0]  ( .D(n3666), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[21][0] ) );
  DFF \registers_reg[20][31]  ( .D(n3665), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][31] ) );
  DFF \registers_reg[20][30]  ( .D(n3664), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][30] ) );
  DFF \registers_reg[20][29]  ( .D(n3663), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][29] ) );
  DFF \registers_reg[20][28]  ( .D(n3662), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][28] ) );
  DFF \registers_reg[20][27]  ( .D(n3661), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][27] ) );
  DFF \registers_reg[20][26]  ( .D(n3660), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][26] ) );
  DFF \registers_reg[20][25]  ( .D(n3659), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][25] ) );
  DFF \registers_reg[20][24]  ( .D(n3658), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][24] ) );
  DFF \registers_reg[20][23]  ( .D(n3657), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][23] ) );
  DFF \registers_reg[20][22]  ( .D(n3656), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][22] ) );
  DFF \registers_reg[20][21]  ( .D(n3655), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][21] ) );
  DFF \registers_reg[20][20]  ( .D(n3654), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][20] ) );
  DFF \registers_reg[20][19]  ( .D(n3653), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][19] ) );
  DFF \registers_reg[20][18]  ( .D(n3652), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][18] ) );
  DFF \registers_reg[20][17]  ( .D(n3651), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][17] ) );
  DFF \registers_reg[20][16]  ( .D(n3650), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][16] ) );
  DFF \registers_reg[20][15]  ( .D(n3649), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][15] ) );
  DFF \registers_reg[20][14]  ( .D(n3648), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][14] ) );
  DFF \registers_reg[20][13]  ( .D(n3647), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][13] ) );
  DFF \registers_reg[20][12]  ( .D(n3646), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][12] ) );
  DFF \registers_reg[20][11]  ( .D(n3645), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][11] ) );
  DFF \registers_reg[20][10]  ( .D(n3644), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][10] ) );
  DFF \registers_reg[20][9]  ( .D(n3643), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][9] ) );
  DFF \registers_reg[20][8]  ( .D(n3642), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][8] ) );
  DFF \registers_reg[20][7]  ( .D(n3641), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][7] ) );
  DFF \registers_reg[20][6]  ( .D(n3640), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][6] ) );
  DFF \registers_reg[20][5]  ( .D(n3639), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][5] ) );
  DFF \registers_reg[20][4]  ( .D(n3638), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][4] ) );
  DFF \registers_reg[20][3]  ( .D(n3637), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][3] ) );
  DFF \registers_reg[20][2]  ( .D(n3636), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][2] ) );
  DFF \registers_reg[20][1]  ( .D(n3635), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][1] ) );
  DFF \registers_reg[20][0]  ( .D(n3634), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[20][0] ) );
  DFF \registers_reg[19][31]  ( .D(n3633), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][31] ) );
  DFF \registers_reg[19][30]  ( .D(n3632), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][30] ) );
  DFF \registers_reg[19][29]  ( .D(n3631), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][29] ) );
  DFF \registers_reg[19][28]  ( .D(n3630), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][28] ) );
  DFF \registers_reg[19][27]  ( .D(n3629), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][27] ) );
  DFF \registers_reg[19][26]  ( .D(n3628), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][26] ) );
  DFF \registers_reg[19][25]  ( .D(n3627), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][25] ) );
  DFF \registers_reg[19][24]  ( .D(n3626), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][24] ) );
  DFF \registers_reg[19][23]  ( .D(n3625), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][23] ) );
  DFF \registers_reg[19][22]  ( .D(n3624), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][22] ) );
  DFF \registers_reg[19][21]  ( .D(n3623), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][21] ) );
  DFF \registers_reg[19][20]  ( .D(n3622), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][20] ) );
  DFF \registers_reg[19][19]  ( .D(n3621), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][19] ) );
  DFF \registers_reg[19][18]  ( .D(n3620), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][18] ) );
  DFF \registers_reg[19][17]  ( .D(n3619), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][17] ) );
  DFF \registers_reg[19][16]  ( .D(n3618), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][16] ) );
  DFF \registers_reg[19][15]  ( .D(n3617), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][15] ) );
  DFF \registers_reg[19][14]  ( .D(n3616), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][14] ) );
  DFF \registers_reg[19][13]  ( .D(n3615), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][13] ) );
  DFF \registers_reg[19][12]  ( .D(n3614), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][12] ) );
  DFF \registers_reg[19][11]  ( .D(n3613), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][11] ) );
  DFF \registers_reg[19][10]  ( .D(n3612), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][10] ) );
  DFF \registers_reg[19][9]  ( .D(n3611), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][9] ) );
  DFF \registers_reg[19][8]  ( .D(n3610), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][8] ) );
  DFF \registers_reg[19][7]  ( .D(n3609), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][7] ) );
  DFF \registers_reg[19][6]  ( .D(n3608), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][6] ) );
  DFF \registers_reg[19][5]  ( .D(n3607), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][5] ) );
  DFF \registers_reg[19][4]  ( .D(n3606), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][4] ) );
  DFF \registers_reg[19][3]  ( .D(n3605), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][3] ) );
  DFF \registers_reg[19][2]  ( .D(n3604), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][2] ) );
  DFF \registers_reg[19][1]  ( .D(n3603), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][1] ) );
  DFF \registers_reg[19][0]  ( .D(n3602), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[19][0] ) );
  DFF \registers_reg[18][31]  ( .D(n3601), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][31] ) );
  DFF \registers_reg[18][30]  ( .D(n3600), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][30] ) );
  DFF \registers_reg[18][29]  ( .D(n3599), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][29] ) );
  DFF \registers_reg[18][28]  ( .D(n3598), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][28] ) );
  DFF \registers_reg[18][27]  ( .D(n3597), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][27] ) );
  DFF \registers_reg[18][26]  ( .D(n3596), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][26] ) );
  DFF \registers_reg[18][25]  ( .D(n3595), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][25] ) );
  DFF \registers_reg[18][24]  ( .D(n3594), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][24] ) );
  DFF \registers_reg[18][23]  ( .D(n3593), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][23] ) );
  DFF \registers_reg[18][22]  ( .D(n3592), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][22] ) );
  DFF \registers_reg[18][21]  ( .D(n3591), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][21] ) );
  DFF \registers_reg[18][20]  ( .D(n3590), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][20] ) );
  DFF \registers_reg[18][19]  ( .D(n3589), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][19] ) );
  DFF \registers_reg[18][18]  ( .D(n3588), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][18] ) );
  DFF \registers_reg[18][17]  ( .D(n3587), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][17] ) );
  DFF \registers_reg[18][16]  ( .D(n3586), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][16] ) );
  DFF \registers_reg[18][15]  ( .D(n3585), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][15] ) );
  DFF \registers_reg[18][14]  ( .D(n3584), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][14] ) );
  DFF \registers_reg[18][13]  ( .D(n3583), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][13] ) );
  DFF \registers_reg[18][12]  ( .D(n3582), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][12] ) );
  DFF \registers_reg[18][11]  ( .D(n3581), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][11] ) );
  DFF \registers_reg[18][10]  ( .D(n3580), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][10] ) );
  DFF \registers_reg[18][9]  ( .D(n3579), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][9] ) );
  DFF \registers_reg[18][8]  ( .D(n3578), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][8] ) );
  DFF \registers_reg[18][7]  ( .D(n3577), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][7] ) );
  DFF \registers_reg[18][6]  ( .D(n3576), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][6] ) );
  DFF \registers_reg[18][5]  ( .D(n3575), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][5] ) );
  DFF \registers_reg[18][4]  ( .D(n3574), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][4] ) );
  DFF \registers_reg[18][3]  ( .D(n3573), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][3] ) );
  DFF \registers_reg[18][2]  ( .D(n3572), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][2] ) );
  DFF \registers_reg[18][1]  ( .D(n3571), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][1] ) );
  DFF \registers_reg[18][0]  ( .D(n3570), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[18][0] ) );
  DFF \registers_reg[17][31]  ( .D(n3569), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][31] ) );
  DFF \registers_reg[17][30]  ( .D(n3568), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][30] ) );
  DFF \registers_reg[17][29]  ( .D(n3567), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][29] ) );
  DFF \registers_reg[17][28]  ( .D(n3566), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][28] ) );
  DFF \registers_reg[17][27]  ( .D(n3565), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][27] ) );
  DFF \registers_reg[17][26]  ( .D(n3564), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][26] ) );
  DFF \registers_reg[17][25]  ( .D(n3563), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][25] ) );
  DFF \registers_reg[17][24]  ( .D(n3562), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][24] ) );
  DFF \registers_reg[17][23]  ( .D(n3561), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][23] ) );
  DFF \registers_reg[17][22]  ( .D(n3560), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][22] ) );
  DFF \registers_reg[17][21]  ( .D(n3559), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][21] ) );
  DFF \registers_reg[17][20]  ( .D(n3558), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][20] ) );
  DFF \registers_reg[17][19]  ( .D(n3557), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][19] ) );
  DFF \registers_reg[17][18]  ( .D(n3556), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][18] ) );
  DFF \registers_reg[17][17]  ( .D(n3555), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][17] ) );
  DFF \registers_reg[17][16]  ( .D(n3554), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][16] ) );
  DFF \registers_reg[17][15]  ( .D(n3553), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][15] ) );
  DFF \registers_reg[17][14]  ( .D(n3552), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][14] ) );
  DFF \registers_reg[17][13]  ( .D(n3551), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][13] ) );
  DFF \registers_reg[17][12]  ( .D(n3550), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][12] ) );
  DFF \registers_reg[17][11]  ( .D(n3549), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][11] ) );
  DFF \registers_reg[17][10]  ( .D(n3548), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][10] ) );
  DFF \registers_reg[17][9]  ( .D(n3547), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][9] ) );
  DFF \registers_reg[17][8]  ( .D(n3546), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][8] ) );
  DFF \registers_reg[17][7]  ( .D(n3545), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][7] ) );
  DFF \registers_reg[17][6]  ( .D(n3544), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][6] ) );
  DFF \registers_reg[17][5]  ( .D(n3543), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][5] ) );
  DFF \registers_reg[17][4]  ( .D(n3542), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][4] ) );
  DFF \registers_reg[17][3]  ( .D(n3541), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][3] ) );
  DFF \registers_reg[17][2]  ( .D(n3540), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][2] ) );
  DFF \registers_reg[17][1]  ( .D(n3539), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][1] ) );
  DFF \registers_reg[17][0]  ( .D(n3538), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[17][0] ) );
  DFF \registers_reg[16][31]  ( .D(n3537), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][31] ) );
  DFF \registers_reg[16][30]  ( .D(n3536), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][30] ) );
  DFF \registers_reg[16][29]  ( .D(n3535), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][29] ) );
  DFF \registers_reg[16][28]  ( .D(n3534), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][28] ) );
  DFF \registers_reg[16][27]  ( .D(n3533), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][27] ) );
  DFF \registers_reg[16][26]  ( .D(n3532), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][26] ) );
  DFF \registers_reg[16][25]  ( .D(n3531), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][25] ) );
  DFF \registers_reg[16][24]  ( .D(n3530), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][24] ) );
  DFF \registers_reg[16][23]  ( .D(n3529), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][23] ) );
  DFF \registers_reg[16][22]  ( .D(n3528), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][22] ) );
  DFF \registers_reg[16][21]  ( .D(n3527), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][21] ) );
  DFF \registers_reg[16][20]  ( .D(n3526), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][20] ) );
  DFF \registers_reg[16][19]  ( .D(n3525), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][19] ) );
  DFF \registers_reg[16][18]  ( .D(n3524), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][18] ) );
  DFF \registers_reg[16][17]  ( .D(n3523), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][17] ) );
  DFF \registers_reg[16][16]  ( .D(n3522), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][16] ) );
  DFF \registers_reg[16][15]  ( .D(n3521), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][15] ) );
  DFF \registers_reg[16][14]  ( .D(n3520), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][14] ) );
  DFF \registers_reg[16][13]  ( .D(n3519), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][13] ) );
  DFF \registers_reg[16][12]  ( .D(n3518), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][12] ) );
  DFF \registers_reg[16][11]  ( .D(n3517), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][11] ) );
  DFF \registers_reg[16][10]  ( .D(n3516), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][10] ) );
  DFF \registers_reg[16][9]  ( .D(n3515), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][9] ) );
  DFF \registers_reg[16][8]  ( .D(n3514), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][8] ) );
  DFF \registers_reg[16][7]  ( .D(n3513), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][7] ) );
  DFF \registers_reg[16][6]  ( .D(n3512), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][6] ) );
  DFF \registers_reg[16][5]  ( .D(n3511), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][5] ) );
  DFF \registers_reg[16][4]  ( .D(n3510), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][4] ) );
  DFF \registers_reg[16][3]  ( .D(n3509), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][3] ) );
  DFF \registers_reg[16][2]  ( .D(n3508), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][2] ) );
  DFF \registers_reg[16][1]  ( .D(n3507), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][1] ) );
  DFF \registers_reg[16][0]  ( .D(n3506), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[16][0] ) );
  DFF \registers_reg[15][31]  ( .D(n3505), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][31] ) );
  DFF \registers_reg[15][30]  ( .D(n3504), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][30] ) );
  DFF \registers_reg[15][29]  ( .D(n3503), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][29] ) );
  DFF \registers_reg[15][28]  ( .D(n3502), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][28] ) );
  DFF \registers_reg[15][27]  ( .D(n3501), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][27] ) );
  DFF \registers_reg[15][26]  ( .D(n3500), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][26] ) );
  DFF \registers_reg[15][25]  ( .D(n3499), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][25] ) );
  DFF \registers_reg[15][24]  ( .D(n3498), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][24] ) );
  DFF \registers_reg[15][23]  ( .D(n3497), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][23] ) );
  DFF \registers_reg[15][22]  ( .D(n3496), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][22] ) );
  DFF \registers_reg[15][21]  ( .D(n3495), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][21] ) );
  DFF \registers_reg[15][20]  ( .D(n3494), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][20] ) );
  DFF \registers_reg[15][19]  ( .D(n3493), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][19] ) );
  DFF \registers_reg[15][18]  ( .D(n3492), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][18] ) );
  DFF \registers_reg[15][17]  ( .D(n3491), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][17] ) );
  DFF \registers_reg[15][16]  ( .D(n3490), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][16] ) );
  DFF \registers_reg[15][15]  ( .D(n3489), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][15] ) );
  DFF \registers_reg[15][14]  ( .D(n3488), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][14] ) );
  DFF \registers_reg[15][13]  ( .D(n3487), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][13] ) );
  DFF \registers_reg[15][12]  ( .D(n3486), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][12] ) );
  DFF \registers_reg[15][11]  ( .D(n3485), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][11] ) );
  DFF \registers_reg[15][10]  ( .D(n3484), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][10] ) );
  DFF \registers_reg[15][9]  ( .D(n3483), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][9] ) );
  DFF \registers_reg[15][8]  ( .D(n3482), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][8] ) );
  DFF \registers_reg[15][7]  ( .D(n3481), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][7] ) );
  DFF \registers_reg[15][6]  ( .D(n3480), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][6] ) );
  DFF \registers_reg[15][5]  ( .D(n3479), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][5] ) );
  DFF \registers_reg[15][4]  ( .D(n3478), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][4] ) );
  DFF \registers_reg[15][3]  ( .D(n3477), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][3] ) );
  DFF \registers_reg[15][2]  ( .D(n3476), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][2] ) );
  DFF \registers_reg[15][1]  ( .D(n3475), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][1] ) );
  DFF \registers_reg[15][0]  ( .D(n3474), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[15][0] ) );
  DFF \registers_reg[14][31]  ( .D(n3473), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][31] ) );
  DFF \registers_reg[14][30]  ( .D(n3472), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][30] ) );
  DFF \registers_reg[14][29]  ( .D(n3471), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][29] ) );
  DFF \registers_reg[14][28]  ( .D(n3470), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][28] ) );
  DFF \registers_reg[14][27]  ( .D(n3469), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][27] ) );
  DFF \registers_reg[14][26]  ( .D(n3468), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][26] ) );
  DFF \registers_reg[14][25]  ( .D(n3467), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][25] ) );
  DFF \registers_reg[14][24]  ( .D(n3466), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][24] ) );
  DFF \registers_reg[14][23]  ( .D(n3465), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][23] ) );
  DFF \registers_reg[14][22]  ( .D(n3464), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][22] ) );
  DFF \registers_reg[14][21]  ( .D(n3463), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][21] ) );
  DFF \registers_reg[14][20]  ( .D(n3462), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][20] ) );
  DFF \registers_reg[14][19]  ( .D(n3461), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][19] ) );
  DFF \registers_reg[14][18]  ( .D(n3460), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][18] ) );
  DFF \registers_reg[14][17]  ( .D(n3459), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][17] ) );
  DFF \registers_reg[14][16]  ( .D(n3458), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][16] ) );
  DFF \registers_reg[14][15]  ( .D(n3457), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][15] ) );
  DFF \registers_reg[14][14]  ( .D(n3456), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][14] ) );
  DFF \registers_reg[14][13]  ( .D(n3455), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][13] ) );
  DFF \registers_reg[14][12]  ( .D(n3454), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][12] ) );
  DFF \registers_reg[14][11]  ( .D(n3453), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][11] ) );
  DFF \registers_reg[14][10]  ( .D(n3452), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][10] ) );
  DFF \registers_reg[14][9]  ( .D(n3451), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][9] ) );
  DFF \registers_reg[14][8]  ( .D(n3450), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][8] ) );
  DFF \registers_reg[14][7]  ( .D(n3449), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][7] ) );
  DFF \registers_reg[14][6]  ( .D(n3448), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][6] ) );
  DFF \registers_reg[14][5]  ( .D(n3447), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][5] ) );
  DFF \registers_reg[14][4]  ( .D(n3446), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][4] ) );
  DFF \registers_reg[14][3]  ( .D(n3445), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][3] ) );
  DFF \registers_reg[14][2]  ( .D(n3444), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][2] ) );
  DFF \registers_reg[14][1]  ( .D(n3443), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][1] ) );
  DFF \registers_reg[14][0]  ( .D(n3442), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[14][0] ) );
  DFF \registers_reg[13][31]  ( .D(n3441), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][31] ) );
  DFF \registers_reg[13][30]  ( .D(n3440), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][30] ) );
  DFF \registers_reg[13][29]  ( .D(n3439), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][29] ) );
  DFF \registers_reg[13][28]  ( .D(n3438), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][28] ) );
  DFF \registers_reg[13][27]  ( .D(n3437), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][27] ) );
  DFF \registers_reg[13][26]  ( .D(n3436), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][26] ) );
  DFF \registers_reg[13][25]  ( .D(n3435), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][25] ) );
  DFF \registers_reg[13][24]  ( .D(n3434), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][24] ) );
  DFF \registers_reg[13][23]  ( .D(n3433), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][23] ) );
  DFF \registers_reg[13][22]  ( .D(n3432), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][22] ) );
  DFF \registers_reg[13][21]  ( .D(n3431), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][21] ) );
  DFF \registers_reg[13][20]  ( .D(n3430), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][20] ) );
  DFF \registers_reg[13][19]  ( .D(n3429), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][19] ) );
  DFF \registers_reg[13][18]  ( .D(n3428), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][18] ) );
  DFF \registers_reg[13][17]  ( .D(n3427), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][17] ) );
  DFF \registers_reg[13][16]  ( .D(n3426), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][16] ) );
  DFF \registers_reg[13][15]  ( .D(n3425), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][15] ) );
  DFF \registers_reg[13][14]  ( .D(n3424), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][14] ) );
  DFF \registers_reg[13][13]  ( .D(n3423), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][13] ) );
  DFF \registers_reg[13][12]  ( .D(n3422), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][12] ) );
  DFF \registers_reg[13][11]  ( .D(n3421), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][11] ) );
  DFF \registers_reg[13][10]  ( .D(n3420), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][10] ) );
  DFF \registers_reg[13][9]  ( .D(n3419), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][9] ) );
  DFF \registers_reg[13][8]  ( .D(n3418), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][8] ) );
  DFF \registers_reg[13][7]  ( .D(n3417), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][7] ) );
  DFF \registers_reg[13][6]  ( .D(n3416), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][6] ) );
  DFF \registers_reg[13][5]  ( .D(n3415), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][5] ) );
  DFF \registers_reg[13][4]  ( .D(n3414), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][4] ) );
  DFF \registers_reg[13][3]  ( .D(n3413), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][3] ) );
  DFF \registers_reg[13][2]  ( .D(n3412), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][2] ) );
  DFF \registers_reg[13][1]  ( .D(n3411), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][1] ) );
  DFF \registers_reg[13][0]  ( .D(n3410), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[13][0] ) );
  DFF \registers_reg[12][31]  ( .D(n3409), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][31] ) );
  DFF \registers_reg[12][30]  ( .D(n3408), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][30] ) );
  DFF \registers_reg[12][29]  ( .D(n3407), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][29] ) );
  DFF \registers_reg[12][28]  ( .D(n3406), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][28] ) );
  DFF \registers_reg[12][27]  ( .D(n3405), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][27] ) );
  DFF \registers_reg[12][26]  ( .D(n3404), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][26] ) );
  DFF \registers_reg[12][25]  ( .D(n3403), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][25] ) );
  DFF \registers_reg[12][24]  ( .D(n3402), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][24] ) );
  DFF \registers_reg[12][23]  ( .D(n3401), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][23] ) );
  DFF \registers_reg[12][22]  ( .D(n3400), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][22] ) );
  DFF \registers_reg[12][21]  ( .D(n3399), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][21] ) );
  DFF \registers_reg[12][20]  ( .D(n3398), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][20] ) );
  DFF \registers_reg[12][19]  ( .D(n3397), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][19] ) );
  DFF \registers_reg[12][18]  ( .D(n3396), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][18] ) );
  DFF \registers_reg[12][17]  ( .D(n3395), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][17] ) );
  DFF \registers_reg[12][16]  ( .D(n3394), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][16] ) );
  DFF \registers_reg[12][15]  ( .D(n3393), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][15] ) );
  DFF \registers_reg[12][14]  ( .D(n3392), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][14] ) );
  DFF \registers_reg[12][13]  ( .D(n3391), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][13] ) );
  DFF \registers_reg[12][12]  ( .D(n3390), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][12] ) );
  DFF \registers_reg[12][11]  ( .D(n3389), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][11] ) );
  DFF \registers_reg[12][10]  ( .D(n3388), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][10] ) );
  DFF \registers_reg[12][9]  ( .D(n3387), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][9] ) );
  DFF \registers_reg[12][8]  ( .D(n3386), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][8] ) );
  DFF \registers_reg[12][7]  ( .D(n3385), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][7] ) );
  DFF \registers_reg[12][6]  ( .D(n3384), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][6] ) );
  DFF \registers_reg[12][5]  ( .D(n3383), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][5] ) );
  DFF \registers_reg[12][4]  ( .D(n3382), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][4] ) );
  DFF \registers_reg[12][3]  ( .D(n3381), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][3] ) );
  DFF \registers_reg[12][2]  ( .D(n3380), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][2] ) );
  DFF \registers_reg[12][1]  ( .D(n3379), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][1] ) );
  DFF \registers_reg[12][0]  ( .D(n3378), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[12][0] ) );
  DFF \registers_reg[11][31]  ( .D(n3377), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][31] ) );
  DFF \registers_reg[11][30]  ( .D(n3376), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][30] ) );
  DFF \registers_reg[11][29]  ( .D(n3375), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][29] ) );
  DFF \registers_reg[11][28]  ( .D(n3374), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][28] ) );
  DFF \registers_reg[11][27]  ( .D(n3373), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][27] ) );
  DFF \registers_reg[11][26]  ( .D(n3372), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][26] ) );
  DFF \registers_reg[11][25]  ( .D(n3371), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][25] ) );
  DFF \registers_reg[11][24]  ( .D(n3370), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][24] ) );
  DFF \registers_reg[11][23]  ( .D(n3369), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][23] ) );
  DFF \registers_reg[11][22]  ( .D(n3368), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][22] ) );
  DFF \registers_reg[11][21]  ( .D(n3367), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][21] ) );
  DFF \registers_reg[11][20]  ( .D(n3366), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][20] ) );
  DFF \registers_reg[11][19]  ( .D(n3365), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][19] ) );
  DFF \registers_reg[11][18]  ( .D(n3364), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][18] ) );
  DFF \registers_reg[11][17]  ( .D(n3363), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][17] ) );
  DFF \registers_reg[11][16]  ( .D(n3362), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][16] ) );
  DFF \registers_reg[11][15]  ( .D(n3361), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][15] ) );
  DFF \registers_reg[11][14]  ( .D(n3360), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][14] ) );
  DFF \registers_reg[11][13]  ( .D(n3359), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][13] ) );
  DFF \registers_reg[11][12]  ( .D(n3358), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][12] ) );
  DFF \registers_reg[11][11]  ( .D(n3357), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][11] ) );
  DFF \registers_reg[11][10]  ( .D(n3356), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][10] ) );
  DFF \registers_reg[11][9]  ( .D(n3355), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][9] ) );
  DFF \registers_reg[11][8]  ( .D(n3354), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][8] ) );
  DFF \registers_reg[11][7]  ( .D(n3353), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][7] ) );
  DFF \registers_reg[11][6]  ( .D(n3352), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][6] ) );
  DFF \registers_reg[11][5]  ( .D(n3351), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][5] ) );
  DFF \registers_reg[11][4]  ( .D(n3350), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][4] ) );
  DFF \registers_reg[11][3]  ( .D(n3349), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][3] ) );
  DFF \registers_reg[11][2]  ( .D(n3348), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][2] ) );
  DFF \registers_reg[11][1]  ( .D(n3347), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][1] ) );
  DFF \registers_reg[11][0]  ( .D(n3346), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[11][0] ) );
  DFF \registers_reg[10][31]  ( .D(n3345), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][31] ) );
  DFF \registers_reg[10][30]  ( .D(n3344), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][30] ) );
  DFF \registers_reg[10][29]  ( .D(n3343), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][29] ) );
  DFF \registers_reg[10][28]  ( .D(n3342), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][28] ) );
  DFF \registers_reg[10][27]  ( .D(n3341), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][27] ) );
  DFF \registers_reg[10][26]  ( .D(n3340), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][26] ) );
  DFF \registers_reg[10][25]  ( .D(n3339), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][25] ) );
  DFF \registers_reg[10][24]  ( .D(n3338), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][24] ) );
  DFF \registers_reg[10][23]  ( .D(n3337), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][23] ) );
  DFF \registers_reg[10][22]  ( .D(n3336), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][22] ) );
  DFF \registers_reg[10][21]  ( .D(n3335), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][21] ) );
  DFF \registers_reg[10][20]  ( .D(n3334), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][20] ) );
  DFF \registers_reg[10][19]  ( .D(n3333), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][19] ) );
  DFF \registers_reg[10][18]  ( .D(n3332), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][18] ) );
  DFF \registers_reg[10][17]  ( .D(n3331), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][17] ) );
  DFF \registers_reg[10][16]  ( .D(n3330), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][16] ) );
  DFF \registers_reg[10][15]  ( .D(n3329), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][15] ) );
  DFF \registers_reg[10][14]  ( .D(n3328), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][14] ) );
  DFF \registers_reg[10][13]  ( .D(n3327), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][13] ) );
  DFF \registers_reg[10][12]  ( .D(n3326), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][12] ) );
  DFF \registers_reg[10][11]  ( .D(n3325), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][11] ) );
  DFF \registers_reg[10][10]  ( .D(n3324), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][10] ) );
  DFF \registers_reg[10][9]  ( .D(n3323), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][9] ) );
  DFF \registers_reg[10][8]  ( .D(n3322), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][8] ) );
  DFF \registers_reg[10][7]  ( .D(n3321), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][7] ) );
  DFF \registers_reg[10][6]  ( .D(n3320), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][6] ) );
  DFF \registers_reg[10][5]  ( .D(n3319), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][5] ) );
  DFF \registers_reg[10][4]  ( .D(n3318), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][4] ) );
  DFF \registers_reg[10][3]  ( .D(n3317), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][3] ) );
  DFF \registers_reg[10][2]  ( .D(n3316), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][2] ) );
  DFF \registers_reg[10][1]  ( .D(n3315), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][1] ) );
  DFF \registers_reg[10][0]  ( .D(n3314), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[10][0] ) );
  DFF \registers_reg[9][31]  ( .D(n3313), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][31] ) );
  DFF \registers_reg[9][30]  ( .D(n3312), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][30] ) );
  DFF \registers_reg[9][29]  ( .D(n3311), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][29] ) );
  DFF \registers_reg[9][28]  ( .D(n3310), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][28] ) );
  DFF \registers_reg[9][27]  ( .D(n3309), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][27] ) );
  DFF \registers_reg[9][26]  ( .D(n3308), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][26] ) );
  DFF \registers_reg[9][25]  ( .D(n3307), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][25] ) );
  DFF \registers_reg[9][24]  ( .D(n3306), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][24] ) );
  DFF \registers_reg[9][23]  ( .D(n3305), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][23] ) );
  DFF \registers_reg[9][22]  ( .D(n3304), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][22] ) );
  DFF \registers_reg[9][21]  ( .D(n3303), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][21] ) );
  DFF \registers_reg[9][20]  ( .D(n3302), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][20] ) );
  DFF \registers_reg[9][19]  ( .D(n3301), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][19] ) );
  DFF \registers_reg[9][18]  ( .D(n3300), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][18] ) );
  DFF \registers_reg[9][17]  ( .D(n3299), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][17] ) );
  DFF \registers_reg[9][16]  ( .D(n3298), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][16] ) );
  DFF \registers_reg[9][15]  ( .D(n3297), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][15] ) );
  DFF \registers_reg[9][14]  ( .D(n3296), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][14] ) );
  DFF \registers_reg[9][13]  ( .D(n3295), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][13] ) );
  DFF \registers_reg[9][12]  ( .D(n3294), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][12] ) );
  DFF \registers_reg[9][11]  ( .D(n3293), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][11] ) );
  DFF \registers_reg[9][10]  ( .D(n3292), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][10] ) );
  DFF \registers_reg[9][9]  ( .D(n3291), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][9] ) );
  DFF \registers_reg[9][8]  ( .D(n3290), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][8] ) );
  DFF \registers_reg[9][7]  ( .D(n3289), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][7] ) );
  DFF \registers_reg[9][6]  ( .D(n3288), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][6] ) );
  DFF \registers_reg[9][5]  ( .D(n3287), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][5] ) );
  DFF \registers_reg[9][4]  ( .D(n3286), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][4] ) );
  DFF \registers_reg[9][3]  ( .D(n3285), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][3] ) );
  DFF \registers_reg[9][2]  ( .D(n3284), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][2] ) );
  DFF \registers_reg[9][1]  ( .D(n3283), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][1] ) );
  DFF \registers_reg[9][0]  ( .D(n3282), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[9][0] ) );
  DFF \registers_reg[8][31]  ( .D(n3281), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][31] ) );
  DFF \registers_reg[8][30]  ( .D(n3280), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][30] ) );
  DFF \registers_reg[8][29]  ( .D(n3279), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][29] ) );
  DFF \registers_reg[8][28]  ( .D(n3278), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][28] ) );
  DFF \registers_reg[8][27]  ( .D(n3277), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][27] ) );
  DFF \registers_reg[8][26]  ( .D(n3276), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][26] ) );
  DFF \registers_reg[8][25]  ( .D(n3275), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][25] ) );
  DFF \registers_reg[8][24]  ( .D(n3274), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][24] ) );
  DFF \registers_reg[8][23]  ( .D(n3273), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][23] ) );
  DFF \registers_reg[8][22]  ( .D(n3272), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][22] ) );
  DFF \registers_reg[8][21]  ( .D(n3271), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][21] ) );
  DFF \registers_reg[8][20]  ( .D(n3270), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][20] ) );
  DFF \registers_reg[8][19]  ( .D(n3269), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][19] ) );
  DFF \registers_reg[8][18]  ( .D(n3268), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][18] ) );
  DFF \registers_reg[8][17]  ( .D(n3267), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][17] ) );
  DFF \registers_reg[8][16]  ( .D(n3266), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][16] ) );
  DFF \registers_reg[8][15]  ( .D(n3265), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][15] ) );
  DFF \registers_reg[8][14]  ( .D(n3264), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][14] ) );
  DFF \registers_reg[8][13]  ( .D(n3263), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][13] ) );
  DFF \registers_reg[8][12]  ( .D(n3262), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][12] ) );
  DFF \registers_reg[8][11]  ( .D(n3261), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][11] ) );
  DFF \registers_reg[8][10]  ( .D(n3260), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][10] ) );
  DFF \registers_reg[8][9]  ( .D(n3259), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][9] ) );
  DFF \registers_reg[8][8]  ( .D(n3258), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][8] ) );
  DFF \registers_reg[8][7]  ( .D(n3257), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][7] ) );
  DFF \registers_reg[8][6]  ( .D(n3256), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][6] ) );
  DFF \registers_reg[8][5]  ( .D(n3255), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][5] ) );
  DFF \registers_reg[8][4]  ( .D(n3254), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][4] ) );
  DFF \registers_reg[8][3]  ( .D(n3253), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][3] ) );
  DFF \registers_reg[8][2]  ( .D(n3252), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][2] ) );
  DFF \registers_reg[8][1]  ( .D(n3251), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][1] ) );
  DFF \registers_reg[8][0]  ( .D(n3250), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[8][0] ) );
  DFF \registers_reg[7][31]  ( .D(n3249), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][31] ) );
  DFF \registers_reg[7][30]  ( .D(n3248), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][30] ) );
  DFF \registers_reg[7][29]  ( .D(n3247), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][29] ) );
  DFF \registers_reg[7][28]  ( .D(n3246), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][28] ) );
  DFF \registers_reg[7][27]  ( .D(n3245), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][27] ) );
  DFF \registers_reg[7][26]  ( .D(n3244), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][26] ) );
  DFF \registers_reg[7][25]  ( .D(n3243), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][25] ) );
  DFF \registers_reg[7][24]  ( .D(n3242), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][24] ) );
  DFF \registers_reg[7][23]  ( .D(n3241), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][23] ) );
  DFF \registers_reg[7][22]  ( .D(n3240), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][22] ) );
  DFF \registers_reg[7][21]  ( .D(n3239), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][21] ) );
  DFF \registers_reg[7][20]  ( .D(n3238), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][20] ) );
  DFF \registers_reg[7][19]  ( .D(n3237), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][19] ) );
  DFF \registers_reg[7][18]  ( .D(n3236), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][18] ) );
  DFF \registers_reg[7][17]  ( .D(n3235), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][17] ) );
  DFF \registers_reg[7][16]  ( .D(n3234), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][16] ) );
  DFF \registers_reg[7][15]  ( .D(n3233), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][15] ) );
  DFF \registers_reg[7][14]  ( .D(n3232), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][14] ) );
  DFF \registers_reg[7][13]  ( .D(n3231), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][13] ) );
  DFF \registers_reg[7][12]  ( .D(n3230), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][12] ) );
  DFF \registers_reg[7][11]  ( .D(n3229), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][11] ) );
  DFF \registers_reg[7][10]  ( .D(n3228), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][10] ) );
  DFF \registers_reg[7][9]  ( .D(n3227), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][9] ) );
  DFF \registers_reg[7][8]  ( .D(n3226), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][8] ) );
  DFF \registers_reg[7][7]  ( .D(n3225), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][7] ) );
  DFF \registers_reg[7][6]  ( .D(n3224), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][6] ) );
  DFF \registers_reg[7][5]  ( .D(n3223), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][5] ) );
  DFF \registers_reg[7][4]  ( .D(n3222), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][4] ) );
  DFF \registers_reg[7][3]  ( .D(n3221), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][3] ) );
  DFF \registers_reg[7][2]  ( .D(n3220), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][2] ) );
  DFF \registers_reg[7][1]  ( .D(n3219), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][1] ) );
  DFF \registers_reg[7][0]  ( .D(n3218), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[7][0] ) );
  DFF \registers_reg[6][31]  ( .D(n3217), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][31] ) );
  DFF \registers_reg[6][30]  ( .D(n3216), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][30] ) );
  DFF \registers_reg[6][29]  ( .D(n3215), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][29] ) );
  DFF \registers_reg[6][28]  ( .D(n3214), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][28] ) );
  DFF \registers_reg[6][27]  ( .D(n3213), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][27] ) );
  DFF \registers_reg[6][26]  ( .D(n3212), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][26] ) );
  DFF \registers_reg[6][25]  ( .D(n3211), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][25] ) );
  DFF \registers_reg[6][24]  ( .D(n3210), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][24] ) );
  DFF \registers_reg[6][23]  ( .D(n3209), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][23] ) );
  DFF \registers_reg[6][22]  ( .D(n3208), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][22] ) );
  DFF \registers_reg[6][21]  ( .D(n3207), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][21] ) );
  DFF \registers_reg[6][20]  ( .D(n3206), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][20] ) );
  DFF \registers_reg[6][19]  ( .D(n3205), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][19] ) );
  DFF \registers_reg[6][18]  ( .D(n3204), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][18] ) );
  DFF \registers_reg[6][17]  ( .D(n3203), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][17] ) );
  DFF \registers_reg[6][16]  ( .D(n3202), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][16] ) );
  DFF \registers_reg[6][15]  ( .D(n3201), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][15] ) );
  DFF \registers_reg[6][14]  ( .D(n3200), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][14] ) );
  DFF \registers_reg[6][13]  ( .D(n3199), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][13] ) );
  DFF \registers_reg[6][12]  ( .D(n3198), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][12] ) );
  DFF \registers_reg[6][11]  ( .D(n3197), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][11] ) );
  DFF \registers_reg[6][10]  ( .D(n3196), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][10] ) );
  DFF \registers_reg[6][9]  ( .D(n3195), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][9] ) );
  DFF \registers_reg[6][8]  ( .D(n3194), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][8] ) );
  DFF \registers_reg[6][7]  ( .D(n3193), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][7] ) );
  DFF \registers_reg[6][6]  ( .D(n3192), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][6] ) );
  DFF \registers_reg[6][5]  ( .D(n3191), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][5] ) );
  DFF \registers_reg[6][4]  ( .D(n3190), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][4] ) );
  DFF \registers_reg[6][3]  ( .D(n3189), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][3] ) );
  DFF \registers_reg[6][2]  ( .D(n3188), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][2] ) );
  DFF \registers_reg[6][1]  ( .D(n3187), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][1] ) );
  DFF \registers_reg[6][0]  ( .D(n3186), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[6][0] ) );
  DFF \registers_reg[5][31]  ( .D(n3185), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][31] ) );
  DFF \registers_reg[5][30]  ( .D(n3184), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][30] ) );
  DFF \registers_reg[5][29]  ( .D(n3183), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][29] ) );
  DFF \registers_reg[5][28]  ( .D(n3182), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][28] ) );
  DFF \registers_reg[5][27]  ( .D(n3181), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][27] ) );
  DFF \registers_reg[5][26]  ( .D(n3180), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][26] ) );
  DFF \registers_reg[5][25]  ( .D(n3179), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][25] ) );
  DFF \registers_reg[5][24]  ( .D(n3178), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][24] ) );
  DFF \registers_reg[5][23]  ( .D(n3177), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][23] ) );
  DFF \registers_reg[5][22]  ( .D(n3176), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][22] ) );
  DFF \registers_reg[5][21]  ( .D(n3175), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][21] ) );
  DFF \registers_reg[5][20]  ( .D(n3174), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][20] ) );
  DFF \registers_reg[5][19]  ( .D(n3173), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][19] ) );
  DFF \registers_reg[5][18]  ( .D(n3172), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][18] ) );
  DFF \registers_reg[5][17]  ( .D(n3171), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][17] ) );
  DFF \registers_reg[5][16]  ( .D(n3170), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][16] ) );
  DFF \registers_reg[5][15]  ( .D(n3169), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][15] ) );
  DFF \registers_reg[5][14]  ( .D(n3168), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][14] ) );
  DFF \registers_reg[5][13]  ( .D(n3167), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][13] ) );
  DFF \registers_reg[5][12]  ( .D(n3166), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][12] ) );
  DFF \registers_reg[5][11]  ( .D(n3165), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][11] ) );
  DFF \registers_reg[5][10]  ( .D(n3164), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][10] ) );
  DFF \registers_reg[5][9]  ( .D(n3163), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][9] ) );
  DFF \registers_reg[5][8]  ( .D(n3162), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][8] ) );
  DFF \registers_reg[5][7]  ( .D(n3161), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][7] ) );
  DFF \registers_reg[5][6]  ( .D(n3160), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][6] ) );
  DFF \registers_reg[5][5]  ( .D(n3159), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][5] ) );
  DFF \registers_reg[5][4]  ( .D(n3158), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][4] ) );
  DFF \registers_reg[5][3]  ( .D(n3157), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][3] ) );
  DFF \registers_reg[5][2]  ( .D(n3156), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][2] ) );
  DFF \registers_reg[5][1]  ( .D(n3155), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][1] ) );
  DFF \registers_reg[5][0]  ( .D(n3154), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[5][0] ) );
  DFF \registers_reg[4][31]  ( .D(n3153), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][31] ) );
  DFF \registers_reg[4][30]  ( .D(n3152), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][30] ) );
  DFF \registers_reg[4][29]  ( .D(n3151), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][29] ) );
  DFF \registers_reg[4][28]  ( .D(n3150), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][28] ) );
  DFF \registers_reg[4][27]  ( .D(n3149), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][27] ) );
  DFF \registers_reg[4][26]  ( .D(n3148), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][26] ) );
  DFF \registers_reg[4][25]  ( .D(n3147), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][25] ) );
  DFF \registers_reg[4][24]  ( .D(n3146), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][24] ) );
  DFF \registers_reg[4][23]  ( .D(n3145), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][23] ) );
  DFF \registers_reg[4][22]  ( .D(n3144), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][22] ) );
  DFF \registers_reg[4][21]  ( .D(n3143), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][21] ) );
  DFF \registers_reg[4][20]  ( .D(n3142), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][20] ) );
  DFF \registers_reg[4][19]  ( .D(n3141), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][19] ) );
  DFF \registers_reg[4][18]  ( .D(n3140), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][18] ) );
  DFF \registers_reg[4][17]  ( .D(n3139), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][17] ) );
  DFF \registers_reg[4][16]  ( .D(n3138), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][16] ) );
  DFF \registers_reg[4][15]  ( .D(n3137), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][15] ) );
  DFF \registers_reg[4][14]  ( .D(n3136), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][14] ) );
  DFF \registers_reg[4][13]  ( .D(n3135), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][13] ) );
  DFF \registers_reg[4][12]  ( .D(n3134), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][12] ) );
  DFF \registers_reg[4][11]  ( .D(n3133), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][11] ) );
  DFF \registers_reg[4][10]  ( .D(n3132), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][10] ) );
  DFF \registers_reg[4][9]  ( .D(n3131), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][9] ) );
  DFF \registers_reg[4][8]  ( .D(n3130), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][8] ) );
  DFF \registers_reg[4][7]  ( .D(n3129), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][7] ) );
  DFF \registers_reg[4][6]  ( .D(n3128), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][6] ) );
  DFF \registers_reg[4][5]  ( .D(n3127), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][5] ) );
  DFF \registers_reg[4][4]  ( .D(n3126), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][4] ) );
  DFF \registers_reg[4][3]  ( .D(n3125), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][3] ) );
  DFF \registers_reg[4][2]  ( .D(n3124), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][2] ) );
  DFF \registers_reg[4][1]  ( .D(n3123), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][1] ) );
  DFF \registers_reg[4][0]  ( .D(n3122), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[4][0] ) );
  DFF \registers_reg[3][31]  ( .D(n3121), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][31] ) );
  DFF \registers_reg[3][30]  ( .D(n3120), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][30] ) );
  DFF \registers_reg[3][29]  ( .D(n3119), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][29] ) );
  DFF \registers_reg[3][28]  ( .D(n3118), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][28] ) );
  DFF \registers_reg[3][27]  ( .D(n3117), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][27] ) );
  DFF \registers_reg[3][26]  ( .D(n3116), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][26] ) );
  DFF \registers_reg[3][25]  ( .D(n3115), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][25] ) );
  DFF \registers_reg[3][24]  ( .D(n3114), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][24] ) );
  DFF \registers_reg[3][23]  ( .D(n3113), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][23] ) );
  DFF \registers_reg[3][22]  ( .D(n3112), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][22] ) );
  DFF \registers_reg[3][21]  ( .D(n3111), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][21] ) );
  DFF \registers_reg[3][20]  ( .D(n3110), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][20] ) );
  DFF \registers_reg[3][19]  ( .D(n3109), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][19] ) );
  DFF \registers_reg[3][18]  ( .D(n3108), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][18] ) );
  DFF \registers_reg[3][17]  ( .D(n3107), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][17] ) );
  DFF \registers_reg[3][16]  ( .D(n3106), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][16] ) );
  DFF \registers_reg[3][15]  ( .D(n3105), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][15] ) );
  DFF \registers_reg[3][14]  ( .D(n3104), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][14] ) );
  DFF \registers_reg[3][13]  ( .D(n3103), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][13] ) );
  DFF \registers_reg[3][12]  ( .D(n3102), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][12] ) );
  DFF \registers_reg[3][11]  ( .D(n3101), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][11] ) );
  DFF \registers_reg[3][10]  ( .D(n3100), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][10] ) );
  DFF \registers_reg[3][9]  ( .D(n3099), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][9] ) );
  DFF \registers_reg[3][8]  ( .D(n3098), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][8] ) );
  DFF \registers_reg[3][7]  ( .D(n3097), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][7] ) );
  DFF \registers_reg[3][6]  ( .D(n3096), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][6] ) );
  DFF \registers_reg[3][5]  ( .D(n3095), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][5] ) );
  DFF \registers_reg[3][4]  ( .D(n3094), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][4] ) );
  DFF \registers_reg[3][3]  ( .D(n3093), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][3] ) );
  DFF \registers_reg[3][2]  ( .D(n3092), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][2] ) );
  DFF \registers_reg[3][1]  ( .D(n3091), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][1] ) );
  DFF \registers_reg[3][0]  ( .D(n3090), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[3][0] ) );
  DFF \registers_reg[2][31]  ( .D(n3089), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][31] ) );
  DFF \registers_reg[2][30]  ( .D(n3088), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][30] ) );
  DFF \registers_reg[2][29]  ( .D(n3087), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][29] ) );
  DFF \registers_reg[2][28]  ( .D(n3086), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][28] ) );
  DFF \registers_reg[2][27]  ( .D(n3085), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][27] ) );
  DFF \registers_reg[2][26]  ( .D(n3084), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][26] ) );
  DFF \registers_reg[2][25]  ( .D(n3083), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][25] ) );
  DFF \registers_reg[2][24]  ( .D(n3082), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][24] ) );
  DFF \registers_reg[2][23]  ( .D(n3081), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][23] ) );
  DFF \registers_reg[2][22]  ( .D(n3080), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][22] ) );
  DFF \registers_reg[2][21]  ( .D(n3079), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][21] ) );
  DFF \registers_reg[2][20]  ( .D(n3078), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][20] ) );
  DFF \registers_reg[2][19]  ( .D(n3077), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][19] ) );
  DFF \registers_reg[2][18]  ( .D(n3076), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][18] ) );
  DFF \registers_reg[2][17]  ( .D(n3075), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][17] ) );
  DFF \registers_reg[2][16]  ( .D(n3074), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][16] ) );
  DFF \registers_reg[2][15]  ( .D(n3073), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][15] ) );
  DFF \registers_reg[2][14]  ( .D(n3072), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][14] ) );
  DFF \registers_reg[2][13]  ( .D(n3071), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][13] ) );
  DFF \registers_reg[2][12]  ( .D(n3070), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][12] ) );
  DFF \registers_reg[2][11]  ( .D(n3069), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][11] ) );
  DFF \registers_reg[2][10]  ( .D(n3068), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][10] ) );
  DFF \registers_reg[2][9]  ( .D(n3067), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][9] ) );
  DFF \registers_reg[2][8]  ( .D(n3066), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][8] ) );
  DFF \registers_reg[2][7]  ( .D(n3065), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][7] ) );
  DFF \registers_reg[2][6]  ( .D(n3064), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][6] ) );
  DFF \registers_reg[2][5]  ( .D(n3063), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][5] ) );
  DFF \registers_reg[2][4]  ( .D(n3062), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][4] ) );
  DFF \registers_reg[2][3]  ( .D(n3061), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][3] ) );
  DFF \registers_reg[2][2]  ( .D(n3060), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][2] ) );
  DFF \registers_reg[2][1]  ( .D(n3059), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][1] ) );
  DFF \registers_reg[2][0]  ( .D(n3058), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[2][0] ) );
  DFF \registers_reg[1][31]  ( .D(n3057), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][31] ) );
  DFF \registers_reg[1][30]  ( .D(n3056), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][30] ) );
  DFF \registers_reg[1][29]  ( .D(n3055), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][29] ) );
  DFF \registers_reg[1][28]  ( .D(n3054), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][28] ) );
  DFF \registers_reg[1][27]  ( .D(n3053), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][27] ) );
  DFF \registers_reg[1][26]  ( .D(n3052), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][26] ) );
  DFF \registers_reg[1][25]  ( .D(n3051), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][25] ) );
  DFF \registers_reg[1][24]  ( .D(n3050), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][24] ) );
  DFF \registers_reg[1][23]  ( .D(n3049), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][23] ) );
  DFF \registers_reg[1][22]  ( .D(n3048), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][22] ) );
  DFF \registers_reg[1][21]  ( .D(n3047), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][21] ) );
  DFF \registers_reg[1][20]  ( .D(n3046), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][20] ) );
  DFF \registers_reg[1][19]  ( .D(n3045), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][19] ) );
  DFF \registers_reg[1][18]  ( .D(n3044), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][18] ) );
  DFF \registers_reg[1][17]  ( .D(n3043), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][17] ) );
  DFF \registers_reg[1][16]  ( .D(n3042), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][16] ) );
  DFF \registers_reg[1][15]  ( .D(n3041), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][15] ) );
  DFF \registers_reg[1][14]  ( .D(n3040), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][14] ) );
  DFF \registers_reg[1][13]  ( .D(n3039), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][13] ) );
  DFF \registers_reg[1][12]  ( .D(n3038), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][12] ) );
  DFF \registers_reg[1][11]  ( .D(n3037), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][11] ) );
  DFF \registers_reg[1][10]  ( .D(n3036), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][10] ) );
  DFF \registers_reg[1][9]  ( .D(n3035), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][9] ) );
  DFF \registers_reg[1][8]  ( .D(n3034), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][8] ) );
  DFF \registers_reg[1][7]  ( .D(n3033), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][7] ) );
  DFF \registers_reg[1][6]  ( .D(n3032), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][6] ) );
  DFF \registers_reg[1][5]  ( .D(n3031), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][5] ) );
  DFF \registers_reg[1][4]  ( .D(n3030), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][4] ) );
  DFF \registers_reg[1][3]  ( .D(n3029), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][3] ) );
  DFF \registers_reg[1][2]  ( .D(n3028), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][2] ) );
  DFF \registers_reg[1][1]  ( .D(n3027), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][1] ) );
  DFF \registers_reg[1][0]  ( .D(n3026), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \registers[1][0] ) );
  MUX U4051 ( .IN0(\registers[30][0] ), .IN1(\registers[31][0] ), .SEL(N9), 
        .F(n4018) );
  MUX U4052 ( .IN0(\registers[28][0] ), .IN1(\registers[29][0] ), .SEL(N9), 
        .F(n4019) );
  MUX U4053 ( .IN0(n4019), .IN1(n4018), .SEL(N10), .F(n4020) );
  MUX U4054 ( .IN0(\registers[26][0] ), .IN1(\registers[27][0] ), .SEL(N9), 
        .F(n4021) );
  MUX U4055 ( .IN0(\registers[24][0] ), .IN1(\registers[25][0] ), .SEL(N9), 
        .F(n4022) );
  MUX U4056 ( .IN0(n4022), .IN1(n4021), .SEL(N10), .F(n4023) );
  MUX U4057 ( .IN0(n4023), .IN1(n4020), .SEL(N11), .F(n4024) );
  MUX U4058 ( .IN0(\registers[22][0] ), .IN1(\registers[23][0] ), .SEL(N9), 
        .F(n4025) );
  MUX U4059 ( .IN0(\registers[20][0] ), .IN1(\registers[21][0] ), .SEL(N9), 
        .F(n4026) );
  MUX U4060 ( .IN0(n4026), .IN1(n4025), .SEL(N10), .F(n4027) );
  MUX U4061 ( .IN0(\registers[18][0] ), .IN1(\registers[19][0] ), .SEL(N9), 
        .F(n4028) );
  MUX U4062 ( .IN0(\registers[16][0] ), .IN1(\registers[17][0] ), .SEL(N9), 
        .F(n4029) );
  MUX U4063 ( .IN0(n4029), .IN1(n4028), .SEL(N10), .F(n4030) );
  MUX U4064 ( .IN0(n4030), .IN1(n4027), .SEL(N11), .F(n4031) );
  MUX U4065 ( .IN0(n4031), .IN1(n4024), .SEL(N12), .F(n4032) );
  MUX U4066 ( .IN0(\registers[14][0] ), .IN1(\registers[15][0] ), .SEL(N9), 
        .F(n4033) );
  MUX U4067 ( .IN0(\registers[12][0] ), .IN1(\registers[13][0] ), .SEL(N9), 
        .F(n4034) );
  MUX U4068 ( .IN0(n4034), .IN1(n4033), .SEL(N10), .F(n4035) );
  MUX U4069 ( .IN0(\registers[10][0] ), .IN1(\registers[11][0] ), .SEL(N9), 
        .F(n4036) );
  MUX U4070 ( .IN0(\registers[8][0] ), .IN1(\registers[9][0] ), .SEL(N9), .F(
        n4037) );
  MUX U4071 ( .IN0(n4037), .IN1(n4036), .SEL(N10), .F(n4038) );
  MUX U4072 ( .IN0(n4038), .IN1(n4035), .SEL(N11), .F(n4039) );
  MUX U4073 ( .IN0(\registers[6][0] ), .IN1(\registers[7][0] ), .SEL(N9), .F(
        n4040) );
  MUX U4074 ( .IN0(\registers[4][0] ), .IN1(\registers[5][0] ), .SEL(N9), .F(
        n4041) );
  MUX U4075 ( .IN0(n4041), .IN1(n4040), .SEL(N10), .F(n4042) );
  MUX U4076 ( .IN0(\registers[2][0] ), .IN1(\registers[3][0] ), .SEL(N9), .F(
        n4043) );
  MUX U4078 ( .IN0(n4044), .IN1(n4043), .SEL(N10), .F(n4045) );
  MUX U4079 ( .IN0(n4045), .IN1(n4042), .SEL(N11), .F(n4046) );
  MUX U4080 ( .IN0(n4046), .IN1(n4039), .SEL(N12), .F(n4047) );
  MUX U4081 ( .IN0(n4047), .IN1(n4032), .SEL(N13), .F(reg_source_out[0]) );
  MUX U4082 ( .IN0(\registers[30][1] ), .IN1(\registers[31][1] ), .SEL(N9), 
        .F(n4048) );
  MUX U4083 ( .IN0(\registers[28][1] ), .IN1(\registers[29][1] ), .SEL(N9), 
        .F(n4049) );
  MUX U4084 ( .IN0(n4049), .IN1(n4048), .SEL(N10), .F(n4050) );
  MUX U4085 ( .IN0(\registers[26][1] ), .IN1(\registers[27][1] ), .SEL(N9), 
        .F(n4051) );
  MUX U4086 ( .IN0(\registers[24][1] ), .IN1(\registers[25][1] ), .SEL(N9), 
        .F(n4052) );
  MUX U4087 ( .IN0(n4052), .IN1(n4051), .SEL(N10), .F(n4053) );
  MUX U4088 ( .IN0(n4053), .IN1(n4050), .SEL(N11), .F(n4054) );
  MUX U4089 ( .IN0(\registers[22][1] ), .IN1(\registers[23][1] ), .SEL(N9), 
        .F(n4055) );
  MUX U4090 ( .IN0(\registers[20][1] ), .IN1(\registers[21][1] ), .SEL(N9), 
        .F(n4056) );
  MUX U4091 ( .IN0(n4056), .IN1(n4055), .SEL(N10), .F(n4057) );
  MUX U4092 ( .IN0(\registers[18][1] ), .IN1(\registers[19][1] ), .SEL(N9), 
        .F(n4058) );
  MUX U4093 ( .IN0(\registers[16][1] ), .IN1(\registers[17][1] ), .SEL(N9), 
        .F(n4059) );
  MUX U4094 ( .IN0(n4059), .IN1(n4058), .SEL(N10), .F(n4060) );
  MUX U4095 ( .IN0(n4060), .IN1(n4057), .SEL(N11), .F(n4061) );
  MUX U4096 ( .IN0(n4061), .IN1(n4054), .SEL(N12), .F(n4062) );
  MUX U4097 ( .IN0(\registers[14][1] ), .IN1(\registers[15][1] ), .SEL(N9), 
        .F(n4063) );
  MUX U4098 ( .IN0(\registers[12][1] ), .IN1(\registers[13][1] ), .SEL(N9), 
        .F(n4064) );
  MUX U4099 ( .IN0(n4064), .IN1(n4063), .SEL(N10), .F(n4065) );
  MUX U4100 ( .IN0(\registers[10][1] ), .IN1(\registers[11][1] ), .SEL(N9), 
        .F(n4066) );
  MUX U4101 ( .IN0(\registers[8][1] ), .IN1(\registers[9][1] ), .SEL(N9), .F(
        n4067) );
  MUX U4102 ( .IN0(n4067), .IN1(n4066), .SEL(N10), .F(n4068) );
  MUX U4103 ( .IN0(n4068), .IN1(n4065), .SEL(N11), .F(n4069) );
  MUX U4104 ( .IN0(\registers[6][1] ), .IN1(\registers[7][1] ), .SEL(N9), .F(
        n4070) );
  MUX U4105 ( .IN0(\registers[4][1] ), .IN1(\registers[5][1] ), .SEL(N9), .F(
        n4071) );
  MUX U4106 ( .IN0(n4071), .IN1(n4070), .SEL(N10), .F(n4072) );
  MUX U4107 ( .IN0(\registers[2][1] ), .IN1(\registers[3][1] ), .SEL(N9), .F(
        n4073) );
  MUX U4109 ( .IN0(n4074), .IN1(n4073), .SEL(N10), .F(n4075) );
  MUX U4110 ( .IN0(n4075), .IN1(n4072), .SEL(N11), .F(n4076) );
  MUX U4111 ( .IN0(n4076), .IN1(n4069), .SEL(N12), .F(n4077) );
  MUX U4112 ( .IN0(n4077), .IN1(n4062), .SEL(N13), .F(reg_source_out[1]) );
  MUX U4113 ( .IN0(\registers[30][2] ), .IN1(\registers[31][2] ), .SEL(N9), 
        .F(n4078) );
  MUX U4114 ( .IN0(\registers[28][2] ), .IN1(\registers[29][2] ), .SEL(N9), 
        .F(n4079) );
  MUX U4115 ( .IN0(n4079), .IN1(n4078), .SEL(N10), .F(n4080) );
  MUX U4116 ( .IN0(\registers[26][2] ), .IN1(\registers[27][2] ), .SEL(N9), 
        .F(n4081) );
  MUX U4117 ( .IN0(\registers[24][2] ), .IN1(\registers[25][2] ), .SEL(N9), 
        .F(n4082) );
  MUX U4118 ( .IN0(n4082), .IN1(n4081), .SEL(N10), .F(n4083) );
  MUX U4119 ( .IN0(n4083), .IN1(n4080), .SEL(N11), .F(n4084) );
  MUX U4120 ( .IN0(\registers[22][2] ), .IN1(\registers[23][2] ), .SEL(N9), 
        .F(n4085) );
  MUX U4121 ( .IN0(\registers[20][2] ), .IN1(\registers[21][2] ), .SEL(N9), 
        .F(n4086) );
  MUX U4122 ( .IN0(n4086), .IN1(n4085), .SEL(N10), .F(n4087) );
  MUX U4123 ( .IN0(\registers[18][2] ), .IN1(\registers[19][2] ), .SEL(N9), 
        .F(n4088) );
  MUX U4124 ( .IN0(\registers[16][2] ), .IN1(\registers[17][2] ), .SEL(N9), 
        .F(n4089) );
  MUX U4125 ( .IN0(n4089), .IN1(n4088), .SEL(N10), .F(n4090) );
  MUX U4126 ( .IN0(n4090), .IN1(n4087), .SEL(N11), .F(n4091) );
  MUX U4127 ( .IN0(n4091), .IN1(n4084), .SEL(N12), .F(n4092) );
  MUX U4128 ( .IN0(\registers[14][2] ), .IN1(\registers[15][2] ), .SEL(N9), 
        .F(n4093) );
  MUX U4129 ( .IN0(\registers[12][2] ), .IN1(\registers[13][2] ), .SEL(N9), 
        .F(n4094) );
  MUX U4130 ( .IN0(n4094), .IN1(n4093), .SEL(N10), .F(n4095) );
  MUX U4131 ( .IN0(\registers[10][2] ), .IN1(\registers[11][2] ), .SEL(N9), 
        .F(n4096) );
  MUX U4132 ( .IN0(\registers[8][2] ), .IN1(\registers[9][2] ), .SEL(N9), .F(
        n4097) );
  MUX U4133 ( .IN0(n4097), .IN1(n4096), .SEL(N10), .F(n4098) );
  MUX U4134 ( .IN0(n4098), .IN1(n4095), .SEL(N11), .F(n4099) );
  MUX U4135 ( .IN0(\registers[6][2] ), .IN1(\registers[7][2] ), .SEL(N9), .F(
        n4100) );
  MUX U4136 ( .IN0(\registers[4][2] ), .IN1(\registers[5][2] ), .SEL(N9), .F(
        n4101) );
  MUX U4137 ( .IN0(n4101), .IN1(n4100), .SEL(N10), .F(n4102) );
  MUX U4138 ( .IN0(\registers[2][2] ), .IN1(\registers[3][2] ), .SEL(N9), .F(
        n4103) );
  MUX U4140 ( .IN0(n4104), .IN1(n4103), .SEL(N10), .F(n4105) );
  MUX U4141 ( .IN0(n4105), .IN1(n4102), .SEL(N11), .F(n4106) );
  MUX U4142 ( .IN0(n4106), .IN1(n4099), .SEL(N12), .F(n4107) );
  MUX U4143 ( .IN0(n4107), .IN1(n4092), .SEL(N13), .F(reg_source_out[2]) );
  MUX U4144 ( .IN0(\registers[30][3] ), .IN1(\registers[31][3] ), .SEL(N9), 
        .F(n4108) );
  MUX U4145 ( .IN0(\registers[28][3] ), .IN1(\registers[29][3] ), .SEL(N9), 
        .F(n4109) );
  MUX U4146 ( .IN0(n4109), .IN1(n4108), .SEL(N10), .F(n4110) );
  MUX U4147 ( .IN0(\registers[26][3] ), .IN1(\registers[27][3] ), .SEL(N9), 
        .F(n4111) );
  MUX U4148 ( .IN0(\registers[24][3] ), .IN1(\registers[25][3] ), .SEL(N9), 
        .F(n4112) );
  MUX U4149 ( .IN0(n4112), .IN1(n4111), .SEL(N10), .F(n4113) );
  MUX U4150 ( .IN0(n4113), .IN1(n4110), .SEL(N11), .F(n4114) );
  MUX U4151 ( .IN0(\registers[22][3] ), .IN1(\registers[23][3] ), .SEL(N9), 
        .F(n4115) );
  MUX U4152 ( .IN0(\registers[20][3] ), .IN1(\registers[21][3] ), .SEL(N9), 
        .F(n4116) );
  MUX U4153 ( .IN0(n4116), .IN1(n4115), .SEL(N10), .F(n4117) );
  MUX U4154 ( .IN0(\registers[18][3] ), .IN1(\registers[19][3] ), .SEL(N9), 
        .F(n4118) );
  MUX U4155 ( .IN0(\registers[16][3] ), .IN1(\registers[17][3] ), .SEL(N9), 
        .F(n4119) );
  MUX U4156 ( .IN0(n4119), .IN1(n4118), .SEL(N10), .F(n4120) );
  MUX U4157 ( .IN0(n4120), .IN1(n4117), .SEL(N11), .F(n4121) );
  MUX U4158 ( .IN0(n4121), .IN1(n4114), .SEL(N12), .F(n4122) );
  MUX U4159 ( .IN0(\registers[14][3] ), .IN1(\registers[15][3] ), .SEL(N9), 
        .F(n4123) );
  MUX U4160 ( .IN0(\registers[12][3] ), .IN1(\registers[13][3] ), .SEL(N9), 
        .F(n4124) );
  MUX U4161 ( .IN0(n4124), .IN1(n4123), .SEL(N10), .F(n4125) );
  MUX U4162 ( .IN0(\registers[10][3] ), .IN1(\registers[11][3] ), .SEL(N9), 
        .F(n4126) );
  MUX U4163 ( .IN0(\registers[8][3] ), .IN1(\registers[9][3] ), .SEL(N9), .F(
        n4127) );
  MUX U4164 ( .IN0(n4127), .IN1(n4126), .SEL(N10), .F(n4128) );
  MUX U4165 ( .IN0(n4128), .IN1(n4125), .SEL(N11), .F(n4129) );
  MUX U4166 ( .IN0(\registers[6][3] ), .IN1(\registers[7][3] ), .SEL(N9), .F(
        n4130) );
  MUX U4167 ( .IN0(\registers[4][3] ), .IN1(\registers[5][3] ), .SEL(N9), .F(
        n4131) );
  MUX U4168 ( .IN0(n4131), .IN1(n4130), .SEL(N10), .F(n4132) );
  MUX U4169 ( .IN0(\registers[2][3] ), .IN1(\registers[3][3] ), .SEL(N9), .F(
        n4133) );
  MUX U4171 ( .IN0(n4134), .IN1(n4133), .SEL(N10), .F(n4135) );
  MUX U4172 ( .IN0(n4135), .IN1(n4132), .SEL(N11), .F(n4136) );
  MUX U4173 ( .IN0(n4136), .IN1(n4129), .SEL(N12), .F(n4137) );
  MUX U4174 ( .IN0(n4137), .IN1(n4122), .SEL(N13), .F(reg_source_out[3]) );
  MUX U4175 ( .IN0(\registers[30][4] ), .IN1(\registers[31][4] ), .SEL(N9), 
        .F(n4138) );
  MUX U4176 ( .IN0(\registers[28][4] ), .IN1(\registers[29][4] ), .SEL(N9), 
        .F(n4139) );
  MUX U4177 ( .IN0(n4139), .IN1(n4138), .SEL(N10), .F(n4140) );
  MUX U4178 ( .IN0(\registers[26][4] ), .IN1(\registers[27][4] ), .SEL(N9), 
        .F(n4141) );
  MUX U4179 ( .IN0(\registers[24][4] ), .IN1(\registers[25][4] ), .SEL(N9), 
        .F(n4142) );
  MUX U4180 ( .IN0(n4142), .IN1(n4141), .SEL(N10), .F(n4143) );
  MUX U4181 ( .IN0(n4143), .IN1(n4140), .SEL(N11), .F(n4144) );
  MUX U4182 ( .IN0(\registers[22][4] ), .IN1(\registers[23][4] ), .SEL(N9), 
        .F(n4145) );
  MUX U4183 ( .IN0(\registers[20][4] ), .IN1(\registers[21][4] ), .SEL(N9), 
        .F(n4146) );
  MUX U4184 ( .IN0(n4146), .IN1(n4145), .SEL(N10), .F(n4147) );
  MUX U4185 ( .IN0(\registers[18][4] ), .IN1(\registers[19][4] ), .SEL(N9), 
        .F(n4148) );
  MUX U4186 ( .IN0(\registers[16][4] ), .IN1(\registers[17][4] ), .SEL(N9), 
        .F(n4149) );
  MUX U4187 ( .IN0(n4149), .IN1(n4148), .SEL(N10), .F(n4150) );
  MUX U4188 ( .IN0(n4150), .IN1(n4147), .SEL(N11), .F(n4151) );
  MUX U4189 ( .IN0(n4151), .IN1(n4144), .SEL(N12), .F(n4152) );
  MUX U4190 ( .IN0(\registers[14][4] ), .IN1(\registers[15][4] ), .SEL(N9), 
        .F(n4153) );
  MUX U4191 ( .IN0(\registers[12][4] ), .IN1(\registers[13][4] ), .SEL(N9), 
        .F(n4154) );
  MUX U4192 ( .IN0(n4154), .IN1(n4153), .SEL(N10), .F(n4155) );
  MUX U4193 ( .IN0(\registers[10][4] ), .IN1(\registers[11][4] ), .SEL(N9), 
        .F(n4156) );
  MUX U4194 ( .IN0(\registers[8][4] ), .IN1(\registers[9][4] ), .SEL(N9), .F(
        n4157) );
  MUX U4195 ( .IN0(n4157), .IN1(n4156), .SEL(N10), .F(n4158) );
  MUX U4196 ( .IN0(n4158), .IN1(n4155), .SEL(N11), .F(n4159) );
  MUX U4197 ( .IN0(\registers[6][4] ), .IN1(\registers[7][4] ), .SEL(N9), .F(
        n4160) );
  MUX U4198 ( .IN0(\registers[4][4] ), .IN1(\registers[5][4] ), .SEL(N9), .F(
        n4161) );
  MUX U4199 ( .IN0(n4161), .IN1(n4160), .SEL(N10), .F(n4162) );
  MUX U4200 ( .IN0(\registers[2][4] ), .IN1(\registers[3][4] ), .SEL(N9), .F(
        n4163) );
  MUX U4202 ( .IN0(n4164), .IN1(n4163), .SEL(N10), .F(n4165) );
  MUX U4203 ( .IN0(n4165), .IN1(n4162), .SEL(N11), .F(n4166) );
  MUX U4204 ( .IN0(n4166), .IN1(n4159), .SEL(N12), .F(n4167) );
  MUX U4205 ( .IN0(n4167), .IN1(n4152), .SEL(N13), .F(reg_source_out[4]) );
  MUX U4206 ( .IN0(\registers[30][5] ), .IN1(\registers[31][5] ), .SEL(N9), 
        .F(n4168) );
  MUX U4207 ( .IN0(\registers[28][5] ), .IN1(\registers[29][5] ), .SEL(N9), 
        .F(n4169) );
  MUX U4208 ( .IN0(n4169), .IN1(n4168), .SEL(N10), .F(n4170) );
  MUX U4209 ( .IN0(\registers[26][5] ), .IN1(\registers[27][5] ), .SEL(N9), 
        .F(n4171) );
  MUX U4210 ( .IN0(\registers[24][5] ), .IN1(\registers[25][5] ), .SEL(N9), 
        .F(n4172) );
  MUX U4211 ( .IN0(n4172), .IN1(n4171), .SEL(N10), .F(n4173) );
  MUX U4212 ( .IN0(n4173), .IN1(n4170), .SEL(N11), .F(n4174) );
  MUX U4213 ( .IN0(\registers[22][5] ), .IN1(\registers[23][5] ), .SEL(N9), 
        .F(n4175) );
  MUX U4214 ( .IN0(\registers[20][5] ), .IN1(\registers[21][5] ), .SEL(N9), 
        .F(n4176) );
  MUX U4215 ( .IN0(n4176), .IN1(n4175), .SEL(N10), .F(n4177) );
  MUX U4216 ( .IN0(\registers[18][5] ), .IN1(\registers[19][5] ), .SEL(N9), 
        .F(n4178) );
  MUX U4217 ( .IN0(\registers[16][5] ), .IN1(\registers[17][5] ), .SEL(N9), 
        .F(n4179) );
  MUX U4218 ( .IN0(n4179), .IN1(n4178), .SEL(N10), .F(n4180) );
  MUX U4219 ( .IN0(n4180), .IN1(n4177), .SEL(N11), .F(n4181) );
  MUX U4220 ( .IN0(n4181), .IN1(n4174), .SEL(N12), .F(n4182) );
  MUX U4221 ( .IN0(\registers[14][5] ), .IN1(\registers[15][5] ), .SEL(N9), 
        .F(n4183) );
  MUX U4222 ( .IN0(\registers[12][5] ), .IN1(\registers[13][5] ), .SEL(N9), 
        .F(n4184) );
  MUX U4223 ( .IN0(n4184), .IN1(n4183), .SEL(N10), .F(n4185) );
  MUX U4224 ( .IN0(\registers[10][5] ), .IN1(\registers[11][5] ), .SEL(N9), 
        .F(n4186) );
  MUX U4225 ( .IN0(\registers[8][5] ), .IN1(\registers[9][5] ), .SEL(N9), .F(
        n4187) );
  MUX U4226 ( .IN0(n4187), .IN1(n4186), .SEL(N10), .F(n4188) );
  MUX U4227 ( .IN0(n4188), .IN1(n4185), .SEL(N11), .F(n4189) );
  MUX U4228 ( .IN0(\registers[6][5] ), .IN1(\registers[7][5] ), .SEL(N9), .F(
        n4190) );
  MUX U4229 ( .IN0(\registers[4][5] ), .IN1(\registers[5][5] ), .SEL(N9), .F(
        n4191) );
  MUX U4230 ( .IN0(n4191), .IN1(n4190), .SEL(N10), .F(n4192) );
  MUX U4231 ( .IN0(\registers[2][5] ), .IN1(\registers[3][5] ), .SEL(N9), .F(
        n4193) );
  MUX U4233 ( .IN0(n4194), .IN1(n4193), .SEL(N10), .F(n4195) );
  MUX U4234 ( .IN0(n4195), .IN1(n4192), .SEL(N11), .F(n4196) );
  MUX U4235 ( .IN0(n4196), .IN1(n4189), .SEL(N12), .F(n4197) );
  MUX U4236 ( .IN0(n4197), .IN1(n4182), .SEL(N13), .F(reg_source_out[5]) );
  MUX U4237 ( .IN0(\registers[30][6] ), .IN1(\registers[31][6] ), .SEL(N9), 
        .F(n4198) );
  MUX U4238 ( .IN0(\registers[28][6] ), .IN1(\registers[29][6] ), .SEL(N9), 
        .F(n4199) );
  MUX U4239 ( .IN0(n4199), .IN1(n4198), .SEL(N10), .F(n4200) );
  MUX U4240 ( .IN0(\registers[26][6] ), .IN1(\registers[27][6] ), .SEL(N9), 
        .F(n4201) );
  MUX U4241 ( .IN0(\registers[24][6] ), .IN1(\registers[25][6] ), .SEL(N9), 
        .F(n4202) );
  MUX U4242 ( .IN0(n4202), .IN1(n4201), .SEL(N10), .F(n4203) );
  MUX U4243 ( .IN0(n4203), .IN1(n4200), .SEL(N11), .F(n4204) );
  MUX U4244 ( .IN0(\registers[22][6] ), .IN1(\registers[23][6] ), .SEL(N9), 
        .F(n4205) );
  MUX U4245 ( .IN0(\registers[20][6] ), .IN1(\registers[21][6] ), .SEL(N9), 
        .F(n4206) );
  MUX U4246 ( .IN0(n4206), .IN1(n4205), .SEL(N10), .F(n4207) );
  MUX U4247 ( .IN0(\registers[18][6] ), .IN1(\registers[19][6] ), .SEL(N9), 
        .F(n4208) );
  MUX U4248 ( .IN0(\registers[16][6] ), .IN1(\registers[17][6] ), .SEL(N9), 
        .F(n4209) );
  MUX U4249 ( .IN0(n4209), .IN1(n4208), .SEL(N10), .F(n4210) );
  MUX U4250 ( .IN0(n4210), .IN1(n4207), .SEL(N11), .F(n4211) );
  MUX U4251 ( .IN0(n4211), .IN1(n4204), .SEL(N12), .F(n4212) );
  MUX U4252 ( .IN0(\registers[14][6] ), .IN1(\registers[15][6] ), .SEL(N9), 
        .F(n4213) );
  MUX U4253 ( .IN0(\registers[12][6] ), .IN1(\registers[13][6] ), .SEL(N9), 
        .F(n4214) );
  MUX U4254 ( .IN0(n4214), .IN1(n4213), .SEL(N10), .F(n4215) );
  MUX U4255 ( .IN0(\registers[10][6] ), .IN1(\registers[11][6] ), .SEL(N9), 
        .F(n4216) );
  MUX U4256 ( .IN0(\registers[8][6] ), .IN1(\registers[9][6] ), .SEL(N9), .F(
        n4217) );
  MUX U4257 ( .IN0(n4217), .IN1(n4216), .SEL(N10), .F(n4218) );
  MUX U4258 ( .IN0(n4218), .IN1(n4215), .SEL(N11), .F(n4219) );
  MUX U4259 ( .IN0(\registers[6][6] ), .IN1(\registers[7][6] ), .SEL(N9), .F(
        n4220) );
  MUX U4260 ( .IN0(\registers[4][6] ), .IN1(\registers[5][6] ), .SEL(N9), .F(
        n4221) );
  MUX U4261 ( .IN0(n4221), .IN1(n4220), .SEL(N10), .F(n4222) );
  MUX U4262 ( .IN0(\registers[2][6] ), .IN1(\registers[3][6] ), .SEL(N9), .F(
        n4223) );
  MUX U4264 ( .IN0(n4224), .IN1(n4223), .SEL(N10), .F(n4225) );
  MUX U4265 ( .IN0(n4225), .IN1(n4222), .SEL(N11), .F(n4226) );
  MUX U4266 ( .IN0(n4226), .IN1(n4219), .SEL(N12), .F(n4227) );
  MUX U4267 ( .IN0(n4227), .IN1(n4212), .SEL(N13), .F(reg_source_out[6]) );
  MUX U4268 ( .IN0(\registers[30][7] ), .IN1(\registers[31][7] ), .SEL(N9), 
        .F(n4228) );
  MUX U4269 ( .IN0(\registers[28][7] ), .IN1(\registers[29][7] ), .SEL(N9), 
        .F(n4229) );
  MUX U4270 ( .IN0(n4229), .IN1(n4228), .SEL(N10), .F(n4230) );
  MUX U4271 ( .IN0(\registers[26][7] ), .IN1(\registers[27][7] ), .SEL(N9), 
        .F(n4231) );
  MUX U4272 ( .IN0(\registers[24][7] ), .IN1(\registers[25][7] ), .SEL(N9), 
        .F(n4232) );
  MUX U4273 ( .IN0(n4232), .IN1(n4231), .SEL(N10), .F(n4233) );
  MUX U4274 ( .IN0(n4233), .IN1(n4230), .SEL(N11), .F(n4234) );
  MUX U4275 ( .IN0(\registers[22][7] ), .IN1(\registers[23][7] ), .SEL(N9), 
        .F(n4235) );
  MUX U4276 ( .IN0(\registers[20][7] ), .IN1(\registers[21][7] ), .SEL(N9), 
        .F(n4236) );
  MUX U4277 ( .IN0(n4236), .IN1(n4235), .SEL(N10), .F(n4237) );
  MUX U4278 ( .IN0(\registers[18][7] ), .IN1(\registers[19][7] ), .SEL(N9), 
        .F(n4238) );
  MUX U4279 ( .IN0(\registers[16][7] ), .IN1(\registers[17][7] ), .SEL(N9), 
        .F(n4239) );
  MUX U4280 ( .IN0(n4239), .IN1(n4238), .SEL(N10), .F(n4240) );
  MUX U4281 ( .IN0(n4240), .IN1(n4237), .SEL(N11), .F(n4241) );
  MUX U4282 ( .IN0(n4241), .IN1(n4234), .SEL(N12), .F(n4242) );
  MUX U4283 ( .IN0(\registers[14][7] ), .IN1(\registers[15][7] ), .SEL(N9), 
        .F(n4243) );
  MUX U4284 ( .IN0(\registers[12][7] ), .IN1(\registers[13][7] ), .SEL(N9), 
        .F(n4244) );
  MUX U4285 ( .IN0(n4244), .IN1(n4243), .SEL(N10), .F(n4245) );
  MUX U4286 ( .IN0(\registers[10][7] ), .IN1(\registers[11][7] ), .SEL(N9), 
        .F(n4246) );
  MUX U4287 ( .IN0(\registers[8][7] ), .IN1(\registers[9][7] ), .SEL(N9), .F(
        n4247) );
  MUX U4288 ( .IN0(n4247), .IN1(n4246), .SEL(N10), .F(n4248) );
  MUX U4289 ( .IN0(n4248), .IN1(n4245), .SEL(N11), .F(n4249) );
  MUX U4290 ( .IN0(\registers[6][7] ), .IN1(\registers[7][7] ), .SEL(N9), .F(
        n4250) );
  MUX U4291 ( .IN0(\registers[4][7] ), .IN1(\registers[5][7] ), .SEL(N9), .F(
        n4251) );
  MUX U4292 ( .IN0(n4251), .IN1(n4250), .SEL(N10), .F(n4252) );
  MUX U4293 ( .IN0(\registers[2][7] ), .IN1(\registers[3][7] ), .SEL(N9), .F(
        n4253) );
  MUX U4295 ( .IN0(n4254), .IN1(n4253), .SEL(N10), .F(n4255) );
  MUX U4296 ( .IN0(n4255), .IN1(n4252), .SEL(N11), .F(n4256) );
  MUX U4297 ( .IN0(n4256), .IN1(n4249), .SEL(N12), .F(n4257) );
  MUX U4298 ( .IN0(n4257), .IN1(n4242), .SEL(N13), .F(reg_source_out[7]) );
  MUX U4299 ( .IN0(\registers[30][8] ), .IN1(\registers[31][8] ), .SEL(N9), 
        .F(n4258) );
  MUX U4300 ( .IN0(\registers[28][8] ), .IN1(\registers[29][8] ), .SEL(N9), 
        .F(n4259) );
  MUX U4301 ( .IN0(n4259), .IN1(n4258), .SEL(N10), .F(n4260) );
  MUX U4302 ( .IN0(\registers[26][8] ), .IN1(\registers[27][8] ), .SEL(N9), 
        .F(n4261) );
  MUX U4303 ( .IN0(\registers[24][8] ), .IN1(\registers[25][8] ), .SEL(N9), 
        .F(n4262) );
  MUX U4304 ( .IN0(n4262), .IN1(n4261), .SEL(N10), .F(n4263) );
  MUX U4305 ( .IN0(n4263), .IN1(n4260), .SEL(N11), .F(n4264) );
  MUX U4306 ( .IN0(\registers[22][8] ), .IN1(\registers[23][8] ), .SEL(N9), 
        .F(n4265) );
  MUX U4307 ( .IN0(\registers[20][8] ), .IN1(\registers[21][8] ), .SEL(N9), 
        .F(n4266) );
  MUX U4308 ( .IN0(n4266), .IN1(n4265), .SEL(N10), .F(n4267) );
  MUX U4309 ( .IN0(\registers[18][8] ), .IN1(\registers[19][8] ), .SEL(N9), 
        .F(n4268) );
  MUX U4310 ( .IN0(\registers[16][8] ), .IN1(\registers[17][8] ), .SEL(N9), 
        .F(n4269) );
  MUX U4311 ( .IN0(n4269), .IN1(n4268), .SEL(N10), .F(n4270) );
  MUX U4312 ( .IN0(n4270), .IN1(n4267), .SEL(N11), .F(n4271) );
  MUX U4313 ( .IN0(n4271), .IN1(n4264), .SEL(N12), .F(n4272) );
  MUX U4314 ( .IN0(\registers[14][8] ), .IN1(\registers[15][8] ), .SEL(N9), 
        .F(n4273) );
  MUX U4315 ( .IN0(\registers[12][8] ), .IN1(\registers[13][8] ), .SEL(N9), 
        .F(n4274) );
  MUX U4316 ( .IN0(n4274), .IN1(n4273), .SEL(N10), .F(n4275) );
  MUX U4317 ( .IN0(\registers[10][8] ), .IN1(\registers[11][8] ), .SEL(N9), 
        .F(n4276) );
  MUX U4318 ( .IN0(\registers[8][8] ), .IN1(\registers[9][8] ), .SEL(N9), .F(
        n4277) );
  MUX U4319 ( .IN0(n4277), .IN1(n4276), .SEL(N10), .F(n4278) );
  MUX U4320 ( .IN0(n4278), .IN1(n4275), .SEL(N11), .F(n4279) );
  MUX U4321 ( .IN0(\registers[6][8] ), .IN1(\registers[7][8] ), .SEL(N9), .F(
        n4280) );
  MUX U4322 ( .IN0(\registers[4][8] ), .IN1(\registers[5][8] ), .SEL(N9), .F(
        n4281) );
  MUX U4323 ( .IN0(n4281), .IN1(n4280), .SEL(N10), .F(n4282) );
  MUX U4324 ( .IN0(\registers[2][8] ), .IN1(\registers[3][8] ), .SEL(N9), .F(
        n4283) );
  MUX U4326 ( .IN0(n4284), .IN1(n4283), .SEL(N10), .F(n4285) );
  MUX U4327 ( .IN0(n4285), .IN1(n4282), .SEL(N11), .F(n4286) );
  MUX U4328 ( .IN0(n4286), .IN1(n4279), .SEL(N12), .F(n4287) );
  MUX U4329 ( .IN0(n4287), .IN1(n4272), .SEL(N13), .F(reg_source_out[8]) );
  MUX U4330 ( .IN0(\registers[30][9] ), .IN1(\registers[31][9] ), .SEL(N9), 
        .F(n4288) );
  MUX U4331 ( .IN0(\registers[28][9] ), .IN1(\registers[29][9] ), .SEL(N9), 
        .F(n4289) );
  MUX U4332 ( .IN0(n4289), .IN1(n4288), .SEL(N10), .F(n4290) );
  MUX U4333 ( .IN0(\registers[26][9] ), .IN1(\registers[27][9] ), .SEL(N9), 
        .F(n4291) );
  MUX U4334 ( .IN0(\registers[24][9] ), .IN1(\registers[25][9] ), .SEL(N9), 
        .F(n4292) );
  MUX U4335 ( .IN0(n4292), .IN1(n4291), .SEL(N10), .F(n4293) );
  MUX U4336 ( .IN0(n4293), .IN1(n4290), .SEL(N11), .F(n4294) );
  MUX U4337 ( .IN0(\registers[22][9] ), .IN1(\registers[23][9] ), .SEL(N9), 
        .F(n4295) );
  MUX U4338 ( .IN0(\registers[20][9] ), .IN1(\registers[21][9] ), .SEL(N9), 
        .F(n4296) );
  MUX U4339 ( .IN0(n4296), .IN1(n4295), .SEL(N10), .F(n4297) );
  MUX U4340 ( .IN0(\registers[18][9] ), .IN1(\registers[19][9] ), .SEL(N9), 
        .F(n4298) );
  MUX U4341 ( .IN0(\registers[16][9] ), .IN1(\registers[17][9] ), .SEL(N9), 
        .F(n4299) );
  MUX U4342 ( .IN0(n4299), .IN1(n4298), .SEL(N10), .F(n4300) );
  MUX U4343 ( .IN0(n4300), .IN1(n4297), .SEL(N11), .F(n4301) );
  MUX U4344 ( .IN0(n4301), .IN1(n4294), .SEL(N12), .F(n4302) );
  MUX U4345 ( .IN0(\registers[14][9] ), .IN1(\registers[15][9] ), .SEL(N9), 
        .F(n4303) );
  MUX U4346 ( .IN0(\registers[12][9] ), .IN1(\registers[13][9] ), .SEL(N9), 
        .F(n4304) );
  MUX U4347 ( .IN0(n4304), .IN1(n4303), .SEL(N10), .F(n4305) );
  MUX U4348 ( .IN0(\registers[10][9] ), .IN1(\registers[11][9] ), .SEL(N9), 
        .F(n4306) );
  MUX U4349 ( .IN0(\registers[8][9] ), .IN1(\registers[9][9] ), .SEL(N9), .F(
        n4307) );
  MUX U4350 ( .IN0(n4307), .IN1(n4306), .SEL(N10), .F(n4308) );
  MUX U4351 ( .IN0(n4308), .IN1(n4305), .SEL(N11), .F(n4309) );
  MUX U4352 ( .IN0(\registers[6][9] ), .IN1(\registers[7][9] ), .SEL(N9), .F(
        n4310) );
  MUX U4353 ( .IN0(\registers[4][9] ), .IN1(\registers[5][9] ), .SEL(N9), .F(
        n4311) );
  MUX U4354 ( .IN0(n4311), .IN1(n4310), .SEL(N10), .F(n4312) );
  MUX U4355 ( .IN0(\registers[2][9] ), .IN1(\registers[3][9] ), .SEL(N9), .F(
        n4313) );
  MUX U4357 ( .IN0(n4314), .IN1(n4313), .SEL(N10), .F(n4315) );
  MUX U4358 ( .IN0(n4315), .IN1(n4312), .SEL(N11), .F(n4316) );
  MUX U4359 ( .IN0(n4316), .IN1(n4309), .SEL(N12), .F(n4317) );
  MUX U4360 ( .IN0(n4317), .IN1(n4302), .SEL(N13), .F(reg_source_out[9]) );
  MUX U4361 ( .IN0(\registers[30][10] ), .IN1(\registers[31][10] ), .SEL(N9), 
        .F(n4318) );
  MUX U4362 ( .IN0(\registers[28][10] ), .IN1(\registers[29][10] ), .SEL(N9), 
        .F(n4319) );
  MUX U4363 ( .IN0(n4319), .IN1(n4318), .SEL(N10), .F(n4320) );
  MUX U4364 ( .IN0(\registers[26][10] ), .IN1(\registers[27][10] ), .SEL(N9), 
        .F(n4321) );
  MUX U4365 ( .IN0(\registers[24][10] ), .IN1(\registers[25][10] ), .SEL(N9), 
        .F(n4322) );
  MUX U4366 ( .IN0(n4322), .IN1(n4321), .SEL(N10), .F(n4323) );
  MUX U4367 ( .IN0(n4323), .IN1(n4320), .SEL(N11), .F(n4324) );
  MUX U4368 ( .IN0(\registers[22][10] ), .IN1(\registers[23][10] ), .SEL(N9), 
        .F(n4325) );
  MUX U4369 ( .IN0(\registers[20][10] ), .IN1(\registers[21][10] ), .SEL(N9), 
        .F(n4326) );
  MUX U4370 ( .IN0(n4326), .IN1(n4325), .SEL(N10), .F(n4327) );
  MUX U4371 ( .IN0(\registers[18][10] ), .IN1(\registers[19][10] ), .SEL(N9), 
        .F(n4328) );
  MUX U4372 ( .IN0(\registers[16][10] ), .IN1(\registers[17][10] ), .SEL(N9), 
        .F(n4329) );
  MUX U4373 ( .IN0(n4329), .IN1(n4328), .SEL(N10), .F(n4330) );
  MUX U4374 ( .IN0(n4330), .IN1(n4327), .SEL(N11), .F(n4331) );
  MUX U4375 ( .IN0(n4331), .IN1(n4324), .SEL(N12), .F(n4332) );
  MUX U4376 ( .IN0(\registers[14][10] ), .IN1(\registers[15][10] ), .SEL(N9), 
        .F(n4333) );
  MUX U4377 ( .IN0(\registers[12][10] ), .IN1(\registers[13][10] ), .SEL(N9), 
        .F(n4334) );
  MUX U4378 ( .IN0(n4334), .IN1(n4333), .SEL(N10), .F(n4335) );
  MUX U4379 ( .IN0(\registers[10][10] ), .IN1(\registers[11][10] ), .SEL(N9), 
        .F(n4336) );
  MUX U4380 ( .IN0(\registers[8][10] ), .IN1(\registers[9][10] ), .SEL(N9), 
        .F(n4337) );
  MUX U4381 ( .IN0(n4337), .IN1(n4336), .SEL(N10), .F(n4338) );
  MUX U4382 ( .IN0(n4338), .IN1(n4335), .SEL(N11), .F(n4339) );
  MUX U4383 ( .IN0(\registers[6][10] ), .IN1(\registers[7][10] ), .SEL(N9), 
        .F(n4340) );
  MUX U4384 ( .IN0(\registers[4][10] ), .IN1(\registers[5][10] ), .SEL(N9), 
        .F(n4341) );
  MUX U4385 ( .IN0(n4341), .IN1(n4340), .SEL(N10), .F(n4342) );
  MUX U4386 ( .IN0(\registers[2][10] ), .IN1(\registers[3][10] ), .SEL(N9), 
        .F(n4343) );
  MUX U4388 ( .IN0(n4344), .IN1(n4343), .SEL(N10), .F(n4345) );
  MUX U4389 ( .IN0(n4345), .IN1(n4342), .SEL(N11), .F(n4346) );
  MUX U4390 ( .IN0(n4346), .IN1(n4339), .SEL(N12), .F(n4347) );
  MUX U4391 ( .IN0(n4347), .IN1(n4332), .SEL(N13), .F(reg_source_out[10]) );
  MUX U4392 ( .IN0(\registers[30][11] ), .IN1(\registers[31][11] ), .SEL(N9), 
        .F(n4348) );
  MUX U4393 ( .IN0(\registers[28][11] ), .IN1(\registers[29][11] ), .SEL(N9), 
        .F(n4349) );
  MUX U4394 ( .IN0(n4349), .IN1(n4348), .SEL(N10), .F(n4350) );
  MUX U4395 ( .IN0(\registers[26][11] ), .IN1(\registers[27][11] ), .SEL(N9), 
        .F(n4351) );
  MUX U4396 ( .IN0(\registers[24][11] ), .IN1(\registers[25][11] ), .SEL(N9), 
        .F(n4352) );
  MUX U4397 ( .IN0(n4352), .IN1(n4351), .SEL(N10), .F(n4353) );
  MUX U4398 ( .IN0(n4353), .IN1(n4350), .SEL(N11), .F(n4354) );
  MUX U4399 ( .IN0(\registers[22][11] ), .IN1(\registers[23][11] ), .SEL(N9), 
        .F(n4355) );
  MUX U4400 ( .IN0(\registers[20][11] ), .IN1(\registers[21][11] ), .SEL(N9), 
        .F(n4356) );
  MUX U4401 ( .IN0(n4356), .IN1(n4355), .SEL(N10), .F(n4357) );
  MUX U4402 ( .IN0(\registers[18][11] ), .IN1(\registers[19][11] ), .SEL(N9), 
        .F(n4358) );
  MUX U4403 ( .IN0(\registers[16][11] ), .IN1(\registers[17][11] ), .SEL(N9), 
        .F(n4359) );
  MUX U4404 ( .IN0(n4359), .IN1(n4358), .SEL(N10), .F(n4360) );
  MUX U4405 ( .IN0(n4360), .IN1(n4357), .SEL(N11), .F(n4361) );
  MUX U4406 ( .IN0(n4361), .IN1(n4354), .SEL(N12), .F(n4362) );
  MUX U4407 ( .IN0(\registers[14][11] ), .IN1(\registers[15][11] ), .SEL(N9), 
        .F(n4363) );
  MUX U4408 ( .IN0(\registers[12][11] ), .IN1(\registers[13][11] ), .SEL(N9), 
        .F(n4364) );
  MUX U4409 ( .IN0(n4364), .IN1(n4363), .SEL(N10), .F(n4365) );
  MUX U4410 ( .IN0(\registers[10][11] ), .IN1(\registers[11][11] ), .SEL(N9), 
        .F(n4366) );
  MUX U4411 ( .IN0(\registers[8][11] ), .IN1(\registers[9][11] ), .SEL(N9), 
        .F(n4367) );
  MUX U4412 ( .IN0(n4367), .IN1(n4366), .SEL(N10), .F(n4368) );
  MUX U4413 ( .IN0(n4368), .IN1(n4365), .SEL(N11), .F(n4369) );
  MUX U4414 ( .IN0(\registers[6][11] ), .IN1(\registers[7][11] ), .SEL(N9), 
        .F(n4370) );
  MUX U4415 ( .IN0(\registers[4][11] ), .IN1(\registers[5][11] ), .SEL(N9), 
        .F(n4371) );
  MUX U4416 ( .IN0(n4371), .IN1(n4370), .SEL(N10), .F(n4372) );
  MUX U4417 ( .IN0(\registers[2][11] ), .IN1(\registers[3][11] ), .SEL(N9), 
        .F(n4373) );
  MUX U4419 ( .IN0(n4374), .IN1(n4373), .SEL(N10), .F(n4375) );
  MUX U4420 ( .IN0(n4375), .IN1(n4372), .SEL(N11), .F(n4376) );
  MUX U4421 ( .IN0(n4376), .IN1(n4369), .SEL(N12), .F(n4377) );
  MUX U4422 ( .IN0(n4377), .IN1(n4362), .SEL(N13), .F(reg_source_out[11]) );
  MUX U4423 ( .IN0(\registers[30][12] ), .IN1(\registers[31][12] ), .SEL(N9), 
        .F(n4378) );
  MUX U4424 ( .IN0(\registers[28][12] ), .IN1(\registers[29][12] ), .SEL(N9), 
        .F(n4379) );
  MUX U4425 ( .IN0(n4379), .IN1(n4378), .SEL(N10), .F(n4380) );
  MUX U4426 ( .IN0(\registers[26][12] ), .IN1(\registers[27][12] ), .SEL(N9), 
        .F(n4381) );
  MUX U4427 ( .IN0(\registers[24][12] ), .IN1(\registers[25][12] ), .SEL(N9), 
        .F(n4382) );
  MUX U4428 ( .IN0(n4382), .IN1(n4381), .SEL(N10), .F(n4383) );
  MUX U4429 ( .IN0(n4383), .IN1(n4380), .SEL(N11), .F(n4384) );
  MUX U4430 ( .IN0(\registers[22][12] ), .IN1(\registers[23][12] ), .SEL(N9), 
        .F(n4385) );
  MUX U4431 ( .IN0(\registers[20][12] ), .IN1(\registers[21][12] ), .SEL(N9), 
        .F(n4386) );
  MUX U4432 ( .IN0(n4386), .IN1(n4385), .SEL(N10), .F(n4387) );
  MUX U4433 ( .IN0(\registers[18][12] ), .IN1(\registers[19][12] ), .SEL(N9), 
        .F(n4388) );
  MUX U4434 ( .IN0(\registers[16][12] ), .IN1(\registers[17][12] ), .SEL(N9), 
        .F(n4389) );
  MUX U4435 ( .IN0(n4389), .IN1(n4388), .SEL(N10), .F(n4390) );
  MUX U4436 ( .IN0(n4390), .IN1(n4387), .SEL(N11), .F(n4391) );
  MUX U4437 ( .IN0(n4391), .IN1(n4384), .SEL(N12), .F(n4392) );
  MUX U4438 ( .IN0(\registers[14][12] ), .IN1(\registers[15][12] ), .SEL(N9), 
        .F(n4393) );
  MUX U4439 ( .IN0(\registers[12][12] ), .IN1(\registers[13][12] ), .SEL(N9), 
        .F(n4394) );
  MUX U4440 ( .IN0(n4394), .IN1(n4393), .SEL(N10), .F(n4395) );
  MUX U4441 ( .IN0(\registers[10][12] ), .IN1(\registers[11][12] ), .SEL(N9), 
        .F(n4396) );
  MUX U4442 ( .IN0(\registers[8][12] ), .IN1(\registers[9][12] ), .SEL(N9), 
        .F(n4397) );
  MUX U4443 ( .IN0(n4397), .IN1(n4396), .SEL(N10), .F(n4398) );
  MUX U4444 ( .IN0(n4398), .IN1(n4395), .SEL(N11), .F(n4399) );
  MUX U4445 ( .IN0(\registers[6][12] ), .IN1(\registers[7][12] ), .SEL(N9), 
        .F(n4400) );
  MUX U4446 ( .IN0(\registers[4][12] ), .IN1(\registers[5][12] ), .SEL(N9), 
        .F(n4401) );
  MUX U4447 ( .IN0(n4401), .IN1(n4400), .SEL(N10), .F(n4402) );
  MUX U4448 ( .IN0(\registers[2][12] ), .IN1(\registers[3][12] ), .SEL(N9), 
        .F(n4403) );
  MUX U4450 ( .IN0(n4404), .IN1(n4403), .SEL(N10), .F(n4405) );
  MUX U4451 ( .IN0(n4405), .IN1(n4402), .SEL(N11), .F(n4406) );
  MUX U4452 ( .IN0(n4406), .IN1(n4399), .SEL(N12), .F(n4407) );
  MUX U4453 ( .IN0(n4407), .IN1(n4392), .SEL(N13), .F(reg_source_out[12]) );
  MUX U4454 ( .IN0(\registers[30][13] ), .IN1(\registers[31][13] ), .SEL(N9), 
        .F(n4408) );
  MUX U4455 ( .IN0(\registers[28][13] ), .IN1(\registers[29][13] ), .SEL(N9), 
        .F(n4409) );
  MUX U4456 ( .IN0(n4409), .IN1(n4408), .SEL(N10), .F(n4410) );
  MUX U4457 ( .IN0(\registers[26][13] ), .IN1(\registers[27][13] ), .SEL(N9), 
        .F(n4411) );
  MUX U4458 ( .IN0(\registers[24][13] ), .IN1(\registers[25][13] ), .SEL(N9), 
        .F(n4412) );
  MUX U4459 ( .IN0(n4412), .IN1(n4411), .SEL(N10), .F(n4413) );
  MUX U4460 ( .IN0(n4413), .IN1(n4410), .SEL(N11), .F(n4414) );
  MUX U4461 ( .IN0(\registers[22][13] ), .IN1(\registers[23][13] ), .SEL(N9), 
        .F(n4415) );
  MUX U4462 ( .IN0(\registers[20][13] ), .IN1(\registers[21][13] ), .SEL(N9), 
        .F(n4416) );
  MUX U4463 ( .IN0(n4416), .IN1(n4415), .SEL(N10), .F(n4417) );
  MUX U4464 ( .IN0(\registers[18][13] ), .IN1(\registers[19][13] ), .SEL(N9), 
        .F(n4418) );
  MUX U4465 ( .IN0(\registers[16][13] ), .IN1(\registers[17][13] ), .SEL(N9), 
        .F(n4419) );
  MUX U4466 ( .IN0(n4419), .IN1(n4418), .SEL(N10), .F(n4420) );
  MUX U4467 ( .IN0(n4420), .IN1(n4417), .SEL(N11), .F(n4421) );
  MUX U4468 ( .IN0(n4421), .IN1(n4414), .SEL(N12), .F(n4422) );
  MUX U4469 ( .IN0(\registers[14][13] ), .IN1(\registers[15][13] ), .SEL(N9), 
        .F(n4423) );
  MUX U4470 ( .IN0(\registers[12][13] ), .IN1(\registers[13][13] ), .SEL(N9), 
        .F(n4424) );
  MUX U4471 ( .IN0(n4424), .IN1(n4423), .SEL(N10), .F(n4425) );
  MUX U4472 ( .IN0(\registers[10][13] ), .IN1(\registers[11][13] ), .SEL(N9), 
        .F(n4426) );
  MUX U4473 ( .IN0(\registers[8][13] ), .IN1(\registers[9][13] ), .SEL(N9), 
        .F(n4427) );
  MUX U4474 ( .IN0(n4427), .IN1(n4426), .SEL(N10), .F(n4428) );
  MUX U4475 ( .IN0(n4428), .IN1(n4425), .SEL(N11), .F(n4429) );
  MUX U4476 ( .IN0(\registers[6][13] ), .IN1(\registers[7][13] ), .SEL(N9), 
        .F(n4430) );
  MUX U4477 ( .IN0(\registers[4][13] ), .IN1(\registers[5][13] ), .SEL(N9), 
        .F(n4431) );
  MUX U4478 ( .IN0(n4431), .IN1(n4430), .SEL(N10), .F(n4432) );
  MUX U4479 ( .IN0(\registers[2][13] ), .IN1(\registers[3][13] ), .SEL(N9), 
        .F(n4433) );
  MUX U4481 ( .IN0(n4434), .IN1(n4433), .SEL(N10), .F(n4435) );
  MUX U4482 ( .IN0(n4435), .IN1(n4432), .SEL(N11), .F(n4436) );
  MUX U4483 ( .IN0(n4436), .IN1(n4429), .SEL(N12), .F(n4437) );
  MUX U4484 ( .IN0(n4437), .IN1(n4422), .SEL(N13), .F(reg_source_out[13]) );
  MUX U4485 ( .IN0(\registers[30][14] ), .IN1(\registers[31][14] ), .SEL(N9), 
        .F(n4438) );
  MUX U4486 ( .IN0(\registers[28][14] ), .IN1(\registers[29][14] ), .SEL(N9), 
        .F(n4439) );
  MUX U4487 ( .IN0(n4439), .IN1(n4438), .SEL(N10), .F(n4440) );
  MUX U4488 ( .IN0(\registers[26][14] ), .IN1(\registers[27][14] ), .SEL(N9), 
        .F(n4441) );
  MUX U4489 ( .IN0(\registers[24][14] ), .IN1(\registers[25][14] ), .SEL(N9), 
        .F(n4442) );
  MUX U4490 ( .IN0(n4442), .IN1(n4441), .SEL(N10), .F(n4443) );
  MUX U4491 ( .IN0(n4443), .IN1(n4440), .SEL(N11), .F(n4444) );
  MUX U4492 ( .IN0(\registers[22][14] ), .IN1(\registers[23][14] ), .SEL(N9), 
        .F(n4445) );
  MUX U4493 ( .IN0(\registers[20][14] ), .IN1(\registers[21][14] ), .SEL(N9), 
        .F(n4446) );
  MUX U4494 ( .IN0(n4446), .IN1(n4445), .SEL(N10), .F(n4447) );
  MUX U4495 ( .IN0(\registers[18][14] ), .IN1(\registers[19][14] ), .SEL(N9), 
        .F(n4448) );
  MUX U4496 ( .IN0(\registers[16][14] ), .IN1(\registers[17][14] ), .SEL(N9), 
        .F(n4449) );
  MUX U4497 ( .IN0(n4449), .IN1(n4448), .SEL(N10), .F(n4450) );
  MUX U4498 ( .IN0(n4450), .IN1(n4447), .SEL(N11), .F(n4451) );
  MUX U4499 ( .IN0(n4451), .IN1(n4444), .SEL(N12), .F(n4452) );
  MUX U4500 ( .IN0(\registers[14][14] ), .IN1(\registers[15][14] ), .SEL(N9), 
        .F(n4453) );
  MUX U4501 ( .IN0(\registers[12][14] ), .IN1(\registers[13][14] ), .SEL(N9), 
        .F(n4454) );
  MUX U4502 ( .IN0(n4454), .IN1(n4453), .SEL(N10), .F(n4455) );
  MUX U4503 ( .IN0(\registers[10][14] ), .IN1(\registers[11][14] ), .SEL(N9), 
        .F(n4456) );
  MUX U4504 ( .IN0(\registers[8][14] ), .IN1(\registers[9][14] ), .SEL(N9), 
        .F(n4457) );
  MUX U4505 ( .IN0(n4457), .IN1(n4456), .SEL(N10), .F(n4458) );
  MUX U4506 ( .IN0(n4458), .IN1(n4455), .SEL(N11), .F(n4459) );
  MUX U4507 ( .IN0(\registers[6][14] ), .IN1(\registers[7][14] ), .SEL(N9), 
        .F(n4460) );
  MUX U4508 ( .IN0(\registers[4][14] ), .IN1(\registers[5][14] ), .SEL(N9), 
        .F(n4461) );
  MUX U4509 ( .IN0(n4461), .IN1(n4460), .SEL(N10), .F(n4462) );
  MUX U4510 ( .IN0(\registers[2][14] ), .IN1(\registers[3][14] ), .SEL(N9), 
        .F(n4463) );
  MUX U4512 ( .IN0(n4464), .IN1(n4463), .SEL(N10), .F(n4465) );
  MUX U4513 ( .IN0(n4465), .IN1(n4462), .SEL(N11), .F(n4466) );
  MUX U4514 ( .IN0(n4466), .IN1(n4459), .SEL(N12), .F(n4467) );
  MUX U4515 ( .IN0(n4467), .IN1(n4452), .SEL(N13), .F(reg_source_out[14]) );
  MUX U4516 ( .IN0(\registers[30][15] ), .IN1(\registers[31][15] ), .SEL(N9), 
        .F(n4468) );
  MUX U4517 ( .IN0(\registers[28][15] ), .IN1(\registers[29][15] ), .SEL(N9), 
        .F(n4469) );
  MUX U4518 ( .IN0(n4469), .IN1(n4468), .SEL(N10), .F(n4470) );
  MUX U4519 ( .IN0(\registers[26][15] ), .IN1(\registers[27][15] ), .SEL(N9), 
        .F(n4471) );
  MUX U4520 ( .IN0(\registers[24][15] ), .IN1(\registers[25][15] ), .SEL(N9), 
        .F(n4472) );
  MUX U4521 ( .IN0(n4472), .IN1(n4471), .SEL(N10), .F(n4473) );
  MUX U4522 ( .IN0(n4473), .IN1(n4470), .SEL(N11), .F(n4474) );
  MUX U4523 ( .IN0(\registers[22][15] ), .IN1(\registers[23][15] ), .SEL(N9), 
        .F(n4475) );
  MUX U4524 ( .IN0(\registers[20][15] ), .IN1(\registers[21][15] ), .SEL(N9), 
        .F(n4476) );
  MUX U4525 ( .IN0(n4476), .IN1(n4475), .SEL(N10), .F(n4477) );
  MUX U4526 ( .IN0(\registers[18][15] ), .IN1(\registers[19][15] ), .SEL(N9), 
        .F(n4478) );
  MUX U4527 ( .IN0(\registers[16][15] ), .IN1(\registers[17][15] ), .SEL(N9), 
        .F(n4479) );
  MUX U4528 ( .IN0(n4479), .IN1(n4478), .SEL(N10), .F(n4480) );
  MUX U4529 ( .IN0(n4480), .IN1(n4477), .SEL(N11), .F(n4481) );
  MUX U4530 ( .IN0(n4481), .IN1(n4474), .SEL(N12), .F(n4482) );
  MUX U4531 ( .IN0(\registers[14][15] ), .IN1(\registers[15][15] ), .SEL(N9), 
        .F(n4483) );
  MUX U4532 ( .IN0(\registers[12][15] ), .IN1(\registers[13][15] ), .SEL(N9), 
        .F(n4484) );
  MUX U4533 ( .IN0(n4484), .IN1(n4483), .SEL(N10), .F(n4485) );
  MUX U4534 ( .IN0(\registers[10][15] ), .IN1(\registers[11][15] ), .SEL(N9), 
        .F(n4486) );
  MUX U4535 ( .IN0(\registers[8][15] ), .IN1(\registers[9][15] ), .SEL(N9), 
        .F(n4487) );
  MUX U4536 ( .IN0(n4487), .IN1(n4486), .SEL(N10), .F(n4488) );
  MUX U4537 ( .IN0(n4488), .IN1(n4485), .SEL(N11), .F(n4489) );
  MUX U4538 ( .IN0(\registers[6][15] ), .IN1(\registers[7][15] ), .SEL(N9), 
        .F(n4490) );
  MUX U4539 ( .IN0(\registers[4][15] ), .IN1(\registers[5][15] ), .SEL(N9), 
        .F(n4491) );
  MUX U4540 ( .IN0(n4491), .IN1(n4490), .SEL(N10), .F(n4492) );
  MUX U4541 ( .IN0(\registers[2][15] ), .IN1(\registers[3][15] ), .SEL(N9), 
        .F(n4493) );
  MUX U4543 ( .IN0(n4494), .IN1(n4493), .SEL(N10), .F(n4495) );
  MUX U4544 ( .IN0(n4495), .IN1(n4492), .SEL(N11), .F(n4496) );
  MUX U4545 ( .IN0(n4496), .IN1(n4489), .SEL(N12), .F(n4497) );
  MUX U4546 ( .IN0(n4497), .IN1(n4482), .SEL(N13), .F(reg_source_out[15]) );
  MUX U4547 ( .IN0(\registers[30][16] ), .IN1(\registers[31][16] ), .SEL(N9), 
        .F(n4498) );
  MUX U4548 ( .IN0(\registers[28][16] ), .IN1(\registers[29][16] ), .SEL(N9), 
        .F(n4499) );
  MUX U4549 ( .IN0(n4499), .IN1(n4498), .SEL(N10), .F(n4500) );
  MUX U4550 ( .IN0(\registers[26][16] ), .IN1(\registers[27][16] ), .SEL(N9), 
        .F(n4501) );
  MUX U4551 ( .IN0(\registers[24][16] ), .IN1(\registers[25][16] ), .SEL(N9), 
        .F(n4502) );
  MUX U4552 ( .IN0(n4502), .IN1(n4501), .SEL(N10), .F(n4503) );
  MUX U4553 ( .IN0(n4503), .IN1(n4500), .SEL(N11), .F(n4504) );
  MUX U4554 ( .IN0(\registers[22][16] ), .IN1(\registers[23][16] ), .SEL(N9), 
        .F(n4505) );
  MUX U4555 ( .IN0(\registers[20][16] ), .IN1(\registers[21][16] ), .SEL(N9), 
        .F(n4506) );
  MUX U4556 ( .IN0(n4506), .IN1(n4505), .SEL(N10), .F(n4507) );
  MUX U4557 ( .IN0(\registers[18][16] ), .IN1(\registers[19][16] ), .SEL(N9), 
        .F(n4508) );
  MUX U4558 ( .IN0(\registers[16][16] ), .IN1(\registers[17][16] ), .SEL(N9), 
        .F(n4509) );
  MUX U4559 ( .IN0(n4509), .IN1(n4508), .SEL(N10), .F(n4510) );
  MUX U4560 ( .IN0(n4510), .IN1(n4507), .SEL(N11), .F(n4511) );
  MUX U4561 ( .IN0(n4511), .IN1(n4504), .SEL(N12), .F(n4512) );
  MUX U4562 ( .IN0(\registers[14][16] ), .IN1(\registers[15][16] ), .SEL(N9), 
        .F(n4513) );
  MUX U4563 ( .IN0(\registers[12][16] ), .IN1(\registers[13][16] ), .SEL(N9), 
        .F(n4514) );
  MUX U4564 ( .IN0(n4514), .IN1(n4513), .SEL(N10), .F(n4515) );
  MUX U4565 ( .IN0(\registers[10][16] ), .IN1(\registers[11][16] ), .SEL(N9), 
        .F(n4516) );
  MUX U4566 ( .IN0(\registers[8][16] ), .IN1(\registers[9][16] ), .SEL(N9), 
        .F(n4517) );
  MUX U4567 ( .IN0(n4517), .IN1(n4516), .SEL(N10), .F(n4518) );
  MUX U4568 ( .IN0(n4518), .IN1(n4515), .SEL(N11), .F(n4519) );
  MUX U4569 ( .IN0(\registers[6][16] ), .IN1(\registers[7][16] ), .SEL(N9), 
        .F(n4520) );
  MUX U4570 ( .IN0(\registers[4][16] ), .IN1(\registers[5][16] ), .SEL(N9), 
        .F(n4521) );
  MUX U4571 ( .IN0(n4521), .IN1(n4520), .SEL(N10), .F(n4522) );
  MUX U4572 ( .IN0(\registers[2][16] ), .IN1(\registers[3][16] ), .SEL(N9), 
        .F(n4523) );
  MUX U4574 ( .IN0(n4524), .IN1(n4523), .SEL(N10), .F(n4525) );
  MUX U4575 ( .IN0(n4525), .IN1(n4522), .SEL(N11), .F(n4526) );
  MUX U4576 ( .IN0(n4526), .IN1(n4519), .SEL(N12), .F(n4527) );
  MUX U4577 ( .IN0(n4527), .IN1(n4512), .SEL(N13), .F(reg_source_out[16]) );
  MUX U4578 ( .IN0(\registers[30][17] ), .IN1(\registers[31][17] ), .SEL(N9), 
        .F(n4528) );
  MUX U4579 ( .IN0(\registers[28][17] ), .IN1(\registers[29][17] ), .SEL(N9), 
        .F(n4529) );
  MUX U4580 ( .IN0(n4529), .IN1(n4528), .SEL(N10), .F(n4530) );
  MUX U4581 ( .IN0(\registers[26][17] ), .IN1(\registers[27][17] ), .SEL(N9), 
        .F(n4531) );
  MUX U4582 ( .IN0(\registers[24][17] ), .IN1(\registers[25][17] ), .SEL(N9), 
        .F(n4532) );
  MUX U4583 ( .IN0(n4532), .IN1(n4531), .SEL(N10), .F(n4533) );
  MUX U4584 ( .IN0(n4533), .IN1(n4530), .SEL(N11), .F(n4534) );
  MUX U4585 ( .IN0(\registers[22][17] ), .IN1(\registers[23][17] ), .SEL(N9), 
        .F(n4535) );
  MUX U4586 ( .IN0(\registers[20][17] ), .IN1(\registers[21][17] ), .SEL(N9), 
        .F(n4536) );
  MUX U4587 ( .IN0(n4536), .IN1(n4535), .SEL(N10), .F(n4537) );
  MUX U4588 ( .IN0(\registers[18][17] ), .IN1(\registers[19][17] ), .SEL(N9), 
        .F(n4538) );
  MUX U4589 ( .IN0(\registers[16][17] ), .IN1(\registers[17][17] ), .SEL(N9), 
        .F(n4539) );
  MUX U4590 ( .IN0(n4539), .IN1(n4538), .SEL(N10), .F(n4540) );
  MUX U4591 ( .IN0(n4540), .IN1(n4537), .SEL(N11), .F(n4541) );
  MUX U4592 ( .IN0(n4541), .IN1(n4534), .SEL(N12), .F(n4542) );
  MUX U4593 ( .IN0(\registers[14][17] ), .IN1(\registers[15][17] ), .SEL(N9), 
        .F(n4543) );
  MUX U4594 ( .IN0(\registers[12][17] ), .IN1(\registers[13][17] ), .SEL(N9), 
        .F(n4544) );
  MUX U4595 ( .IN0(n4544), .IN1(n4543), .SEL(N10), .F(n4545) );
  MUX U4596 ( .IN0(\registers[10][17] ), .IN1(\registers[11][17] ), .SEL(N9), 
        .F(n4546) );
  MUX U4597 ( .IN0(\registers[8][17] ), .IN1(\registers[9][17] ), .SEL(N9), 
        .F(n4547) );
  MUX U4598 ( .IN0(n4547), .IN1(n4546), .SEL(N10), .F(n4548) );
  MUX U4599 ( .IN0(n4548), .IN1(n4545), .SEL(N11), .F(n4549) );
  MUX U4600 ( .IN0(\registers[6][17] ), .IN1(\registers[7][17] ), .SEL(N9), 
        .F(n4550) );
  MUX U4601 ( .IN0(\registers[4][17] ), .IN1(\registers[5][17] ), .SEL(N9), 
        .F(n4551) );
  MUX U4602 ( .IN0(n4551), .IN1(n4550), .SEL(N10), .F(n4552) );
  MUX U4603 ( .IN0(\registers[2][17] ), .IN1(\registers[3][17] ), .SEL(N9), 
        .F(n4553) );
  MUX U4605 ( .IN0(n4554), .IN1(n4553), .SEL(N10), .F(n4555) );
  MUX U4606 ( .IN0(n4555), .IN1(n4552), .SEL(N11), .F(n4556) );
  MUX U4607 ( .IN0(n4556), .IN1(n4549), .SEL(N12), .F(n4557) );
  MUX U4608 ( .IN0(n4557), .IN1(n4542), .SEL(N13), .F(reg_source_out[17]) );
  MUX U4609 ( .IN0(\registers[30][18] ), .IN1(\registers[31][18] ), .SEL(N9), 
        .F(n4558) );
  MUX U4610 ( .IN0(\registers[28][18] ), .IN1(\registers[29][18] ), .SEL(N9), 
        .F(n4559) );
  MUX U4611 ( .IN0(n4559), .IN1(n4558), .SEL(N10), .F(n4560) );
  MUX U4612 ( .IN0(\registers[26][18] ), .IN1(\registers[27][18] ), .SEL(N9), 
        .F(n4561) );
  MUX U4613 ( .IN0(\registers[24][18] ), .IN1(\registers[25][18] ), .SEL(N9), 
        .F(n4562) );
  MUX U4614 ( .IN0(n4562), .IN1(n4561), .SEL(N10), .F(n4563) );
  MUX U4615 ( .IN0(n4563), .IN1(n4560), .SEL(N11), .F(n4564) );
  MUX U4616 ( .IN0(\registers[22][18] ), .IN1(\registers[23][18] ), .SEL(N9), 
        .F(n4565) );
  MUX U4617 ( .IN0(\registers[20][18] ), .IN1(\registers[21][18] ), .SEL(N9), 
        .F(n4566) );
  MUX U4618 ( .IN0(n4566), .IN1(n4565), .SEL(N10), .F(n4567) );
  MUX U4619 ( .IN0(\registers[18][18] ), .IN1(\registers[19][18] ), .SEL(N9), 
        .F(n4568) );
  MUX U4620 ( .IN0(\registers[16][18] ), .IN1(\registers[17][18] ), .SEL(N9), 
        .F(n4569) );
  MUX U4621 ( .IN0(n4569), .IN1(n4568), .SEL(N10), .F(n4570) );
  MUX U4622 ( .IN0(n4570), .IN1(n4567), .SEL(N11), .F(n4571) );
  MUX U4623 ( .IN0(n4571), .IN1(n4564), .SEL(N12), .F(n4572) );
  MUX U4624 ( .IN0(\registers[14][18] ), .IN1(\registers[15][18] ), .SEL(N9), 
        .F(n4573) );
  MUX U4625 ( .IN0(\registers[12][18] ), .IN1(\registers[13][18] ), .SEL(N9), 
        .F(n4574) );
  MUX U4626 ( .IN0(n4574), .IN1(n4573), .SEL(N10), .F(n4575) );
  MUX U4627 ( .IN0(\registers[10][18] ), .IN1(\registers[11][18] ), .SEL(N9), 
        .F(n4576) );
  MUX U4628 ( .IN0(\registers[8][18] ), .IN1(\registers[9][18] ), .SEL(N9), 
        .F(n4577) );
  MUX U4629 ( .IN0(n4577), .IN1(n4576), .SEL(N10), .F(n4578) );
  MUX U4630 ( .IN0(n4578), .IN1(n4575), .SEL(N11), .F(n4579) );
  MUX U4631 ( .IN0(\registers[6][18] ), .IN1(\registers[7][18] ), .SEL(N9), 
        .F(n4580) );
  MUX U4632 ( .IN0(\registers[4][18] ), .IN1(\registers[5][18] ), .SEL(N9), 
        .F(n4581) );
  MUX U4633 ( .IN0(n4581), .IN1(n4580), .SEL(N10), .F(n4582) );
  MUX U4634 ( .IN0(\registers[2][18] ), .IN1(\registers[3][18] ), .SEL(N9), 
        .F(n4583) );
  MUX U4636 ( .IN0(n4584), .IN1(n4583), .SEL(N10), .F(n4585) );
  MUX U4637 ( .IN0(n4585), .IN1(n4582), .SEL(N11), .F(n4586) );
  MUX U4638 ( .IN0(n4586), .IN1(n4579), .SEL(N12), .F(n4587) );
  MUX U4639 ( .IN0(n4587), .IN1(n4572), .SEL(N13), .F(reg_source_out[18]) );
  MUX U4640 ( .IN0(\registers[30][19] ), .IN1(\registers[31][19] ), .SEL(N9), 
        .F(n4588) );
  MUX U4641 ( .IN0(\registers[28][19] ), .IN1(\registers[29][19] ), .SEL(N9), 
        .F(n4589) );
  MUX U4642 ( .IN0(n4589), .IN1(n4588), .SEL(N10), .F(n4590) );
  MUX U4643 ( .IN0(\registers[26][19] ), .IN1(\registers[27][19] ), .SEL(N9), 
        .F(n4591) );
  MUX U4644 ( .IN0(\registers[24][19] ), .IN1(\registers[25][19] ), .SEL(N9), 
        .F(n4592) );
  MUX U4645 ( .IN0(n4592), .IN1(n4591), .SEL(N10), .F(n4593) );
  MUX U4646 ( .IN0(n4593), .IN1(n4590), .SEL(N11), .F(n4594) );
  MUX U4647 ( .IN0(\registers[22][19] ), .IN1(\registers[23][19] ), .SEL(N9), 
        .F(n4595) );
  MUX U4648 ( .IN0(\registers[20][19] ), .IN1(\registers[21][19] ), .SEL(N9), 
        .F(n4596) );
  MUX U4649 ( .IN0(n4596), .IN1(n4595), .SEL(N10), .F(n4597) );
  MUX U4650 ( .IN0(\registers[18][19] ), .IN1(\registers[19][19] ), .SEL(N9), 
        .F(n4598) );
  MUX U4651 ( .IN0(\registers[16][19] ), .IN1(\registers[17][19] ), .SEL(N9), 
        .F(n4599) );
  MUX U4652 ( .IN0(n4599), .IN1(n4598), .SEL(N10), .F(n4600) );
  MUX U4653 ( .IN0(n4600), .IN1(n4597), .SEL(N11), .F(n4601) );
  MUX U4654 ( .IN0(n4601), .IN1(n4594), .SEL(N12), .F(n4602) );
  MUX U4655 ( .IN0(\registers[14][19] ), .IN1(\registers[15][19] ), .SEL(N9), 
        .F(n4603) );
  MUX U4656 ( .IN0(\registers[12][19] ), .IN1(\registers[13][19] ), .SEL(N9), 
        .F(n4604) );
  MUX U4657 ( .IN0(n4604), .IN1(n4603), .SEL(N10), .F(n4605) );
  MUX U4658 ( .IN0(\registers[10][19] ), .IN1(\registers[11][19] ), .SEL(N9), 
        .F(n4606) );
  MUX U4659 ( .IN0(\registers[8][19] ), .IN1(\registers[9][19] ), .SEL(N9), 
        .F(n4607) );
  MUX U4660 ( .IN0(n4607), .IN1(n4606), .SEL(N10), .F(n4608) );
  MUX U4661 ( .IN0(n4608), .IN1(n4605), .SEL(N11), .F(n4609) );
  MUX U4662 ( .IN0(\registers[6][19] ), .IN1(\registers[7][19] ), .SEL(N9), 
        .F(n4610) );
  MUX U4663 ( .IN0(\registers[4][19] ), .IN1(\registers[5][19] ), .SEL(N9), 
        .F(n4611) );
  MUX U4664 ( .IN0(n4611), .IN1(n4610), .SEL(N10), .F(n4612) );
  MUX U4665 ( .IN0(\registers[2][19] ), .IN1(\registers[3][19] ), .SEL(N9), 
        .F(n4613) );
  MUX U4667 ( .IN0(n4614), .IN1(n4613), .SEL(N10), .F(n4615) );
  MUX U4668 ( .IN0(n4615), .IN1(n4612), .SEL(N11), .F(n4616) );
  MUX U4669 ( .IN0(n4616), .IN1(n4609), .SEL(N12), .F(n4617) );
  MUX U4670 ( .IN0(n4617), .IN1(n4602), .SEL(N13), .F(reg_source_out[19]) );
  MUX U4671 ( .IN0(\registers[30][20] ), .IN1(\registers[31][20] ), .SEL(N9), 
        .F(n4618) );
  MUX U4672 ( .IN0(\registers[28][20] ), .IN1(\registers[29][20] ), .SEL(N9), 
        .F(n4619) );
  MUX U4673 ( .IN0(n4619), .IN1(n4618), .SEL(N10), .F(n4620) );
  MUX U4674 ( .IN0(\registers[26][20] ), .IN1(\registers[27][20] ), .SEL(N9), 
        .F(n4621) );
  MUX U4675 ( .IN0(\registers[24][20] ), .IN1(\registers[25][20] ), .SEL(N9), 
        .F(n4622) );
  MUX U4676 ( .IN0(n4622), .IN1(n4621), .SEL(N10), .F(n4623) );
  MUX U4677 ( .IN0(n4623), .IN1(n4620), .SEL(N11), .F(n4624) );
  MUX U4678 ( .IN0(\registers[22][20] ), .IN1(\registers[23][20] ), .SEL(N9), 
        .F(n4625) );
  MUX U4679 ( .IN0(\registers[20][20] ), .IN1(\registers[21][20] ), .SEL(N9), 
        .F(n4626) );
  MUX U4680 ( .IN0(n4626), .IN1(n4625), .SEL(N10), .F(n4627) );
  MUX U4681 ( .IN0(\registers[18][20] ), .IN1(\registers[19][20] ), .SEL(N9), 
        .F(n4628) );
  MUX U4682 ( .IN0(\registers[16][20] ), .IN1(\registers[17][20] ), .SEL(N9), 
        .F(n4629) );
  MUX U4683 ( .IN0(n4629), .IN1(n4628), .SEL(N10), .F(n4630) );
  MUX U4684 ( .IN0(n4630), .IN1(n4627), .SEL(N11), .F(n4631) );
  MUX U4685 ( .IN0(n4631), .IN1(n4624), .SEL(N12), .F(n4632) );
  MUX U4686 ( .IN0(\registers[14][20] ), .IN1(\registers[15][20] ), .SEL(N9), 
        .F(n4633) );
  MUX U4687 ( .IN0(\registers[12][20] ), .IN1(\registers[13][20] ), .SEL(N9), 
        .F(n4634) );
  MUX U4688 ( .IN0(n4634), .IN1(n4633), .SEL(N10), .F(n4635) );
  MUX U4689 ( .IN0(\registers[10][20] ), .IN1(\registers[11][20] ), .SEL(N9), 
        .F(n4636) );
  MUX U4690 ( .IN0(\registers[8][20] ), .IN1(\registers[9][20] ), .SEL(N9), 
        .F(n4637) );
  MUX U4691 ( .IN0(n4637), .IN1(n4636), .SEL(N10), .F(n4638) );
  MUX U4692 ( .IN0(n4638), .IN1(n4635), .SEL(N11), .F(n4639) );
  MUX U4693 ( .IN0(\registers[6][20] ), .IN1(\registers[7][20] ), .SEL(N9), 
        .F(n4640) );
  MUX U4694 ( .IN0(\registers[4][20] ), .IN1(\registers[5][20] ), .SEL(N9), 
        .F(n4641) );
  MUX U4695 ( .IN0(n4641), .IN1(n4640), .SEL(N10), .F(n4642) );
  MUX U4696 ( .IN0(\registers[2][20] ), .IN1(\registers[3][20] ), .SEL(N9), 
        .F(n4643) );
  MUX U4698 ( .IN0(n4644), .IN1(n4643), .SEL(N10), .F(n4645) );
  MUX U4699 ( .IN0(n4645), .IN1(n4642), .SEL(N11), .F(n4646) );
  MUX U4700 ( .IN0(n4646), .IN1(n4639), .SEL(N12), .F(n4647) );
  MUX U4701 ( .IN0(n4647), .IN1(n4632), .SEL(N13), .F(reg_source_out[20]) );
  MUX U4702 ( .IN0(\registers[30][21] ), .IN1(\registers[31][21] ), .SEL(N9), 
        .F(n4648) );
  MUX U4703 ( .IN0(\registers[28][21] ), .IN1(\registers[29][21] ), .SEL(N9), 
        .F(n4649) );
  MUX U4704 ( .IN0(n4649), .IN1(n4648), .SEL(N10), .F(n4650) );
  MUX U4705 ( .IN0(\registers[26][21] ), .IN1(\registers[27][21] ), .SEL(N9), 
        .F(n4651) );
  MUX U4706 ( .IN0(\registers[24][21] ), .IN1(\registers[25][21] ), .SEL(N9), 
        .F(n4652) );
  MUX U4707 ( .IN0(n4652), .IN1(n4651), .SEL(N10), .F(n4653) );
  MUX U4708 ( .IN0(n4653), .IN1(n4650), .SEL(N11), .F(n4654) );
  MUX U4709 ( .IN0(\registers[22][21] ), .IN1(\registers[23][21] ), .SEL(N9), 
        .F(n4655) );
  MUX U4710 ( .IN0(\registers[20][21] ), .IN1(\registers[21][21] ), .SEL(N9), 
        .F(n4656) );
  MUX U4711 ( .IN0(n4656), .IN1(n4655), .SEL(N10), .F(n4657) );
  MUX U4712 ( .IN0(\registers[18][21] ), .IN1(\registers[19][21] ), .SEL(N9), 
        .F(n4658) );
  MUX U4713 ( .IN0(\registers[16][21] ), .IN1(\registers[17][21] ), .SEL(N9), 
        .F(n4659) );
  MUX U4714 ( .IN0(n4659), .IN1(n4658), .SEL(N10), .F(n4660) );
  MUX U4715 ( .IN0(n4660), .IN1(n4657), .SEL(N11), .F(n4661) );
  MUX U4716 ( .IN0(n4661), .IN1(n4654), .SEL(N12), .F(n4662) );
  MUX U4717 ( .IN0(\registers[14][21] ), .IN1(\registers[15][21] ), .SEL(N9), 
        .F(n4663) );
  MUX U4718 ( .IN0(\registers[12][21] ), .IN1(\registers[13][21] ), .SEL(N9), 
        .F(n4664) );
  MUX U4719 ( .IN0(n4664), .IN1(n4663), .SEL(N10), .F(n4665) );
  MUX U4720 ( .IN0(\registers[10][21] ), .IN1(\registers[11][21] ), .SEL(N9), 
        .F(n4666) );
  MUX U4721 ( .IN0(\registers[8][21] ), .IN1(\registers[9][21] ), .SEL(N9), 
        .F(n4667) );
  MUX U4722 ( .IN0(n4667), .IN1(n4666), .SEL(N10), .F(n4668) );
  MUX U4723 ( .IN0(n4668), .IN1(n4665), .SEL(N11), .F(n4669) );
  MUX U4724 ( .IN0(\registers[6][21] ), .IN1(\registers[7][21] ), .SEL(N9), 
        .F(n4670) );
  MUX U4725 ( .IN0(\registers[4][21] ), .IN1(\registers[5][21] ), .SEL(N9), 
        .F(n4671) );
  MUX U4726 ( .IN0(n4671), .IN1(n4670), .SEL(N10), .F(n4672) );
  MUX U4727 ( .IN0(\registers[2][21] ), .IN1(\registers[3][21] ), .SEL(N9), 
        .F(n4673) );
  MUX U4729 ( .IN0(n4674), .IN1(n4673), .SEL(N10), .F(n4675) );
  MUX U4730 ( .IN0(n4675), .IN1(n4672), .SEL(N11), .F(n4676) );
  MUX U4731 ( .IN0(n4676), .IN1(n4669), .SEL(N12), .F(n4677) );
  MUX U4732 ( .IN0(n4677), .IN1(n4662), .SEL(N13), .F(reg_source_out[21]) );
  MUX U4733 ( .IN0(\registers[30][22] ), .IN1(\registers[31][22] ), .SEL(N9), 
        .F(n4678) );
  MUX U4734 ( .IN0(\registers[28][22] ), .IN1(\registers[29][22] ), .SEL(N9), 
        .F(n4679) );
  MUX U4735 ( .IN0(n4679), .IN1(n4678), .SEL(N10), .F(n4680) );
  MUX U4736 ( .IN0(\registers[26][22] ), .IN1(\registers[27][22] ), .SEL(N9), 
        .F(n4681) );
  MUX U4737 ( .IN0(\registers[24][22] ), .IN1(\registers[25][22] ), .SEL(N9), 
        .F(n4682) );
  MUX U4738 ( .IN0(n4682), .IN1(n4681), .SEL(N10), .F(n4683) );
  MUX U4739 ( .IN0(n4683), .IN1(n4680), .SEL(N11), .F(n4684) );
  MUX U4740 ( .IN0(\registers[22][22] ), .IN1(\registers[23][22] ), .SEL(N9), 
        .F(n4685) );
  MUX U4741 ( .IN0(\registers[20][22] ), .IN1(\registers[21][22] ), .SEL(N9), 
        .F(n4686) );
  MUX U4742 ( .IN0(n4686), .IN1(n4685), .SEL(N10), .F(n4687) );
  MUX U4743 ( .IN0(\registers[18][22] ), .IN1(\registers[19][22] ), .SEL(N9), 
        .F(n4688) );
  MUX U4744 ( .IN0(\registers[16][22] ), .IN1(\registers[17][22] ), .SEL(N9), 
        .F(n4689) );
  MUX U4745 ( .IN0(n4689), .IN1(n4688), .SEL(N10), .F(n4690) );
  MUX U4746 ( .IN0(n4690), .IN1(n4687), .SEL(N11), .F(n4691) );
  MUX U4747 ( .IN0(n4691), .IN1(n4684), .SEL(N12), .F(n4692) );
  MUX U4748 ( .IN0(\registers[14][22] ), .IN1(\registers[15][22] ), .SEL(N9), 
        .F(n4693) );
  MUX U4749 ( .IN0(\registers[12][22] ), .IN1(\registers[13][22] ), .SEL(N9), 
        .F(n4694) );
  MUX U4750 ( .IN0(n4694), .IN1(n4693), .SEL(N10), .F(n4695) );
  MUX U4751 ( .IN0(\registers[10][22] ), .IN1(\registers[11][22] ), .SEL(N9), 
        .F(n4696) );
  MUX U4752 ( .IN0(\registers[8][22] ), .IN1(\registers[9][22] ), .SEL(N9), 
        .F(n4697) );
  MUX U4753 ( .IN0(n4697), .IN1(n4696), .SEL(N10), .F(n4698) );
  MUX U4754 ( .IN0(n4698), .IN1(n4695), .SEL(N11), .F(n4699) );
  MUX U4755 ( .IN0(\registers[6][22] ), .IN1(\registers[7][22] ), .SEL(N9), 
        .F(n4700) );
  MUX U4756 ( .IN0(\registers[4][22] ), .IN1(\registers[5][22] ), .SEL(N9), 
        .F(n4701) );
  MUX U4757 ( .IN0(n4701), .IN1(n4700), .SEL(N10), .F(n4702) );
  MUX U4758 ( .IN0(\registers[2][22] ), .IN1(\registers[3][22] ), .SEL(N9), 
        .F(n4703) );
  MUX U4760 ( .IN0(n4704), .IN1(n4703), .SEL(N10), .F(n4705) );
  MUX U4761 ( .IN0(n4705), .IN1(n4702), .SEL(N11), .F(n4706) );
  MUX U4762 ( .IN0(n4706), .IN1(n4699), .SEL(N12), .F(n4707) );
  MUX U4763 ( .IN0(n4707), .IN1(n4692), .SEL(N13), .F(reg_source_out[22]) );
  MUX U4764 ( .IN0(\registers[30][23] ), .IN1(\registers[31][23] ), .SEL(N9), 
        .F(n4708) );
  MUX U4765 ( .IN0(\registers[28][23] ), .IN1(\registers[29][23] ), .SEL(N9), 
        .F(n4709) );
  MUX U4766 ( .IN0(n4709), .IN1(n4708), .SEL(N10), .F(n4710) );
  MUX U4767 ( .IN0(\registers[26][23] ), .IN1(\registers[27][23] ), .SEL(N9), 
        .F(n4711) );
  MUX U4768 ( .IN0(\registers[24][23] ), .IN1(\registers[25][23] ), .SEL(N9), 
        .F(n4712) );
  MUX U4769 ( .IN0(n4712), .IN1(n4711), .SEL(N10), .F(n4713) );
  MUX U4770 ( .IN0(n4713), .IN1(n4710), .SEL(N11), .F(n4714) );
  MUX U4771 ( .IN0(\registers[22][23] ), .IN1(\registers[23][23] ), .SEL(N9), 
        .F(n4715) );
  MUX U4772 ( .IN0(\registers[20][23] ), .IN1(\registers[21][23] ), .SEL(N9), 
        .F(n4716) );
  MUX U4773 ( .IN0(n4716), .IN1(n4715), .SEL(N10), .F(n4717) );
  MUX U4774 ( .IN0(\registers[18][23] ), .IN1(\registers[19][23] ), .SEL(N9), 
        .F(n4718) );
  MUX U4775 ( .IN0(\registers[16][23] ), .IN1(\registers[17][23] ), .SEL(N9), 
        .F(n4719) );
  MUX U4776 ( .IN0(n4719), .IN1(n4718), .SEL(N10), .F(n4720) );
  MUX U4777 ( .IN0(n4720), .IN1(n4717), .SEL(N11), .F(n4721) );
  MUX U4778 ( .IN0(n4721), .IN1(n4714), .SEL(N12), .F(n4722) );
  MUX U4779 ( .IN0(\registers[14][23] ), .IN1(\registers[15][23] ), .SEL(N9), 
        .F(n4723) );
  MUX U4780 ( .IN0(\registers[12][23] ), .IN1(\registers[13][23] ), .SEL(N9), 
        .F(n4724) );
  MUX U4781 ( .IN0(n4724), .IN1(n4723), .SEL(N10), .F(n4725) );
  MUX U4782 ( .IN0(\registers[10][23] ), .IN1(\registers[11][23] ), .SEL(N9), 
        .F(n4726) );
  MUX U4783 ( .IN0(\registers[8][23] ), .IN1(\registers[9][23] ), .SEL(N9), 
        .F(n4727) );
  MUX U4784 ( .IN0(n4727), .IN1(n4726), .SEL(N10), .F(n4728) );
  MUX U4785 ( .IN0(n4728), .IN1(n4725), .SEL(N11), .F(n4729) );
  MUX U4786 ( .IN0(\registers[6][23] ), .IN1(\registers[7][23] ), .SEL(N9), 
        .F(n4730) );
  MUX U4787 ( .IN0(\registers[4][23] ), .IN1(\registers[5][23] ), .SEL(N9), 
        .F(n4731) );
  MUX U4788 ( .IN0(n4731), .IN1(n4730), .SEL(N10), .F(n4732) );
  MUX U4789 ( .IN0(\registers[2][23] ), .IN1(\registers[3][23] ), .SEL(N9), 
        .F(n4733) );
  MUX U4791 ( .IN0(n4734), .IN1(n4733), .SEL(N10), .F(n4735) );
  MUX U4792 ( .IN0(n4735), .IN1(n4732), .SEL(N11), .F(n4736) );
  MUX U4793 ( .IN0(n4736), .IN1(n4729), .SEL(N12), .F(n4737) );
  MUX U4794 ( .IN0(n4737), .IN1(n4722), .SEL(N13), .F(reg_source_out[23]) );
  MUX U4795 ( .IN0(\registers[30][24] ), .IN1(\registers[31][24] ), .SEL(N9), 
        .F(n4738) );
  MUX U4796 ( .IN0(\registers[28][24] ), .IN1(\registers[29][24] ), .SEL(N9), 
        .F(n4739) );
  MUX U4797 ( .IN0(n4739), .IN1(n4738), .SEL(N10), .F(n4740) );
  MUX U4798 ( .IN0(\registers[26][24] ), .IN1(\registers[27][24] ), .SEL(N9), 
        .F(n4741) );
  MUX U4799 ( .IN0(\registers[24][24] ), .IN1(\registers[25][24] ), .SEL(N9), 
        .F(n4742) );
  MUX U4800 ( .IN0(n4742), .IN1(n4741), .SEL(N10), .F(n4743) );
  MUX U4801 ( .IN0(n4743), .IN1(n4740), .SEL(N11), .F(n4744) );
  MUX U4802 ( .IN0(\registers[22][24] ), .IN1(\registers[23][24] ), .SEL(N9), 
        .F(n4745) );
  MUX U4803 ( .IN0(\registers[20][24] ), .IN1(\registers[21][24] ), .SEL(N9), 
        .F(n4746) );
  MUX U4804 ( .IN0(n4746), .IN1(n4745), .SEL(N10), .F(n4747) );
  MUX U4805 ( .IN0(\registers[18][24] ), .IN1(\registers[19][24] ), .SEL(N9), 
        .F(n4748) );
  MUX U4806 ( .IN0(\registers[16][24] ), .IN1(\registers[17][24] ), .SEL(N9), 
        .F(n4749) );
  MUX U4807 ( .IN0(n4749), .IN1(n4748), .SEL(N10), .F(n4750) );
  MUX U4808 ( .IN0(n4750), .IN1(n4747), .SEL(N11), .F(n4751) );
  MUX U4809 ( .IN0(n4751), .IN1(n4744), .SEL(N12), .F(n4752) );
  MUX U4810 ( .IN0(\registers[14][24] ), .IN1(\registers[15][24] ), .SEL(N9), 
        .F(n4753) );
  MUX U4811 ( .IN0(\registers[12][24] ), .IN1(\registers[13][24] ), .SEL(N9), 
        .F(n4754) );
  MUX U4812 ( .IN0(n4754), .IN1(n4753), .SEL(N10), .F(n4755) );
  MUX U4813 ( .IN0(\registers[10][24] ), .IN1(\registers[11][24] ), .SEL(N9), 
        .F(n4756) );
  MUX U4814 ( .IN0(\registers[8][24] ), .IN1(\registers[9][24] ), .SEL(N9), 
        .F(n4757) );
  MUX U4815 ( .IN0(n4757), .IN1(n4756), .SEL(N10), .F(n4758) );
  MUX U4816 ( .IN0(n4758), .IN1(n4755), .SEL(N11), .F(n4759) );
  MUX U4817 ( .IN0(\registers[6][24] ), .IN1(\registers[7][24] ), .SEL(N9), 
        .F(n4760) );
  MUX U4818 ( .IN0(\registers[4][24] ), .IN1(\registers[5][24] ), .SEL(N9), 
        .F(n4761) );
  MUX U4819 ( .IN0(n4761), .IN1(n4760), .SEL(N10), .F(n4762) );
  MUX U4820 ( .IN0(\registers[2][24] ), .IN1(\registers[3][24] ), .SEL(N9), 
        .F(n4763) );
  MUX U4822 ( .IN0(n4764), .IN1(n4763), .SEL(N10), .F(n4765) );
  MUX U4823 ( .IN0(n4765), .IN1(n4762), .SEL(N11), .F(n4766) );
  MUX U4824 ( .IN0(n4766), .IN1(n4759), .SEL(N12), .F(n4767) );
  MUX U4825 ( .IN0(n4767), .IN1(n4752), .SEL(N13), .F(reg_source_out[24]) );
  MUX U4826 ( .IN0(\registers[30][25] ), .IN1(\registers[31][25] ), .SEL(N9), 
        .F(n4768) );
  MUX U4827 ( .IN0(\registers[28][25] ), .IN1(\registers[29][25] ), .SEL(N9), 
        .F(n4769) );
  MUX U4828 ( .IN0(n4769), .IN1(n4768), .SEL(N10), .F(n4770) );
  MUX U4829 ( .IN0(\registers[26][25] ), .IN1(\registers[27][25] ), .SEL(N9), 
        .F(n4771) );
  MUX U4830 ( .IN0(\registers[24][25] ), .IN1(\registers[25][25] ), .SEL(N9), 
        .F(n4772) );
  MUX U4831 ( .IN0(n4772), .IN1(n4771), .SEL(N10), .F(n4773) );
  MUX U4832 ( .IN0(n4773), .IN1(n4770), .SEL(N11), .F(n4774) );
  MUX U4833 ( .IN0(\registers[22][25] ), .IN1(\registers[23][25] ), .SEL(N9), 
        .F(n4775) );
  MUX U4834 ( .IN0(\registers[20][25] ), .IN1(\registers[21][25] ), .SEL(N9), 
        .F(n4776) );
  MUX U4835 ( .IN0(n4776), .IN1(n4775), .SEL(N10), .F(n4777) );
  MUX U4836 ( .IN0(\registers[18][25] ), .IN1(\registers[19][25] ), .SEL(N9), 
        .F(n4778) );
  MUX U4837 ( .IN0(\registers[16][25] ), .IN1(\registers[17][25] ), .SEL(N9), 
        .F(n4779) );
  MUX U4838 ( .IN0(n4779), .IN1(n4778), .SEL(N10), .F(n4780) );
  MUX U4839 ( .IN0(n4780), .IN1(n4777), .SEL(N11), .F(n4781) );
  MUX U4840 ( .IN0(n4781), .IN1(n4774), .SEL(N12), .F(n4782) );
  MUX U4841 ( .IN0(\registers[14][25] ), .IN1(\registers[15][25] ), .SEL(N9), 
        .F(n4783) );
  MUX U4842 ( .IN0(\registers[12][25] ), .IN1(\registers[13][25] ), .SEL(N9), 
        .F(n4784) );
  MUX U4843 ( .IN0(n4784), .IN1(n4783), .SEL(N10), .F(n4785) );
  MUX U4844 ( .IN0(\registers[10][25] ), .IN1(\registers[11][25] ), .SEL(N9), 
        .F(n4786) );
  MUX U4845 ( .IN0(\registers[8][25] ), .IN1(\registers[9][25] ), .SEL(N9), 
        .F(n4787) );
  MUX U4846 ( .IN0(n4787), .IN1(n4786), .SEL(N10), .F(n4788) );
  MUX U4847 ( .IN0(n4788), .IN1(n4785), .SEL(N11), .F(n4789) );
  MUX U4848 ( .IN0(\registers[6][25] ), .IN1(\registers[7][25] ), .SEL(N9), 
        .F(n4790) );
  MUX U4849 ( .IN0(\registers[4][25] ), .IN1(\registers[5][25] ), .SEL(N9), 
        .F(n4791) );
  MUX U4850 ( .IN0(n4791), .IN1(n4790), .SEL(N10), .F(n4792) );
  MUX U4851 ( .IN0(\registers[2][25] ), .IN1(\registers[3][25] ), .SEL(N9), 
        .F(n4793) );
  MUX U4853 ( .IN0(n4794), .IN1(n4793), .SEL(N10), .F(n4795) );
  MUX U4854 ( .IN0(n4795), .IN1(n4792), .SEL(N11), .F(n4796) );
  MUX U4855 ( .IN0(n4796), .IN1(n4789), .SEL(N12), .F(n4797) );
  MUX U4856 ( .IN0(n4797), .IN1(n4782), .SEL(N13), .F(reg_source_out[25]) );
  MUX U4857 ( .IN0(\registers[30][26] ), .IN1(\registers[31][26] ), .SEL(N9), 
        .F(n4798) );
  MUX U4858 ( .IN0(\registers[28][26] ), .IN1(\registers[29][26] ), .SEL(N9), 
        .F(n4799) );
  MUX U4859 ( .IN0(n4799), .IN1(n4798), .SEL(N10), .F(n4800) );
  MUX U4860 ( .IN0(\registers[26][26] ), .IN1(\registers[27][26] ), .SEL(N9), 
        .F(n4801) );
  MUX U4861 ( .IN0(\registers[24][26] ), .IN1(\registers[25][26] ), .SEL(N9), 
        .F(n4802) );
  MUX U4862 ( .IN0(n4802), .IN1(n4801), .SEL(N10), .F(n4803) );
  MUX U4863 ( .IN0(n4803), .IN1(n4800), .SEL(N11), .F(n4804) );
  MUX U4864 ( .IN0(\registers[22][26] ), .IN1(\registers[23][26] ), .SEL(N9), 
        .F(n4805) );
  MUX U4865 ( .IN0(\registers[20][26] ), .IN1(\registers[21][26] ), .SEL(N9), 
        .F(n4806) );
  MUX U4866 ( .IN0(n4806), .IN1(n4805), .SEL(N10), .F(n4807) );
  MUX U4867 ( .IN0(\registers[18][26] ), .IN1(\registers[19][26] ), .SEL(N9), 
        .F(n4808) );
  MUX U4868 ( .IN0(\registers[16][26] ), .IN1(\registers[17][26] ), .SEL(N9), 
        .F(n4809) );
  MUX U4869 ( .IN0(n4809), .IN1(n4808), .SEL(N10), .F(n4810) );
  MUX U4870 ( .IN0(n4810), .IN1(n4807), .SEL(N11), .F(n4811) );
  MUX U4871 ( .IN0(n4811), .IN1(n4804), .SEL(N12), .F(n4812) );
  MUX U4872 ( .IN0(\registers[14][26] ), .IN1(\registers[15][26] ), .SEL(N9), 
        .F(n4813) );
  MUX U4873 ( .IN0(\registers[12][26] ), .IN1(\registers[13][26] ), .SEL(N9), 
        .F(n4814) );
  MUX U4874 ( .IN0(n4814), .IN1(n4813), .SEL(N10), .F(n4815) );
  MUX U4875 ( .IN0(\registers[10][26] ), .IN1(\registers[11][26] ), .SEL(N9), 
        .F(n4816) );
  MUX U4876 ( .IN0(\registers[8][26] ), .IN1(\registers[9][26] ), .SEL(N9), 
        .F(n4817) );
  MUX U4877 ( .IN0(n4817), .IN1(n4816), .SEL(N10), .F(n4818) );
  MUX U4878 ( .IN0(n4818), .IN1(n4815), .SEL(N11), .F(n4819) );
  MUX U4879 ( .IN0(\registers[6][26] ), .IN1(\registers[7][26] ), .SEL(N9), 
        .F(n4820) );
  MUX U4880 ( .IN0(\registers[4][26] ), .IN1(\registers[5][26] ), .SEL(N9), 
        .F(n4821) );
  MUX U4881 ( .IN0(n4821), .IN1(n4820), .SEL(N10), .F(n4822) );
  MUX U4882 ( .IN0(\registers[2][26] ), .IN1(\registers[3][26] ), .SEL(N9), 
        .F(n4823) );
  MUX U4884 ( .IN0(n4824), .IN1(n4823), .SEL(N10), .F(n4825) );
  MUX U4885 ( .IN0(n4825), .IN1(n4822), .SEL(N11), .F(n4826) );
  MUX U4886 ( .IN0(n4826), .IN1(n4819), .SEL(N12), .F(n4827) );
  MUX U4887 ( .IN0(n4827), .IN1(n4812), .SEL(N13), .F(reg_source_out[26]) );
  MUX U4888 ( .IN0(\registers[30][27] ), .IN1(\registers[31][27] ), .SEL(N9), 
        .F(n4828) );
  MUX U4889 ( .IN0(\registers[28][27] ), .IN1(\registers[29][27] ), .SEL(N9), 
        .F(n4829) );
  MUX U4890 ( .IN0(n4829), .IN1(n4828), .SEL(N10), .F(n4830) );
  MUX U4891 ( .IN0(\registers[26][27] ), .IN1(\registers[27][27] ), .SEL(N9), 
        .F(n4831) );
  MUX U4892 ( .IN0(\registers[24][27] ), .IN1(\registers[25][27] ), .SEL(N9), 
        .F(n4832) );
  MUX U4893 ( .IN0(n4832), .IN1(n4831), .SEL(N10), .F(n4833) );
  MUX U4894 ( .IN0(n4833), .IN1(n4830), .SEL(N11), .F(n4834) );
  MUX U4895 ( .IN0(\registers[22][27] ), .IN1(\registers[23][27] ), .SEL(N9), 
        .F(n4835) );
  MUX U4896 ( .IN0(\registers[20][27] ), .IN1(\registers[21][27] ), .SEL(N9), 
        .F(n4836) );
  MUX U4897 ( .IN0(n4836), .IN1(n4835), .SEL(N10), .F(n4837) );
  MUX U4898 ( .IN0(\registers[18][27] ), .IN1(\registers[19][27] ), .SEL(N9), 
        .F(n4838) );
  MUX U4899 ( .IN0(\registers[16][27] ), .IN1(\registers[17][27] ), .SEL(N9), 
        .F(n4839) );
  MUX U4900 ( .IN0(n4839), .IN1(n4838), .SEL(N10), .F(n4840) );
  MUX U4901 ( .IN0(n4840), .IN1(n4837), .SEL(N11), .F(n4841) );
  MUX U4902 ( .IN0(n4841), .IN1(n4834), .SEL(N12), .F(n4842) );
  MUX U4903 ( .IN0(\registers[14][27] ), .IN1(\registers[15][27] ), .SEL(N9), 
        .F(n4843) );
  MUX U4904 ( .IN0(\registers[12][27] ), .IN1(\registers[13][27] ), .SEL(N9), 
        .F(n4844) );
  MUX U4905 ( .IN0(n4844), .IN1(n4843), .SEL(N10), .F(n4845) );
  MUX U4906 ( .IN0(\registers[10][27] ), .IN1(\registers[11][27] ), .SEL(N9), 
        .F(n4846) );
  MUX U4907 ( .IN0(\registers[8][27] ), .IN1(\registers[9][27] ), .SEL(N9), 
        .F(n4847) );
  MUX U4908 ( .IN0(n4847), .IN1(n4846), .SEL(N10), .F(n4848) );
  MUX U4909 ( .IN0(n4848), .IN1(n4845), .SEL(N11), .F(n4849) );
  MUX U4910 ( .IN0(\registers[6][27] ), .IN1(\registers[7][27] ), .SEL(N9), 
        .F(n4850) );
  MUX U4911 ( .IN0(\registers[4][27] ), .IN1(\registers[5][27] ), .SEL(N9), 
        .F(n4851) );
  MUX U4912 ( .IN0(n4851), .IN1(n4850), .SEL(N10), .F(n4852) );
  MUX U4913 ( .IN0(\registers[2][27] ), .IN1(\registers[3][27] ), .SEL(N9), 
        .F(n4853) );
  MUX U4915 ( .IN0(n4854), .IN1(n4853), .SEL(N10), .F(n4855) );
  MUX U4916 ( .IN0(n4855), .IN1(n4852), .SEL(N11), .F(n4856) );
  MUX U4917 ( .IN0(n4856), .IN1(n4849), .SEL(N12), .F(n4857) );
  MUX U4918 ( .IN0(n4857), .IN1(n4842), .SEL(N13), .F(reg_source_out[27]) );
  MUX U4919 ( .IN0(\registers[30][28] ), .IN1(\registers[31][28] ), .SEL(N9), 
        .F(n4858) );
  MUX U4920 ( .IN0(\registers[28][28] ), .IN1(\registers[29][28] ), .SEL(N9), 
        .F(n4859) );
  MUX U4921 ( .IN0(n4859), .IN1(n4858), .SEL(N10), .F(n4860) );
  MUX U4922 ( .IN0(\registers[26][28] ), .IN1(\registers[27][28] ), .SEL(N9), 
        .F(n4861) );
  MUX U4923 ( .IN0(\registers[24][28] ), .IN1(\registers[25][28] ), .SEL(N9), 
        .F(n4862) );
  MUX U4924 ( .IN0(n4862), .IN1(n4861), .SEL(N10), .F(n4863) );
  MUX U4925 ( .IN0(n4863), .IN1(n4860), .SEL(N11), .F(n4864) );
  MUX U4926 ( .IN0(\registers[22][28] ), .IN1(\registers[23][28] ), .SEL(N9), 
        .F(n4865) );
  MUX U4927 ( .IN0(\registers[20][28] ), .IN1(\registers[21][28] ), .SEL(N9), 
        .F(n4866) );
  MUX U4928 ( .IN0(n4866), .IN1(n4865), .SEL(N10), .F(n4867) );
  MUX U4929 ( .IN0(\registers[18][28] ), .IN1(\registers[19][28] ), .SEL(N9), 
        .F(n4868) );
  MUX U4930 ( .IN0(\registers[16][28] ), .IN1(\registers[17][28] ), .SEL(N9), 
        .F(n4869) );
  MUX U4931 ( .IN0(n4869), .IN1(n4868), .SEL(N10), .F(n4870) );
  MUX U4932 ( .IN0(n4870), .IN1(n4867), .SEL(N11), .F(n4871) );
  MUX U4933 ( .IN0(n4871), .IN1(n4864), .SEL(N12), .F(n4872) );
  MUX U4934 ( .IN0(\registers[14][28] ), .IN1(\registers[15][28] ), .SEL(N9), 
        .F(n4873) );
  MUX U4935 ( .IN0(\registers[12][28] ), .IN1(\registers[13][28] ), .SEL(N9), 
        .F(n4874) );
  MUX U4936 ( .IN0(n4874), .IN1(n4873), .SEL(N10), .F(n4875) );
  MUX U4937 ( .IN0(\registers[10][28] ), .IN1(\registers[11][28] ), .SEL(N9), 
        .F(n4876) );
  MUX U4938 ( .IN0(\registers[8][28] ), .IN1(\registers[9][28] ), .SEL(N9), 
        .F(n4877) );
  MUX U4939 ( .IN0(n4877), .IN1(n4876), .SEL(N10), .F(n4878) );
  MUX U4940 ( .IN0(n4878), .IN1(n4875), .SEL(N11), .F(n4879) );
  MUX U4941 ( .IN0(\registers[6][28] ), .IN1(\registers[7][28] ), .SEL(N9), 
        .F(n4880) );
  MUX U4942 ( .IN0(\registers[4][28] ), .IN1(\registers[5][28] ), .SEL(N9), 
        .F(n4881) );
  MUX U4943 ( .IN0(n4881), .IN1(n4880), .SEL(N10), .F(n4882) );
  MUX U4944 ( .IN0(\registers[2][28] ), .IN1(\registers[3][28] ), .SEL(N9), 
        .F(n4883) );
  MUX U4946 ( .IN0(n4884), .IN1(n4883), .SEL(N10), .F(n4885) );
  MUX U4947 ( .IN0(n4885), .IN1(n4882), .SEL(N11), .F(n4886) );
  MUX U4948 ( .IN0(n4886), .IN1(n4879), .SEL(N12), .F(n4887) );
  MUX U4949 ( .IN0(n4887), .IN1(n4872), .SEL(N13), .F(reg_source_out[28]) );
  MUX U4950 ( .IN0(\registers[30][29] ), .IN1(\registers[31][29] ), .SEL(N9), 
        .F(n4888) );
  MUX U4951 ( .IN0(\registers[28][29] ), .IN1(\registers[29][29] ), .SEL(N9), 
        .F(n4889) );
  MUX U4952 ( .IN0(n4889), .IN1(n4888), .SEL(N10), .F(n4890) );
  MUX U4953 ( .IN0(\registers[26][29] ), .IN1(\registers[27][29] ), .SEL(N9), 
        .F(n4891) );
  MUX U4954 ( .IN0(\registers[24][29] ), .IN1(\registers[25][29] ), .SEL(N9), 
        .F(n4892) );
  MUX U4955 ( .IN0(n4892), .IN1(n4891), .SEL(N10), .F(n4893) );
  MUX U4956 ( .IN0(n4893), .IN1(n4890), .SEL(N11), .F(n4894) );
  MUX U4957 ( .IN0(\registers[22][29] ), .IN1(\registers[23][29] ), .SEL(N9), 
        .F(n4895) );
  MUX U4958 ( .IN0(\registers[20][29] ), .IN1(\registers[21][29] ), .SEL(N9), 
        .F(n4896) );
  MUX U4959 ( .IN0(n4896), .IN1(n4895), .SEL(N10), .F(n4897) );
  MUX U4960 ( .IN0(\registers[18][29] ), .IN1(\registers[19][29] ), .SEL(N9), 
        .F(n4898) );
  MUX U4961 ( .IN0(\registers[16][29] ), .IN1(\registers[17][29] ), .SEL(N9), 
        .F(n4899) );
  MUX U4962 ( .IN0(n4899), .IN1(n4898), .SEL(N10), .F(n4900) );
  MUX U4963 ( .IN0(n4900), .IN1(n4897), .SEL(N11), .F(n4901) );
  MUX U4964 ( .IN0(n4901), .IN1(n4894), .SEL(N12), .F(n4902) );
  MUX U4965 ( .IN0(\registers[14][29] ), .IN1(\registers[15][29] ), .SEL(N9), 
        .F(n4903) );
  MUX U4966 ( .IN0(\registers[12][29] ), .IN1(\registers[13][29] ), .SEL(N9), 
        .F(n4904) );
  MUX U4967 ( .IN0(n4904), .IN1(n4903), .SEL(N10), .F(n4905) );
  MUX U4968 ( .IN0(\registers[10][29] ), .IN1(\registers[11][29] ), .SEL(N9), 
        .F(n4906) );
  MUX U4969 ( .IN0(\registers[8][29] ), .IN1(\registers[9][29] ), .SEL(N9), 
        .F(n4907) );
  MUX U4970 ( .IN0(n4907), .IN1(n4906), .SEL(N10), .F(n4908) );
  MUX U4971 ( .IN0(n4908), .IN1(n4905), .SEL(N11), .F(n4909) );
  MUX U4972 ( .IN0(\registers[6][29] ), .IN1(\registers[7][29] ), .SEL(N9), 
        .F(n4910) );
  MUX U4973 ( .IN0(\registers[4][29] ), .IN1(\registers[5][29] ), .SEL(N9), 
        .F(n4911) );
  MUX U4974 ( .IN0(n4911), .IN1(n4910), .SEL(N10), .F(n4912) );
  MUX U4975 ( .IN0(\registers[2][29] ), .IN1(\registers[3][29] ), .SEL(N9), 
        .F(n4913) );
  MUX U4977 ( .IN0(n4914), .IN1(n4913), .SEL(N10), .F(n4915) );
  MUX U4978 ( .IN0(n4915), .IN1(n4912), .SEL(N11), .F(n4916) );
  MUX U4979 ( .IN0(n4916), .IN1(n4909), .SEL(N12), .F(n4917) );
  MUX U4980 ( .IN0(n4917), .IN1(n4902), .SEL(N13), .F(reg_source_out[29]) );
  MUX U4981 ( .IN0(\registers[30][30] ), .IN1(\registers[31][30] ), .SEL(N9), 
        .F(n4918) );
  MUX U4982 ( .IN0(\registers[28][30] ), .IN1(\registers[29][30] ), .SEL(N9), 
        .F(n4919) );
  MUX U4983 ( .IN0(n4919), .IN1(n4918), .SEL(N10), .F(n4920) );
  MUX U4984 ( .IN0(\registers[26][30] ), .IN1(\registers[27][30] ), .SEL(N9), 
        .F(n4921) );
  MUX U4985 ( .IN0(\registers[24][30] ), .IN1(\registers[25][30] ), .SEL(N9), 
        .F(n4922) );
  MUX U4986 ( .IN0(n4922), .IN1(n4921), .SEL(N10), .F(n4923) );
  MUX U4987 ( .IN0(n4923), .IN1(n4920), .SEL(N11), .F(n4924) );
  MUX U4988 ( .IN0(\registers[22][30] ), .IN1(\registers[23][30] ), .SEL(N9), 
        .F(n4925) );
  MUX U4989 ( .IN0(\registers[20][30] ), .IN1(\registers[21][30] ), .SEL(N9), 
        .F(n4926) );
  MUX U4990 ( .IN0(n4926), .IN1(n4925), .SEL(N10), .F(n4927) );
  MUX U4991 ( .IN0(\registers[18][30] ), .IN1(\registers[19][30] ), .SEL(N9), 
        .F(n4928) );
  MUX U4992 ( .IN0(\registers[16][30] ), .IN1(\registers[17][30] ), .SEL(N9), 
        .F(n4929) );
  MUX U4993 ( .IN0(n4929), .IN1(n4928), .SEL(N10), .F(n4930) );
  MUX U4994 ( .IN0(n4930), .IN1(n4927), .SEL(N11), .F(n4931) );
  MUX U4995 ( .IN0(n4931), .IN1(n4924), .SEL(N12), .F(n4932) );
  MUX U4996 ( .IN0(\registers[14][30] ), .IN1(\registers[15][30] ), .SEL(N9), 
        .F(n4933) );
  MUX U4997 ( .IN0(\registers[12][30] ), .IN1(\registers[13][30] ), .SEL(N9), 
        .F(n4934) );
  MUX U4998 ( .IN0(n4934), .IN1(n4933), .SEL(N10), .F(n4935) );
  MUX U4999 ( .IN0(\registers[10][30] ), .IN1(\registers[11][30] ), .SEL(N9), 
        .F(n4936) );
  MUX U5000 ( .IN0(\registers[8][30] ), .IN1(\registers[9][30] ), .SEL(N9), 
        .F(n4937) );
  MUX U5001 ( .IN0(n4937), .IN1(n4936), .SEL(N10), .F(n4938) );
  MUX U5002 ( .IN0(n4938), .IN1(n4935), .SEL(N11), .F(n4939) );
  MUX U5003 ( .IN0(\registers[6][30] ), .IN1(\registers[7][30] ), .SEL(N9), 
        .F(n4940) );
  MUX U5004 ( .IN0(\registers[4][30] ), .IN1(\registers[5][30] ), .SEL(N9), 
        .F(n4941) );
  MUX U5005 ( .IN0(n4941), .IN1(n4940), .SEL(N10), .F(n4942) );
  MUX U5006 ( .IN0(\registers[2][30] ), .IN1(\registers[3][30] ), .SEL(N9), 
        .F(n4943) );
  MUX U5008 ( .IN0(n4944), .IN1(n4943), .SEL(N10), .F(n4945) );
  MUX U5009 ( .IN0(n4945), .IN1(n4942), .SEL(N11), .F(n4946) );
  MUX U5010 ( .IN0(n4946), .IN1(n4939), .SEL(N12), .F(n4947) );
  MUX U5011 ( .IN0(n4947), .IN1(n4932), .SEL(N13), .F(reg_source_out[30]) );
  MUX U5012 ( .IN0(\registers[30][31] ), .IN1(\registers[31][31] ), .SEL(N9), 
        .F(n4948) );
  MUX U5013 ( .IN0(\registers[28][31] ), .IN1(\registers[29][31] ), .SEL(N9), 
        .F(n4949) );
  MUX U5014 ( .IN0(n4949), .IN1(n4948), .SEL(N10), .F(n4950) );
  MUX U5015 ( .IN0(\registers[26][31] ), .IN1(\registers[27][31] ), .SEL(N9), 
        .F(n4951) );
  MUX U5016 ( .IN0(\registers[24][31] ), .IN1(\registers[25][31] ), .SEL(N9), 
        .F(n4952) );
  MUX U5017 ( .IN0(n4952), .IN1(n4951), .SEL(N10), .F(n4953) );
  MUX U5018 ( .IN0(n4953), .IN1(n4950), .SEL(N11), .F(n4954) );
  MUX U5019 ( .IN0(\registers[22][31] ), .IN1(\registers[23][31] ), .SEL(N9), 
        .F(n4955) );
  MUX U5020 ( .IN0(\registers[20][31] ), .IN1(\registers[21][31] ), .SEL(N9), 
        .F(n4956) );
  MUX U5021 ( .IN0(n4956), .IN1(n4955), .SEL(N10), .F(n4957) );
  MUX U5022 ( .IN0(\registers[18][31] ), .IN1(\registers[19][31] ), .SEL(N9), 
        .F(n4958) );
  MUX U5023 ( .IN0(\registers[16][31] ), .IN1(\registers[17][31] ), .SEL(N9), 
        .F(n4959) );
  MUX U5024 ( .IN0(n4959), .IN1(n4958), .SEL(N10), .F(n4960) );
  MUX U5025 ( .IN0(n4960), .IN1(n4957), .SEL(N11), .F(n4961) );
  MUX U5026 ( .IN0(n4961), .IN1(n4954), .SEL(N12), .F(n4962) );
  MUX U5027 ( .IN0(\registers[14][31] ), .IN1(\registers[15][31] ), .SEL(N9), 
        .F(n4963) );
  MUX U5028 ( .IN0(\registers[12][31] ), .IN1(\registers[13][31] ), .SEL(N9), 
        .F(n4964) );
  MUX U5029 ( .IN0(n4964), .IN1(n4963), .SEL(N10), .F(n4965) );
  MUX U5030 ( .IN0(\registers[10][31] ), .IN1(\registers[11][31] ), .SEL(N9), 
        .F(n4966) );
  MUX U5031 ( .IN0(\registers[8][31] ), .IN1(\registers[9][31] ), .SEL(N9), 
        .F(n4967) );
  MUX U5032 ( .IN0(n4967), .IN1(n4966), .SEL(N10), .F(n4968) );
  MUX U5033 ( .IN0(n4968), .IN1(n4965), .SEL(N11), .F(n4969) );
  MUX U5034 ( .IN0(\registers[6][31] ), .IN1(\registers[7][31] ), .SEL(N9), 
        .F(n4970) );
  MUX U5035 ( .IN0(\registers[4][31] ), .IN1(\registers[5][31] ), .SEL(N9), 
        .F(n4971) );
  MUX U5036 ( .IN0(n4971), .IN1(n4970), .SEL(N10), .F(n4972) );
  MUX U5037 ( .IN0(\registers[2][31] ), .IN1(\registers[3][31] ), .SEL(N9), 
        .F(n4973) );
  MUX U5039 ( .IN0(n4974), .IN1(n4973), .SEL(N10), .F(n4975) );
  MUX U5040 ( .IN0(n4975), .IN1(n4972), .SEL(N11), .F(n4976) );
  MUX U5041 ( .IN0(n4976), .IN1(n4969), .SEL(N12), .F(n4977) );
  MUX U5042 ( .IN0(n4977), .IN1(n4962), .SEL(N13), .F(reg_source_out[31]) );
  MUX U5043 ( .IN0(\registers[30][0] ), .IN1(\registers[31][0] ), .SEL(N14), 
        .F(n4978) );
  MUX U5044 ( .IN0(\registers[28][0] ), .IN1(\registers[29][0] ), .SEL(N14), 
        .F(n4979) );
  MUX U5045 ( .IN0(n4979), .IN1(n4978), .SEL(N15), .F(n4980) );
  MUX U5046 ( .IN0(\registers[26][0] ), .IN1(\registers[27][0] ), .SEL(N14), 
        .F(n4981) );
  MUX U5047 ( .IN0(\registers[24][0] ), .IN1(\registers[25][0] ), .SEL(N14), 
        .F(n4982) );
  MUX U5048 ( .IN0(n4982), .IN1(n4981), .SEL(N15), .F(n4983) );
  MUX U5049 ( .IN0(n4983), .IN1(n4980), .SEL(N16), .F(n4984) );
  MUX U5050 ( .IN0(\registers[22][0] ), .IN1(\registers[23][0] ), .SEL(N14), 
        .F(n4985) );
  MUX U5051 ( .IN0(\registers[20][0] ), .IN1(\registers[21][0] ), .SEL(N14), 
        .F(n4986) );
  MUX U5052 ( .IN0(n4986), .IN1(n4985), .SEL(N15), .F(n4987) );
  MUX U5053 ( .IN0(\registers[18][0] ), .IN1(\registers[19][0] ), .SEL(N14), 
        .F(n4988) );
  MUX U5054 ( .IN0(\registers[16][0] ), .IN1(\registers[17][0] ), .SEL(N14), 
        .F(n4989) );
  MUX U5055 ( .IN0(n4989), .IN1(n4988), .SEL(N15), .F(n4990) );
  MUX U5056 ( .IN0(n4990), .IN1(n4987), .SEL(N16), .F(n4991) );
  MUX U5057 ( .IN0(n4991), .IN1(n4984), .SEL(N17), .F(n4992) );
  MUX U5058 ( .IN0(\registers[14][0] ), .IN1(\registers[15][0] ), .SEL(N14), 
        .F(n4993) );
  MUX U5059 ( .IN0(\registers[12][0] ), .IN1(\registers[13][0] ), .SEL(N14), 
        .F(n4994) );
  MUX U5060 ( .IN0(n4994), .IN1(n4993), .SEL(N15), .F(n4995) );
  MUX U5061 ( .IN0(\registers[10][0] ), .IN1(\registers[11][0] ), .SEL(N14), 
        .F(n4996) );
  MUX U5062 ( .IN0(\registers[8][0] ), .IN1(\registers[9][0] ), .SEL(N14), .F(
        n4997) );
  MUX U5063 ( .IN0(n4997), .IN1(n4996), .SEL(N15), .F(n4998) );
  MUX U5064 ( .IN0(n4998), .IN1(n4995), .SEL(N16), .F(n4999) );
  MUX U5065 ( .IN0(\registers[6][0] ), .IN1(\registers[7][0] ), .SEL(N14), .F(
        n5000) );
  MUX U5066 ( .IN0(\registers[4][0] ), .IN1(\registers[5][0] ), .SEL(N14), .F(
        n5001) );
  MUX U5067 ( .IN0(n5001), .IN1(n5000), .SEL(N15), .F(n5002) );
  MUX U5068 ( .IN0(\registers[2][0] ), .IN1(\registers[3][0] ), .SEL(N14), .F(
        n5003) );
  MUX U5070 ( .IN0(n5004), .IN1(n5003), .SEL(N15), .F(n5005) );
  MUX U5071 ( .IN0(n5005), .IN1(n5002), .SEL(N16), .F(n5006) );
  MUX U5072 ( .IN0(n5006), .IN1(n4999), .SEL(N17), .F(n5007) );
  MUX U5073 ( .IN0(n5007), .IN1(n4992), .SEL(N18), .F(reg_target_out[0]) );
  MUX U5074 ( .IN0(\registers[30][1] ), .IN1(\registers[31][1] ), .SEL(N14), 
        .F(n5008) );
  MUX U5075 ( .IN0(\registers[28][1] ), .IN1(\registers[29][1] ), .SEL(N14), 
        .F(n5009) );
  MUX U5076 ( .IN0(n5009), .IN1(n5008), .SEL(N15), .F(n5010) );
  MUX U5077 ( .IN0(\registers[26][1] ), .IN1(\registers[27][1] ), .SEL(N14), 
        .F(n5011) );
  MUX U5078 ( .IN0(\registers[24][1] ), .IN1(\registers[25][1] ), .SEL(N14), 
        .F(n5012) );
  MUX U5079 ( .IN0(n5012), .IN1(n5011), .SEL(N15), .F(n5013) );
  MUX U5080 ( .IN0(n5013), .IN1(n5010), .SEL(N16), .F(n5014) );
  MUX U5081 ( .IN0(\registers[22][1] ), .IN1(\registers[23][1] ), .SEL(N14), 
        .F(n5015) );
  MUX U5082 ( .IN0(\registers[20][1] ), .IN1(\registers[21][1] ), .SEL(N14), 
        .F(n5016) );
  MUX U5083 ( .IN0(n5016), .IN1(n5015), .SEL(N15), .F(n5017) );
  MUX U5084 ( .IN0(\registers[18][1] ), .IN1(\registers[19][1] ), .SEL(N14), 
        .F(n5018) );
  MUX U5085 ( .IN0(\registers[16][1] ), .IN1(\registers[17][1] ), .SEL(N14), 
        .F(n5019) );
  MUX U5086 ( .IN0(n5019), .IN1(n5018), .SEL(N15), .F(n5020) );
  MUX U5087 ( .IN0(n5020), .IN1(n5017), .SEL(N16), .F(n5021) );
  MUX U5088 ( .IN0(n5021), .IN1(n5014), .SEL(N17), .F(n5022) );
  MUX U5089 ( .IN0(\registers[14][1] ), .IN1(\registers[15][1] ), .SEL(N14), 
        .F(n5023) );
  MUX U5090 ( .IN0(\registers[12][1] ), .IN1(\registers[13][1] ), .SEL(N14), 
        .F(n5024) );
  MUX U5091 ( .IN0(n5024), .IN1(n5023), .SEL(N15), .F(n5025) );
  MUX U5092 ( .IN0(\registers[10][1] ), .IN1(\registers[11][1] ), .SEL(N14), 
        .F(n5026) );
  MUX U5093 ( .IN0(\registers[8][1] ), .IN1(\registers[9][1] ), .SEL(N14), .F(
        n5027) );
  MUX U5094 ( .IN0(n5027), .IN1(n5026), .SEL(N15), .F(n5028) );
  MUX U5095 ( .IN0(n5028), .IN1(n5025), .SEL(N16), .F(n5029) );
  MUX U5096 ( .IN0(\registers[6][1] ), .IN1(\registers[7][1] ), .SEL(N14), .F(
        n5030) );
  MUX U5097 ( .IN0(\registers[4][1] ), .IN1(\registers[5][1] ), .SEL(N14), .F(
        n5031) );
  MUX U5098 ( .IN0(n5031), .IN1(n5030), .SEL(N15), .F(n5032) );
  MUX U5099 ( .IN0(\registers[2][1] ), .IN1(\registers[3][1] ), .SEL(N14), .F(
        n5033) );
  MUX U5101 ( .IN0(n5034), .IN1(n5033), .SEL(N15), .F(n5035) );
  MUX U5102 ( .IN0(n5035), .IN1(n5032), .SEL(N16), .F(n5036) );
  MUX U5103 ( .IN0(n5036), .IN1(n5029), .SEL(N17), .F(n5037) );
  MUX U5104 ( .IN0(n5037), .IN1(n5022), .SEL(N18), .F(reg_target_out[1]) );
  MUX U5105 ( .IN0(\registers[30][2] ), .IN1(\registers[31][2] ), .SEL(N14), 
        .F(n5038) );
  MUX U5106 ( .IN0(\registers[28][2] ), .IN1(\registers[29][2] ), .SEL(N14), 
        .F(n5039) );
  MUX U5107 ( .IN0(n5039), .IN1(n5038), .SEL(N15), .F(n5040) );
  MUX U5108 ( .IN0(\registers[26][2] ), .IN1(\registers[27][2] ), .SEL(N14), 
        .F(n5041) );
  MUX U5109 ( .IN0(\registers[24][2] ), .IN1(\registers[25][2] ), .SEL(N14), 
        .F(n5042) );
  MUX U5110 ( .IN0(n5042), .IN1(n5041), .SEL(N15), .F(n5043) );
  MUX U5111 ( .IN0(n5043), .IN1(n5040), .SEL(N16), .F(n5044) );
  MUX U5112 ( .IN0(\registers[22][2] ), .IN1(\registers[23][2] ), .SEL(N14), 
        .F(n5045) );
  MUX U5113 ( .IN0(\registers[20][2] ), .IN1(\registers[21][2] ), .SEL(N14), 
        .F(n5046) );
  MUX U5114 ( .IN0(n5046), .IN1(n5045), .SEL(N15), .F(n5047) );
  MUX U5115 ( .IN0(\registers[18][2] ), .IN1(\registers[19][2] ), .SEL(N14), 
        .F(n5048) );
  MUX U5116 ( .IN0(\registers[16][2] ), .IN1(\registers[17][2] ), .SEL(N14), 
        .F(n5049) );
  MUX U5117 ( .IN0(n5049), .IN1(n5048), .SEL(N15), .F(n5050) );
  MUX U5118 ( .IN0(n5050), .IN1(n5047), .SEL(N16), .F(n5051) );
  MUX U5119 ( .IN0(n5051), .IN1(n5044), .SEL(N17), .F(n5052) );
  MUX U5120 ( .IN0(\registers[14][2] ), .IN1(\registers[15][2] ), .SEL(N14), 
        .F(n5053) );
  MUX U5121 ( .IN0(\registers[12][2] ), .IN1(\registers[13][2] ), .SEL(N14), 
        .F(n5054) );
  MUX U5122 ( .IN0(n5054), .IN1(n5053), .SEL(N15), .F(n5055) );
  MUX U5123 ( .IN0(\registers[10][2] ), .IN1(\registers[11][2] ), .SEL(N14), 
        .F(n5056) );
  MUX U5124 ( .IN0(\registers[8][2] ), .IN1(\registers[9][2] ), .SEL(N14), .F(
        n5057) );
  MUX U5125 ( .IN0(n5057), .IN1(n5056), .SEL(N15), .F(n5058) );
  MUX U5126 ( .IN0(n5058), .IN1(n5055), .SEL(N16), .F(n5059) );
  MUX U5127 ( .IN0(\registers[6][2] ), .IN1(\registers[7][2] ), .SEL(N14), .F(
        n5060) );
  MUX U5128 ( .IN0(\registers[4][2] ), .IN1(\registers[5][2] ), .SEL(N14), .F(
        n5061) );
  MUX U5129 ( .IN0(n5061), .IN1(n5060), .SEL(N15), .F(n5062) );
  MUX U5130 ( .IN0(\registers[2][2] ), .IN1(\registers[3][2] ), .SEL(N14), .F(
        n5063) );
  MUX U5132 ( .IN0(n5064), .IN1(n5063), .SEL(N15), .F(n5065) );
  MUX U5133 ( .IN0(n5065), .IN1(n5062), .SEL(N16), .F(n5066) );
  MUX U5134 ( .IN0(n5066), .IN1(n5059), .SEL(N17), .F(n5067) );
  MUX U5135 ( .IN0(n5067), .IN1(n5052), .SEL(N18), .F(reg_target_out[2]) );
  MUX U5136 ( .IN0(\registers[30][3] ), .IN1(\registers[31][3] ), .SEL(N14), 
        .F(n5068) );
  MUX U5137 ( .IN0(\registers[28][3] ), .IN1(\registers[29][3] ), .SEL(N14), 
        .F(n5069) );
  MUX U5138 ( .IN0(n5069), .IN1(n5068), .SEL(N15), .F(n5070) );
  MUX U5139 ( .IN0(\registers[26][3] ), .IN1(\registers[27][3] ), .SEL(N14), 
        .F(n5071) );
  MUX U5140 ( .IN0(\registers[24][3] ), .IN1(\registers[25][3] ), .SEL(N14), 
        .F(n5072) );
  MUX U5141 ( .IN0(n5072), .IN1(n5071), .SEL(N15), .F(n5073) );
  MUX U5142 ( .IN0(n5073), .IN1(n5070), .SEL(N16), .F(n5074) );
  MUX U5143 ( .IN0(\registers[22][3] ), .IN1(\registers[23][3] ), .SEL(N14), 
        .F(n5075) );
  MUX U5144 ( .IN0(\registers[20][3] ), .IN1(\registers[21][3] ), .SEL(N14), 
        .F(n5076) );
  MUX U5145 ( .IN0(n5076), .IN1(n5075), .SEL(N15), .F(n5077) );
  MUX U5146 ( .IN0(\registers[18][3] ), .IN1(\registers[19][3] ), .SEL(N14), 
        .F(n5078) );
  MUX U5147 ( .IN0(\registers[16][3] ), .IN1(\registers[17][3] ), .SEL(N14), 
        .F(n5079) );
  MUX U5148 ( .IN0(n5079), .IN1(n5078), .SEL(N15), .F(n5080) );
  MUX U5149 ( .IN0(n5080), .IN1(n5077), .SEL(N16), .F(n5081) );
  MUX U5150 ( .IN0(n5081), .IN1(n5074), .SEL(N17), .F(n5082) );
  MUX U5151 ( .IN0(\registers[14][3] ), .IN1(\registers[15][3] ), .SEL(N14), 
        .F(n5083) );
  MUX U5152 ( .IN0(\registers[12][3] ), .IN1(\registers[13][3] ), .SEL(N14), 
        .F(n5084) );
  MUX U5153 ( .IN0(n5084), .IN1(n5083), .SEL(N15), .F(n5085) );
  MUX U5154 ( .IN0(\registers[10][3] ), .IN1(\registers[11][3] ), .SEL(N14), 
        .F(n5086) );
  MUX U5155 ( .IN0(\registers[8][3] ), .IN1(\registers[9][3] ), .SEL(N14), .F(
        n5087) );
  MUX U5156 ( .IN0(n5087), .IN1(n5086), .SEL(N15), .F(n5088) );
  MUX U5157 ( .IN0(n5088), .IN1(n5085), .SEL(N16), .F(n5089) );
  MUX U5158 ( .IN0(\registers[6][3] ), .IN1(\registers[7][3] ), .SEL(N14), .F(
        n5090) );
  MUX U5159 ( .IN0(\registers[4][3] ), .IN1(\registers[5][3] ), .SEL(N14), .F(
        n5091) );
  MUX U5160 ( .IN0(n5091), .IN1(n5090), .SEL(N15), .F(n5092) );
  MUX U5161 ( .IN0(\registers[2][3] ), .IN1(\registers[3][3] ), .SEL(N14), .F(
        n5093) );
  MUX U5163 ( .IN0(n5094), .IN1(n5093), .SEL(N15), .F(n5095) );
  MUX U5164 ( .IN0(n5095), .IN1(n5092), .SEL(N16), .F(n5096) );
  MUX U5165 ( .IN0(n5096), .IN1(n5089), .SEL(N17), .F(n5097) );
  MUX U5166 ( .IN0(n5097), .IN1(n5082), .SEL(N18), .F(reg_target_out[3]) );
  MUX U5167 ( .IN0(\registers[30][4] ), .IN1(\registers[31][4] ), .SEL(N14), 
        .F(n5098) );
  MUX U5168 ( .IN0(\registers[28][4] ), .IN1(\registers[29][4] ), .SEL(N14), 
        .F(n5099) );
  MUX U5169 ( .IN0(n5099), .IN1(n5098), .SEL(N15), .F(n5100) );
  MUX U5170 ( .IN0(\registers[26][4] ), .IN1(\registers[27][4] ), .SEL(N14), 
        .F(n5101) );
  MUX U5171 ( .IN0(\registers[24][4] ), .IN1(\registers[25][4] ), .SEL(N14), 
        .F(n5102) );
  MUX U5172 ( .IN0(n5102), .IN1(n5101), .SEL(N15), .F(n5103) );
  MUX U5173 ( .IN0(n5103), .IN1(n5100), .SEL(N16), .F(n5104) );
  MUX U5174 ( .IN0(\registers[22][4] ), .IN1(\registers[23][4] ), .SEL(N14), 
        .F(n5105) );
  MUX U5175 ( .IN0(\registers[20][4] ), .IN1(\registers[21][4] ), .SEL(N14), 
        .F(n5106) );
  MUX U5176 ( .IN0(n5106), .IN1(n5105), .SEL(N15), .F(n5107) );
  MUX U5177 ( .IN0(\registers[18][4] ), .IN1(\registers[19][4] ), .SEL(N14), 
        .F(n5108) );
  MUX U5178 ( .IN0(\registers[16][4] ), .IN1(\registers[17][4] ), .SEL(N14), 
        .F(n5109) );
  MUX U5179 ( .IN0(n5109), .IN1(n5108), .SEL(N15), .F(n5110) );
  MUX U5180 ( .IN0(n5110), .IN1(n5107), .SEL(N16), .F(n5111) );
  MUX U5181 ( .IN0(n5111), .IN1(n5104), .SEL(N17), .F(n5112) );
  MUX U5182 ( .IN0(\registers[14][4] ), .IN1(\registers[15][4] ), .SEL(N14), 
        .F(n5113) );
  MUX U5183 ( .IN0(\registers[12][4] ), .IN1(\registers[13][4] ), .SEL(N14), 
        .F(n5114) );
  MUX U5184 ( .IN0(n5114), .IN1(n5113), .SEL(N15), .F(n5115) );
  MUX U5185 ( .IN0(\registers[10][4] ), .IN1(\registers[11][4] ), .SEL(N14), 
        .F(n5116) );
  MUX U5186 ( .IN0(\registers[8][4] ), .IN1(\registers[9][4] ), .SEL(N14), .F(
        n5117) );
  MUX U5187 ( .IN0(n5117), .IN1(n5116), .SEL(N15), .F(n5118) );
  MUX U5188 ( .IN0(n5118), .IN1(n5115), .SEL(N16), .F(n5119) );
  MUX U5189 ( .IN0(\registers[6][4] ), .IN1(\registers[7][4] ), .SEL(N14), .F(
        n5120) );
  MUX U5190 ( .IN0(\registers[4][4] ), .IN1(\registers[5][4] ), .SEL(N14), .F(
        n5121) );
  MUX U5191 ( .IN0(n5121), .IN1(n5120), .SEL(N15), .F(n5122) );
  MUX U5192 ( .IN0(\registers[2][4] ), .IN1(\registers[3][4] ), .SEL(N14), .F(
        n5123) );
  MUX U5194 ( .IN0(n5124), .IN1(n5123), .SEL(N15), .F(n5125) );
  MUX U5195 ( .IN0(n5125), .IN1(n5122), .SEL(N16), .F(n5126) );
  MUX U5196 ( .IN0(n5126), .IN1(n5119), .SEL(N17), .F(n5127) );
  MUX U5197 ( .IN0(n5127), .IN1(n5112), .SEL(N18), .F(reg_target_out[4]) );
  MUX U5198 ( .IN0(\registers[30][5] ), .IN1(\registers[31][5] ), .SEL(N14), 
        .F(n5128) );
  MUX U5199 ( .IN0(\registers[28][5] ), .IN1(\registers[29][5] ), .SEL(N14), 
        .F(n5129) );
  MUX U5200 ( .IN0(n5129), .IN1(n5128), .SEL(N15), .F(n5130) );
  MUX U5201 ( .IN0(\registers[26][5] ), .IN1(\registers[27][5] ), .SEL(N14), 
        .F(n5131) );
  MUX U5202 ( .IN0(\registers[24][5] ), .IN1(\registers[25][5] ), .SEL(N14), 
        .F(n5132) );
  MUX U5203 ( .IN0(n5132), .IN1(n5131), .SEL(N15), .F(n5133) );
  MUX U5204 ( .IN0(n5133), .IN1(n5130), .SEL(N16), .F(n5134) );
  MUX U5205 ( .IN0(\registers[22][5] ), .IN1(\registers[23][5] ), .SEL(N14), 
        .F(n5135) );
  MUX U5206 ( .IN0(\registers[20][5] ), .IN1(\registers[21][5] ), .SEL(N14), 
        .F(n5136) );
  MUX U5207 ( .IN0(n5136), .IN1(n5135), .SEL(N15), .F(n5137) );
  MUX U5208 ( .IN0(\registers[18][5] ), .IN1(\registers[19][5] ), .SEL(N14), 
        .F(n5138) );
  MUX U5209 ( .IN0(\registers[16][5] ), .IN1(\registers[17][5] ), .SEL(N14), 
        .F(n5139) );
  MUX U5210 ( .IN0(n5139), .IN1(n5138), .SEL(N15), .F(n5140) );
  MUX U5211 ( .IN0(n5140), .IN1(n5137), .SEL(N16), .F(n5141) );
  MUX U5212 ( .IN0(n5141), .IN1(n5134), .SEL(N17), .F(n5142) );
  MUX U5213 ( .IN0(\registers[14][5] ), .IN1(\registers[15][5] ), .SEL(N14), 
        .F(n5143) );
  MUX U5214 ( .IN0(\registers[12][5] ), .IN1(\registers[13][5] ), .SEL(N14), 
        .F(n5144) );
  MUX U5215 ( .IN0(n5144), .IN1(n5143), .SEL(N15), .F(n5145) );
  MUX U5216 ( .IN0(\registers[10][5] ), .IN1(\registers[11][5] ), .SEL(N14), 
        .F(n5146) );
  MUX U5217 ( .IN0(\registers[8][5] ), .IN1(\registers[9][5] ), .SEL(N14), .F(
        n5147) );
  MUX U5218 ( .IN0(n5147), .IN1(n5146), .SEL(N15), .F(n5148) );
  MUX U5219 ( .IN0(n5148), .IN1(n5145), .SEL(N16), .F(n5149) );
  MUX U5220 ( .IN0(\registers[6][5] ), .IN1(\registers[7][5] ), .SEL(N14), .F(
        n5150) );
  MUX U5221 ( .IN0(\registers[4][5] ), .IN1(\registers[5][5] ), .SEL(N14), .F(
        n5151) );
  MUX U5222 ( .IN0(n5151), .IN1(n5150), .SEL(N15), .F(n5152) );
  MUX U5223 ( .IN0(\registers[2][5] ), .IN1(\registers[3][5] ), .SEL(N14), .F(
        n5153) );
  MUX U5225 ( .IN0(n5154), .IN1(n5153), .SEL(N15), .F(n5155) );
  MUX U5226 ( .IN0(n5155), .IN1(n5152), .SEL(N16), .F(n5156) );
  MUX U5227 ( .IN0(n5156), .IN1(n5149), .SEL(N17), .F(n5157) );
  MUX U5228 ( .IN0(n5157), .IN1(n5142), .SEL(N18), .F(reg_target_out[5]) );
  MUX U5229 ( .IN0(\registers[30][6] ), .IN1(\registers[31][6] ), .SEL(N14), 
        .F(n5158) );
  MUX U5230 ( .IN0(\registers[28][6] ), .IN1(\registers[29][6] ), .SEL(N14), 
        .F(n5159) );
  MUX U5231 ( .IN0(n5159), .IN1(n5158), .SEL(N15), .F(n5160) );
  MUX U5232 ( .IN0(\registers[26][6] ), .IN1(\registers[27][6] ), .SEL(N14), 
        .F(n5161) );
  MUX U5233 ( .IN0(\registers[24][6] ), .IN1(\registers[25][6] ), .SEL(N14), 
        .F(n5162) );
  MUX U5234 ( .IN0(n5162), .IN1(n5161), .SEL(N15), .F(n5163) );
  MUX U5235 ( .IN0(n5163), .IN1(n5160), .SEL(N16), .F(n5164) );
  MUX U5236 ( .IN0(\registers[22][6] ), .IN1(\registers[23][6] ), .SEL(N14), 
        .F(n5165) );
  MUX U5237 ( .IN0(\registers[20][6] ), .IN1(\registers[21][6] ), .SEL(N14), 
        .F(n5166) );
  MUX U5238 ( .IN0(n5166), .IN1(n5165), .SEL(N15), .F(n5167) );
  MUX U5239 ( .IN0(\registers[18][6] ), .IN1(\registers[19][6] ), .SEL(N14), 
        .F(n5168) );
  MUX U5240 ( .IN0(\registers[16][6] ), .IN1(\registers[17][6] ), .SEL(N14), 
        .F(n5169) );
  MUX U5241 ( .IN0(n5169), .IN1(n5168), .SEL(N15), .F(n5170) );
  MUX U5242 ( .IN0(n5170), .IN1(n5167), .SEL(N16), .F(n5171) );
  MUX U5243 ( .IN0(n5171), .IN1(n5164), .SEL(N17), .F(n5172) );
  MUX U5244 ( .IN0(\registers[14][6] ), .IN1(\registers[15][6] ), .SEL(N14), 
        .F(n5173) );
  MUX U5245 ( .IN0(\registers[12][6] ), .IN1(\registers[13][6] ), .SEL(N14), 
        .F(n5174) );
  MUX U5246 ( .IN0(n5174), .IN1(n5173), .SEL(N15), .F(n5175) );
  MUX U5247 ( .IN0(\registers[10][6] ), .IN1(\registers[11][6] ), .SEL(N14), 
        .F(n5176) );
  MUX U5248 ( .IN0(\registers[8][6] ), .IN1(\registers[9][6] ), .SEL(N14), .F(
        n5177) );
  MUX U5249 ( .IN0(n5177), .IN1(n5176), .SEL(N15), .F(n5178) );
  MUX U5250 ( .IN0(n5178), .IN1(n5175), .SEL(N16), .F(n5179) );
  MUX U5251 ( .IN0(\registers[6][6] ), .IN1(\registers[7][6] ), .SEL(N14), .F(
        n5180) );
  MUX U5252 ( .IN0(\registers[4][6] ), .IN1(\registers[5][6] ), .SEL(N14), .F(
        n5181) );
  MUX U5253 ( .IN0(n5181), .IN1(n5180), .SEL(N15), .F(n5182) );
  MUX U5254 ( .IN0(\registers[2][6] ), .IN1(\registers[3][6] ), .SEL(N14), .F(
        n5183) );
  MUX U5256 ( .IN0(n5184), .IN1(n5183), .SEL(N15), .F(n5185) );
  MUX U5257 ( .IN0(n5185), .IN1(n5182), .SEL(N16), .F(n5186) );
  MUX U5258 ( .IN0(n5186), .IN1(n5179), .SEL(N17), .F(n5187) );
  MUX U5259 ( .IN0(n5187), .IN1(n5172), .SEL(N18), .F(reg_target_out[6]) );
  MUX U5260 ( .IN0(\registers[30][7] ), .IN1(\registers[31][7] ), .SEL(N14), 
        .F(n5188) );
  MUX U5261 ( .IN0(\registers[28][7] ), .IN1(\registers[29][7] ), .SEL(N14), 
        .F(n5189) );
  MUX U5262 ( .IN0(n5189), .IN1(n5188), .SEL(N15), .F(n5190) );
  MUX U5263 ( .IN0(\registers[26][7] ), .IN1(\registers[27][7] ), .SEL(N14), 
        .F(n5191) );
  MUX U5264 ( .IN0(\registers[24][7] ), .IN1(\registers[25][7] ), .SEL(N14), 
        .F(n5192) );
  MUX U5265 ( .IN0(n5192), .IN1(n5191), .SEL(N15), .F(n5193) );
  MUX U5266 ( .IN0(n5193), .IN1(n5190), .SEL(N16), .F(n5194) );
  MUX U5267 ( .IN0(\registers[22][7] ), .IN1(\registers[23][7] ), .SEL(N14), 
        .F(n5195) );
  MUX U5268 ( .IN0(\registers[20][7] ), .IN1(\registers[21][7] ), .SEL(N14), 
        .F(n5196) );
  MUX U5269 ( .IN0(n5196), .IN1(n5195), .SEL(N15), .F(n5197) );
  MUX U5270 ( .IN0(\registers[18][7] ), .IN1(\registers[19][7] ), .SEL(N14), 
        .F(n5198) );
  MUX U5271 ( .IN0(\registers[16][7] ), .IN1(\registers[17][7] ), .SEL(N14), 
        .F(n5199) );
  MUX U5272 ( .IN0(n5199), .IN1(n5198), .SEL(N15), .F(n5200) );
  MUX U5273 ( .IN0(n5200), .IN1(n5197), .SEL(N16), .F(n5201) );
  MUX U5274 ( .IN0(n5201), .IN1(n5194), .SEL(N17), .F(n5202) );
  MUX U5275 ( .IN0(\registers[14][7] ), .IN1(\registers[15][7] ), .SEL(N14), 
        .F(n5203) );
  MUX U5276 ( .IN0(\registers[12][7] ), .IN1(\registers[13][7] ), .SEL(N14), 
        .F(n5204) );
  MUX U5277 ( .IN0(n5204), .IN1(n5203), .SEL(N15), .F(n5205) );
  MUX U5278 ( .IN0(\registers[10][7] ), .IN1(\registers[11][7] ), .SEL(N14), 
        .F(n5206) );
  MUX U5279 ( .IN0(\registers[8][7] ), .IN1(\registers[9][7] ), .SEL(N14), .F(
        n5207) );
  MUX U5280 ( .IN0(n5207), .IN1(n5206), .SEL(N15), .F(n5208) );
  MUX U5281 ( .IN0(n5208), .IN1(n5205), .SEL(N16), .F(n5209) );
  MUX U5282 ( .IN0(\registers[6][7] ), .IN1(\registers[7][7] ), .SEL(N14), .F(
        n5210) );
  MUX U5283 ( .IN0(\registers[4][7] ), .IN1(\registers[5][7] ), .SEL(N14), .F(
        n5211) );
  MUX U5284 ( .IN0(n5211), .IN1(n5210), .SEL(N15), .F(n5212) );
  MUX U5285 ( .IN0(\registers[2][7] ), .IN1(\registers[3][7] ), .SEL(N14), .F(
        n5213) );
  MUX U5287 ( .IN0(n5214), .IN1(n5213), .SEL(N15), .F(n5215) );
  MUX U5288 ( .IN0(n5215), .IN1(n5212), .SEL(N16), .F(n5216) );
  MUX U5289 ( .IN0(n5216), .IN1(n5209), .SEL(N17), .F(n5217) );
  MUX U5290 ( .IN0(n5217), .IN1(n5202), .SEL(N18), .F(reg_target_out[7]) );
  MUX U5291 ( .IN0(\registers[30][8] ), .IN1(\registers[31][8] ), .SEL(N14), 
        .F(n5218) );
  MUX U5292 ( .IN0(\registers[28][8] ), .IN1(\registers[29][8] ), .SEL(N14), 
        .F(n5219) );
  MUX U5293 ( .IN0(n5219), .IN1(n5218), .SEL(N15), .F(n5220) );
  MUX U5294 ( .IN0(\registers[26][8] ), .IN1(\registers[27][8] ), .SEL(N14), 
        .F(n5221) );
  MUX U5295 ( .IN0(\registers[24][8] ), .IN1(\registers[25][8] ), .SEL(N14), 
        .F(n5222) );
  MUX U5296 ( .IN0(n5222), .IN1(n5221), .SEL(N15), .F(n5223) );
  MUX U5297 ( .IN0(n5223), .IN1(n5220), .SEL(N16), .F(n5224) );
  MUX U5298 ( .IN0(\registers[22][8] ), .IN1(\registers[23][8] ), .SEL(N14), 
        .F(n5225) );
  MUX U5299 ( .IN0(\registers[20][8] ), .IN1(\registers[21][8] ), .SEL(N14), 
        .F(n5226) );
  MUX U5300 ( .IN0(n5226), .IN1(n5225), .SEL(N15), .F(n5227) );
  MUX U5301 ( .IN0(\registers[18][8] ), .IN1(\registers[19][8] ), .SEL(N14), 
        .F(n5228) );
  MUX U5302 ( .IN0(\registers[16][8] ), .IN1(\registers[17][8] ), .SEL(N14), 
        .F(n5229) );
  MUX U5303 ( .IN0(n5229), .IN1(n5228), .SEL(N15), .F(n5230) );
  MUX U5304 ( .IN0(n5230), .IN1(n5227), .SEL(N16), .F(n5231) );
  MUX U5305 ( .IN0(n5231), .IN1(n5224), .SEL(N17), .F(n5232) );
  MUX U5306 ( .IN0(\registers[14][8] ), .IN1(\registers[15][8] ), .SEL(N14), 
        .F(n5233) );
  MUX U5307 ( .IN0(\registers[12][8] ), .IN1(\registers[13][8] ), .SEL(N14), 
        .F(n5234) );
  MUX U5308 ( .IN0(n5234), .IN1(n5233), .SEL(N15), .F(n5235) );
  MUX U5309 ( .IN0(\registers[10][8] ), .IN1(\registers[11][8] ), .SEL(N14), 
        .F(n5236) );
  MUX U5310 ( .IN0(\registers[8][8] ), .IN1(\registers[9][8] ), .SEL(N14), .F(
        n5237) );
  MUX U5311 ( .IN0(n5237), .IN1(n5236), .SEL(N15), .F(n5238) );
  MUX U5312 ( .IN0(n5238), .IN1(n5235), .SEL(N16), .F(n5239) );
  MUX U5313 ( .IN0(\registers[6][8] ), .IN1(\registers[7][8] ), .SEL(N14), .F(
        n5240) );
  MUX U5314 ( .IN0(\registers[4][8] ), .IN1(\registers[5][8] ), .SEL(N14), .F(
        n5241) );
  MUX U5315 ( .IN0(n5241), .IN1(n5240), .SEL(N15), .F(n5242) );
  MUX U5316 ( .IN0(\registers[2][8] ), .IN1(\registers[3][8] ), .SEL(N14), .F(
        n5243) );
  MUX U5318 ( .IN0(n5244), .IN1(n5243), .SEL(N15), .F(n5245) );
  MUX U5319 ( .IN0(n5245), .IN1(n5242), .SEL(N16), .F(n5246) );
  MUX U5320 ( .IN0(n5246), .IN1(n5239), .SEL(N17), .F(n5247) );
  MUX U5321 ( .IN0(n5247), .IN1(n5232), .SEL(N18), .F(reg_target_out[8]) );
  MUX U5322 ( .IN0(\registers[30][9] ), .IN1(\registers[31][9] ), .SEL(N14), 
        .F(n5248) );
  MUX U5323 ( .IN0(\registers[28][9] ), .IN1(\registers[29][9] ), .SEL(N14), 
        .F(n5249) );
  MUX U5324 ( .IN0(n5249), .IN1(n5248), .SEL(N15), .F(n5250) );
  MUX U5325 ( .IN0(\registers[26][9] ), .IN1(\registers[27][9] ), .SEL(N14), 
        .F(n5251) );
  MUX U5326 ( .IN0(\registers[24][9] ), .IN1(\registers[25][9] ), .SEL(N14), 
        .F(n5252) );
  MUX U5327 ( .IN0(n5252), .IN1(n5251), .SEL(N15), .F(n5253) );
  MUX U5328 ( .IN0(n5253), .IN1(n5250), .SEL(N16), .F(n5254) );
  MUX U5329 ( .IN0(\registers[22][9] ), .IN1(\registers[23][9] ), .SEL(N14), 
        .F(n5255) );
  MUX U5330 ( .IN0(\registers[20][9] ), .IN1(\registers[21][9] ), .SEL(N14), 
        .F(n5256) );
  MUX U5331 ( .IN0(n5256), .IN1(n5255), .SEL(N15), .F(n5257) );
  MUX U5332 ( .IN0(\registers[18][9] ), .IN1(\registers[19][9] ), .SEL(N14), 
        .F(n5258) );
  MUX U5333 ( .IN0(\registers[16][9] ), .IN1(\registers[17][9] ), .SEL(N14), 
        .F(n5259) );
  MUX U5334 ( .IN0(n5259), .IN1(n5258), .SEL(N15), .F(n5260) );
  MUX U5335 ( .IN0(n5260), .IN1(n5257), .SEL(N16), .F(n5261) );
  MUX U5336 ( .IN0(n5261), .IN1(n5254), .SEL(N17), .F(n5262) );
  MUX U5337 ( .IN0(\registers[14][9] ), .IN1(\registers[15][9] ), .SEL(N14), 
        .F(n5263) );
  MUX U5338 ( .IN0(\registers[12][9] ), .IN1(\registers[13][9] ), .SEL(N14), 
        .F(n5264) );
  MUX U5339 ( .IN0(n5264), .IN1(n5263), .SEL(N15), .F(n5265) );
  MUX U5340 ( .IN0(\registers[10][9] ), .IN1(\registers[11][9] ), .SEL(N14), 
        .F(n5266) );
  MUX U5341 ( .IN0(\registers[8][9] ), .IN1(\registers[9][9] ), .SEL(N14), .F(
        n5267) );
  MUX U5342 ( .IN0(n5267), .IN1(n5266), .SEL(N15), .F(n5268) );
  MUX U5343 ( .IN0(n5268), .IN1(n5265), .SEL(N16), .F(n5269) );
  MUX U5344 ( .IN0(\registers[6][9] ), .IN1(\registers[7][9] ), .SEL(N14), .F(
        n5270) );
  MUX U5345 ( .IN0(\registers[4][9] ), .IN1(\registers[5][9] ), .SEL(N14), .F(
        n5271) );
  MUX U5346 ( .IN0(n5271), .IN1(n5270), .SEL(N15), .F(n5272) );
  MUX U5347 ( .IN0(\registers[2][9] ), .IN1(\registers[3][9] ), .SEL(N14), .F(
        n5273) );
  MUX U5349 ( .IN0(n5274), .IN1(n5273), .SEL(N15), .F(n5275) );
  MUX U5350 ( .IN0(n5275), .IN1(n5272), .SEL(N16), .F(n5276) );
  MUX U5351 ( .IN0(n5276), .IN1(n5269), .SEL(N17), .F(n5277) );
  MUX U5352 ( .IN0(n5277), .IN1(n5262), .SEL(N18), .F(reg_target_out[9]) );
  MUX U5353 ( .IN0(\registers[30][10] ), .IN1(\registers[31][10] ), .SEL(N14), 
        .F(n5278) );
  MUX U5354 ( .IN0(\registers[28][10] ), .IN1(\registers[29][10] ), .SEL(N14), 
        .F(n5279) );
  MUX U5355 ( .IN0(n5279), .IN1(n5278), .SEL(N15), .F(n5280) );
  MUX U5356 ( .IN0(\registers[26][10] ), .IN1(\registers[27][10] ), .SEL(N14), 
        .F(n5281) );
  MUX U5357 ( .IN0(\registers[24][10] ), .IN1(\registers[25][10] ), .SEL(N14), 
        .F(n5282) );
  MUX U5358 ( .IN0(n5282), .IN1(n5281), .SEL(N15), .F(n5283) );
  MUX U5359 ( .IN0(n5283), .IN1(n5280), .SEL(N16), .F(n5284) );
  MUX U5360 ( .IN0(\registers[22][10] ), .IN1(\registers[23][10] ), .SEL(N14), 
        .F(n5285) );
  MUX U5361 ( .IN0(\registers[20][10] ), .IN1(\registers[21][10] ), .SEL(N14), 
        .F(n5286) );
  MUX U5362 ( .IN0(n5286), .IN1(n5285), .SEL(N15), .F(n5287) );
  MUX U5363 ( .IN0(\registers[18][10] ), .IN1(\registers[19][10] ), .SEL(N14), 
        .F(n5288) );
  MUX U5364 ( .IN0(\registers[16][10] ), .IN1(\registers[17][10] ), .SEL(N14), 
        .F(n5289) );
  MUX U5365 ( .IN0(n5289), .IN1(n5288), .SEL(N15), .F(n5290) );
  MUX U5366 ( .IN0(n5290), .IN1(n5287), .SEL(N16), .F(n5291) );
  MUX U5367 ( .IN0(n5291), .IN1(n5284), .SEL(N17), .F(n5292) );
  MUX U5368 ( .IN0(\registers[14][10] ), .IN1(\registers[15][10] ), .SEL(N14), 
        .F(n5293) );
  MUX U5369 ( .IN0(\registers[12][10] ), .IN1(\registers[13][10] ), .SEL(N14), 
        .F(n5294) );
  MUX U5370 ( .IN0(n5294), .IN1(n5293), .SEL(N15), .F(n5295) );
  MUX U5371 ( .IN0(\registers[10][10] ), .IN1(\registers[11][10] ), .SEL(N14), 
        .F(n5296) );
  MUX U5372 ( .IN0(\registers[8][10] ), .IN1(\registers[9][10] ), .SEL(N14), 
        .F(n5297) );
  MUX U5373 ( .IN0(n5297), .IN1(n5296), .SEL(N15), .F(n5298) );
  MUX U5374 ( .IN0(n5298), .IN1(n5295), .SEL(N16), .F(n5299) );
  MUX U5375 ( .IN0(\registers[6][10] ), .IN1(\registers[7][10] ), .SEL(N14), 
        .F(n5300) );
  MUX U5376 ( .IN0(\registers[4][10] ), .IN1(\registers[5][10] ), .SEL(N14), 
        .F(n5301) );
  MUX U5377 ( .IN0(n5301), .IN1(n5300), .SEL(N15), .F(n5302) );
  MUX U5378 ( .IN0(\registers[2][10] ), .IN1(\registers[3][10] ), .SEL(N14), 
        .F(n5303) );
  MUX U5380 ( .IN0(n5304), .IN1(n5303), .SEL(N15), .F(n5305) );
  MUX U5381 ( .IN0(n5305), .IN1(n5302), .SEL(N16), .F(n5306) );
  MUX U5382 ( .IN0(n5306), .IN1(n5299), .SEL(N17), .F(n5307) );
  MUX U5383 ( .IN0(n5307), .IN1(n5292), .SEL(N18), .F(reg_target_out[10]) );
  MUX U5384 ( .IN0(\registers[30][11] ), .IN1(\registers[31][11] ), .SEL(N14), 
        .F(n5308) );
  MUX U5385 ( .IN0(\registers[28][11] ), .IN1(\registers[29][11] ), .SEL(N14), 
        .F(n5309) );
  MUX U5386 ( .IN0(n5309), .IN1(n5308), .SEL(N15), .F(n5310) );
  MUX U5387 ( .IN0(\registers[26][11] ), .IN1(\registers[27][11] ), .SEL(N14), 
        .F(n5311) );
  MUX U5388 ( .IN0(\registers[24][11] ), .IN1(\registers[25][11] ), .SEL(N14), 
        .F(n5312) );
  MUX U5389 ( .IN0(n5312), .IN1(n5311), .SEL(N15), .F(n5313) );
  MUX U5390 ( .IN0(n5313), .IN1(n5310), .SEL(N16), .F(n5314) );
  MUX U5391 ( .IN0(\registers[22][11] ), .IN1(\registers[23][11] ), .SEL(N14), 
        .F(n5315) );
  MUX U5392 ( .IN0(\registers[20][11] ), .IN1(\registers[21][11] ), .SEL(N14), 
        .F(n5316) );
  MUX U5393 ( .IN0(n5316), .IN1(n5315), .SEL(N15), .F(n5317) );
  MUX U5394 ( .IN0(\registers[18][11] ), .IN1(\registers[19][11] ), .SEL(N14), 
        .F(n5318) );
  MUX U5395 ( .IN0(\registers[16][11] ), .IN1(\registers[17][11] ), .SEL(N14), 
        .F(n5319) );
  MUX U5396 ( .IN0(n5319), .IN1(n5318), .SEL(N15), .F(n5320) );
  MUX U5397 ( .IN0(n5320), .IN1(n5317), .SEL(N16), .F(n5321) );
  MUX U5398 ( .IN0(n5321), .IN1(n5314), .SEL(N17), .F(n5322) );
  MUX U5399 ( .IN0(\registers[14][11] ), .IN1(\registers[15][11] ), .SEL(N14), 
        .F(n5323) );
  MUX U5400 ( .IN0(\registers[12][11] ), .IN1(\registers[13][11] ), .SEL(N14), 
        .F(n5324) );
  MUX U5401 ( .IN0(n5324), .IN1(n5323), .SEL(N15), .F(n5325) );
  MUX U5402 ( .IN0(\registers[10][11] ), .IN1(\registers[11][11] ), .SEL(N14), 
        .F(n5326) );
  MUX U5403 ( .IN0(\registers[8][11] ), .IN1(\registers[9][11] ), .SEL(N14), 
        .F(n5327) );
  MUX U5404 ( .IN0(n5327), .IN1(n5326), .SEL(N15), .F(n5328) );
  MUX U5405 ( .IN0(n5328), .IN1(n5325), .SEL(N16), .F(n5329) );
  MUX U5406 ( .IN0(\registers[6][11] ), .IN1(\registers[7][11] ), .SEL(N14), 
        .F(n5330) );
  MUX U5407 ( .IN0(\registers[4][11] ), .IN1(\registers[5][11] ), .SEL(N14), 
        .F(n5331) );
  MUX U5408 ( .IN0(n5331), .IN1(n5330), .SEL(N15), .F(n5332) );
  MUX U5409 ( .IN0(\registers[2][11] ), .IN1(\registers[3][11] ), .SEL(N14), 
        .F(n5333) );
  MUX U5411 ( .IN0(n5334), .IN1(n5333), .SEL(N15), .F(n5335) );
  MUX U5412 ( .IN0(n5335), .IN1(n5332), .SEL(N16), .F(n5336) );
  MUX U5413 ( .IN0(n5336), .IN1(n5329), .SEL(N17), .F(n5337) );
  MUX U5414 ( .IN0(n5337), .IN1(n5322), .SEL(N18), .F(reg_target_out[11]) );
  MUX U5415 ( .IN0(\registers[30][12] ), .IN1(\registers[31][12] ), .SEL(N14), 
        .F(n5338) );
  MUX U5416 ( .IN0(\registers[28][12] ), .IN1(\registers[29][12] ), .SEL(N14), 
        .F(n5339) );
  MUX U5417 ( .IN0(n5339), .IN1(n5338), .SEL(N15), .F(n5340) );
  MUX U5418 ( .IN0(\registers[26][12] ), .IN1(\registers[27][12] ), .SEL(N14), 
        .F(n5341) );
  MUX U5419 ( .IN0(\registers[24][12] ), .IN1(\registers[25][12] ), .SEL(N14), 
        .F(n5342) );
  MUX U5420 ( .IN0(n5342), .IN1(n5341), .SEL(N15), .F(n5343) );
  MUX U5421 ( .IN0(n5343), .IN1(n5340), .SEL(N16), .F(n5344) );
  MUX U5422 ( .IN0(\registers[22][12] ), .IN1(\registers[23][12] ), .SEL(N14), 
        .F(n5345) );
  MUX U5423 ( .IN0(\registers[20][12] ), .IN1(\registers[21][12] ), .SEL(N14), 
        .F(n5346) );
  MUX U5424 ( .IN0(n5346), .IN1(n5345), .SEL(N15), .F(n5347) );
  MUX U5425 ( .IN0(\registers[18][12] ), .IN1(\registers[19][12] ), .SEL(N14), 
        .F(n5348) );
  MUX U5426 ( .IN0(\registers[16][12] ), .IN1(\registers[17][12] ), .SEL(N14), 
        .F(n5349) );
  MUX U5427 ( .IN0(n5349), .IN1(n5348), .SEL(N15), .F(n5350) );
  MUX U5428 ( .IN0(n5350), .IN1(n5347), .SEL(N16), .F(n5351) );
  MUX U5429 ( .IN0(n5351), .IN1(n5344), .SEL(N17), .F(n5352) );
  MUX U5430 ( .IN0(\registers[14][12] ), .IN1(\registers[15][12] ), .SEL(N14), 
        .F(n5353) );
  MUX U5431 ( .IN0(\registers[12][12] ), .IN1(\registers[13][12] ), .SEL(N14), 
        .F(n5354) );
  MUX U5432 ( .IN0(n5354), .IN1(n5353), .SEL(N15), .F(n5355) );
  MUX U5433 ( .IN0(\registers[10][12] ), .IN1(\registers[11][12] ), .SEL(N14), 
        .F(n5356) );
  MUX U5434 ( .IN0(\registers[8][12] ), .IN1(\registers[9][12] ), .SEL(N14), 
        .F(n5357) );
  MUX U5435 ( .IN0(n5357), .IN1(n5356), .SEL(N15), .F(n5358) );
  MUX U5436 ( .IN0(n5358), .IN1(n5355), .SEL(N16), .F(n5359) );
  MUX U5437 ( .IN0(\registers[6][12] ), .IN1(\registers[7][12] ), .SEL(N14), 
        .F(n5360) );
  MUX U5438 ( .IN0(\registers[4][12] ), .IN1(\registers[5][12] ), .SEL(N14), 
        .F(n5361) );
  MUX U5439 ( .IN0(n5361), .IN1(n5360), .SEL(N15), .F(n5362) );
  MUX U5440 ( .IN0(\registers[2][12] ), .IN1(\registers[3][12] ), .SEL(N14), 
        .F(n5363) );
  MUX U5442 ( .IN0(n5364), .IN1(n5363), .SEL(N15), .F(n5365) );
  MUX U5443 ( .IN0(n5365), .IN1(n5362), .SEL(N16), .F(n5366) );
  MUX U5444 ( .IN0(n5366), .IN1(n5359), .SEL(N17), .F(n5367) );
  MUX U5445 ( .IN0(n5367), .IN1(n5352), .SEL(N18), .F(reg_target_out[12]) );
  MUX U5446 ( .IN0(\registers[30][13] ), .IN1(\registers[31][13] ), .SEL(N14), 
        .F(n5368) );
  MUX U5447 ( .IN0(\registers[28][13] ), .IN1(\registers[29][13] ), .SEL(N14), 
        .F(n5369) );
  MUX U5448 ( .IN0(n5369), .IN1(n5368), .SEL(N15), .F(n5370) );
  MUX U5449 ( .IN0(\registers[26][13] ), .IN1(\registers[27][13] ), .SEL(N14), 
        .F(n5371) );
  MUX U5450 ( .IN0(\registers[24][13] ), .IN1(\registers[25][13] ), .SEL(N14), 
        .F(n5372) );
  MUX U5451 ( .IN0(n5372), .IN1(n5371), .SEL(N15), .F(n5373) );
  MUX U5452 ( .IN0(n5373), .IN1(n5370), .SEL(N16), .F(n5374) );
  MUX U5453 ( .IN0(\registers[22][13] ), .IN1(\registers[23][13] ), .SEL(N14), 
        .F(n5375) );
  MUX U5454 ( .IN0(\registers[20][13] ), .IN1(\registers[21][13] ), .SEL(N14), 
        .F(n5376) );
  MUX U5455 ( .IN0(n5376), .IN1(n5375), .SEL(N15), .F(n5377) );
  MUX U5456 ( .IN0(\registers[18][13] ), .IN1(\registers[19][13] ), .SEL(N14), 
        .F(n5378) );
  MUX U5457 ( .IN0(\registers[16][13] ), .IN1(\registers[17][13] ), .SEL(N14), 
        .F(n5379) );
  MUX U5458 ( .IN0(n5379), .IN1(n5378), .SEL(N15), .F(n5380) );
  MUX U5459 ( .IN0(n5380), .IN1(n5377), .SEL(N16), .F(n5381) );
  MUX U5460 ( .IN0(n5381), .IN1(n5374), .SEL(N17), .F(n5382) );
  MUX U5461 ( .IN0(\registers[14][13] ), .IN1(\registers[15][13] ), .SEL(N14), 
        .F(n5383) );
  MUX U5462 ( .IN0(\registers[12][13] ), .IN1(\registers[13][13] ), .SEL(N14), 
        .F(n5384) );
  MUX U5463 ( .IN0(n5384), .IN1(n5383), .SEL(N15), .F(n5385) );
  MUX U5464 ( .IN0(\registers[10][13] ), .IN1(\registers[11][13] ), .SEL(N14), 
        .F(n5386) );
  MUX U5465 ( .IN0(\registers[8][13] ), .IN1(\registers[9][13] ), .SEL(N14), 
        .F(n5387) );
  MUX U5466 ( .IN0(n5387), .IN1(n5386), .SEL(N15), .F(n5388) );
  MUX U5467 ( .IN0(n5388), .IN1(n5385), .SEL(N16), .F(n5389) );
  MUX U5468 ( .IN0(\registers[6][13] ), .IN1(\registers[7][13] ), .SEL(N14), 
        .F(n5390) );
  MUX U5469 ( .IN0(\registers[4][13] ), .IN1(\registers[5][13] ), .SEL(N14), 
        .F(n5391) );
  MUX U5470 ( .IN0(n5391), .IN1(n5390), .SEL(N15), .F(n5392) );
  MUX U5471 ( .IN0(\registers[2][13] ), .IN1(\registers[3][13] ), .SEL(N14), 
        .F(n5393) );
  MUX U5473 ( .IN0(n5394), .IN1(n5393), .SEL(N15), .F(n5395) );
  MUX U5474 ( .IN0(n5395), .IN1(n5392), .SEL(N16), .F(n5396) );
  MUX U5475 ( .IN0(n5396), .IN1(n5389), .SEL(N17), .F(n5397) );
  MUX U5476 ( .IN0(n5397), .IN1(n5382), .SEL(N18), .F(reg_target_out[13]) );
  MUX U5477 ( .IN0(\registers[30][14] ), .IN1(\registers[31][14] ), .SEL(N14), 
        .F(n5398) );
  MUX U5478 ( .IN0(\registers[28][14] ), .IN1(\registers[29][14] ), .SEL(N14), 
        .F(n5399) );
  MUX U5479 ( .IN0(n5399), .IN1(n5398), .SEL(N15), .F(n5400) );
  MUX U5480 ( .IN0(\registers[26][14] ), .IN1(\registers[27][14] ), .SEL(N14), 
        .F(n5401) );
  MUX U5481 ( .IN0(\registers[24][14] ), .IN1(\registers[25][14] ), .SEL(N14), 
        .F(n5402) );
  MUX U5482 ( .IN0(n5402), .IN1(n5401), .SEL(N15), .F(n5403) );
  MUX U5483 ( .IN0(n5403), .IN1(n5400), .SEL(N16), .F(n5404) );
  MUX U5484 ( .IN0(\registers[22][14] ), .IN1(\registers[23][14] ), .SEL(N14), 
        .F(n5405) );
  MUX U5485 ( .IN0(\registers[20][14] ), .IN1(\registers[21][14] ), .SEL(N14), 
        .F(n5406) );
  MUX U5486 ( .IN0(n5406), .IN1(n5405), .SEL(N15), .F(n5407) );
  MUX U5487 ( .IN0(\registers[18][14] ), .IN1(\registers[19][14] ), .SEL(N14), 
        .F(n5408) );
  MUX U5488 ( .IN0(\registers[16][14] ), .IN1(\registers[17][14] ), .SEL(N14), 
        .F(n5409) );
  MUX U5489 ( .IN0(n5409), .IN1(n5408), .SEL(N15), .F(n5410) );
  MUX U5490 ( .IN0(n5410), .IN1(n5407), .SEL(N16), .F(n5411) );
  MUX U5491 ( .IN0(n5411), .IN1(n5404), .SEL(N17), .F(n5412) );
  MUX U5492 ( .IN0(\registers[14][14] ), .IN1(\registers[15][14] ), .SEL(N14), 
        .F(n5413) );
  MUX U5493 ( .IN0(\registers[12][14] ), .IN1(\registers[13][14] ), .SEL(N14), 
        .F(n5414) );
  MUX U5494 ( .IN0(n5414), .IN1(n5413), .SEL(N15), .F(n5415) );
  MUX U5495 ( .IN0(\registers[10][14] ), .IN1(\registers[11][14] ), .SEL(N14), 
        .F(n5416) );
  MUX U5496 ( .IN0(\registers[8][14] ), .IN1(\registers[9][14] ), .SEL(N14), 
        .F(n5417) );
  MUX U5497 ( .IN0(n5417), .IN1(n5416), .SEL(N15), .F(n5418) );
  MUX U5498 ( .IN0(n5418), .IN1(n5415), .SEL(N16), .F(n5419) );
  MUX U5499 ( .IN0(\registers[6][14] ), .IN1(\registers[7][14] ), .SEL(N14), 
        .F(n5420) );
  MUX U5500 ( .IN0(\registers[4][14] ), .IN1(\registers[5][14] ), .SEL(N14), 
        .F(n5421) );
  MUX U5501 ( .IN0(n5421), .IN1(n5420), .SEL(N15), .F(n5422) );
  MUX U5502 ( .IN0(\registers[2][14] ), .IN1(\registers[3][14] ), .SEL(N14), 
        .F(n5423) );
  MUX U5504 ( .IN0(n5424), .IN1(n5423), .SEL(N15), .F(n5425) );
  MUX U5505 ( .IN0(n5425), .IN1(n5422), .SEL(N16), .F(n5426) );
  MUX U5506 ( .IN0(n5426), .IN1(n5419), .SEL(N17), .F(n5427) );
  MUX U5507 ( .IN0(n5427), .IN1(n5412), .SEL(N18), .F(reg_target_out[14]) );
  MUX U5508 ( .IN0(\registers[30][15] ), .IN1(\registers[31][15] ), .SEL(N14), 
        .F(n5428) );
  MUX U5509 ( .IN0(\registers[28][15] ), .IN1(\registers[29][15] ), .SEL(N14), 
        .F(n5429) );
  MUX U5510 ( .IN0(n5429), .IN1(n5428), .SEL(N15), .F(n5430) );
  MUX U5511 ( .IN0(\registers[26][15] ), .IN1(\registers[27][15] ), .SEL(N14), 
        .F(n5431) );
  MUX U5512 ( .IN0(\registers[24][15] ), .IN1(\registers[25][15] ), .SEL(N14), 
        .F(n5432) );
  MUX U5513 ( .IN0(n5432), .IN1(n5431), .SEL(N15), .F(n5433) );
  MUX U5514 ( .IN0(n5433), .IN1(n5430), .SEL(N16), .F(n5434) );
  MUX U5515 ( .IN0(\registers[22][15] ), .IN1(\registers[23][15] ), .SEL(N14), 
        .F(n5435) );
  MUX U5516 ( .IN0(\registers[20][15] ), .IN1(\registers[21][15] ), .SEL(N14), 
        .F(n5436) );
  MUX U5517 ( .IN0(n5436), .IN1(n5435), .SEL(N15), .F(n5437) );
  MUX U5518 ( .IN0(\registers[18][15] ), .IN1(\registers[19][15] ), .SEL(N14), 
        .F(n5438) );
  MUX U5519 ( .IN0(\registers[16][15] ), .IN1(\registers[17][15] ), .SEL(N14), 
        .F(n5439) );
  MUX U5520 ( .IN0(n5439), .IN1(n5438), .SEL(N15), .F(n5440) );
  MUX U5521 ( .IN0(n5440), .IN1(n5437), .SEL(N16), .F(n5441) );
  MUX U5522 ( .IN0(n5441), .IN1(n5434), .SEL(N17), .F(n5442) );
  MUX U5523 ( .IN0(\registers[14][15] ), .IN1(\registers[15][15] ), .SEL(N14), 
        .F(n5443) );
  MUX U5524 ( .IN0(\registers[12][15] ), .IN1(\registers[13][15] ), .SEL(N14), 
        .F(n5444) );
  MUX U5525 ( .IN0(n5444), .IN1(n5443), .SEL(N15), .F(n5445) );
  MUX U5526 ( .IN0(\registers[10][15] ), .IN1(\registers[11][15] ), .SEL(N14), 
        .F(n5446) );
  MUX U5527 ( .IN0(\registers[8][15] ), .IN1(\registers[9][15] ), .SEL(N14), 
        .F(n5447) );
  MUX U5528 ( .IN0(n5447), .IN1(n5446), .SEL(N15), .F(n5448) );
  MUX U5529 ( .IN0(n5448), .IN1(n5445), .SEL(N16), .F(n5449) );
  MUX U5530 ( .IN0(\registers[6][15] ), .IN1(\registers[7][15] ), .SEL(N14), 
        .F(n5450) );
  MUX U5531 ( .IN0(\registers[4][15] ), .IN1(\registers[5][15] ), .SEL(N14), 
        .F(n5451) );
  MUX U5532 ( .IN0(n5451), .IN1(n5450), .SEL(N15), .F(n5452) );
  MUX U5533 ( .IN0(\registers[2][15] ), .IN1(\registers[3][15] ), .SEL(N14), 
        .F(n5453) );
  MUX U5535 ( .IN0(n5454), .IN1(n5453), .SEL(N15), .F(n5455) );
  MUX U5536 ( .IN0(n5455), .IN1(n5452), .SEL(N16), .F(n5456) );
  MUX U5537 ( .IN0(n5456), .IN1(n5449), .SEL(N17), .F(n5457) );
  MUX U5538 ( .IN0(n5457), .IN1(n5442), .SEL(N18), .F(reg_target_out[15]) );
  MUX U5539 ( .IN0(\registers[30][16] ), .IN1(\registers[31][16] ), .SEL(N14), 
        .F(n5458) );
  MUX U5540 ( .IN0(\registers[28][16] ), .IN1(\registers[29][16] ), .SEL(N14), 
        .F(n5459) );
  MUX U5541 ( .IN0(n5459), .IN1(n5458), .SEL(N15), .F(n5460) );
  MUX U5542 ( .IN0(\registers[26][16] ), .IN1(\registers[27][16] ), .SEL(N14), 
        .F(n5461) );
  MUX U5543 ( .IN0(\registers[24][16] ), .IN1(\registers[25][16] ), .SEL(N14), 
        .F(n5462) );
  MUX U5544 ( .IN0(n5462), .IN1(n5461), .SEL(N15), .F(n5463) );
  MUX U5545 ( .IN0(n5463), .IN1(n5460), .SEL(N16), .F(n5464) );
  MUX U5546 ( .IN0(\registers[22][16] ), .IN1(\registers[23][16] ), .SEL(N14), 
        .F(n5465) );
  MUX U5547 ( .IN0(\registers[20][16] ), .IN1(\registers[21][16] ), .SEL(N14), 
        .F(n5466) );
  MUX U5548 ( .IN0(n5466), .IN1(n5465), .SEL(N15), .F(n5467) );
  MUX U5549 ( .IN0(\registers[18][16] ), .IN1(\registers[19][16] ), .SEL(N14), 
        .F(n5468) );
  MUX U5550 ( .IN0(\registers[16][16] ), .IN1(\registers[17][16] ), .SEL(N14), 
        .F(n5469) );
  MUX U5551 ( .IN0(n5469), .IN1(n5468), .SEL(N15), .F(n5470) );
  MUX U5552 ( .IN0(n5470), .IN1(n5467), .SEL(N16), .F(n5471) );
  MUX U5553 ( .IN0(n5471), .IN1(n5464), .SEL(N17), .F(n5472) );
  MUX U5554 ( .IN0(\registers[14][16] ), .IN1(\registers[15][16] ), .SEL(N14), 
        .F(n5473) );
  MUX U5555 ( .IN0(\registers[12][16] ), .IN1(\registers[13][16] ), .SEL(N14), 
        .F(n5474) );
  MUX U5556 ( .IN0(n5474), .IN1(n5473), .SEL(N15), .F(n5475) );
  MUX U5557 ( .IN0(\registers[10][16] ), .IN1(\registers[11][16] ), .SEL(N14), 
        .F(n5476) );
  MUX U5558 ( .IN0(\registers[8][16] ), .IN1(\registers[9][16] ), .SEL(N14), 
        .F(n5477) );
  MUX U5559 ( .IN0(n5477), .IN1(n5476), .SEL(N15), .F(n5478) );
  MUX U5560 ( .IN0(n5478), .IN1(n5475), .SEL(N16), .F(n5479) );
  MUX U5561 ( .IN0(\registers[6][16] ), .IN1(\registers[7][16] ), .SEL(N14), 
        .F(n5480) );
  MUX U5562 ( .IN0(\registers[4][16] ), .IN1(\registers[5][16] ), .SEL(N14), 
        .F(n5481) );
  MUX U5563 ( .IN0(n5481), .IN1(n5480), .SEL(N15), .F(n5482) );
  MUX U5564 ( .IN0(\registers[2][16] ), .IN1(\registers[3][16] ), .SEL(N14), 
        .F(n5483) );
  MUX U5566 ( .IN0(n5484), .IN1(n5483), .SEL(N15), .F(n5485) );
  MUX U5567 ( .IN0(n5485), .IN1(n5482), .SEL(N16), .F(n5486) );
  MUX U5568 ( .IN0(n5486), .IN1(n5479), .SEL(N17), .F(n5487) );
  MUX U5569 ( .IN0(n5487), .IN1(n5472), .SEL(N18), .F(reg_target_out[16]) );
  MUX U5570 ( .IN0(\registers[30][17] ), .IN1(\registers[31][17] ), .SEL(N14), 
        .F(n5488) );
  MUX U5571 ( .IN0(\registers[28][17] ), .IN1(\registers[29][17] ), .SEL(N14), 
        .F(n5489) );
  MUX U5572 ( .IN0(n5489), .IN1(n5488), .SEL(N15), .F(n5490) );
  MUX U5573 ( .IN0(\registers[26][17] ), .IN1(\registers[27][17] ), .SEL(N14), 
        .F(n5491) );
  MUX U5574 ( .IN0(\registers[24][17] ), .IN1(\registers[25][17] ), .SEL(N14), 
        .F(n5492) );
  MUX U5575 ( .IN0(n5492), .IN1(n5491), .SEL(N15), .F(n5493) );
  MUX U5576 ( .IN0(n5493), .IN1(n5490), .SEL(N16), .F(n5494) );
  MUX U5577 ( .IN0(\registers[22][17] ), .IN1(\registers[23][17] ), .SEL(N14), 
        .F(n5495) );
  MUX U5578 ( .IN0(\registers[20][17] ), .IN1(\registers[21][17] ), .SEL(N14), 
        .F(n5496) );
  MUX U5579 ( .IN0(n5496), .IN1(n5495), .SEL(N15), .F(n5497) );
  MUX U5580 ( .IN0(\registers[18][17] ), .IN1(\registers[19][17] ), .SEL(N14), 
        .F(n5498) );
  MUX U5581 ( .IN0(\registers[16][17] ), .IN1(\registers[17][17] ), .SEL(N14), 
        .F(n5499) );
  MUX U5582 ( .IN0(n5499), .IN1(n5498), .SEL(N15), .F(n5500) );
  MUX U5583 ( .IN0(n5500), .IN1(n5497), .SEL(N16), .F(n5501) );
  MUX U5584 ( .IN0(n5501), .IN1(n5494), .SEL(N17), .F(n5502) );
  MUX U5585 ( .IN0(\registers[14][17] ), .IN1(\registers[15][17] ), .SEL(N14), 
        .F(n5503) );
  MUX U5586 ( .IN0(\registers[12][17] ), .IN1(\registers[13][17] ), .SEL(N14), 
        .F(n5504) );
  MUX U5587 ( .IN0(n5504), .IN1(n5503), .SEL(N15), .F(n5505) );
  MUX U5588 ( .IN0(\registers[10][17] ), .IN1(\registers[11][17] ), .SEL(N14), 
        .F(n5506) );
  MUX U5589 ( .IN0(\registers[8][17] ), .IN1(\registers[9][17] ), .SEL(N14), 
        .F(n5507) );
  MUX U5590 ( .IN0(n5507), .IN1(n5506), .SEL(N15), .F(n5508) );
  MUX U5591 ( .IN0(n5508), .IN1(n5505), .SEL(N16), .F(n5509) );
  MUX U5592 ( .IN0(\registers[6][17] ), .IN1(\registers[7][17] ), .SEL(N14), 
        .F(n5510) );
  MUX U5593 ( .IN0(\registers[4][17] ), .IN1(\registers[5][17] ), .SEL(N14), 
        .F(n5511) );
  MUX U5594 ( .IN0(n5511), .IN1(n5510), .SEL(N15), .F(n5512) );
  MUX U5595 ( .IN0(\registers[2][17] ), .IN1(\registers[3][17] ), .SEL(N14), 
        .F(n5513) );
  MUX U5597 ( .IN0(n5514), .IN1(n5513), .SEL(N15), .F(n5515) );
  MUX U5598 ( .IN0(n5515), .IN1(n5512), .SEL(N16), .F(n5516) );
  MUX U5599 ( .IN0(n5516), .IN1(n5509), .SEL(N17), .F(n5517) );
  MUX U5600 ( .IN0(n5517), .IN1(n5502), .SEL(N18), .F(reg_target_out[17]) );
  MUX U5601 ( .IN0(\registers[30][18] ), .IN1(\registers[31][18] ), .SEL(N14), 
        .F(n5518) );
  MUX U5602 ( .IN0(\registers[28][18] ), .IN1(\registers[29][18] ), .SEL(N14), 
        .F(n5519) );
  MUX U5603 ( .IN0(n5519), .IN1(n5518), .SEL(N15), .F(n5520) );
  MUX U5604 ( .IN0(\registers[26][18] ), .IN1(\registers[27][18] ), .SEL(N14), 
        .F(n5521) );
  MUX U5605 ( .IN0(\registers[24][18] ), .IN1(\registers[25][18] ), .SEL(N14), 
        .F(n5522) );
  MUX U5606 ( .IN0(n5522), .IN1(n5521), .SEL(N15), .F(n5523) );
  MUX U5607 ( .IN0(n5523), .IN1(n5520), .SEL(N16), .F(n5524) );
  MUX U5608 ( .IN0(\registers[22][18] ), .IN1(\registers[23][18] ), .SEL(N14), 
        .F(n5525) );
  MUX U5609 ( .IN0(\registers[20][18] ), .IN1(\registers[21][18] ), .SEL(N14), 
        .F(n5526) );
  MUX U5610 ( .IN0(n5526), .IN1(n5525), .SEL(N15), .F(n5527) );
  MUX U5611 ( .IN0(\registers[18][18] ), .IN1(\registers[19][18] ), .SEL(N14), 
        .F(n5528) );
  MUX U5612 ( .IN0(\registers[16][18] ), .IN1(\registers[17][18] ), .SEL(N14), 
        .F(n5529) );
  MUX U5613 ( .IN0(n5529), .IN1(n5528), .SEL(N15), .F(n5530) );
  MUX U5614 ( .IN0(n5530), .IN1(n5527), .SEL(N16), .F(n5531) );
  MUX U5615 ( .IN0(n5531), .IN1(n5524), .SEL(N17), .F(n5532) );
  MUX U5616 ( .IN0(\registers[14][18] ), .IN1(\registers[15][18] ), .SEL(N14), 
        .F(n5533) );
  MUX U5617 ( .IN0(\registers[12][18] ), .IN1(\registers[13][18] ), .SEL(N14), 
        .F(n5534) );
  MUX U5618 ( .IN0(n5534), .IN1(n5533), .SEL(N15), .F(n5535) );
  MUX U5619 ( .IN0(\registers[10][18] ), .IN1(\registers[11][18] ), .SEL(N14), 
        .F(n5536) );
  MUX U5620 ( .IN0(\registers[8][18] ), .IN1(\registers[9][18] ), .SEL(N14), 
        .F(n5537) );
  MUX U5621 ( .IN0(n5537), .IN1(n5536), .SEL(N15), .F(n5538) );
  MUX U5622 ( .IN0(n5538), .IN1(n5535), .SEL(N16), .F(n5539) );
  MUX U5623 ( .IN0(\registers[6][18] ), .IN1(\registers[7][18] ), .SEL(N14), 
        .F(n5540) );
  MUX U5624 ( .IN0(\registers[4][18] ), .IN1(\registers[5][18] ), .SEL(N14), 
        .F(n5541) );
  MUX U5625 ( .IN0(n5541), .IN1(n5540), .SEL(N15), .F(n5542) );
  MUX U5626 ( .IN0(\registers[2][18] ), .IN1(\registers[3][18] ), .SEL(N14), 
        .F(n5543) );
  MUX U5628 ( .IN0(n5544), .IN1(n5543), .SEL(N15), .F(n5545) );
  MUX U5629 ( .IN0(n5545), .IN1(n5542), .SEL(N16), .F(n5546) );
  MUX U5630 ( .IN0(n5546), .IN1(n5539), .SEL(N17), .F(n5547) );
  MUX U5631 ( .IN0(n5547), .IN1(n5532), .SEL(N18), .F(reg_target_out[18]) );
  MUX U5632 ( .IN0(\registers[30][19] ), .IN1(\registers[31][19] ), .SEL(N14), 
        .F(n5548) );
  MUX U5633 ( .IN0(\registers[28][19] ), .IN1(\registers[29][19] ), .SEL(N14), 
        .F(n5549) );
  MUX U5634 ( .IN0(n5549), .IN1(n5548), .SEL(N15), .F(n5550) );
  MUX U5635 ( .IN0(\registers[26][19] ), .IN1(\registers[27][19] ), .SEL(N14), 
        .F(n5551) );
  MUX U5636 ( .IN0(\registers[24][19] ), .IN1(\registers[25][19] ), .SEL(N14), 
        .F(n5552) );
  MUX U5637 ( .IN0(n5552), .IN1(n5551), .SEL(N15), .F(n5553) );
  MUX U5638 ( .IN0(n5553), .IN1(n5550), .SEL(N16), .F(n5554) );
  MUX U5639 ( .IN0(\registers[22][19] ), .IN1(\registers[23][19] ), .SEL(N14), 
        .F(n5555) );
  MUX U5640 ( .IN0(\registers[20][19] ), .IN1(\registers[21][19] ), .SEL(N14), 
        .F(n5556) );
  MUX U5641 ( .IN0(n5556), .IN1(n5555), .SEL(N15), .F(n5557) );
  MUX U5642 ( .IN0(\registers[18][19] ), .IN1(\registers[19][19] ), .SEL(N14), 
        .F(n5558) );
  MUX U5643 ( .IN0(\registers[16][19] ), .IN1(\registers[17][19] ), .SEL(N14), 
        .F(n5559) );
  MUX U5644 ( .IN0(n5559), .IN1(n5558), .SEL(N15), .F(n5560) );
  MUX U5645 ( .IN0(n5560), .IN1(n5557), .SEL(N16), .F(n5561) );
  MUX U5646 ( .IN0(n5561), .IN1(n5554), .SEL(N17), .F(n5562) );
  MUX U5647 ( .IN0(\registers[14][19] ), .IN1(\registers[15][19] ), .SEL(N14), 
        .F(n5563) );
  MUX U5648 ( .IN0(\registers[12][19] ), .IN1(\registers[13][19] ), .SEL(N14), 
        .F(n5564) );
  MUX U5649 ( .IN0(n5564), .IN1(n5563), .SEL(N15), .F(n5565) );
  MUX U5650 ( .IN0(\registers[10][19] ), .IN1(\registers[11][19] ), .SEL(N14), 
        .F(n5566) );
  MUX U5651 ( .IN0(\registers[8][19] ), .IN1(\registers[9][19] ), .SEL(N14), 
        .F(n5567) );
  MUX U5652 ( .IN0(n5567), .IN1(n5566), .SEL(N15), .F(n5568) );
  MUX U5653 ( .IN0(n5568), .IN1(n5565), .SEL(N16), .F(n5569) );
  MUX U5654 ( .IN0(\registers[6][19] ), .IN1(\registers[7][19] ), .SEL(N14), 
        .F(n5570) );
  MUX U5655 ( .IN0(\registers[4][19] ), .IN1(\registers[5][19] ), .SEL(N14), 
        .F(n5571) );
  MUX U5656 ( .IN0(n5571), .IN1(n5570), .SEL(N15), .F(n5572) );
  MUX U5657 ( .IN0(\registers[2][19] ), .IN1(\registers[3][19] ), .SEL(N14), 
        .F(n5573) );
  MUX U5659 ( .IN0(n5574), .IN1(n5573), .SEL(N15), .F(n5575) );
  MUX U5660 ( .IN0(n5575), .IN1(n5572), .SEL(N16), .F(n5576) );
  MUX U5661 ( .IN0(n5576), .IN1(n5569), .SEL(N17), .F(n5577) );
  MUX U5662 ( .IN0(n5577), .IN1(n5562), .SEL(N18), .F(reg_target_out[19]) );
  MUX U5663 ( .IN0(\registers[30][20] ), .IN1(\registers[31][20] ), .SEL(N14), 
        .F(n5578) );
  MUX U5664 ( .IN0(\registers[28][20] ), .IN1(\registers[29][20] ), .SEL(N14), 
        .F(n5579) );
  MUX U5665 ( .IN0(n5579), .IN1(n5578), .SEL(N15), .F(n5580) );
  MUX U5666 ( .IN0(\registers[26][20] ), .IN1(\registers[27][20] ), .SEL(N14), 
        .F(n5581) );
  MUX U5667 ( .IN0(\registers[24][20] ), .IN1(\registers[25][20] ), .SEL(N14), 
        .F(n5582) );
  MUX U5668 ( .IN0(n5582), .IN1(n5581), .SEL(N15), .F(n5583) );
  MUX U5669 ( .IN0(n5583), .IN1(n5580), .SEL(N16), .F(n5584) );
  MUX U5670 ( .IN0(\registers[22][20] ), .IN1(\registers[23][20] ), .SEL(N14), 
        .F(n5585) );
  MUX U5671 ( .IN0(\registers[20][20] ), .IN1(\registers[21][20] ), .SEL(N14), 
        .F(n5586) );
  MUX U5672 ( .IN0(n5586), .IN1(n5585), .SEL(N15), .F(n5587) );
  MUX U5673 ( .IN0(\registers[18][20] ), .IN1(\registers[19][20] ), .SEL(N14), 
        .F(n5588) );
  MUX U5674 ( .IN0(\registers[16][20] ), .IN1(\registers[17][20] ), .SEL(N14), 
        .F(n5589) );
  MUX U5675 ( .IN0(n5589), .IN1(n5588), .SEL(N15), .F(n5590) );
  MUX U5676 ( .IN0(n5590), .IN1(n5587), .SEL(N16), .F(n5591) );
  MUX U5677 ( .IN0(n5591), .IN1(n5584), .SEL(N17), .F(n5592) );
  MUX U5678 ( .IN0(\registers[14][20] ), .IN1(\registers[15][20] ), .SEL(N14), 
        .F(n5593) );
  MUX U5679 ( .IN0(\registers[12][20] ), .IN1(\registers[13][20] ), .SEL(N14), 
        .F(n5594) );
  MUX U5680 ( .IN0(n5594), .IN1(n5593), .SEL(N15), .F(n5595) );
  MUX U5681 ( .IN0(\registers[10][20] ), .IN1(\registers[11][20] ), .SEL(N14), 
        .F(n5596) );
  MUX U5682 ( .IN0(\registers[8][20] ), .IN1(\registers[9][20] ), .SEL(N14), 
        .F(n5597) );
  MUX U5683 ( .IN0(n5597), .IN1(n5596), .SEL(N15), .F(n5598) );
  MUX U5684 ( .IN0(n5598), .IN1(n5595), .SEL(N16), .F(n5599) );
  MUX U5685 ( .IN0(\registers[6][20] ), .IN1(\registers[7][20] ), .SEL(N14), 
        .F(n5600) );
  MUX U5686 ( .IN0(\registers[4][20] ), .IN1(\registers[5][20] ), .SEL(N14), 
        .F(n5601) );
  MUX U5687 ( .IN0(n5601), .IN1(n5600), .SEL(N15), .F(n5602) );
  MUX U5688 ( .IN0(\registers[2][20] ), .IN1(\registers[3][20] ), .SEL(N14), 
        .F(n5603) );
  MUX U5690 ( .IN0(n5604), .IN1(n5603), .SEL(N15), .F(n5605) );
  MUX U5691 ( .IN0(n5605), .IN1(n5602), .SEL(N16), .F(n5606) );
  MUX U5692 ( .IN0(n5606), .IN1(n5599), .SEL(N17), .F(n5607) );
  MUX U5693 ( .IN0(n5607), .IN1(n5592), .SEL(N18), .F(reg_target_out[20]) );
  MUX U5694 ( .IN0(\registers[30][21] ), .IN1(\registers[31][21] ), .SEL(N14), 
        .F(n5608) );
  MUX U5695 ( .IN0(\registers[28][21] ), .IN1(\registers[29][21] ), .SEL(N14), 
        .F(n5609) );
  MUX U5696 ( .IN0(n5609), .IN1(n5608), .SEL(N15), .F(n5610) );
  MUX U5697 ( .IN0(\registers[26][21] ), .IN1(\registers[27][21] ), .SEL(N14), 
        .F(n5611) );
  MUX U5698 ( .IN0(\registers[24][21] ), .IN1(\registers[25][21] ), .SEL(N14), 
        .F(n5612) );
  MUX U5699 ( .IN0(n5612), .IN1(n5611), .SEL(N15), .F(n5613) );
  MUX U5700 ( .IN0(n5613), .IN1(n5610), .SEL(N16), .F(n5614) );
  MUX U5701 ( .IN0(\registers[22][21] ), .IN1(\registers[23][21] ), .SEL(N14), 
        .F(n5615) );
  MUX U5702 ( .IN0(\registers[20][21] ), .IN1(\registers[21][21] ), .SEL(N14), 
        .F(n5616) );
  MUX U5703 ( .IN0(n5616), .IN1(n5615), .SEL(N15), .F(n5617) );
  MUX U5704 ( .IN0(\registers[18][21] ), .IN1(\registers[19][21] ), .SEL(N14), 
        .F(n5618) );
  MUX U5705 ( .IN0(\registers[16][21] ), .IN1(\registers[17][21] ), .SEL(N14), 
        .F(n5619) );
  MUX U5706 ( .IN0(n5619), .IN1(n5618), .SEL(N15), .F(n5620) );
  MUX U5707 ( .IN0(n5620), .IN1(n5617), .SEL(N16), .F(n5621) );
  MUX U5708 ( .IN0(n5621), .IN1(n5614), .SEL(N17), .F(n5622) );
  MUX U5709 ( .IN0(\registers[14][21] ), .IN1(\registers[15][21] ), .SEL(N14), 
        .F(n5623) );
  MUX U5710 ( .IN0(\registers[12][21] ), .IN1(\registers[13][21] ), .SEL(N14), 
        .F(n5624) );
  MUX U5711 ( .IN0(n5624), .IN1(n5623), .SEL(N15), .F(n5625) );
  MUX U5712 ( .IN0(\registers[10][21] ), .IN1(\registers[11][21] ), .SEL(N14), 
        .F(n5626) );
  MUX U5713 ( .IN0(\registers[8][21] ), .IN1(\registers[9][21] ), .SEL(N14), 
        .F(n5627) );
  MUX U5714 ( .IN0(n5627), .IN1(n5626), .SEL(N15), .F(n5628) );
  MUX U5715 ( .IN0(n5628), .IN1(n5625), .SEL(N16), .F(n5629) );
  MUX U5716 ( .IN0(\registers[6][21] ), .IN1(\registers[7][21] ), .SEL(N14), 
        .F(n5630) );
  MUX U5717 ( .IN0(\registers[4][21] ), .IN1(\registers[5][21] ), .SEL(N14), 
        .F(n5631) );
  MUX U5718 ( .IN0(n5631), .IN1(n5630), .SEL(N15), .F(n5632) );
  MUX U5719 ( .IN0(\registers[2][21] ), .IN1(\registers[3][21] ), .SEL(N14), 
        .F(n5633) );
  MUX U5721 ( .IN0(n5634), .IN1(n5633), .SEL(N15), .F(n5635) );
  MUX U5722 ( .IN0(n5635), .IN1(n5632), .SEL(N16), .F(n5636) );
  MUX U5723 ( .IN0(n5636), .IN1(n5629), .SEL(N17), .F(n5637) );
  MUX U5724 ( .IN0(n5637), .IN1(n5622), .SEL(N18), .F(reg_target_out[21]) );
  MUX U5725 ( .IN0(\registers[30][22] ), .IN1(\registers[31][22] ), .SEL(N14), 
        .F(n5638) );
  MUX U5726 ( .IN0(\registers[28][22] ), .IN1(\registers[29][22] ), .SEL(N14), 
        .F(n5639) );
  MUX U5727 ( .IN0(n5639), .IN1(n5638), .SEL(N15), .F(n5640) );
  MUX U5728 ( .IN0(\registers[26][22] ), .IN1(\registers[27][22] ), .SEL(N14), 
        .F(n5641) );
  MUX U5729 ( .IN0(\registers[24][22] ), .IN1(\registers[25][22] ), .SEL(N14), 
        .F(n5642) );
  MUX U5730 ( .IN0(n5642), .IN1(n5641), .SEL(N15), .F(n5643) );
  MUX U5731 ( .IN0(n5643), .IN1(n5640), .SEL(N16), .F(n5644) );
  MUX U5732 ( .IN0(\registers[22][22] ), .IN1(\registers[23][22] ), .SEL(N14), 
        .F(n5645) );
  MUX U5733 ( .IN0(\registers[20][22] ), .IN1(\registers[21][22] ), .SEL(N14), 
        .F(n5646) );
  MUX U5734 ( .IN0(n5646), .IN1(n5645), .SEL(N15), .F(n5647) );
  MUX U5735 ( .IN0(\registers[18][22] ), .IN1(\registers[19][22] ), .SEL(N14), 
        .F(n5648) );
  MUX U5736 ( .IN0(\registers[16][22] ), .IN1(\registers[17][22] ), .SEL(N14), 
        .F(n5649) );
  MUX U5737 ( .IN0(n5649), .IN1(n5648), .SEL(N15), .F(n5650) );
  MUX U5738 ( .IN0(n5650), .IN1(n5647), .SEL(N16), .F(n5651) );
  MUX U5739 ( .IN0(n5651), .IN1(n5644), .SEL(N17), .F(n5652) );
  MUX U5740 ( .IN0(\registers[14][22] ), .IN1(\registers[15][22] ), .SEL(N14), 
        .F(n5653) );
  MUX U5741 ( .IN0(\registers[12][22] ), .IN1(\registers[13][22] ), .SEL(N14), 
        .F(n5654) );
  MUX U5742 ( .IN0(n5654), .IN1(n5653), .SEL(N15), .F(n5655) );
  MUX U5743 ( .IN0(\registers[10][22] ), .IN1(\registers[11][22] ), .SEL(N14), 
        .F(n5656) );
  MUX U5744 ( .IN0(\registers[8][22] ), .IN1(\registers[9][22] ), .SEL(N14), 
        .F(n5657) );
  MUX U5745 ( .IN0(n5657), .IN1(n5656), .SEL(N15), .F(n5658) );
  MUX U5746 ( .IN0(n5658), .IN1(n5655), .SEL(N16), .F(n5659) );
  MUX U5747 ( .IN0(\registers[6][22] ), .IN1(\registers[7][22] ), .SEL(N14), 
        .F(n5660) );
  MUX U5748 ( .IN0(\registers[4][22] ), .IN1(\registers[5][22] ), .SEL(N14), 
        .F(n5661) );
  MUX U5749 ( .IN0(n5661), .IN1(n5660), .SEL(N15), .F(n5662) );
  MUX U5750 ( .IN0(\registers[2][22] ), .IN1(\registers[3][22] ), .SEL(N14), 
        .F(n5663) );
  MUX U5752 ( .IN0(n5664), .IN1(n5663), .SEL(N15), .F(n5665) );
  MUX U5753 ( .IN0(n5665), .IN1(n5662), .SEL(N16), .F(n5666) );
  MUX U5754 ( .IN0(n5666), .IN1(n5659), .SEL(N17), .F(n5667) );
  MUX U5755 ( .IN0(n5667), .IN1(n5652), .SEL(N18), .F(reg_target_out[22]) );
  MUX U5756 ( .IN0(\registers[30][23] ), .IN1(\registers[31][23] ), .SEL(N14), 
        .F(n5668) );
  MUX U5757 ( .IN0(\registers[28][23] ), .IN1(\registers[29][23] ), .SEL(N14), 
        .F(n5669) );
  MUX U5758 ( .IN0(n5669), .IN1(n5668), .SEL(N15), .F(n5670) );
  MUX U5759 ( .IN0(\registers[26][23] ), .IN1(\registers[27][23] ), .SEL(N14), 
        .F(n5671) );
  MUX U5760 ( .IN0(\registers[24][23] ), .IN1(\registers[25][23] ), .SEL(N14), 
        .F(n5672) );
  MUX U5761 ( .IN0(n5672), .IN1(n5671), .SEL(N15), .F(n5673) );
  MUX U5762 ( .IN0(n5673), .IN1(n5670), .SEL(N16), .F(n5674) );
  MUX U5763 ( .IN0(\registers[22][23] ), .IN1(\registers[23][23] ), .SEL(N14), 
        .F(n5675) );
  MUX U5764 ( .IN0(\registers[20][23] ), .IN1(\registers[21][23] ), .SEL(N14), 
        .F(n5676) );
  MUX U5765 ( .IN0(n5676), .IN1(n5675), .SEL(N15), .F(n5677) );
  MUX U5766 ( .IN0(\registers[18][23] ), .IN1(\registers[19][23] ), .SEL(N14), 
        .F(n5678) );
  MUX U5767 ( .IN0(\registers[16][23] ), .IN1(\registers[17][23] ), .SEL(N14), 
        .F(n5679) );
  MUX U5768 ( .IN0(n5679), .IN1(n5678), .SEL(N15), .F(n5680) );
  MUX U5769 ( .IN0(n5680), .IN1(n5677), .SEL(N16), .F(n5681) );
  MUX U5770 ( .IN0(n5681), .IN1(n5674), .SEL(N17), .F(n5682) );
  MUX U5771 ( .IN0(\registers[14][23] ), .IN1(\registers[15][23] ), .SEL(N14), 
        .F(n5683) );
  MUX U5772 ( .IN0(\registers[12][23] ), .IN1(\registers[13][23] ), .SEL(N14), 
        .F(n5684) );
  MUX U5773 ( .IN0(n5684), .IN1(n5683), .SEL(N15), .F(n5685) );
  MUX U5774 ( .IN0(\registers[10][23] ), .IN1(\registers[11][23] ), .SEL(N14), 
        .F(n5686) );
  MUX U5775 ( .IN0(\registers[8][23] ), .IN1(\registers[9][23] ), .SEL(N14), 
        .F(n5687) );
  MUX U5776 ( .IN0(n5687), .IN1(n5686), .SEL(N15), .F(n5688) );
  MUX U5777 ( .IN0(n5688), .IN1(n5685), .SEL(N16), .F(n5689) );
  MUX U5778 ( .IN0(\registers[6][23] ), .IN1(\registers[7][23] ), .SEL(N14), 
        .F(n5690) );
  MUX U5779 ( .IN0(\registers[4][23] ), .IN1(\registers[5][23] ), .SEL(N14), 
        .F(n5691) );
  MUX U5780 ( .IN0(n5691), .IN1(n5690), .SEL(N15), .F(n5692) );
  MUX U5781 ( .IN0(\registers[2][23] ), .IN1(\registers[3][23] ), .SEL(N14), 
        .F(n5693) );
  MUX U5783 ( .IN0(n5694), .IN1(n5693), .SEL(N15), .F(n5695) );
  MUX U5784 ( .IN0(n5695), .IN1(n5692), .SEL(N16), .F(n5696) );
  MUX U5785 ( .IN0(n5696), .IN1(n5689), .SEL(N17), .F(n5697) );
  MUX U5786 ( .IN0(n5697), .IN1(n5682), .SEL(N18), .F(reg_target_out[23]) );
  MUX U5787 ( .IN0(\registers[30][24] ), .IN1(\registers[31][24] ), .SEL(N14), 
        .F(n5698) );
  MUX U5788 ( .IN0(\registers[28][24] ), .IN1(\registers[29][24] ), .SEL(N14), 
        .F(n5699) );
  MUX U5789 ( .IN0(n5699), .IN1(n5698), .SEL(N15), .F(n5700) );
  MUX U5790 ( .IN0(\registers[26][24] ), .IN1(\registers[27][24] ), .SEL(N14), 
        .F(n5701) );
  MUX U5791 ( .IN0(\registers[24][24] ), .IN1(\registers[25][24] ), .SEL(N14), 
        .F(n5702) );
  MUX U5792 ( .IN0(n5702), .IN1(n5701), .SEL(N15), .F(n5703) );
  MUX U5793 ( .IN0(n5703), .IN1(n5700), .SEL(N16), .F(n5704) );
  MUX U5794 ( .IN0(\registers[22][24] ), .IN1(\registers[23][24] ), .SEL(N14), 
        .F(n5705) );
  MUX U5795 ( .IN0(\registers[20][24] ), .IN1(\registers[21][24] ), .SEL(N14), 
        .F(n5706) );
  MUX U5796 ( .IN0(n5706), .IN1(n5705), .SEL(N15), .F(n5707) );
  MUX U5797 ( .IN0(\registers[18][24] ), .IN1(\registers[19][24] ), .SEL(N14), 
        .F(n5708) );
  MUX U5798 ( .IN0(\registers[16][24] ), .IN1(\registers[17][24] ), .SEL(N14), 
        .F(n5709) );
  MUX U5799 ( .IN0(n5709), .IN1(n5708), .SEL(N15), .F(n5710) );
  MUX U5800 ( .IN0(n5710), .IN1(n5707), .SEL(N16), .F(n5711) );
  MUX U5801 ( .IN0(n5711), .IN1(n5704), .SEL(N17), .F(n5712) );
  MUX U5802 ( .IN0(\registers[14][24] ), .IN1(\registers[15][24] ), .SEL(N14), 
        .F(n5713) );
  MUX U5803 ( .IN0(\registers[12][24] ), .IN1(\registers[13][24] ), .SEL(N14), 
        .F(n5714) );
  MUX U5804 ( .IN0(n5714), .IN1(n5713), .SEL(N15), .F(n5715) );
  MUX U5805 ( .IN0(\registers[10][24] ), .IN1(\registers[11][24] ), .SEL(N14), 
        .F(n5716) );
  MUX U5806 ( .IN0(\registers[8][24] ), .IN1(\registers[9][24] ), .SEL(N14), 
        .F(n5717) );
  MUX U5807 ( .IN0(n5717), .IN1(n5716), .SEL(N15), .F(n5718) );
  MUX U5808 ( .IN0(n5718), .IN1(n5715), .SEL(N16), .F(n5719) );
  MUX U5809 ( .IN0(\registers[6][24] ), .IN1(\registers[7][24] ), .SEL(N14), 
        .F(n5720) );
  MUX U5810 ( .IN0(\registers[4][24] ), .IN1(\registers[5][24] ), .SEL(N14), 
        .F(n5721) );
  MUX U5811 ( .IN0(n5721), .IN1(n5720), .SEL(N15), .F(n5722) );
  MUX U5812 ( .IN0(\registers[2][24] ), .IN1(\registers[3][24] ), .SEL(N14), 
        .F(n5723) );
  MUX U5814 ( .IN0(n5724), .IN1(n5723), .SEL(N15), .F(n5725) );
  MUX U5815 ( .IN0(n5725), .IN1(n5722), .SEL(N16), .F(n5726) );
  MUX U5816 ( .IN0(n5726), .IN1(n5719), .SEL(N17), .F(n5727) );
  MUX U5817 ( .IN0(n5727), .IN1(n5712), .SEL(N18), .F(reg_target_out[24]) );
  MUX U5818 ( .IN0(\registers[30][25] ), .IN1(\registers[31][25] ), .SEL(N14), 
        .F(n5728) );
  MUX U5819 ( .IN0(\registers[28][25] ), .IN1(\registers[29][25] ), .SEL(N14), 
        .F(n5729) );
  MUX U5820 ( .IN0(n5729), .IN1(n5728), .SEL(N15), .F(n5730) );
  MUX U5821 ( .IN0(\registers[26][25] ), .IN1(\registers[27][25] ), .SEL(N14), 
        .F(n5731) );
  MUX U5822 ( .IN0(\registers[24][25] ), .IN1(\registers[25][25] ), .SEL(N14), 
        .F(n5732) );
  MUX U5823 ( .IN0(n5732), .IN1(n5731), .SEL(N15), .F(n5733) );
  MUX U5824 ( .IN0(n5733), .IN1(n5730), .SEL(N16), .F(n5734) );
  MUX U5825 ( .IN0(\registers[22][25] ), .IN1(\registers[23][25] ), .SEL(N14), 
        .F(n5735) );
  MUX U5826 ( .IN0(\registers[20][25] ), .IN1(\registers[21][25] ), .SEL(N14), 
        .F(n5736) );
  MUX U5827 ( .IN0(n5736), .IN1(n5735), .SEL(N15), .F(n5737) );
  MUX U5828 ( .IN0(\registers[18][25] ), .IN1(\registers[19][25] ), .SEL(N14), 
        .F(n5738) );
  MUX U5829 ( .IN0(\registers[16][25] ), .IN1(\registers[17][25] ), .SEL(N14), 
        .F(n5739) );
  MUX U5830 ( .IN0(n5739), .IN1(n5738), .SEL(N15), .F(n5740) );
  MUX U5831 ( .IN0(n5740), .IN1(n5737), .SEL(N16), .F(n5741) );
  MUX U5832 ( .IN0(n5741), .IN1(n5734), .SEL(N17), .F(n5742) );
  MUX U5833 ( .IN0(\registers[14][25] ), .IN1(\registers[15][25] ), .SEL(N14), 
        .F(n5743) );
  MUX U5834 ( .IN0(\registers[12][25] ), .IN1(\registers[13][25] ), .SEL(N14), 
        .F(n5744) );
  MUX U5835 ( .IN0(n5744), .IN1(n5743), .SEL(N15), .F(n5745) );
  MUX U5836 ( .IN0(\registers[10][25] ), .IN1(\registers[11][25] ), .SEL(N14), 
        .F(n5746) );
  MUX U5837 ( .IN0(\registers[8][25] ), .IN1(\registers[9][25] ), .SEL(N14), 
        .F(n5747) );
  MUX U5838 ( .IN0(n5747), .IN1(n5746), .SEL(N15), .F(n5748) );
  MUX U5839 ( .IN0(n5748), .IN1(n5745), .SEL(N16), .F(n5749) );
  MUX U5840 ( .IN0(\registers[6][25] ), .IN1(\registers[7][25] ), .SEL(N14), 
        .F(n5750) );
  MUX U5841 ( .IN0(\registers[4][25] ), .IN1(\registers[5][25] ), .SEL(N14), 
        .F(n5751) );
  MUX U5842 ( .IN0(n5751), .IN1(n5750), .SEL(N15), .F(n5752) );
  MUX U5843 ( .IN0(\registers[2][25] ), .IN1(\registers[3][25] ), .SEL(N14), 
        .F(n5753) );
  MUX U5845 ( .IN0(n5754), .IN1(n5753), .SEL(N15), .F(n5755) );
  MUX U5846 ( .IN0(n5755), .IN1(n5752), .SEL(N16), .F(n5756) );
  MUX U5847 ( .IN0(n5756), .IN1(n5749), .SEL(N17), .F(n5757) );
  MUX U5848 ( .IN0(n5757), .IN1(n5742), .SEL(N18), .F(reg_target_out[25]) );
  MUX U5849 ( .IN0(\registers[30][26] ), .IN1(\registers[31][26] ), .SEL(N14), 
        .F(n5758) );
  MUX U5850 ( .IN0(\registers[28][26] ), .IN1(\registers[29][26] ), .SEL(N14), 
        .F(n5759) );
  MUX U5851 ( .IN0(n5759), .IN1(n5758), .SEL(N15), .F(n5760) );
  MUX U5852 ( .IN0(\registers[26][26] ), .IN1(\registers[27][26] ), .SEL(N14), 
        .F(n5761) );
  MUX U5853 ( .IN0(\registers[24][26] ), .IN1(\registers[25][26] ), .SEL(N14), 
        .F(n5762) );
  MUX U5854 ( .IN0(n5762), .IN1(n5761), .SEL(N15), .F(n5763) );
  MUX U5855 ( .IN0(n5763), .IN1(n5760), .SEL(N16), .F(n5764) );
  MUX U5856 ( .IN0(\registers[22][26] ), .IN1(\registers[23][26] ), .SEL(N14), 
        .F(n5765) );
  MUX U5857 ( .IN0(\registers[20][26] ), .IN1(\registers[21][26] ), .SEL(N14), 
        .F(n5766) );
  MUX U5858 ( .IN0(n5766), .IN1(n5765), .SEL(N15), .F(n5767) );
  MUX U5859 ( .IN0(\registers[18][26] ), .IN1(\registers[19][26] ), .SEL(N14), 
        .F(n5768) );
  MUX U5860 ( .IN0(\registers[16][26] ), .IN1(\registers[17][26] ), .SEL(N14), 
        .F(n5769) );
  MUX U5861 ( .IN0(n5769), .IN1(n5768), .SEL(N15), .F(n5770) );
  MUX U5862 ( .IN0(n5770), .IN1(n5767), .SEL(N16), .F(n5771) );
  MUX U5863 ( .IN0(n5771), .IN1(n5764), .SEL(N17), .F(n5772) );
  MUX U5864 ( .IN0(\registers[14][26] ), .IN1(\registers[15][26] ), .SEL(N14), 
        .F(n5773) );
  MUX U5865 ( .IN0(\registers[12][26] ), .IN1(\registers[13][26] ), .SEL(N14), 
        .F(n5774) );
  MUX U5866 ( .IN0(n5774), .IN1(n5773), .SEL(N15), .F(n5775) );
  MUX U5867 ( .IN0(\registers[10][26] ), .IN1(\registers[11][26] ), .SEL(N14), 
        .F(n5776) );
  MUX U5868 ( .IN0(\registers[8][26] ), .IN1(\registers[9][26] ), .SEL(N14), 
        .F(n5777) );
  MUX U5869 ( .IN0(n5777), .IN1(n5776), .SEL(N15), .F(n5778) );
  MUX U5870 ( .IN0(n5778), .IN1(n5775), .SEL(N16), .F(n5779) );
  MUX U5871 ( .IN0(\registers[6][26] ), .IN1(\registers[7][26] ), .SEL(N14), 
        .F(n5780) );
  MUX U5872 ( .IN0(\registers[4][26] ), .IN1(\registers[5][26] ), .SEL(N14), 
        .F(n5781) );
  MUX U5873 ( .IN0(n5781), .IN1(n5780), .SEL(N15), .F(n5782) );
  MUX U5874 ( .IN0(\registers[2][26] ), .IN1(\registers[3][26] ), .SEL(N14), 
        .F(n5783) );
  MUX U5876 ( .IN0(n5784), .IN1(n5783), .SEL(N15), .F(n5785) );
  MUX U5877 ( .IN0(n5785), .IN1(n5782), .SEL(N16), .F(n5786) );
  MUX U5878 ( .IN0(n5786), .IN1(n5779), .SEL(N17), .F(n5787) );
  MUX U5879 ( .IN0(n5787), .IN1(n5772), .SEL(N18), .F(reg_target_out[26]) );
  MUX U5880 ( .IN0(\registers[30][27] ), .IN1(\registers[31][27] ), .SEL(N14), 
        .F(n5788) );
  MUX U5881 ( .IN0(\registers[28][27] ), .IN1(\registers[29][27] ), .SEL(N14), 
        .F(n5789) );
  MUX U5882 ( .IN0(n5789), .IN1(n5788), .SEL(N15), .F(n5790) );
  MUX U5883 ( .IN0(\registers[26][27] ), .IN1(\registers[27][27] ), .SEL(N14), 
        .F(n5791) );
  MUX U5884 ( .IN0(\registers[24][27] ), .IN1(\registers[25][27] ), .SEL(N14), 
        .F(n5792) );
  MUX U5885 ( .IN0(n5792), .IN1(n5791), .SEL(N15), .F(n5793) );
  MUX U5886 ( .IN0(n5793), .IN1(n5790), .SEL(N16), .F(n5794) );
  MUX U5887 ( .IN0(\registers[22][27] ), .IN1(\registers[23][27] ), .SEL(N14), 
        .F(n5795) );
  MUX U5888 ( .IN0(\registers[20][27] ), .IN1(\registers[21][27] ), .SEL(N14), 
        .F(n5796) );
  MUX U5889 ( .IN0(n5796), .IN1(n5795), .SEL(N15), .F(n5797) );
  MUX U5890 ( .IN0(\registers[18][27] ), .IN1(\registers[19][27] ), .SEL(N14), 
        .F(n5798) );
  MUX U5891 ( .IN0(\registers[16][27] ), .IN1(\registers[17][27] ), .SEL(N14), 
        .F(n5799) );
  MUX U5892 ( .IN0(n5799), .IN1(n5798), .SEL(N15), .F(n5800) );
  MUX U5893 ( .IN0(n5800), .IN1(n5797), .SEL(N16), .F(n5801) );
  MUX U5894 ( .IN0(n5801), .IN1(n5794), .SEL(N17), .F(n5802) );
  MUX U5895 ( .IN0(\registers[14][27] ), .IN1(\registers[15][27] ), .SEL(N14), 
        .F(n5803) );
  MUX U5896 ( .IN0(\registers[12][27] ), .IN1(\registers[13][27] ), .SEL(N14), 
        .F(n5804) );
  MUX U5897 ( .IN0(n5804), .IN1(n5803), .SEL(N15), .F(n5805) );
  MUX U5898 ( .IN0(\registers[10][27] ), .IN1(\registers[11][27] ), .SEL(N14), 
        .F(n5806) );
  MUX U5899 ( .IN0(\registers[8][27] ), .IN1(\registers[9][27] ), .SEL(N14), 
        .F(n5807) );
  MUX U5900 ( .IN0(n5807), .IN1(n5806), .SEL(N15), .F(n5808) );
  MUX U5901 ( .IN0(n5808), .IN1(n5805), .SEL(N16), .F(n5809) );
  MUX U5902 ( .IN0(\registers[6][27] ), .IN1(\registers[7][27] ), .SEL(N14), 
        .F(n5810) );
  MUX U5903 ( .IN0(\registers[4][27] ), .IN1(\registers[5][27] ), .SEL(N14), 
        .F(n5811) );
  MUX U5904 ( .IN0(n5811), .IN1(n5810), .SEL(N15), .F(n5812) );
  MUX U5905 ( .IN0(\registers[2][27] ), .IN1(\registers[3][27] ), .SEL(N14), 
        .F(n5813) );
  MUX U5907 ( .IN0(n5814), .IN1(n5813), .SEL(N15), .F(n5815) );
  MUX U5908 ( .IN0(n5815), .IN1(n5812), .SEL(N16), .F(n5816) );
  MUX U5909 ( .IN0(n5816), .IN1(n5809), .SEL(N17), .F(n5817) );
  MUX U5910 ( .IN0(n5817), .IN1(n5802), .SEL(N18), .F(reg_target_out[27]) );
  MUX U5911 ( .IN0(\registers[30][28] ), .IN1(\registers[31][28] ), .SEL(N14), 
        .F(n5818) );
  MUX U5912 ( .IN0(\registers[28][28] ), .IN1(\registers[29][28] ), .SEL(N14), 
        .F(n5819) );
  MUX U5913 ( .IN0(n5819), .IN1(n5818), .SEL(N15), .F(n5820) );
  MUX U5914 ( .IN0(\registers[26][28] ), .IN1(\registers[27][28] ), .SEL(N14), 
        .F(n5821) );
  MUX U5915 ( .IN0(\registers[24][28] ), .IN1(\registers[25][28] ), .SEL(N14), 
        .F(n5822) );
  MUX U5916 ( .IN0(n5822), .IN1(n5821), .SEL(N15), .F(n5823) );
  MUX U5917 ( .IN0(n5823), .IN1(n5820), .SEL(N16), .F(n5824) );
  MUX U5918 ( .IN0(\registers[22][28] ), .IN1(\registers[23][28] ), .SEL(N14), 
        .F(n5825) );
  MUX U5919 ( .IN0(\registers[20][28] ), .IN1(\registers[21][28] ), .SEL(N14), 
        .F(n5826) );
  MUX U5920 ( .IN0(n5826), .IN1(n5825), .SEL(N15), .F(n5827) );
  MUX U5921 ( .IN0(\registers[18][28] ), .IN1(\registers[19][28] ), .SEL(N14), 
        .F(n5828) );
  MUX U5922 ( .IN0(\registers[16][28] ), .IN1(\registers[17][28] ), .SEL(N14), 
        .F(n5829) );
  MUX U5923 ( .IN0(n5829), .IN1(n5828), .SEL(N15), .F(n5830) );
  MUX U5924 ( .IN0(n5830), .IN1(n5827), .SEL(N16), .F(n5831) );
  MUX U5925 ( .IN0(n5831), .IN1(n5824), .SEL(N17), .F(n5832) );
  MUX U5926 ( .IN0(\registers[14][28] ), .IN1(\registers[15][28] ), .SEL(N14), 
        .F(n5833) );
  MUX U5927 ( .IN0(\registers[12][28] ), .IN1(\registers[13][28] ), .SEL(N14), 
        .F(n5834) );
  MUX U5928 ( .IN0(n5834), .IN1(n5833), .SEL(N15), .F(n5835) );
  MUX U5929 ( .IN0(\registers[10][28] ), .IN1(\registers[11][28] ), .SEL(N14), 
        .F(n5836) );
  MUX U5930 ( .IN0(\registers[8][28] ), .IN1(\registers[9][28] ), .SEL(N14), 
        .F(n5837) );
  MUX U5931 ( .IN0(n5837), .IN1(n5836), .SEL(N15), .F(n5838) );
  MUX U5932 ( .IN0(n5838), .IN1(n5835), .SEL(N16), .F(n5839) );
  MUX U5933 ( .IN0(\registers[6][28] ), .IN1(\registers[7][28] ), .SEL(N14), 
        .F(n5840) );
  MUX U5934 ( .IN0(\registers[4][28] ), .IN1(\registers[5][28] ), .SEL(N14), 
        .F(n5841) );
  MUX U5935 ( .IN0(n5841), .IN1(n5840), .SEL(N15), .F(n5842) );
  MUX U5936 ( .IN0(\registers[2][28] ), .IN1(\registers[3][28] ), .SEL(N14), 
        .F(n5843) );
  MUX U5938 ( .IN0(n5844), .IN1(n5843), .SEL(N15), .F(n5845) );
  MUX U5939 ( .IN0(n5845), .IN1(n5842), .SEL(N16), .F(n5846) );
  MUX U5940 ( .IN0(n5846), .IN1(n5839), .SEL(N17), .F(n5847) );
  MUX U5941 ( .IN0(n5847), .IN1(n5832), .SEL(N18), .F(reg_target_out[28]) );
  MUX U5942 ( .IN0(\registers[30][29] ), .IN1(\registers[31][29] ), .SEL(N14), 
        .F(n5848) );
  MUX U5943 ( .IN0(\registers[28][29] ), .IN1(\registers[29][29] ), .SEL(N14), 
        .F(n5849) );
  MUX U5944 ( .IN0(n5849), .IN1(n5848), .SEL(N15), .F(n5850) );
  MUX U5945 ( .IN0(\registers[26][29] ), .IN1(\registers[27][29] ), .SEL(N14), 
        .F(n5851) );
  MUX U5946 ( .IN0(\registers[24][29] ), .IN1(\registers[25][29] ), .SEL(N14), 
        .F(n5852) );
  MUX U5947 ( .IN0(n5852), .IN1(n5851), .SEL(N15), .F(n5853) );
  MUX U5948 ( .IN0(n5853), .IN1(n5850), .SEL(N16), .F(n5854) );
  MUX U5949 ( .IN0(\registers[22][29] ), .IN1(\registers[23][29] ), .SEL(N14), 
        .F(n5855) );
  MUX U5950 ( .IN0(\registers[20][29] ), .IN1(\registers[21][29] ), .SEL(N14), 
        .F(n5856) );
  MUX U5951 ( .IN0(n5856), .IN1(n5855), .SEL(N15), .F(n5857) );
  MUX U5952 ( .IN0(\registers[18][29] ), .IN1(\registers[19][29] ), .SEL(N14), 
        .F(n5858) );
  MUX U5953 ( .IN0(\registers[16][29] ), .IN1(\registers[17][29] ), .SEL(N14), 
        .F(n5859) );
  MUX U5954 ( .IN0(n5859), .IN1(n5858), .SEL(N15), .F(n5860) );
  MUX U5955 ( .IN0(n5860), .IN1(n5857), .SEL(N16), .F(n5861) );
  MUX U5956 ( .IN0(n5861), .IN1(n5854), .SEL(N17), .F(n5862) );
  MUX U5957 ( .IN0(\registers[14][29] ), .IN1(\registers[15][29] ), .SEL(N14), 
        .F(n5863) );
  MUX U5958 ( .IN0(\registers[12][29] ), .IN1(\registers[13][29] ), .SEL(N14), 
        .F(n5864) );
  MUX U5959 ( .IN0(n5864), .IN1(n5863), .SEL(N15), .F(n5865) );
  MUX U5960 ( .IN0(\registers[10][29] ), .IN1(\registers[11][29] ), .SEL(N14), 
        .F(n5866) );
  MUX U5961 ( .IN0(\registers[8][29] ), .IN1(\registers[9][29] ), .SEL(N14), 
        .F(n5867) );
  MUX U5962 ( .IN0(n5867), .IN1(n5866), .SEL(N15), .F(n5868) );
  MUX U5963 ( .IN0(n5868), .IN1(n5865), .SEL(N16), .F(n5869) );
  MUX U5964 ( .IN0(\registers[6][29] ), .IN1(\registers[7][29] ), .SEL(N14), 
        .F(n5870) );
  MUX U5965 ( .IN0(\registers[4][29] ), .IN1(\registers[5][29] ), .SEL(N14), 
        .F(n5871) );
  MUX U5966 ( .IN0(n5871), .IN1(n5870), .SEL(N15), .F(n5872) );
  MUX U5967 ( .IN0(\registers[2][29] ), .IN1(\registers[3][29] ), .SEL(N14), 
        .F(n5873) );
  MUX U5969 ( .IN0(n5874), .IN1(n5873), .SEL(N15), .F(n5875) );
  MUX U5970 ( .IN0(n5875), .IN1(n5872), .SEL(N16), .F(n5876) );
  MUX U5971 ( .IN0(n5876), .IN1(n5869), .SEL(N17), .F(n5877) );
  MUX U5972 ( .IN0(n5877), .IN1(n5862), .SEL(N18), .F(reg_target_out[29]) );
  MUX U5973 ( .IN0(\registers[30][30] ), .IN1(\registers[31][30] ), .SEL(N14), 
        .F(n5878) );
  MUX U5974 ( .IN0(\registers[28][30] ), .IN1(\registers[29][30] ), .SEL(N14), 
        .F(n5879) );
  MUX U5975 ( .IN0(n5879), .IN1(n5878), .SEL(N15), .F(n5880) );
  MUX U5976 ( .IN0(\registers[26][30] ), .IN1(\registers[27][30] ), .SEL(N14), 
        .F(n5881) );
  MUX U5977 ( .IN0(\registers[24][30] ), .IN1(\registers[25][30] ), .SEL(N14), 
        .F(n5882) );
  MUX U5978 ( .IN0(n5882), .IN1(n5881), .SEL(N15), .F(n5883) );
  MUX U5979 ( .IN0(n5883), .IN1(n5880), .SEL(N16), .F(n5884) );
  MUX U5980 ( .IN0(\registers[22][30] ), .IN1(\registers[23][30] ), .SEL(N14), 
        .F(n5885) );
  MUX U5981 ( .IN0(\registers[20][30] ), .IN1(\registers[21][30] ), .SEL(N14), 
        .F(n5886) );
  MUX U5982 ( .IN0(n5886), .IN1(n5885), .SEL(N15), .F(n5887) );
  MUX U5983 ( .IN0(\registers[18][30] ), .IN1(\registers[19][30] ), .SEL(N14), 
        .F(n5888) );
  MUX U5984 ( .IN0(\registers[16][30] ), .IN1(\registers[17][30] ), .SEL(N14), 
        .F(n5889) );
  MUX U5985 ( .IN0(n5889), .IN1(n5888), .SEL(N15), .F(n5890) );
  MUX U5986 ( .IN0(n5890), .IN1(n5887), .SEL(N16), .F(n5891) );
  MUX U5987 ( .IN0(n5891), .IN1(n5884), .SEL(N17), .F(n5892) );
  MUX U5988 ( .IN0(\registers[14][30] ), .IN1(\registers[15][30] ), .SEL(N14), 
        .F(n5893) );
  MUX U5989 ( .IN0(\registers[12][30] ), .IN1(\registers[13][30] ), .SEL(N14), 
        .F(n5894) );
  MUX U5990 ( .IN0(n5894), .IN1(n5893), .SEL(N15), .F(n5895) );
  MUX U5991 ( .IN0(\registers[10][30] ), .IN1(\registers[11][30] ), .SEL(N14), 
        .F(n5896) );
  MUX U5992 ( .IN0(\registers[8][30] ), .IN1(\registers[9][30] ), .SEL(N14), 
        .F(n5897) );
  MUX U5993 ( .IN0(n5897), .IN1(n5896), .SEL(N15), .F(n5898) );
  MUX U5994 ( .IN0(n5898), .IN1(n5895), .SEL(N16), .F(n5899) );
  MUX U5995 ( .IN0(\registers[6][30] ), .IN1(\registers[7][30] ), .SEL(N14), 
        .F(n5900) );
  MUX U5996 ( .IN0(\registers[4][30] ), .IN1(\registers[5][30] ), .SEL(N14), 
        .F(n5901) );
  MUX U5997 ( .IN0(n5901), .IN1(n5900), .SEL(N15), .F(n5902) );
  MUX U5998 ( .IN0(\registers[2][30] ), .IN1(\registers[3][30] ), .SEL(N14), 
        .F(n5903) );
  MUX U6000 ( .IN0(n5904), .IN1(n5903), .SEL(N15), .F(n5905) );
  MUX U6001 ( .IN0(n5905), .IN1(n5902), .SEL(N16), .F(n5906) );
  MUX U6002 ( .IN0(n5906), .IN1(n5899), .SEL(N17), .F(n5907) );
  MUX U6003 ( .IN0(n5907), .IN1(n5892), .SEL(N18), .F(reg_target_out[30]) );
  MUX U6004 ( .IN0(\registers[30][31] ), .IN1(\registers[31][31] ), .SEL(N14), 
        .F(n5908) );
  MUX U6005 ( .IN0(\registers[28][31] ), .IN1(\registers[29][31] ), .SEL(N14), 
        .F(n5909) );
  MUX U6006 ( .IN0(n5909), .IN1(n5908), .SEL(N15), .F(n5910) );
  MUX U6007 ( .IN0(\registers[26][31] ), .IN1(\registers[27][31] ), .SEL(N14), 
        .F(n5911) );
  MUX U6008 ( .IN0(\registers[24][31] ), .IN1(\registers[25][31] ), .SEL(N14), 
        .F(n5912) );
  MUX U6009 ( .IN0(n5912), .IN1(n5911), .SEL(N15), .F(n5913) );
  MUX U6010 ( .IN0(n5913), .IN1(n5910), .SEL(N16), .F(n5914) );
  MUX U6011 ( .IN0(\registers[22][31] ), .IN1(\registers[23][31] ), .SEL(N14), 
        .F(n5915) );
  MUX U6012 ( .IN0(\registers[20][31] ), .IN1(\registers[21][31] ), .SEL(N14), 
        .F(n5916) );
  MUX U6013 ( .IN0(n5916), .IN1(n5915), .SEL(N15), .F(n5917) );
  MUX U6014 ( .IN0(\registers[18][31] ), .IN1(\registers[19][31] ), .SEL(N14), 
        .F(n5918) );
  MUX U6015 ( .IN0(\registers[16][31] ), .IN1(\registers[17][31] ), .SEL(N14), 
        .F(n5919) );
  MUX U6016 ( .IN0(n5919), .IN1(n5918), .SEL(N15), .F(n5920) );
  MUX U6017 ( .IN0(n5920), .IN1(n5917), .SEL(N16), .F(n5921) );
  MUX U6018 ( .IN0(n5921), .IN1(n5914), .SEL(N17), .F(n5922) );
  MUX U6019 ( .IN0(\registers[14][31] ), .IN1(\registers[15][31] ), .SEL(N14), 
        .F(n5923) );
  MUX U6020 ( .IN0(\registers[12][31] ), .IN1(\registers[13][31] ), .SEL(N14), 
        .F(n5924) );
  MUX U6021 ( .IN0(n5924), .IN1(n5923), .SEL(N15), .F(n5925) );
  MUX U6022 ( .IN0(\registers[10][31] ), .IN1(\registers[11][31] ), .SEL(N14), 
        .F(n5926) );
  MUX U6023 ( .IN0(\registers[8][31] ), .IN1(\registers[9][31] ), .SEL(N14), 
        .F(n5927) );
  MUX U6024 ( .IN0(n5927), .IN1(n5926), .SEL(N15), .F(n5928) );
  MUX U6025 ( .IN0(n5928), .IN1(n5925), .SEL(N16), .F(n5929) );
  MUX U6026 ( .IN0(\registers[6][31] ), .IN1(\registers[7][31] ), .SEL(N14), 
        .F(n5930) );
  MUX U6027 ( .IN0(\registers[4][31] ), .IN1(\registers[5][31] ), .SEL(N14), 
        .F(n5931) );
  MUX U6028 ( .IN0(n5931), .IN1(n5930), .SEL(N15), .F(n5932) );
  MUX U6029 ( .IN0(\registers[2][31] ), .IN1(\registers[3][31] ), .SEL(N14), 
        .F(n5933) );
  MUX U6031 ( .IN0(n5934), .IN1(n5933), .SEL(N15), .F(n5935) );
  MUX U6032 ( .IN0(n5935), .IN1(n5932), .SEL(N16), .F(n5936) );
  MUX U6033 ( .IN0(n5936), .IN1(n5929), .SEL(N17), .F(n5937) );
  MUX U6034 ( .IN0(n5937), .IN1(n5922), .SEL(N18), .F(reg_target_out[31]) );
  AND U6035 ( .A(N14), .B(\registers[1][0] ), .Z(n5004) );
  AND U6036 ( .A(N9), .B(\registers[1][0] ), .Z(n4044) );
  AND U6037 ( .A(N14), .B(\registers[1][1] ), .Z(n5034) );
  AND U6038 ( .A(N9), .B(\registers[1][1] ), .Z(n4074) );
  AND U6039 ( .A(N14), .B(\registers[1][2] ), .Z(n5064) );
  AND U6040 ( .A(N9), .B(\registers[1][2] ), .Z(n4104) );
  AND U6041 ( .A(N14), .B(\registers[1][3] ), .Z(n5094) );
  AND U6042 ( .A(N9), .B(\registers[1][3] ), .Z(n4134) );
  AND U6043 ( .A(N14), .B(\registers[1][4] ), .Z(n5124) );
  AND U6044 ( .A(N9), .B(\registers[1][4] ), .Z(n4164) );
  AND U6045 ( .A(N14), .B(\registers[1][5] ), .Z(n5154) );
  AND U6046 ( .A(N9), .B(\registers[1][5] ), .Z(n4194) );
  AND U6047 ( .A(N14), .B(\registers[1][6] ), .Z(n5184) );
  AND U6048 ( .A(N9), .B(\registers[1][6] ), .Z(n4224) );
  AND U6049 ( .A(N14), .B(\registers[1][7] ), .Z(n5214) );
  AND U6050 ( .A(N9), .B(\registers[1][7] ), .Z(n4254) );
  AND U6051 ( .A(N14), .B(\registers[1][8] ), .Z(n5244) );
  AND U6052 ( .A(N9), .B(\registers[1][8] ), .Z(n4284) );
  AND U6053 ( .A(N14), .B(\registers[1][9] ), .Z(n5274) );
  AND U6054 ( .A(N9), .B(\registers[1][9] ), .Z(n4314) );
  AND U6055 ( .A(N14), .B(\registers[1][10] ), .Z(n5304) );
  AND U6056 ( .A(N9), .B(\registers[1][10] ), .Z(n4344) );
  AND U6057 ( .A(N14), .B(\registers[1][11] ), .Z(n5334) );
  AND U6058 ( .A(N9), .B(\registers[1][11] ), .Z(n4374) );
  AND U6059 ( .A(N14), .B(\registers[1][12] ), .Z(n5364) );
  AND U6060 ( .A(N9), .B(\registers[1][12] ), .Z(n4404) );
  AND U6061 ( .A(N14), .B(\registers[1][13] ), .Z(n5394) );
  AND U6062 ( .A(N9), .B(\registers[1][13] ), .Z(n4434) );
  AND U6063 ( .A(N14), .B(\registers[1][14] ), .Z(n5424) );
  AND U6064 ( .A(N9), .B(\registers[1][14] ), .Z(n4464) );
  AND U6065 ( .A(N14), .B(\registers[1][15] ), .Z(n5454) );
  AND U6066 ( .A(N9), .B(\registers[1][15] ), .Z(n4494) );
  AND U6067 ( .A(N14), .B(\registers[1][16] ), .Z(n5484) );
  AND U6068 ( .A(N9), .B(\registers[1][16] ), .Z(n4524) );
  AND U6069 ( .A(N14), .B(\registers[1][17] ), .Z(n5514) );
  AND U6070 ( .A(N9), .B(\registers[1][17] ), .Z(n4554) );
  AND U6071 ( .A(N14), .B(\registers[1][18] ), .Z(n5544) );
  AND U6072 ( .A(N9), .B(\registers[1][18] ), .Z(n4584) );
  AND U6073 ( .A(N14), .B(\registers[1][19] ), .Z(n5574) );
  AND U6074 ( .A(N9), .B(\registers[1][19] ), .Z(n4614) );
  AND U6075 ( .A(N14), .B(\registers[1][20] ), .Z(n5604) );
  AND U6076 ( .A(N9), .B(\registers[1][20] ), .Z(n4644) );
  AND U6077 ( .A(N14), .B(\registers[1][21] ), .Z(n5634) );
  AND U6078 ( .A(N9), .B(\registers[1][21] ), .Z(n4674) );
  AND U6079 ( .A(N14), .B(\registers[1][22] ), .Z(n5664) );
  AND U6080 ( .A(N9), .B(\registers[1][22] ), .Z(n4704) );
  AND U6081 ( .A(N14), .B(\registers[1][23] ), .Z(n5694) );
  AND U6082 ( .A(N9), .B(\registers[1][23] ), .Z(n4734) );
  AND U6083 ( .A(N14), .B(\registers[1][24] ), .Z(n5724) );
  AND U6084 ( .A(N9), .B(\registers[1][24] ), .Z(n4764) );
  AND U6085 ( .A(N14), .B(\registers[1][25] ), .Z(n5754) );
  AND U6086 ( .A(N9), .B(\registers[1][25] ), .Z(n4794) );
  AND U6087 ( .A(N14), .B(\registers[1][26] ), .Z(n5784) );
  AND U6088 ( .A(N9), .B(\registers[1][26] ), .Z(n4824) );
  AND U6089 ( .A(N14), .B(\registers[1][27] ), .Z(n5814) );
  AND U6090 ( .A(N9), .B(\registers[1][27] ), .Z(n4854) );
  AND U6091 ( .A(N14), .B(\registers[1][28] ), .Z(n5844) );
  AND U6092 ( .A(N9), .B(\registers[1][28] ), .Z(n4884) );
  AND U6093 ( .A(N14), .B(\registers[1][29] ), .Z(n5874) );
  AND U6094 ( .A(N9), .B(\registers[1][29] ), .Z(n4914) );
  AND U6095 ( .A(N14), .B(\registers[1][30] ), .Z(n5904) );
  AND U6096 ( .A(N9), .B(\registers[1][30] ), .Z(n4944) );
  AND U6097 ( .A(N14), .B(\registers[1][31] ), .Z(n5934) );
  AND U6098 ( .A(N9), .B(\registers[1][31] ), .Z(n4974) );
  MUX U6099 ( .IN0(reg_dest_new[31]), .IN1(\registers[31][31] ), .SEL(n5938), 
        .F(n4017) );
  MUX U6100 ( .IN0(reg_dest_new[30]), .IN1(\registers[31][30] ), .SEL(n5938), 
        .F(n4016) );
  MUX U6101 ( .IN0(reg_dest_new[29]), .IN1(\registers[31][29] ), .SEL(n5938), 
        .F(n4015) );
  MUX U6102 ( .IN0(reg_dest_new[28]), .IN1(\registers[31][28] ), .SEL(n5938), 
        .F(n4014) );
  MUX U6103 ( .IN0(reg_dest_new[27]), .IN1(\registers[31][27] ), .SEL(n5938), 
        .F(n4013) );
  MUX U6104 ( .IN0(reg_dest_new[26]), .IN1(\registers[31][26] ), .SEL(n5938), 
        .F(n4012) );
  MUX U6105 ( .IN0(reg_dest_new[25]), .IN1(\registers[31][25] ), .SEL(n5938), 
        .F(n4011) );
  MUX U6106 ( .IN0(reg_dest_new[24]), .IN1(\registers[31][24] ), .SEL(n5938), 
        .F(n4010) );
  MUX U6107 ( .IN0(reg_dest_new[23]), .IN1(\registers[31][23] ), .SEL(n5938), 
        .F(n4009) );
  MUX U6108 ( .IN0(reg_dest_new[22]), .IN1(\registers[31][22] ), .SEL(n5938), 
        .F(n4008) );
  MUX U6109 ( .IN0(reg_dest_new[21]), .IN1(\registers[31][21] ), .SEL(n5938), 
        .F(n4007) );
  MUX U6110 ( .IN0(reg_dest_new[20]), .IN1(\registers[31][20] ), .SEL(n5938), 
        .F(n4006) );
  MUX U6111 ( .IN0(reg_dest_new[19]), .IN1(\registers[31][19] ), .SEL(n5938), 
        .F(n4005) );
  MUX U6112 ( .IN0(reg_dest_new[18]), .IN1(\registers[31][18] ), .SEL(n5938), 
        .F(n4004) );
  MUX U6113 ( .IN0(reg_dest_new[17]), .IN1(\registers[31][17] ), .SEL(n5938), 
        .F(n4003) );
  MUX U6114 ( .IN0(reg_dest_new[16]), .IN1(\registers[31][16] ), .SEL(n5938), 
        .F(n4002) );
  MUX U6115 ( .IN0(reg_dest_new[15]), .IN1(\registers[31][15] ), .SEL(n5938), 
        .F(n4001) );
  MUX U6116 ( .IN0(reg_dest_new[14]), .IN1(\registers[31][14] ), .SEL(n5938), 
        .F(n4000) );
  MUX U6117 ( .IN0(reg_dest_new[13]), .IN1(\registers[31][13] ), .SEL(n5938), 
        .F(n3999) );
  MUX U6118 ( .IN0(reg_dest_new[12]), .IN1(\registers[31][12] ), .SEL(n5938), 
        .F(n3998) );
  MUX U6119 ( .IN0(reg_dest_new[11]), .IN1(\registers[31][11] ), .SEL(n5938), 
        .F(n3997) );
  MUX U6120 ( .IN0(reg_dest_new[10]), .IN1(\registers[31][10] ), .SEL(n5938), 
        .F(n3996) );
  MUX U6121 ( .IN0(reg_dest_new[9]), .IN1(\registers[31][9] ), .SEL(n5938), 
        .F(n3995) );
  MUX U6122 ( .IN0(reg_dest_new[8]), .IN1(\registers[31][8] ), .SEL(n5938), 
        .F(n3994) );
  MUX U6123 ( .IN0(reg_dest_new[7]), .IN1(\registers[31][7] ), .SEL(n5938), 
        .F(n3993) );
  MUX U6124 ( .IN0(reg_dest_new[6]), .IN1(\registers[31][6] ), .SEL(n5938), 
        .F(n3992) );
  MUX U6125 ( .IN0(reg_dest_new[5]), .IN1(\registers[31][5] ), .SEL(n5938), 
        .F(n3991) );
  MUX U6126 ( .IN0(reg_dest_new[4]), .IN1(\registers[31][4] ), .SEL(n5938), 
        .F(n3990) );
  MUX U6127 ( .IN0(reg_dest_new[3]), .IN1(\registers[31][3] ), .SEL(n5938), 
        .F(n3989) );
  MUX U6128 ( .IN0(reg_dest_new[2]), .IN1(\registers[31][2] ), .SEL(n5938), 
        .F(n3988) );
  IV U6129 ( .A(n5939), .Z(n5938) );
  MUX U6130 ( .IN0(\registers[31][1] ), .IN1(reg_dest_new[1]), .SEL(n5939), 
        .F(n3987) );
  MUX U6131 ( .IN0(\registers[31][0] ), .IN1(reg_dest_new[0]), .SEL(n5939), 
        .F(n3986) );
  NOR U6132 ( .A(n5940), .B(n5941), .Z(n5939) );
  MUX U6133 ( .IN0(reg_dest_new[31]), .IN1(\registers[30][31] ), .SEL(n5942), 
        .F(n3985) );
  MUX U6134 ( .IN0(reg_dest_new[30]), .IN1(\registers[30][30] ), .SEL(n5942), 
        .F(n3984) );
  MUX U6135 ( .IN0(reg_dest_new[29]), .IN1(\registers[30][29] ), .SEL(n5942), 
        .F(n3983) );
  MUX U6136 ( .IN0(reg_dest_new[28]), .IN1(\registers[30][28] ), .SEL(n5942), 
        .F(n3982) );
  MUX U6137 ( .IN0(reg_dest_new[27]), .IN1(\registers[30][27] ), .SEL(n5942), 
        .F(n3981) );
  MUX U6138 ( .IN0(reg_dest_new[26]), .IN1(\registers[30][26] ), .SEL(n5942), 
        .F(n3980) );
  MUX U6139 ( .IN0(reg_dest_new[25]), .IN1(\registers[30][25] ), .SEL(n5942), 
        .F(n3979) );
  MUX U6140 ( .IN0(reg_dest_new[24]), .IN1(\registers[30][24] ), .SEL(n5942), 
        .F(n3978) );
  MUX U6141 ( .IN0(reg_dest_new[23]), .IN1(\registers[30][23] ), .SEL(n5942), 
        .F(n3977) );
  MUX U6142 ( .IN0(reg_dest_new[22]), .IN1(\registers[30][22] ), .SEL(n5942), 
        .F(n3976) );
  MUX U6143 ( .IN0(reg_dest_new[21]), .IN1(\registers[30][21] ), .SEL(n5942), 
        .F(n3975) );
  MUX U6144 ( .IN0(reg_dest_new[20]), .IN1(\registers[30][20] ), .SEL(n5942), 
        .F(n3974) );
  MUX U6145 ( .IN0(reg_dest_new[19]), .IN1(\registers[30][19] ), .SEL(n5942), 
        .F(n3973) );
  MUX U6146 ( .IN0(reg_dest_new[18]), .IN1(\registers[30][18] ), .SEL(n5942), 
        .F(n3972) );
  MUX U6147 ( .IN0(reg_dest_new[17]), .IN1(\registers[30][17] ), .SEL(n5942), 
        .F(n3971) );
  MUX U6148 ( .IN0(reg_dest_new[16]), .IN1(\registers[30][16] ), .SEL(n5942), 
        .F(n3970) );
  MUX U6149 ( .IN0(reg_dest_new[15]), .IN1(\registers[30][15] ), .SEL(n5942), 
        .F(n3969) );
  MUX U6150 ( .IN0(reg_dest_new[14]), .IN1(\registers[30][14] ), .SEL(n5942), 
        .F(n3968) );
  MUX U6151 ( .IN0(reg_dest_new[13]), .IN1(\registers[30][13] ), .SEL(n5942), 
        .F(n3967) );
  MUX U6152 ( .IN0(reg_dest_new[12]), .IN1(\registers[30][12] ), .SEL(n5942), 
        .F(n3966) );
  MUX U6153 ( .IN0(reg_dest_new[11]), .IN1(\registers[30][11] ), .SEL(n5942), 
        .F(n3965) );
  MUX U6154 ( .IN0(reg_dest_new[10]), .IN1(\registers[30][10] ), .SEL(n5942), 
        .F(n3964) );
  MUX U6155 ( .IN0(reg_dest_new[9]), .IN1(\registers[30][9] ), .SEL(n5942), 
        .F(n3963) );
  MUX U6156 ( .IN0(reg_dest_new[8]), .IN1(\registers[30][8] ), .SEL(n5942), 
        .F(n3962) );
  MUX U6157 ( .IN0(reg_dest_new[7]), .IN1(\registers[30][7] ), .SEL(n5942), 
        .F(n3961) );
  MUX U6158 ( .IN0(reg_dest_new[6]), .IN1(\registers[30][6] ), .SEL(n5942), 
        .F(n3960) );
  MUX U6159 ( .IN0(reg_dest_new[5]), .IN1(\registers[30][5] ), .SEL(n5942), 
        .F(n3959) );
  MUX U6160 ( .IN0(reg_dest_new[4]), .IN1(\registers[30][4] ), .SEL(n5942), 
        .F(n3958) );
  MUX U6161 ( .IN0(reg_dest_new[3]), .IN1(\registers[30][3] ), .SEL(n5942), 
        .F(n3957) );
  MUX U6162 ( .IN0(reg_dest_new[2]), .IN1(\registers[30][2] ), .SEL(n5942), 
        .F(n3956) );
  IV U6163 ( .A(n5943), .Z(n5942) );
  MUX U6164 ( .IN0(\registers[30][1] ), .IN1(reg_dest_new[1]), .SEL(n5943), 
        .F(n3955) );
  MUX U6165 ( .IN0(\registers[30][0] ), .IN1(reg_dest_new[0]), .SEL(n5943), 
        .F(n3954) );
  NOR U6166 ( .A(n5944), .B(n5940), .Z(n5943) );
  MUX U6167 ( .IN0(reg_dest_new[31]), .IN1(\registers[29][31] ), .SEL(n5945), 
        .F(n3953) );
  MUX U6168 ( .IN0(reg_dest_new[30]), .IN1(\registers[29][30] ), .SEL(n5945), 
        .F(n3952) );
  MUX U6169 ( .IN0(reg_dest_new[29]), .IN1(\registers[29][29] ), .SEL(n5945), 
        .F(n3951) );
  MUX U6170 ( .IN0(reg_dest_new[28]), .IN1(\registers[29][28] ), .SEL(n5945), 
        .F(n3950) );
  MUX U6171 ( .IN0(reg_dest_new[27]), .IN1(\registers[29][27] ), .SEL(n5945), 
        .F(n3949) );
  MUX U6172 ( .IN0(reg_dest_new[26]), .IN1(\registers[29][26] ), .SEL(n5945), 
        .F(n3948) );
  MUX U6173 ( .IN0(reg_dest_new[25]), .IN1(\registers[29][25] ), .SEL(n5945), 
        .F(n3947) );
  MUX U6174 ( .IN0(reg_dest_new[24]), .IN1(\registers[29][24] ), .SEL(n5945), 
        .F(n3946) );
  MUX U6175 ( .IN0(reg_dest_new[23]), .IN1(\registers[29][23] ), .SEL(n5945), 
        .F(n3945) );
  MUX U6176 ( .IN0(reg_dest_new[22]), .IN1(\registers[29][22] ), .SEL(n5945), 
        .F(n3944) );
  MUX U6177 ( .IN0(reg_dest_new[21]), .IN1(\registers[29][21] ), .SEL(n5945), 
        .F(n3943) );
  MUX U6178 ( .IN0(reg_dest_new[20]), .IN1(\registers[29][20] ), .SEL(n5945), 
        .F(n3942) );
  MUX U6179 ( .IN0(reg_dest_new[19]), .IN1(\registers[29][19] ), .SEL(n5945), 
        .F(n3941) );
  MUX U6180 ( .IN0(reg_dest_new[18]), .IN1(\registers[29][18] ), .SEL(n5945), 
        .F(n3940) );
  MUX U6181 ( .IN0(reg_dest_new[17]), .IN1(\registers[29][17] ), .SEL(n5945), 
        .F(n3939) );
  MUX U6182 ( .IN0(reg_dest_new[16]), .IN1(\registers[29][16] ), .SEL(n5945), 
        .F(n3938) );
  MUX U6183 ( .IN0(reg_dest_new[15]), .IN1(\registers[29][15] ), .SEL(n5945), 
        .F(n3937) );
  MUX U6184 ( .IN0(reg_dest_new[14]), .IN1(\registers[29][14] ), .SEL(n5945), 
        .F(n3936) );
  MUX U6185 ( .IN0(reg_dest_new[13]), .IN1(\registers[29][13] ), .SEL(n5945), 
        .F(n3935) );
  MUX U6186 ( .IN0(reg_dest_new[12]), .IN1(\registers[29][12] ), .SEL(n5945), 
        .F(n3934) );
  MUX U6187 ( .IN0(reg_dest_new[11]), .IN1(\registers[29][11] ), .SEL(n5945), 
        .F(n3933) );
  MUX U6188 ( .IN0(reg_dest_new[10]), .IN1(\registers[29][10] ), .SEL(n5945), 
        .F(n3932) );
  MUX U6189 ( .IN0(reg_dest_new[9]), .IN1(\registers[29][9] ), .SEL(n5945), 
        .F(n3931) );
  MUX U6190 ( .IN0(reg_dest_new[8]), .IN1(\registers[29][8] ), .SEL(n5945), 
        .F(n3930) );
  MUX U6191 ( .IN0(reg_dest_new[7]), .IN1(\registers[29][7] ), .SEL(n5945), 
        .F(n3929) );
  MUX U6192 ( .IN0(reg_dest_new[6]), .IN1(\registers[29][6] ), .SEL(n5945), 
        .F(n3928) );
  MUX U6193 ( .IN0(reg_dest_new[5]), .IN1(\registers[29][5] ), .SEL(n5945), 
        .F(n3927) );
  MUX U6194 ( .IN0(reg_dest_new[4]), .IN1(\registers[29][4] ), .SEL(n5945), 
        .F(n3926) );
  MUX U6195 ( .IN0(reg_dest_new[3]), .IN1(\registers[29][3] ), .SEL(n5945), 
        .F(n3925) );
  MUX U6196 ( .IN0(reg_dest_new[2]), .IN1(\registers[29][2] ), .SEL(n5945), 
        .F(n3924) );
  IV U6197 ( .A(n5946), .Z(n5945) );
  MUX U6198 ( .IN0(\registers[29][1] ), .IN1(reg_dest_new[1]), .SEL(n5946), 
        .F(n3923) );
  MUX U6199 ( .IN0(\registers[29][0] ), .IN1(reg_dest_new[0]), .SEL(n5946), 
        .F(n3922) );
  NOR U6200 ( .A(n5947), .B(n5940), .Z(n5946) );
  MUX U6201 ( .IN0(reg_dest_new[31]), .IN1(\registers[28][31] ), .SEL(n5948), 
        .F(n3921) );
  MUX U6202 ( .IN0(reg_dest_new[30]), .IN1(\registers[28][30] ), .SEL(n5948), 
        .F(n3920) );
  MUX U6203 ( .IN0(reg_dest_new[29]), .IN1(\registers[28][29] ), .SEL(n5948), 
        .F(n3919) );
  MUX U6204 ( .IN0(reg_dest_new[28]), .IN1(\registers[28][28] ), .SEL(n5948), 
        .F(n3918) );
  MUX U6205 ( .IN0(reg_dest_new[27]), .IN1(\registers[28][27] ), .SEL(n5948), 
        .F(n3917) );
  MUX U6206 ( .IN0(reg_dest_new[26]), .IN1(\registers[28][26] ), .SEL(n5948), 
        .F(n3916) );
  MUX U6207 ( .IN0(reg_dest_new[25]), .IN1(\registers[28][25] ), .SEL(n5948), 
        .F(n3915) );
  MUX U6208 ( .IN0(reg_dest_new[24]), .IN1(\registers[28][24] ), .SEL(n5948), 
        .F(n3914) );
  MUX U6209 ( .IN0(reg_dest_new[23]), .IN1(\registers[28][23] ), .SEL(n5948), 
        .F(n3913) );
  MUX U6210 ( .IN0(reg_dest_new[22]), .IN1(\registers[28][22] ), .SEL(n5948), 
        .F(n3912) );
  MUX U6211 ( .IN0(reg_dest_new[21]), .IN1(\registers[28][21] ), .SEL(n5948), 
        .F(n3911) );
  MUX U6212 ( .IN0(reg_dest_new[20]), .IN1(\registers[28][20] ), .SEL(n5948), 
        .F(n3910) );
  MUX U6213 ( .IN0(reg_dest_new[19]), .IN1(\registers[28][19] ), .SEL(n5948), 
        .F(n3909) );
  MUX U6214 ( .IN0(reg_dest_new[18]), .IN1(\registers[28][18] ), .SEL(n5948), 
        .F(n3908) );
  MUX U6215 ( .IN0(reg_dest_new[17]), .IN1(\registers[28][17] ), .SEL(n5948), 
        .F(n3907) );
  MUX U6216 ( .IN0(reg_dest_new[16]), .IN1(\registers[28][16] ), .SEL(n5948), 
        .F(n3906) );
  MUX U6217 ( .IN0(reg_dest_new[15]), .IN1(\registers[28][15] ), .SEL(n5948), 
        .F(n3905) );
  MUX U6218 ( .IN0(reg_dest_new[14]), .IN1(\registers[28][14] ), .SEL(n5948), 
        .F(n3904) );
  MUX U6219 ( .IN0(reg_dest_new[13]), .IN1(\registers[28][13] ), .SEL(n5948), 
        .F(n3903) );
  MUX U6220 ( .IN0(reg_dest_new[12]), .IN1(\registers[28][12] ), .SEL(n5948), 
        .F(n3902) );
  MUX U6221 ( .IN0(reg_dest_new[11]), .IN1(\registers[28][11] ), .SEL(n5948), 
        .F(n3901) );
  MUX U6222 ( .IN0(reg_dest_new[10]), .IN1(\registers[28][10] ), .SEL(n5948), 
        .F(n3900) );
  MUX U6223 ( .IN0(reg_dest_new[9]), .IN1(\registers[28][9] ), .SEL(n5948), 
        .F(n3899) );
  MUX U6224 ( .IN0(reg_dest_new[8]), .IN1(\registers[28][8] ), .SEL(n5948), 
        .F(n3898) );
  MUX U6225 ( .IN0(reg_dest_new[7]), .IN1(\registers[28][7] ), .SEL(n5948), 
        .F(n3897) );
  MUX U6226 ( .IN0(reg_dest_new[6]), .IN1(\registers[28][6] ), .SEL(n5948), 
        .F(n3896) );
  MUX U6227 ( .IN0(reg_dest_new[5]), .IN1(\registers[28][5] ), .SEL(n5948), 
        .F(n3895) );
  MUX U6228 ( .IN0(reg_dest_new[4]), .IN1(\registers[28][4] ), .SEL(n5948), 
        .F(n3894) );
  MUX U6229 ( .IN0(reg_dest_new[3]), .IN1(\registers[28][3] ), .SEL(n5948), 
        .F(n3893) );
  MUX U6230 ( .IN0(reg_dest_new[2]), .IN1(\registers[28][2] ), .SEL(n5948), 
        .F(n3892) );
  IV U6231 ( .A(n5949), .Z(n5948) );
  MUX U6232 ( .IN0(\registers[28][1] ), .IN1(reg_dest_new[1]), .SEL(n5949), 
        .F(n3891) );
  MUX U6233 ( .IN0(\registers[28][0] ), .IN1(reg_dest_new[0]), .SEL(n5949), 
        .F(n3890) );
  NOR U6234 ( .A(n5950), .B(n5940), .Z(n5949) );
  MUX U6235 ( .IN0(reg_dest_new[31]), .IN1(\registers[27][31] ), .SEL(n5951), 
        .F(n3889) );
  MUX U6236 ( .IN0(reg_dest_new[30]), .IN1(\registers[27][30] ), .SEL(n5951), 
        .F(n3888) );
  MUX U6237 ( .IN0(reg_dest_new[29]), .IN1(\registers[27][29] ), .SEL(n5951), 
        .F(n3887) );
  MUX U6238 ( .IN0(reg_dest_new[28]), .IN1(\registers[27][28] ), .SEL(n5951), 
        .F(n3886) );
  MUX U6239 ( .IN0(reg_dest_new[27]), .IN1(\registers[27][27] ), .SEL(n5951), 
        .F(n3885) );
  MUX U6240 ( .IN0(reg_dest_new[26]), .IN1(\registers[27][26] ), .SEL(n5951), 
        .F(n3884) );
  MUX U6241 ( .IN0(reg_dest_new[25]), .IN1(\registers[27][25] ), .SEL(n5951), 
        .F(n3883) );
  MUX U6242 ( .IN0(reg_dest_new[24]), .IN1(\registers[27][24] ), .SEL(n5951), 
        .F(n3882) );
  MUX U6243 ( .IN0(reg_dest_new[23]), .IN1(\registers[27][23] ), .SEL(n5951), 
        .F(n3881) );
  MUX U6244 ( .IN0(reg_dest_new[22]), .IN1(\registers[27][22] ), .SEL(n5951), 
        .F(n3880) );
  MUX U6245 ( .IN0(reg_dest_new[21]), .IN1(\registers[27][21] ), .SEL(n5951), 
        .F(n3879) );
  MUX U6246 ( .IN0(reg_dest_new[20]), .IN1(\registers[27][20] ), .SEL(n5951), 
        .F(n3878) );
  MUX U6247 ( .IN0(reg_dest_new[19]), .IN1(\registers[27][19] ), .SEL(n5951), 
        .F(n3877) );
  MUX U6248 ( .IN0(reg_dest_new[18]), .IN1(\registers[27][18] ), .SEL(n5951), 
        .F(n3876) );
  MUX U6249 ( .IN0(reg_dest_new[17]), .IN1(\registers[27][17] ), .SEL(n5951), 
        .F(n3875) );
  MUX U6250 ( .IN0(reg_dest_new[16]), .IN1(\registers[27][16] ), .SEL(n5951), 
        .F(n3874) );
  MUX U6251 ( .IN0(reg_dest_new[15]), .IN1(\registers[27][15] ), .SEL(n5951), 
        .F(n3873) );
  MUX U6252 ( .IN0(reg_dest_new[14]), .IN1(\registers[27][14] ), .SEL(n5951), 
        .F(n3872) );
  MUX U6253 ( .IN0(reg_dest_new[13]), .IN1(\registers[27][13] ), .SEL(n5951), 
        .F(n3871) );
  MUX U6254 ( .IN0(reg_dest_new[12]), .IN1(\registers[27][12] ), .SEL(n5951), 
        .F(n3870) );
  MUX U6255 ( .IN0(reg_dest_new[11]), .IN1(\registers[27][11] ), .SEL(n5951), 
        .F(n3869) );
  MUX U6256 ( .IN0(reg_dest_new[10]), .IN1(\registers[27][10] ), .SEL(n5951), 
        .F(n3868) );
  MUX U6257 ( .IN0(reg_dest_new[9]), .IN1(\registers[27][9] ), .SEL(n5951), 
        .F(n3867) );
  MUX U6258 ( .IN0(reg_dest_new[8]), .IN1(\registers[27][8] ), .SEL(n5951), 
        .F(n3866) );
  MUX U6259 ( .IN0(reg_dest_new[7]), .IN1(\registers[27][7] ), .SEL(n5951), 
        .F(n3865) );
  MUX U6260 ( .IN0(reg_dest_new[6]), .IN1(\registers[27][6] ), .SEL(n5951), 
        .F(n3864) );
  MUX U6261 ( .IN0(reg_dest_new[5]), .IN1(\registers[27][5] ), .SEL(n5951), 
        .F(n3863) );
  MUX U6262 ( .IN0(reg_dest_new[4]), .IN1(\registers[27][4] ), .SEL(n5951), 
        .F(n3862) );
  MUX U6263 ( .IN0(reg_dest_new[3]), .IN1(\registers[27][3] ), .SEL(n5951), 
        .F(n3861) );
  MUX U6264 ( .IN0(reg_dest_new[2]), .IN1(\registers[27][2] ), .SEL(n5951), 
        .F(n3860) );
  IV U6265 ( .A(n5952), .Z(n5951) );
  MUX U6266 ( .IN0(\registers[27][1] ), .IN1(reg_dest_new[1]), .SEL(n5952), 
        .F(n3859) );
  MUX U6267 ( .IN0(\registers[27][0] ), .IN1(reg_dest_new[0]), .SEL(n5952), 
        .F(n3858) );
  NOR U6268 ( .A(n5953), .B(n5940), .Z(n5952) );
  MUX U6269 ( .IN0(reg_dest_new[31]), .IN1(\registers[26][31] ), .SEL(n5954), 
        .F(n3857) );
  MUX U6270 ( .IN0(reg_dest_new[30]), .IN1(\registers[26][30] ), .SEL(n5954), 
        .F(n3856) );
  MUX U6271 ( .IN0(reg_dest_new[29]), .IN1(\registers[26][29] ), .SEL(n5954), 
        .F(n3855) );
  MUX U6272 ( .IN0(reg_dest_new[28]), .IN1(\registers[26][28] ), .SEL(n5954), 
        .F(n3854) );
  MUX U6273 ( .IN0(reg_dest_new[27]), .IN1(\registers[26][27] ), .SEL(n5954), 
        .F(n3853) );
  MUX U6274 ( .IN0(reg_dest_new[26]), .IN1(\registers[26][26] ), .SEL(n5954), 
        .F(n3852) );
  MUX U6275 ( .IN0(reg_dest_new[25]), .IN1(\registers[26][25] ), .SEL(n5954), 
        .F(n3851) );
  MUX U6276 ( .IN0(reg_dest_new[24]), .IN1(\registers[26][24] ), .SEL(n5954), 
        .F(n3850) );
  MUX U6277 ( .IN0(reg_dest_new[23]), .IN1(\registers[26][23] ), .SEL(n5954), 
        .F(n3849) );
  MUX U6278 ( .IN0(reg_dest_new[22]), .IN1(\registers[26][22] ), .SEL(n5954), 
        .F(n3848) );
  MUX U6279 ( .IN0(reg_dest_new[21]), .IN1(\registers[26][21] ), .SEL(n5954), 
        .F(n3847) );
  MUX U6280 ( .IN0(reg_dest_new[20]), .IN1(\registers[26][20] ), .SEL(n5954), 
        .F(n3846) );
  MUX U6281 ( .IN0(reg_dest_new[19]), .IN1(\registers[26][19] ), .SEL(n5954), 
        .F(n3845) );
  MUX U6282 ( .IN0(reg_dest_new[18]), .IN1(\registers[26][18] ), .SEL(n5954), 
        .F(n3844) );
  MUX U6283 ( .IN0(reg_dest_new[17]), .IN1(\registers[26][17] ), .SEL(n5954), 
        .F(n3843) );
  MUX U6284 ( .IN0(reg_dest_new[16]), .IN1(\registers[26][16] ), .SEL(n5954), 
        .F(n3842) );
  MUX U6285 ( .IN0(reg_dest_new[15]), .IN1(\registers[26][15] ), .SEL(n5954), 
        .F(n3841) );
  MUX U6286 ( .IN0(reg_dest_new[14]), .IN1(\registers[26][14] ), .SEL(n5954), 
        .F(n3840) );
  MUX U6287 ( .IN0(reg_dest_new[13]), .IN1(\registers[26][13] ), .SEL(n5954), 
        .F(n3839) );
  MUX U6288 ( .IN0(reg_dest_new[12]), .IN1(\registers[26][12] ), .SEL(n5954), 
        .F(n3838) );
  MUX U6289 ( .IN0(reg_dest_new[11]), .IN1(\registers[26][11] ), .SEL(n5954), 
        .F(n3837) );
  MUX U6290 ( .IN0(reg_dest_new[10]), .IN1(\registers[26][10] ), .SEL(n5954), 
        .F(n3836) );
  MUX U6291 ( .IN0(reg_dest_new[9]), .IN1(\registers[26][9] ), .SEL(n5954), 
        .F(n3835) );
  MUX U6292 ( .IN0(reg_dest_new[8]), .IN1(\registers[26][8] ), .SEL(n5954), 
        .F(n3834) );
  MUX U6293 ( .IN0(reg_dest_new[7]), .IN1(\registers[26][7] ), .SEL(n5954), 
        .F(n3833) );
  MUX U6294 ( .IN0(reg_dest_new[6]), .IN1(\registers[26][6] ), .SEL(n5954), 
        .F(n3832) );
  MUX U6295 ( .IN0(reg_dest_new[5]), .IN1(\registers[26][5] ), .SEL(n5954), 
        .F(n3831) );
  MUX U6296 ( .IN0(reg_dest_new[4]), .IN1(\registers[26][4] ), .SEL(n5954), 
        .F(n3830) );
  MUX U6297 ( .IN0(reg_dest_new[3]), .IN1(\registers[26][3] ), .SEL(n5954), 
        .F(n3829) );
  MUX U6298 ( .IN0(reg_dest_new[2]), .IN1(\registers[26][2] ), .SEL(n5954), 
        .F(n3828) );
  IV U6299 ( .A(n5955), .Z(n5954) );
  MUX U6300 ( .IN0(\registers[26][1] ), .IN1(reg_dest_new[1]), .SEL(n5955), 
        .F(n3827) );
  MUX U6301 ( .IN0(\registers[26][0] ), .IN1(reg_dest_new[0]), .SEL(n5955), 
        .F(n3826) );
  NOR U6302 ( .A(n5956), .B(n5940), .Z(n5955) );
  MUX U6303 ( .IN0(reg_dest_new[31]), .IN1(\registers[25][31] ), .SEL(n5957), 
        .F(n3825) );
  MUX U6304 ( .IN0(reg_dest_new[30]), .IN1(\registers[25][30] ), .SEL(n5957), 
        .F(n3824) );
  MUX U6305 ( .IN0(reg_dest_new[29]), .IN1(\registers[25][29] ), .SEL(n5957), 
        .F(n3823) );
  MUX U6306 ( .IN0(reg_dest_new[28]), .IN1(\registers[25][28] ), .SEL(n5957), 
        .F(n3822) );
  MUX U6307 ( .IN0(reg_dest_new[27]), .IN1(\registers[25][27] ), .SEL(n5957), 
        .F(n3821) );
  MUX U6308 ( .IN0(reg_dest_new[26]), .IN1(\registers[25][26] ), .SEL(n5957), 
        .F(n3820) );
  MUX U6309 ( .IN0(reg_dest_new[25]), .IN1(\registers[25][25] ), .SEL(n5957), 
        .F(n3819) );
  MUX U6310 ( .IN0(reg_dest_new[24]), .IN1(\registers[25][24] ), .SEL(n5957), 
        .F(n3818) );
  MUX U6311 ( .IN0(reg_dest_new[23]), .IN1(\registers[25][23] ), .SEL(n5957), 
        .F(n3817) );
  MUX U6312 ( .IN0(reg_dest_new[22]), .IN1(\registers[25][22] ), .SEL(n5957), 
        .F(n3816) );
  MUX U6313 ( .IN0(reg_dest_new[21]), .IN1(\registers[25][21] ), .SEL(n5957), 
        .F(n3815) );
  MUX U6314 ( .IN0(reg_dest_new[20]), .IN1(\registers[25][20] ), .SEL(n5957), 
        .F(n3814) );
  MUX U6315 ( .IN0(reg_dest_new[19]), .IN1(\registers[25][19] ), .SEL(n5957), 
        .F(n3813) );
  MUX U6316 ( .IN0(reg_dest_new[18]), .IN1(\registers[25][18] ), .SEL(n5957), 
        .F(n3812) );
  MUX U6317 ( .IN0(reg_dest_new[17]), .IN1(\registers[25][17] ), .SEL(n5957), 
        .F(n3811) );
  MUX U6318 ( .IN0(reg_dest_new[16]), .IN1(\registers[25][16] ), .SEL(n5957), 
        .F(n3810) );
  MUX U6319 ( .IN0(reg_dest_new[15]), .IN1(\registers[25][15] ), .SEL(n5957), 
        .F(n3809) );
  MUX U6320 ( .IN0(reg_dest_new[14]), .IN1(\registers[25][14] ), .SEL(n5957), 
        .F(n3808) );
  MUX U6321 ( .IN0(reg_dest_new[13]), .IN1(\registers[25][13] ), .SEL(n5957), 
        .F(n3807) );
  MUX U6322 ( .IN0(reg_dest_new[12]), .IN1(\registers[25][12] ), .SEL(n5957), 
        .F(n3806) );
  MUX U6323 ( .IN0(reg_dest_new[11]), .IN1(\registers[25][11] ), .SEL(n5957), 
        .F(n3805) );
  MUX U6324 ( .IN0(reg_dest_new[10]), .IN1(\registers[25][10] ), .SEL(n5957), 
        .F(n3804) );
  MUX U6325 ( .IN0(reg_dest_new[9]), .IN1(\registers[25][9] ), .SEL(n5957), 
        .F(n3803) );
  MUX U6326 ( .IN0(reg_dest_new[8]), .IN1(\registers[25][8] ), .SEL(n5957), 
        .F(n3802) );
  MUX U6327 ( .IN0(reg_dest_new[7]), .IN1(\registers[25][7] ), .SEL(n5957), 
        .F(n3801) );
  MUX U6328 ( .IN0(reg_dest_new[6]), .IN1(\registers[25][6] ), .SEL(n5957), 
        .F(n3800) );
  MUX U6329 ( .IN0(reg_dest_new[5]), .IN1(\registers[25][5] ), .SEL(n5957), 
        .F(n3799) );
  MUX U6330 ( .IN0(reg_dest_new[4]), .IN1(\registers[25][4] ), .SEL(n5957), 
        .F(n3798) );
  MUX U6331 ( .IN0(reg_dest_new[3]), .IN1(\registers[25][3] ), .SEL(n5957), 
        .F(n3797) );
  MUX U6332 ( .IN0(reg_dest_new[2]), .IN1(\registers[25][2] ), .SEL(n5957), 
        .F(n3796) );
  IV U6333 ( .A(n5958), .Z(n5957) );
  MUX U6334 ( .IN0(\registers[25][1] ), .IN1(reg_dest_new[1]), .SEL(n5958), 
        .F(n3795) );
  MUX U6335 ( .IN0(\registers[25][0] ), .IN1(reg_dest_new[0]), .SEL(n5958), 
        .F(n3794) );
  NOR U6336 ( .A(n5959), .B(n5940), .Z(n5958) );
  MUX U6337 ( .IN0(reg_dest_new[31]), .IN1(\registers[24][31] ), .SEL(n5960), 
        .F(n3793) );
  MUX U6338 ( .IN0(reg_dest_new[30]), .IN1(\registers[24][30] ), .SEL(n5960), 
        .F(n3792) );
  MUX U6339 ( .IN0(reg_dest_new[29]), .IN1(\registers[24][29] ), .SEL(n5960), 
        .F(n3791) );
  MUX U6340 ( .IN0(reg_dest_new[28]), .IN1(\registers[24][28] ), .SEL(n5960), 
        .F(n3790) );
  MUX U6341 ( .IN0(reg_dest_new[27]), .IN1(\registers[24][27] ), .SEL(n5960), 
        .F(n3789) );
  MUX U6342 ( .IN0(reg_dest_new[26]), .IN1(\registers[24][26] ), .SEL(n5960), 
        .F(n3788) );
  MUX U6343 ( .IN0(reg_dest_new[25]), .IN1(\registers[24][25] ), .SEL(n5960), 
        .F(n3787) );
  MUX U6344 ( .IN0(reg_dest_new[24]), .IN1(\registers[24][24] ), .SEL(n5960), 
        .F(n3786) );
  MUX U6345 ( .IN0(reg_dest_new[23]), .IN1(\registers[24][23] ), .SEL(n5960), 
        .F(n3785) );
  MUX U6346 ( .IN0(reg_dest_new[22]), .IN1(\registers[24][22] ), .SEL(n5960), 
        .F(n3784) );
  MUX U6347 ( .IN0(reg_dest_new[21]), .IN1(\registers[24][21] ), .SEL(n5960), 
        .F(n3783) );
  MUX U6348 ( .IN0(reg_dest_new[20]), .IN1(\registers[24][20] ), .SEL(n5960), 
        .F(n3782) );
  MUX U6349 ( .IN0(reg_dest_new[19]), .IN1(\registers[24][19] ), .SEL(n5960), 
        .F(n3781) );
  MUX U6350 ( .IN0(reg_dest_new[18]), .IN1(\registers[24][18] ), .SEL(n5960), 
        .F(n3780) );
  MUX U6351 ( .IN0(reg_dest_new[17]), .IN1(\registers[24][17] ), .SEL(n5960), 
        .F(n3779) );
  MUX U6352 ( .IN0(reg_dest_new[16]), .IN1(\registers[24][16] ), .SEL(n5960), 
        .F(n3778) );
  MUX U6353 ( .IN0(reg_dest_new[15]), .IN1(\registers[24][15] ), .SEL(n5960), 
        .F(n3777) );
  MUX U6354 ( .IN0(reg_dest_new[14]), .IN1(\registers[24][14] ), .SEL(n5960), 
        .F(n3776) );
  MUX U6355 ( .IN0(reg_dest_new[13]), .IN1(\registers[24][13] ), .SEL(n5960), 
        .F(n3775) );
  MUX U6356 ( .IN0(reg_dest_new[12]), .IN1(\registers[24][12] ), .SEL(n5960), 
        .F(n3774) );
  MUX U6357 ( .IN0(reg_dest_new[11]), .IN1(\registers[24][11] ), .SEL(n5960), 
        .F(n3773) );
  MUX U6358 ( .IN0(reg_dest_new[10]), .IN1(\registers[24][10] ), .SEL(n5960), 
        .F(n3772) );
  MUX U6359 ( .IN0(reg_dest_new[9]), .IN1(\registers[24][9] ), .SEL(n5960), 
        .F(n3771) );
  MUX U6360 ( .IN0(reg_dest_new[8]), .IN1(\registers[24][8] ), .SEL(n5960), 
        .F(n3770) );
  MUX U6361 ( .IN0(reg_dest_new[7]), .IN1(\registers[24][7] ), .SEL(n5960), 
        .F(n3769) );
  MUX U6362 ( .IN0(reg_dest_new[6]), .IN1(\registers[24][6] ), .SEL(n5960), 
        .F(n3768) );
  MUX U6363 ( .IN0(reg_dest_new[5]), .IN1(\registers[24][5] ), .SEL(n5960), 
        .F(n3767) );
  MUX U6364 ( .IN0(reg_dest_new[4]), .IN1(\registers[24][4] ), .SEL(n5960), 
        .F(n3766) );
  MUX U6365 ( .IN0(reg_dest_new[3]), .IN1(\registers[24][3] ), .SEL(n5960), 
        .F(n3765) );
  MUX U6366 ( .IN0(reg_dest_new[2]), .IN1(\registers[24][2] ), .SEL(n5960), 
        .F(n3764) );
  IV U6367 ( .A(n5961), .Z(n5960) );
  MUX U6368 ( .IN0(\registers[24][1] ), .IN1(reg_dest_new[1]), .SEL(n5961), 
        .F(n3763) );
  MUX U6369 ( .IN0(\registers[24][0] ), .IN1(reg_dest_new[0]), .SEL(n5961), 
        .F(n3762) );
  NOR U6370 ( .A(n5962), .B(n5940), .Z(n5961) );
  NANDN U6371 ( .A(n5963), .B(rd_index[4]), .Z(n5940) );
  MUX U6372 ( .IN0(reg_dest_new[31]), .IN1(\registers[23][31] ), .SEL(n5964), 
        .F(n3761) );
  MUX U6373 ( .IN0(reg_dest_new[30]), .IN1(\registers[23][30] ), .SEL(n5964), 
        .F(n3760) );
  MUX U6374 ( .IN0(reg_dest_new[29]), .IN1(\registers[23][29] ), .SEL(n5964), 
        .F(n3759) );
  MUX U6375 ( .IN0(reg_dest_new[28]), .IN1(\registers[23][28] ), .SEL(n5964), 
        .F(n3758) );
  MUX U6376 ( .IN0(reg_dest_new[27]), .IN1(\registers[23][27] ), .SEL(n5964), 
        .F(n3757) );
  MUX U6377 ( .IN0(reg_dest_new[26]), .IN1(\registers[23][26] ), .SEL(n5964), 
        .F(n3756) );
  MUX U6378 ( .IN0(reg_dest_new[25]), .IN1(\registers[23][25] ), .SEL(n5964), 
        .F(n3755) );
  MUX U6379 ( .IN0(reg_dest_new[24]), .IN1(\registers[23][24] ), .SEL(n5964), 
        .F(n3754) );
  MUX U6380 ( .IN0(reg_dest_new[23]), .IN1(\registers[23][23] ), .SEL(n5964), 
        .F(n3753) );
  MUX U6381 ( .IN0(reg_dest_new[22]), .IN1(\registers[23][22] ), .SEL(n5964), 
        .F(n3752) );
  MUX U6382 ( .IN0(reg_dest_new[21]), .IN1(\registers[23][21] ), .SEL(n5964), 
        .F(n3751) );
  MUX U6383 ( .IN0(reg_dest_new[20]), .IN1(\registers[23][20] ), .SEL(n5964), 
        .F(n3750) );
  MUX U6384 ( .IN0(reg_dest_new[19]), .IN1(\registers[23][19] ), .SEL(n5964), 
        .F(n3749) );
  MUX U6385 ( .IN0(reg_dest_new[18]), .IN1(\registers[23][18] ), .SEL(n5964), 
        .F(n3748) );
  MUX U6386 ( .IN0(reg_dest_new[17]), .IN1(\registers[23][17] ), .SEL(n5964), 
        .F(n3747) );
  MUX U6387 ( .IN0(reg_dest_new[16]), .IN1(\registers[23][16] ), .SEL(n5964), 
        .F(n3746) );
  MUX U6388 ( .IN0(reg_dest_new[15]), .IN1(\registers[23][15] ), .SEL(n5964), 
        .F(n3745) );
  MUX U6389 ( .IN0(reg_dest_new[14]), .IN1(\registers[23][14] ), .SEL(n5964), 
        .F(n3744) );
  MUX U6390 ( .IN0(reg_dest_new[13]), .IN1(\registers[23][13] ), .SEL(n5964), 
        .F(n3743) );
  MUX U6391 ( .IN0(reg_dest_new[12]), .IN1(\registers[23][12] ), .SEL(n5964), 
        .F(n3742) );
  MUX U6392 ( .IN0(reg_dest_new[11]), .IN1(\registers[23][11] ), .SEL(n5964), 
        .F(n3741) );
  MUX U6393 ( .IN0(reg_dest_new[10]), .IN1(\registers[23][10] ), .SEL(n5964), 
        .F(n3740) );
  MUX U6394 ( .IN0(reg_dest_new[9]), .IN1(\registers[23][9] ), .SEL(n5964), 
        .F(n3739) );
  MUX U6395 ( .IN0(reg_dest_new[8]), .IN1(\registers[23][8] ), .SEL(n5964), 
        .F(n3738) );
  MUX U6396 ( .IN0(reg_dest_new[7]), .IN1(\registers[23][7] ), .SEL(n5964), 
        .F(n3737) );
  MUX U6397 ( .IN0(reg_dest_new[6]), .IN1(\registers[23][6] ), .SEL(n5964), 
        .F(n3736) );
  MUX U6398 ( .IN0(reg_dest_new[5]), .IN1(\registers[23][5] ), .SEL(n5964), 
        .F(n3735) );
  MUX U6399 ( .IN0(reg_dest_new[4]), .IN1(\registers[23][4] ), .SEL(n5964), 
        .F(n3734) );
  MUX U6400 ( .IN0(reg_dest_new[3]), .IN1(\registers[23][3] ), .SEL(n5964), 
        .F(n3733) );
  MUX U6401 ( .IN0(reg_dest_new[2]), .IN1(\registers[23][2] ), .SEL(n5964), 
        .F(n3732) );
  IV U6402 ( .A(n5965), .Z(n5964) );
  MUX U6403 ( .IN0(\registers[23][1] ), .IN1(reg_dest_new[1]), .SEL(n5965), 
        .F(n3731) );
  MUX U6404 ( .IN0(\registers[23][0] ), .IN1(reg_dest_new[0]), .SEL(n5965), 
        .F(n3730) );
  NOR U6405 ( .A(n5966), .B(n5941), .Z(n5965) );
  MUX U6406 ( .IN0(reg_dest_new[31]), .IN1(\registers[22][31] ), .SEL(n5967), 
        .F(n3729) );
  MUX U6407 ( .IN0(reg_dest_new[30]), .IN1(\registers[22][30] ), .SEL(n5967), 
        .F(n3728) );
  MUX U6408 ( .IN0(reg_dest_new[29]), .IN1(\registers[22][29] ), .SEL(n5967), 
        .F(n3727) );
  MUX U6409 ( .IN0(reg_dest_new[28]), .IN1(\registers[22][28] ), .SEL(n5967), 
        .F(n3726) );
  MUX U6410 ( .IN0(reg_dest_new[27]), .IN1(\registers[22][27] ), .SEL(n5967), 
        .F(n3725) );
  MUX U6411 ( .IN0(reg_dest_new[26]), .IN1(\registers[22][26] ), .SEL(n5967), 
        .F(n3724) );
  MUX U6412 ( .IN0(reg_dest_new[25]), .IN1(\registers[22][25] ), .SEL(n5967), 
        .F(n3723) );
  MUX U6413 ( .IN0(reg_dest_new[24]), .IN1(\registers[22][24] ), .SEL(n5967), 
        .F(n3722) );
  MUX U6414 ( .IN0(reg_dest_new[23]), .IN1(\registers[22][23] ), .SEL(n5967), 
        .F(n3721) );
  MUX U6415 ( .IN0(reg_dest_new[22]), .IN1(\registers[22][22] ), .SEL(n5967), 
        .F(n3720) );
  MUX U6416 ( .IN0(reg_dest_new[21]), .IN1(\registers[22][21] ), .SEL(n5967), 
        .F(n3719) );
  MUX U6417 ( .IN0(reg_dest_new[20]), .IN1(\registers[22][20] ), .SEL(n5967), 
        .F(n3718) );
  MUX U6418 ( .IN0(reg_dest_new[19]), .IN1(\registers[22][19] ), .SEL(n5967), 
        .F(n3717) );
  MUX U6419 ( .IN0(reg_dest_new[18]), .IN1(\registers[22][18] ), .SEL(n5967), 
        .F(n3716) );
  MUX U6420 ( .IN0(reg_dest_new[17]), .IN1(\registers[22][17] ), .SEL(n5967), 
        .F(n3715) );
  MUX U6421 ( .IN0(reg_dest_new[16]), .IN1(\registers[22][16] ), .SEL(n5967), 
        .F(n3714) );
  MUX U6422 ( .IN0(reg_dest_new[15]), .IN1(\registers[22][15] ), .SEL(n5967), 
        .F(n3713) );
  MUX U6423 ( .IN0(reg_dest_new[14]), .IN1(\registers[22][14] ), .SEL(n5967), 
        .F(n3712) );
  MUX U6424 ( .IN0(reg_dest_new[13]), .IN1(\registers[22][13] ), .SEL(n5967), 
        .F(n3711) );
  MUX U6425 ( .IN0(reg_dest_new[12]), .IN1(\registers[22][12] ), .SEL(n5967), 
        .F(n3710) );
  MUX U6426 ( .IN0(reg_dest_new[11]), .IN1(\registers[22][11] ), .SEL(n5967), 
        .F(n3709) );
  MUX U6427 ( .IN0(reg_dest_new[10]), .IN1(\registers[22][10] ), .SEL(n5967), 
        .F(n3708) );
  MUX U6428 ( .IN0(reg_dest_new[9]), .IN1(\registers[22][9] ), .SEL(n5967), 
        .F(n3707) );
  MUX U6429 ( .IN0(reg_dest_new[8]), .IN1(\registers[22][8] ), .SEL(n5967), 
        .F(n3706) );
  MUX U6430 ( .IN0(reg_dest_new[7]), .IN1(\registers[22][7] ), .SEL(n5967), 
        .F(n3705) );
  MUX U6431 ( .IN0(reg_dest_new[6]), .IN1(\registers[22][6] ), .SEL(n5967), 
        .F(n3704) );
  MUX U6432 ( .IN0(reg_dest_new[5]), .IN1(\registers[22][5] ), .SEL(n5967), 
        .F(n3703) );
  MUX U6433 ( .IN0(reg_dest_new[4]), .IN1(\registers[22][4] ), .SEL(n5967), 
        .F(n3702) );
  MUX U6434 ( .IN0(reg_dest_new[3]), .IN1(\registers[22][3] ), .SEL(n5967), 
        .F(n3701) );
  MUX U6435 ( .IN0(reg_dest_new[2]), .IN1(\registers[22][2] ), .SEL(n5967), 
        .F(n3700) );
  IV U6436 ( .A(n5968), .Z(n5967) );
  MUX U6437 ( .IN0(\registers[22][1] ), .IN1(reg_dest_new[1]), .SEL(n5968), 
        .F(n3699) );
  MUX U6438 ( .IN0(\registers[22][0] ), .IN1(reg_dest_new[0]), .SEL(n5968), 
        .F(n3698) );
  NOR U6439 ( .A(n5966), .B(n5944), .Z(n5968) );
  MUX U6440 ( .IN0(reg_dest_new[31]), .IN1(\registers[21][31] ), .SEL(n5969), 
        .F(n3697) );
  MUX U6441 ( .IN0(reg_dest_new[30]), .IN1(\registers[21][30] ), .SEL(n5969), 
        .F(n3696) );
  MUX U6442 ( .IN0(reg_dest_new[29]), .IN1(\registers[21][29] ), .SEL(n5969), 
        .F(n3695) );
  MUX U6443 ( .IN0(reg_dest_new[28]), .IN1(\registers[21][28] ), .SEL(n5969), 
        .F(n3694) );
  MUX U6444 ( .IN0(reg_dest_new[27]), .IN1(\registers[21][27] ), .SEL(n5969), 
        .F(n3693) );
  MUX U6445 ( .IN0(reg_dest_new[26]), .IN1(\registers[21][26] ), .SEL(n5969), 
        .F(n3692) );
  MUX U6446 ( .IN0(reg_dest_new[25]), .IN1(\registers[21][25] ), .SEL(n5969), 
        .F(n3691) );
  MUX U6447 ( .IN0(reg_dest_new[24]), .IN1(\registers[21][24] ), .SEL(n5969), 
        .F(n3690) );
  MUX U6448 ( .IN0(reg_dest_new[23]), .IN1(\registers[21][23] ), .SEL(n5969), 
        .F(n3689) );
  MUX U6449 ( .IN0(reg_dest_new[22]), .IN1(\registers[21][22] ), .SEL(n5969), 
        .F(n3688) );
  MUX U6450 ( .IN0(reg_dest_new[21]), .IN1(\registers[21][21] ), .SEL(n5969), 
        .F(n3687) );
  MUX U6451 ( .IN0(reg_dest_new[20]), .IN1(\registers[21][20] ), .SEL(n5969), 
        .F(n3686) );
  MUX U6452 ( .IN0(reg_dest_new[19]), .IN1(\registers[21][19] ), .SEL(n5969), 
        .F(n3685) );
  MUX U6453 ( .IN0(reg_dest_new[18]), .IN1(\registers[21][18] ), .SEL(n5969), 
        .F(n3684) );
  MUX U6454 ( .IN0(reg_dest_new[17]), .IN1(\registers[21][17] ), .SEL(n5969), 
        .F(n3683) );
  MUX U6455 ( .IN0(reg_dest_new[16]), .IN1(\registers[21][16] ), .SEL(n5969), 
        .F(n3682) );
  MUX U6456 ( .IN0(reg_dest_new[15]), .IN1(\registers[21][15] ), .SEL(n5969), 
        .F(n3681) );
  MUX U6457 ( .IN0(reg_dest_new[14]), .IN1(\registers[21][14] ), .SEL(n5969), 
        .F(n3680) );
  MUX U6458 ( .IN0(reg_dest_new[13]), .IN1(\registers[21][13] ), .SEL(n5969), 
        .F(n3679) );
  MUX U6459 ( .IN0(reg_dest_new[12]), .IN1(\registers[21][12] ), .SEL(n5969), 
        .F(n3678) );
  MUX U6460 ( .IN0(reg_dest_new[11]), .IN1(\registers[21][11] ), .SEL(n5969), 
        .F(n3677) );
  MUX U6461 ( .IN0(reg_dest_new[10]), .IN1(\registers[21][10] ), .SEL(n5969), 
        .F(n3676) );
  MUX U6462 ( .IN0(reg_dest_new[9]), .IN1(\registers[21][9] ), .SEL(n5969), 
        .F(n3675) );
  MUX U6463 ( .IN0(reg_dest_new[8]), .IN1(\registers[21][8] ), .SEL(n5969), 
        .F(n3674) );
  MUX U6464 ( .IN0(reg_dest_new[7]), .IN1(\registers[21][7] ), .SEL(n5969), 
        .F(n3673) );
  MUX U6465 ( .IN0(reg_dest_new[6]), .IN1(\registers[21][6] ), .SEL(n5969), 
        .F(n3672) );
  MUX U6466 ( .IN0(reg_dest_new[5]), .IN1(\registers[21][5] ), .SEL(n5969), 
        .F(n3671) );
  MUX U6467 ( .IN0(reg_dest_new[4]), .IN1(\registers[21][4] ), .SEL(n5969), 
        .F(n3670) );
  MUX U6468 ( .IN0(reg_dest_new[3]), .IN1(\registers[21][3] ), .SEL(n5969), 
        .F(n3669) );
  MUX U6469 ( .IN0(reg_dest_new[2]), .IN1(\registers[21][2] ), .SEL(n5969), 
        .F(n3668) );
  IV U6470 ( .A(n5970), .Z(n5969) );
  MUX U6471 ( .IN0(\registers[21][1] ), .IN1(reg_dest_new[1]), .SEL(n5970), 
        .F(n3667) );
  MUX U6472 ( .IN0(\registers[21][0] ), .IN1(reg_dest_new[0]), .SEL(n5970), 
        .F(n3666) );
  NOR U6473 ( .A(n5966), .B(n5947), .Z(n5970) );
  MUX U6474 ( .IN0(reg_dest_new[31]), .IN1(\registers[20][31] ), .SEL(n5971), 
        .F(n3665) );
  MUX U6475 ( .IN0(reg_dest_new[30]), .IN1(\registers[20][30] ), .SEL(n5971), 
        .F(n3664) );
  MUX U6476 ( .IN0(reg_dest_new[29]), .IN1(\registers[20][29] ), .SEL(n5971), 
        .F(n3663) );
  MUX U6477 ( .IN0(reg_dest_new[28]), .IN1(\registers[20][28] ), .SEL(n5971), 
        .F(n3662) );
  MUX U6478 ( .IN0(reg_dest_new[27]), .IN1(\registers[20][27] ), .SEL(n5971), 
        .F(n3661) );
  MUX U6479 ( .IN0(reg_dest_new[26]), .IN1(\registers[20][26] ), .SEL(n5971), 
        .F(n3660) );
  MUX U6480 ( .IN0(reg_dest_new[25]), .IN1(\registers[20][25] ), .SEL(n5971), 
        .F(n3659) );
  MUX U6481 ( .IN0(reg_dest_new[24]), .IN1(\registers[20][24] ), .SEL(n5971), 
        .F(n3658) );
  MUX U6482 ( .IN0(reg_dest_new[23]), .IN1(\registers[20][23] ), .SEL(n5971), 
        .F(n3657) );
  MUX U6483 ( .IN0(reg_dest_new[22]), .IN1(\registers[20][22] ), .SEL(n5971), 
        .F(n3656) );
  MUX U6484 ( .IN0(reg_dest_new[21]), .IN1(\registers[20][21] ), .SEL(n5971), 
        .F(n3655) );
  MUX U6485 ( .IN0(reg_dest_new[20]), .IN1(\registers[20][20] ), .SEL(n5971), 
        .F(n3654) );
  MUX U6486 ( .IN0(reg_dest_new[19]), .IN1(\registers[20][19] ), .SEL(n5971), 
        .F(n3653) );
  MUX U6487 ( .IN0(reg_dest_new[18]), .IN1(\registers[20][18] ), .SEL(n5971), 
        .F(n3652) );
  MUX U6488 ( .IN0(reg_dest_new[17]), .IN1(\registers[20][17] ), .SEL(n5971), 
        .F(n3651) );
  MUX U6489 ( .IN0(reg_dest_new[16]), .IN1(\registers[20][16] ), .SEL(n5971), 
        .F(n3650) );
  MUX U6490 ( .IN0(reg_dest_new[15]), .IN1(\registers[20][15] ), .SEL(n5971), 
        .F(n3649) );
  MUX U6491 ( .IN0(reg_dest_new[14]), .IN1(\registers[20][14] ), .SEL(n5971), 
        .F(n3648) );
  MUX U6492 ( .IN0(reg_dest_new[13]), .IN1(\registers[20][13] ), .SEL(n5971), 
        .F(n3647) );
  MUX U6493 ( .IN0(reg_dest_new[12]), .IN1(\registers[20][12] ), .SEL(n5971), 
        .F(n3646) );
  MUX U6494 ( .IN0(reg_dest_new[11]), .IN1(\registers[20][11] ), .SEL(n5971), 
        .F(n3645) );
  MUX U6495 ( .IN0(reg_dest_new[10]), .IN1(\registers[20][10] ), .SEL(n5971), 
        .F(n3644) );
  MUX U6496 ( .IN0(reg_dest_new[9]), .IN1(\registers[20][9] ), .SEL(n5971), 
        .F(n3643) );
  MUX U6497 ( .IN0(reg_dest_new[8]), .IN1(\registers[20][8] ), .SEL(n5971), 
        .F(n3642) );
  MUX U6498 ( .IN0(reg_dest_new[7]), .IN1(\registers[20][7] ), .SEL(n5971), 
        .F(n3641) );
  MUX U6499 ( .IN0(reg_dest_new[6]), .IN1(\registers[20][6] ), .SEL(n5971), 
        .F(n3640) );
  MUX U6500 ( .IN0(reg_dest_new[5]), .IN1(\registers[20][5] ), .SEL(n5971), 
        .F(n3639) );
  MUX U6501 ( .IN0(reg_dest_new[4]), .IN1(\registers[20][4] ), .SEL(n5971), 
        .F(n3638) );
  MUX U6502 ( .IN0(reg_dest_new[3]), .IN1(\registers[20][3] ), .SEL(n5971), 
        .F(n3637) );
  MUX U6503 ( .IN0(reg_dest_new[2]), .IN1(\registers[20][2] ), .SEL(n5971), 
        .F(n3636) );
  IV U6504 ( .A(n5972), .Z(n5971) );
  MUX U6505 ( .IN0(\registers[20][1] ), .IN1(reg_dest_new[1]), .SEL(n5972), 
        .F(n3635) );
  MUX U6506 ( .IN0(\registers[20][0] ), .IN1(reg_dest_new[0]), .SEL(n5972), 
        .F(n3634) );
  NOR U6507 ( .A(n5966), .B(n5950), .Z(n5972) );
  MUX U6508 ( .IN0(reg_dest_new[31]), .IN1(\registers[19][31] ), .SEL(n5973), 
        .F(n3633) );
  MUX U6509 ( .IN0(reg_dest_new[30]), .IN1(\registers[19][30] ), .SEL(n5973), 
        .F(n3632) );
  MUX U6510 ( .IN0(reg_dest_new[29]), .IN1(\registers[19][29] ), .SEL(n5973), 
        .F(n3631) );
  MUX U6511 ( .IN0(reg_dest_new[28]), .IN1(\registers[19][28] ), .SEL(n5973), 
        .F(n3630) );
  MUX U6512 ( .IN0(reg_dest_new[27]), .IN1(\registers[19][27] ), .SEL(n5973), 
        .F(n3629) );
  MUX U6513 ( .IN0(reg_dest_new[26]), .IN1(\registers[19][26] ), .SEL(n5973), 
        .F(n3628) );
  MUX U6514 ( .IN0(reg_dest_new[25]), .IN1(\registers[19][25] ), .SEL(n5973), 
        .F(n3627) );
  MUX U6515 ( .IN0(reg_dest_new[24]), .IN1(\registers[19][24] ), .SEL(n5973), 
        .F(n3626) );
  MUX U6516 ( .IN0(reg_dest_new[23]), .IN1(\registers[19][23] ), .SEL(n5973), 
        .F(n3625) );
  MUX U6517 ( .IN0(reg_dest_new[22]), .IN1(\registers[19][22] ), .SEL(n5973), 
        .F(n3624) );
  MUX U6518 ( .IN0(reg_dest_new[21]), .IN1(\registers[19][21] ), .SEL(n5973), 
        .F(n3623) );
  MUX U6519 ( .IN0(reg_dest_new[20]), .IN1(\registers[19][20] ), .SEL(n5973), 
        .F(n3622) );
  MUX U6520 ( .IN0(reg_dest_new[19]), .IN1(\registers[19][19] ), .SEL(n5973), 
        .F(n3621) );
  MUX U6521 ( .IN0(reg_dest_new[18]), .IN1(\registers[19][18] ), .SEL(n5973), 
        .F(n3620) );
  MUX U6522 ( .IN0(reg_dest_new[17]), .IN1(\registers[19][17] ), .SEL(n5973), 
        .F(n3619) );
  MUX U6523 ( .IN0(reg_dest_new[16]), .IN1(\registers[19][16] ), .SEL(n5973), 
        .F(n3618) );
  MUX U6524 ( .IN0(reg_dest_new[15]), .IN1(\registers[19][15] ), .SEL(n5973), 
        .F(n3617) );
  MUX U6525 ( .IN0(reg_dest_new[14]), .IN1(\registers[19][14] ), .SEL(n5973), 
        .F(n3616) );
  MUX U6526 ( .IN0(reg_dest_new[13]), .IN1(\registers[19][13] ), .SEL(n5973), 
        .F(n3615) );
  MUX U6527 ( .IN0(reg_dest_new[12]), .IN1(\registers[19][12] ), .SEL(n5973), 
        .F(n3614) );
  MUX U6528 ( .IN0(reg_dest_new[11]), .IN1(\registers[19][11] ), .SEL(n5973), 
        .F(n3613) );
  MUX U6529 ( .IN0(reg_dest_new[10]), .IN1(\registers[19][10] ), .SEL(n5973), 
        .F(n3612) );
  MUX U6530 ( .IN0(reg_dest_new[9]), .IN1(\registers[19][9] ), .SEL(n5973), 
        .F(n3611) );
  MUX U6531 ( .IN0(reg_dest_new[8]), .IN1(\registers[19][8] ), .SEL(n5973), 
        .F(n3610) );
  MUX U6532 ( .IN0(reg_dest_new[7]), .IN1(\registers[19][7] ), .SEL(n5973), 
        .F(n3609) );
  MUX U6533 ( .IN0(reg_dest_new[6]), .IN1(\registers[19][6] ), .SEL(n5973), 
        .F(n3608) );
  MUX U6534 ( .IN0(reg_dest_new[5]), .IN1(\registers[19][5] ), .SEL(n5973), 
        .F(n3607) );
  MUX U6535 ( .IN0(reg_dest_new[4]), .IN1(\registers[19][4] ), .SEL(n5973), 
        .F(n3606) );
  MUX U6536 ( .IN0(reg_dest_new[3]), .IN1(\registers[19][3] ), .SEL(n5973), 
        .F(n3605) );
  MUX U6537 ( .IN0(reg_dest_new[2]), .IN1(\registers[19][2] ), .SEL(n5973), 
        .F(n3604) );
  IV U6538 ( .A(n5974), .Z(n5973) );
  MUX U6539 ( .IN0(\registers[19][1] ), .IN1(reg_dest_new[1]), .SEL(n5974), 
        .F(n3603) );
  MUX U6540 ( .IN0(\registers[19][0] ), .IN1(reg_dest_new[0]), .SEL(n5974), 
        .F(n3602) );
  NOR U6541 ( .A(n5966), .B(n5953), .Z(n5974) );
  MUX U6542 ( .IN0(reg_dest_new[31]), .IN1(\registers[18][31] ), .SEL(n5975), 
        .F(n3601) );
  MUX U6543 ( .IN0(reg_dest_new[30]), .IN1(\registers[18][30] ), .SEL(n5975), 
        .F(n3600) );
  MUX U6544 ( .IN0(reg_dest_new[29]), .IN1(\registers[18][29] ), .SEL(n5975), 
        .F(n3599) );
  MUX U6545 ( .IN0(reg_dest_new[28]), .IN1(\registers[18][28] ), .SEL(n5975), 
        .F(n3598) );
  MUX U6546 ( .IN0(reg_dest_new[27]), .IN1(\registers[18][27] ), .SEL(n5975), 
        .F(n3597) );
  MUX U6547 ( .IN0(reg_dest_new[26]), .IN1(\registers[18][26] ), .SEL(n5975), 
        .F(n3596) );
  MUX U6548 ( .IN0(reg_dest_new[25]), .IN1(\registers[18][25] ), .SEL(n5975), 
        .F(n3595) );
  MUX U6549 ( .IN0(reg_dest_new[24]), .IN1(\registers[18][24] ), .SEL(n5975), 
        .F(n3594) );
  MUX U6550 ( .IN0(reg_dest_new[23]), .IN1(\registers[18][23] ), .SEL(n5975), 
        .F(n3593) );
  MUX U6551 ( .IN0(reg_dest_new[22]), .IN1(\registers[18][22] ), .SEL(n5975), 
        .F(n3592) );
  MUX U6552 ( .IN0(reg_dest_new[21]), .IN1(\registers[18][21] ), .SEL(n5975), 
        .F(n3591) );
  MUX U6553 ( .IN0(reg_dest_new[20]), .IN1(\registers[18][20] ), .SEL(n5975), 
        .F(n3590) );
  MUX U6554 ( .IN0(reg_dest_new[19]), .IN1(\registers[18][19] ), .SEL(n5975), 
        .F(n3589) );
  MUX U6555 ( .IN0(reg_dest_new[18]), .IN1(\registers[18][18] ), .SEL(n5975), 
        .F(n3588) );
  MUX U6556 ( .IN0(reg_dest_new[17]), .IN1(\registers[18][17] ), .SEL(n5975), 
        .F(n3587) );
  MUX U6557 ( .IN0(reg_dest_new[16]), .IN1(\registers[18][16] ), .SEL(n5975), 
        .F(n3586) );
  MUX U6558 ( .IN0(reg_dest_new[15]), .IN1(\registers[18][15] ), .SEL(n5975), 
        .F(n3585) );
  MUX U6559 ( .IN0(reg_dest_new[14]), .IN1(\registers[18][14] ), .SEL(n5975), 
        .F(n3584) );
  MUX U6560 ( .IN0(reg_dest_new[13]), .IN1(\registers[18][13] ), .SEL(n5975), 
        .F(n3583) );
  MUX U6561 ( .IN0(reg_dest_new[12]), .IN1(\registers[18][12] ), .SEL(n5975), 
        .F(n3582) );
  MUX U6562 ( .IN0(reg_dest_new[11]), .IN1(\registers[18][11] ), .SEL(n5975), 
        .F(n3581) );
  MUX U6563 ( .IN0(reg_dest_new[10]), .IN1(\registers[18][10] ), .SEL(n5975), 
        .F(n3580) );
  MUX U6564 ( .IN0(reg_dest_new[9]), .IN1(\registers[18][9] ), .SEL(n5975), 
        .F(n3579) );
  MUX U6565 ( .IN0(reg_dest_new[8]), .IN1(\registers[18][8] ), .SEL(n5975), 
        .F(n3578) );
  MUX U6566 ( .IN0(reg_dest_new[7]), .IN1(\registers[18][7] ), .SEL(n5975), 
        .F(n3577) );
  MUX U6567 ( .IN0(reg_dest_new[6]), .IN1(\registers[18][6] ), .SEL(n5975), 
        .F(n3576) );
  MUX U6568 ( .IN0(reg_dest_new[5]), .IN1(\registers[18][5] ), .SEL(n5975), 
        .F(n3575) );
  MUX U6569 ( .IN0(reg_dest_new[4]), .IN1(\registers[18][4] ), .SEL(n5975), 
        .F(n3574) );
  MUX U6570 ( .IN0(reg_dest_new[3]), .IN1(\registers[18][3] ), .SEL(n5975), 
        .F(n3573) );
  MUX U6571 ( .IN0(reg_dest_new[2]), .IN1(\registers[18][2] ), .SEL(n5975), 
        .F(n3572) );
  IV U6572 ( .A(n5976), .Z(n5975) );
  MUX U6573 ( .IN0(\registers[18][1] ), .IN1(reg_dest_new[1]), .SEL(n5976), 
        .F(n3571) );
  MUX U6574 ( .IN0(\registers[18][0] ), .IN1(reg_dest_new[0]), .SEL(n5976), 
        .F(n3570) );
  NOR U6575 ( .A(n5966), .B(n5956), .Z(n5976) );
  MUX U6576 ( .IN0(reg_dest_new[31]), .IN1(\registers[17][31] ), .SEL(n5977), 
        .F(n3569) );
  MUX U6577 ( .IN0(reg_dest_new[30]), .IN1(\registers[17][30] ), .SEL(n5977), 
        .F(n3568) );
  MUX U6578 ( .IN0(reg_dest_new[29]), .IN1(\registers[17][29] ), .SEL(n5977), 
        .F(n3567) );
  MUX U6579 ( .IN0(reg_dest_new[28]), .IN1(\registers[17][28] ), .SEL(n5977), 
        .F(n3566) );
  MUX U6580 ( .IN0(reg_dest_new[27]), .IN1(\registers[17][27] ), .SEL(n5977), 
        .F(n3565) );
  MUX U6581 ( .IN0(reg_dest_new[26]), .IN1(\registers[17][26] ), .SEL(n5977), 
        .F(n3564) );
  MUX U6582 ( .IN0(reg_dest_new[25]), .IN1(\registers[17][25] ), .SEL(n5977), 
        .F(n3563) );
  MUX U6583 ( .IN0(reg_dest_new[24]), .IN1(\registers[17][24] ), .SEL(n5977), 
        .F(n3562) );
  MUX U6584 ( .IN0(reg_dest_new[23]), .IN1(\registers[17][23] ), .SEL(n5977), 
        .F(n3561) );
  MUX U6585 ( .IN0(reg_dest_new[22]), .IN1(\registers[17][22] ), .SEL(n5977), 
        .F(n3560) );
  MUX U6586 ( .IN0(reg_dest_new[21]), .IN1(\registers[17][21] ), .SEL(n5977), 
        .F(n3559) );
  MUX U6587 ( .IN0(reg_dest_new[20]), .IN1(\registers[17][20] ), .SEL(n5977), 
        .F(n3558) );
  MUX U6588 ( .IN0(reg_dest_new[19]), .IN1(\registers[17][19] ), .SEL(n5977), 
        .F(n3557) );
  MUX U6589 ( .IN0(reg_dest_new[18]), .IN1(\registers[17][18] ), .SEL(n5977), 
        .F(n3556) );
  MUX U6590 ( .IN0(reg_dest_new[17]), .IN1(\registers[17][17] ), .SEL(n5977), 
        .F(n3555) );
  MUX U6591 ( .IN0(reg_dest_new[16]), .IN1(\registers[17][16] ), .SEL(n5977), 
        .F(n3554) );
  MUX U6592 ( .IN0(reg_dest_new[15]), .IN1(\registers[17][15] ), .SEL(n5977), 
        .F(n3553) );
  MUX U6593 ( .IN0(reg_dest_new[14]), .IN1(\registers[17][14] ), .SEL(n5977), 
        .F(n3552) );
  MUX U6594 ( .IN0(reg_dest_new[13]), .IN1(\registers[17][13] ), .SEL(n5977), 
        .F(n3551) );
  MUX U6595 ( .IN0(reg_dest_new[12]), .IN1(\registers[17][12] ), .SEL(n5977), 
        .F(n3550) );
  MUX U6596 ( .IN0(reg_dest_new[11]), .IN1(\registers[17][11] ), .SEL(n5977), 
        .F(n3549) );
  MUX U6597 ( .IN0(reg_dest_new[10]), .IN1(\registers[17][10] ), .SEL(n5977), 
        .F(n3548) );
  MUX U6598 ( .IN0(reg_dest_new[9]), .IN1(\registers[17][9] ), .SEL(n5977), 
        .F(n3547) );
  MUX U6599 ( .IN0(reg_dest_new[8]), .IN1(\registers[17][8] ), .SEL(n5977), 
        .F(n3546) );
  MUX U6600 ( .IN0(reg_dest_new[7]), .IN1(\registers[17][7] ), .SEL(n5977), 
        .F(n3545) );
  MUX U6601 ( .IN0(reg_dest_new[6]), .IN1(\registers[17][6] ), .SEL(n5977), 
        .F(n3544) );
  MUX U6602 ( .IN0(reg_dest_new[5]), .IN1(\registers[17][5] ), .SEL(n5977), 
        .F(n3543) );
  MUX U6603 ( .IN0(reg_dest_new[4]), .IN1(\registers[17][4] ), .SEL(n5977), 
        .F(n3542) );
  MUX U6604 ( .IN0(reg_dest_new[3]), .IN1(\registers[17][3] ), .SEL(n5977), 
        .F(n3541) );
  MUX U6605 ( .IN0(reg_dest_new[2]), .IN1(\registers[17][2] ), .SEL(n5977), 
        .F(n3540) );
  IV U6606 ( .A(n5978), .Z(n5977) );
  MUX U6607 ( .IN0(\registers[17][1] ), .IN1(reg_dest_new[1]), .SEL(n5978), 
        .F(n3539) );
  MUX U6608 ( .IN0(\registers[17][0] ), .IN1(reg_dest_new[0]), .SEL(n5978), 
        .F(n3538) );
  NOR U6609 ( .A(n5966), .B(n5959), .Z(n5978) );
  MUX U6610 ( .IN0(reg_dest_new[31]), .IN1(\registers[16][31] ), .SEL(n5979), 
        .F(n3537) );
  MUX U6611 ( .IN0(reg_dest_new[30]), .IN1(\registers[16][30] ), .SEL(n5979), 
        .F(n3536) );
  MUX U6612 ( .IN0(reg_dest_new[29]), .IN1(\registers[16][29] ), .SEL(n5979), 
        .F(n3535) );
  MUX U6613 ( .IN0(reg_dest_new[28]), .IN1(\registers[16][28] ), .SEL(n5979), 
        .F(n3534) );
  MUX U6614 ( .IN0(reg_dest_new[27]), .IN1(\registers[16][27] ), .SEL(n5979), 
        .F(n3533) );
  MUX U6615 ( .IN0(reg_dest_new[26]), .IN1(\registers[16][26] ), .SEL(n5979), 
        .F(n3532) );
  MUX U6616 ( .IN0(reg_dest_new[25]), .IN1(\registers[16][25] ), .SEL(n5979), 
        .F(n3531) );
  MUX U6617 ( .IN0(reg_dest_new[24]), .IN1(\registers[16][24] ), .SEL(n5979), 
        .F(n3530) );
  MUX U6618 ( .IN0(reg_dest_new[23]), .IN1(\registers[16][23] ), .SEL(n5979), 
        .F(n3529) );
  MUX U6619 ( .IN0(reg_dest_new[22]), .IN1(\registers[16][22] ), .SEL(n5979), 
        .F(n3528) );
  MUX U6620 ( .IN0(reg_dest_new[21]), .IN1(\registers[16][21] ), .SEL(n5979), 
        .F(n3527) );
  MUX U6621 ( .IN0(reg_dest_new[20]), .IN1(\registers[16][20] ), .SEL(n5979), 
        .F(n3526) );
  MUX U6622 ( .IN0(reg_dest_new[19]), .IN1(\registers[16][19] ), .SEL(n5979), 
        .F(n3525) );
  MUX U6623 ( .IN0(reg_dest_new[18]), .IN1(\registers[16][18] ), .SEL(n5979), 
        .F(n3524) );
  MUX U6624 ( .IN0(reg_dest_new[17]), .IN1(\registers[16][17] ), .SEL(n5979), 
        .F(n3523) );
  MUX U6625 ( .IN0(reg_dest_new[16]), .IN1(\registers[16][16] ), .SEL(n5979), 
        .F(n3522) );
  MUX U6626 ( .IN0(reg_dest_new[15]), .IN1(\registers[16][15] ), .SEL(n5979), 
        .F(n3521) );
  MUX U6627 ( .IN0(reg_dest_new[14]), .IN1(\registers[16][14] ), .SEL(n5979), 
        .F(n3520) );
  MUX U6628 ( .IN0(reg_dest_new[13]), .IN1(\registers[16][13] ), .SEL(n5979), 
        .F(n3519) );
  MUX U6629 ( .IN0(reg_dest_new[12]), .IN1(\registers[16][12] ), .SEL(n5979), 
        .F(n3518) );
  MUX U6630 ( .IN0(reg_dest_new[11]), .IN1(\registers[16][11] ), .SEL(n5979), 
        .F(n3517) );
  MUX U6631 ( .IN0(reg_dest_new[10]), .IN1(\registers[16][10] ), .SEL(n5979), 
        .F(n3516) );
  MUX U6632 ( .IN0(reg_dest_new[9]), .IN1(\registers[16][9] ), .SEL(n5979), 
        .F(n3515) );
  MUX U6633 ( .IN0(reg_dest_new[8]), .IN1(\registers[16][8] ), .SEL(n5979), 
        .F(n3514) );
  MUX U6634 ( .IN0(reg_dest_new[7]), .IN1(\registers[16][7] ), .SEL(n5979), 
        .F(n3513) );
  MUX U6635 ( .IN0(reg_dest_new[6]), .IN1(\registers[16][6] ), .SEL(n5979), 
        .F(n3512) );
  MUX U6636 ( .IN0(reg_dest_new[5]), .IN1(\registers[16][5] ), .SEL(n5979), 
        .F(n3511) );
  MUX U6637 ( .IN0(reg_dest_new[4]), .IN1(\registers[16][4] ), .SEL(n5979), 
        .F(n3510) );
  MUX U6638 ( .IN0(reg_dest_new[3]), .IN1(\registers[16][3] ), .SEL(n5979), 
        .F(n3509) );
  MUX U6639 ( .IN0(reg_dest_new[2]), .IN1(\registers[16][2] ), .SEL(n5979), 
        .F(n3508) );
  IV U6640 ( .A(n5980), .Z(n5979) );
  MUX U6641 ( .IN0(\registers[16][1] ), .IN1(reg_dest_new[1]), .SEL(n5980), 
        .F(n3507) );
  MUX U6642 ( .IN0(\registers[16][0] ), .IN1(reg_dest_new[0]), .SEL(n5980), 
        .F(n3506) );
  NOR U6643 ( .A(n5962), .B(n5966), .Z(n5980) );
  NANDN U6644 ( .A(rd_index[3]), .B(rd_index[4]), .Z(n5966) );
  MUX U6645 ( .IN0(reg_dest_new[31]), .IN1(\registers[15][31] ), .SEL(n5981), 
        .F(n3505) );
  MUX U6646 ( .IN0(reg_dest_new[30]), .IN1(\registers[15][30] ), .SEL(n5981), 
        .F(n3504) );
  MUX U6647 ( .IN0(reg_dest_new[29]), .IN1(\registers[15][29] ), .SEL(n5981), 
        .F(n3503) );
  MUX U6648 ( .IN0(reg_dest_new[28]), .IN1(\registers[15][28] ), .SEL(n5981), 
        .F(n3502) );
  MUX U6649 ( .IN0(reg_dest_new[27]), .IN1(\registers[15][27] ), .SEL(n5981), 
        .F(n3501) );
  MUX U6650 ( .IN0(reg_dest_new[26]), .IN1(\registers[15][26] ), .SEL(n5981), 
        .F(n3500) );
  MUX U6651 ( .IN0(reg_dest_new[25]), .IN1(\registers[15][25] ), .SEL(n5981), 
        .F(n3499) );
  MUX U6652 ( .IN0(reg_dest_new[24]), .IN1(\registers[15][24] ), .SEL(n5981), 
        .F(n3498) );
  MUX U6653 ( .IN0(reg_dest_new[23]), .IN1(\registers[15][23] ), .SEL(n5981), 
        .F(n3497) );
  MUX U6654 ( .IN0(reg_dest_new[22]), .IN1(\registers[15][22] ), .SEL(n5981), 
        .F(n3496) );
  MUX U6655 ( .IN0(reg_dest_new[21]), .IN1(\registers[15][21] ), .SEL(n5981), 
        .F(n3495) );
  MUX U6656 ( .IN0(reg_dest_new[20]), .IN1(\registers[15][20] ), .SEL(n5981), 
        .F(n3494) );
  MUX U6657 ( .IN0(reg_dest_new[19]), .IN1(\registers[15][19] ), .SEL(n5981), 
        .F(n3493) );
  MUX U6658 ( .IN0(reg_dest_new[18]), .IN1(\registers[15][18] ), .SEL(n5981), 
        .F(n3492) );
  MUX U6659 ( .IN0(reg_dest_new[17]), .IN1(\registers[15][17] ), .SEL(n5981), 
        .F(n3491) );
  MUX U6660 ( .IN0(reg_dest_new[16]), .IN1(\registers[15][16] ), .SEL(n5981), 
        .F(n3490) );
  MUX U6661 ( .IN0(reg_dest_new[15]), .IN1(\registers[15][15] ), .SEL(n5981), 
        .F(n3489) );
  MUX U6662 ( .IN0(reg_dest_new[14]), .IN1(\registers[15][14] ), .SEL(n5981), 
        .F(n3488) );
  MUX U6663 ( .IN0(reg_dest_new[13]), .IN1(\registers[15][13] ), .SEL(n5981), 
        .F(n3487) );
  MUX U6664 ( .IN0(reg_dest_new[12]), .IN1(\registers[15][12] ), .SEL(n5981), 
        .F(n3486) );
  MUX U6665 ( .IN0(reg_dest_new[11]), .IN1(\registers[15][11] ), .SEL(n5981), 
        .F(n3485) );
  MUX U6666 ( .IN0(reg_dest_new[10]), .IN1(\registers[15][10] ), .SEL(n5981), 
        .F(n3484) );
  MUX U6667 ( .IN0(reg_dest_new[9]), .IN1(\registers[15][9] ), .SEL(n5981), 
        .F(n3483) );
  MUX U6668 ( .IN0(reg_dest_new[8]), .IN1(\registers[15][8] ), .SEL(n5981), 
        .F(n3482) );
  MUX U6669 ( .IN0(reg_dest_new[7]), .IN1(\registers[15][7] ), .SEL(n5981), 
        .F(n3481) );
  MUX U6670 ( .IN0(reg_dest_new[6]), .IN1(\registers[15][6] ), .SEL(n5981), 
        .F(n3480) );
  MUX U6671 ( .IN0(reg_dest_new[5]), .IN1(\registers[15][5] ), .SEL(n5981), 
        .F(n3479) );
  MUX U6672 ( .IN0(reg_dest_new[4]), .IN1(\registers[15][4] ), .SEL(n5981), 
        .F(n3478) );
  MUX U6673 ( .IN0(reg_dest_new[3]), .IN1(\registers[15][3] ), .SEL(n5981), 
        .F(n3477) );
  MUX U6674 ( .IN0(reg_dest_new[2]), .IN1(\registers[15][2] ), .SEL(n5981), 
        .F(n3476) );
  IV U6675 ( .A(n5982), .Z(n5981) );
  MUX U6676 ( .IN0(\registers[15][1] ), .IN1(reg_dest_new[1]), .SEL(n5982), 
        .F(n3475) );
  MUX U6677 ( .IN0(\registers[15][0] ), .IN1(reg_dest_new[0]), .SEL(n5982), 
        .F(n3474) );
  NOR U6678 ( .A(n5983), .B(n5941), .Z(n5982) );
  MUX U6679 ( .IN0(reg_dest_new[31]), .IN1(\registers[14][31] ), .SEL(n5984), 
        .F(n3473) );
  MUX U6680 ( .IN0(reg_dest_new[30]), .IN1(\registers[14][30] ), .SEL(n5984), 
        .F(n3472) );
  MUX U6681 ( .IN0(reg_dest_new[29]), .IN1(\registers[14][29] ), .SEL(n5984), 
        .F(n3471) );
  MUX U6682 ( .IN0(reg_dest_new[28]), .IN1(\registers[14][28] ), .SEL(n5984), 
        .F(n3470) );
  MUX U6683 ( .IN0(reg_dest_new[27]), .IN1(\registers[14][27] ), .SEL(n5984), 
        .F(n3469) );
  MUX U6684 ( .IN0(reg_dest_new[26]), .IN1(\registers[14][26] ), .SEL(n5984), 
        .F(n3468) );
  MUX U6685 ( .IN0(reg_dest_new[25]), .IN1(\registers[14][25] ), .SEL(n5984), 
        .F(n3467) );
  MUX U6686 ( .IN0(reg_dest_new[24]), .IN1(\registers[14][24] ), .SEL(n5984), 
        .F(n3466) );
  MUX U6687 ( .IN0(reg_dest_new[23]), .IN1(\registers[14][23] ), .SEL(n5984), 
        .F(n3465) );
  MUX U6688 ( .IN0(reg_dest_new[22]), .IN1(\registers[14][22] ), .SEL(n5984), 
        .F(n3464) );
  MUX U6689 ( .IN0(reg_dest_new[21]), .IN1(\registers[14][21] ), .SEL(n5984), 
        .F(n3463) );
  MUX U6690 ( .IN0(reg_dest_new[20]), .IN1(\registers[14][20] ), .SEL(n5984), 
        .F(n3462) );
  MUX U6691 ( .IN0(reg_dest_new[19]), .IN1(\registers[14][19] ), .SEL(n5984), 
        .F(n3461) );
  MUX U6692 ( .IN0(reg_dest_new[18]), .IN1(\registers[14][18] ), .SEL(n5984), 
        .F(n3460) );
  MUX U6693 ( .IN0(reg_dest_new[17]), .IN1(\registers[14][17] ), .SEL(n5984), 
        .F(n3459) );
  MUX U6694 ( .IN0(reg_dest_new[16]), .IN1(\registers[14][16] ), .SEL(n5984), 
        .F(n3458) );
  MUX U6695 ( .IN0(reg_dest_new[15]), .IN1(\registers[14][15] ), .SEL(n5984), 
        .F(n3457) );
  MUX U6696 ( .IN0(reg_dest_new[14]), .IN1(\registers[14][14] ), .SEL(n5984), 
        .F(n3456) );
  MUX U6697 ( .IN0(reg_dest_new[13]), .IN1(\registers[14][13] ), .SEL(n5984), 
        .F(n3455) );
  MUX U6698 ( .IN0(reg_dest_new[12]), .IN1(\registers[14][12] ), .SEL(n5984), 
        .F(n3454) );
  MUX U6699 ( .IN0(reg_dest_new[11]), .IN1(\registers[14][11] ), .SEL(n5984), 
        .F(n3453) );
  MUX U6700 ( .IN0(reg_dest_new[10]), .IN1(\registers[14][10] ), .SEL(n5984), 
        .F(n3452) );
  MUX U6701 ( .IN0(reg_dest_new[9]), .IN1(\registers[14][9] ), .SEL(n5984), 
        .F(n3451) );
  MUX U6702 ( .IN0(reg_dest_new[8]), .IN1(\registers[14][8] ), .SEL(n5984), 
        .F(n3450) );
  MUX U6703 ( .IN0(reg_dest_new[7]), .IN1(\registers[14][7] ), .SEL(n5984), 
        .F(n3449) );
  MUX U6704 ( .IN0(reg_dest_new[6]), .IN1(\registers[14][6] ), .SEL(n5984), 
        .F(n3448) );
  MUX U6705 ( .IN0(reg_dest_new[5]), .IN1(\registers[14][5] ), .SEL(n5984), 
        .F(n3447) );
  MUX U6706 ( .IN0(reg_dest_new[4]), .IN1(\registers[14][4] ), .SEL(n5984), 
        .F(n3446) );
  MUX U6707 ( .IN0(reg_dest_new[3]), .IN1(\registers[14][3] ), .SEL(n5984), 
        .F(n3445) );
  MUX U6708 ( .IN0(reg_dest_new[2]), .IN1(\registers[14][2] ), .SEL(n5984), 
        .F(n3444) );
  IV U6709 ( .A(n5985), .Z(n5984) );
  MUX U6710 ( .IN0(\registers[14][1] ), .IN1(reg_dest_new[1]), .SEL(n5985), 
        .F(n3443) );
  MUX U6711 ( .IN0(\registers[14][0] ), .IN1(reg_dest_new[0]), .SEL(n5985), 
        .F(n3442) );
  NOR U6712 ( .A(n5983), .B(n5944), .Z(n5985) );
  MUX U6713 ( .IN0(reg_dest_new[31]), .IN1(\registers[13][31] ), .SEL(n5986), 
        .F(n3441) );
  MUX U6714 ( .IN0(reg_dest_new[30]), .IN1(\registers[13][30] ), .SEL(n5986), 
        .F(n3440) );
  MUX U6715 ( .IN0(reg_dest_new[29]), .IN1(\registers[13][29] ), .SEL(n5986), 
        .F(n3439) );
  MUX U6716 ( .IN0(reg_dest_new[28]), .IN1(\registers[13][28] ), .SEL(n5986), 
        .F(n3438) );
  MUX U6717 ( .IN0(reg_dest_new[27]), .IN1(\registers[13][27] ), .SEL(n5986), 
        .F(n3437) );
  MUX U6718 ( .IN0(reg_dest_new[26]), .IN1(\registers[13][26] ), .SEL(n5986), 
        .F(n3436) );
  MUX U6719 ( .IN0(reg_dest_new[25]), .IN1(\registers[13][25] ), .SEL(n5986), 
        .F(n3435) );
  MUX U6720 ( .IN0(reg_dest_new[24]), .IN1(\registers[13][24] ), .SEL(n5986), 
        .F(n3434) );
  MUX U6721 ( .IN0(reg_dest_new[23]), .IN1(\registers[13][23] ), .SEL(n5986), 
        .F(n3433) );
  MUX U6722 ( .IN0(reg_dest_new[22]), .IN1(\registers[13][22] ), .SEL(n5986), 
        .F(n3432) );
  MUX U6723 ( .IN0(reg_dest_new[21]), .IN1(\registers[13][21] ), .SEL(n5986), 
        .F(n3431) );
  MUX U6724 ( .IN0(reg_dest_new[20]), .IN1(\registers[13][20] ), .SEL(n5986), 
        .F(n3430) );
  MUX U6725 ( .IN0(reg_dest_new[19]), .IN1(\registers[13][19] ), .SEL(n5986), 
        .F(n3429) );
  MUX U6726 ( .IN0(reg_dest_new[18]), .IN1(\registers[13][18] ), .SEL(n5986), 
        .F(n3428) );
  MUX U6727 ( .IN0(reg_dest_new[17]), .IN1(\registers[13][17] ), .SEL(n5986), 
        .F(n3427) );
  MUX U6728 ( .IN0(reg_dest_new[16]), .IN1(\registers[13][16] ), .SEL(n5986), 
        .F(n3426) );
  MUX U6729 ( .IN0(reg_dest_new[15]), .IN1(\registers[13][15] ), .SEL(n5986), 
        .F(n3425) );
  MUX U6730 ( .IN0(reg_dest_new[14]), .IN1(\registers[13][14] ), .SEL(n5986), 
        .F(n3424) );
  MUX U6731 ( .IN0(reg_dest_new[13]), .IN1(\registers[13][13] ), .SEL(n5986), 
        .F(n3423) );
  MUX U6732 ( .IN0(reg_dest_new[12]), .IN1(\registers[13][12] ), .SEL(n5986), 
        .F(n3422) );
  MUX U6733 ( .IN0(reg_dest_new[11]), .IN1(\registers[13][11] ), .SEL(n5986), 
        .F(n3421) );
  MUX U6734 ( .IN0(reg_dest_new[10]), .IN1(\registers[13][10] ), .SEL(n5986), 
        .F(n3420) );
  MUX U6735 ( .IN0(reg_dest_new[9]), .IN1(\registers[13][9] ), .SEL(n5986), 
        .F(n3419) );
  MUX U6736 ( .IN0(reg_dest_new[8]), .IN1(\registers[13][8] ), .SEL(n5986), 
        .F(n3418) );
  MUX U6737 ( .IN0(reg_dest_new[7]), .IN1(\registers[13][7] ), .SEL(n5986), 
        .F(n3417) );
  MUX U6738 ( .IN0(reg_dest_new[6]), .IN1(\registers[13][6] ), .SEL(n5986), 
        .F(n3416) );
  MUX U6739 ( .IN0(reg_dest_new[5]), .IN1(\registers[13][5] ), .SEL(n5986), 
        .F(n3415) );
  MUX U6740 ( .IN0(reg_dest_new[4]), .IN1(\registers[13][4] ), .SEL(n5986), 
        .F(n3414) );
  MUX U6741 ( .IN0(reg_dest_new[3]), .IN1(\registers[13][3] ), .SEL(n5986), 
        .F(n3413) );
  MUX U6742 ( .IN0(reg_dest_new[2]), .IN1(\registers[13][2] ), .SEL(n5986), 
        .F(n3412) );
  IV U6743 ( .A(n5987), .Z(n5986) );
  MUX U6744 ( .IN0(\registers[13][1] ), .IN1(reg_dest_new[1]), .SEL(n5987), 
        .F(n3411) );
  MUX U6745 ( .IN0(\registers[13][0] ), .IN1(reg_dest_new[0]), .SEL(n5987), 
        .F(n3410) );
  NOR U6746 ( .A(n5983), .B(n5947), .Z(n5987) );
  MUX U6747 ( .IN0(reg_dest_new[31]), .IN1(\registers[12][31] ), .SEL(n5988), 
        .F(n3409) );
  MUX U6748 ( .IN0(reg_dest_new[30]), .IN1(\registers[12][30] ), .SEL(n5988), 
        .F(n3408) );
  MUX U6749 ( .IN0(reg_dest_new[29]), .IN1(\registers[12][29] ), .SEL(n5988), 
        .F(n3407) );
  MUX U6750 ( .IN0(reg_dest_new[28]), .IN1(\registers[12][28] ), .SEL(n5988), 
        .F(n3406) );
  MUX U6751 ( .IN0(reg_dest_new[27]), .IN1(\registers[12][27] ), .SEL(n5988), 
        .F(n3405) );
  MUX U6752 ( .IN0(reg_dest_new[26]), .IN1(\registers[12][26] ), .SEL(n5988), 
        .F(n3404) );
  MUX U6753 ( .IN0(reg_dest_new[25]), .IN1(\registers[12][25] ), .SEL(n5988), 
        .F(n3403) );
  MUX U6754 ( .IN0(reg_dest_new[24]), .IN1(\registers[12][24] ), .SEL(n5988), 
        .F(n3402) );
  MUX U6755 ( .IN0(reg_dest_new[23]), .IN1(\registers[12][23] ), .SEL(n5988), 
        .F(n3401) );
  MUX U6756 ( .IN0(reg_dest_new[22]), .IN1(\registers[12][22] ), .SEL(n5988), 
        .F(n3400) );
  MUX U6757 ( .IN0(reg_dest_new[21]), .IN1(\registers[12][21] ), .SEL(n5988), 
        .F(n3399) );
  MUX U6758 ( .IN0(reg_dest_new[20]), .IN1(\registers[12][20] ), .SEL(n5988), 
        .F(n3398) );
  MUX U6759 ( .IN0(reg_dest_new[19]), .IN1(\registers[12][19] ), .SEL(n5988), 
        .F(n3397) );
  MUX U6760 ( .IN0(reg_dest_new[18]), .IN1(\registers[12][18] ), .SEL(n5988), 
        .F(n3396) );
  MUX U6761 ( .IN0(reg_dest_new[17]), .IN1(\registers[12][17] ), .SEL(n5988), 
        .F(n3395) );
  MUX U6762 ( .IN0(reg_dest_new[16]), .IN1(\registers[12][16] ), .SEL(n5988), 
        .F(n3394) );
  MUX U6763 ( .IN0(reg_dest_new[15]), .IN1(\registers[12][15] ), .SEL(n5988), 
        .F(n3393) );
  MUX U6764 ( .IN0(reg_dest_new[14]), .IN1(\registers[12][14] ), .SEL(n5988), 
        .F(n3392) );
  MUX U6765 ( .IN0(reg_dest_new[13]), .IN1(\registers[12][13] ), .SEL(n5988), 
        .F(n3391) );
  MUX U6766 ( .IN0(reg_dest_new[12]), .IN1(\registers[12][12] ), .SEL(n5988), 
        .F(n3390) );
  MUX U6767 ( .IN0(reg_dest_new[11]), .IN1(\registers[12][11] ), .SEL(n5988), 
        .F(n3389) );
  MUX U6768 ( .IN0(reg_dest_new[10]), .IN1(\registers[12][10] ), .SEL(n5988), 
        .F(n3388) );
  MUX U6769 ( .IN0(reg_dest_new[9]), .IN1(\registers[12][9] ), .SEL(n5988), 
        .F(n3387) );
  MUX U6770 ( .IN0(reg_dest_new[8]), .IN1(\registers[12][8] ), .SEL(n5988), 
        .F(n3386) );
  MUX U6771 ( .IN0(reg_dest_new[7]), .IN1(\registers[12][7] ), .SEL(n5988), 
        .F(n3385) );
  MUX U6772 ( .IN0(reg_dest_new[6]), .IN1(\registers[12][6] ), .SEL(n5988), 
        .F(n3384) );
  MUX U6773 ( .IN0(reg_dest_new[5]), .IN1(\registers[12][5] ), .SEL(n5988), 
        .F(n3383) );
  MUX U6774 ( .IN0(reg_dest_new[4]), .IN1(\registers[12][4] ), .SEL(n5988), 
        .F(n3382) );
  MUX U6775 ( .IN0(reg_dest_new[3]), .IN1(\registers[12][3] ), .SEL(n5988), 
        .F(n3381) );
  MUX U6776 ( .IN0(reg_dest_new[2]), .IN1(\registers[12][2] ), .SEL(n5988), 
        .F(n3380) );
  IV U6777 ( .A(n5989), .Z(n5988) );
  MUX U6778 ( .IN0(\registers[12][1] ), .IN1(reg_dest_new[1]), .SEL(n5989), 
        .F(n3379) );
  MUX U6779 ( .IN0(\registers[12][0] ), .IN1(reg_dest_new[0]), .SEL(n5989), 
        .F(n3378) );
  NOR U6780 ( .A(n5983), .B(n5950), .Z(n5989) );
  MUX U6781 ( .IN0(reg_dest_new[31]), .IN1(\registers[11][31] ), .SEL(n5990), 
        .F(n3377) );
  MUX U6782 ( .IN0(reg_dest_new[30]), .IN1(\registers[11][30] ), .SEL(n5990), 
        .F(n3376) );
  MUX U6783 ( .IN0(reg_dest_new[29]), .IN1(\registers[11][29] ), .SEL(n5990), 
        .F(n3375) );
  MUX U6784 ( .IN0(reg_dest_new[28]), .IN1(\registers[11][28] ), .SEL(n5990), 
        .F(n3374) );
  MUX U6785 ( .IN0(reg_dest_new[27]), .IN1(\registers[11][27] ), .SEL(n5990), 
        .F(n3373) );
  MUX U6786 ( .IN0(reg_dest_new[26]), .IN1(\registers[11][26] ), .SEL(n5990), 
        .F(n3372) );
  MUX U6787 ( .IN0(reg_dest_new[25]), .IN1(\registers[11][25] ), .SEL(n5990), 
        .F(n3371) );
  MUX U6788 ( .IN0(reg_dest_new[24]), .IN1(\registers[11][24] ), .SEL(n5990), 
        .F(n3370) );
  MUX U6789 ( .IN0(reg_dest_new[23]), .IN1(\registers[11][23] ), .SEL(n5990), 
        .F(n3369) );
  MUX U6790 ( .IN0(reg_dest_new[22]), .IN1(\registers[11][22] ), .SEL(n5990), 
        .F(n3368) );
  MUX U6791 ( .IN0(reg_dest_new[21]), .IN1(\registers[11][21] ), .SEL(n5990), 
        .F(n3367) );
  MUX U6792 ( .IN0(reg_dest_new[20]), .IN1(\registers[11][20] ), .SEL(n5990), 
        .F(n3366) );
  MUX U6793 ( .IN0(reg_dest_new[19]), .IN1(\registers[11][19] ), .SEL(n5990), 
        .F(n3365) );
  MUX U6794 ( .IN0(reg_dest_new[18]), .IN1(\registers[11][18] ), .SEL(n5990), 
        .F(n3364) );
  MUX U6795 ( .IN0(reg_dest_new[17]), .IN1(\registers[11][17] ), .SEL(n5990), 
        .F(n3363) );
  MUX U6796 ( .IN0(reg_dest_new[16]), .IN1(\registers[11][16] ), .SEL(n5990), 
        .F(n3362) );
  MUX U6797 ( .IN0(reg_dest_new[15]), .IN1(\registers[11][15] ), .SEL(n5990), 
        .F(n3361) );
  MUX U6798 ( .IN0(reg_dest_new[14]), .IN1(\registers[11][14] ), .SEL(n5990), 
        .F(n3360) );
  MUX U6799 ( .IN0(reg_dest_new[13]), .IN1(\registers[11][13] ), .SEL(n5990), 
        .F(n3359) );
  MUX U6800 ( .IN0(reg_dest_new[12]), .IN1(\registers[11][12] ), .SEL(n5990), 
        .F(n3358) );
  MUX U6801 ( .IN0(reg_dest_new[11]), .IN1(\registers[11][11] ), .SEL(n5990), 
        .F(n3357) );
  MUX U6802 ( .IN0(reg_dest_new[10]), .IN1(\registers[11][10] ), .SEL(n5990), 
        .F(n3356) );
  MUX U6803 ( .IN0(reg_dest_new[9]), .IN1(\registers[11][9] ), .SEL(n5990), 
        .F(n3355) );
  MUX U6804 ( .IN0(reg_dest_new[8]), .IN1(\registers[11][8] ), .SEL(n5990), 
        .F(n3354) );
  MUX U6805 ( .IN0(reg_dest_new[7]), .IN1(\registers[11][7] ), .SEL(n5990), 
        .F(n3353) );
  MUX U6806 ( .IN0(reg_dest_new[6]), .IN1(\registers[11][6] ), .SEL(n5990), 
        .F(n3352) );
  MUX U6807 ( .IN0(reg_dest_new[5]), .IN1(\registers[11][5] ), .SEL(n5990), 
        .F(n3351) );
  MUX U6808 ( .IN0(reg_dest_new[4]), .IN1(\registers[11][4] ), .SEL(n5990), 
        .F(n3350) );
  MUX U6809 ( .IN0(reg_dest_new[3]), .IN1(\registers[11][3] ), .SEL(n5990), 
        .F(n3349) );
  MUX U6810 ( .IN0(reg_dest_new[2]), .IN1(\registers[11][2] ), .SEL(n5990), 
        .F(n3348) );
  IV U6811 ( .A(n5991), .Z(n5990) );
  MUX U6812 ( .IN0(\registers[11][1] ), .IN1(reg_dest_new[1]), .SEL(n5991), 
        .F(n3347) );
  MUX U6813 ( .IN0(\registers[11][0] ), .IN1(reg_dest_new[0]), .SEL(n5991), 
        .F(n3346) );
  NOR U6814 ( .A(n5983), .B(n5953), .Z(n5991) );
  MUX U6815 ( .IN0(reg_dest_new[31]), .IN1(\registers[10][31] ), .SEL(n5992), 
        .F(n3345) );
  MUX U6816 ( .IN0(reg_dest_new[30]), .IN1(\registers[10][30] ), .SEL(n5992), 
        .F(n3344) );
  MUX U6817 ( .IN0(reg_dest_new[29]), .IN1(\registers[10][29] ), .SEL(n5992), 
        .F(n3343) );
  MUX U6818 ( .IN0(reg_dest_new[28]), .IN1(\registers[10][28] ), .SEL(n5992), 
        .F(n3342) );
  MUX U6819 ( .IN0(reg_dest_new[27]), .IN1(\registers[10][27] ), .SEL(n5992), 
        .F(n3341) );
  MUX U6820 ( .IN0(reg_dest_new[26]), .IN1(\registers[10][26] ), .SEL(n5992), 
        .F(n3340) );
  MUX U6821 ( .IN0(reg_dest_new[25]), .IN1(\registers[10][25] ), .SEL(n5992), 
        .F(n3339) );
  MUX U6822 ( .IN0(reg_dest_new[24]), .IN1(\registers[10][24] ), .SEL(n5992), 
        .F(n3338) );
  MUX U6823 ( .IN0(reg_dest_new[23]), .IN1(\registers[10][23] ), .SEL(n5992), 
        .F(n3337) );
  MUX U6824 ( .IN0(reg_dest_new[22]), .IN1(\registers[10][22] ), .SEL(n5992), 
        .F(n3336) );
  MUX U6825 ( .IN0(reg_dest_new[21]), .IN1(\registers[10][21] ), .SEL(n5992), 
        .F(n3335) );
  MUX U6826 ( .IN0(reg_dest_new[20]), .IN1(\registers[10][20] ), .SEL(n5992), 
        .F(n3334) );
  MUX U6827 ( .IN0(reg_dest_new[19]), .IN1(\registers[10][19] ), .SEL(n5992), 
        .F(n3333) );
  MUX U6828 ( .IN0(reg_dest_new[18]), .IN1(\registers[10][18] ), .SEL(n5992), 
        .F(n3332) );
  MUX U6829 ( .IN0(reg_dest_new[17]), .IN1(\registers[10][17] ), .SEL(n5992), 
        .F(n3331) );
  MUX U6830 ( .IN0(reg_dest_new[16]), .IN1(\registers[10][16] ), .SEL(n5992), 
        .F(n3330) );
  MUX U6831 ( .IN0(reg_dest_new[15]), .IN1(\registers[10][15] ), .SEL(n5992), 
        .F(n3329) );
  MUX U6832 ( .IN0(reg_dest_new[14]), .IN1(\registers[10][14] ), .SEL(n5992), 
        .F(n3328) );
  MUX U6833 ( .IN0(reg_dest_new[13]), .IN1(\registers[10][13] ), .SEL(n5992), 
        .F(n3327) );
  MUX U6834 ( .IN0(reg_dest_new[12]), .IN1(\registers[10][12] ), .SEL(n5992), 
        .F(n3326) );
  MUX U6835 ( .IN0(reg_dest_new[11]), .IN1(\registers[10][11] ), .SEL(n5992), 
        .F(n3325) );
  MUX U6836 ( .IN0(reg_dest_new[10]), .IN1(\registers[10][10] ), .SEL(n5992), 
        .F(n3324) );
  MUX U6837 ( .IN0(reg_dest_new[9]), .IN1(\registers[10][9] ), .SEL(n5992), 
        .F(n3323) );
  MUX U6838 ( .IN0(reg_dest_new[8]), .IN1(\registers[10][8] ), .SEL(n5992), 
        .F(n3322) );
  MUX U6839 ( .IN0(reg_dest_new[7]), .IN1(\registers[10][7] ), .SEL(n5992), 
        .F(n3321) );
  MUX U6840 ( .IN0(reg_dest_new[6]), .IN1(\registers[10][6] ), .SEL(n5992), 
        .F(n3320) );
  MUX U6841 ( .IN0(reg_dest_new[5]), .IN1(\registers[10][5] ), .SEL(n5992), 
        .F(n3319) );
  MUX U6842 ( .IN0(reg_dest_new[4]), .IN1(\registers[10][4] ), .SEL(n5992), 
        .F(n3318) );
  MUX U6843 ( .IN0(reg_dest_new[3]), .IN1(\registers[10][3] ), .SEL(n5992), 
        .F(n3317) );
  MUX U6844 ( .IN0(reg_dest_new[2]), .IN1(\registers[10][2] ), .SEL(n5992), 
        .F(n3316) );
  IV U6845 ( .A(n5993), .Z(n5992) );
  MUX U6846 ( .IN0(\registers[10][1] ), .IN1(reg_dest_new[1]), .SEL(n5993), 
        .F(n3315) );
  MUX U6847 ( .IN0(\registers[10][0] ), .IN1(reg_dest_new[0]), .SEL(n5993), 
        .F(n3314) );
  NOR U6848 ( .A(n5983), .B(n5956), .Z(n5993) );
  MUX U6849 ( .IN0(reg_dest_new[31]), .IN1(\registers[9][31] ), .SEL(n5994), 
        .F(n3313) );
  MUX U6850 ( .IN0(reg_dest_new[30]), .IN1(\registers[9][30] ), .SEL(n5994), 
        .F(n3312) );
  MUX U6851 ( .IN0(reg_dest_new[29]), .IN1(\registers[9][29] ), .SEL(n5994), 
        .F(n3311) );
  MUX U6852 ( .IN0(reg_dest_new[28]), .IN1(\registers[9][28] ), .SEL(n5994), 
        .F(n3310) );
  MUX U6853 ( .IN0(reg_dest_new[27]), .IN1(\registers[9][27] ), .SEL(n5994), 
        .F(n3309) );
  MUX U6854 ( .IN0(reg_dest_new[26]), .IN1(\registers[9][26] ), .SEL(n5994), 
        .F(n3308) );
  MUX U6855 ( .IN0(reg_dest_new[25]), .IN1(\registers[9][25] ), .SEL(n5994), 
        .F(n3307) );
  MUX U6856 ( .IN0(reg_dest_new[24]), .IN1(\registers[9][24] ), .SEL(n5994), 
        .F(n3306) );
  MUX U6857 ( .IN0(reg_dest_new[23]), .IN1(\registers[9][23] ), .SEL(n5994), 
        .F(n3305) );
  MUX U6858 ( .IN0(reg_dest_new[22]), .IN1(\registers[9][22] ), .SEL(n5994), 
        .F(n3304) );
  MUX U6859 ( .IN0(reg_dest_new[21]), .IN1(\registers[9][21] ), .SEL(n5994), 
        .F(n3303) );
  MUX U6860 ( .IN0(reg_dest_new[20]), .IN1(\registers[9][20] ), .SEL(n5994), 
        .F(n3302) );
  MUX U6861 ( .IN0(reg_dest_new[19]), .IN1(\registers[9][19] ), .SEL(n5994), 
        .F(n3301) );
  MUX U6862 ( .IN0(reg_dest_new[18]), .IN1(\registers[9][18] ), .SEL(n5994), 
        .F(n3300) );
  MUX U6863 ( .IN0(reg_dest_new[17]), .IN1(\registers[9][17] ), .SEL(n5994), 
        .F(n3299) );
  MUX U6864 ( .IN0(reg_dest_new[16]), .IN1(\registers[9][16] ), .SEL(n5994), 
        .F(n3298) );
  MUX U6865 ( .IN0(reg_dest_new[15]), .IN1(\registers[9][15] ), .SEL(n5994), 
        .F(n3297) );
  MUX U6866 ( .IN0(reg_dest_new[14]), .IN1(\registers[9][14] ), .SEL(n5994), 
        .F(n3296) );
  MUX U6867 ( .IN0(reg_dest_new[13]), .IN1(\registers[9][13] ), .SEL(n5994), 
        .F(n3295) );
  MUX U6868 ( .IN0(reg_dest_new[12]), .IN1(\registers[9][12] ), .SEL(n5994), 
        .F(n3294) );
  MUX U6869 ( .IN0(reg_dest_new[11]), .IN1(\registers[9][11] ), .SEL(n5994), 
        .F(n3293) );
  MUX U6870 ( .IN0(reg_dest_new[10]), .IN1(\registers[9][10] ), .SEL(n5994), 
        .F(n3292) );
  MUX U6871 ( .IN0(reg_dest_new[9]), .IN1(\registers[9][9] ), .SEL(n5994), .F(
        n3291) );
  MUX U6872 ( .IN0(reg_dest_new[8]), .IN1(\registers[9][8] ), .SEL(n5994), .F(
        n3290) );
  MUX U6873 ( .IN0(reg_dest_new[7]), .IN1(\registers[9][7] ), .SEL(n5994), .F(
        n3289) );
  MUX U6874 ( .IN0(reg_dest_new[6]), .IN1(\registers[9][6] ), .SEL(n5994), .F(
        n3288) );
  MUX U6875 ( .IN0(reg_dest_new[5]), .IN1(\registers[9][5] ), .SEL(n5994), .F(
        n3287) );
  MUX U6876 ( .IN0(reg_dest_new[4]), .IN1(\registers[9][4] ), .SEL(n5994), .F(
        n3286) );
  MUX U6877 ( .IN0(reg_dest_new[3]), .IN1(\registers[9][3] ), .SEL(n5994), .F(
        n3285) );
  MUX U6878 ( .IN0(reg_dest_new[2]), .IN1(\registers[9][2] ), .SEL(n5994), .F(
        n3284) );
  IV U6879 ( .A(n5995), .Z(n5994) );
  MUX U6880 ( .IN0(\registers[9][1] ), .IN1(reg_dest_new[1]), .SEL(n5995), .F(
        n3283) );
  MUX U6881 ( .IN0(\registers[9][0] ), .IN1(reg_dest_new[0]), .SEL(n5995), .F(
        n3282) );
  NOR U6882 ( .A(n5983), .B(n5959), .Z(n5995) );
  MUX U6883 ( .IN0(reg_dest_new[31]), .IN1(\registers[8][31] ), .SEL(n5996), 
        .F(n3281) );
  MUX U6884 ( .IN0(reg_dest_new[30]), .IN1(\registers[8][30] ), .SEL(n5996), 
        .F(n3280) );
  MUX U6885 ( .IN0(reg_dest_new[29]), .IN1(\registers[8][29] ), .SEL(n5996), 
        .F(n3279) );
  MUX U6886 ( .IN0(reg_dest_new[28]), .IN1(\registers[8][28] ), .SEL(n5996), 
        .F(n3278) );
  MUX U6887 ( .IN0(reg_dest_new[27]), .IN1(\registers[8][27] ), .SEL(n5996), 
        .F(n3277) );
  MUX U6888 ( .IN0(reg_dest_new[26]), .IN1(\registers[8][26] ), .SEL(n5996), 
        .F(n3276) );
  MUX U6889 ( .IN0(reg_dest_new[25]), .IN1(\registers[8][25] ), .SEL(n5996), 
        .F(n3275) );
  MUX U6890 ( .IN0(reg_dest_new[24]), .IN1(\registers[8][24] ), .SEL(n5996), 
        .F(n3274) );
  MUX U6891 ( .IN0(reg_dest_new[23]), .IN1(\registers[8][23] ), .SEL(n5996), 
        .F(n3273) );
  MUX U6892 ( .IN0(reg_dest_new[22]), .IN1(\registers[8][22] ), .SEL(n5996), 
        .F(n3272) );
  MUX U6893 ( .IN0(reg_dest_new[21]), .IN1(\registers[8][21] ), .SEL(n5996), 
        .F(n3271) );
  MUX U6894 ( .IN0(reg_dest_new[20]), .IN1(\registers[8][20] ), .SEL(n5996), 
        .F(n3270) );
  MUX U6895 ( .IN0(reg_dest_new[19]), .IN1(\registers[8][19] ), .SEL(n5996), 
        .F(n3269) );
  MUX U6896 ( .IN0(reg_dest_new[18]), .IN1(\registers[8][18] ), .SEL(n5996), 
        .F(n3268) );
  MUX U6897 ( .IN0(reg_dest_new[17]), .IN1(\registers[8][17] ), .SEL(n5996), 
        .F(n3267) );
  MUX U6898 ( .IN0(reg_dest_new[16]), .IN1(\registers[8][16] ), .SEL(n5996), 
        .F(n3266) );
  MUX U6899 ( .IN0(reg_dest_new[15]), .IN1(\registers[8][15] ), .SEL(n5996), 
        .F(n3265) );
  MUX U6900 ( .IN0(reg_dest_new[14]), .IN1(\registers[8][14] ), .SEL(n5996), 
        .F(n3264) );
  MUX U6901 ( .IN0(reg_dest_new[13]), .IN1(\registers[8][13] ), .SEL(n5996), 
        .F(n3263) );
  MUX U6902 ( .IN0(reg_dest_new[12]), .IN1(\registers[8][12] ), .SEL(n5996), 
        .F(n3262) );
  MUX U6903 ( .IN0(reg_dest_new[11]), .IN1(\registers[8][11] ), .SEL(n5996), 
        .F(n3261) );
  MUX U6904 ( .IN0(reg_dest_new[10]), .IN1(\registers[8][10] ), .SEL(n5996), 
        .F(n3260) );
  MUX U6905 ( .IN0(reg_dest_new[9]), .IN1(\registers[8][9] ), .SEL(n5996), .F(
        n3259) );
  MUX U6906 ( .IN0(reg_dest_new[8]), .IN1(\registers[8][8] ), .SEL(n5996), .F(
        n3258) );
  MUX U6907 ( .IN0(reg_dest_new[7]), .IN1(\registers[8][7] ), .SEL(n5996), .F(
        n3257) );
  MUX U6908 ( .IN0(reg_dest_new[6]), .IN1(\registers[8][6] ), .SEL(n5996), .F(
        n3256) );
  MUX U6909 ( .IN0(reg_dest_new[5]), .IN1(\registers[8][5] ), .SEL(n5996), .F(
        n3255) );
  MUX U6910 ( .IN0(reg_dest_new[4]), .IN1(\registers[8][4] ), .SEL(n5996), .F(
        n3254) );
  MUX U6911 ( .IN0(reg_dest_new[3]), .IN1(\registers[8][3] ), .SEL(n5996), .F(
        n3253) );
  MUX U6912 ( .IN0(reg_dest_new[2]), .IN1(\registers[8][2] ), .SEL(n5996), .F(
        n3252) );
  IV U6913 ( .A(n5997), .Z(n5996) );
  MUX U6914 ( .IN0(\registers[8][1] ), .IN1(reg_dest_new[1]), .SEL(n5997), .F(
        n3251) );
  MUX U6915 ( .IN0(\registers[8][0] ), .IN1(reg_dest_new[0]), .SEL(n5997), .F(
        n3250) );
  NOR U6916 ( .A(n5983), .B(n5962), .Z(n5997) );
  OR U6917 ( .A(rd_index[2]), .B(n5998), .Z(n5962) );
  OR U6918 ( .A(rd_index[4]), .B(n5963), .Z(n5983) );
  IV U6919 ( .A(rd_index[3]), .Z(n5963) );
  MUX U6920 ( .IN0(reg_dest_new[31]), .IN1(\registers[7][31] ), .SEL(n5999), 
        .F(n3249) );
  MUX U6921 ( .IN0(reg_dest_new[30]), .IN1(\registers[7][30] ), .SEL(n5999), 
        .F(n3248) );
  MUX U6922 ( .IN0(reg_dest_new[29]), .IN1(\registers[7][29] ), .SEL(n5999), 
        .F(n3247) );
  MUX U6923 ( .IN0(reg_dest_new[28]), .IN1(\registers[7][28] ), .SEL(n5999), 
        .F(n3246) );
  MUX U6924 ( .IN0(reg_dest_new[27]), .IN1(\registers[7][27] ), .SEL(n5999), 
        .F(n3245) );
  MUX U6925 ( .IN0(reg_dest_new[26]), .IN1(\registers[7][26] ), .SEL(n5999), 
        .F(n3244) );
  MUX U6926 ( .IN0(reg_dest_new[25]), .IN1(\registers[7][25] ), .SEL(n5999), 
        .F(n3243) );
  MUX U6927 ( .IN0(reg_dest_new[24]), .IN1(\registers[7][24] ), .SEL(n5999), 
        .F(n3242) );
  MUX U6928 ( .IN0(reg_dest_new[23]), .IN1(\registers[7][23] ), .SEL(n5999), 
        .F(n3241) );
  MUX U6929 ( .IN0(reg_dest_new[22]), .IN1(\registers[7][22] ), .SEL(n5999), 
        .F(n3240) );
  MUX U6930 ( .IN0(reg_dest_new[21]), .IN1(\registers[7][21] ), .SEL(n5999), 
        .F(n3239) );
  MUX U6931 ( .IN0(reg_dest_new[20]), .IN1(\registers[7][20] ), .SEL(n5999), 
        .F(n3238) );
  MUX U6932 ( .IN0(reg_dest_new[19]), .IN1(\registers[7][19] ), .SEL(n5999), 
        .F(n3237) );
  MUX U6933 ( .IN0(reg_dest_new[18]), .IN1(\registers[7][18] ), .SEL(n5999), 
        .F(n3236) );
  MUX U6934 ( .IN0(reg_dest_new[17]), .IN1(\registers[7][17] ), .SEL(n5999), 
        .F(n3235) );
  MUX U6935 ( .IN0(reg_dest_new[16]), .IN1(\registers[7][16] ), .SEL(n5999), 
        .F(n3234) );
  MUX U6936 ( .IN0(reg_dest_new[15]), .IN1(\registers[7][15] ), .SEL(n5999), 
        .F(n3233) );
  MUX U6937 ( .IN0(reg_dest_new[14]), .IN1(\registers[7][14] ), .SEL(n5999), 
        .F(n3232) );
  MUX U6938 ( .IN0(reg_dest_new[13]), .IN1(\registers[7][13] ), .SEL(n5999), 
        .F(n3231) );
  MUX U6939 ( .IN0(reg_dest_new[12]), .IN1(\registers[7][12] ), .SEL(n5999), 
        .F(n3230) );
  MUX U6940 ( .IN0(reg_dest_new[11]), .IN1(\registers[7][11] ), .SEL(n5999), 
        .F(n3229) );
  MUX U6941 ( .IN0(reg_dest_new[10]), .IN1(\registers[7][10] ), .SEL(n5999), 
        .F(n3228) );
  MUX U6942 ( .IN0(reg_dest_new[9]), .IN1(\registers[7][9] ), .SEL(n5999), .F(
        n3227) );
  MUX U6943 ( .IN0(reg_dest_new[8]), .IN1(\registers[7][8] ), .SEL(n5999), .F(
        n3226) );
  MUX U6944 ( .IN0(reg_dest_new[7]), .IN1(\registers[7][7] ), .SEL(n5999), .F(
        n3225) );
  MUX U6945 ( .IN0(reg_dest_new[6]), .IN1(\registers[7][6] ), .SEL(n5999), .F(
        n3224) );
  MUX U6946 ( .IN0(reg_dest_new[5]), .IN1(\registers[7][5] ), .SEL(n5999), .F(
        n3223) );
  MUX U6947 ( .IN0(reg_dest_new[4]), .IN1(\registers[7][4] ), .SEL(n5999), .F(
        n3222) );
  MUX U6948 ( .IN0(reg_dest_new[3]), .IN1(\registers[7][3] ), .SEL(n5999), .F(
        n3221) );
  MUX U6949 ( .IN0(reg_dest_new[2]), .IN1(\registers[7][2] ), .SEL(n5999), .F(
        n3220) );
  IV U6950 ( .A(n6000), .Z(n5999) );
  MUX U6951 ( .IN0(\registers[7][1] ), .IN1(reg_dest_new[1]), .SEL(n6000), .F(
        n3219) );
  MUX U6952 ( .IN0(\registers[7][0] ), .IN1(reg_dest_new[0]), .SEL(n6000), .F(
        n3218) );
  NOR U6953 ( .A(n6001), .B(n5941), .Z(n6000) );
  NANDN U6954 ( .A(n6002), .B(rd_index[2]), .Z(n5941) );
  MUX U6955 ( .IN0(reg_dest_new[31]), .IN1(\registers[6][31] ), .SEL(n6003), 
        .F(n3217) );
  MUX U6956 ( .IN0(reg_dest_new[30]), .IN1(\registers[6][30] ), .SEL(n6003), 
        .F(n3216) );
  MUX U6957 ( .IN0(reg_dest_new[29]), .IN1(\registers[6][29] ), .SEL(n6003), 
        .F(n3215) );
  MUX U6958 ( .IN0(reg_dest_new[28]), .IN1(\registers[6][28] ), .SEL(n6003), 
        .F(n3214) );
  MUX U6959 ( .IN0(reg_dest_new[27]), .IN1(\registers[6][27] ), .SEL(n6003), 
        .F(n3213) );
  MUX U6960 ( .IN0(reg_dest_new[26]), .IN1(\registers[6][26] ), .SEL(n6003), 
        .F(n3212) );
  MUX U6961 ( .IN0(reg_dest_new[25]), .IN1(\registers[6][25] ), .SEL(n6003), 
        .F(n3211) );
  MUX U6962 ( .IN0(reg_dest_new[24]), .IN1(\registers[6][24] ), .SEL(n6003), 
        .F(n3210) );
  MUX U6963 ( .IN0(reg_dest_new[23]), .IN1(\registers[6][23] ), .SEL(n6003), 
        .F(n3209) );
  MUX U6964 ( .IN0(reg_dest_new[22]), .IN1(\registers[6][22] ), .SEL(n6003), 
        .F(n3208) );
  MUX U6965 ( .IN0(reg_dest_new[21]), .IN1(\registers[6][21] ), .SEL(n6003), 
        .F(n3207) );
  MUX U6966 ( .IN0(reg_dest_new[20]), .IN1(\registers[6][20] ), .SEL(n6003), 
        .F(n3206) );
  MUX U6967 ( .IN0(reg_dest_new[19]), .IN1(\registers[6][19] ), .SEL(n6003), 
        .F(n3205) );
  MUX U6968 ( .IN0(reg_dest_new[18]), .IN1(\registers[6][18] ), .SEL(n6003), 
        .F(n3204) );
  MUX U6969 ( .IN0(reg_dest_new[17]), .IN1(\registers[6][17] ), .SEL(n6003), 
        .F(n3203) );
  MUX U6970 ( .IN0(reg_dest_new[16]), .IN1(\registers[6][16] ), .SEL(n6003), 
        .F(n3202) );
  MUX U6971 ( .IN0(reg_dest_new[15]), .IN1(\registers[6][15] ), .SEL(n6003), 
        .F(n3201) );
  MUX U6972 ( .IN0(reg_dest_new[14]), .IN1(\registers[6][14] ), .SEL(n6003), 
        .F(n3200) );
  MUX U6973 ( .IN0(reg_dest_new[13]), .IN1(\registers[6][13] ), .SEL(n6003), 
        .F(n3199) );
  MUX U6974 ( .IN0(reg_dest_new[12]), .IN1(\registers[6][12] ), .SEL(n6003), 
        .F(n3198) );
  MUX U6975 ( .IN0(reg_dest_new[11]), .IN1(\registers[6][11] ), .SEL(n6003), 
        .F(n3197) );
  MUX U6976 ( .IN0(reg_dest_new[10]), .IN1(\registers[6][10] ), .SEL(n6003), 
        .F(n3196) );
  MUX U6977 ( .IN0(reg_dest_new[9]), .IN1(\registers[6][9] ), .SEL(n6003), .F(
        n3195) );
  MUX U6978 ( .IN0(reg_dest_new[8]), .IN1(\registers[6][8] ), .SEL(n6003), .F(
        n3194) );
  MUX U6979 ( .IN0(reg_dest_new[7]), .IN1(\registers[6][7] ), .SEL(n6003), .F(
        n3193) );
  MUX U6980 ( .IN0(reg_dest_new[6]), .IN1(\registers[6][6] ), .SEL(n6003), .F(
        n3192) );
  MUX U6981 ( .IN0(reg_dest_new[5]), .IN1(\registers[6][5] ), .SEL(n6003), .F(
        n3191) );
  MUX U6982 ( .IN0(reg_dest_new[4]), .IN1(\registers[6][4] ), .SEL(n6003), .F(
        n3190) );
  MUX U6983 ( .IN0(reg_dest_new[3]), .IN1(\registers[6][3] ), .SEL(n6003), .F(
        n3189) );
  MUX U6984 ( .IN0(reg_dest_new[2]), .IN1(\registers[6][2] ), .SEL(n6003), .F(
        n3188) );
  IV U6985 ( .A(n6004), .Z(n6003) );
  MUX U6986 ( .IN0(\registers[6][1] ), .IN1(reg_dest_new[1]), .SEL(n6004), .F(
        n3187) );
  MUX U6987 ( .IN0(\registers[6][0] ), .IN1(reg_dest_new[0]), .SEL(n6004), .F(
        n3186) );
  NOR U6988 ( .A(n6001), .B(n5944), .Z(n6004) );
  NANDN U6989 ( .A(n6005), .B(rd_index[2]), .Z(n5944) );
  MUX U6990 ( .IN0(reg_dest_new[31]), .IN1(\registers[5][31] ), .SEL(n6006), 
        .F(n3185) );
  MUX U6991 ( .IN0(reg_dest_new[30]), .IN1(\registers[5][30] ), .SEL(n6006), 
        .F(n3184) );
  MUX U6992 ( .IN0(reg_dest_new[29]), .IN1(\registers[5][29] ), .SEL(n6006), 
        .F(n3183) );
  MUX U6993 ( .IN0(reg_dest_new[28]), .IN1(\registers[5][28] ), .SEL(n6006), 
        .F(n3182) );
  MUX U6994 ( .IN0(reg_dest_new[27]), .IN1(\registers[5][27] ), .SEL(n6006), 
        .F(n3181) );
  MUX U6995 ( .IN0(reg_dest_new[26]), .IN1(\registers[5][26] ), .SEL(n6006), 
        .F(n3180) );
  MUX U6996 ( .IN0(reg_dest_new[25]), .IN1(\registers[5][25] ), .SEL(n6006), 
        .F(n3179) );
  MUX U6997 ( .IN0(reg_dest_new[24]), .IN1(\registers[5][24] ), .SEL(n6006), 
        .F(n3178) );
  MUX U6998 ( .IN0(reg_dest_new[23]), .IN1(\registers[5][23] ), .SEL(n6006), 
        .F(n3177) );
  MUX U6999 ( .IN0(reg_dest_new[22]), .IN1(\registers[5][22] ), .SEL(n6006), 
        .F(n3176) );
  MUX U7000 ( .IN0(reg_dest_new[21]), .IN1(\registers[5][21] ), .SEL(n6006), 
        .F(n3175) );
  MUX U7001 ( .IN0(reg_dest_new[20]), .IN1(\registers[5][20] ), .SEL(n6006), 
        .F(n3174) );
  MUX U7002 ( .IN0(reg_dest_new[19]), .IN1(\registers[5][19] ), .SEL(n6006), 
        .F(n3173) );
  MUX U7003 ( .IN0(reg_dest_new[18]), .IN1(\registers[5][18] ), .SEL(n6006), 
        .F(n3172) );
  MUX U7004 ( .IN0(reg_dest_new[17]), .IN1(\registers[5][17] ), .SEL(n6006), 
        .F(n3171) );
  MUX U7005 ( .IN0(reg_dest_new[16]), .IN1(\registers[5][16] ), .SEL(n6006), 
        .F(n3170) );
  MUX U7006 ( .IN0(reg_dest_new[15]), .IN1(\registers[5][15] ), .SEL(n6006), 
        .F(n3169) );
  MUX U7007 ( .IN0(reg_dest_new[14]), .IN1(\registers[5][14] ), .SEL(n6006), 
        .F(n3168) );
  MUX U7008 ( .IN0(reg_dest_new[13]), .IN1(\registers[5][13] ), .SEL(n6006), 
        .F(n3167) );
  MUX U7009 ( .IN0(reg_dest_new[12]), .IN1(\registers[5][12] ), .SEL(n6006), 
        .F(n3166) );
  MUX U7010 ( .IN0(reg_dest_new[11]), .IN1(\registers[5][11] ), .SEL(n6006), 
        .F(n3165) );
  MUX U7011 ( .IN0(reg_dest_new[10]), .IN1(\registers[5][10] ), .SEL(n6006), 
        .F(n3164) );
  MUX U7012 ( .IN0(reg_dest_new[9]), .IN1(\registers[5][9] ), .SEL(n6006), .F(
        n3163) );
  MUX U7013 ( .IN0(reg_dest_new[8]), .IN1(\registers[5][8] ), .SEL(n6006), .F(
        n3162) );
  MUX U7014 ( .IN0(reg_dest_new[7]), .IN1(\registers[5][7] ), .SEL(n6006), .F(
        n3161) );
  MUX U7015 ( .IN0(reg_dest_new[6]), .IN1(\registers[5][6] ), .SEL(n6006), .F(
        n3160) );
  MUX U7016 ( .IN0(reg_dest_new[5]), .IN1(\registers[5][5] ), .SEL(n6006), .F(
        n3159) );
  MUX U7017 ( .IN0(reg_dest_new[4]), .IN1(\registers[5][4] ), .SEL(n6006), .F(
        n3158) );
  MUX U7018 ( .IN0(reg_dest_new[3]), .IN1(\registers[5][3] ), .SEL(n6006), .F(
        n3157) );
  MUX U7019 ( .IN0(reg_dest_new[2]), .IN1(\registers[5][2] ), .SEL(n6006), .F(
        n3156) );
  IV U7020 ( .A(n6007), .Z(n6006) );
  MUX U7021 ( .IN0(\registers[5][1] ), .IN1(reg_dest_new[1]), .SEL(n6007), .F(
        n3155) );
  MUX U7022 ( .IN0(\registers[5][0] ), .IN1(reg_dest_new[0]), .SEL(n6007), .F(
        n3154) );
  NOR U7023 ( .A(n6001), .B(n5947), .Z(n6007) );
  NANDN U7024 ( .A(n6008), .B(rd_index[2]), .Z(n5947) );
  MUX U7025 ( .IN0(reg_dest_new[31]), .IN1(\registers[4][31] ), .SEL(n6009), 
        .F(n3153) );
  MUX U7026 ( .IN0(reg_dest_new[30]), .IN1(\registers[4][30] ), .SEL(n6009), 
        .F(n3152) );
  MUX U7027 ( .IN0(reg_dest_new[29]), .IN1(\registers[4][29] ), .SEL(n6009), 
        .F(n3151) );
  MUX U7028 ( .IN0(reg_dest_new[28]), .IN1(\registers[4][28] ), .SEL(n6009), 
        .F(n3150) );
  MUX U7029 ( .IN0(reg_dest_new[27]), .IN1(\registers[4][27] ), .SEL(n6009), 
        .F(n3149) );
  MUX U7030 ( .IN0(reg_dest_new[26]), .IN1(\registers[4][26] ), .SEL(n6009), 
        .F(n3148) );
  MUX U7031 ( .IN0(reg_dest_new[25]), .IN1(\registers[4][25] ), .SEL(n6009), 
        .F(n3147) );
  MUX U7032 ( .IN0(reg_dest_new[24]), .IN1(\registers[4][24] ), .SEL(n6009), 
        .F(n3146) );
  MUX U7033 ( .IN0(reg_dest_new[23]), .IN1(\registers[4][23] ), .SEL(n6009), 
        .F(n3145) );
  MUX U7034 ( .IN0(reg_dest_new[22]), .IN1(\registers[4][22] ), .SEL(n6009), 
        .F(n3144) );
  MUX U7035 ( .IN0(reg_dest_new[21]), .IN1(\registers[4][21] ), .SEL(n6009), 
        .F(n3143) );
  MUX U7036 ( .IN0(reg_dest_new[20]), .IN1(\registers[4][20] ), .SEL(n6009), 
        .F(n3142) );
  MUX U7037 ( .IN0(reg_dest_new[19]), .IN1(\registers[4][19] ), .SEL(n6009), 
        .F(n3141) );
  MUX U7038 ( .IN0(reg_dest_new[18]), .IN1(\registers[4][18] ), .SEL(n6009), 
        .F(n3140) );
  MUX U7039 ( .IN0(reg_dest_new[17]), .IN1(\registers[4][17] ), .SEL(n6009), 
        .F(n3139) );
  MUX U7040 ( .IN0(reg_dest_new[16]), .IN1(\registers[4][16] ), .SEL(n6009), 
        .F(n3138) );
  MUX U7041 ( .IN0(reg_dest_new[15]), .IN1(\registers[4][15] ), .SEL(n6009), 
        .F(n3137) );
  MUX U7042 ( .IN0(reg_dest_new[14]), .IN1(\registers[4][14] ), .SEL(n6009), 
        .F(n3136) );
  MUX U7043 ( .IN0(reg_dest_new[13]), .IN1(\registers[4][13] ), .SEL(n6009), 
        .F(n3135) );
  MUX U7044 ( .IN0(reg_dest_new[12]), .IN1(\registers[4][12] ), .SEL(n6009), 
        .F(n3134) );
  MUX U7045 ( .IN0(reg_dest_new[11]), .IN1(\registers[4][11] ), .SEL(n6009), 
        .F(n3133) );
  MUX U7046 ( .IN0(reg_dest_new[10]), .IN1(\registers[4][10] ), .SEL(n6009), 
        .F(n3132) );
  MUX U7047 ( .IN0(reg_dest_new[9]), .IN1(\registers[4][9] ), .SEL(n6009), .F(
        n3131) );
  MUX U7048 ( .IN0(reg_dest_new[8]), .IN1(\registers[4][8] ), .SEL(n6009), .F(
        n3130) );
  MUX U7049 ( .IN0(reg_dest_new[7]), .IN1(\registers[4][7] ), .SEL(n6009), .F(
        n3129) );
  MUX U7050 ( .IN0(reg_dest_new[6]), .IN1(\registers[4][6] ), .SEL(n6009), .F(
        n3128) );
  MUX U7051 ( .IN0(reg_dest_new[5]), .IN1(\registers[4][5] ), .SEL(n6009), .F(
        n3127) );
  MUX U7052 ( .IN0(reg_dest_new[4]), .IN1(\registers[4][4] ), .SEL(n6009), .F(
        n3126) );
  MUX U7053 ( .IN0(reg_dest_new[3]), .IN1(\registers[4][3] ), .SEL(n6009), .F(
        n3125) );
  MUX U7054 ( .IN0(reg_dest_new[2]), .IN1(\registers[4][2] ), .SEL(n6009), .F(
        n3124) );
  IV U7055 ( .A(n6010), .Z(n6009) );
  MUX U7056 ( .IN0(\registers[4][1] ), .IN1(reg_dest_new[1]), .SEL(n6010), .F(
        n3123) );
  MUX U7057 ( .IN0(\registers[4][0] ), .IN1(reg_dest_new[0]), .SEL(n6010), .F(
        n3122) );
  NOR U7058 ( .A(n6001), .B(n5950), .Z(n6010) );
  NANDN U7059 ( .A(n5998), .B(rd_index[2]), .Z(n5950) );
  OR U7060 ( .A(rd_index[1]), .B(rd_index[0]), .Z(n5998) );
  MUX U7061 ( .IN0(reg_dest_new[31]), .IN1(\registers[3][31] ), .SEL(n6011), 
        .F(n3121) );
  MUX U7062 ( .IN0(reg_dest_new[30]), .IN1(\registers[3][30] ), .SEL(n6011), 
        .F(n3120) );
  MUX U7063 ( .IN0(reg_dest_new[29]), .IN1(\registers[3][29] ), .SEL(n6011), 
        .F(n3119) );
  MUX U7064 ( .IN0(reg_dest_new[28]), .IN1(\registers[3][28] ), .SEL(n6011), 
        .F(n3118) );
  MUX U7065 ( .IN0(reg_dest_new[27]), .IN1(\registers[3][27] ), .SEL(n6011), 
        .F(n3117) );
  MUX U7066 ( .IN0(reg_dest_new[26]), .IN1(\registers[3][26] ), .SEL(n6011), 
        .F(n3116) );
  MUX U7067 ( .IN0(reg_dest_new[25]), .IN1(\registers[3][25] ), .SEL(n6011), 
        .F(n3115) );
  MUX U7068 ( .IN0(reg_dest_new[24]), .IN1(\registers[3][24] ), .SEL(n6011), 
        .F(n3114) );
  MUX U7069 ( .IN0(reg_dest_new[23]), .IN1(\registers[3][23] ), .SEL(n6011), 
        .F(n3113) );
  MUX U7070 ( .IN0(reg_dest_new[22]), .IN1(\registers[3][22] ), .SEL(n6011), 
        .F(n3112) );
  MUX U7071 ( .IN0(reg_dest_new[21]), .IN1(\registers[3][21] ), .SEL(n6011), 
        .F(n3111) );
  MUX U7072 ( .IN0(reg_dest_new[20]), .IN1(\registers[3][20] ), .SEL(n6011), 
        .F(n3110) );
  MUX U7073 ( .IN0(reg_dest_new[19]), .IN1(\registers[3][19] ), .SEL(n6011), 
        .F(n3109) );
  MUX U7074 ( .IN0(reg_dest_new[18]), .IN1(\registers[3][18] ), .SEL(n6011), 
        .F(n3108) );
  MUX U7075 ( .IN0(reg_dest_new[17]), .IN1(\registers[3][17] ), .SEL(n6011), 
        .F(n3107) );
  MUX U7076 ( .IN0(reg_dest_new[16]), .IN1(\registers[3][16] ), .SEL(n6011), 
        .F(n3106) );
  MUX U7077 ( .IN0(reg_dest_new[15]), .IN1(\registers[3][15] ), .SEL(n6011), 
        .F(n3105) );
  MUX U7078 ( .IN0(reg_dest_new[14]), .IN1(\registers[3][14] ), .SEL(n6011), 
        .F(n3104) );
  MUX U7079 ( .IN0(reg_dest_new[13]), .IN1(\registers[3][13] ), .SEL(n6011), 
        .F(n3103) );
  MUX U7080 ( .IN0(reg_dest_new[12]), .IN1(\registers[3][12] ), .SEL(n6011), 
        .F(n3102) );
  MUX U7081 ( .IN0(reg_dest_new[11]), .IN1(\registers[3][11] ), .SEL(n6011), 
        .F(n3101) );
  MUX U7082 ( .IN0(reg_dest_new[10]), .IN1(\registers[3][10] ), .SEL(n6011), 
        .F(n3100) );
  MUX U7083 ( .IN0(reg_dest_new[9]), .IN1(\registers[3][9] ), .SEL(n6011), .F(
        n3099) );
  MUX U7084 ( .IN0(reg_dest_new[8]), .IN1(\registers[3][8] ), .SEL(n6011), .F(
        n3098) );
  MUX U7085 ( .IN0(reg_dest_new[7]), .IN1(\registers[3][7] ), .SEL(n6011), .F(
        n3097) );
  MUX U7086 ( .IN0(reg_dest_new[6]), .IN1(\registers[3][6] ), .SEL(n6011), .F(
        n3096) );
  MUX U7087 ( .IN0(reg_dest_new[5]), .IN1(\registers[3][5] ), .SEL(n6011), .F(
        n3095) );
  MUX U7088 ( .IN0(reg_dest_new[4]), .IN1(\registers[3][4] ), .SEL(n6011), .F(
        n3094) );
  MUX U7089 ( .IN0(reg_dest_new[3]), .IN1(\registers[3][3] ), .SEL(n6011), .F(
        n3093) );
  MUX U7090 ( .IN0(reg_dest_new[2]), .IN1(\registers[3][2] ), .SEL(n6011), .F(
        n3092) );
  IV U7091 ( .A(n6012), .Z(n6011) );
  MUX U7092 ( .IN0(\registers[3][1] ), .IN1(reg_dest_new[1]), .SEL(n6012), .F(
        n3091) );
  MUX U7093 ( .IN0(\registers[3][0] ), .IN1(reg_dest_new[0]), .SEL(n6012), .F(
        n3090) );
  NOR U7094 ( .A(n6001), .B(n5953), .Z(n6012) );
  OR U7095 ( .A(rd_index[2]), .B(n6002), .Z(n5953) );
  NANDN U7096 ( .A(n6013), .B(rd_index[1]), .Z(n6002) );
  MUX U7097 ( .IN0(reg_dest_new[31]), .IN1(\registers[2][31] ), .SEL(n6014), 
        .F(n3089) );
  MUX U7098 ( .IN0(reg_dest_new[30]), .IN1(\registers[2][30] ), .SEL(n6014), 
        .F(n3088) );
  MUX U7099 ( .IN0(reg_dest_new[29]), .IN1(\registers[2][29] ), .SEL(n6014), 
        .F(n3087) );
  MUX U7100 ( .IN0(reg_dest_new[28]), .IN1(\registers[2][28] ), .SEL(n6014), 
        .F(n3086) );
  MUX U7101 ( .IN0(reg_dest_new[27]), .IN1(\registers[2][27] ), .SEL(n6014), 
        .F(n3085) );
  MUX U7102 ( .IN0(reg_dest_new[26]), .IN1(\registers[2][26] ), .SEL(n6014), 
        .F(n3084) );
  MUX U7103 ( .IN0(reg_dest_new[25]), .IN1(\registers[2][25] ), .SEL(n6014), 
        .F(n3083) );
  MUX U7104 ( .IN0(reg_dest_new[24]), .IN1(\registers[2][24] ), .SEL(n6014), 
        .F(n3082) );
  MUX U7105 ( .IN0(reg_dest_new[23]), .IN1(\registers[2][23] ), .SEL(n6014), 
        .F(n3081) );
  MUX U7106 ( .IN0(reg_dest_new[22]), .IN1(\registers[2][22] ), .SEL(n6014), 
        .F(n3080) );
  MUX U7107 ( .IN0(reg_dest_new[21]), .IN1(\registers[2][21] ), .SEL(n6014), 
        .F(n3079) );
  MUX U7108 ( .IN0(reg_dest_new[20]), .IN1(\registers[2][20] ), .SEL(n6014), 
        .F(n3078) );
  MUX U7109 ( .IN0(reg_dest_new[19]), .IN1(\registers[2][19] ), .SEL(n6014), 
        .F(n3077) );
  MUX U7110 ( .IN0(reg_dest_new[18]), .IN1(\registers[2][18] ), .SEL(n6014), 
        .F(n3076) );
  MUX U7111 ( .IN0(reg_dest_new[17]), .IN1(\registers[2][17] ), .SEL(n6014), 
        .F(n3075) );
  MUX U7112 ( .IN0(reg_dest_new[16]), .IN1(\registers[2][16] ), .SEL(n6014), 
        .F(n3074) );
  MUX U7113 ( .IN0(reg_dest_new[15]), .IN1(\registers[2][15] ), .SEL(n6014), 
        .F(n3073) );
  MUX U7114 ( .IN0(reg_dest_new[14]), .IN1(\registers[2][14] ), .SEL(n6014), 
        .F(n3072) );
  MUX U7115 ( .IN0(reg_dest_new[13]), .IN1(\registers[2][13] ), .SEL(n6014), 
        .F(n3071) );
  MUX U7116 ( .IN0(reg_dest_new[12]), .IN1(\registers[2][12] ), .SEL(n6014), 
        .F(n3070) );
  MUX U7117 ( .IN0(reg_dest_new[11]), .IN1(\registers[2][11] ), .SEL(n6014), 
        .F(n3069) );
  MUX U7118 ( .IN0(reg_dest_new[10]), .IN1(\registers[2][10] ), .SEL(n6014), 
        .F(n3068) );
  MUX U7119 ( .IN0(reg_dest_new[9]), .IN1(\registers[2][9] ), .SEL(n6014), .F(
        n3067) );
  MUX U7120 ( .IN0(reg_dest_new[8]), .IN1(\registers[2][8] ), .SEL(n6014), .F(
        n3066) );
  MUX U7121 ( .IN0(reg_dest_new[7]), .IN1(\registers[2][7] ), .SEL(n6014), .F(
        n3065) );
  MUX U7122 ( .IN0(reg_dest_new[6]), .IN1(\registers[2][6] ), .SEL(n6014), .F(
        n3064) );
  MUX U7123 ( .IN0(reg_dest_new[5]), .IN1(\registers[2][5] ), .SEL(n6014), .F(
        n3063) );
  MUX U7124 ( .IN0(reg_dest_new[4]), .IN1(\registers[2][4] ), .SEL(n6014), .F(
        n3062) );
  MUX U7125 ( .IN0(reg_dest_new[3]), .IN1(\registers[2][3] ), .SEL(n6014), .F(
        n3061) );
  MUX U7126 ( .IN0(reg_dest_new[2]), .IN1(\registers[2][2] ), .SEL(n6014), .F(
        n3060) );
  IV U7127 ( .A(n6015), .Z(n6014) );
  MUX U7128 ( .IN0(\registers[2][1] ), .IN1(reg_dest_new[1]), .SEL(n6015), .F(
        n3059) );
  MUX U7129 ( .IN0(\registers[2][0] ), .IN1(reg_dest_new[0]), .SEL(n6015), .F(
        n3058) );
  NOR U7130 ( .A(n6001), .B(n5956), .Z(n6015) );
  OR U7131 ( .A(rd_index[2]), .B(n6005), .Z(n5956) );
  NANDN U7132 ( .A(rd_index[0]), .B(rd_index[1]), .Z(n6005) );
  MUX U7133 ( .IN0(reg_dest_new[31]), .IN1(\registers[1][31] ), .SEL(n6016), 
        .F(n3057) );
  MUX U7134 ( .IN0(reg_dest_new[30]), .IN1(\registers[1][30] ), .SEL(n6016), 
        .F(n3056) );
  MUX U7135 ( .IN0(reg_dest_new[29]), .IN1(\registers[1][29] ), .SEL(n6016), 
        .F(n3055) );
  MUX U7136 ( .IN0(reg_dest_new[28]), .IN1(\registers[1][28] ), .SEL(n6016), 
        .F(n3054) );
  MUX U7137 ( .IN0(reg_dest_new[27]), .IN1(\registers[1][27] ), .SEL(n6016), 
        .F(n3053) );
  MUX U7138 ( .IN0(reg_dest_new[26]), .IN1(\registers[1][26] ), .SEL(n6016), 
        .F(n3052) );
  MUX U7139 ( .IN0(reg_dest_new[25]), .IN1(\registers[1][25] ), .SEL(n6016), 
        .F(n3051) );
  MUX U7140 ( .IN0(reg_dest_new[24]), .IN1(\registers[1][24] ), .SEL(n6016), 
        .F(n3050) );
  MUX U7141 ( .IN0(reg_dest_new[23]), .IN1(\registers[1][23] ), .SEL(n6016), 
        .F(n3049) );
  MUX U7142 ( .IN0(reg_dest_new[22]), .IN1(\registers[1][22] ), .SEL(n6016), 
        .F(n3048) );
  MUX U7143 ( .IN0(reg_dest_new[21]), .IN1(\registers[1][21] ), .SEL(n6016), 
        .F(n3047) );
  MUX U7144 ( .IN0(reg_dest_new[20]), .IN1(\registers[1][20] ), .SEL(n6016), 
        .F(n3046) );
  MUX U7145 ( .IN0(reg_dest_new[19]), .IN1(\registers[1][19] ), .SEL(n6016), 
        .F(n3045) );
  MUX U7146 ( .IN0(reg_dest_new[18]), .IN1(\registers[1][18] ), .SEL(n6016), 
        .F(n3044) );
  MUX U7147 ( .IN0(reg_dest_new[17]), .IN1(\registers[1][17] ), .SEL(n6016), 
        .F(n3043) );
  MUX U7148 ( .IN0(reg_dest_new[16]), .IN1(\registers[1][16] ), .SEL(n6016), 
        .F(n3042) );
  MUX U7149 ( .IN0(reg_dest_new[15]), .IN1(\registers[1][15] ), .SEL(n6016), 
        .F(n3041) );
  MUX U7150 ( .IN0(reg_dest_new[14]), .IN1(\registers[1][14] ), .SEL(n6016), 
        .F(n3040) );
  MUX U7151 ( .IN0(reg_dest_new[13]), .IN1(\registers[1][13] ), .SEL(n6016), 
        .F(n3039) );
  MUX U7152 ( .IN0(reg_dest_new[12]), .IN1(\registers[1][12] ), .SEL(n6016), 
        .F(n3038) );
  MUX U7153 ( .IN0(reg_dest_new[11]), .IN1(\registers[1][11] ), .SEL(n6016), 
        .F(n3037) );
  MUX U7154 ( .IN0(reg_dest_new[10]), .IN1(\registers[1][10] ), .SEL(n6016), 
        .F(n3036) );
  MUX U7155 ( .IN0(reg_dest_new[9]), .IN1(\registers[1][9] ), .SEL(n6016), .F(
        n3035) );
  MUX U7156 ( .IN0(reg_dest_new[8]), .IN1(\registers[1][8] ), .SEL(n6016), .F(
        n3034) );
  MUX U7157 ( .IN0(reg_dest_new[7]), .IN1(\registers[1][7] ), .SEL(n6016), .F(
        n3033) );
  MUX U7158 ( .IN0(reg_dest_new[6]), .IN1(\registers[1][6] ), .SEL(n6016), .F(
        n3032) );
  MUX U7159 ( .IN0(reg_dest_new[5]), .IN1(\registers[1][5] ), .SEL(n6016), .F(
        n3031) );
  MUX U7160 ( .IN0(reg_dest_new[4]), .IN1(\registers[1][4] ), .SEL(n6016), .F(
        n3030) );
  MUX U7161 ( .IN0(reg_dest_new[3]), .IN1(\registers[1][3] ), .SEL(n6016), .F(
        n3029) );
  MUX U7162 ( .IN0(reg_dest_new[2]), .IN1(\registers[1][2] ), .SEL(n6016), .F(
        n3028) );
  IV U7163 ( .A(n6017), .Z(n6016) );
  MUX U7164 ( .IN0(\registers[1][1] ), .IN1(reg_dest_new[1]), .SEL(n6017), .F(
        n3027) );
  MUX U7165 ( .IN0(\registers[1][0] ), .IN1(reg_dest_new[0]), .SEL(n6017), .F(
        n3026) );
  NOR U7166 ( .A(n6001), .B(n5959), .Z(n6017) );
  OR U7167 ( .A(rd_index[2]), .B(n6008), .Z(n5959) );
  OR U7168 ( .A(rd_index[1]), .B(n6013), .Z(n6008) );
  IV U7169 ( .A(rd_index[0]), .Z(n6013) );
  OR U7170 ( .A(rd_index[4]), .B(rd_index[3]), .Z(n6001) );
endmodule

