
module sum_N16384_CC4 ( clk, rst, a, b, c );
  input [4095:0] a;
  input [4095:0] b;
  output [4095:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U5 ( .B(n4), .A(n5), .Z(n2) );
  XOR U6 ( .A(b[4095]), .B(n3), .Z(n4) );
  XNOR U7 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U8 ( .A(b[99]), .B(n7), .Z(c[99]) );
  XNOR U9 ( .A(b[999]), .B(n8), .Z(c[999]) );
  XNOR U10 ( .A(b[998]), .B(n9), .Z(c[998]) );
  XNOR U11 ( .A(b[997]), .B(n10), .Z(c[997]) );
  XNOR U12 ( .A(b[996]), .B(n11), .Z(c[996]) );
  XNOR U13 ( .A(b[995]), .B(n12), .Z(c[995]) );
  XNOR U14 ( .A(b[994]), .B(n13), .Z(c[994]) );
  XNOR U15 ( .A(b[993]), .B(n14), .Z(c[993]) );
  XNOR U16 ( .A(b[992]), .B(n15), .Z(c[992]) );
  XNOR U17 ( .A(b[991]), .B(n16), .Z(c[991]) );
  XNOR U18 ( .A(b[990]), .B(n17), .Z(c[990]) );
  XNOR U19 ( .A(b[98]), .B(n18), .Z(c[98]) );
  XNOR U20 ( .A(b[989]), .B(n19), .Z(c[989]) );
  XNOR U21 ( .A(b[988]), .B(n20), .Z(c[988]) );
  XNOR U22 ( .A(b[987]), .B(n21), .Z(c[987]) );
  XNOR U23 ( .A(b[986]), .B(n22), .Z(c[986]) );
  XNOR U24 ( .A(b[985]), .B(n23), .Z(c[985]) );
  XNOR U25 ( .A(b[984]), .B(n24), .Z(c[984]) );
  XNOR U26 ( .A(b[983]), .B(n25), .Z(c[983]) );
  XNOR U27 ( .A(b[982]), .B(n26), .Z(c[982]) );
  XNOR U28 ( .A(b[981]), .B(n27), .Z(c[981]) );
  XNOR U29 ( .A(b[980]), .B(n28), .Z(c[980]) );
  XNOR U30 ( .A(b[97]), .B(n29), .Z(c[97]) );
  XNOR U31 ( .A(b[979]), .B(n30), .Z(c[979]) );
  XNOR U32 ( .A(b[978]), .B(n31), .Z(c[978]) );
  XNOR U33 ( .A(b[977]), .B(n32), .Z(c[977]) );
  XNOR U34 ( .A(b[976]), .B(n33), .Z(c[976]) );
  XNOR U35 ( .A(b[975]), .B(n34), .Z(c[975]) );
  XNOR U36 ( .A(b[974]), .B(n35), .Z(c[974]) );
  XNOR U37 ( .A(b[973]), .B(n36), .Z(c[973]) );
  XNOR U38 ( .A(b[972]), .B(n37), .Z(c[972]) );
  XNOR U39 ( .A(b[971]), .B(n38), .Z(c[971]) );
  XNOR U40 ( .A(b[970]), .B(n39), .Z(c[970]) );
  XNOR U41 ( .A(b[96]), .B(n40), .Z(c[96]) );
  XNOR U42 ( .A(b[969]), .B(n41), .Z(c[969]) );
  XNOR U43 ( .A(b[968]), .B(n42), .Z(c[968]) );
  XNOR U44 ( .A(b[967]), .B(n43), .Z(c[967]) );
  XNOR U45 ( .A(b[966]), .B(n44), .Z(c[966]) );
  XNOR U46 ( .A(b[965]), .B(n45), .Z(c[965]) );
  XNOR U47 ( .A(b[964]), .B(n46), .Z(c[964]) );
  XNOR U48 ( .A(b[963]), .B(n47), .Z(c[963]) );
  XNOR U49 ( .A(b[962]), .B(n48), .Z(c[962]) );
  XNOR U50 ( .A(b[961]), .B(n49), .Z(c[961]) );
  XNOR U51 ( .A(b[960]), .B(n50), .Z(c[960]) );
  XNOR U52 ( .A(b[95]), .B(n51), .Z(c[95]) );
  XNOR U53 ( .A(b[959]), .B(n52), .Z(c[959]) );
  XNOR U54 ( .A(b[958]), .B(n53), .Z(c[958]) );
  XNOR U55 ( .A(b[957]), .B(n54), .Z(c[957]) );
  XNOR U56 ( .A(b[956]), .B(n55), .Z(c[956]) );
  XNOR U57 ( .A(b[955]), .B(n56), .Z(c[955]) );
  XNOR U58 ( .A(b[954]), .B(n57), .Z(c[954]) );
  XNOR U59 ( .A(b[953]), .B(n58), .Z(c[953]) );
  XNOR U60 ( .A(b[952]), .B(n59), .Z(c[952]) );
  XNOR U61 ( .A(b[951]), .B(n60), .Z(c[951]) );
  XNOR U62 ( .A(b[950]), .B(n61), .Z(c[950]) );
  XNOR U63 ( .A(b[94]), .B(n62), .Z(c[94]) );
  XNOR U64 ( .A(b[949]), .B(n63), .Z(c[949]) );
  XNOR U65 ( .A(b[948]), .B(n64), .Z(c[948]) );
  XNOR U66 ( .A(b[947]), .B(n65), .Z(c[947]) );
  XNOR U67 ( .A(b[946]), .B(n66), .Z(c[946]) );
  XNOR U68 ( .A(b[945]), .B(n67), .Z(c[945]) );
  XNOR U69 ( .A(b[944]), .B(n68), .Z(c[944]) );
  XNOR U70 ( .A(b[943]), .B(n69), .Z(c[943]) );
  XNOR U71 ( .A(b[942]), .B(n70), .Z(c[942]) );
  XNOR U72 ( .A(b[941]), .B(n71), .Z(c[941]) );
  XNOR U73 ( .A(b[940]), .B(n72), .Z(c[940]) );
  XNOR U74 ( .A(b[93]), .B(n73), .Z(c[93]) );
  XNOR U75 ( .A(b[939]), .B(n74), .Z(c[939]) );
  XNOR U76 ( .A(b[938]), .B(n75), .Z(c[938]) );
  XNOR U77 ( .A(b[937]), .B(n76), .Z(c[937]) );
  XNOR U78 ( .A(b[936]), .B(n77), .Z(c[936]) );
  XNOR U79 ( .A(b[935]), .B(n78), .Z(c[935]) );
  XNOR U80 ( .A(b[934]), .B(n79), .Z(c[934]) );
  XNOR U81 ( .A(b[933]), .B(n80), .Z(c[933]) );
  XNOR U82 ( .A(b[932]), .B(n81), .Z(c[932]) );
  XNOR U83 ( .A(b[931]), .B(n82), .Z(c[931]) );
  XNOR U84 ( .A(b[930]), .B(n83), .Z(c[930]) );
  XNOR U85 ( .A(b[92]), .B(n84), .Z(c[92]) );
  XNOR U86 ( .A(b[929]), .B(n85), .Z(c[929]) );
  XNOR U87 ( .A(b[928]), .B(n86), .Z(c[928]) );
  XNOR U88 ( .A(b[927]), .B(n87), .Z(c[927]) );
  XNOR U89 ( .A(b[926]), .B(n88), .Z(c[926]) );
  XNOR U90 ( .A(b[925]), .B(n89), .Z(c[925]) );
  XNOR U91 ( .A(b[924]), .B(n90), .Z(c[924]) );
  XNOR U92 ( .A(b[923]), .B(n91), .Z(c[923]) );
  XNOR U93 ( .A(b[922]), .B(n92), .Z(c[922]) );
  XNOR U94 ( .A(b[921]), .B(n93), .Z(c[921]) );
  XNOR U95 ( .A(b[920]), .B(n94), .Z(c[920]) );
  XNOR U96 ( .A(b[91]), .B(n95), .Z(c[91]) );
  XNOR U97 ( .A(b[919]), .B(n96), .Z(c[919]) );
  XNOR U98 ( .A(b[918]), .B(n97), .Z(c[918]) );
  XNOR U99 ( .A(b[917]), .B(n98), .Z(c[917]) );
  XNOR U100 ( .A(b[916]), .B(n99), .Z(c[916]) );
  XNOR U101 ( .A(b[915]), .B(n100), .Z(c[915]) );
  XNOR U102 ( .A(b[914]), .B(n101), .Z(c[914]) );
  XNOR U103 ( .A(b[913]), .B(n102), .Z(c[913]) );
  XNOR U104 ( .A(b[912]), .B(n103), .Z(c[912]) );
  XNOR U105 ( .A(b[911]), .B(n104), .Z(c[911]) );
  XNOR U106 ( .A(b[910]), .B(n105), .Z(c[910]) );
  XNOR U107 ( .A(b[90]), .B(n106), .Z(c[90]) );
  XNOR U108 ( .A(b[909]), .B(n107), .Z(c[909]) );
  XNOR U109 ( .A(b[908]), .B(n108), .Z(c[908]) );
  XNOR U110 ( .A(b[907]), .B(n109), .Z(c[907]) );
  XNOR U111 ( .A(b[906]), .B(n110), .Z(c[906]) );
  XNOR U112 ( .A(b[905]), .B(n111), .Z(c[905]) );
  XNOR U113 ( .A(b[904]), .B(n112), .Z(c[904]) );
  XNOR U114 ( .A(b[903]), .B(n113), .Z(c[903]) );
  XNOR U115 ( .A(b[902]), .B(n114), .Z(c[902]) );
  XNOR U116 ( .A(b[901]), .B(n115), .Z(c[901]) );
  XNOR U117 ( .A(b[900]), .B(n116), .Z(c[900]) );
  XNOR U118 ( .A(b[8]), .B(n117), .Z(c[8]) );
  XNOR U119 ( .A(b[89]), .B(n118), .Z(c[89]) );
  XNOR U120 ( .A(b[899]), .B(n119), .Z(c[899]) );
  XNOR U121 ( .A(b[898]), .B(n120), .Z(c[898]) );
  XNOR U122 ( .A(b[897]), .B(n121), .Z(c[897]) );
  XNOR U123 ( .A(b[896]), .B(n122), .Z(c[896]) );
  XNOR U124 ( .A(b[895]), .B(n123), .Z(c[895]) );
  XNOR U125 ( .A(b[894]), .B(n124), .Z(c[894]) );
  XNOR U126 ( .A(b[893]), .B(n125), .Z(c[893]) );
  XNOR U127 ( .A(b[892]), .B(n126), .Z(c[892]) );
  XNOR U128 ( .A(b[891]), .B(n127), .Z(c[891]) );
  XNOR U129 ( .A(b[890]), .B(n128), .Z(c[890]) );
  XNOR U130 ( .A(b[88]), .B(n129), .Z(c[88]) );
  XNOR U131 ( .A(b[889]), .B(n130), .Z(c[889]) );
  XNOR U132 ( .A(b[888]), .B(n131), .Z(c[888]) );
  XNOR U133 ( .A(b[887]), .B(n132), .Z(c[887]) );
  XNOR U134 ( .A(b[886]), .B(n133), .Z(c[886]) );
  XNOR U135 ( .A(b[885]), .B(n134), .Z(c[885]) );
  XNOR U136 ( .A(b[884]), .B(n135), .Z(c[884]) );
  XNOR U137 ( .A(b[883]), .B(n136), .Z(c[883]) );
  XNOR U138 ( .A(b[882]), .B(n137), .Z(c[882]) );
  XNOR U139 ( .A(b[881]), .B(n138), .Z(c[881]) );
  XNOR U140 ( .A(b[880]), .B(n139), .Z(c[880]) );
  XNOR U141 ( .A(b[87]), .B(n140), .Z(c[87]) );
  XNOR U142 ( .A(b[879]), .B(n141), .Z(c[879]) );
  XNOR U143 ( .A(b[878]), .B(n142), .Z(c[878]) );
  XNOR U144 ( .A(b[877]), .B(n143), .Z(c[877]) );
  XNOR U145 ( .A(b[876]), .B(n144), .Z(c[876]) );
  XNOR U146 ( .A(b[875]), .B(n145), .Z(c[875]) );
  XNOR U147 ( .A(b[874]), .B(n146), .Z(c[874]) );
  XNOR U148 ( .A(b[873]), .B(n147), .Z(c[873]) );
  XNOR U149 ( .A(b[872]), .B(n148), .Z(c[872]) );
  XNOR U150 ( .A(b[871]), .B(n149), .Z(c[871]) );
  XNOR U151 ( .A(b[870]), .B(n150), .Z(c[870]) );
  XNOR U152 ( .A(b[86]), .B(n151), .Z(c[86]) );
  XNOR U153 ( .A(b[869]), .B(n152), .Z(c[869]) );
  XNOR U154 ( .A(b[868]), .B(n153), .Z(c[868]) );
  XNOR U155 ( .A(b[867]), .B(n154), .Z(c[867]) );
  XNOR U156 ( .A(b[866]), .B(n155), .Z(c[866]) );
  XNOR U157 ( .A(b[865]), .B(n156), .Z(c[865]) );
  XNOR U158 ( .A(b[864]), .B(n157), .Z(c[864]) );
  XNOR U159 ( .A(b[863]), .B(n158), .Z(c[863]) );
  XNOR U160 ( .A(b[862]), .B(n159), .Z(c[862]) );
  XNOR U161 ( .A(b[861]), .B(n160), .Z(c[861]) );
  XNOR U162 ( .A(b[860]), .B(n161), .Z(c[860]) );
  XNOR U163 ( .A(b[85]), .B(n162), .Z(c[85]) );
  XNOR U164 ( .A(b[859]), .B(n163), .Z(c[859]) );
  XNOR U165 ( .A(b[858]), .B(n164), .Z(c[858]) );
  XNOR U166 ( .A(b[857]), .B(n165), .Z(c[857]) );
  XNOR U167 ( .A(b[856]), .B(n166), .Z(c[856]) );
  XNOR U168 ( .A(b[855]), .B(n167), .Z(c[855]) );
  XNOR U169 ( .A(b[854]), .B(n168), .Z(c[854]) );
  XNOR U170 ( .A(b[853]), .B(n169), .Z(c[853]) );
  XNOR U171 ( .A(b[852]), .B(n170), .Z(c[852]) );
  XNOR U172 ( .A(b[851]), .B(n171), .Z(c[851]) );
  XNOR U173 ( .A(b[850]), .B(n172), .Z(c[850]) );
  XNOR U174 ( .A(b[84]), .B(n173), .Z(c[84]) );
  XNOR U175 ( .A(b[849]), .B(n174), .Z(c[849]) );
  XNOR U176 ( .A(b[848]), .B(n175), .Z(c[848]) );
  XNOR U177 ( .A(b[847]), .B(n176), .Z(c[847]) );
  XNOR U178 ( .A(b[846]), .B(n177), .Z(c[846]) );
  XNOR U179 ( .A(b[845]), .B(n178), .Z(c[845]) );
  XNOR U180 ( .A(b[844]), .B(n179), .Z(c[844]) );
  XNOR U181 ( .A(b[843]), .B(n180), .Z(c[843]) );
  XNOR U182 ( .A(b[842]), .B(n181), .Z(c[842]) );
  XNOR U183 ( .A(b[841]), .B(n182), .Z(c[841]) );
  XNOR U184 ( .A(b[840]), .B(n183), .Z(c[840]) );
  XNOR U185 ( .A(b[83]), .B(n184), .Z(c[83]) );
  XNOR U186 ( .A(b[839]), .B(n185), .Z(c[839]) );
  XNOR U187 ( .A(b[838]), .B(n186), .Z(c[838]) );
  XNOR U188 ( .A(b[837]), .B(n187), .Z(c[837]) );
  XNOR U189 ( .A(b[836]), .B(n188), .Z(c[836]) );
  XNOR U190 ( .A(b[835]), .B(n189), .Z(c[835]) );
  XNOR U191 ( .A(b[834]), .B(n190), .Z(c[834]) );
  XNOR U192 ( .A(b[833]), .B(n191), .Z(c[833]) );
  XNOR U193 ( .A(b[832]), .B(n192), .Z(c[832]) );
  XNOR U194 ( .A(b[831]), .B(n193), .Z(c[831]) );
  XNOR U195 ( .A(b[830]), .B(n194), .Z(c[830]) );
  XNOR U196 ( .A(b[82]), .B(n195), .Z(c[82]) );
  XNOR U197 ( .A(b[829]), .B(n196), .Z(c[829]) );
  XNOR U198 ( .A(b[828]), .B(n197), .Z(c[828]) );
  XNOR U199 ( .A(b[827]), .B(n198), .Z(c[827]) );
  XNOR U200 ( .A(b[826]), .B(n199), .Z(c[826]) );
  XNOR U201 ( .A(b[825]), .B(n200), .Z(c[825]) );
  XNOR U202 ( .A(b[824]), .B(n201), .Z(c[824]) );
  XNOR U203 ( .A(b[823]), .B(n202), .Z(c[823]) );
  XNOR U204 ( .A(b[822]), .B(n203), .Z(c[822]) );
  XNOR U205 ( .A(b[821]), .B(n204), .Z(c[821]) );
  XNOR U206 ( .A(b[820]), .B(n205), .Z(c[820]) );
  XNOR U207 ( .A(b[81]), .B(n206), .Z(c[81]) );
  XNOR U208 ( .A(b[819]), .B(n207), .Z(c[819]) );
  XNOR U209 ( .A(b[818]), .B(n208), .Z(c[818]) );
  XNOR U210 ( .A(b[817]), .B(n209), .Z(c[817]) );
  XNOR U211 ( .A(b[816]), .B(n210), .Z(c[816]) );
  XNOR U212 ( .A(b[815]), .B(n211), .Z(c[815]) );
  XNOR U213 ( .A(b[814]), .B(n212), .Z(c[814]) );
  XNOR U214 ( .A(b[813]), .B(n213), .Z(c[813]) );
  XNOR U215 ( .A(b[812]), .B(n214), .Z(c[812]) );
  XNOR U216 ( .A(b[811]), .B(n215), .Z(c[811]) );
  XNOR U217 ( .A(b[810]), .B(n216), .Z(c[810]) );
  XNOR U218 ( .A(b[80]), .B(n217), .Z(c[80]) );
  XNOR U219 ( .A(b[809]), .B(n218), .Z(c[809]) );
  XNOR U220 ( .A(b[808]), .B(n219), .Z(c[808]) );
  XNOR U221 ( .A(b[807]), .B(n220), .Z(c[807]) );
  XNOR U222 ( .A(b[806]), .B(n221), .Z(c[806]) );
  XNOR U223 ( .A(b[805]), .B(n222), .Z(c[805]) );
  XNOR U224 ( .A(b[804]), .B(n223), .Z(c[804]) );
  XNOR U225 ( .A(b[803]), .B(n224), .Z(c[803]) );
  XNOR U226 ( .A(b[802]), .B(n225), .Z(c[802]) );
  XNOR U227 ( .A(b[801]), .B(n226), .Z(c[801]) );
  XNOR U228 ( .A(b[800]), .B(n227), .Z(c[800]) );
  XNOR U229 ( .A(b[7]), .B(n228), .Z(c[7]) );
  XNOR U230 ( .A(b[79]), .B(n229), .Z(c[79]) );
  XNOR U231 ( .A(b[799]), .B(n230), .Z(c[799]) );
  XNOR U232 ( .A(b[798]), .B(n231), .Z(c[798]) );
  XNOR U233 ( .A(b[797]), .B(n232), .Z(c[797]) );
  XNOR U234 ( .A(b[796]), .B(n233), .Z(c[796]) );
  XNOR U235 ( .A(b[795]), .B(n234), .Z(c[795]) );
  XNOR U236 ( .A(b[794]), .B(n235), .Z(c[794]) );
  XNOR U237 ( .A(b[793]), .B(n236), .Z(c[793]) );
  XNOR U238 ( .A(b[792]), .B(n237), .Z(c[792]) );
  XNOR U239 ( .A(b[791]), .B(n238), .Z(c[791]) );
  XNOR U240 ( .A(b[790]), .B(n239), .Z(c[790]) );
  XNOR U241 ( .A(b[78]), .B(n240), .Z(c[78]) );
  XNOR U242 ( .A(b[789]), .B(n241), .Z(c[789]) );
  XNOR U243 ( .A(b[788]), .B(n242), .Z(c[788]) );
  XNOR U244 ( .A(b[787]), .B(n243), .Z(c[787]) );
  XNOR U245 ( .A(b[786]), .B(n244), .Z(c[786]) );
  XNOR U246 ( .A(b[785]), .B(n245), .Z(c[785]) );
  XNOR U247 ( .A(b[784]), .B(n246), .Z(c[784]) );
  XNOR U248 ( .A(b[783]), .B(n247), .Z(c[783]) );
  XNOR U249 ( .A(b[782]), .B(n248), .Z(c[782]) );
  XNOR U250 ( .A(b[781]), .B(n249), .Z(c[781]) );
  XNOR U251 ( .A(b[780]), .B(n250), .Z(c[780]) );
  XNOR U252 ( .A(b[77]), .B(n251), .Z(c[77]) );
  XNOR U253 ( .A(b[779]), .B(n252), .Z(c[779]) );
  XNOR U254 ( .A(b[778]), .B(n253), .Z(c[778]) );
  XNOR U255 ( .A(b[777]), .B(n254), .Z(c[777]) );
  XNOR U256 ( .A(b[776]), .B(n255), .Z(c[776]) );
  XNOR U257 ( .A(b[775]), .B(n256), .Z(c[775]) );
  XNOR U258 ( .A(b[774]), .B(n257), .Z(c[774]) );
  XNOR U259 ( .A(b[773]), .B(n258), .Z(c[773]) );
  XNOR U260 ( .A(b[772]), .B(n259), .Z(c[772]) );
  XNOR U261 ( .A(b[771]), .B(n260), .Z(c[771]) );
  XNOR U262 ( .A(b[770]), .B(n261), .Z(c[770]) );
  XNOR U263 ( .A(b[76]), .B(n262), .Z(c[76]) );
  XNOR U264 ( .A(b[769]), .B(n263), .Z(c[769]) );
  XNOR U265 ( .A(b[768]), .B(n264), .Z(c[768]) );
  XNOR U266 ( .A(b[767]), .B(n265), .Z(c[767]) );
  XNOR U267 ( .A(b[766]), .B(n266), .Z(c[766]) );
  XNOR U268 ( .A(b[765]), .B(n267), .Z(c[765]) );
  XNOR U269 ( .A(b[764]), .B(n268), .Z(c[764]) );
  XNOR U270 ( .A(b[763]), .B(n269), .Z(c[763]) );
  XNOR U271 ( .A(b[762]), .B(n270), .Z(c[762]) );
  XNOR U272 ( .A(b[761]), .B(n271), .Z(c[761]) );
  XNOR U273 ( .A(b[760]), .B(n272), .Z(c[760]) );
  XNOR U274 ( .A(b[75]), .B(n273), .Z(c[75]) );
  XNOR U275 ( .A(b[759]), .B(n274), .Z(c[759]) );
  XNOR U276 ( .A(b[758]), .B(n275), .Z(c[758]) );
  XNOR U277 ( .A(b[757]), .B(n276), .Z(c[757]) );
  XNOR U278 ( .A(b[756]), .B(n277), .Z(c[756]) );
  XNOR U279 ( .A(b[755]), .B(n278), .Z(c[755]) );
  XNOR U280 ( .A(b[754]), .B(n279), .Z(c[754]) );
  XNOR U281 ( .A(b[753]), .B(n280), .Z(c[753]) );
  XNOR U282 ( .A(b[752]), .B(n281), .Z(c[752]) );
  XNOR U283 ( .A(b[751]), .B(n282), .Z(c[751]) );
  XNOR U284 ( .A(b[750]), .B(n283), .Z(c[750]) );
  XNOR U285 ( .A(b[74]), .B(n284), .Z(c[74]) );
  XNOR U286 ( .A(b[749]), .B(n285), .Z(c[749]) );
  XNOR U287 ( .A(b[748]), .B(n286), .Z(c[748]) );
  XNOR U288 ( .A(b[747]), .B(n287), .Z(c[747]) );
  XNOR U289 ( .A(b[746]), .B(n288), .Z(c[746]) );
  XNOR U290 ( .A(b[745]), .B(n289), .Z(c[745]) );
  XNOR U291 ( .A(b[744]), .B(n290), .Z(c[744]) );
  XNOR U292 ( .A(b[743]), .B(n291), .Z(c[743]) );
  XNOR U293 ( .A(b[742]), .B(n292), .Z(c[742]) );
  XNOR U294 ( .A(b[741]), .B(n293), .Z(c[741]) );
  XNOR U295 ( .A(b[740]), .B(n294), .Z(c[740]) );
  XNOR U296 ( .A(b[73]), .B(n295), .Z(c[73]) );
  XNOR U297 ( .A(b[739]), .B(n296), .Z(c[739]) );
  XNOR U298 ( .A(b[738]), .B(n297), .Z(c[738]) );
  XNOR U299 ( .A(b[737]), .B(n298), .Z(c[737]) );
  XNOR U300 ( .A(b[736]), .B(n299), .Z(c[736]) );
  XNOR U301 ( .A(b[735]), .B(n300), .Z(c[735]) );
  XNOR U302 ( .A(b[734]), .B(n301), .Z(c[734]) );
  XNOR U303 ( .A(b[733]), .B(n302), .Z(c[733]) );
  XNOR U304 ( .A(b[732]), .B(n303), .Z(c[732]) );
  XNOR U305 ( .A(b[731]), .B(n304), .Z(c[731]) );
  XNOR U306 ( .A(b[730]), .B(n305), .Z(c[730]) );
  XNOR U307 ( .A(b[72]), .B(n306), .Z(c[72]) );
  XNOR U308 ( .A(b[729]), .B(n307), .Z(c[729]) );
  XNOR U309 ( .A(b[728]), .B(n308), .Z(c[728]) );
  XNOR U310 ( .A(b[727]), .B(n309), .Z(c[727]) );
  XNOR U311 ( .A(b[726]), .B(n310), .Z(c[726]) );
  XNOR U312 ( .A(b[725]), .B(n311), .Z(c[725]) );
  XNOR U313 ( .A(b[724]), .B(n312), .Z(c[724]) );
  XNOR U314 ( .A(b[723]), .B(n313), .Z(c[723]) );
  XNOR U315 ( .A(b[722]), .B(n314), .Z(c[722]) );
  XNOR U316 ( .A(b[721]), .B(n315), .Z(c[721]) );
  XNOR U317 ( .A(b[720]), .B(n316), .Z(c[720]) );
  XNOR U318 ( .A(b[71]), .B(n317), .Z(c[71]) );
  XNOR U319 ( .A(b[719]), .B(n318), .Z(c[719]) );
  XNOR U320 ( .A(b[718]), .B(n319), .Z(c[718]) );
  XNOR U321 ( .A(b[717]), .B(n320), .Z(c[717]) );
  XNOR U322 ( .A(b[716]), .B(n321), .Z(c[716]) );
  XNOR U323 ( .A(b[715]), .B(n322), .Z(c[715]) );
  XNOR U324 ( .A(b[714]), .B(n323), .Z(c[714]) );
  XNOR U325 ( .A(b[713]), .B(n324), .Z(c[713]) );
  XNOR U326 ( .A(b[712]), .B(n325), .Z(c[712]) );
  XNOR U327 ( .A(b[711]), .B(n326), .Z(c[711]) );
  XNOR U328 ( .A(b[710]), .B(n327), .Z(c[710]) );
  XNOR U329 ( .A(b[70]), .B(n328), .Z(c[70]) );
  XNOR U330 ( .A(b[709]), .B(n329), .Z(c[709]) );
  XNOR U331 ( .A(b[708]), .B(n330), .Z(c[708]) );
  XNOR U332 ( .A(b[707]), .B(n331), .Z(c[707]) );
  XNOR U333 ( .A(b[706]), .B(n332), .Z(c[706]) );
  XNOR U334 ( .A(b[705]), .B(n333), .Z(c[705]) );
  XNOR U335 ( .A(b[704]), .B(n334), .Z(c[704]) );
  XNOR U336 ( .A(b[703]), .B(n335), .Z(c[703]) );
  XNOR U337 ( .A(b[702]), .B(n336), .Z(c[702]) );
  XNOR U338 ( .A(b[701]), .B(n337), .Z(c[701]) );
  XNOR U339 ( .A(b[700]), .B(n338), .Z(c[700]) );
  XNOR U340 ( .A(b[6]), .B(n339), .Z(c[6]) );
  XNOR U341 ( .A(b[69]), .B(n340), .Z(c[69]) );
  XNOR U342 ( .A(b[699]), .B(n341), .Z(c[699]) );
  XNOR U343 ( .A(b[698]), .B(n342), .Z(c[698]) );
  XNOR U344 ( .A(b[697]), .B(n343), .Z(c[697]) );
  XNOR U345 ( .A(b[696]), .B(n344), .Z(c[696]) );
  XNOR U346 ( .A(b[695]), .B(n345), .Z(c[695]) );
  XNOR U347 ( .A(b[694]), .B(n346), .Z(c[694]) );
  XNOR U348 ( .A(b[693]), .B(n347), .Z(c[693]) );
  XNOR U349 ( .A(b[692]), .B(n348), .Z(c[692]) );
  XNOR U350 ( .A(b[691]), .B(n349), .Z(c[691]) );
  XNOR U351 ( .A(b[690]), .B(n350), .Z(c[690]) );
  XNOR U352 ( .A(b[68]), .B(n351), .Z(c[68]) );
  XNOR U353 ( .A(b[689]), .B(n352), .Z(c[689]) );
  XNOR U354 ( .A(b[688]), .B(n353), .Z(c[688]) );
  XNOR U355 ( .A(b[687]), .B(n354), .Z(c[687]) );
  XNOR U356 ( .A(b[686]), .B(n355), .Z(c[686]) );
  XNOR U357 ( .A(b[685]), .B(n356), .Z(c[685]) );
  XNOR U358 ( .A(b[684]), .B(n357), .Z(c[684]) );
  XNOR U359 ( .A(b[683]), .B(n358), .Z(c[683]) );
  XNOR U360 ( .A(b[682]), .B(n359), .Z(c[682]) );
  XNOR U361 ( .A(b[681]), .B(n360), .Z(c[681]) );
  XNOR U362 ( .A(b[680]), .B(n361), .Z(c[680]) );
  XNOR U363 ( .A(b[67]), .B(n362), .Z(c[67]) );
  XNOR U364 ( .A(b[679]), .B(n363), .Z(c[679]) );
  XNOR U365 ( .A(b[678]), .B(n364), .Z(c[678]) );
  XNOR U366 ( .A(b[677]), .B(n365), .Z(c[677]) );
  XNOR U367 ( .A(b[676]), .B(n366), .Z(c[676]) );
  XNOR U368 ( .A(b[675]), .B(n367), .Z(c[675]) );
  XNOR U369 ( .A(b[674]), .B(n368), .Z(c[674]) );
  XNOR U370 ( .A(b[673]), .B(n369), .Z(c[673]) );
  XNOR U371 ( .A(b[672]), .B(n370), .Z(c[672]) );
  XNOR U372 ( .A(b[671]), .B(n371), .Z(c[671]) );
  XNOR U373 ( .A(b[670]), .B(n372), .Z(c[670]) );
  XNOR U374 ( .A(b[66]), .B(n373), .Z(c[66]) );
  XNOR U375 ( .A(b[669]), .B(n374), .Z(c[669]) );
  XNOR U376 ( .A(b[668]), .B(n375), .Z(c[668]) );
  XNOR U377 ( .A(b[667]), .B(n376), .Z(c[667]) );
  XNOR U378 ( .A(b[666]), .B(n377), .Z(c[666]) );
  XNOR U379 ( .A(b[665]), .B(n378), .Z(c[665]) );
  XNOR U380 ( .A(b[664]), .B(n379), .Z(c[664]) );
  XNOR U381 ( .A(b[663]), .B(n380), .Z(c[663]) );
  XNOR U382 ( .A(b[662]), .B(n381), .Z(c[662]) );
  XNOR U383 ( .A(b[661]), .B(n382), .Z(c[661]) );
  XNOR U384 ( .A(b[660]), .B(n383), .Z(c[660]) );
  XNOR U385 ( .A(b[65]), .B(n384), .Z(c[65]) );
  XNOR U386 ( .A(b[659]), .B(n385), .Z(c[659]) );
  XNOR U387 ( .A(b[658]), .B(n386), .Z(c[658]) );
  XNOR U388 ( .A(b[657]), .B(n387), .Z(c[657]) );
  XNOR U389 ( .A(b[656]), .B(n388), .Z(c[656]) );
  XNOR U390 ( .A(b[655]), .B(n389), .Z(c[655]) );
  XNOR U391 ( .A(b[654]), .B(n390), .Z(c[654]) );
  XNOR U392 ( .A(b[653]), .B(n391), .Z(c[653]) );
  XNOR U393 ( .A(b[652]), .B(n392), .Z(c[652]) );
  XNOR U394 ( .A(b[651]), .B(n393), .Z(c[651]) );
  XNOR U395 ( .A(b[650]), .B(n394), .Z(c[650]) );
  XNOR U396 ( .A(b[64]), .B(n395), .Z(c[64]) );
  XNOR U397 ( .A(b[649]), .B(n396), .Z(c[649]) );
  XNOR U398 ( .A(b[648]), .B(n397), .Z(c[648]) );
  XNOR U399 ( .A(b[647]), .B(n398), .Z(c[647]) );
  XNOR U400 ( .A(b[646]), .B(n399), .Z(c[646]) );
  XNOR U401 ( .A(b[645]), .B(n400), .Z(c[645]) );
  XNOR U402 ( .A(b[644]), .B(n401), .Z(c[644]) );
  XNOR U403 ( .A(b[643]), .B(n402), .Z(c[643]) );
  XNOR U404 ( .A(b[642]), .B(n403), .Z(c[642]) );
  XNOR U405 ( .A(b[641]), .B(n404), .Z(c[641]) );
  XNOR U406 ( .A(b[640]), .B(n405), .Z(c[640]) );
  XNOR U407 ( .A(b[63]), .B(n406), .Z(c[63]) );
  XNOR U408 ( .A(b[639]), .B(n407), .Z(c[639]) );
  XNOR U409 ( .A(b[638]), .B(n408), .Z(c[638]) );
  XNOR U410 ( .A(b[637]), .B(n409), .Z(c[637]) );
  XNOR U411 ( .A(b[636]), .B(n410), .Z(c[636]) );
  XNOR U412 ( .A(b[635]), .B(n411), .Z(c[635]) );
  XNOR U413 ( .A(b[634]), .B(n412), .Z(c[634]) );
  XNOR U414 ( .A(b[633]), .B(n413), .Z(c[633]) );
  XNOR U415 ( .A(b[632]), .B(n414), .Z(c[632]) );
  XNOR U416 ( .A(b[631]), .B(n415), .Z(c[631]) );
  XNOR U417 ( .A(b[630]), .B(n416), .Z(c[630]) );
  XNOR U418 ( .A(b[62]), .B(n417), .Z(c[62]) );
  XNOR U419 ( .A(b[629]), .B(n418), .Z(c[629]) );
  XNOR U420 ( .A(b[628]), .B(n419), .Z(c[628]) );
  XNOR U421 ( .A(b[627]), .B(n420), .Z(c[627]) );
  XNOR U422 ( .A(b[626]), .B(n421), .Z(c[626]) );
  XNOR U423 ( .A(b[625]), .B(n422), .Z(c[625]) );
  XNOR U424 ( .A(b[624]), .B(n423), .Z(c[624]) );
  XNOR U425 ( .A(b[623]), .B(n424), .Z(c[623]) );
  XNOR U426 ( .A(b[622]), .B(n425), .Z(c[622]) );
  XNOR U427 ( .A(b[621]), .B(n426), .Z(c[621]) );
  XNOR U428 ( .A(b[620]), .B(n427), .Z(c[620]) );
  XNOR U429 ( .A(b[61]), .B(n428), .Z(c[61]) );
  XNOR U430 ( .A(b[619]), .B(n429), .Z(c[619]) );
  XNOR U431 ( .A(b[618]), .B(n430), .Z(c[618]) );
  XNOR U432 ( .A(b[617]), .B(n431), .Z(c[617]) );
  XNOR U433 ( .A(b[616]), .B(n432), .Z(c[616]) );
  XNOR U434 ( .A(b[615]), .B(n433), .Z(c[615]) );
  XNOR U435 ( .A(b[614]), .B(n434), .Z(c[614]) );
  XNOR U436 ( .A(b[613]), .B(n435), .Z(c[613]) );
  XNOR U437 ( .A(b[612]), .B(n436), .Z(c[612]) );
  XNOR U438 ( .A(b[611]), .B(n437), .Z(c[611]) );
  XNOR U439 ( .A(b[610]), .B(n438), .Z(c[610]) );
  XNOR U440 ( .A(b[60]), .B(n439), .Z(c[60]) );
  XNOR U441 ( .A(b[609]), .B(n440), .Z(c[609]) );
  XNOR U442 ( .A(b[608]), .B(n441), .Z(c[608]) );
  XNOR U443 ( .A(b[607]), .B(n442), .Z(c[607]) );
  XNOR U444 ( .A(b[606]), .B(n443), .Z(c[606]) );
  XNOR U445 ( .A(b[605]), .B(n444), .Z(c[605]) );
  XNOR U446 ( .A(b[604]), .B(n445), .Z(c[604]) );
  XNOR U447 ( .A(b[603]), .B(n446), .Z(c[603]) );
  XNOR U448 ( .A(b[602]), .B(n447), .Z(c[602]) );
  XNOR U449 ( .A(b[601]), .B(n448), .Z(c[601]) );
  XNOR U450 ( .A(b[600]), .B(n449), .Z(c[600]) );
  XNOR U451 ( .A(b[5]), .B(n450), .Z(c[5]) );
  XNOR U452 ( .A(b[59]), .B(n451), .Z(c[59]) );
  XNOR U453 ( .A(b[599]), .B(n452), .Z(c[599]) );
  XNOR U454 ( .A(b[598]), .B(n453), .Z(c[598]) );
  XNOR U455 ( .A(b[597]), .B(n454), .Z(c[597]) );
  XNOR U456 ( .A(b[596]), .B(n455), .Z(c[596]) );
  XNOR U457 ( .A(b[595]), .B(n456), .Z(c[595]) );
  XNOR U458 ( .A(b[594]), .B(n457), .Z(c[594]) );
  XNOR U459 ( .A(b[593]), .B(n458), .Z(c[593]) );
  XNOR U460 ( .A(b[592]), .B(n459), .Z(c[592]) );
  XNOR U461 ( .A(b[591]), .B(n460), .Z(c[591]) );
  XNOR U462 ( .A(b[590]), .B(n461), .Z(c[590]) );
  XNOR U463 ( .A(b[58]), .B(n462), .Z(c[58]) );
  XNOR U464 ( .A(b[589]), .B(n463), .Z(c[589]) );
  XNOR U465 ( .A(b[588]), .B(n464), .Z(c[588]) );
  XNOR U466 ( .A(b[587]), .B(n465), .Z(c[587]) );
  XNOR U467 ( .A(b[586]), .B(n466), .Z(c[586]) );
  XNOR U468 ( .A(b[585]), .B(n467), .Z(c[585]) );
  XNOR U469 ( .A(b[584]), .B(n468), .Z(c[584]) );
  XNOR U470 ( .A(b[583]), .B(n469), .Z(c[583]) );
  XNOR U471 ( .A(b[582]), .B(n470), .Z(c[582]) );
  XNOR U472 ( .A(b[581]), .B(n471), .Z(c[581]) );
  XNOR U473 ( .A(b[580]), .B(n472), .Z(c[580]) );
  XNOR U474 ( .A(b[57]), .B(n473), .Z(c[57]) );
  XNOR U475 ( .A(b[579]), .B(n474), .Z(c[579]) );
  XNOR U476 ( .A(b[578]), .B(n475), .Z(c[578]) );
  XNOR U477 ( .A(b[577]), .B(n476), .Z(c[577]) );
  XNOR U478 ( .A(b[576]), .B(n477), .Z(c[576]) );
  XNOR U479 ( .A(b[575]), .B(n478), .Z(c[575]) );
  XNOR U480 ( .A(b[574]), .B(n479), .Z(c[574]) );
  XNOR U481 ( .A(b[573]), .B(n480), .Z(c[573]) );
  XNOR U482 ( .A(b[572]), .B(n481), .Z(c[572]) );
  XNOR U483 ( .A(b[571]), .B(n482), .Z(c[571]) );
  XNOR U484 ( .A(b[570]), .B(n483), .Z(c[570]) );
  XNOR U485 ( .A(b[56]), .B(n484), .Z(c[56]) );
  XNOR U486 ( .A(b[569]), .B(n485), .Z(c[569]) );
  XNOR U487 ( .A(b[568]), .B(n486), .Z(c[568]) );
  XNOR U488 ( .A(b[567]), .B(n487), .Z(c[567]) );
  XNOR U489 ( .A(b[566]), .B(n488), .Z(c[566]) );
  XNOR U490 ( .A(b[565]), .B(n489), .Z(c[565]) );
  XNOR U491 ( .A(b[564]), .B(n490), .Z(c[564]) );
  XNOR U492 ( .A(b[563]), .B(n491), .Z(c[563]) );
  XNOR U493 ( .A(b[562]), .B(n492), .Z(c[562]) );
  XNOR U494 ( .A(b[561]), .B(n493), .Z(c[561]) );
  XNOR U495 ( .A(b[560]), .B(n494), .Z(c[560]) );
  XNOR U496 ( .A(b[55]), .B(n495), .Z(c[55]) );
  XNOR U497 ( .A(b[559]), .B(n496), .Z(c[559]) );
  XNOR U498 ( .A(b[558]), .B(n497), .Z(c[558]) );
  XNOR U499 ( .A(b[557]), .B(n498), .Z(c[557]) );
  XNOR U500 ( .A(b[556]), .B(n499), .Z(c[556]) );
  XNOR U501 ( .A(b[555]), .B(n500), .Z(c[555]) );
  XNOR U502 ( .A(b[554]), .B(n501), .Z(c[554]) );
  XNOR U503 ( .A(b[553]), .B(n502), .Z(c[553]) );
  XNOR U504 ( .A(b[552]), .B(n503), .Z(c[552]) );
  XNOR U505 ( .A(b[551]), .B(n504), .Z(c[551]) );
  XNOR U506 ( .A(b[550]), .B(n505), .Z(c[550]) );
  XNOR U507 ( .A(b[54]), .B(n506), .Z(c[54]) );
  XNOR U508 ( .A(b[549]), .B(n507), .Z(c[549]) );
  XNOR U509 ( .A(b[548]), .B(n508), .Z(c[548]) );
  XNOR U510 ( .A(b[547]), .B(n509), .Z(c[547]) );
  XNOR U511 ( .A(b[546]), .B(n510), .Z(c[546]) );
  XNOR U512 ( .A(b[545]), .B(n511), .Z(c[545]) );
  XNOR U513 ( .A(b[544]), .B(n512), .Z(c[544]) );
  XNOR U514 ( .A(b[543]), .B(n513), .Z(c[543]) );
  XNOR U515 ( .A(b[542]), .B(n514), .Z(c[542]) );
  XNOR U516 ( .A(b[541]), .B(n515), .Z(c[541]) );
  XNOR U517 ( .A(b[540]), .B(n516), .Z(c[540]) );
  XNOR U518 ( .A(b[53]), .B(n517), .Z(c[53]) );
  XNOR U519 ( .A(b[539]), .B(n518), .Z(c[539]) );
  XNOR U520 ( .A(b[538]), .B(n519), .Z(c[538]) );
  XNOR U521 ( .A(b[537]), .B(n520), .Z(c[537]) );
  XNOR U522 ( .A(b[536]), .B(n521), .Z(c[536]) );
  XNOR U523 ( .A(b[535]), .B(n522), .Z(c[535]) );
  XNOR U524 ( .A(b[534]), .B(n523), .Z(c[534]) );
  XNOR U525 ( .A(b[533]), .B(n524), .Z(c[533]) );
  XNOR U526 ( .A(b[532]), .B(n525), .Z(c[532]) );
  XNOR U527 ( .A(b[531]), .B(n526), .Z(c[531]) );
  XNOR U528 ( .A(b[530]), .B(n527), .Z(c[530]) );
  XNOR U529 ( .A(b[52]), .B(n528), .Z(c[52]) );
  XNOR U530 ( .A(b[529]), .B(n529), .Z(c[529]) );
  XNOR U531 ( .A(b[528]), .B(n530), .Z(c[528]) );
  XNOR U532 ( .A(b[527]), .B(n531), .Z(c[527]) );
  XNOR U533 ( .A(b[526]), .B(n532), .Z(c[526]) );
  XNOR U534 ( .A(b[525]), .B(n533), .Z(c[525]) );
  XNOR U535 ( .A(b[524]), .B(n534), .Z(c[524]) );
  XNOR U536 ( .A(b[523]), .B(n535), .Z(c[523]) );
  XNOR U537 ( .A(b[522]), .B(n536), .Z(c[522]) );
  XNOR U538 ( .A(b[521]), .B(n537), .Z(c[521]) );
  XNOR U539 ( .A(b[520]), .B(n538), .Z(c[520]) );
  XNOR U540 ( .A(b[51]), .B(n539), .Z(c[51]) );
  XNOR U541 ( .A(b[519]), .B(n540), .Z(c[519]) );
  XNOR U542 ( .A(b[518]), .B(n541), .Z(c[518]) );
  XNOR U543 ( .A(b[517]), .B(n542), .Z(c[517]) );
  XNOR U544 ( .A(b[516]), .B(n543), .Z(c[516]) );
  XNOR U545 ( .A(b[515]), .B(n544), .Z(c[515]) );
  XNOR U546 ( .A(b[514]), .B(n545), .Z(c[514]) );
  XNOR U547 ( .A(b[513]), .B(n546), .Z(c[513]) );
  XNOR U548 ( .A(b[512]), .B(n547), .Z(c[512]) );
  XNOR U549 ( .A(b[511]), .B(n548), .Z(c[511]) );
  XNOR U550 ( .A(b[510]), .B(n549), .Z(c[510]) );
  XNOR U551 ( .A(b[50]), .B(n550), .Z(c[50]) );
  XNOR U552 ( .A(b[509]), .B(n551), .Z(c[509]) );
  XNOR U553 ( .A(b[508]), .B(n552), .Z(c[508]) );
  XNOR U554 ( .A(b[507]), .B(n553), .Z(c[507]) );
  XNOR U555 ( .A(b[506]), .B(n554), .Z(c[506]) );
  XNOR U556 ( .A(b[505]), .B(n555), .Z(c[505]) );
  XNOR U557 ( .A(b[504]), .B(n556), .Z(c[504]) );
  XNOR U558 ( .A(b[503]), .B(n557), .Z(c[503]) );
  XNOR U559 ( .A(b[502]), .B(n558), .Z(c[502]) );
  XNOR U560 ( .A(b[501]), .B(n559), .Z(c[501]) );
  XNOR U561 ( .A(b[500]), .B(n560), .Z(c[500]) );
  XNOR U562 ( .A(b[4]), .B(n561), .Z(c[4]) );
  XNOR U563 ( .A(b[49]), .B(n562), .Z(c[49]) );
  XNOR U564 ( .A(b[499]), .B(n563), .Z(c[499]) );
  XNOR U565 ( .A(b[498]), .B(n564), .Z(c[498]) );
  XNOR U566 ( .A(b[497]), .B(n565), .Z(c[497]) );
  XNOR U567 ( .A(b[496]), .B(n566), .Z(c[496]) );
  XNOR U568 ( .A(b[495]), .B(n567), .Z(c[495]) );
  XNOR U569 ( .A(b[494]), .B(n568), .Z(c[494]) );
  XNOR U570 ( .A(b[493]), .B(n569), .Z(c[493]) );
  XNOR U571 ( .A(b[492]), .B(n570), .Z(c[492]) );
  XNOR U572 ( .A(b[491]), .B(n571), .Z(c[491]) );
  XNOR U573 ( .A(b[490]), .B(n572), .Z(c[490]) );
  XNOR U574 ( .A(b[48]), .B(n573), .Z(c[48]) );
  XNOR U575 ( .A(b[489]), .B(n574), .Z(c[489]) );
  XNOR U576 ( .A(b[488]), .B(n575), .Z(c[488]) );
  XNOR U577 ( .A(b[487]), .B(n576), .Z(c[487]) );
  XNOR U578 ( .A(b[486]), .B(n577), .Z(c[486]) );
  XNOR U579 ( .A(b[485]), .B(n578), .Z(c[485]) );
  XNOR U580 ( .A(b[484]), .B(n579), .Z(c[484]) );
  XNOR U581 ( .A(b[483]), .B(n580), .Z(c[483]) );
  XNOR U582 ( .A(b[482]), .B(n581), .Z(c[482]) );
  XNOR U583 ( .A(b[481]), .B(n582), .Z(c[481]) );
  XNOR U584 ( .A(b[480]), .B(n583), .Z(c[480]) );
  XNOR U585 ( .A(b[47]), .B(n584), .Z(c[47]) );
  XNOR U586 ( .A(b[479]), .B(n585), .Z(c[479]) );
  XNOR U587 ( .A(b[478]), .B(n586), .Z(c[478]) );
  XNOR U588 ( .A(b[477]), .B(n587), .Z(c[477]) );
  XNOR U589 ( .A(b[476]), .B(n588), .Z(c[476]) );
  XNOR U590 ( .A(b[475]), .B(n589), .Z(c[475]) );
  XNOR U591 ( .A(b[474]), .B(n590), .Z(c[474]) );
  XNOR U592 ( .A(b[473]), .B(n591), .Z(c[473]) );
  XNOR U593 ( .A(b[472]), .B(n592), .Z(c[472]) );
  XNOR U594 ( .A(b[471]), .B(n593), .Z(c[471]) );
  XNOR U595 ( .A(b[470]), .B(n594), .Z(c[470]) );
  XNOR U596 ( .A(b[46]), .B(n595), .Z(c[46]) );
  XNOR U597 ( .A(b[469]), .B(n596), .Z(c[469]) );
  XNOR U598 ( .A(b[468]), .B(n597), .Z(c[468]) );
  XNOR U599 ( .A(b[467]), .B(n598), .Z(c[467]) );
  XNOR U600 ( .A(b[466]), .B(n599), .Z(c[466]) );
  XNOR U601 ( .A(b[465]), .B(n600), .Z(c[465]) );
  XNOR U602 ( .A(b[464]), .B(n601), .Z(c[464]) );
  XNOR U603 ( .A(b[463]), .B(n602), .Z(c[463]) );
  XNOR U604 ( .A(b[462]), .B(n603), .Z(c[462]) );
  XNOR U605 ( .A(b[461]), .B(n604), .Z(c[461]) );
  XNOR U606 ( .A(b[460]), .B(n605), .Z(c[460]) );
  XNOR U607 ( .A(b[45]), .B(n606), .Z(c[45]) );
  XNOR U608 ( .A(b[459]), .B(n607), .Z(c[459]) );
  XNOR U609 ( .A(b[458]), .B(n608), .Z(c[458]) );
  XNOR U610 ( .A(b[457]), .B(n609), .Z(c[457]) );
  XNOR U611 ( .A(b[456]), .B(n610), .Z(c[456]) );
  XNOR U612 ( .A(b[455]), .B(n611), .Z(c[455]) );
  XNOR U613 ( .A(b[454]), .B(n612), .Z(c[454]) );
  XNOR U614 ( .A(b[453]), .B(n613), .Z(c[453]) );
  XNOR U615 ( .A(b[452]), .B(n614), .Z(c[452]) );
  XNOR U616 ( .A(b[451]), .B(n615), .Z(c[451]) );
  XNOR U617 ( .A(b[450]), .B(n616), .Z(c[450]) );
  XNOR U618 ( .A(b[44]), .B(n617), .Z(c[44]) );
  XNOR U619 ( .A(b[449]), .B(n618), .Z(c[449]) );
  XNOR U620 ( .A(b[448]), .B(n619), .Z(c[448]) );
  XNOR U621 ( .A(b[447]), .B(n620), .Z(c[447]) );
  XNOR U622 ( .A(b[446]), .B(n621), .Z(c[446]) );
  XNOR U623 ( .A(b[445]), .B(n622), .Z(c[445]) );
  XNOR U624 ( .A(b[444]), .B(n623), .Z(c[444]) );
  XNOR U625 ( .A(b[443]), .B(n624), .Z(c[443]) );
  XNOR U626 ( .A(b[442]), .B(n625), .Z(c[442]) );
  XNOR U627 ( .A(b[441]), .B(n626), .Z(c[441]) );
  XNOR U628 ( .A(b[440]), .B(n627), .Z(c[440]) );
  XNOR U629 ( .A(b[43]), .B(n628), .Z(c[43]) );
  XNOR U630 ( .A(b[439]), .B(n629), .Z(c[439]) );
  XNOR U631 ( .A(b[438]), .B(n630), .Z(c[438]) );
  XNOR U632 ( .A(b[437]), .B(n631), .Z(c[437]) );
  XNOR U633 ( .A(b[436]), .B(n632), .Z(c[436]) );
  XNOR U634 ( .A(b[435]), .B(n633), .Z(c[435]) );
  XNOR U635 ( .A(b[434]), .B(n634), .Z(c[434]) );
  XNOR U636 ( .A(b[433]), .B(n635), .Z(c[433]) );
  XNOR U637 ( .A(b[432]), .B(n636), .Z(c[432]) );
  XNOR U638 ( .A(b[431]), .B(n637), .Z(c[431]) );
  XNOR U639 ( .A(b[430]), .B(n638), .Z(c[430]) );
  XNOR U640 ( .A(b[42]), .B(n639), .Z(c[42]) );
  XNOR U641 ( .A(b[429]), .B(n640), .Z(c[429]) );
  XNOR U642 ( .A(b[428]), .B(n641), .Z(c[428]) );
  XNOR U643 ( .A(b[427]), .B(n642), .Z(c[427]) );
  XNOR U644 ( .A(b[426]), .B(n643), .Z(c[426]) );
  XNOR U645 ( .A(b[425]), .B(n644), .Z(c[425]) );
  XNOR U646 ( .A(b[424]), .B(n645), .Z(c[424]) );
  XNOR U647 ( .A(b[423]), .B(n646), .Z(c[423]) );
  XNOR U648 ( .A(b[422]), .B(n647), .Z(c[422]) );
  XNOR U649 ( .A(b[421]), .B(n648), .Z(c[421]) );
  XNOR U650 ( .A(b[420]), .B(n649), .Z(c[420]) );
  XNOR U651 ( .A(b[41]), .B(n650), .Z(c[41]) );
  XNOR U652 ( .A(b[419]), .B(n651), .Z(c[419]) );
  XNOR U653 ( .A(b[418]), .B(n652), .Z(c[418]) );
  XNOR U654 ( .A(b[417]), .B(n653), .Z(c[417]) );
  XNOR U655 ( .A(b[416]), .B(n654), .Z(c[416]) );
  XNOR U656 ( .A(b[415]), .B(n655), .Z(c[415]) );
  XNOR U657 ( .A(b[414]), .B(n656), .Z(c[414]) );
  XNOR U658 ( .A(b[413]), .B(n657), .Z(c[413]) );
  XNOR U659 ( .A(b[412]), .B(n658), .Z(c[412]) );
  XNOR U660 ( .A(b[411]), .B(n659), .Z(c[411]) );
  XNOR U661 ( .A(b[410]), .B(n660), .Z(c[410]) );
  XNOR U662 ( .A(b[40]), .B(n661), .Z(c[40]) );
  XNOR U663 ( .A(b[409]), .B(n662), .Z(c[409]) );
  XNOR U664 ( .A(b[4095]), .B(n5), .Z(c[4095]) );
  XNOR U665 ( .A(a[4095]), .B(n3), .Z(n5) );
  XNOR U666 ( .A(n663), .B(n664), .Z(n3) );
  ANDN U667 ( .B(n665), .A(n666), .Z(n663) );
  XNOR U668 ( .A(b[4094]), .B(n664), .Z(n665) );
  XNOR U669 ( .A(b[4094]), .B(n666), .Z(c[4094]) );
  XNOR U670 ( .A(a[4094]), .B(n667), .Z(n666) );
  IV U671 ( .A(n664), .Z(n667) );
  XOR U672 ( .A(n668), .B(n669), .Z(n664) );
  ANDN U673 ( .B(n670), .A(n671), .Z(n668) );
  XNOR U674 ( .A(b[4093]), .B(n669), .Z(n670) );
  XNOR U675 ( .A(b[4093]), .B(n671), .Z(c[4093]) );
  XNOR U676 ( .A(a[4093]), .B(n672), .Z(n671) );
  IV U677 ( .A(n669), .Z(n672) );
  XOR U678 ( .A(n673), .B(n674), .Z(n669) );
  ANDN U679 ( .B(n675), .A(n676), .Z(n673) );
  XNOR U680 ( .A(b[4092]), .B(n674), .Z(n675) );
  XNOR U681 ( .A(b[4092]), .B(n676), .Z(c[4092]) );
  XNOR U682 ( .A(a[4092]), .B(n677), .Z(n676) );
  IV U683 ( .A(n674), .Z(n677) );
  XOR U684 ( .A(n678), .B(n679), .Z(n674) );
  ANDN U685 ( .B(n680), .A(n681), .Z(n678) );
  XNOR U686 ( .A(b[4091]), .B(n679), .Z(n680) );
  XNOR U687 ( .A(b[4091]), .B(n681), .Z(c[4091]) );
  XNOR U688 ( .A(a[4091]), .B(n682), .Z(n681) );
  IV U689 ( .A(n679), .Z(n682) );
  XOR U690 ( .A(n683), .B(n684), .Z(n679) );
  ANDN U691 ( .B(n685), .A(n686), .Z(n683) );
  XNOR U692 ( .A(b[4090]), .B(n684), .Z(n685) );
  XNOR U693 ( .A(b[4090]), .B(n686), .Z(c[4090]) );
  XNOR U694 ( .A(a[4090]), .B(n687), .Z(n686) );
  IV U695 ( .A(n684), .Z(n687) );
  XOR U696 ( .A(n688), .B(n689), .Z(n684) );
  ANDN U697 ( .B(n690), .A(n691), .Z(n688) );
  XNOR U698 ( .A(b[4089]), .B(n689), .Z(n690) );
  XNOR U699 ( .A(b[408]), .B(n692), .Z(c[408]) );
  XNOR U700 ( .A(b[4089]), .B(n691), .Z(c[4089]) );
  XNOR U701 ( .A(a[4089]), .B(n693), .Z(n691) );
  IV U702 ( .A(n689), .Z(n693) );
  XOR U703 ( .A(n694), .B(n695), .Z(n689) );
  ANDN U704 ( .B(n696), .A(n697), .Z(n694) );
  XNOR U705 ( .A(b[4088]), .B(n695), .Z(n696) );
  XNOR U706 ( .A(b[4088]), .B(n697), .Z(c[4088]) );
  XNOR U707 ( .A(a[4088]), .B(n698), .Z(n697) );
  IV U708 ( .A(n695), .Z(n698) );
  XOR U709 ( .A(n699), .B(n700), .Z(n695) );
  ANDN U710 ( .B(n701), .A(n702), .Z(n699) );
  XNOR U711 ( .A(b[4087]), .B(n700), .Z(n701) );
  XNOR U712 ( .A(b[4087]), .B(n702), .Z(c[4087]) );
  XNOR U713 ( .A(a[4087]), .B(n703), .Z(n702) );
  IV U714 ( .A(n700), .Z(n703) );
  XOR U715 ( .A(n704), .B(n705), .Z(n700) );
  ANDN U716 ( .B(n706), .A(n707), .Z(n704) );
  XNOR U717 ( .A(b[4086]), .B(n705), .Z(n706) );
  XNOR U718 ( .A(b[4086]), .B(n707), .Z(c[4086]) );
  XNOR U719 ( .A(a[4086]), .B(n708), .Z(n707) );
  IV U720 ( .A(n705), .Z(n708) );
  XOR U721 ( .A(n709), .B(n710), .Z(n705) );
  ANDN U722 ( .B(n711), .A(n712), .Z(n709) );
  XNOR U723 ( .A(b[4085]), .B(n710), .Z(n711) );
  XNOR U724 ( .A(b[4085]), .B(n712), .Z(c[4085]) );
  XNOR U725 ( .A(a[4085]), .B(n713), .Z(n712) );
  IV U726 ( .A(n710), .Z(n713) );
  XOR U727 ( .A(n714), .B(n715), .Z(n710) );
  ANDN U728 ( .B(n716), .A(n717), .Z(n714) );
  XNOR U729 ( .A(b[4084]), .B(n715), .Z(n716) );
  XNOR U730 ( .A(b[4084]), .B(n717), .Z(c[4084]) );
  XNOR U731 ( .A(a[4084]), .B(n718), .Z(n717) );
  IV U732 ( .A(n715), .Z(n718) );
  XOR U733 ( .A(n719), .B(n720), .Z(n715) );
  ANDN U734 ( .B(n721), .A(n722), .Z(n719) );
  XNOR U735 ( .A(b[4083]), .B(n720), .Z(n721) );
  XNOR U736 ( .A(b[4083]), .B(n722), .Z(c[4083]) );
  XNOR U737 ( .A(a[4083]), .B(n723), .Z(n722) );
  IV U738 ( .A(n720), .Z(n723) );
  XOR U739 ( .A(n724), .B(n725), .Z(n720) );
  ANDN U740 ( .B(n726), .A(n727), .Z(n724) );
  XNOR U741 ( .A(b[4082]), .B(n725), .Z(n726) );
  XNOR U742 ( .A(b[4082]), .B(n727), .Z(c[4082]) );
  XNOR U743 ( .A(a[4082]), .B(n728), .Z(n727) );
  IV U744 ( .A(n725), .Z(n728) );
  XOR U745 ( .A(n729), .B(n730), .Z(n725) );
  ANDN U746 ( .B(n731), .A(n732), .Z(n729) );
  XNOR U747 ( .A(b[4081]), .B(n730), .Z(n731) );
  XNOR U748 ( .A(b[4081]), .B(n732), .Z(c[4081]) );
  XNOR U749 ( .A(a[4081]), .B(n733), .Z(n732) );
  IV U750 ( .A(n730), .Z(n733) );
  XOR U751 ( .A(n734), .B(n735), .Z(n730) );
  ANDN U752 ( .B(n736), .A(n737), .Z(n734) );
  XNOR U753 ( .A(b[4080]), .B(n735), .Z(n736) );
  XNOR U754 ( .A(b[4080]), .B(n737), .Z(c[4080]) );
  XNOR U755 ( .A(a[4080]), .B(n738), .Z(n737) );
  IV U756 ( .A(n735), .Z(n738) );
  XOR U757 ( .A(n739), .B(n740), .Z(n735) );
  ANDN U758 ( .B(n741), .A(n742), .Z(n739) );
  XNOR U759 ( .A(b[4079]), .B(n740), .Z(n741) );
  XNOR U760 ( .A(b[407]), .B(n743), .Z(c[407]) );
  XNOR U761 ( .A(b[4079]), .B(n742), .Z(c[4079]) );
  XNOR U762 ( .A(a[4079]), .B(n744), .Z(n742) );
  IV U763 ( .A(n740), .Z(n744) );
  XOR U764 ( .A(n745), .B(n746), .Z(n740) );
  ANDN U765 ( .B(n747), .A(n748), .Z(n745) );
  XNOR U766 ( .A(b[4078]), .B(n746), .Z(n747) );
  XNOR U767 ( .A(b[4078]), .B(n748), .Z(c[4078]) );
  XNOR U768 ( .A(a[4078]), .B(n749), .Z(n748) );
  IV U769 ( .A(n746), .Z(n749) );
  XOR U770 ( .A(n750), .B(n751), .Z(n746) );
  ANDN U771 ( .B(n752), .A(n753), .Z(n750) );
  XNOR U772 ( .A(b[4077]), .B(n751), .Z(n752) );
  XNOR U773 ( .A(b[4077]), .B(n753), .Z(c[4077]) );
  XNOR U774 ( .A(a[4077]), .B(n754), .Z(n753) );
  IV U775 ( .A(n751), .Z(n754) );
  XOR U776 ( .A(n755), .B(n756), .Z(n751) );
  ANDN U777 ( .B(n757), .A(n758), .Z(n755) );
  XNOR U778 ( .A(b[4076]), .B(n756), .Z(n757) );
  XNOR U779 ( .A(b[4076]), .B(n758), .Z(c[4076]) );
  XNOR U780 ( .A(a[4076]), .B(n759), .Z(n758) );
  IV U781 ( .A(n756), .Z(n759) );
  XOR U782 ( .A(n760), .B(n761), .Z(n756) );
  ANDN U783 ( .B(n762), .A(n763), .Z(n760) );
  XNOR U784 ( .A(b[4075]), .B(n761), .Z(n762) );
  XNOR U785 ( .A(b[4075]), .B(n763), .Z(c[4075]) );
  XNOR U786 ( .A(a[4075]), .B(n764), .Z(n763) );
  IV U787 ( .A(n761), .Z(n764) );
  XOR U788 ( .A(n765), .B(n766), .Z(n761) );
  ANDN U789 ( .B(n767), .A(n768), .Z(n765) );
  XNOR U790 ( .A(b[4074]), .B(n766), .Z(n767) );
  XNOR U791 ( .A(b[4074]), .B(n768), .Z(c[4074]) );
  XNOR U792 ( .A(a[4074]), .B(n769), .Z(n768) );
  IV U793 ( .A(n766), .Z(n769) );
  XOR U794 ( .A(n770), .B(n771), .Z(n766) );
  ANDN U795 ( .B(n772), .A(n773), .Z(n770) );
  XNOR U796 ( .A(b[4073]), .B(n771), .Z(n772) );
  XNOR U797 ( .A(b[4073]), .B(n773), .Z(c[4073]) );
  XNOR U798 ( .A(a[4073]), .B(n774), .Z(n773) );
  IV U799 ( .A(n771), .Z(n774) );
  XOR U800 ( .A(n775), .B(n776), .Z(n771) );
  ANDN U801 ( .B(n777), .A(n778), .Z(n775) );
  XNOR U802 ( .A(b[4072]), .B(n776), .Z(n777) );
  XNOR U803 ( .A(b[4072]), .B(n778), .Z(c[4072]) );
  XNOR U804 ( .A(a[4072]), .B(n779), .Z(n778) );
  IV U805 ( .A(n776), .Z(n779) );
  XOR U806 ( .A(n780), .B(n781), .Z(n776) );
  ANDN U807 ( .B(n782), .A(n783), .Z(n780) );
  XNOR U808 ( .A(b[4071]), .B(n781), .Z(n782) );
  XNOR U809 ( .A(b[4071]), .B(n783), .Z(c[4071]) );
  XNOR U810 ( .A(a[4071]), .B(n784), .Z(n783) );
  IV U811 ( .A(n781), .Z(n784) );
  XOR U812 ( .A(n785), .B(n786), .Z(n781) );
  ANDN U813 ( .B(n787), .A(n788), .Z(n785) );
  XNOR U814 ( .A(b[4070]), .B(n786), .Z(n787) );
  XNOR U815 ( .A(b[4070]), .B(n788), .Z(c[4070]) );
  XNOR U816 ( .A(a[4070]), .B(n789), .Z(n788) );
  IV U817 ( .A(n786), .Z(n789) );
  XOR U818 ( .A(n790), .B(n791), .Z(n786) );
  ANDN U819 ( .B(n792), .A(n793), .Z(n790) );
  XNOR U820 ( .A(b[4069]), .B(n791), .Z(n792) );
  XNOR U821 ( .A(b[406]), .B(n794), .Z(c[406]) );
  XNOR U822 ( .A(b[4069]), .B(n793), .Z(c[4069]) );
  XNOR U823 ( .A(a[4069]), .B(n795), .Z(n793) );
  IV U824 ( .A(n791), .Z(n795) );
  XOR U825 ( .A(n796), .B(n797), .Z(n791) );
  ANDN U826 ( .B(n798), .A(n799), .Z(n796) );
  XNOR U827 ( .A(b[4068]), .B(n797), .Z(n798) );
  XNOR U828 ( .A(b[4068]), .B(n799), .Z(c[4068]) );
  XNOR U829 ( .A(a[4068]), .B(n800), .Z(n799) );
  IV U830 ( .A(n797), .Z(n800) );
  XOR U831 ( .A(n801), .B(n802), .Z(n797) );
  ANDN U832 ( .B(n803), .A(n804), .Z(n801) );
  XNOR U833 ( .A(b[4067]), .B(n802), .Z(n803) );
  XNOR U834 ( .A(b[4067]), .B(n804), .Z(c[4067]) );
  XNOR U835 ( .A(a[4067]), .B(n805), .Z(n804) );
  IV U836 ( .A(n802), .Z(n805) );
  XOR U837 ( .A(n806), .B(n807), .Z(n802) );
  ANDN U838 ( .B(n808), .A(n809), .Z(n806) );
  XNOR U839 ( .A(b[4066]), .B(n807), .Z(n808) );
  XNOR U840 ( .A(b[4066]), .B(n809), .Z(c[4066]) );
  XNOR U841 ( .A(a[4066]), .B(n810), .Z(n809) );
  IV U842 ( .A(n807), .Z(n810) );
  XOR U843 ( .A(n811), .B(n812), .Z(n807) );
  ANDN U844 ( .B(n813), .A(n814), .Z(n811) );
  XNOR U845 ( .A(b[4065]), .B(n812), .Z(n813) );
  XNOR U846 ( .A(b[4065]), .B(n814), .Z(c[4065]) );
  XNOR U847 ( .A(a[4065]), .B(n815), .Z(n814) );
  IV U848 ( .A(n812), .Z(n815) );
  XOR U849 ( .A(n816), .B(n817), .Z(n812) );
  ANDN U850 ( .B(n818), .A(n819), .Z(n816) );
  XNOR U851 ( .A(b[4064]), .B(n817), .Z(n818) );
  XNOR U852 ( .A(b[4064]), .B(n819), .Z(c[4064]) );
  XNOR U853 ( .A(a[4064]), .B(n820), .Z(n819) );
  IV U854 ( .A(n817), .Z(n820) );
  XOR U855 ( .A(n821), .B(n822), .Z(n817) );
  ANDN U856 ( .B(n823), .A(n824), .Z(n821) );
  XNOR U857 ( .A(b[4063]), .B(n822), .Z(n823) );
  XNOR U858 ( .A(b[4063]), .B(n824), .Z(c[4063]) );
  XNOR U859 ( .A(a[4063]), .B(n825), .Z(n824) );
  IV U860 ( .A(n822), .Z(n825) );
  XOR U861 ( .A(n826), .B(n827), .Z(n822) );
  ANDN U862 ( .B(n828), .A(n829), .Z(n826) );
  XNOR U863 ( .A(b[4062]), .B(n827), .Z(n828) );
  XNOR U864 ( .A(b[4062]), .B(n829), .Z(c[4062]) );
  XNOR U865 ( .A(a[4062]), .B(n830), .Z(n829) );
  IV U866 ( .A(n827), .Z(n830) );
  XOR U867 ( .A(n831), .B(n832), .Z(n827) );
  ANDN U868 ( .B(n833), .A(n834), .Z(n831) );
  XNOR U869 ( .A(b[4061]), .B(n832), .Z(n833) );
  XNOR U870 ( .A(b[4061]), .B(n834), .Z(c[4061]) );
  XNOR U871 ( .A(a[4061]), .B(n835), .Z(n834) );
  IV U872 ( .A(n832), .Z(n835) );
  XOR U873 ( .A(n836), .B(n837), .Z(n832) );
  ANDN U874 ( .B(n838), .A(n839), .Z(n836) );
  XNOR U875 ( .A(b[4060]), .B(n837), .Z(n838) );
  XNOR U876 ( .A(b[4060]), .B(n839), .Z(c[4060]) );
  XNOR U877 ( .A(a[4060]), .B(n840), .Z(n839) );
  IV U878 ( .A(n837), .Z(n840) );
  XOR U879 ( .A(n841), .B(n842), .Z(n837) );
  ANDN U880 ( .B(n843), .A(n844), .Z(n841) );
  XNOR U881 ( .A(b[4059]), .B(n842), .Z(n843) );
  XNOR U882 ( .A(b[405]), .B(n845), .Z(c[405]) );
  XNOR U883 ( .A(b[4059]), .B(n844), .Z(c[4059]) );
  XNOR U884 ( .A(a[4059]), .B(n846), .Z(n844) );
  IV U885 ( .A(n842), .Z(n846) );
  XOR U886 ( .A(n847), .B(n848), .Z(n842) );
  ANDN U887 ( .B(n849), .A(n850), .Z(n847) );
  XNOR U888 ( .A(b[4058]), .B(n848), .Z(n849) );
  XNOR U889 ( .A(b[4058]), .B(n850), .Z(c[4058]) );
  XNOR U890 ( .A(a[4058]), .B(n851), .Z(n850) );
  IV U891 ( .A(n848), .Z(n851) );
  XOR U892 ( .A(n852), .B(n853), .Z(n848) );
  ANDN U893 ( .B(n854), .A(n855), .Z(n852) );
  XNOR U894 ( .A(b[4057]), .B(n853), .Z(n854) );
  XNOR U895 ( .A(b[4057]), .B(n855), .Z(c[4057]) );
  XNOR U896 ( .A(a[4057]), .B(n856), .Z(n855) );
  IV U897 ( .A(n853), .Z(n856) );
  XOR U898 ( .A(n857), .B(n858), .Z(n853) );
  ANDN U899 ( .B(n859), .A(n860), .Z(n857) );
  XNOR U900 ( .A(b[4056]), .B(n858), .Z(n859) );
  XNOR U901 ( .A(b[4056]), .B(n860), .Z(c[4056]) );
  XNOR U902 ( .A(a[4056]), .B(n861), .Z(n860) );
  IV U903 ( .A(n858), .Z(n861) );
  XOR U904 ( .A(n862), .B(n863), .Z(n858) );
  ANDN U905 ( .B(n864), .A(n865), .Z(n862) );
  XNOR U906 ( .A(b[4055]), .B(n863), .Z(n864) );
  XNOR U907 ( .A(b[4055]), .B(n865), .Z(c[4055]) );
  XNOR U908 ( .A(a[4055]), .B(n866), .Z(n865) );
  IV U909 ( .A(n863), .Z(n866) );
  XOR U910 ( .A(n867), .B(n868), .Z(n863) );
  ANDN U911 ( .B(n869), .A(n870), .Z(n867) );
  XNOR U912 ( .A(b[4054]), .B(n868), .Z(n869) );
  XNOR U913 ( .A(b[4054]), .B(n870), .Z(c[4054]) );
  XNOR U914 ( .A(a[4054]), .B(n871), .Z(n870) );
  IV U915 ( .A(n868), .Z(n871) );
  XOR U916 ( .A(n872), .B(n873), .Z(n868) );
  ANDN U917 ( .B(n874), .A(n875), .Z(n872) );
  XNOR U918 ( .A(b[4053]), .B(n873), .Z(n874) );
  XNOR U919 ( .A(b[4053]), .B(n875), .Z(c[4053]) );
  XNOR U920 ( .A(a[4053]), .B(n876), .Z(n875) );
  IV U921 ( .A(n873), .Z(n876) );
  XOR U922 ( .A(n877), .B(n878), .Z(n873) );
  ANDN U923 ( .B(n879), .A(n880), .Z(n877) );
  XNOR U924 ( .A(b[4052]), .B(n878), .Z(n879) );
  XNOR U925 ( .A(b[4052]), .B(n880), .Z(c[4052]) );
  XNOR U926 ( .A(a[4052]), .B(n881), .Z(n880) );
  IV U927 ( .A(n878), .Z(n881) );
  XOR U928 ( .A(n882), .B(n883), .Z(n878) );
  ANDN U929 ( .B(n884), .A(n885), .Z(n882) );
  XNOR U930 ( .A(b[4051]), .B(n883), .Z(n884) );
  XNOR U931 ( .A(b[4051]), .B(n885), .Z(c[4051]) );
  XNOR U932 ( .A(a[4051]), .B(n886), .Z(n885) );
  IV U933 ( .A(n883), .Z(n886) );
  XOR U934 ( .A(n887), .B(n888), .Z(n883) );
  ANDN U935 ( .B(n889), .A(n890), .Z(n887) );
  XNOR U936 ( .A(b[4050]), .B(n888), .Z(n889) );
  XNOR U937 ( .A(b[4050]), .B(n890), .Z(c[4050]) );
  XNOR U938 ( .A(a[4050]), .B(n891), .Z(n890) );
  IV U939 ( .A(n888), .Z(n891) );
  XOR U940 ( .A(n892), .B(n893), .Z(n888) );
  ANDN U941 ( .B(n894), .A(n895), .Z(n892) );
  XNOR U942 ( .A(b[4049]), .B(n893), .Z(n894) );
  XNOR U943 ( .A(b[404]), .B(n896), .Z(c[404]) );
  XNOR U944 ( .A(b[4049]), .B(n895), .Z(c[4049]) );
  XNOR U945 ( .A(a[4049]), .B(n897), .Z(n895) );
  IV U946 ( .A(n893), .Z(n897) );
  XOR U947 ( .A(n898), .B(n899), .Z(n893) );
  ANDN U948 ( .B(n900), .A(n901), .Z(n898) );
  XNOR U949 ( .A(b[4048]), .B(n899), .Z(n900) );
  XNOR U950 ( .A(b[4048]), .B(n901), .Z(c[4048]) );
  XNOR U951 ( .A(a[4048]), .B(n902), .Z(n901) );
  IV U952 ( .A(n899), .Z(n902) );
  XOR U953 ( .A(n903), .B(n904), .Z(n899) );
  ANDN U954 ( .B(n905), .A(n906), .Z(n903) );
  XNOR U955 ( .A(b[4047]), .B(n904), .Z(n905) );
  XNOR U956 ( .A(b[4047]), .B(n906), .Z(c[4047]) );
  XNOR U957 ( .A(a[4047]), .B(n907), .Z(n906) );
  IV U958 ( .A(n904), .Z(n907) );
  XOR U959 ( .A(n908), .B(n909), .Z(n904) );
  ANDN U960 ( .B(n910), .A(n911), .Z(n908) );
  XNOR U961 ( .A(b[4046]), .B(n909), .Z(n910) );
  XNOR U962 ( .A(b[4046]), .B(n911), .Z(c[4046]) );
  XNOR U963 ( .A(a[4046]), .B(n912), .Z(n911) );
  IV U964 ( .A(n909), .Z(n912) );
  XOR U965 ( .A(n913), .B(n914), .Z(n909) );
  ANDN U966 ( .B(n915), .A(n916), .Z(n913) );
  XNOR U967 ( .A(b[4045]), .B(n914), .Z(n915) );
  XNOR U968 ( .A(b[4045]), .B(n916), .Z(c[4045]) );
  XNOR U969 ( .A(a[4045]), .B(n917), .Z(n916) );
  IV U970 ( .A(n914), .Z(n917) );
  XOR U971 ( .A(n918), .B(n919), .Z(n914) );
  ANDN U972 ( .B(n920), .A(n921), .Z(n918) );
  XNOR U973 ( .A(b[4044]), .B(n919), .Z(n920) );
  XNOR U974 ( .A(b[4044]), .B(n921), .Z(c[4044]) );
  XNOR U975 ( .A(a[4044]), .B(n922), .Z(n921) );
  IV U976 ( .A(n919), .Z(n922) );
  XOR U977 ( .A(n923), .B(n924), .Z(n919) );
  ANDN U978 ( .B(n925), .A(n926), .Z(n923) );
  XNOR U979 ( .A(b[4043]), .B(n924), .Z(n925) );
  XNOR U980 ( .A(b[4043]), .B(n926), .Z(c[4043]) );
  XNOR U981 ( .A(a[4043]), .B(n927), .Z(n926) );
  IV U982 ( .A(n924), .Z(n927) );
  XOR U983 ( .A(n928), .B(n929), .Z(n924) );
  ANDN U984 ( .B(n930), .A(n931), .Z(n928) );
  XNOR U985 ( .A(b[4042]), .B(n929), .Z(n930) );
  XNOR U986 ( .A(b[4042]), .B(n931), .Z(c[4042]) );
  XNOR U987 ( .A(a[4042]), .B(n932), .Z(n931) );
  IV U988 ( .A(n929), .Z(n932) );
  XOR U989 ( .A(n933), .B(n934), .Z(n929) );
  ANDN U990 ( .B(n935), .A(n936), .Z(n933) );
  XNOR U991 ( .A(b[4041]), .B(n934), .Z(n935) );
  XNOR U992 ( .A(b[4041]), .B(n936), .Z(c[4041]) );
  XNOR U993 ( .A(a[4041]), .B(n937), .Z(n936) );
  IV U994 ( .A(n934), .Z(n937) );
  XOR U995 ( .A(n938), .B(n939), .Z(n934) );
  ANDN U996 ( .B(n940), .A(n941), .Z(n938) );
  XNOR U997 ( .A(b[4040]), .B(n939), .Z(n940) );
  XNOR U998 ( .A(b[4040]), .B(n941), .Z(c[4040]) );
  XNOR U999 ( .A(a[4040]), .B(n942), .Z(n941) );
  IV U1000 ( .A(n939), .Z(n942) );
  XOR U1001 ( .A(n943), .B(n944), .Z(n939) );
  ANDN U1002 ( .B(n945), .A(n946), .Z(n943) );
  XNOR U1003 ( .A(b[4039]), .B(n944), .Z(n945) );
  XNOR U1004 ( .A(b[403]), .B(n947), .Z(c[403]) );
  XNOR U1005 ( .A(b[4039]), .B(n946), .Z(c[4039]) );
  XNOR U1006 ( .A(a[4039]), .B(n948), .Z(n946) );
  IV U1007 ( .A(n944), .Z(n948) );
  XOR U1008 ( .A(n949), .B(n950), .Z(n944) );
  ANDN U1009 ( .B(n951), .A(n952), .Z(n949) );
  XNOR U1010 ( .A(b[4038]), .B(n950), .Z(n951) );
  XNOR U1011 ( .A(b[4038]), .B(n952), .Z(c[4038]) );
  XNOR U1012 ( .A(a[4038]), .B(n953), .Z(n952) );
  IV U1013 ( .A(n950), .Z(n953) );
  XOR U1014 ( .A(n954), .B(n955), .Z(n950) );
  ANDN U1015 ( .B(n956), .A(n957), .Z(n954) );
  XNOR U1016 ( .A(b[4037]), .B(n955), .Z(n956) );
  XNOR U1017 ( .A(b[4037]), .B(n957), .Z(c[4037]) );
  XNOR U1018 ( .A(a[4037]), .B(n958), .Z(n957) );
  IV U1019 ( .A(n955), .Z(n958) );
  XOR U1020 ( .A(n959), .B(n960), .Z(n955) );
  ANDN U1021 ( .B(n961), .A(n962), .Z(n959) );
  XNOR U1022 ( .A(b[4036]), .B(n960), .Z(n961) );
  XNOR U1023 ( .A(b[4036]), .B(n962), .Z(c[4036]) );
  XNOR U1024 ( .A(a[4036]), .B(n963), .Z(n962) );
  IV U1025 ( .A(n960), .Z(n963) );
  XOR U1026 ( .A(n964), .B(n965), .Z(n960) );
  ANDN U1027 ( .B(n966), .A(n967), .Z(n964) );
  XNOR U1028 ( .A(b[4035]), .B(n965), .Z(n966) );
  XNOR U1029 ( .A(b[4035]), .B(n967), .Z(c[4035]) );
  XNOR U1030 ( .A(a[4035]), .B(n968), .Z(n967) );
  IV U1031 ( .A(n965), .Z(n968) );
  XOR U1032 ( .A(n969), .B(n970), .Z(n965) );
  ANDN U1033 ( .B(n971), .A(n972), .Z(n969) );
  XNOR U1034 ( .A(b[4034]), .B(n970), .Z(n971) );
  XNOR U1035 ( .A(b[4034]), .B(n972), .Z(c[4034]) );
  XNOR U1036 ( .A(a[4034]), .B(n973), .Z(n972) );
  IV U1037 ( .A(n970), .Z(n973) );
  XOR U1038 ( .A(n974), .B(n975), .Z(n970) );
  ANDN U1039 ( .B(n976), .A(n977), .Z(n974) );
  XNOR U1040 ( .A(b[4033]), .B(n975), .Z(n976) );
  XNOR U1041 ( .A(b[4033]), .B(n977), .Z(c[4033]) );
  XNOR U1042 ( .A(a[4033]), .B(n978), .Z(n977) );
  IV U1043 ( .A(n975), .Z(n978) );
  XOR U1044 ( .A(n979), .B(n980), .Z(n975) );
  ANDN U1045 ( .B(n981), .A(n982), .Z(n979) );
  XNOR U1046 ( .A(b[4032]), .B(n980), .Z(n981) );
  XNOR U1047 ( .A(b[4032]), .B(n982), .Z(c[4032]) );
  XNOR U1048 ( .A(a[4032]), .B(n983), .Z(n982) );
  IV U1049 ( .A(n980), .Z(n983) );
  XOR U1050 ( .A(n984), .B(n985), .Z(n980) );
  ANDN U1051 ( .B(n986), .A(n987), .Z(n984) );
  XNOR U1052 ( .A(b[4031]), .B(n985), .Z(n986) );
  XNOR U1053 ( .A(b[4031]), .B(n987), .Z(c[4031]) );
  XNOR U1054 ( .A(a[4031]), .B(n988), .Z(n987) );
  IV U1055 ( .A(n985), .Z(n988) );
  XOR U1056 ( .A(n989), .B(n990), .Z(n985) );
  ANDN U1057 ( .B(n991), .A(n992), .Z(n989) );
  XNOR U1058 ( .A(b[4030]), .B(n990), .Z(n991) );
  XNOR U1059 ( .A(b[4030]), .B(n992), .Z(c[4030]) );
  XNOR U1060 ( .A(a[4030]), .B(n993), .Z(n992) );
  IV U1061 ( .A(n990), .Z(n993) );
  XOR U1062 ( .A(n994), .B(n995), .Z(n990) );
  ANDN U1063 ( .B(n996), .A(n997), .Z(n994) );
  XNOR U1064 ( .A(b[4029]), .B(n995), .Z(n996) );
  XNOR U1065 ( .A(b[402]), .B(n998), .Z(c[402]) );
  XNOR U1066 ( .A(b[4029]), .B(n997), .Z(c[4029]) );
  XNOR U1067 ( .A(a[4029]), .B(n999), .Z(n997) );
  IV U1068 ( .A(n995), .Z(n999) );
  XOR U1069 ( .A(n1000), .B(n1001), .Z(n995) );
  ANDN U1070 ( .B(n1002), .A(n1003), .Z(n1000) );
  XNOR U1071 ( .A(b[4028]), .B(n1001), .Z(n1002) );
  XNOR U1072 ( .A(b[4028]), .B(n1003), .Z(c[4028]) );
  XNOR U1073 ( .A(a[4028]), .B(n1004), .Z(n1003) );
  IV U1074 ( .A(n1001), .Z(n1004) );
  XOR U1075 ( .A(n1005), .B(n1006), .Z(n1001) );
  ANDN U1076 ( .B(n1007), .A(n1008), .Z(n1005) );
  XNOR U1077 ( .A(b[4027]), .B(n1006), .Z(n1007) );
  XNOR U1078 ( .A(b[4027]), .B(n1008), .Z(c[4027]) );
  XNOR U1079 ( .A(a[4027]), .B(n1009), .Z(n1008) );
  IV U1080 ( .A(n1006), .Z(n1009) );
  XOR U1081 ( .A(n1010), .B(n1011), .Z(n1006) );
  ANDN U1082 ( .B(n1012), .A(n1013), .Z(n1010) );
  XNOR U1083 ( .A(b[4026]), .B(n1011), .Z(n1012) );
  XNOR U1084 ( .A(b[4026]), .B(n1013), .Z(c[4026]) );
  XNOR U1085 ( .A(a[4026]), .B(n1014), .Z(n1013) );
  IV U1086 ( .A(n1011), .Z(n1014) );
  XOR U1087 ( .A(n1015), .B(n1016), .Z(n1011) );
  ANDN U1088 ( .B(n1017), .A(n1018), .Z(n1015) );
  XNOR U1089 ( .A(b[4025]), .B(n1016), .Z(n1017) );
  XNOR U1090 ( .A(b[4025]), .B(n1018), .Z(c[4025]) );
  XNOR U1091 ( .A(a[4025]), .B(n1019), .Z(n1018) );
  IV U1092 ( .A(n1016), .Z(n1019) );
  XOR U1093 ( .A(n1020), .B(n1021), .Z(n1016) );
  ANDN U1094 ( .B(n1022), .A(n1023), .Z(n1020) );
  XNOR U1095 ( .A(b[4024]), .B(n1021), .Z(n1022) );
  XNOR U1096 ( .A(b[4024]), .B(n1023), .Z(c[4024]) );
  XNOR U1097 ( .A(a[4024]), .B(n1024), .Z(n1023) );
  IV U1098 ( .A(n1021), .Z(n1024) );
  XOR U1099 ( .A(n1025), .B(n1026), .Z(n1021) );
  ANDN U1100 ( .B(n1027), .A(n1028), .Z(n1025) );
  XNOR U1101 ( .A(b[4023]), .B(n1026), .Z(n1027) );
  XNOR U1102 ( .A(b[4023]), .B(n1028), .Z(c[4023]) );
  XNOR U1103 ( .A(a[4023]), .B(n1029), .Z(n1028) );
  IV U1104 ( .A(n1026), .Z(n1029) );
  XOR U1105 ( .A(n1030), .B(n1031), .Z(n1026) );
  ANDN U1106 ( .B(n1032), .A(n1033), .Z(n1030) );
  XNOR U1107 ( .A(b[4022]), .B(n1031), .Z(n1032) );
  XNOR U1108 ( .A(b[4022]), .B(n1033), .Z(c[4022]) );
  XNOR U1109 ( .A(a[4022]), .B(n1034), .Z(n1033) );
  IV U1110 ( .A(n1031), .Z(n1034) );
  XOR U1111 ( .A(n1035), .B(n1036), .Z(n1031) );
  ANDN U1112 ( .B(n1037), .A(n1038), .Z(n1035) );
  XNOR U1113 ( .A(b[4021]), .B(n1036), .Z(n1037) );
  XNOR U1114 ( .A(b[4021]), .B(n1038), .Z(c[4021]) );
  XNOR U1115 ( .A(a[4021]), .B(n1039), .Z(n1038) );
  IV U1116 ( .A(n1036), .Z(n1039) );
  XOR U1117 ( .A(n1040), .B(n1041), .Z(n1036) );
  ANDN U1118 ( .B(n1042), .A(n1043), .Z(n1040) );
  XNOR U1119 ( .A(b[4020]), .B(n1041), .Z(n1042) );
  XNOR U1120 ( .A(b[4020]), .B(n1043), .Z(c[4020]) );
  XNOR U1121 ( .A(a[4020]), .B(n1044), .Z(n1043) );
  IV U1122 ( .A(n1041), .Z(n1044) );
  XOR U1123 ( .A(n1045), .B(n1046), .Z(n1041) );
  ANDN U1124 ( .B(n1047), .A(n1048), .Z(n1045) );
  XNOR U1125 ( .A(b[4019]), .B(n1046), .Z(n1047) );
  XNOR U1126 ( .A(b[401]), .B(n1049), .Z(c[401]) );
  XNOR U1127 ( .A(b[4019]), .B(n1048), .Z(c[4019]) );
  XNOR U1128 ( .A(a[4019]), .B(n1050), .Z(n1048) );
  IV U1129 ( .A(n1046), .Z(n1050) );
  XOR U1130 ( .A(n1051), .B(n1052), .Z(n1046) );
  ANDN U1131 ( .B(n1053), .A(n1054), .Z(n1051) );
  XNOR U1132 ( .A(b[4018]), .B(n1052), .Z(n1053) );
  XNOR U1133 ( .A(b[4018]), .B(n1054), .Z(c[4018]) );
  XNOR U1134 ( .A(a[4018]), .B(n1055), .Z(n1054) );
  IV U1135 ( .A(n1052), .Z(n1055) );
  XOR U1136 ( .A(n1056), .B(n1057), .Z(n1052) );
  ANDN U1137 ( .B(n1058), .A(n1059), .Z(n1056) );
  XNOR U1138 ( .A(b[4017]), .B(n1057), .Z(n1058) );
  XNOR U1139 ( .A(b[4017]), .B(n1059), .Z(c[4017]) );
  XNOR U1140 ( .A(a[4017]), .B(n1060), .Z(n1059) );
  IV U1141 ( .A(n1057), .Z(n1060) );
  XOR U1142 ( .A(n1061), .B(n1062), .Z(n1057) );
  ANDN U1143 ( .B(n1063), .A(n1064), .Z(n1061) );
  XNOR U1144 ( .A(b[4016]), .B(n1062), .Z(n1063) );
  XNOR U1145 ( .A(b[4016]), .B(n1064), .Z(c[4016]) );
  XNOR U1146 ( .A(a[4016]), .B(n1065), .Z(n1064) );
  IV U1147 ( .A(n1062), .Z(n1065) );
  XOR U1148 ( .A(n1066), .B(n1067), .Z(n1062) );
  ANDN U1149 ( .B(n1068), .A(n1069), .Z(n1066) );
  XNOR U1150 ( .A(b[4015]), .B(n1067), .Z(n1068) );
  XNOR U1151 ( .A(b[4015]), .B(n1069), .Z(c[4015]) );
  XNOR U1152 ( .A(a[4015]), .B(n1070), .Z(n1069) );
  IV U1153 ( .A(n1067), .Z(n1070) );
  XOR U1154 ( .A(n1071), .B(n1072), .Z(n1067) );
  ANDN U1155 ( .B(n1073), .A(n1074), .Z(n1071) );
  XNOR U1156 ( .A(b[4014]), .B(n1072), .Z(n1073) );
  XNOR U1157 ( .A(b[4014]), .B(n1074), .Z(c[4014]) );
  XNOR U1158 ( .A(a[4014]), .B(n1075), .Z(n1074) );
  IV U1159 ( .A(n1072), .Z(n1075) );
  XOR U1160 ( .A(n1076), .B(n1077), .Z(n1072) );
  ANDN U1161 ( .B(n1078), .A(n1079), .Z(n1076) );
  XNOR U1162 ( .A(b[4013]), .B(n1077), .Z(n1078) );
  XNOR U1163 ( .A(b[4013]), .B(n1079), .Z(c[4013]) );
  XNOR U1164 ( .A(a[4013]), .B(n1080), .Z(n1079) );
  IV U1165 ( .A(n1077), .Z(n1080) );
  XOR U1166 ( .A(n1081), .B(n1082), .Z(n1077) );
  ANDN U1167 ( .B(n1083), .A(n1084), .Z(n1081) );
  XNOR U1168 ( .A(b[4012]), .B(n1082), .Z(n1083) );
  XNOR U1169 ( .A(b[4012]), .B(n1084), .Z(c[4012]) );
  XNOR U1170 ( .A(a[4012]), .B(n1085), .Z(n1084) );
  IV U1171 ( .A(n1082), .Z(n1085) );
  XOR U1172 ( .A(n1086), .B(n1087), .Z(n1082) );
  ANDN U1173 ( .B(n1088), .A(n1089), .Z(n1086) );
  XNOR U1174 ( .A(b[4011]), .B(n1087), .Z(n1088) );
  XNOR U1175 ( .A(b[4011]), .B(n1089), .Z(c[4011]) );
  XNOR U1176 ( .A(a[4011]), .B(n1090), .Z(n1089) );
  IV U1177 ( .A(n1087), .Z(n1090) );
  XOR U1178 ( .A(n1091), .B(n1092), .Z(n1087) );
  ANDN U1179 ( .B(n1093), .A(n1094), .Z(n1091) );
  XNOR U1180 ( .A(b[4010]), .B(n1092), .Z(n1093) );
  XNOR U1181 ( .A(b[4010]), .B(n1094), .Z(c[4010]) );
  XNOR U1182 ( .A(a[4010]), .B(n1095), .Z(n1094) );
  IV U1183 ( .A(n1092), .Z(n1095) );
  XOR U1184 ( .A(n1096), .B(n1097), .Z(n1092) );
  ANDN U1185 ( .B(n1098), .A(n1099), .Z(n1096) );
  XNOR U1186 ( .A(b[4009]), .B(n1097), .Z(n1098) );
  XNOR U1187 ( .A(b[400]), .B(n1100), .Z(c[400]) );
  XNOR U1188 ( .A(b[4009]), .B(n1099), .Z(c[4009]) );
  XNOR U1189 ( .A(a[4009]), .B(n1101), .Z(n1099) );
  IV U1190 ( .A(n1097), .Z(n1101) );
  XOR U1191 ( .A(n1102), .B(n1103), .Z(n1097) );
  ANDN U1192 ( .B(n1104), .A(n1105), .Z(n1102) );
  XNOR U1193 ( .A(b[4008]), .B(n1103), .Z(n1104) );
  XNOR U1194 ( .A(b[4008]), .B(n1105), .Z(c[4008]) );
  XNOR U1195 ( .A(a[4008]), .B(n1106), .Z(n1105) );
  IV U1196 ( .A(n1103), .Z(n1106) );
  XOR U1197 ( .A(n1107), .B(n1108), .Z(n1103) );
  ANDN U1198 ( .B(n1109), .A(n1110), .Z(n1107) );
  XNOR U1199 ( .A(b[4007]), .B(n1108), .Z(n1109) );
  XNOR U1200 ( .A(b[4007]), .B(n1110), .Z(c[4007]) );
  XNOR U1201 ( .A(a[4007]), .B(n1111), .Z(n1110) );
  IV U1202 ( .A(n1108), .Z(n1111) );
  XOR U1203 ( .A(n1112), .B(n1113), .Z(n1108) );
  ANDN U1204 ( .B(n1114), .A(n1115), .Z(n1112) );
  XNOR U1205 ( .A(b[4006]), .B(n1113), .Z(n1114) );
  XNOR U1206 ( .A(b[4006]), .B(n1115), .Z(c[4006]) );
  XNOR U1207 ( .A(a[4006]), .B(n1116), .Z(n1115) );
  IV U1208 ( .A(n1113), .Z(n1116) );
  XOR U1209 ( .A(n1117), .B(n1118), .Z(n1113) );
  ANDN U1210 ( .B(n1119), .A(n1120), .Z(n1117) );
  XNOR U1211 ( .A(b[4005]), .B(n1118), .Z(n1119) );
  XNOR U1212 ( .A(b[4005]), .B(n1120), .Z(c[4005]) );
  XNOR U1213 ( .A(a[4005]), .B(n1121), .Z(n1120) );
  IV U1214 ( .A(n1118), .Z(n1121) );
  XOR U1215 ( .A(n1122), .B(n1123), .Z(n1118) );
  ANDN U1216 ( .B(n1124), .A(n1125), .Z(n1122) );
  XNOR U1217 ( .A(b[4004]), .B(n1123), .Z(n1124) );
  XNOR U1218 ( .A(b[4004]), .B(n1125), .Z(c[4004]) );
  XNOR U1219 ( .A(a[4004]), .B(n1126), .Z(n1125) );
  IV U1220 ( .A(n1123), .Z(n1126) );
  XOR U1221 ( .A(n1127), .B(n1128), .Z(n1123) );
  ANDN U1222 ( .B(n1129), .A(n1130), .Z(n1127) );
  XNOR U1223 ( .A(b[4003]), .B(n1128), .Z(n1129) );
  XNOR U1224 ( .A(b[4003]), .B(n1130), .Z(c[4003]) );
  XNOR U1225 ( .A(a[4003]), .B(n1131), .Z(n1130) );
  IV U1226 ( .A(n1128), .Z(n1131) );
  XOR U1227 ( .A(n1132), .B(n1133), .Z(n1128) );
  ANDN U1228 ( .B(n1134), .A(n1135), .Z(n1132) );
  XNOR U1229 ( .A(b[4002]), .B(n1133), .Z(n1134) );
  XNOR U1230 ( .A(b[4002]), .B(n1135), .Z(c[4002]) );
  XNOR U1231 ( .A(a[4002]), .B(n1136), .Z(n1135) );
  IV U1232 ( .A(n1133), .Z(n1136) );
  XOR U1233 ( .A(n1137), .B(n1138), .Z(n1133) );
  ANDN U1234 ( .B(n1139), .A(n1140), .Z(n1137) );
  XNOR U1235 ( .A(b[4001]), .B(n1138), .Z(n1139) );
  XNOR U1236 ( .A(b[4001]), .B(n1140), .Z(c[4001]) );
  XNOR U1237 ( .A(a[4001]), .B(n1141), .Z(n1140) );
  IV U1238 ( .A(n1138), .Z(n1141) );
  XOR U1239 ( .A(n1142), .B(n1143), .Z(n1138) );
  ANDN U1240 ( .B(n1144), .A(n1145), .Z(n1142) );
  XNOR U1241 ( .A(b[4000]), .B(n1143), .Z(n1144) );
  XNOR U1242 ( .A(b[4000]), .B(n1145), .Z(c[4000]) );
  XNOR U1243 ( .A(a[4000]), .B(n1146), .Z(n1145) );
  IV U1244 ( .A(n1143), .Z(n1146) );
  XOR U1245 ( .A(n1147), .B(n1148), .Z(n1143) );
  ANDN U1246 ( .B(n1149), .A(n1150), .Z(n1147) );
  XNOR U1247 ( .A(b[3999]), .B(n1148), .Z(n1149) );
  XNOR U1248 ( .A(b[3]), .B(n1151), .Z(c[3]) );
  XNOR U1249 ( .A(b[39]), .B(n1152), .Z(c[39]) );
  XNOR U1250 ( .A(b[399]), .B(n1153), .Z(c[399]) );
  XNOR U1251 ( .A(b[3999]), .B(n1150), .Z(c[3999]) );
  XNOR U1252 ( .A(a[3999]), .B(n1154), .Z(n1150) );
  IV U1253 ( .A(n1148), .Z(n1154) );
  XOR U1254 ( .A(n1155), .B(n1156), .Z(n1148) );
  ANDN U1255 ( .B(n1157), .A(n1158), .Z(n1155) );
  XNOR U1256 ( .A(b[3998]), .B(n1156), .Z(n1157) );
  XNOR U1257 ( .A(b[3998]), .B(n1158), .Z(c[3998]) );
  XNOR U1258 ( .A(a[3998]), .B(n1159), .Z(n1158) );
  IV U1259 ( .A(n1156), .Z(n1159) );
  XOR U1260 ( .A(n1160), .B(n1161), .Z(n1156) );
  ANDN U1261 ( .B(n1162), .A(n1163), .Z(n1160) );
  XNOR U1262 ( .A(b[3997]), .B(n1161), .Z(n1162) );
  XNOR U1263 ( .A(b[3997]), .B(n1163), .Z(c[3997]) );
  XNOR U1264 ( .A(a[3997]), .B(n1164), .Z(n1163) );
  IV U1265 ( .A(n1161), .Z(n1164) );
  XOR U1266 ( .A(n1165), .B(n1166), .Z(n1161) );
  ANDN U1267 ( .B(n1167), .A(n1168), .Z(n1165) );
  XNOR U1268 ( .A(b[3996]), .B(n1166), .Z(n1167) );
  XNOR U1269 ( .A(b[3996]), .B(n1168), .Z(c[3996]) );
  XNOR U1270 ( .A(a[3996]), .B(n1169), .Z(n1168) );
  IV U1271 ( .A(n1166), .Z(n1169) );
  XOR U1272 ( .A(n1170), .B(n1171), .Z(n1166) );
  ANDN U1273 ( .B(n1172), .A(n1173), .Z(n1170) );
  XNOR U1274 ( .A(b[3995]), .B(n1171), .Z(n1172) );
  XNOR U1275 ( .A(b[3995]), .B(n1173), .Z(c[3995]) );
  XNOR U1276 ( .A(a[3995]), .B(n1174), .Z(n1173) );
  IV U1277 ( .A(n1171), .Z(n1174) );
  XOR U1278 ( .A(n1175), .B(n1176), .Z(n1171) );
  ANDN U1279 ( .B(n1177), .A(n1178), .Z(n1175) );
  XNOR U1280 ( .A(b[3994]), .B(n1176), .Z(n1177) );
  XNOR U1281 ( .A(b[3994]), .B(n1178), .Z(c[3994]) );
  XNOR U1282 ( .A(a[3994]), .B(n1179), .Z(n1178) );
  IV U1283 ( .A(n1176), .Z(n1179) );
  XOR U1284 ( .A(n1180), .B(n1181), .Z(n1176) );
  ANDN U1285 ( .B(n1182), .A(n1183), .Z(n1180) );
  XNOR U1286 ( .A(b[3993]), .B(n1181), .Z(n1182) );
  XNOR U1287 ( .A(b[3993]), .B(n1183), .Z(c[3993]) );
  XNOR U1288 ( .A(a[3993]), .B(n1184), .Z(n1183) );
  IV U1289 ( .A(n1181), .Z(n1184) );
  XOR U1290 ( .A(n1185), .B(n1186), .Z(n1181) );
  ANDN U1291 ( .B(n1187), .A(n1188), .Z(n1185) );
  XNOR U1292 ( .A(b[3992]), .B(n1186), .Z(n1187) );
  XNOR U1293 ( .A(b[3992]), .B(n1188), .Z(c[3992]) );
  XNOR U1294 ( .A(a[3992]), .B(n1189), .Z(n1188) );
  IV U1295 ( .A(n1186), .Z(n1189) );
  XOR U1296 ( .A(n1190), .B(n1191), .Z(n1186) );
  ANDN U1297 ( .B(n1192), .A(n1193), .Z(n1190) );
  XNOR U1298 ( .A(b[3991]), .B(n1191), .Z(n1192) );
  XNOR U1299 ( .A(b[3991]), .B(n1193), .Z(c[3991]) );
  XNOR U1300 ( .A(a[3991]), .B(n1194), .Z(n1193) );
  IV U1301 ( .A(n1191), .Z(n1194) );
  XOR U1302 ( .A(n1195), .B(n1196), .Z(n1191) );
  ANDN U1303 ( .B(n1197), .A(n1198), .Z(n1195) );
  XNOR U1304 ( .A(b[3990]), .B(n1196), .Z(n1197) );
  XNOR U1305 ( .A(b[3990]), .B(n1198), .Z(c[3990]) );
  XNOR U1306 ( .A(a[3990]), .B(n1199), .Z(n1198) );
  IV U1307 ( .A(n1196), .Z(n1199) );
  XOR U1308 ( .A(n1200), .B(n1201), .Z(n1196) );
  ANDN U1309 ( .B(n1202), .A(n1203), .Z(n1200) );
  XNOR U1310 ( .A(b[3989]), .B(n1201), .Z(n1202) );
  XNOR U1311 ( .A(b[398]), .B(n1204), .Z(c[398]) );
  XNOR U1312 ( .A(b[3989]), .B(n1203), .Z(c[3989]) );
  XNOR U1313 ( .A(a[3989]), .B(n1205), .Z(n1203) );
  IV U1314 ( .A(n1201), .Z(n1205) );
  XOR U1315 ( .A(n1206), .B(n1207), .Z(n1201) );
  ANDN U1316 ( .B(n1208), .A(n1209), .Z(n1206) );
  XNOR U1317 ( .A(b[3988]), .B(n1207), .Z(n1208) );
  XNOR U1318 ( .A(b[3988]), .B(n1209), .Z(c[3988]) );
  XNOR U1319 ( .A(a[3988]), .B(n1210), .Z(n1209) );
  IV U1320 ( .A(n1207), .Z(n1210) );
  XOR U1321 ( .A(n1211), .B(n1212), .Z(n1207) );
  ANDN U1322 ( .B(n1213), .A(n1214), .Z(n1211) );
  XNOR U1323 ( .A(b[3987]), .B(n1212), .Z(n1213) );
  XNOR U1324 ( .A(b[3987]), .B(n1214), .Z(c[3987]) );
  XNOR U1325 ( .A(a[3987]), .B(n1215), .Z(n1214) );
  IV U1326 ( .A(n1212), .Z(n1215) );
  XOR U1327 ( .A(n1216), .B(n1217), .Z(n1212) );
  ANDN U1328 ( .B(n1218), .A(n1219), .Z(n1216) );
  XNOR U1329 ( .A(b[3986]), .B(n1217), .Z(n1218) );
  XNOR U1330 ( .A(b[3986]), .B(n1219), .Z(c[3986]) );
  XNOR U1331 ( .A(a[3986]), .B(n1220), .Z(n1219) );
  IV U1332 ( .A(n1217), .Z(n1220) );
  XOR U1333 ( .A(n1221), .B(n1222), .Z(n1217) );
  ANDN U1334 ( .B(n1223), .A(n1224), .Z(n1221) );
  XNOR U1335 ( .A(b[3985]), .B(n1222), .Z(n1223) );
  XNOR U1336 ( .A(b[3985]), .B(n1224), .Z(c[3985]) );
  XNOR U1337 ( .A(a[3985]), .B(n1225), .Z(n1224) );
  IV U1338 ( .A(n1222), .Z(n1225) );
  XOR U1339 ( .A(n1226), .B(n1227), .Z(n1222) );
  ANDN U1340 ( .B(n1228), .A(n1229), .Z(n1226) );
  XNOR U1341 ( .A(b[3984]), .B(n1227), .Z(n1228) );
  XNOR U1342 ( .A(b[3984]), .B(n1229), .Z(c[3984]) );
  XNOR U1343 ( .A(a[3984]), .B(n1230), .Z(n1229) );
  IV U1344 ( .A(n1227), .Z(n1230) );
  XOR U1345 ( .A(n1231), .B(n1232), .Z(n1227) );
  ANDN U1346 ( .B(n1233), .A(n1234), .Z(n1231) );
  XNOR U1347 ( .A(b[3983]), .B(n1232), .Z(n1233) );
  XNOR U1348 ( .A(b[3983]), .B(n1234), .Z(c[3983]) );
  XNOR U1349 ( .A(a[3983]), .B(n1235), .Z(n1234) );
  IV U1350 ( .A(n1232), .Z(n1235) );
  XOR U1351 ( .A(n1236), .B(n1237), .Z(n1232) );
  ANDN U1352 ( .B(n1238), .A(n1239), .Z(n1236) );
  XNOR U1353 ( .A(b[3982]), .B(n1237), .Z(n1238) );
  XNOR U1354 ( .A(b[3982]), .B(n1239), .Z(c[3982]) );
  XNOR U1355 ( .A(a[3982]), .B(n1240), .Z(n1239) );
  IV U1356 ( .A(n1237), .Z(n1240) );
  XOR U1357 ( .A(n1241), .B(n1242), .Z(n1237) );
  ANDN U1358 ( .B(n1243), .A(n1244), .Z(n1241) );
  XNOR U1359 ( .A(b[3981]), .B(n1242), .Z(n1243) );
  XNOR U1360 ( .A(b[3981]), .B(n1244), .Z(c[3981]) );
  XNOR U1361 ( .A(a[3981]), .B(n1245), .Z(n1244) );
  IV U1362 ( .A(n1242), .Z(n1245) );
  XOR U1363 ( .A(n1246), .B(n1247), .Z(n1242) );
  ANDN U1364 ( .B(n1248), .A(n1249), .Z(n1246) );
  XNOR U1365 ( .A(b[3980]), .B(n1247), .Z(n1248) );
  XNOR U1366 ( .A(b[3980]), .B(n1249), .Z(c[3980]) );
  XNOR U1367 ( .A(a[3980]), .B(n1250), .Z(n1249) );
  IV U1368 ( .A(n1247), .Z(n1250) );
  XOR U1369 ( .A(n1251), .B(n1252), .Z(n1247) );
  ANDN U1370 ( .B(n1253), .A(n1254), .Z(n1251) );
  XNOR U1371 ( .A(b[3979]), .B(n1252), .Z(n1253) );
  XNOR U1372 ( .A(b[397]), .B(n1255), .Z(c[397]) );
  XNOR U1373 ( .A(b[3979]), .B(n1254), .Z(c[3979]) );
  XNOR U1374 ( .A(a[3979]), .B(n1256), .Z(n1254) );
  IV U1375 ( .A(n1252), .Z(n1256) );
  XOR U1376 ( .A(n1257), .B(n1258), .Z(n1252) );
  ANDN U1377 ( .B(n1259), .A(n1260), .Z(n1257) );
  XNOR U1378 ( .A(b[3978]), .B(n1258), .Z(n1259) );
  XNOR U1379 ( .A(b[3978]), .B(n1260), .Z(c[3978]) );
  XNOR U1380 ( .A(a[3978]), .B(n1261), .Z(n1260) );
  IV U1381 ( .A(n1258), .Z(n1261) );
  XOR U1382 ( .A(n1262), .B(n1263), .Z(n1258) );
  ANDN U1383 ( .B(n1264), .A(n1265), .Z(n1262) );
  XNOR U1384 ( .A(b[3977]), .B(n1263), .Z(n1264) );
  XNOR U1385 ( .A(b[3977]), .B(n1265), .Z(c[3977]) );
  XNOR U1386 ( .A(a[3977]), .B(n1266), .Z(n1265) );
  IV U1387 ( .A(n1263), .Z(n1266) );
  XOR U1388 ( .A(n1267), .B(n1268), .Z(n1263) );
  ANDN U1389 ( .B(n1269), .A(n1270), .Z(n1267) );
  XNOR U1390 ( .A(b[3976]), .B(n1268), .Z(n1269) );
  XNOR U1391 ( .A(b[3976]), .B(n1270), .Z(c[3976]) );
  XNOR U1392 ( .A(a[3976]), .B(n1271), .Z(n1270) );
  IV U1393 ( .A(n1268), .Z(n1271) );
  XOR U1394 ( .A(n1272), .B(n1273), .Z(n1268) );
  ANDN U1395 ( .B(n1274), .A(n1275), .Z(n1272) );
  XNOR U1396 ( .A(b[3975]), .B(n1273), .Z(n1274) );
  XNOR U1397 ( .A(b[3975]), .B(n1275), .Z(c[3975]) );
  XNOR U1398 ( .A(a[3975]), .B(n1276), .Z(n1275) );
  IV U1399 ( .A(n1273), .Z(n1276) );
  XOR U1400 ( .A(n1277), .B(n1278), .Z(n1273) );
  ANDN U1401 ( .B(n1279), .A(n1280), .Z(n1277) );
  XNOR U1402 ( .A(b[3974]), .B(n1278), .Z(n1279) );
  XNOR U1403 ( .A(b[3974]), .B(n1280), .Z(c[3974]) );
  XNOR U1404 ( .A(a[3974]), .B(n1281), .Z(n1280) );
  IV U1405 ( .A(n1278), .Z(n1281) );
  XOR U1406 ( .A(n1282), .B(n1283), .Z(n1278) );
  ANDN U1407 ( .B(n1284), .A(n1285), .Z(n1282) );
  XNOR U1408 ( .A(b[3973]), .B(n1283), .Z(n1284) );
  XNOR U1409 ( .A(b[3973]), .B(n1285), .Z(c[3973]) );
  XNOR U1410 ( .A(a[3973]), .B(n1286), .Z(n1285) );
  IV U1411 ( .A(n1283), .Z(n1286) );
  XOR U1412 ( .A(n1287), .B(n1288), .Z(n1283) );
  ANDN U1413 ( .B(n1289), .A(n1290), .Z(n1287) );
  XNOR U1414 ( .A(b[3972]), .B(n1288), .Z(n1289) );
  XNOR U1415 ( .A(b[3972]), .B(n1290), .Z(c[3972]) );
  XNOR U1416 ( .A(a[3972]), .B(n1291), .Z(n1290) );
  IV U1417 ( .A(n1288), .Z(n1291) );
  XOR U1418 ( .A(n1292), .B(n1293), .Z(n1288) );
  ANDN U1419 ( .B(n1294), .A(n1295), .Z(n1292) );
  XNOR U1420 ( .A(b[3971]), .B(n1293), .Z(n1294) );
  XNOR U1421 ( .A(b[3971]), .B(n1295), .Z(c[3971]) );
  XNOR U1422 ( .A(a[3971]), .B(n1296), .Z(n1295) );
  IV U1423 ( .A(n1293), .Z(n1296) );
  XOR U1424 ( .A(n1297), .B(n1298), .Z(n1293) );
  ANDN U1425 ( .B(n1299), .A(n1300), .Z(n1297) );
  XNOR U1426 ( .A(b[3970]), .B(n1298), .Z(n1299) );
  XNOR U1427 ( .A(b[3970]), .B(n1300), .Z(c[3970]) );
  XNOR U1428 ( .A(a[3970]), .B(n1301), .Z(n1300) );
  IV U1429 ( .A(n1298), .Z(n1301) );
  XOR U1430 ( .A(n1302), .B(n1303), .Z(n1298) );
  ANDN U1431 ( .B(n1304), .A(n1305), .Z(n1302) );
  XNOR U1432 ( .A(b[3969]), .B(n1303), .Z(n1304) );
  XNOR U1433 ( .A(b[396]), .B(n1306), .Z(c[396]) );
  XNOR U1434 ( .A(b[3969]), .B(n1305), .Z(c[3969]) );
  XNOR U1435 ( .A(a[3969]), .B(n1307), .Z(n1305) );
  IV U1436 ( .A(n1303), .Z(n1307) );
  XOR U1437 ( .A(n1308), .B(n1309), .Z(n1303) );
  ANDN U1438 ( .B(n1310), .A(n1311), .Z(n1308) );
  XNOR U1439 ( .A(b[3968]), .B(n1309), .Z(n1310) );
  XNOR U1440 ( .A(b[3968]), .B(n1311), .Z(c[3968]) );
  XNOR U1441 ( .A(a[3968]), .B(n1312), .Z(n1311) );
  IV U1442 ( .A(n1309), .Z(n1312) );
  XOR U1443 ( .A(n1313), .B(n1314), .Z(n1309) );
  ANDN U1444 ( .B(n1315), .A(n1316), .Z(n1313) );
  XNOR U1445 ( .A(b[3967]), .B(n1314), .Z(n1315) );
  XNOR U1446 ( .A(b[3967]), .B(n1316), .Z(c[3967]) );
  XNOR U1447 ( .A(a[3967]), .B(n1317), .Z(n1316) );
  IV U1448 ( .A(n1314), .Z(n1317) );
  XOR U1449 ( .A(n1318), .B(n1319), .Z(n1314) );
  ANDN U1450 ( .B(n1320), .A(n1321), .Z(n1318) );
  XNOR U1451 ( .A(b[3966]), .B(n1319), .Z(n1320) );
  XNOR U1452 ( .A(b[3966]), .B(n1321), .Z(c[3966]) );
  XNOR U1453 ( .A(a[3966]), .B(n1322), .Z(n1321) );
  IV U1454 ( .A(n1319), .Z(n1322) );
  XOR U1455 ( .A(n1323), .B(n1324), .Z(n1319) );
  ANDN U1456 ( .B(n1325), .A(n1326), .Z(n1323) );
  XNOR U1457 ( .A(b[3965]), .B(n1324), .Z(n1325) );
  XNOR U1458 ( .A(b[3965]), .B(n1326), .Z(c[3965]) );
  XNOR U1459 ( .A(a[3965]), .B(n1327), .Z(n1326) );
  IV U1460 ( .A(n1324), .Z(n1327) );
  XOR U1461 ( .A(n1328), .B(n1329), .Z(n1324) );
  ANDN U1462 ( .B(n1330), .A(n1331), .Z(n1328) );
  XNOR U1463 ( .A(b[3964]), .B(n1329), .Z(n1330) );
  XNOR U1464 ( .A(b[3964]), .B(n1331), .Z(c[3964]) );
  XNOR U1465 ( .A(a[3964]), .B(n1332), .Z(n1331) );
  IV U1466 ( .A(n1329), .Z(n1332) );
  XOR U1467 ( .A(n1333), .B(n1334), .Z(n1329) );
  ANDN U1468 ( .B(n1335), .A(n1336), .Z(n1333) );
  XNOR U1469 ( .A(b[3963]), .B(n1334), .Z(n1335) );
  XNOR U1470 ( .A(b[3963]), .B(n1336), .Z(c[3963]) );
  XNOR U1471 ( .A(a[3963]), .B(n1337), .Z(n1336) );
  IV U1472 ( .A(n1334), .Z(n1337) );
  XOR U1473 ( .A(n1338), .B(n1339), .Z(n1334) );
  ANDN U1474 ( .B(n1340), .A(n1341), .Z(n1338) );
  XNOR U1475 ( .A(b[3962]), .B(n1339), .Z(n1340) );
  XNOR U1476 ( .A(b[3962]), .B(n1341), .Z(c[3962]) );
  XNOR U1477 ( .A(a[3962]), .B(n1342), .Z(n1341) );
  IV U1478 ( .A(n1339), .Z(n1342) );
  XOR U1479 ( .A(n1343), .B(n1344), .Z(n1339) );
  ANDN U1480 ( .B(n1345), .A(n1346), .Z(n1343) );
  XNOR U1481 ( .A(b[3961]), .B(n1344), .Z(n1345) );
  XNOR U1482 ( .A(b[3961]), .B(n1346), .Z(c[3961]) );
  XNOR U1483 ( .A(a[3961]), .B(n1347), .Z(n1346) );
  IV U1484 ( .A(n1344), .Z(n1347) );
  XOR U1485 ( .A(n1348), .B(n1349), .Z(n1344) );
  ANDN U1486 ( .B(n1350), .A(n1351), .Z(n1348) );
  XNOR U1487 ( .A(b[3960]), .B(n1349), .Z(n1350) );
  XNOR U1488 ( .A(b[3960]), .B(n1351), .Z(c[3960]) );
  XNOR U1489 ( .A(a[3960]), .B(n1352), .Z(n1351) );
  IV U1490 ( .A(n1349), .Z(n1352) );
  XOR U1491 ( .A(n1353), .B(n1354), .Z(n1349) );
  ANDN U1492 ( .B(n1355), .A(n1356), .Z(n1353) );
  XNOR U1493 ( .A(b[3959]), .B(n1354), .Z(n1355) );
  XNOR U1494 ( .A(b[395]), .B(n1357), .Z(c[395]) );
  XNOR U1495 ( .A(b[3959]), .B(n1356), .Z(c[3959]) );
  XNOR U1496 ( .A(a[3959]), .B(n1358), .Z(n1356) );
  IV U1497 ( .A(n1354), .Z(n1358) );
  XOR U1498 ( .A(n1359), .B(n1360), .Z(n1354) );
  ANDN U1499 ( .B(n1361), .A(n1362), .Z(n1359) );
  XNOR U1500 ( .A(b[3958]), .B(n1360), .Z(n1361) );
  XNOR U1501 ( .A(b[3958]), .B(n1362), .Z(c[3958]) );
  XNOR U1502 ( .A(a[3958]), .B(n1363), .Z(n1362) );
  IV U1503 ( .A(n1360), .Z(n1363) );
  XOR U1504 ( .A(n1364), .B(n1365), .Z(n1360) );
  ANDN U1505 ( .B(n1366), .A(n1367), .Z(n1364) );
  XNOR U1506 ( .A(b[3957]), .B(n1365), .Z(n1366) );
  XNOR U1507 ( .A(b[3957]), .B(n1367), .Z(c[3957]) );
  XNOR U1508 ( .A(a[3957]), .B(n1368), .Z(n1367) );
  IV U1509 ( .A(n1365), .Z(n1368) );
  XOR U1510 ( .A(n1369), .B(n1370), .Z(n1365) );
  ANDN U1511 ( .B(n1371), .A(n1372), .Z(n1369) );
  XNOR U1512 ( .A(b[3956]), .B(n1370), .Z(n1371) );
  XNOR U1513 ( .A(b[3956]), .B(n1372), .Z(c[3956]) );
  XNOR U1514 ( .A(a[3956]), .B(n1373), .Z(n1372) );
  IV U1515 ( .A(n1370), .Z(n1373) );
  XOR U1516 ( .A(n1374), .B(n1375), .Z(n1370) );
  ANDN U1517 ( .B(n1376), .A(n1377), .Z(n1374) );
  XNOR U1518 ( .A(b[3955]), .B(n1375), .Z(n1376) );
  XNOR U1519 ( .A(b[3955]), .B(n1377), .Z(c[3955]) );
  XNOR U1520 ( .A(a[3955]), .B(n1378), .Z(n1377) );
  IV U1521 ( .A(n1375), .Z(n1378) );
  XOR U1522 ( .A(n1379), .B(n1380), .Z(n1375) );
  ANDN U1523 ( .B(n1381), .A(n1382), .Z(n1379) );
  XNOR U1524 ( .A(b[3954]), .B(n1380), .Z(n1381) );
  XNOR U1525 ( .A(b[3954]), .B(n1382), .Z(c[3954]) );
  XNOR U1526 ( .A(a[3954]), .B(n1383), .Z(n1382) );
  IV U1527 ( .A(n1380), .Z(n1383) );
  XOR U1528 ( .A(n1384), .B(n1385), .Z(n1380) );
  ANDN U1529 ( .B(n1386), .A(n1387), .Z(n1384) );
  XNOR U1530 ( .A(b[3953]), .B(n1385), .Z(n1386) );
  XNOR U1531 ( .A(b[3953]), .B(n1387), .Z(c[3953]) );
  XNOR U1532 ( .A(a[3953]), .B(n1388), .Z(n1387) );
  IV U1533 ( .A(n1385), .Z(n1388) );
  XOR U1534 ( .A(n1389), .B(n1390), .Z(n1385) );
  ANDN U1535 ( .B(n1391), .A(n1392), .Z(n1389) );
  XNOR U1536 ( .A(b[3952]), .B(n1390), .Z(n1391) );
  XNOR U1537 ( .A(b[3952]), .B(n1392), .Z(c[3952]) );
  XNOR U1538 ( .A(a[3952]), .B(n1393), .Z(n1392) );
  IV U1539 ( .A(n1390), .Z(n1393) );
  XOR U1540 ( .A(n1394), .B(n1395), .Z(n1390) );
  ANDN U1541 ( .B(n1396), .A(n1397), .Z(n1394) );
  XNOR U1542 ( .A(b[3951]), .B(n1395), .Z(n1396) );
  XNOR U1543 ( .A(b[3951]), .B(n1397), .Z(c[3951]) );
  XNOR U1544 ( .A(a[3951]), .B(n1398), .Z(n1397) );
  IV U1545 ( .A(n1395), .Z(n1398) );
  XOR U1546 ( .A(n1399), .B(n1400), .Z(n1395) );
  ANDN U1547 ( .B(n1401), .A(n1402), .Z(n1399) );
  XNOR U1548 ( .A(b[3950]), .B(n1400), .Z(n1401) );
  XNOR U1549 ( .A(b[3950]), .B(n1402), .Z(c[3950]) );
  XNOR U1550 ( .A(a[3950]), .B(n1403), .Z(n1402) );
  IV U1551 ( .A(n1400), .Z(n1403) );
  XOR U1552 ( .A(n1404), .B(n1405), .Z(n1400) );
  ANDN U1553 ( .B(n1406), .A(n1407), .Z(n1404) );
  XNOR U1554 ( .A(b[3949]), .B(n1405), .Z(n1406) );
  XNOR U1555 ( .A(b[394]), .B(n1408), .Z(c[394]) );
  XNOR U1556 ( .A(b[3949]), .B(n1407), .Z(c[3949]) );
  XNOR U1557 ( .A(a[3949]), .B(n1409), .Z(n1407) );
  IV U1558 ( .A(n1405), .Z(n1409) );
  XOR U1559 ( .A(n1410), .B(n1411), .Z(n1405) );
  ANDN U1560 ( .B(n1412), .A(n1413), .Z(n1410) );
  XNOR U1561 ( .A(b[3948]), .B(n1411), .Z(n1412) );
  XNOR U1562 ( .A(b[3948]), .B(n1413), .Z(c[3948]) );
  XNOR U1563 ( .A(a[3948]), .B(n1414), .Z(n1413) );
  IV U1564 ( .A(n1411), .Z(n1414) );
  XOR U1565 ( .A(n1415), .B(n1416), .Z(n1411) );
  ANDN U1566 ( .B(n1417), .A(n1418), .Z(n1415) );
  XNOR U1567 ( .A(b[3947]), .B(n1416), .Z(n1417) );
  XNOR U1568 ( .A(b[3947]), .B(n1418), .Z(c[3947]) );
  XNOR U1569 ( .A(a[3947]), .B(n1419), .Z(n1418) );
  IV U1570 ( .A(n1416), .Z(n1419) );
  XOR U1571 ( .A(n1420), .B(n1421), .Z(n1416) );
  ANDN U1572 ( .B(n1422), .A(n1423), .Z(n1420) );
  XNOR U1573 ( .A(b[3946]), .B(n1421), .Z(n1422) );
  XNOR U1574 ( .A(b[3946]), .B(n1423), .Z(c[3946]) );
  XNOR U1575 ( .A(a[3946]), .B(n1424), .Z(n1423) );
  IV U1576 ( .A(n1421), .Z(n1424) );
  XOR U1577 ( .A(n1425), .B(n1426), .Z(n1421) );
  ANDN U1578 ( .B(n1427), .A(n1428), .Z(n1425) );
  XNOR U1579 ( .A(b[3945]), .B(n1426), .Z(n1427) );
  XNOR U1580 ( .A(b[3945]), .B(n1428), .Z(c[3945]) );
  XNOR U1581 ( .A(a[3945]), .B(n1429), .Z(n1428) );
  IV U1582 ( .A(n1426), .Z(n1429) );
  XOR U1583 ( .A(n1430), .B(n1431), .Z(n1426) );
  ANDN U1584 ( .B(n1432), .A(n1433), .Z(n1430) );
  XNOR U1585 ( .A(b[3944]), .B(n1431), .Z(n1432) );
  XNOR U1586 ( .A(b[3944]), .B(n1433), .Z(c[3944]) );
  XNOR U1587 ( .A(a[3944]), .B(n1434), .Z(n1433) );
  IV U1588 ( .A(n1431), .Z(n1434) );
  XOR U1589 ( .A(n1435), .B(n1436), .Z(n1431) );
  ANDN U1590 ( .B(n1437), .A(n1438), .Z(n1435) );
  XNOR U1591 ( .A(b[3943]), .B(n1436), .Z(n1437) );
  XNOR U1592 ( .A(b[3943]), .B(n1438), .Z(c[3943]) );
  XNOR U1593 ( .A(a[3943]), .B(n1439), .Z(n1438) );
  IV U1594 ( .A(n1436), .Z(n1439) );
  XOR U1595 ( .A(n1440), .B(n1441), .Z(n1436) );
  ANDN U1596 ( .B(n1442), .A(n1443), .Z(n1440) );
  XNOR U1597 ( .A(b[3942]), .B(n1441), .Z(n1442) );
  XNOR U1598 ( .A(b[3942]), .B(n1443), .Z(c[3942]) );
  XNOR U1599 ( .A(a[3942]), .B(n1444), .Z(n1443) );
  IV U1600 ( .A(n1441), .Z(n1444) );
  XOR U1601 ( .A(n1445), .B(n1446), .Z(n1441) );
  ANDN U1602 ( .B(n1447), .A(n1448), .Z(n1445) );
  XNOR U1603 ( .A(b[3941]), .B(n1446), .Z(n1447) );
  XNOR U1604 ( .A(b[3941]), .B(n1448), .Z(c[3941]) );
  XNOR U1605 ( .A(a[3941]), .B(n1449), .Z(n1448) );
  IV U1606 ( .A(n1446), .Z(n1449) );
  XOR U1607 ( .A(n1450), .B(n1451), .Z(n1446) );
  ANDN U1608 ( .B(n1452), .A(n1453), .Z(n1450) );
  XNOR U1609 ( .A(b[3940]), .B(n1451), .Z(n1452) );
  XNOR U1610 ( .A(b[3940]), .B(n1453), .Z(c[3940]) );
  XNOR U1611 ( .A(a[3940]), .B(n1454), .Z(n1453) );
  IV U1612 ( .A(n1451), .Z(n1454) );
  XOR U1613 ( .A(n1455), .B(n1456), .Z(n1451) );
  ANDN U1614 ( .B(n1457), .A(n1458), .Z(n1455) );
  XNOR U1615 ( .A(b[3939]), .B(n1456), .Z(n1457) );
  XNOR U1616 ( .A(b[393]), .B(n1459), .Z(c[393]) );
  XNOR U1617 ( .A(b[3939]), .B(n1458), .Z(c[3939]) );
  XNOR U1618 ( .A(a[3939]), .B(n1460), .Z(n1458) );
  IV U1619 ( .A(n1456), .Z(n1460) );
  XOR U1620 ( .A(n1461), .B(n1462), .Z(n1456) );
  ANDN U1621 ( .B(n1463), .A(n1464), .Z(n1461) );
  XNOR U1622 ( .A(b[3938]), .B(n1462), .Z(n1463) );
  XNOR U1623 ( .A(b[3938]), .B(n1464), .Z(c[3938]) );
  XNOR U1624 ( .A(a[3938]), .B(n1465), .Z(n1464) );
  IV U1625 ( .A(n1462), .Z(n1465) );
  XOR U1626 ( .A(n1466), .B(n1467), .Z(n1462) );
  ANDN U1627 ( .B(n1468), .A(n1469), .Z(n1466) );
  XNOR U1628 ( .A(b[3937]), .B(n1467), .Z(n1468) );
  XNOR U1629 ( .A(b[3937]), .B(n1469), .Z(c[3937]) );
  XNOR U1630 ( .A(a[3937]), .B(n1470), .Z(n1469) );
  IV U1631 ( .A(n1467), .Z(n1470) );
  XOR U1632 ( .A(n1471), .B(n1472), .Z(n1467) );
  ANDN U1633 ( .B(n1473), .A(n1474), .Z(n1471) );
  XNOR U1634 ( .A(b[3936]), .B(n1472), .Z(n1473) );
  XNOR U1635 ( .A(b[3936]), .B(n1474), .Z(c[3936]) );
  XNOR U1636 ( .A(a[3936]), .B(n1475), .Z(n1474) );
  IV U1637 ( .A(n1472), .Z(n1475) );
  XOR U1638 ( .A(n1476), .B(n1477), .Z(n1472) );
  ANDN U1639 ( .B(n1478), .A(n1479), .Z(n1476) );
  XNOR U1640 ( .A(b[3935]), .B(n1477), .Z(n1478) );
  XNOR U1641 ( .A(b[3935]), .B(n1479), .Z(c[3935]) );
  XNOR U1642 ( .A(a[3935]), .B(n1480), .Z(n1479) );
  IV U1643 ( .A(n1477), .Z(n1480) );
  XOR U1644 ( .A(n1481), .B(n1482), .Z(n1477) );
  ANDN U1645 ( .B(n1483), .A(n1484), .Z(n1481) );
  XNOR U1646 ( .A(b[3934]), .B(n1482), .Z(n1483) );
  XNOR U1647 ( .A(b[3934]), .B(n1484), .Z(c[3934]) );
  XNOR U1648 ( .A(a[3934]), .B(n1485), .Z(n1484) );
  IV U1649 ( .A(n1482), .Z(n1485) );
  XOR U1650 ( .A(n1486), .B(n1487), .Z(n1482) );
  ANDN U1651 ( .B(n1488), .A(n1489), .Z(n1486) );
  XNOR U1652 ( .A(b[3933]), .B(n1487), .Z(n1488) );
  XNOR U1653 ( .A(b[3933]), .B(n1489), .Z(c[3933]) );
  XNOR U1654 ( .A(a[3933]), .B(n1490), .Z(n1489) );
  IV U1655 ( .A(n1487), .Z(n1490) );
  XOR U1656 ( .A(n1491), .B(n1492), .Z(n1487) );
  ANDN U1657 ( .B(n1493), .A(n1494), .Z(n1491) );
  XNOR U1658 ( .A(b[3932]), .B(n1492), .Z(n1493) );
  XNOR U1659 ( .A(b[3932]), .B(n1494), .Z(c[3932]) );
  XNOR U1660 ( .A(a[3932]), .B(n1495), .Z(n1494) );
  IV U1661 ( .A(n1492), .Z(n1495) );
  XOR U1662 ( .A(n1496), .B(n1497), .Z(n1492) );
  ANDN U1663 ( .B(n1498), .A(n1499), .Z(n1496) );
  XNOR U1664 ( .A(b[3931]), .B(n1497), .Z(n1498) );
  XNOR U1665 ( .A(b[3931]), .B(n1499), .Z(c[3931]) );
  XNOR U1666 ( .A(a[3931]), .B(n1500), .Z(n1499) );
  IV U1667 ( .A(n1497), .Z(n1500) );
  XOR U1668 ( .A(n1501), .B(n1502), .Z(n1497) );
  ANDN U1669 ( .B(n1503), .A(n1504), .Z(n1501) );
  XNOR U1670 ( .A(b[3930]), .B(n1502), .Z(n1503) );
  XNOR U1671 ( .A(b[3930]), .B(n1504), .Z(c[3930]) );
  XNOR U1672 ( .A(a[3930]), .B(n1505), .Z(n1504) );
  IV U1673 ( .A(n1502), .Z(n1505) );
  XOR U1674 ( .A(n1506), .B(n1507), .Z(n1502) );
  ANDN U1675 ( .B(n1508), .A(n1509), .Z(n1506) );
  XNOR U1676 ( .A(b[3929]), .B(n1507), .Z(n1508) );
  XNOR U1677 ( .A(b[392]), .B(n1510), .Z(c[392]) );
  XNOR U1678 ( .A(b[3929]), .B(n1509), .Z(c[3929]) );
  XNOR U1679 ( .A(a[3929]), .B(n1511), .Z(n1509) );
  IV U1680 ( .A(n1507), .Z(n1511) );
  XOR U1681 ( .A(n1512), .B(n1513), .Z(n1507) );
  ANDN U1682 ( .B(n1514), .A(n1515), .Z(n1512) );
  XNOR U1683 ( .A(b[3928]), .B(n1513), .Z(n1514) );
  XNOR U1684 ( .A(b[3928]), .B(n1515), .Z(c[3928]) );
  XNOR U1685 ( .A(a[3928]), .B(n1516), .Z(n1515) );
  IV U1686 ( .A(n1513), .Z(n1516) );
  XOR U1687 ( .A(n1517), .B(n1518), .Z(n1513) );
  ANDN U1688 ( .B(n1519), .A(n1520), .Z(n1517) );
  XNOR U1689 ( .A(b[3927]), .B(n1518), .Z(n1519) );
  XNOR U1690 ( .A(b[3927]), .B(n1520), .Z(c[3927]) );
  XNOR U1691 ( .A(a[3927]), .B(n1521), .Z(n1520) );
  IV U1692 ( .A(n1518), .Z(n1521) );
  XOR U1693 ( .A(n1522), .B(n1523), .Z(n1518) );
  ANDN U1694 ( .B(n1524), .A(n1525), .Z(n1522) );
  XNOR U1695 ( .A(b[3926]), .B(n1523), .Z(n1524) );
  XNOR U1696 ( .A(b[3926]), .B(n1525), .Z(c[3926]) );
  XNOR U1697 ( .A(a[3926]), .B(n1526), .Z(n1525) );
  IV U1698 ( .A(n1523), .Z(n1526) );
  XOR U1699 ( .A(n1527), .B(n1528), .Z(n1523) );
  ANDN U1700 ( .B(n1529), .A(n1530), .Z(n1527) );
  XNOR U1701 ( .A(b[3925]), .B(n1528), .Z(n1529) );
  XNOR U1702 ( .A(b[3925]), .B(n1530), .Z(c[3925]) );
  XNOR U1703 ( .A(a[3925]), .B(n1531), .Z(n1530) );
  IV U1704 ( .A(n1528), .Z(n1531) );
  XOR U1705 ( .A(n1532), .B(n1533), .Z(n1528) );
  ANDN U1706 ( .B(n1534), .A(n1535), .Z(n1532) );
  XNOR U1707 ( .A(b[3924]), .B(n1533), .Z(n1534) );
  XNOR U1708 ( .A(b[3924]), .B(n1535), .Z(c[3924]) );
  XNOR U1709 ( .A(a[3924]), .B(n1536), .Z(n1535) );
  IV U1710 ( .A(n1533), .Z(n1536) );
  XOR U1711 ( .A(n1537), .B(n1538), .Z(n1533) );
  ANDN U1712 ( .B(n1539), .A(n1540), .Z(n1537) );
  XNOR U1713 ( .A(b[3923]), .B(n1538), .Z(n1539) );
  XNOR U1714 ( .A(b[3923]), .B(n1540), .Z(c[3923]) );
  XNOR U1715 ( .A(a[3923]), .B(n1541), .Z(n1540) );
  IV U1716 ( .A(n1538), .Z(n1541) );
  XOR U1717 ( .A(n1542), .B(n1543), .Z(n1538) );
  ANDN U1718 ( .B(n1544), .A(n1545), .Z(n1542) );
  XNOR U1719 ( .A(b[3922]), .B(n1543), .Z(n1544) );
  XNOR U1720 ( .A(b[3922]), .B(n1545), .Z(c[3922]) );
  XNOR U1721 ( .A(a[3922]), .B(n1546), .Z(n1545) );
  IV U1722 ( .A(n1543), .Z(n1546) );
  XOR U1723 ( .A(n1547), .B(n1548), .Z(n1543) );
  ANDN U1724 ( .B(n1549), .A(n1550), .Z(n1547) );
  XNOR U1725 ( .A(b[3921]), .B(n1548), .Z(n1549) );
  XNOR U1726 ( .A(b[3921]), .B(n1550), .Z(c[3921]) );
  XNOR U1727 ( .A(a[3921]), .B(n1551), .Z(n1550) );
  IV U1728 ( .A(n1548), .Z(n1551) );
  XOR U1729 ( .A(n1552), .B(n1553), .Z(n1548) );
  ANDN U1730 ( .B(n1554), .A(n1555), .Z(n1552) );
  XNOR U1731 ( .A(b[3920]), .B(n1553), .Z(n1554) );
  XNOR U1732 ( .A(b[3920]), .B(n1555), .Z(c[3920]) );
  XNOR U1733 ( .A(a[3920]), .B(n1556), .Z(n1555) );
  IV U1734 ( .A(n1553), .Z(n1556) );
  XOR U1735 ( .A(n1557), .B(n1558), .Z(n1553) );
  ANDN U1736 ( .B(n1559), .A(n1560), .Z(n1557) );
  XNOR U1737 ( .A(b[3919]), .B(n1558), .Z(n1559) );
  XNOR U1738 ( .A(b[391]), .B(n1561), .Z(c[391]) );
  XNOR U1739 ( .A(b[3919]), .B(n1560), .Z(c[3919]) );
  XNOR U1740 ( .A(a[3919]), .B(n1562), .Z(n1560) );
  IV U1741 ( .A(n1558), .Z(n1562) );
  XOR U1742 ( .A(n1563), .B(n1564), .Z(n1558) );
  ANDN U1743 ( .B(n1565), .A(n1566), .Z(n1563) );
  XNOR U1744 ( .A(b[3918]), .B(n1564), .Z(n1565) );
  XNOR U1745 ( .A(b[3918]), .B(n1566), .Z(c[3918]) );
  XNOR U1746 ( .A(a[3918]), .B(n1567), .Z(n1566) );
  IV U1747 ( .A(n1564), .Z(n1567) );
  XOR U1748 ( .A(n1568), .B(n1569), .Z(n1564) );
  ANDN U1749 ( .B(n1570), .A(n1571), .Z(n1568) );
  XNOR U1750 ( .A(b[3917]), .B(n1569), .Z(n1570) );
  XNOR U1751 ( .A(b[3917]), .B(n1571), .Z(c[3917]) );
  XNOR U1752 ( .A(a[3917]), .B(n1572), .Z(n1571) );
  IV U1753 ( .A(n1569), .Z(n1572) );
  XOR U1754 ( .A(n1573), .B(n1574), .Z(n1569) );
  ANDN U1755 ( .B(n1575), .A(n1576), .Z(n1573) );
  XNOR U1756 ( .A(b[3916]), .B(n1574), .Z(n1575) );
  XNOR U1757 ( .A(b[3916]), .B(n1576), .Z(c[3916]) );
  XNOR U1758 ( .A(a[3916]), .B(n1577), .Z(n1576) );
  IV U1759 ( .A(n1574), .Z(n1577) );
  XOR U1760 ( .A(n1578), .B(n1579), .Z(n1574) );
  ANDN U1761 ( .B(n1580), .A(n1581), .Z(n1578) );
  XNOR U1762 ( .A(b[3915]), .B(n1579), .Z(n1580) );
  XNOR U1763 ( .A(b[3915]), .B(n1581), .Z(c[3915]) );
  XNOR U1764 ( .A(a[3915]), .B(n1582), .Z(n1581) );
  IV U1765 ( .A(n1579), .Z(n1582) );
  XOR U1766 ( .A(n1583), .B(n1584), .Z(n1579) );
  ANDN U1767 ( .B(n1585), .A(n1586), .Z(n1583) );
  XNOR U1768 ( .A(b[3914]), .B(n1584), .Z(n1585) );
  XNOR U1769 ( .A(b[3914]), .B(n1586), .Z(c[3914]) );
  XNOR U1770 ( .A(a[3914]), .B(n1587), .Z(n1586) );
  IV U1771 ( .A(n1584), .Z(n1587) );
  XOR U1772 ( .A(n1588), .B(n1589), .Z(n1584) );
  ANDN U1773 ( .B(n1590), .A(n1591), .Z(n1588) );
  XNOR U1774 ( .A(b[3913]), .B(n1589), .Z(n1590) );
  XNOR U1775 ( .A(b[3913]), .B(n1591), .Z(c[3913]) );
  XNOR U1776 ( .A(a[3913]), .B(n1592), .Z(n1591) );
  IV U1777 ( .A(n1589), .Z(n1592) );
  XOR U1778 ( .A(n1593), .B(n1594), .Z(n1589) );
  ANDN U1779 ( .B(n1595), .A(n1596), .Z(n1593) );
  XNOR U1780 ( .A(b[3912]), .B(n1594), .Z(n1595) );
  XNOR U1781 ( .A(b[3912]), .B(n1596), .Z(c[3912]) );
  XNOR U1782 ( .A(a[3912]), .B(n1597), .Z(n1596) );
  IV U1783 ( .A(n1594), .Z(n1597) );
  XOR U1784 ( .A(n1598), .B(n1599), .Z(n1594) );
  ANDN U1785 ( .B(n1600), .A(n1601), .Z(n1598) );
  XNOR U1786 ( .A(b[3911]), .B(n1599), .Z(n1600) );
  XNOR U1787 ( .A(b[3911]), .B(n1601), .Z(c[3911]) );
  XNOR U1788 ( .A(a[3911]), .B(n1602), .Z(n1601) );
  IV U1789 ( .A(n1599), .Z(n1602) );
  XOR U1790 ( .A(n1603), .B(n1604), .Z(n1599) );
  ANDN U1791 ( .B(n1605), .A(n1606), .Z(n1603) );
  XNOR U1792 ( .A(b[3910]), .B(n1604), .Z(n1605) );
  XNOR U1793 ( .A(b[3910]), .B(n1606), .Z(c[3910]) );
  XNOR U1794 ( .A(a[3910]), .B(n1607), .Z(n1606) );
  IV U1795 ( .A(n1604), .Z(n1607) );
  XOR U1796 ( .A(n1608), .B(n1609), .Z(n1604) );
  ANDN U1797 ( .B(n1610), .A(n1611), .Z(n1608) );
  XNOR U1798 ( .A(b[3909]), .B(n1609), .Z(n1610) );
  XNOR U1799 ( .A(b[390]), .B(n1612), .Z(c[390]) );
  XNOR U1800 ( .A(b[3909]), .B(n1611), .Z(c[3909]) );
  XNOR U1801 ( .A(a[3909]), .B(n1613), .Z(n1611) );
  IV U1802 ( .A(n1609), .Z(n1613) );
  XOR U1803 ( .A(n1614), .B(n1615), .Z(n1609) );
  ANDN U1804 ( .B(n1616), .A(n1617), .Z(n1614) );
  XNOR U1805 ( .A(b[3908]), .B(n1615), .Z(n1616) );
  XNOR U1806 ( .A(b[3908]), .B(n1617), .Z(c[3908]) );
  XNOR U1807 ( .A(a[3908]), .B(n1618), .Z(n1617) );
  IV U1808 ( .A(n1615), .Z(n1618) );
  XOR U1809 ( .A(n1619), .B(n1620), .Z(n1615) );
  ANDN U1810 ( .B(n1621), .A(n1622), .Z(n1619) );
  XNOR U1811 ( .A(b[3907]), .B(n1620), .Z(n1621) );
  XNOR U1812 ( .A(b[3907]), .B(n1622), .Z(c[3907]) );
  XNOR U1813 ( .A(a[3907]), .B(n1623), .Z(n1622) );
  IV U1814 ( .A(n1620), .Z(n1623) );
  XOR U1815 ( .A(n1624), .B(n1625), .Z(n1620) );
  ANDN U1816 ( .B(n1626), .A(n1627), .Z(n1624) );
  XNOR U1817 ( .A(b[3906]), .B(n1625), .Z(n1626) );
  XNOR U1818 ( .A(b[3906]), .B(n1627), .Z(c[3906]) );
  XNOR U1819 ( .A(a[3906]), .B(n1628), .Z(n1627) );
  IV U1820 ( .A(n1625), .Z(n1628) );
  XOR U1821 ( .A(n1629), .B(n1630), .Z(n1625) );
  ANDN U1822 ( .B(n1631), .A(n1632), .Z(n1629) );
  XNOR U1823 ( .A(b[3905]), .B(n1630), .Z(n1631) );
  XNOR U1824 ( .A(b[3905]), .B(n1632), .Z(c[3905]) );
  XNOR U1825 ( .A(a[3905]), .B(n1633), .Z(n1632) );
  IV U1826 ( .A(n1630), .Z(n1633) );
  XOR U1827 ( .A(n1634), .B(n1635), .Z(n1630) );
  ANDN U1828 ( .B(n1636), .A(n1637), .Z(n1634) );
  XNOR U1829 ( .A(b[3904]), .B(n1635), .Z(n1636) );
  XNOR U1830 ( .A(b[3904]), .B(n1637), .Z(c[3904]) );
  XNOR U1831 ( .A(a[3904]), .B(n1638), .Z(n1637) );
  IV U1832 ( .A(n1635), .Z(n1638) );
  XOR U1833 ( .A(n1639), .B(n1640), .Z(n1635) );
  ANDN U1834 ( .B(n1641), .A(n1642), .Z(n1639) );
  XNOR U1835 ( .A(b[3903]), .B(n1640), .Z(n1641) );
  XNOR U1836 ( .A(b[3903]), .B(n1642), .Z(c[3903]) );
  XNOR U1837 ( .A(a[3903]), .B(n1643), .Z(n1642) );
  IV U1838 ( .A(n1640), .Z(n1643) );
  XOR U1839 ( .A(n1644), .B(n1645), .Z(n1640) );
  ANDN U1840 ( .B(n1646), .A(n1647), .Z(n1644) );
  XNOR U1841 ( .A(b[3902]), .B(n1645), .Z(n1646) );
  XNOR U1842 ( .A(b[3902]), .B(n1647), .Z(c[3902]) );
  XNOR U1843 ( .A(a[3902]), .B(n1648), .Z(n1647) );
  IV U1844 ( .A(n1645), .Z(n1648) );
  XOR U1845 ( .A(n1649), .B(n1650), .Z(n1645) );
  ANDN U1846 ( .B(n1651), .A(n1652), .Z(n1649) );
  XNOR U1847 ( .A(b[3901]), .B(n1650), .Z(n1651) );
  XNOR U1848 ( .A(b[3901]), .B(n1652), .Z(c[3901]) );
  XNOR U1849 ( .A(a[3901]), .B(n1653), .Z(n1652) );
  IV U1850 ( .A(n1650), .Z(n1653) );
  XOR U1851 ( .A(n1654), .B(n1655), .Z(n1650) );
  ANDN U1852 ( .B(n1656), .A(n1657), .Z(n1654) );
  XNOR U1853 ( .A(b[3900]), .B(n1655), .Z(n1656) );
  XNOR U1854 ( .A(b[3900]), .B(n1657), .Z(c[3900]) );
  XNOR U1855 ( .A(a[3900]), .B(n1658), .Z(n1657) );
  IV U1856 ( .A(n1655), .Z(n1658) );
  XOR U1857 ( .A(n1659), .B(n1660), .Z(n1655) );
  ANDN U1858 ( .B(n1661), .A(n1662), .Z(n1659) );
  XNOR U1859 ( .A(b[3899]), .B(n1660), .Z(n1661) );
  XNOR U1860 ( .A(b[38]), .B(n1663), .Z(c[38]) );
  XNOR U1861 ( .A(b[389]), .B(n1664), .Z(c[389]) );
  XNOR U1862 ( .A(b[3899]), .B(n1662), .Z(c[3899]) );
  XNOR U1863 ( .A(a[3899]), .B(n1665), .Z(n1662) );
  IV U1864 ( .A(n1660), .Z(n1665) );
  XOR U1865 ( .A(n1666), .B(n1667), .Z(n1660) );
  ANDN U1866 ( .B(n1668), .A(n1669), .Z(n1666) );
  XNOR U1867 ( .A(b[3898]), .B(n1667), .Z(n1668) );
  XNOR U1868 ( .A(b[3898]), .B(n1669), .Z(c[3898]) );
  XNOR U1869 ( .A(a[3898]), .B(n1670), .Z(n1669) );
  IV U1870 ( .A(n1667), .Z(n1670) );
  XOR U1871 ( .A(n1671), .B(n1672), .Z(n1667) );
  ANDN U1872 ( .B(n1673), .A(n1674), .Z(n1671) );
  XNOR U1873 ( .A(b[3897]), .B(n1672), .Z(n1673) );
  XNOR U1874 ( .A(b[3897]), .B(n1674), .Z(c[3897]) );
  XNOR U1875 ( .A(a[3897]), .B(n1675), .Z(n1674) );
  IV U1876 ( .A(n1672), .Z(n1675) );
  XOR U1877 ( .A(n1676), .B(n1677), .Z(n1672) );
  ANDN U1878 ( .B(n1678), .A(n1679), .Z(n1676) );
  XNOR U1879 ( .A(b[3896]), .B(n1677), .Z(n1678) );
  XNOR U1880 ( .A(b[3896]), .B(n1679), .Z(c[3896]) );
  XNOR U1881 ( .A(a[3896]), .B(n1680), .Z(n1679) );
  IV U1882 ( .A(n1677), .Z(n1680) );
  XOR U1883 ( .A(n1681), .B(n1682), .Z(n1677) );
  ANDN U1884 ( .B(n1683), .A(n1684), .Z(n1681) );
  XNOR U1885 ( .A(b[3895]), .B(n1682), .Z(n1683) );
  XNOR U1886 ( .A(b[3895]), .B(n1684), .Z(c[3895]) );
  XNOR U1887 ( .A(a[3895]), .B(n1685), .Z(n1684) );
  IV U1888 ( .A(n1682), .Z(n1685) );
  XOR U1889 ( .A(n1686), .B(n1687), .Z(n1682) );
  ANDN U1890 ( .B(n1688), .A(n1689), .Z(n1686) );
  XNOR U1891 ( .A(b[3894]), .B(n1687), .Z(n1688) );
  XNOR U1892 ( .A(b[3894]), .B(n1689), .Z(c[3894]) );
  XNOR U1893 ( .A(a[3894]), .B(n1690), .Z(n1689) );
  IV U1894 ( .A(n1687), .Z(n1690) );
  XOR U1895 ( .A(n1691), .B(n1692), .Z(n1687) );
  ANDN U1896 ( .B(n1693), .A(n1694), .Z(n1691) );
  XNOR U1897 ( .A(b[3893]), .B(n1692), .Z(n1693) );
  XNOR U1898 ( .A(b[3893]), .B(n1694), .Z(c[3893]) );
  XNOR U1899 ( .A(a[3893]), .B(n1695), .Z(n1694) );
  IV U1900 ( .A(n1692), .Z(n1695) );
  XOR U1901 ( .A(n1696), .B(n1697), .Z(n1692) );
  ANDN U1902 ( .B(n1698), .A(n1699), .Z(n1696) );
  XNOR U1903 ( .A(b[3892]), .B(n1697), .Z(n1698) );
  XNOR U1904 ( .A(b[3892]), .B(n1699), .Z(c[3892]) );
  XNOR U1905 ( .A(a[3892]), .B(n1700), .Z(n1699) );
  IV U1906 ( .A(n1697), .Z(n1700) );
  XOR U1907 ( .A(n1701), .B(n1702), .Z(n1697) );
  ANDN U1908 ( .B(n1703), .A(n1704), .Z(n1701) );
  XNOR U1909 ( .A(b[3891]), .B(n1702), .Z(n1703) );
  XNOR U1910 ( .A(b[3891]), .B(n1704), .Z(c[3891]) );
  XNOR U1911 ( .A(a[3891]), .B(n1705), .Z(n1704) );
  IV U1912 ( .A(n1702), .Z(n1705) );
  XOR U1913 ( .A(n1706), .B(n1707), .Z(n1702) );
  ANDN U1914 ( .B(n1708), .A(n1709), .Z(n1706) );
  XNOR U1915 ( .A(b[3890]), .B(n1707), .Z(n1708) );
  XNOR U1916 ( .A(b[3890]), .B(n1709), .Z(c[3890]) );
  XNOR U1917 ( .A(a[3890]), .B(n1710), .Z(n1709) );
  IV U1918 ( .A(n1707), .Z(n1710) );
  XOR U1919 ( .A(n1711), .B(n1712), .Z(n1707) );
  ANDN U1920 ( .B(n1713), .A(n1714), .Z(n1711) );
  XNOR U1921 ( .A(b[3889]), .B(n1712), .Z(n1713) );
  XNOR U1922 ( .A(b[388]), .B(n1715), .Z(c[388]) );
  XNOR U1923 ( .A(b[3889]), .B(n1714), .Z(c[3889]) );
  XNOR U1924 ( .A(a[3889]), .B(n1716), .Z(n1714) );
  IV U1925 ( .A(n1712), .Z(n1716) );
  XOR U1926 ( .A(n1717), .B(n1718), .Z(n1712) );
  ANDN U1927 ( .B(n1719), .A(n1720), .Z(n1717) );
  XNOR U1928 ( .A(b[3888]), .B(n1718), .Z(n1719) );
  XNOR U1929 ( .A(b[3888]), .B(n1720), .Z(c[3888]) );
  XNOR U1930 ( .A(a[3888]), .B(n1721), .Z(n1720) );
  IV U1931 ( .A(n1718), .Z(n1721) );
  XOR U1932 ( .A(n1722), .B(n1723), .Z(n1718) );
  ANDN U1933 ( .B(n1724), .A(n1725), .Z(n1722) );
  XNOR U1934 ( .A(b[3887]), .B(n1723), .Z(n1724) );
  XNOR U1935 ( .A(b[3887]), .B(n1725), .Z(c[3887]) );
  XNOR U1936 ( .A(a[3887]), .B(n1726), .Z(n1725) );
  IV U1937 ( .A(n1723), .Z(n1726) );
  XOR U1938 ( .A(n1727), .B(n1728), .Z(n1723) );
  ANDN U1939 ( .B(n1729), .A(n1730), .Z(n1727) );
  XNOR U1940 ( .A(b[3886]), .B(n1728), .Z(n1729) );
  XNOR U1941 ( .A(b[3886]), .B(n1730), .Z(c[3886]) );
  XNOR U1942 ( .A(a[3886]), .B(n1731), .Z(n1730) );
  IV U1943 ( .A(n1728), .Z(n1731) );
  XOR U1944 ( .A(n1732), .B(n1733), .Z(n1728) );
  ANDN U1945 ( .B(n1734), .A(n1735), .Z(n1732) );
  XNOR U1946 ( .A(b[3885]), .B(n1733), .Z(n1734) );
  XNOR U1947 ( .A(b[3885]), .B(n1735), .Z(c[3885]) );
  XNOR U1948 ( .A(a[3885]), .B(n1736), .Z(n1735) );
  IV U1949 ( .A(n1733), .Z(n1736) );
  XOR U1950 ( .A(n1737), .B(n1738), .Z(n1733) );
  ANDN U1951 ( .B(n1739), .A(n1740), .Z(n1737) );
  XNOR U1952 ( .A(b[3884]), .B(n1738), .Z(n1739) );
  XNOR U1953 ( .A(b[3884]), .B(n1740), .Z(c[3884]) );
  XNOR U1954 ( .A(a[3884]), .B(n1741), .Z(n1740) );
  IV U1955 ( .A(n1738), .Z(n1741) );
  XOR U1956 ( .A(n1742), .B(n1743), .Z(n1738) );
  ANDN U1957 ( .B(n1744), .A(n1745), .Z(n1742) );
  XNOR U1958 ( .A(b[3883]), .B(n1743), .Z(n1744) );
  XNOR U1959 ( .A(b[3883]), .B(n1745), .Z(c[3883]) );
  XNOR U1960 ( .A(a[3883]), .B(n1746), .Z(n1745) );
  IV U1961 ( .A(n1743), .Z(n1746) );
  XOR U1962 ( .A(n1747), .B(n1748), .Z(n1743) );
  ANDN U1963 ( .B(n1749), .A(n1750), .Z(n1747) );
  XNOR U1964 ( .A(b[3882]), .B(n1748), .Z(n1749) );
  XNOR U1965 ( .A(b[3882]), .B(n1750), .Z(c[3882]) );
  XNOR U1966 ( .A(a[3882]), .B(n1751), .Z(n1750) );
  IV U1967 ( .A(n1748), .Z(n1751) );
  XOR U1968 ( .A(n1752), .B(n1753), .Z(n1748) );
  ANDN U1969 ( .B(n1754), .A(n1755), .Z(n1752) );
  XNOR U1970 ( .A(b[3881]), .B(n1753), .Z(n1754) );
  XNOR U1971 ( .A(b[3881]), .B(n1755), .Z(c[3881]) );
  XNOR U1972 ( .A(a[3881]), .B(n1756), .Z(n1755) );
  IV U1973 ( .A(n1753), .Z(n1756) );
  XOR U1974 ( .A(n1757), .B(n1758), .Z(n1753) );
  ANDN U1975 ( .B(n1759), .A(n1760), .Z(n1757) );
  XNOR U1976 ( .A(b[3880]), .B(n1758), .Z(n1759) );
  XNOR U1977 ( .A(b[3880]), .B(n1760), .Z(c[3880]) );
  XNOR U1978 ( .A(a[3880]), .B(n1761), .Z(n1760) );
  IV U1979 ( .A(n1758), .Z(n1761) );
  XOR U1980 ( .A(n1762), .B(n1763), .Z(n1758) );
  ANDN U1981 ( .B(n1764), .A(n1765), .Z(n1762) );
  XNOR U1982 ( .A(b[3879]), .B(n1763), .Z(n1764) );
  XNOR U1983 ( .A(b[387]), .B(n1766), .Z(c[387]) );
  XNOR U1984 ( .A(b[3879]), .B(n1765), .Z(c[3879]) );
  XNOR U1985 ( .A(a[3879]), .B(n1767), .Z(n1765) );
  IV U1986 ( .A(n1763), .Z(n1767) );
  XOR U1987 ( .A(n1768), .B(n1769), .Z(n1763) );
  ANDN U1988 ( .B(n1770), .A(n1771), .Z(n1768) );
  XNOR U1989 ( .A(b[3878]), .B(n1769), .Z(n1770) );
  XNOR U1990 ( .A(b[3878]), .B(n1771), .Z(c[3878]) );
  XNOR U1991 ( .A(a[3878]), .B(n1772), .Z(n1771) );
  IV U1992 ( .A(n1769), .Z(n1772) );
  XOR U1993 ( .A(n1773), .B(n1774), .Z(n1769) );
  ANDN U1994 ( .B(n1775), .A(n1776), .Z(n1773) );
  XNOR U1995 ( .A(b[3877]), .B(n1774), .Z(n1775) );
  XNOR U1996 ( .A(b[3877]), .B(n1776), .Z(c[3877]) );
  XNOR U1997 ( .A(a[3877]), .B(n1777), .Z(n1776) );
  IV U1998 ( .A(n1774), .Z(n1777) );
  XOR U1999 ( .A(n1778), .B(n1779), .Z(n1774) );
  ANDN U2000 ( .B(n1780), .A(n1781), .Z(n1778) );
  XNOR U2001 ( .A(b[3876]), .B(n1779), .Z(n1780) );
  XNOR U2002 ( .A(b[3876]), .B(n1781), .Z(c[3876]) );
  XNOR U2003 ( .A(a[3876]), .B(n1782), .Z(n1781) );
  IV U2004 ( .A(n1779), .Z(n1782) );
  XOR U2005 ( .A(n1783), .B(n1784), .Z(n1779) );
  ANDN U2006 ( .B(n1785), .A(n1786), .Z(n1783) );
  XNOR U2007 ( .A(b[3875]), .B(n1784), .Z(n1785) );
  XNOR U2008 ( .A(b[3875]), .B(n1786), .Z(c[3875]) );
  XNOR U2009 ( .A(a[3875]), .B(n1787), .Z(n1786) );
  IV U2010 ( .A(n1784), .Z(n1787) );
  XOR U2011 ( .A(n1788), .B(n1789), .Z(n1784) );
  ANDN U2012 ( .B(n1790), .A(n1791), .Z(n1788) );
  XNOR U2013 ( .A(b[3874]), .B(n1789), .Z(n1790) );
  XNOR U2014 ( .A(b[3874]), .B(n1791), .Z(c[3874]) );
  XNOR U2015 ( .A(a[3874]), .B(n1792), .Z(n1791) );
  IV U2016 ( .A(n1789), .Z(n1792) );
  XOR U2017 ( .A(n1793), .B(n1794), .Z(n1789) );
  ANDN U2018 ( .B(n1795), .A(n1796), .Z(n1793) );
  XNOR U2019 ( .A(b[3873]), .B(n1794), .Z(n1795) );
  XNOR U2020 ( .A(b[3873]), .B(n1796), .Z(c[3873]) );
  XNOR U2021 ( .A(a[3873]), .B(n1797), .Z(n1796) );
  IV U2022 ( .A(n1794), .Z(n1797) );
  XOR U2023 ( .A(n1798), .B(n1799), .Z(n1794) );
  ANDN U2024 ( .B(n1800), .A(n1801), .Z(n1798) );
  XNOR U2025 ( .A(b[3872]), .B(n1799), .Z(n1800) );
  XNOR U2026 ( .A(b[3872]), .B(n1801), .Z(c[3872]) );
  XNOR U2027 ( .A(a[3872]), .B(n1802), .Z(n1801) );
  IV U2028 ( .A(n1799), .Z(n1802) );
  XOR U2029 ( .A(n1803), .B(n1804), .Z(n1799) );
  ANDN U2030 ( .B(n1805), .A(n1806), .Z(n1803) );
  XNOR U2031 ( .A(b[3871]), .B(n1804), .Z(n1805) );
  XNOR U2032 ( .A(b[3871]), .B(n1806), .Z(c[3871]) );
  XNOR U2033 ( .A(a[3871]), .B(n1807), .Z(n1806) );
  IV U2034 ( .A(n1804), .Z(n1807) );
  XOR U2035 ( .A(n1808), .B(n1809), .Z(n1804) );
  ANDN U2036 ( .B(n1810), .A(n1811), .Z(n1808) );
  XNOR U2037 ( .A(b[3870]), .B(n1809), .Z(n1810) );
  XNOR U2038 ( .A(b[3870]), .B(n1811), .Z(c[3870]) );
  XNOR U2039 ( .A(a[3870]), .B(n1812), .Z(n1811) );
  IV U2040 ( .A(n1809), .Z(n1812) );
  XOR U2041 ( .A(n1813), .B(n1814), .Z(n1809) );
  ANDN U2042 ( .B(n1815), .A(n1816), .Z(n1813) );
  XNOR U2043 ( .A(b[3869]), .B(n1814), .Z(n1815) );
  XNOR U2044 ( .A(b[386]), .B(n1817), .Z(c[386]) );
  XNOR U2045 ( .A(b[3869]), .B(n1816), .Z(c[3869]) );
  XNOR U2046 ( .A(a[3869]), .B(n1818), .Z(n1816) );
  IV U2047 ( .A(n1814), .Z(n1818) );
  XOR U2048 ( .A(n1819), .B(n1820), .Z(n1814) );
  ANDN U2049 ( .B(n1821), .A(n1822), .Z(n1819) );
  XNOR U2050 ( .A(b[3868]), .B(n1820), .Z(n1821) );
  XNOR U2051 ( .A(b[3868]), .B(n1822), .Z(c[3868]) );
  XNOR U2052 ( .A(a[3868]), .B(n1823), .Z(n1822) );
  IV U2053 ( .A(n1820), .Z(n1823) );
  XOR U2054 ( .A(n1824), .B(n1825), .Z(n1820) );
  ANDN U2055 ( .B(n1826), .A(n1827), .Z(n1824) );
  XNOR U2056 ( .A(b[3867]), .B(n1825), .Z(n1826) );
  XNOR U2057 ( .A(b[3867]), .B(n1827), .Z(c[3867]) );
  XNOR U2058 ( .A(a[3867]), .B(n1828), .Z(n1827) );
  IV U2059 ( .A(n1825), .Z(n1828) );
  XOR U2060 ( .A(n1829), .B(n1830), .Z(n1825) );
  ANDN U2061 ( .B(n1831), .A(n1832), .Z(n1829) );
  XNOR U2062 ( .A(b[3866]), .B(n1830), .Z(n1831) );
  XNOR U2063 ( .A(b[3866]), .B(n1832), .Z(c[3866]) );
  XNOR U2064 ( .A(a[3866]), .B(n1833), .Z(n1832) );
  IV U2065 ( .A(n1830), .Z(n1833) );
  XOR U2066 ( .A(n1834), .B(n1835), .Z(n1830) );
  ANDN U2067 ( .B(n1836), .A(n1837), .Z(n1834) );
  XNOR U2068 ( .A(b[3865]), .B(n1835), .Z(n1836) );
  XNOR U2069 ( .A(b[3865]), .B(n1837), .Z(c[3865]) );
  XNOR U2070 ( .A(a[3865]), .B(n1838), .Z(n1837) );
  IV U2071 ( .A(n1835), .Z(n1838) );
  XOR U2072 ( .A(n1839), .B(n1840), .Z(n1835) );
  ANDN U2073 ( .B(n1841), .A(n1842), .Z(n1839) );
  XNOR U2074 ( .A(b[3864]), .B(n1840), .Z(n1841) );
  XNOR U2075 ( .A(b[3864]), .B(n1842), .Z(c[3864]) );
  XNOR U2076 ( .A(a[3864]), .B(n1843), .Z(n1842) );
  IV U2077 ( .A(n1840), .Z(n1843) );
  XOR U2078 ( .A(n1844), .B(n1845), .Z(n1840) );
  ANDN U2079 ( .B(n1846), .A(n1847), .Z(n1844) );
  XNOR U2080 ( .A(b[3863]), .B(n1845), .Z(n1846) );
  XNOR U2081 ( .A(b[3863]), .B(n1847), .Z(c[3863]) );
  XNOR U2082 ( .A(a[3863]), .B(n1848), .Z(n1847) );
  IV U2083 ( .A(n1845), .Z(n1848) );
  XOR U2084 ( .A(n1849), .B(n1850), .Z(n1845) );
  ANDN U2085 ( .B(n1851), .A(n1852), .Z(n1849) );
  XNOR U2086 ( .A(b[3862]), .B(n1850), .Z(n1851) );
  XNOR U2087 ( .A(b[3862]), .B(n1852), .Z(c[3862]) );
  XNOR U2088 ( .A(a[3862]), .B(n1853), .Z(n1852) );
  IV U2089 ( .A(n1850), .Z(n1853) );
  XOR U2090 ( .A(n1854), .B(n1855), .Z(n1850) );
  ANDN U2091 ( .B(n1856), .A(n1857), .Z(n1854) );
  XNOR U2092 ( .A(b[3861]), .B(n1855), .Z(n1856) );
  XNOR U2093 ( .A(b[3861]), .B(n1857), .Z(c[3861]) );
  XNOR U2094 ( .A(a[3861]), .B(n1858), .Z(n1857) );
  IV U2095 ( .A(n1855), .Z(n1858) );
  XOR U2096 ( .A(n1859), .B(n1860), .Z(n1855) );
  ANDN U2097 ( .B(n1861), .A(n1862), .Z(n1859) );
  XNOR U2098 ( .A(b[3860]), .B(n1860), .Z(n1861) );
  XNOR U2099 ( .A(b[3860]), .B(n1862), .Z(c[3860]) );
  XNOR U2100 ( .A(a[3860]), .B(n1863), .Z(n1862) );
  IV U2101 ( .A(n1860), .Z(n1863) );
  XOR U2102 ( .A(n1864), .B(n1865), .Z(n1860) );
  ANDN U2103 ( .B(n1866), .A(n1867), .Z(n1864) );
  XNOR U2104 ( .A(b[3859]), .B(n1865), .Z(n1866) );
  XNOR U2105 ( .A(b[385]), .B(n1868), .Z(c[385]) );
  XNOR U2106 ( .A(b[3859]), .B(n1867), .Z(c[3859]) );
  XNOR U2107 ( .A(a[3859]), .B(n1869), .Z(n1867) );
  IV U2108 ( .A(n1865), .Z(n1869) );
  XOR U2109 ( .A(n1870), .B(n1871), .Z(n1865) );
  ANDN U2110 ( .B(n1872), .A(n1873), .Z(n1870) );
  XNOR U2111 ( .A(b[3858]), .B(n1871), .Z(n1872) );
  XNOR U2112 ( .A(b[3858]), .B(n1873), .Z(c[3858]) );
  XNOR U2113 ( .A(a[3858]), .B(n1874), .Z(n1873) );
  IV U2114 ( .A(n1871), .Z(n1874) );
  XOR U2115 ( .A(n1875), .B(n1876), .Z(n1871) );
  ANDN U2116 ( .B(n1877), .A(n1878), .Z(n1875) );
  XNOR U2117 ( .A(b[3857]), .B(n1876), .Z(n1877) );
  XNOR U2118 ( .A(b[3857]), .B(n1878), .Z(c[3857]) );
  XNOR U2119 ( .A(a[3857]), .B(n1879), .Z(n1878) );
  IV U2120 ( .A(n1876), .Z(n1879) );
  XOR U2121 ( .A(n1880), .B(n1881), .Z(n1876) );
  ANDN U2122 ( .B(n1882), .A(n1883), .Z(n1880) );
  XNOR U2123 ( .A(b[3856]), .B(n1881), .Z(n1882) );
  XNOR U2124 ( .A(b[3856]), .B(n1883), .Z(c[3856]) );
  XNOR U2125 ( .A(a[3856]), .B(n1884), .Z(n1883) );
  IV U2126 ( .A(n1881), .Z(n1884) );
  XOR U2127 ( .A(n1885), .B(n1886), .Z(n1881) );
  ANDN U2128 ( .B(n1887), .A(n1888), .Z(n1885) );
  XNOR U2129 ( .A(b[3855]), .B(n1886), .Z(n1887) );
  XNOR U2130 ( .A(b[3855]), .B(n1888), .Z(c[3855]) );
  XNOR U2131 ( .A(a[3855]), .B(n1889), .Z(n1888) );
  IV U2132 ( .A(n1886), .Z(n1889) );
  XOR U2133 ( .A(n1890), .B(n1891), .Z(n1886) );
  ANDN U2134 ( .B(n1892), .A(n1893), .Z(n1890) );
  XNOR U2135 ( .A(b[3854]), .B(n1891), .Z(n1892) );
  XNOR U2136 ( .A(b[3854]), .B(n1893), .Z(c[3854]) );
  XNOR U2137 ( .A(a[3854]), .B(n1894), .Z(n1893) );
  IV U2138 ( .A(n1891), .Z(n1894) );
  XOR U2139 ( .A(n1895), .B(n1896), .Z(n1891) );
  ANDN U2140 ( .B(n1897), .A(n1898), .Z(n1895) );
  XNOR U2141 ( .A(b[3853]), .B(n1896), .Z(n1897) );
  XNOR U2142 ( .A(b[3853]), .B(n1898), .Z(c[3853]) );
  XNOR U2143 ( .A(a[3853]), .B(n1899), .Z(n1898) );
  IV U2144 ( .A(n1896), .Z(n1899) );
  XOR U2145 ( .A(n1900), .B(n1901), .Z(n1896) );
  ANDN U2146 ( .B(n1902), .A(n1903), .Z(n1900) );
  XNOR U2147 ( .A(b[3852]), .B(n1901), .Z(n1902) );
  XNOR U2148 ( .A(b[3852]), .B(n1903), .Z(c[3852]) );
  XNOR U2149 ( .A(a[3852]), .B(n1904), .Z(n1903) );
  IV U2150 ( .A(n1901), .Z(n1904) );
  XOR U2151 ( .A(n1905), .B(n1906), .Z(n1901) );
  ANDN U2152 ( .B(n1907), .A(n1908), .Z(n1905) );
  XNOR U2153 ( .A(b[3851]), .B(n1906), .Z(n1907) );
  XNOR U2154 ( .A(b[3851]), .B(n1908), .Z(c[3851]) );
  XNOR U2155 ( .A(a[3851]), .B(n1909), .Z(n1908) );
  IV U2156 ( .A(n1906), .Z(n1909) );
  XOR U2157 ( .A(n1910), .B(n1911), .Z(n1906) );
  ANDN U2158 ( .B(n1912), .A(n1913), .Z(n1910) );
  XNOR U2159 ( .A(b[3850]), .B(n1911), .Z(n1912) );
  XNOR U2160 ( .A(b[3850]), .B(n1913), .Z(c[3850]) );
  XNOR U2161 ( .A(a[3850]), .B(n1914), .Z(n1913) );
  IV U2162 ( .A(n1911), .Z(n1914) );
  XOR U2163 ( .A(n1915), .B(n1916), .Z(n1911) );
  ANDN U2164 ( .B(n1917), .A(n1918), .Z(n1915) );
  XNOR U2165 ( .A(b[3849]), .B(n1916), .Z(n1917) );
  XNOR U2166 ( .A(b[384]), .B(n1919), .Z(c[384]) );
  XNOR U2167 ( .A(b[3849]), .B(n1918), .Z(c[3849]) );
  XNOR U2168 ( .A(a[3849]), .B(n1920), .Z(n1918) );
  IV U2169 ( .A(n1916), .Z(n1920) );
  XOR U2170 ( .A(n1921), .B(n1922), .Z(n1916) );
  ANDN U2171 ( .B(n1923), .A(n1924), .Z(n1921) );
  XNOR U2172 ( .A(b[3848]), .B(n1922), .Z(n1923) );
  XNOR U2173 ( .A(b[3848]), .B(n1924), .Z(c[3848]) );
  XNOR U2174 ( .A(a[3848]), .B(n1925), .Z(n1924) );
  IV U2175 ( .A(n1922), .Z(n1925) );
  XOR U2176 ( .A(n1926), .B(n1927), .Z(n1922) );
  ANDN U2177 ( .B(n1928), .A(n1929), .Z(n1926) );
  XNOR U2178 ( .A(b[3847]), .B(n1927), .Z(n1928) );
  XNOR U2179 ( .A(b[3847]), .B(n1929), .Z(c[3847]) );
  XNOR U2180 ( .A(a[3847]), .B(n1930), .Z(n1929) );
  IV U2181 ( .A(n1927), .Z(n1930) );
  XOR U2182 ( .A(n1931), .B(n1932), .Z(n1927) );
  ANDN U2183 ( .B(n1933), .A(n1934), .Z(n1931) );
  XNOR U2184 ( .A(b[3846]), .B(n1932), .Z(n1933) );
  XNOR U2185 ( .A(b[3846]), .B(n1934), .Z(c[3846]) );
  XNOR U2186 ( .A(a[3846]), .B(n1935), .Z(n1934) );
  IV U2187 ( .A(n1932), .Z(n1935) );
  XOR U2188 ( .A(n1936), .B(n1937), .Z(n1932) );
  ANDN U2189 ( .B(n1938), .A(n1939), .Z(n1936) );
  XNOR U2190 ( .A(b[3845]), .B(n1937), .Z(n1938) );
  XNOR U2191 ( .A(b[3845]), .B(n1939), .Z(c[3845]) );
  XNOR U2192 ( .A(a[3845]), .B(n1940), .Z(n1939) );
  IV U2193 ( .A(n1937), .Z(n1940) );
  XOR U2194 ( .A(n1941), .B(n1942), .Z(n1937) );
  ANDN U2195 ( .B(n1943), .A(n1944), .Z(n1941) );
  XNOR U2196 ( .A(b[3844]), .B(n1942), .Z(n1943) );
  XNOR U2197 ( .A(b[3844]), .B(n1944), .Z(c[3844]) );
  XNOR U2198 ( .A(a[3844]), .B(n1945), .Z(n1944) );
  IV U2199 ( .A(n1942), .Z(n1945) );
  XOR U2200 ( .A(n1946), .B(n1947), .Z(n1942) );
  ANDN U2201 ( .B(n1948), .A(n1949), .Z(n1946) );
  XNOR U2202 ( .A(b[3843]), .B(n1947), .Z(n1948) );
  XNOR U2203 ( .A(b[3843]), .B(n1949), .Z(c[3843]) );
  XNOR U2204 ( .A(a[3843]), .B(n1950), .Z(n1949) );
  IV U2205 ( .A(n1947), .Z(n1950) );
  XOR U2206 ( .A(n1951), .B(n1952), .Z(n1947) );
  ANDN U2207 ( .B(n1953), .A(n1954), .Z(n1951) );
  XNOR U2208 ( .A(b[3842]), .B(n1952), .Z(n1953) );
  XNOR U2209 ( .A(b[3842]), .B(n1954), .Z(c[3842]) );
  XNOR U2210 ( .A(a[3842]), .B(n1955), .Z(n1954) );
  IV U2211 ( .A(n1952), .Z(n1955) );
  XOR U2212 ( .A(n1956), .B(n1957), .Z(n1952) );
  ANDN U2213 ( .B(n1958), .A(n1959), .Z(n1956) );
  XNOR U2214 ( .A(b[3841]), .B(n1957), .Z(n1958) );
  XNOR U2215 ( .A(b[3841]), .B(n1959), .Z(c[3841]) );
  XNOR U2216 ( .A(a[3841]), .B(n1960), .Z(n1959) );
  IV U2217 ( .A(n1957), .Z(n1960) );
  XOR U2218 ( .A(n1961), .B(n1962), .Z(n1957) );
  ANDN U2219 ( .B(n1963), .A(n1964), .Z(n1961) );
  XNOR U2220 ( .A(b[3840]), .B(n1962), .Z(n1963) );
  XNOR U2221 ( .A(b[3840]), .B(n1964), .Z(c[3840]) );
  XNOR U2222 ( .A(a[3840]), .B(n1965), .Z(n1964) );
  IV U2223 ( .A(n1962), .Z(n1965) );
  XOR U2224 ( .A(n1966), .B(n1967), .Z(n1962) );
  ANDN U2225 ( .B(n1968), .A(n1969), .Z(n1966) );
  XNOR U2226 ( .A(b[3839]), .B(n1967), .Z(n1968) );
  XNOR U2227 ( .A(b[383]), .B(n1970), .Z(c[383]) );
  XNOR U2228 ( .A(b[3839]), .B(n1969), .Z(c[3839]) );
  XNOR U2229 ( .A(a[3839]), .B(n1971), .Z(n1969) );
  IV U2230 ( .A(n1967), .Z(n1971) );
  XOR U2231 ( .A(n1972), .B(n1973), .Z(n1967) );
  ANDN U2232 ( .B(n1974), .A(n1975), .Z(n1972) );
  XNOR U2233 ( .A(b[3838]), .B(n1973), .Z(n1974) );
  XNOR U2234 ( .A(b[3838]), .B(n1975), .Z(c[3838]) );
  XNOR U2235 ( .A(a[3838]), .B(n1976), .Z(n1975) );
  IV U2236 ( .A(n1973), .Z(n1976) );
  XOR U2237 ( .A(n1977), .B(n1978), .Z(n1973) );
  ANDN U2238 ( .B(n1979), .A(n1980), .Z(n1977) );
  XNOR U2239 ( .A(b[3837]), .B(n1978), .Z(n1979) );
  XNOR U2240 ( .A(b[3837]), .B(n1980), .Z(c[3837]) );
  XNOR U2241 ( .A(a[3837]), .B(n1981), .Z(n1980) );
  IV U2242 ( .A(n1978), .Z(n1981) );
  XOR U2243 ( .A(n1982), .B(n1983), .Z(n1978) );
  ANDN U2244 ( .B(n1984), .A(n1985), .Z(n1982) );
  XNOR U2245 ( .A(b[3836]), .B(n1983), .Z(n1984) );
  XNOR U2246 ( .A(b[3836]), .B(n1985), .Z(c[3836]) );
  XNOR U2247 ( .A(a[3836]), .B(n1986), .Z(n1985) );
  IV U2248 ( .A(n1983), .Z(n1986) );
  XOR U2249 ( .A(n1987), .B(n1988), .Z(n1983) );
  ANDN U2250 ( .B(n1989), .A(n1990), .Z(n1987) );
  XNOR U2251 ( .A(b[3835]), .B(n1988), .Z(n1989) );
  XNOR U2252 ( .A(b[3835]), .B(n1990), .Z(c[3835]) );
  XNOR U2253 ( .A(a[3835]), .B(n1991), .Z(n1990) );
  IV U2254 ( .A(n1988), .Z(n1991) );
  XOR U2255 ( .A(n1992), .B(n1993), .Z(n1988) );
  ANDN U2256 ( .B(n1994), .A(n1995), .Z(n1992) );
  XNOR U2257 ( .A(b[3834]), .B(n1993), .Z(n1994) );
  XNOR U2258 ( .A(b[3834]), .B(n1995), .Z(c[3834]) );
  XNOR U2259 ( .A(a[3834]), .B(n1996), .Z(n1995) );
  IV U2260 ( .A(n1993), .Z(n1996) );
  XOR U2261 ( .A(n1997), .B(n1998), .Z(n1993) );
  ANDN U2262 ( .B(n1999), .A(n2000), .Z(n1997) );
  XNOR U2263 ( .A(b[3833]), .B(n1998), .Z(n1999) );
  XNOR U2264 ( .A(b[3833]), .B(n2000), .Z(c[3833]) );
  XNOR U2265 ( .A(a[3833]), .B(n2001), .Z(n2000) );
  IV U2266 ( .A(n1998), .Z(n2001) );
  XOR U2267 ( .A(n2002), .B(n2003), .Z(n1998) );
  ANDN U2268 ( .B(n2004), .A(n2005), .Z(n2002) );
  XNOR U2269 ( .A(b[3832]), .B(n2003), .Z(n2004) );
  XNOR U2270 ( .A(b[3832]), .B(n2005), .Z(c[3832]) );
  XNOR U2271 ( .A(a[3832]), .B(n2006), .Z(n2005) );
  IV U2272 ( .A(n2003), .Z(n2006) );
  XOR U2273 ( .A(n2007), .B(n2008), .Z(n2003) );
  ANDN U2274 ( .B(n2009), .A(n2010), .Z(n2007) );
  XNOR U2275 ( .A(b[3831]), .B(n2008), .Z(n2009) );
  XNOR U2276 ( .A(b[3831]), .B(n2010), .Z(c[3831]) );
  XNOR U2277 ( .A(a[3831]), .B(n2011), .Z(n2010) );
  IV U2278 ( .A(n2008), .Z(n2011) );
  XOR U2279 ( .A(n2012), .B(n2013), .Z(n2008) );
  ANDN U2280 ( .B(n2014), .A(n2015), .Z(n2012) );
  XNOR U2281 ( .A(b[3830]), .B(n2013), .Z(n2014) );
  XNOR U2282 ( .A(b[3830]), .B(n2015), .Z(c[3830]) );
  XNOR U2283 ( .A(a[3830]), .B(n2016), .Z(n2015) );
  IV U2284 ( .A(n2013), .Z(n2016) );
  XOR U2285 ( .A(n2017), .B(n2018), .Z(n2013) );
  ANDN U2286 ( .B(n2019), .A(n2020), .Z(n2017) );
  XNOR U2287 ( .A(b[3829]), .B(n2018), .Z(n2019) );
  XNOR U2288 ( .A(b[382]), .B(n2021), .Z(c[382]) );
  XNOR U2289 ( .A(b[3829]), .B(n2020), .Z(c[3829]) );
  XNOR U2290 ( .A(a[3829]), .B(n2022), .Z(n2020) );
  IV U2291 ( .A(n2018), .Z(n2022) );
  XOR U2292 ( .A(n2023), .B(n2024), .Z(n2018) );
  ANDN U2293 ( .B(n2025), .A(n2026), .Z(n2023) );
  XNOR U2294 ( .A(b[3828]), .B(n2024), .Z(n2025) );
  XNOR U2295 ( .A(b[3828]), .B(n2026), .Z(c[3828]) );
  XNOR U2296 ( .A(a[3828]), .B(n2027), .Z(n2026) );
  IV U2297 ( .A(n2024), .Z(n2027) );
  XOR U2298 ( .A(n2028), .B(n2029), .Z(n2024) );
  ANDN U2299 ( .B(n2030), .A(n2031), .Z(n2028) );
  XNOR U2300 ( .A(b[3827]), .B(n2029), .Z(n2030) );
  XNOR U2301 ( .A(b[3827]), .B(n2031), .Z(c[3827]) );
  XNOR U2302 ( .A(a[3827]), .B(n2032), .Z(n2031) );
  IV U2303 ( .A(n2029), .Z(n2032) );
  XOR U2304 ( .A(n2033), .B(n2034), .Z(n2029) );
  ANDN U2305 ( .B(n2035), .A(n2036), .Z(n2033) );
  XNOR U2306 ( .A(b[3826]), .B(n2034), .Z(n2035) );
  XNOR U2307 ( .A(b[3826]), .B(n2036), .Z(c[3826]) );
  XNOR U2308 ( .A(a[3826]), .B(n2037), .Z(n2036) );
  IV U2309 ( .A(n2034), .Z(n2037) );
  XOR U2310 ( .A(n2038), .B(n2039), .Z(n2034) );
  ANDN U2311 ( .B(n2040), .A(n2041), .Z(n2038) );
  XNOR U2312 ( .A(b[3825]), .B(n2039), .Z(n2040) );
  XNOR U2313 ( .A(b[3825]), .B(n2041), .Z(c[3825]) );
  XNOR U2314 ( .A(a[3825]), .B(n2042), .Z(n2041) );
  IV U2315 ( .A(n2039), .Z(n2042) );
  XOR U2316 ( .A(n2043), .B(n2044), .Z(n2039) );
  ANDN U2317 ( .B(n2045), .A(n2046), .Z(n2043) );
  XNOR U2318 ( .A(b[3824]), .B(n2044), .Z(n2045) );
  XNOR U2319 ( .A(b[3824]), .B(n2046), .Z(c[3824]) );
  XNOR U2320 ( .A(a[3824]), .B(n2047), .Z(n2046) );
  IV U2321 ( .A(n2044), .Z(n2047) );
  XOR U2322 ( .A(n2048), .B(n2049), .Z(n2044) );
  ANDN U2323 ( .B(n2050), .A(n2051), .Z(n2048) );
  XNOR U2324 ( .A(b[3823]), .B(n2049), .Z(n2050) );
  XNOR U2325 ( .A(b[3823]), .B(n2051), .Z(c[3823]) );
  XNOR U2326 ( .A(a[3823]), .B(n2052), .Z(n2051) );
  IV U2327 ( .A(n2049), .Z(n2052) );
  XOR U2328 ( .A(n2053), .B(n2054), .Z(n2049) );
  ANDN U2329 ( .B(n2055), .A(n2056), .Z(n2053) );
  XNOR U2330 ( .A(b[3822]), .B(n2054), .Z(n2055) );
  XNOR U2331 ( .A(b[3822]), .B(n2056), .Z(c[3822]) );
  XNOR U2332 ( .A(a[3822]), .B(n2057), .Z(n2056) );
  IV U2333 ( .A(n2054), .Z(n2057) );
  XOR U2334 ( .A(n2058), .B(n2059), .Z(n2054) );
  ANDN U2335 ( .B(n2060), .A(n2061), .Z(n2058) );
  XNOR U2336 ( .A(b[3821]), .B(n2059), .Z(n2060) );
  XNOR U2337 ( .A(b[3821]), .B(n2061), .Z(c[3821]) );
  XNOR U2338 ( .A(a[3821]), .B(n2062), .Z(n2061) );
  IV U2339 ( .A(n2059), .Z(n2062) );
  XOR U2340 ( .A(n2063), .B(n2064), .Z(n2059) );
  ANDN U2341 ( .B(n2065), .A(n2066), .Z(n2063) );
  XNOR U2342 ( .A(b[3820]), .B(n2064), .Z(n2065) );
  XNOR U2343 ( .A(b[3820]), .B(n2066), .Z(c[3820]) );
  XNOR U2344 ( .A(a[3820]), .B(n2067), .Z(n2066) );
  IV U2345 ( .A(n2064), .Z(n2067) );
  XOR U2346 ( .A(n2068), .B(n2069), .Z(n2064) );
  ANDN U2347 ( .B(n2070), .A(n2071), .Z(n2068) );
  XNOR U2348 ( .A(b[3819]), .B(n2069), .Z(n2070) );
  XNOR U2349 ( .A(b[381]), .B(n2072), .Z(c[381]) );
  XNOR U2350 ( .A(b[3819]), .B(n2071), .Z(c[3819]) );
  XNOR U2351 ( .A(a[3819]), .B(n2073), .Z(n2071) );
  IV U2352 ( .A(n2069), .Z(n2073) );
  XOR U2353 ( .A(n2074), .B(n2075), .Z(n2069) );
  ANDN U2354 ( .B(n2076), .A(n2077), .Z(n2074) );
  XNOR U2355 ( .A(b[3818]), .B(n2075), .Z(n2076) );
  XNOR U2356 ( .A(b[3818]), .B(n2077), .Z(c[3818]) );
  XNOR U2357 ( .A(a[3818]), .B(n2078), .Z(n2077) );
  IV U2358 ( .A(n2075), .Z(n2078) );
  XOR U2359 ( .A(n2079), .B(n2080), .Z(n2075) );
  ANDN U2360 ( .B(n2081), .A(n2082), .Z(n2079) );
  XNOR U2361 ( .A(b[3817]), .B(n2080), .Z(n2081) );
  XNOR U2362 ( .A(b[3817]), .B(n2082), .Z(c[3817]) );
  XNOR U2363 ( .A(a[3817]), .B(n2083), .Z(n2082) );
  IV U2364 ( .A(n2080), .Z(n2083) );
  XOR U2365 ( .A(n2084), .B(n2085), .Z(n2080) );
  ANDN U2366 ( .B(n2086), .A(n2087), .Z(n2084) );
  XNOR U2367 ( .A(b[3816]), .B(n2085), .Z(n2086) );
  XNOR U2368 ( .A(b[3816]), .B(n2087), .Z(c[3816]) );
  XNOR U2369 ( .A(a[3816]), .B(n2088), .Z(n2087) );
  IV U2370 ( .A(n2085), .Z(n2088) );
  XOR U2371 ( .A(n2089), .B(n2090), .Z(n2085) );
  ANDN U2372 ( .B(n2091), .A(n2092), .Z(n2089) );
  XNOR U2373 ( .A(b[3815]), .B(n2090), .Z(n2091) );
  XNOR U2374 ( .A(b[3815]), .B(n2092), .Z(c[3815]) );
  XNOR U2375 ( .A(a[3815]), .B(n2093), .Z(n2092) );
  IV U2376 ( .A(n2090), .Z(n2093) );
  XOR U2377 ( .A(n2094), .B(n2095), .Z(n2090) );
  ANDN U2378 ( .B(n2096), .A(n2097), .Z(n2094) );
  XNOR U2379 ( .A(b[3814]), .B(n2095), .Z(n2096) );
  XNOR U2380 ( .A(b[3814]), .B(n2097), .Z(c[3814]) );
  XNOR U2381 ( .A(a[3814]), .B(n2098), .Z(n2097) );
  IV U2382 ( .A(n2095), .Z(n2098) );
  XOR U2383 ( .A(n2099), .B(n2100), .Z(n2095) );
  ANDN U2384 ( .B(n2101), .A(n2102), .Z(n2099) );
  XNOR U2385 ( .A(b[3813]), .B(n2100), .Z(n2101) );
  XNOR U2386 ( .A(b[3813]), .B(n2102), .Z(c[3813]) );
  XNOR U2387 ( .A(a[3813]), .B(n2103), .Z(n2102) );
  IV U2388 ( .A(n2100), .Z(n2103) );
  XOR U2389 ( .A(n2104), .B(n2105), .Z(n2100) );
  ANDN U2390 ( .B(n2106), .A(n2107), .Z(n2104) );
  XNOR U2391 ( .A(b[3812]), .B(n2105), .Z(n2106) );
  XNOR U2392 ( .A(b[3812]), .B(n2107), .Z(c[3812]) );
  XNOR U2393 ( .A(a[3812]), .B(n2108), .Z(n2107) );
  IV U2394 ( .A(n2105), .Z(n2108) );
  XOR U2395 ( .A(n2109), .B(n2110), .Z(n2105) );
  ANDN U2396 ( .B(n2111), .A(n2112), .Z(n2109) );
  XNOR U2397 ( .A(b[3811]), .B(n2110), .Z(n2111) );
  XNOR U2398 ( .A(b[3811]), .B(n2112), .Z(c[3811]) );
  XNOR U2399 ( .A(a[3811]), .B(n2113), .Z(n2112) );
  IV U2400 ( .A(n2110), .Z(n2113) );
  XOR U2401 ( .A(n2114), .B(n2115), .Z(n2110) );
  ANDN U2402 ( .B(n2116), .A(n2117), .Z(n2114) );
  XNOR U2403 ( .A(b[3810]), .B(n2115), .Z(n2116) );
  XNOR U2404 ( .A(b[3810]), .B(n2117), .Z(c[3810]) );
  XNOR U2405 ( .A(a[3810]), .B(n2118), .Z(n2117) );
  IV U2406 ( .A(n2115), .Z(n2118) );
  XOR U2407 ( .A(n2119), .B(n2120), .Z(n2115) );
  ANDN U2408 ( .B(n2121), .A(n2122), .Z(n2119) );
  XNOR U2409 ( .A(b[3809]), .B(n2120), .Z(n2121) );
  XNOR U2410 ( .A(b[380]), .B(n2123), .Z(c[380]) );
  XNOR U2411 ( .A(b[3809]), .B(n2122), .Z(c[3809]) );
  XNOR U2412 ( .A(a[3809]), .B(n2124), .Z(n2122) );
  IV U2413 ( .A(n2120), .Z(n2124) );
  XOR U2414 ( .A(n2125), .B(n2126), .Z(n2120) );
  ANDN U2415 ( .B(n2127), .A(n2128), .Z(n2125) );
  XNOR U2416 ( .A(b[3808]), .B(n2126), .Z(n2127) );
  XNOR U2417 ( .A(b[3808]), .B(n2128), .Z(c[3808]) );
  XNOR U2418 ( .A(a[3808]), .B(n2129), .Z(n2128) );
  IV U2419 ( .A(n2126), .Z(n2129) );
  XOR U2420 ( .A(n2130), .B(n2131), .Z(n2126) );
  ANDN U2421 ( .B(n2132), .A(n2133), .Z(n2130) );
  XNOR U2422 ( .A(b[3807]), .B(n2131), .Z(n2132) );
  XNOR U2423 ( .A(b[3807]), .B(n2133), .Z(c[3807]) );
  XNOR U2424 ( .A(a[3807]), .B(n2134), .Z(n2133) );
  IV U2425 ( .A(n2131), .Z(n2134) );
  XOR U2426 ( .A(n2135), .B(n2136), .Z(n2131) );
  ANDN U2427 ( .B(n2137), .A(n2138), .Z(n2135) );
  XNOR U2428 ( .A(b[3806]), .B(n2136), .Z(n2137) );
  XNOR U2429 ( .A(b[3806]), .B(n2138), .Z(c[3806]) );
  XNOR U2430 ( .A(a[3806]), .B(n2139), .Z(n2138) );
  IV U2431 ( .A(n2136), .Z(n2139) );
  XOR U2432 ( .A(n2140), .B(n2141), .Z(n2136) );
  ANDN U2433 ( .B(n2142), .A(n2143), .Z(n2140) );
  XNOR U2434 ( .A(b[3805]), .B(n2141), .Z(n2142) );
  XNOR U2435 ( .A(b[3805]), .B(n2143), .Z(c[3805]) );
  XNOR U2436 ( .A(a[3805]), .B(n2144), .Z(n2143) );
  IV U2437 ( .A(n2141), .Z(n2144) );
  XOR U2438 ( .A(n2145), .B(n2146), .Z(n2141) );
  ANDN U2439 ( .B(n2147), .A(n2148), .Z(n2145) );
  XNOR U2440 ( .A(b[3804]), .B(n2146), .Z(n2147) );
  XNOR U2441 ( .A(b[3804]), .B(n2148), .Z(c[3804]) );
  XNOR U2442 ( .A(a[3804]), .B(n2149), .Z(n2148) );
  IV U2443 ( .A(n2146), .Z(n2149) );
  XOR U2444 ( .A(n2150), .B(n2151), .Z(n2146) );
  ANDN U2445 ( .B(n2152), .A(n2153), .Z(n2150) );
  XNOR U2446 ( .A(b[3803]), .B(n2151), .Z(n2152) );
  XNOR U2447 ( .A(b[3803]), .B(n2153), .Z(c[3803]) );
  XNOR U2448 ( .A(a[3803]), .B(n2154), .Z(n2153) );
  IV U2449 ( .A(n2151), .Z(n2154) );
  XOR U2450 ( .A(n2155), .B(n2156), .Z(n2151) );
  ANDN U2451 ( .B(n2157), .A(n2158), .Z(n2155) );
  XNOR U2452 ( .A(b[3802]), .B(n2156), .Z(n2157) );
  XNOR U2453 ( .A(b[3802]), .B(n2158), .Z(c[3802]) );
  XNOR U2454 ( .A(a[3802]), .B(n2159), .Z(n2158) );
  IV U2455 ( .A(n2156), .Z(n2159) );
  XOR U2456 ( .A(n2160), .B(n2161), .Z(n2156) );
  ANDN U2457 ( .B(n2162), .A(n2163), .Z(n2160) );
  XNOR U2458 ( .A(b[3801]), .B(n2161), .Z(n2162) );
  XNOR U2459 ( .A(b[3801]), .B(n2163), .Z(c[3801]) );
  XNOR U2460 ( .A(a[3801]), .B(n2164), .Z(n2163) );
  IV U2461 ( .A(n2161), .Z(n2164) );
  XOR U2462 ( .A(n2165), .B(n2166), .Z(n2161) );
  ANDN U2463 ( .B(n2167), .A(n2168), .Z(n2165) );
  XNOR U2464 ( .A(b[3800]), .B(n2166), .Z(n2167) );
  XNOR U2465 ( .A(b[3800]), .B(n2168), .Z(c[3800]) );
  XNOR U2466 ( .A(a[3800]), .B(n2169), .Z(n2168) );
  IV U2467 ( .A(n2166), .Z(n2169) );
  XOR U2468 ( .A(n2170), .B(n2171), .Z(n2166) );
  ANDN U2469 ( .B(n2172), .A(n2173), .Z(n2170) );
  XNOR U2470 ( .A(b[3799]), .B(n2171), .Z(n2172) );
  XNOR U2471 ( .A(b[37]), .B(n2174), .Z(c[37]) );
  XNOR U2472 ( .A(b[379]), .B(n2175), .Z(c[379]) );
  XNOR U2473 ( .A(b[3799]), .B(n2173), .Z(c[3799]) );
  XNOR U2474 ( .A(a[3799]), .B(n2176), .Z(n2173) );
  IV U2475 ( .A(n2171), .Z(n2176) );
  XOR U2476 ( .A(n2177), .B(n2178), .Z(n2171) );
  ANDN U2477 ( .B(n2179), .A(n2180), .Z(n2177) );
  XNOR U2478 ( .A(b[3798]), .B(n2178), .Z(n2179) );
  XNOR U2479 ( .A(b[3798]), .B(n2180), .Z(c[3798]) );
  XNOR U2480 ( .A(a[3798]), .B(n2181), .Z(n2180) );
  IV U2481 ( .A(n2178), .Z(n2181) );
  XOR U2482 ( .A(n2182), .B(n2183), .Z(n2178) );
  ANDN U2483 ( .B(n2184), .A(n2185), .Z(n2182) );
  XNOR U2484 ( .A(b[3797]), .B(n2183), .Z(n2184) );
  XNOR U2485 ( .A(b[3797]), .B(n2185), .Z(c[3797]) );
  XNOR U2486 ( .A(a[3797]), .B(n2186), .Z(n2185) );
  IV U2487 ( .A(n2183), .Z(n2186) );
  XOR U2488 ( .A(n2187), .B(n2188), .Z(n2183) );
  ANDN U2489 ( .B(n2189), .A(n2190), .Z(n2187) );
  XNOR U2490 ( .A(b[3796]), .B(n2188), .Z(n2189) );
  XNOR U2491 ( .A(b[3796]), .B(n2190), .Z(c[3796]) );
  XNOR U2492 ( .A(a[3796]), .B(n2191), .Z(n2190) );
  IV U2493 ( .A(n2188), .Z(n2191) );
  XOR U2494 ( .A(n2192), .B(n2193), .Z(n2188) );
  ANDN U2495 ( .B(n2194), .A(n2195), .Z(n2192) );
  XNOR U2496 ( .A(b[3795]), .B(n2193), .Z(n2194) );
  XNOR U2497 ( .A(b[3795]), .B(n2195), .Z(c[3795]) );
  XNOR U2498 ( .A(a[3795]), .B(n2196), .Z(n2195) );
  IV U2499 ( .A(n2193), .Z(n2196) );
  XOR U2500 ( .A(n2197), .B(n2198), .Z(n2193) );
  ANDN U2501 ( .B(n2199), .A(n2200), .Z(n2197) );
  XNOR U2502 ( .A(b[3794]), .B(n2198), .Z(n2199) );
  XNOR U2503 ( .A(b[3794]), .B(n2200), .Z(c[3794]) );
  XNOR U2504 ( .A(a[3794]), .B(n2201), .Z(n2200) );
  IV U2505 ( .A(n2198), .Z(n2201) );
  XOR U2506 ( .A(n2202), .B(n2203), .Z(n2198) );
  ANDN U2507 ( .B(n2204), .A(n2205), .Z(n2202) );
  XNOR U2508 ( .A(b[3793]), .B(n2203), .Z(n2204) );
  XNOR U2509 ( .A(b[3793]), .B(n2205), .Z(c[3793]) );
  XNOR U2510 ( .A(a[3793]), .B(n2206), .Z(n2205) );
  IV U2511 ( .A(n2203), .Z(n2206) );
  XOR U2512 ( .A(n2207), .B(n2208), .Z(n2203) );
  ANDN U2513 ( .B(n2209), .A(n2210), .Z(n2207) );
  XNOR U2514 ( .A(b[3792]), .B(n2208), .Z(n2209) );
  XNOR U2515 ( .A(b[3792]), .B(n2210), .Z(c[3792]) );
  XNOR U2516 ( .A(a[3792]), .B(n2211), .Z(n2210) );
  IV U2517 ( .A(n2208), .Z(n2211) );
  XOR U2518 ( .A(n2212), .B(n2213), .Z(n2208) );
  ANDN U2519 ( .B(n2214), .A(n2215), .Z(n2212) );
  XNOR U2520 ( .A(b[3791]), .B(n2213), .Z(n2214) );
  XNOR U2521 ( .A(b[3791]), .B(n2215), .Z(c[3791]) );
  XNOR U2522 ( .A(a[3791]), .B(n2216), .Z(n2215) );
  IV U2523 ( .A(n2213), .Z(n2216) );
  XOR U2524 ( .A(n2217), .B(n2218), .Z(n2213) );
  ANDN U2525 ( .B(n2219), .A(n2220), .Z(n2217) );
  XNOR U2526 ( .A(b[3790]), .B(n2218), .Z(n2219) );
  XNOR U2527 ( .A(b[3790]), .B(n2220), .Z(c[3790]) );
  XNOR U2528 ( .A(a[3790]), .B(n2221), .Z(n2220) );
  IV U2529 ( .A(n2218), .Z(n2221) );
  XOR U2530 ( .A(n2222), .B(n2223), .Z(n2218) );
  ANDN U2531 ( .B(n2224), .A(n2225), .Z(n2222) );
  XNOR U2532 ( .A(b[3789]), .B(n2223), .Z(n2224) );
  XNOR U2533 ( .A(b[378]), .B(n2226), .Z(c[378]) );
  XNOR U2534 ( .A(b[3789]), .B(n2225), .Z(c[3789]) );
  XNOR U2535 ( .A(a[3789]), .B(n2227), .Z(n2225) );
  IV U2536 ( .A(n2223), .Z(n2227) );
  XOR U2537 ( .A(n2228), .B(n2229), .Z(n2223) );
  ANDN U2538 ( .B(n2230), .A(n2231), .Z(n2228) );
  XNOR U2539 ( .A(b[3788]), .B(n2229), .Z(n2230) );
  XNOR U2540 ( .A(b[3788]), .B(n2231), .Z(c[3788]) );
  XNOR U2541 ( .A(a[3788]), .B(n2232), .Z(n2231) );
  IV U2542 ( .A(n2229), .Z(n2232) );
  XOR U2543 ( .A(n2233), .B(n2234), .Z(n2229) );
  ANDN U2544 ( .B(n2235), .A(n2236), .Z(n2233) );
  XNOR U2545 ( .A(b[3787]), .B(n2234), .Z(n2235) );
  XNOR U2546 ( .A(b[3787]), .B(n2236), .Z(c[3787]) );
  XNOR U2547 ( .A(a[3787]), .B(n2237), .Z(n2236) );
  IV U2548 ( .A(n2234), .Z(n2237) );
  XOR U2549 ( .A(n2238), .B(n2239), .Z(n2234) );
  ANDN U2550 ( .B(n2240), .A(n2241), .Z(n2238) );
  XNOR U2551 ( .A(b[3786]), .B(n2239), .Z(n2240) );
  XNOR U2552 ( .A(b[3786]), .B(n2241), .Z(c[3786]) );
  XNOR U2553 ( .A(a[3786]), .B(n2242), .Z(n2241) );
  IV U2554 ( .A(n2239), .Z(n2242) );
  XOR U2555 ( .A(n2243), .B(n2244), .Z(n2239) );
  ANDN U2556 ( .B(n2245), .A(n2246), .Z(n2243) );
  XNOR U2557 ( .A(b[3785]), .B(n2244), .Z(n2245) );
  XNOR U2558 ( .A(b[3785]), .B(n2246), .Z(c[3785]) );
  XNOR U2559 ( .A(a[3785]), .B(n2247), .Z(n2246) );
  IV U2560 ( .A(n2244), .Z(n2247) );
  XOR U2561 ( .A(n2248), .B(n2249), .Z(n2244) );
  ANDN U2562 ( .B(n2250), .A(n2251), .Z(n2248) );
  XNOR U2563 ( .A(b[3784]), .B(n2249), .Z(n2250) );
  XNOR U2564 ( .A(b[3784]), .B(n2251), .Z(c[3784]) );
  XNOR U2565 ( .A(a[3784]), .B(n2252), .Z(n2251) );
  IV U2566 ( .A(n2249), .Z(n2252) );
  XOR U2567 ( .A(n2253), .B(n2254), .Z(n2249) );
  ANDN U2568 ( .B(n2255), .A(n2256), .Z(n2253) );
  XNOR U2569 ( .A(b[3783]), .B(n2254), .Z(n2255) );
  XNOR U2570 ( .A(b[3783]), .B(n2256), .Z(c[3783]) );
  XNOR U2571 ( .A(a[3783]), .B(n2257), .Z(n2256) );
  IV U2572 ( .A(n2254), .Z(n2257) );
  XOR U2573 ( .A(n2258), .B(n2259), .Z(n2254) );
  ANDN U2574 ( .B(n2260), .A(n2261), .Z(n2258) );
  XNOR U2575 ( .A(b[3782]), .B(n2259), .Z(n2260) );
  XNOR U2576 ( .A(b[3782]), .B(n2261), .Z(c[3782]) );
  XNOR U2577 ( .A(a[3782]), .B(n2262), .Z(n2261) );
  IV U2578 ( .A(n2259), .Z(n2262) );
  XOR U2579 ( .A(n2263), .B(n2264), .Z(n2259) );
  ANDN U2580 ( .B(n2265), .A(n2266), .Z(n2263) );
  XNOR U2581 ( .A(b[3781]), .B(n2264), .Z(n2265) );
  XNOR U2582 ( .A(b[3781]), .B(n2266), .Z(c[3781]) );
  XNOR U2583 ( .A(a[3781]), .B(n2267), .Z(n2266) );
  IV U2584 ( .A(n2264), .Z(n2267) );
  XOR U2585 ( .A(n2268), .B(n2269), .Z(n2264) );
  ANDN U2586 ( .B(n2270), .A(n2271), .Z(n2268) );
  XNOR U2587 ( .A(b[3780]), .B(n2269), .Z(n2270) );
  XNOR U2588 ( .A(b[3780]), .B(n2271), .Z(c[3780]) );
  XNOR U2589 ( .A(a[3780]), .B(n2272), .Z(n2271) );
  IV U2590 ( .A(n2269), .Z(n2272) );
  XOR U2591 ( .A(n2273), .B(n2274), .Z(n2269) );
  ANDN U2592 ( .B(n2275), .A(n2276), .Z(n2273) );
  XNOR U2593 ( .A(b[3779]), .B(n2274), .Z(n2275) );
  XNOR U2594 ( .A(b[377]), .B(n2277), .Z(c[377]) );
  XNOR U2595 ( .A(b[3779]), .B(n2276), .Z(c[3779]) );
  XNOR U2596 ( .A(a[3779]), .B(n2278), .Z(n2276) );
  IV U2597 ( .A(n2274), .Z(n2278) );
  XOR U2598 ( .A(n2279), .B(n2280), .Z(n2274) );
  ANDN U2599 ( .B(n2281), .A(n2282), .Z(n2279) );
  XNOR U2600 ( .A(b[3778]), .B(n2280), .Z(n2281) );
  XNOR U2601 ( .A(b[3778]), .B(n2282), .Z(c[3778]) );
  XNOR U2602 ( .A(a[3778]), .B(n2283), .Z(n2282) );
  IV U2603 ( .A(n2280), .Z(n2283) );
  XOR U2604 ( .A(n2284), .B(n2285), .Z(n2280) );
  ANDN U2605 ( .B(n2286), .A(n2287), .Z(n2284) );
  XNOR U2606 ( .A(b[3777]), .B(n2285), .Z(n2286) );
  XNOR U2607 ( .A(b[3777]), .B(n2287), .Z(c[3777]) );
  XNOR U2608 ( .A(a[3777]), .B(n2288), .Z(n2287) );
  IV U2609 ( .A(n2285), .Z(n2288) );
  XOR U2610 ( .A(n2289), .B(n2290), .Z(n2285) );
  ANDN U2611 ( .B(n2291), .A(n2292), .Z(n2289) );
  XNOR U2612 ( .A(b[3776]), .B(n2290), .Z(n2291) );
  XNOR U2613 ( .A(b[3776]), .B(n2292), .Z(c[3776]) );
  XNOR U2614 ( .A(a[3776]), .B(n2293), .Z(n2292) );
  IV U2615 ( .A(n2290), .Z(n2293) );
  XOR U2616 ( .A(n2294), .B(n2295), .Z(n2290) );
  ANDN U2617 ( .B(n2296), .A(n2297), .Z(n2294) );
  XNOR U2618 ( .A(b[3775]), .B(n2295), .Z(n2296) );
  XNOR U2619 ( .A(b[3775]), .B(n2297), .Z(c[3775]) );
  XNOR U2620 ( .A(a[3775]), .B(n2298), .Z(n2297) );
  IV U2621 ( .A(n2295), .Z(n2298) );
  XOR U2622 ( .A(n2299), .B(n2300), .Z(n2295) );
  ANDN U2623 ( .B(n2301), .A(n2302), .Z(n2299) );
  XNOR U2624 ( .A(b[3774]), .B(n2300), .Z(n2301) );
  XNOR U2625 ( .A(b[3774]), .B(n2302), .Z(c[3774]) );
  XNOR U2626 ( .A(a[3774]), .B(n2303), .Z(n2302) );
  IV U2627 ( .A(n2300), .Z(n2303) );
  XOR U2628 ( .A(n2304), .B(n2305), .Z(n2300) );
  ANDN U2629 ( .B(n2306), .A(n2307), .Z(n2304) );
  XNOR U2630 ( .A(b[3773]), .B(n2305), .Z(n2306) );
  XNOR U2631 ( .A(b[3773]), .B(n2307), .Z(c[3773]) );
  XNOR U2632 ( .A(a[3773]), .B(n2308), .Z(n2307) );
  IV U2633 ( .A(n2305), .Z(n2308) );
  XOR U2634 ( .A(n2309), .B(n2310), .Z(n2305) );
  ANDN U2635 ( .B(n2311), .A(n2312), .Z(n2309) );
  XNOR U2636 ( .A(b[3772]), .B(n2310), .Z(n2311) );
  XNOR U2637 ( .A(b[3772]), .B(n2312), .Z(c[3772]) );
  XNOR U2638 ( .A(a[3772]), .B(n2313), .Z(n2312) );
  IV U2639 ( .A(n2310), .Z(n2313) );
  XOR U2640 ( .A(n2314), .B(n2315), .Z(n2310) );
  ANDN U2641 ( .B(n2316), .A(n2317), .Z(n2314) );
  XNOR U2642 ( .A(b[3771]), .B(n2315), .Z(n2316) );
  XNOR U2643 ( .A(b[3771]), .B(n2317), .Z(c[3771]) );
  XNOR U2644 ( .A(a[3771]), .B(n2318), .Z(n2317) );
  IV U2645 ( .A(n2315), .Z(n2318) );
  XOR U2646 ( .A(n2319), .B(n2320), .Z(n2315) );
  ANDN U2647 ( .B(n2321), .A(n2322), .Z(n2319) );
  XNOR U2648 ( .A(b[3770]), .B(n2320), .Z(n2321) );
  XNOR U2649 ( .A(b[3770]), .B(n2322), .Z(c[3770]) );
  XNOR U2650 ( .A(a[3770]), .B(n2323), .Z(n2322) );
  IV U2651 ( .A(n2320), .Z(n2323) );
  XOR U2652 ( .A(n2324), .B(n2325), .Z(n2320) );
  ANDN U2653 ( .B(n2326), .A(n2327), .Z(n2324) );
  XNOR U2654 ( .A(b[3769]), .B(n2325), .Z(n2326) );
  XNOR U2655 ( .A(b[376]), .B(n2328), .Z(c[376]) );
  XNOR U2656 ( .A(b[3769]), .B(n2327), .Z(c[3769]) );
  XNOR U2657 ( .A(a[3769]), .B(n2329), .Z(n2327) );
  IV U2658 ( .A(n2325), .Z(n2329) );
  XOR U2659 ( .A(n2330), .B(n2331), .Z(n2325) );
  ANDN U2660 ( .B(n2332), .A(n2333), .Z(n2330) );
  XNOR U2661 ( .A(b[3768]), .B(n2331), .Z(n2332) );
  XNOR U2662 ( .A(b[3768]), .B(n2333), .Z(c[3768]) );
  XNOR U2663 ( .A(a[3768]), .B(n2334), .Z(n2333) );
  IV U2664 ( .A(n2331), .Z(n2334) );
  XOR U2665 ( .A(n2335), .B(n2336), .Z(n2331) );
  ANDN U2666 ( .B(n2337), .A(n2338), .Z(n2335) );
  XNOR U2667 ( .A(b[3767]), .B(n2336), .Z(n2337) );
  XNOR U2668 ( .A(b[3767]), .B(n2338), .Z(c[3767]) );
  XNOR U2669 ( .A(a[3767]), .B(n2339), .Z(n2338) );
  IV U2670 ( .A(n2336), .Z(n2339) );
  XOR U2671 ( .A(n2340), .B(n2341), .Z(n2336) );
  ANDN U2672 ( .B(n2342), .A(n2343), .Z(n2340) );
  XNOR U2673 ( .A(b[3766]), .B(n2341), .Z(n2342) );
  XNOR U2674 ( .A(b[3766]), .B(n2343), .Z(c[3766]) );
  XNOR U2675 ( .A(a[3766]), .B(n2344), .Z(n2343) );
  IV U2676 ( .A(n2341), .Z(n2344) );
  XOR U2677 ( .A(n2345), .B(n2346), .Z(n2341) );
  ANDN U2678 ( .B(n2347), .A(n2348), .Z(n2345) );
  XNOR U2679 ( .A(b[3765]), .B(n2346), .Z(n2347) );
  XNOR U2680 ( .A(b[3765]), .B(n2348), .Z(c[3765]) );
  XNOR U2681 ( .A(a[3765]), .B(n2349), .Z(n2348) );
  IV U2682 ( .A(n2346), .Z(n2349) );
  XOR U2683 ( .A(n2350), .B(n2351), .Z(n2346) );
  ANDN U2684 ( .B(n2352), .A(n2353), .Z(n2350) );
  XNOR U2685 ( .A(b[3764]), .B(n2351), .Z(n2352) );
  XNOR U2686 ( .A(b[3764]), .B(n2353), .Z(c[3764]) );
  XNOR U2687 ( .A(a[3764]), .B(n2354), .Z(n2353) );
  IV U2688 ( .A(n2351), .Z(n2354) );
  XOR U2689 ( .A(n2355), .B(n2356), .Z(n2351) );
  ANDN U2690 ( .B(n2357), .A(n2358), .Z(n2355) );
  XNOR U2691 ( .A(b[3763]), .B(n2356), .Z(n2357) );
  XNOR U2692 ( .A(b[3763]), .B(n2358), .Z(c[3763]) );
  XNOR U2693 ( .A(a[3763]), .B(n2359), .Z(n2358) );
  IV U2694 ( .A(n2356), .Z(n2359) );
  XOR U2695 ( .A(n2360), .B(n2361), .Z(n2356) );
  ANDN U2696 ( .B(n2362), .A(n2363), .Z(n2360) );
  XNOR U2697 ( .A(b[3762]), .B(n2361), .Z(n2362) );
  XNOR U2698 ( .A(b[3762]), .B(n2363), .Z(c[3762]) );
  XNOR U2699 ( .A(a[3762]), .B(n2364), .Z(n2363) );
  IV U2700 ( .A(n2361), .Z(n2364) );
  XOR U2701 ( .A(n2365), .B(n2366), .Z(n2361) );
  ANDN U2702 ( .B(n2367), .A(n2368), .Z(n2365) );
  XNOR U2703 ( .A(b[3761]), .B(n2366), .Z(n2367) );
  XNOR U2704 ( .A(b[3761]), .B(n2368), .Z(c[3761]) );
  XNOR U2705 ( .A(a[3761]), .B(n2369), .Z(n2368) );
  IV U2706 ( .A(n2366), .Z(n2369) );
  XOR U2707 ( .A(n2370), .B(n2371), .Z(n2366) );
  ANDN U2708 ( .B(n2372), .A(n2373), .Z(n2370) );
  XNOR U2709 ( .A(b[3760]), .B(n2371), .Z(n2372) );
  XNOR U2710 ( .A(b[3760]), .B(n2373), .Z(c[3760]) );
  XNOR U2711 ( .A(a[3760]), .B(n2374), .Z(n2373) );
  IV U2712 ( .A(n2371), .Z(n2374) );
  XOR U2713 ( .A(n2375), .B(n2376), .Z(n2371) );
  ANDN U2714 ( .B(n2377), .A(n2378), .Z(n2375) );
  XNOR U2715 ( .A(b[3759]), .B(n2376), .Z(n2377) );
  XNOR U2716 ( .A(b[375]), .B(n2379), .Z(c[375]) );
  XNOR U2717 ( .A(b[3759]), .B(n2378), .Z(c[3759]) );
  XNOR U2718 ( .A(a[3759]), .B(n2380), .Z(n2378) );
  IV U2719 ( .A(n2376), .Z(n2380) );
  XOR U2720 ( .A(n2381), .B(n2382), .Z(n2376) );
  ANDN U2721 ( .B(n2383), .A(n2384), .Z(n2381) );
  XNOR U2722 ( .A(b[3758]), .B(n2382), .Z(n2383) );
  XNOR U2723 ( .A(b[3758]), .B(n2384), .Z(c[3758]) );
  XNOR U2724 ( .A(a[3758]), .B(n2385), .Z(n2384) );
  IV U2725 ( .A(n2382), .Z(n2385) );
  XOR U2726 ( .A(n2386), .B(n2387), .Z(n2382) );
  ANDN U2727 ( .B(n2388), .A(n2389), .Z(n2386) );
  XNOR U2728 ( .A(b[3757]), .B(n2387), .Z(n2388) );
  XNOR U2729 ( .A(b[3757]), .B(n2389), .Z(c[3757]) );
  XNOR U2730 ( .A(a[3757]), .B(n2390), .Z(n2389) );
  IV U2731 ( .A(n2387), .Z(n2390) );
  XOR U2732 ( .A(n2391), .B(n2392), .Z(n2387) );
  ANDN U2733 ( .B(n2393), .A(n2394), .Z(n2391) );
  XNOR U2734 ( .A(b[3756]), .B(n2392), .Z(n2393) );
  XNOR U2735 ( .A(b[3756]), .B(n2394), .Z(c[3756]) );
  XNOR U2736 ( .A(a[3756]), .B(n2395), .Z(n2394) );
  IV U2737 ( .A(n2392), .Z(n2395) );
  XOR U2738 ( .A(n2396), .B(n2397), .Z(n2392) );
  ANDN U2739 ( .B(n2398), .A(n2399), .Z(n2396) );
  XNOR U2740 ( .A(b[3755]), .B(n2397), .Z(n2398) );
  XNOR U2741 ( .A(b[3755]), .B(n2399), .Z(c[3755]) );
  XNOR U2742 ( .A(a[3755]), .B(n2400), .Z(n2399) );
  IV U2743 ( .A(n2397), .Z(n2400) );
  XOR U2744 ( .A(n2401), .B(n2402), .Z(n2397) );
  ANDN U2745 ( .B(n2403), .A(n2404), .Z(n2401) );
  XNOR U2746 ( .A(b[3754]), .B(n2402), .Z(n2403) );
  XNOR U2747 ( .A(b[3754]), .B(n2404), .Z(c[3754]) );
  XNOR U2748 ( .A(a[3754]), .B(n2405), .Z(n2404) );
  IV U2749 ( .A(n2402), .Z(n2405) );
  XOR U2750 ( .A(n2406), .B(n2407), .Z(n2402) );
  ANDN U2751 ( .B(n2408), .A(n2409), .Z(n2406) );
  XNOR U2752 ( .A(b[3753]), .B(n2407), .Z(n2408) );
  XNOR U2753 ( .A(b[3753]), .B(n2409), .Z(c[3753]) );
  XNOR U2754 ( .A(a[3753]), .B(n2410), .Z(n2409) );
  IV U2755 ( .A(n2407), .Z(n2410) );
  XOR U2756 ( .A(n2411), .B(n2412), .Z(n2407) );
  ANDN U2757 ( .B(n2413), .A(n2414), .Z(n2411) );
  XNOR U2758 ( .A(b[3752]), .B(n2412), .Z(n2413) );
  XNOR U2759 ( .A(b[3752]), .B(n2414), .Z(c[3752]) );
  XNOR U2760 ( .A(a[3752]), .B(n2415), .Z(n2414) );
  IV U2761 ( .A(n2412), .Z(n2415) );
  XOR U2762 ( .A(n2416), .B(n2417), .Z(n2412) );
  ANDN U2763 ( .B(n2418), .A(n2419), .Z(n2416) );
  XNOR U2764 ( .A(b[3751]), .B(n2417), .Z(n2418) );
  XNOR U2765 ( .A(b[3751]), .B(n2419), .Z(c[3751]) );
  XNOR U2766 ( .A(a[3751]), .B(n2420), .Z(n2419) );
  IV U2767 ( .A(n2417), .Z(n2420) );
  XOR U2768 ( .A(n2421), .B(n2422), .Z(n2417) );
  ANDN U2769 ( .B(n2423), .A(n2424), .Z(n2421) );
  XNOR U2770 ( .A(b[3750]), .B(n2422), .Z(n2423) );
  XNOR U2771 ( .A(b[3750]), .B(n2424), .Z(c[3750]) );
  XNOR U2772 ( .A(a[3750]), .B(n2425), .Z(n2424) );
  IV U2773 ( .A(n2422), .Z(n2425) );
  XOR U2774 ( .A(n2426), .B(n2427), .Z(n2422) );
  ANDN U2775 ( .B(n2428), .A(n2429), .Z(n2426) );
  XNOR U2776 ( .A(b[3749]), .B(n2427), .Z(n2428) );
  XNOR U2777 ( .A(b[374]), .B(n2430), .Z(c[374]) );
  XNOR U2778 ( .A(b[3749]), .B(n2429), .Z(c[3749]) );
  XNOR U2779 ( .A(a[3749]), .B(n2431), .Z(n2429) );
  IV U2780 ( .A(n2427), .Z(n2431) );
  XOR U2781 ( .A(n2432), .B(n2433), .Z(n2427) );
  ANDN U2782 ( .B(n2434), .A(n2435), .Z(n2432) );
  XNOR U2783 ( .A(b[3748]), .B(n2433), .Z(n2434) );
  XNOR U2784 ( .A(b[3748]), .B(n2435), .Z(c[3748]) );
  XNOR U2785 ( .A(a[3748]), .B(n2436), .Z(n2435) );
  IV U2786 ( .A(n2433), .Z(n2436) );
  XOR U2787 ( .A(n2437), .B(n2438), .Z(n2433) );
  ANDN U2788 ( .B(n2439), .A(n2440), .Z(n2437) );
  XNOR U2789 ( .A(b[3747]), .B(n2438), .Z(n2439) );
  XNOR U2790 ( .A(b[3747]), .B(n2440), .Z(c[3747]) );
  XNOR U2791 ( .A(a[3747]), .B(n2441), .Z(n2440) );
  IV U2792 ( .A(n2438), .Z(n2441) );
  XOR U2793 ( .A(n2442), .B(n2443), .Z(n2438) );
  ANDN U2794 ( .B(n2444), .A(n2445), .Z(n2442) );
  XNOR U2795 ( .A(b[3746]), .B(n2443), .Z(n2444) );
  XNOR U2796 ( .A(b[3746]), .B(n2445), .Z(c[3746]) );
  XNOR U2797 ( .A(a[3746]), .B(n2446), .Z(n2445) );
  IV U2798 ( .A(n2443), .Z(n2446) );
  XOR U2799 ( .A(n2447), .B(n2448), .Z(n2443) );
  ANDN U2800 ( .B(n2449), .A(n2450), .Z(n2447) );
  XNOR U2801 ( .A(b[3745]), .B(n2448), .Z(n2449) );
  XNOR U2802 ( .A(b[3745]), .B(n2450), .Z(c[3745]) );
  XNOR U2803 ( .A(a[3745]), .B(n2451), .Z(n2450) );
  IV U2804 ( .A(n2448), .Z(n2451) );
  XOR U2805 ( .A(n2452), .B(n2453), .Z(n2448) );
  ANDN U2806 ( .B(n2454), .A(n2455), .Z(n2452) );
  XNOR U2807 ( .A(b[3744]), .B(n2453), .Z(n2454) );
  XNOR U2808 ( .A(b[3744]), .B(n2455), .Z(c[3744]) );
  XNOR U2809 ( .A(a[3744]), .B(n2456), .Z(n2455) );
  IV U2810 ( .A(n2453), .Z(n2456) );
  XOR U2811 ( .A(n2457), .B(n2458), .Z(n2453) );
  ANDN U2812 ( .B(n2459), .A(n2460), .Z(n2457) );
  XNOR U2813 ( .A(b[3743]), .B(n2458), .Z(n2459) );
  XNOR U2814 ( .A(b[3743]), .B(n2460), .Z(c[3743]) );
  XNOR U2815 ( .A(a[3743]), .B(n2461), .Z(n2460) );
  IV U2816 ( .A(n2458), .Z(n2461) );
  XOR U2817 ( .A(n2462), .B(n2463), .Z(n2458) );
  ANDN U2818 ( .B(n2464), .A(n2465), .Z(n2462) );
  XNOR U2819 ( .A(b[3742]), .B(n2463), .Z(n2464) );
  XNOR U2820 ( .A(b[3742]), .B(n2465), .Z(c[3742]) );
  XNOR U2821 ( .A(a[3742]), .B(n2466), .Z(n2465) );
  IV U2822 ( .A(n2463), .Z(n2466) );
  XOR U2823 ( .A(n2467), .B(n2468), .Z(n2463) );
  ANDN U2824 ( .B(n2469), .A(n2470), .Z(n2467) );
  XNOR U2825 ( .A(b[3741]), .B(n2468), .Z(n2469) );
  XNOR U2826 ( .A(b[3741]), .B(n2470), .Z(c[3741]) );
  XNOR U2827 ( .A(a[3741]), .B(n2471), .Z(n2470) );
  IV U2828 ( .A(n2468), .Z(n2471) );
  XOR U2829 ( .A(n2472), .B(n2473), .Z(n2468) );
  ANDN U2830 ( .B(n2474), .A(n2475), .Z(n2472) );
  XNOR U2831 ( .A(b[3740]), .B(n2473), .Z(n2474) );
  XNOR U2832 ( .A(b[3740]), .B(n2475), .Z(c[3740]) );
  XNOR U2833 ( .A(a[3740]), .B(n2476), .Z(n2475) );
  IV U2834 ( .A(n2473), .Z(n2476) );
  XOR U2835 ( .A(n2477), .B(n2478), .Z(n2473) );
  ANDN U2836 ( .B(n2479), .A(n2480), .Z(n2477) );
  XNOR U2837 ( .A(b[3739]), .B(n2478), .Z(n2479) );
  XNOR U2838 ( .A(b[373]), .B(n2481), .Z(c[373]) );
  XNOR U2839 ( .A(b[3739]), .B(n2480), .Z(c[3739]) );
  XNOR U2840 ( .A(a[3739]), .B(n2482), .Z(n2480) );
  IV U2841 ( .A(n2478), .Z(n2482) );
  XOR U2842 ( .A(n2483), .B(n2484), .Z(n2478) );
  ANDN U2843 ( .B(n2485), .A(n2486), .Z(n2483) );
  XNOR U2844 ( .A(b[3738]), .B(n2484), .Z(n2485) );
  XNOR U2845 ( .A(b[3738]), .B(n2486), .Z(c[3738]) );
  XNOR U2846 ( .A(a[3738]), .B(n2487), .Z(n2486) );
  IV U2847 ( .A(n2484), .Z(n2487) );
  XOR U2848 ( .A(n2488), .B(n2489), .Z(n2484) );
  ANDN U2849 ( .B(n2490), .A(n2491), .Z(n2488) );
  XNOR U2850 ( .A(b[3737]), .B(n2489), .Z(n2490) );
  XNOR U2851 ( .A(b[3737]), .B(n2491), .Z(c[3737]) );
  XNOR U2852 ( .A(a[3737]), .B(n2492), .Z(n2491) );
  IV U2853 ( .A(n2489), .Z(n2492) );
  XOR U2854 ( .A(n2493), .B(n2494), .Z(n2489) );
  ANDN U2855 ( .B(n2495), .A(n2496), .Z(n2493) );
  XNOR U2856 ( .A(b[3736]), .B(n2494), .Z(n2495) );
  XNOR U2857 ( .A(b[3736]), .B(n2496), .Z(c[3736]) );
  XNOR U2858 ( .A(a[3736]), .B(n2497), .Z(n2496) );
  IV U2859 ( .A(n2494), .Z(n2497) );
  XOR U2860 ( .A(n2498), .B(n2499), .Z(n2494) );
  ANDN U2861 ( .B(n2500), .A(n2501), .Z(n2498) );
  XNOR U2862 ( .A(b[3735]), .B(n2499), .Z(n2500) );
  XNOR U2863 ( .A(b[3735]), .B(n2501), .Z(c[3735]) );
  XNOR U2864 ( .A(a[3735]), .B(n2502), .Z(n2501) );
  IV U2865 ( .A(n2499), .Z(n2502) );
  XOR U2866 ( .A(n2503), .B(n2504), .Z(n2499) );
  ANDN U2867 ( .B(n2505), .A(n2506), .Z(n2503) );
  XNOR U2868 ( .A(b[3734]), .B(n2504), .Z(n2505) );
  XNOR U2869 ( .A(b[3734]), .B(n2506), .Z(c[3734]) );
  XNOR U2870 ( .A(a[3734]), .B(n2507), .Z(n2506) );
  IV U2871 ( .A(n2504), .Z(n2507) );
  XOR U2872 ( .A(n2508), .B(n2509), .Z(n2504) );
  ANDN U2873 ( .B(n2510), .A(n2511), .Z(n2508) );
  XNOR U2874 ( .A(b[3733]), .B(n2509), .Z(n2510) );
  XNOR U2875 ( .A(b[3733]), .B(n2511), .Z(c[3733]) );
  XNOR U2876 ( .A(a[3733]), .B(n2512), .Z(n2511) );
  IV U2877 ( .A(n2509), .Z(n2512) );
  XOR U2878 ( .A(n2513), .B(n2514), .Z(n2509) );
  ANDN U2879 ( .B(n2515), .A(n2516), .Z(n2513) );
  XNOR U2880 ( .A(b[3732]), .B(n2514), .Z(n2515) );
  XNOR U2881 ( .A(b[3732]), .B(n2516), .Z(c[3732]) );
  XNOR U2882 ( .A(a[3732]), .B(n2517), .Z(n2516) );
  IV U2883 ( .A(n2514), .Z(n2517) );
  XOR U2884 ( .A(n2518), .B(n2519), .Z(n2514) );
  ANDN U2885 ( .B(n2520), .A(n2521), .Z(n2518) );
  XNOR U2886 ( .A(b[3731]), .B(n2519), .Z(n2520) );
  XNOR U2887 ( .A(b[3731]), .B(n2521), .Z(c[3731]) );
  XNOR U2888 ( .A(a[3731]), .B(n2522), .Z(n2521) );
  IV U2889 ( .A(n2519), .Z(n2522) );
  XOR U2890 ( .A(n2523), .B(n2524), .Z(n2519) );
  ANDN U2891 ( .B(n2525), .A(n2526), .Z(n2523) );
  XNOR U2892 ( .A(b[3730]), .B(n2524), .Z(n2525) );
  XNOR U2893 ( .A(b[3730]), .B(n2526), .Z(c[3730]) );
  XNOR U2894 ( .A(a[3730]), .B(n2527), .Z(n2526) );
  IV U2895 ( .A(n2524), .Z(n2527) );
  XOR U2896 ( .A(n2528), .B(n2529), .Z(n2524) );
  ANDN U2897 ( .B(n2530), .A(n2531), .Z(n2528) );
  XNOR U2898 ( .A(b[3729]), .B(n2529), .Z(n2530) );
  XNOR U2899 ( .A(b[372]), .B(n2532), .Z(c[372]) );
  XNOR U2900 ( .A(b[3729]), .B(n2531), .Z(c[3729]) );
  XNOR U2901 ( .A(a[3729]), .B(n2533), .Z(n2531) );
  IV U2902 ( .A(n2529), .Z(n2533) );
  XOR U2903 ( .A(n2534), .B(n2535), .Z(n2529) );
  ANDN U2904 ( .B(n2536), .A(n2537), .Z(n2534) );
  XNOR U2905 ( .A(b[3728]), .B(n2535), .Z(n2536) );
  XNOR U2906 ( .A(b[3728]), .B(n2537), .Z(c[3728]) );
  XNOR U2907 ( .A(a[3728]), .B(n2538), .Z(n2537) );
  IV U2908 ( .A(n2535), .Z(n2538) );
  XOR U2909 ( .A(n2539), .B(n2540), .Z(n2535) );
  ANDN U2910 ( .B(n2541), .A(n2542), .Z(n2539) );
  XNOR U2911 ( .A(b[3727]), .B(n2540), .Z(n2541) );
  XNOR U2912 ( .A(b[3727]), .B(n2542), .Z(c[3727]) );
  XNOR U2913 ( .A(a[3727]), .B(n2543), .Z(n2542) );
  IV U2914 ( .A(n2540), .Z(n2543) );
  XOR U2915 ( .A(n2544), .B(n2545), .Z(n2540) );
  ANDN U2916 ( .B(n2546), .A(n2547), .Z(n2544) );
  XNOR U2917 ( .A(b[3726]), .B(n2545), .Z(n2546) );
  XNOR U2918 ( .A(b[3726]), .B(n2547), .Z(c[3726]) );
  XNOR U2919 ( .A(a[3726]), .B(n2548), .Z(n2547) );
  IV U2920 ( .A(n2545), .Z(n2548) );
  XOR U2921 ( .A(n2549), .B(n2550), .Z(n2545) );
  ANDN U2922 ( .B(n2551), .A(n2552), .Z(n2549) );
  XNOR U2923 ( .A(b[3725]), .B(n2550), .Z(n2551) );
  XNOR U2924 ( .A(b[3725]), .B(n2552), .Z(c[3725]) );
  XNOR U2925 ( .A(a[3725]), .B(n2553), .Z(n2552) );
  IV U2926 ( .A(n2550), .Z(n2553) );
  XOR U2927 ( .A(n2554), .B(n2555), .Z(n2550) );
  ANDN U2928 ( .B(n2556), .A(n2557), .Z(n2554) );
  XNOR U2929 ( .A(b[3724]), .B(n2555), .Z(n2556) );
  XNOR U2930 ( .A(b[3724]), .B(n2557), .Z(c[3724]) );
  XNOR U2931 ( .A(a[3724]), .B(n2558), .Z(n2557) );
  IV U2932 ( .A(n2555), .Z(n2558) );
  XOR U2933 ( .A(n2559), .B(n2560), .Z(n2555) );
  ANDN U2934 ( .B(n2561), .A(n2562), .Z(n2559) );
  XNOR U2935 ( .A(b[3723]), .B(n2560), .Z(n2561) );
  XNOR U2936 ( .A(b[3723]), .B(n2562), .Z(c[3723]) );
  XNOR U2937 ( .A(a[3723]), .B(n2563), .Z(n2562) );
  IV U2938 ( .A(n2560), .Z(n2563) );
  XOR U2939 ( .A(n2564), .B(n2565), .Z(n2560) );
  ANDN U2940 ( .B(n2566), .A(n2567), .Z(n2564) );
  XNOR U2941 ( .A(b[3722]), .B(n2565), .Z(n2566) );
  XNOR U2942 ( .A(b[3722]), .B(n2567), .Z(c[3722]) );
  XNOR U2943 ( .A(a[3722]), .B(n2568), .Z(n2567) );
  IV U2944 ( .A(n2565), .Z(n2568) );
  XOR U2945 ( .A(n2569), .B(n2570), .Z(n2565) );
  ANDN U2946 ( .B(n2571), .A(n2572), .Z(n2569) );
  XNOR U2947 ( .A(b[3721]), .B(n2570), .Z(n2571) );
  XNOR U2948 ( .A(b[3721]), .B(n2572), .Z(c[3721]) );
  XNOR U2949 ( .A(a[3721]), .B(n2573), .Z(n2572) );
  IV U2950 ( .A(n2570), .Z(n2573) );
  XOR U2951 ( .A(n2574), .B(n2575), .Z(n2570) );
  ANDN U2952 ( .B(n2576), .A(n2577), .Z(n2574) );
  XNOR U2953 ( .A(b[3720]), .B(n2575), .Z(n2576) );
  XNOR U2954 ( .A(b[3720]), .B(n2577), .Z(c[3720]) );
  XNOR U2955 ( .A(a[3720]), .B(n2578), .Z(n2577) );
  IV U2956 ( .A(n2575), .Z(n2578) );
  XOR U2957 ( .A(n2579), .B(n2580), .Z(n2575) );
  ANDN U2958 ( .B(n2581), .A(n2582), .Z(n2579) );
  XNOR U2959 ( .A(b[3719]), .B(n2580), .Z(n2581) );
  XNOR U2960 ( .A(b[371]), .B(n2583), .Z(c[371]) );
  XNOR U2961 ( .A(b[3719]), .B(n2582), .Z(c[3719]) );
  XNOR U2962 ( .A(a[3719]), .B(n2584), .Z(n2582) );
  IV U2963 ( .A(n2580), .Z(n2584) );
  XOR U2964 ( .A(n2585), .B(n2586), .Z(n2580) );
  ANDN U2965 ( .B(n2587), .A(n2588), .Z(n2585) );
  XNOR U2966 ( .A(b[3718]), .B(n2586), .Z(n2587) );
  XNOR U2967 ( .A(b[3718]), .B(n2588), .Z(c[3718]) );
  XNOR U2968 ( .A(a[3718]), .B(n2589), .Z(n2588) );
  IV U2969 ( .A(n2586), .Z(n2589) );
  XOR U2970 ( .A(n2590), .B(n2591), .Z(n2586) );
  ANDN U2971 ( .B(n2592), .A(n2593), .Z(n2590) );
  XNOR U2972 ( .A(b[3717]), .B(n2591), .Z(n2592) );
  XNOR U2973 ( .A(b[3717]), .B(n2593), .Z(c[3717]) );
  XNOR U2974 ( .A(a[3717]), .B(n2594), .Z(n2593) );
  IV U2975 ( .A(n2591), .Z(n2594) );
  XOR U2976 ( .A(n2595), .B(n2596), .Z(n2591) );
  ANDN U2977 ( .B(n2597), .A(n2598), .Z(n2595) );
  XNOR U2978 ( .A(b[3716]), .B(n2596), .Z(n2597) );
  XNOR U2979 ( .A(b[3716]), .B(n2598), .Z(c[3716]) );
  XNOR U2980 ( .A(a[3716]), .B(n2599), .Z(n2598) );
  IV U2981 ( .A(n2596), .Z(n2599) );
  XOR U2982 ( .A(n2600), .B(n2601), .Z(n2596) );
  ANDN U2983 ( .B(n2602), .A(n2603), .Z(n2600) );
  XNOR U2984 ( .A(b[3715]), .B(n2601), .Z(n2602) );
  XNOR U2985 ( .A(b[3715]), .B(n2603), .Z(c[3715]) );
  XNOR U2986 ( .A(a[3715]), .B(n2604), .Z(n2603) );
  IV U2987 ( .A(n2601), .Z(n2604) );
  XOR U2988 ( .A(n2605), .B(n2606), .Z(n2601) );
  ANDN U2989 ( .B(n2607), .A(n2608), .Z(n2605) );
  XNOR U2990 ( .A(b[3714]), .B(n2606), .Z(n2607) );
  XNOR U2991 ( .A(b[3714]), .B(n2608), .Z(c[3714]) );
  XNOR U2992 ( .A(a[3714]), .B(n2609), .Z(n2608) );
  IV U2993 ( .A(n2606), .Z(n2609) );
  XOR U2994 ( .A(n2610), .B(n2611), .Z(n2606) );
  ANDN U2995 ( .B(n2612), .A(n2613), .Z(n2610) );
  XNOR U2996 ( .A(b[3713]), .B(n2611), .Z(n2612) );
  XNOR U2997 ( .A(b[3713]), .B(n2613), .Z(c[3713]) );
  XNOR U2998 ( .A(a[3713]), .B(n2614), .Z(n2613) );
  IV U2999 ( .A(n2611), .Z(n2614) );
  XOR U3000 ( .A(n2615), .B(n2616), .Z(n2611) );
  ANDN U3001 ( .B(n2617), .A(n2618), .Z(n2615) );
  XNOR U3002 ( .A(b[3712]), .B(n2616), .Z(n2617) );
  XNOR U3003 ( .A(b[3712]), .B(n2618), .Z(c[3712]) );
  XNOR U3004 ( .A(a[3712]), .B(n2619), .Z(n2618) );
  IV U3005 ( .A(n2616), .Z(n2619) );
  XOR U3006 ( .A(n2620), .B(n2621), .Z(n2616) );
  ANDN U3007 ( .B(n2622), .A(n2623), .Z(n2620) );
  XNOR U3008 ( .A(b[3711]), .B(n2621), .Z(n2622) );
  XNOR U3009 ( .A(b[3711]), .B(n2623), .Z(c[3711]) );
  XNOR U3010 ( .A(a[3711]), .B(n2624), .Z(n2623) );
  IV U3011 ( .A(n2621), .Z(n2624) );
  XOR U3012 ( .A(n2625), .B(n2626), .Z(n2621) );
  ANDN U3013 ( .B(n2627), .A(n2628), .Z(n2625) );
  XNOR U3014 ( .A(b[3710]), .B(n2626), .Z(n2627) );
  XNOR U3015 ( .A(b[3710]), .B(n2628), .Z(c[3710]) );
  XNOR U3016 ( .A(a[3710]), .B(n2629), .Z(n2628) );
  IV U3017 ( .A(n2626), .Z(n2629) );
  XOR U3018 ( .A(n2630), .B(n2631), .Z(n2626) );
  ANDN U3019 ( .B(n2632), .A(n2633), .Z(n2630) );
  XNOR U3020 ( .A(b[3709]), .B(n2631), .Z(n2632) );
  XNOR U3021 ( .A(b[370]), .B(n2634), .Z(c[370]) );
  XNOR U3022 ( .A(b[3709]), .B(n2633), .Z(c[3709]) );
  XNOR U3023 ( .A(a[3709]), .B(n2635), .Z(n2633) );
  IV U3024 ( .A(n2631), .Z(n2635) );
  XOR U3025 ( .A(n2636), .B(n2637), .Z(n2631) );
  ANDN U3026 ( .B(n2638), .A(n2639), .Z(n2636) );
  XNOR U3027 ( .A(b[3708]), .B(n2637), .Z(n2638) );
  XNOR U3028 ( .A(b[3708]), .B(n2639), .Z(c[3708]) );
  XNOR U3029 ( .A(a[3708]), .B(n2640), .Z(n2639) );
  IV U3030 ( .A(n2637), .Z(n2640) );
  XOR U3031 ( .A(n2641), .B(n2642), .Z(n2637) );
  ANDN U3032 ( .B(n2643), .A(n2644), .Z(n2641) );
  XNOR U3033 ( .A(b[3707]), .B(n2642), .Z(n2643) );
  XNOR U3034 ( .A(b[3707]), .B(n2644), .Z(c[3707]) );
  XNOR U3035 ( .A(a[3707]), .B(n2645), .Z(n2644) );
  IV U3036 ( .A(n2642), .Z(n2645) );
  XOR U3037 ( .A(n2646), .B(n2647), .Z(n2642) );
  ANDN U3038 ( .B(n2648), .A(n2649), .Z(n2646) );
  XNOR U3039 ( .A(b[3706]), .B(n2647), .Z(n2648) );
  XNOR U3040 ( .A(b[3706]), .B(n2649), .Z(c[3706]) );
  XNOR U3041 ( .A(a[3706]), .B(n2650), .Z(n2649) );
  IV U3042 ( .A(n2647), .Z(n2650) );
  XOR U3043 ( .A(n2651), .B(n2652), .Z(n2647) );
  ANDN U3044 ( .B(n2653), .A(n2654), .Z(n2651) );
  XNOR U3045 ( .A(b[3705]), .B(n2652), .Z(n2653) );
  XNOR U3046 ( .A(b[3705]), .B(n2654), .Z(c[3705]) );
  XNOR U3047 ( .A(a[3705]), .B(n2655), .Z(n2654) );
  IV U3048 ( .A(n2652), .Z(n2655) );
  XOR U3049 ( .A(n2656), .B(n2657), .Z(n2652) );
  ANDN U3050 ( .B(n2658), .A(n2659), .Z(n2656) );
  XNOR U3051 ( .A(b[3704]), .B(n2657), .Z(n2658) );
  XNOR U3052 ( .A(b[3704]), .B(n2659), .Z(c[3704]) );
  XNOR U3053 ( .A(a[3704]), .B(n2660), .Z(n2659) );
  IV U3054 ( .A(n2657), .Z(n2660) );
  XOR U3055 ( .A(n2661), .B(n2662), .Z(n2657) );
  ANDN U3056 ( .B(n2663), .A(n2664), .Z(n2661) );
  XNOR U3057 ( .A(b[3703]), .B(n2662), .Z(n2663) );
  XNOR U3058 ( .A(b[3703]), .B(n2664), .Z(c[3703]) );
  XNOR U3059 ( .A(a[3703]), .B(n2665), .Z(n2664) );
  IV U3060 ( .A(n2662), .Z(n2665) );
  XOR U3061 ( .A(n2666), .B(n2667), .Z(n2662) );
  ANDN U3062 ( .B(n2668), .A(n2669), .Z(n2666) );
  XNOR U3063 ( .A(b[3702]), .B(n2667), .Z(n2668) );
  XNOR U3064 ( .A(b[3702]), .B(n2669), .Z(c[3702]) );
  XNOR U3065 ( .A(a[3702]), .B(n2670), .Z(n2669) );
  IV U3066 ( .A(n2667), .Z(n2670) );
  XOR U3067 ( .A(n2671), .B(n2672), .Z(n2667) );
  ANDN U3068 ( .B(n2673), .A(n2674), .Z(n2671) );
  XNOR U3069 ( .A(b[3701]), .B(n2672), .Z(n2673) );
  XNOR U3070 ( .A(b[3701]), .B(n2674), .Z(c[3701]) );
  XNOR U3071 ( .A(a[3701]), .B(n2675), .Z(n2674) );
  IV U3072 ( .A(n2672), .Z(n2675) );
  XOR U3073 ( .A(n2676), .B(n2677), .Z(n2672) );
  ANDN U3074 ( .B(n2678), .A(n2679), .Z(n2676) );
  XNOR U3075 ( .A(b[3700]), .B(n2677), .Z(n2678) );
  XNOR U3076 ( .A(b[3700]), .B(n2679), .Z(c[3700]) );
  XNOR U3077 ( .A(a[3700]), .B(n2680), .Z(n2679) );
  IV U3078 ( .A(n2677), .Z(n2680) );
  XOR U3079 ( .A(n2681), .B(n2682), .Z(n2677) );
  ANDN U3080 ( .B(n2683), .A(n2684), .Z(n2681) );
  XNOR U3081 ( .A(b[3699]), .B(n2682), .Z(n2683) );
  XNOR U3082 ( .A(b[36]), .B(n2685), .Z(c[36]) );
  XNOR U3083 ( .A(b[369]), .B(n2686), .Z(c[369]) );
  XNOR U3084 ( .A(b[3699]), .B(n2684), .Z(c[3699]) );
  XNOR U3085 ( .A(a[3699]), .B(n2687), .Z(n2684) );
  IV U3086 ( .A(n2682), .Z(n2687) );
  XOR U3087 ( .A(n2688), .B(n2689), .Z(n2682) );
  ANDN U3088 ( .B(n2690), .A(n2691), .Z(n2688) );
  XNOR U3089 ( .A(b[3698]), .B(n2689), .Z(n2690) );
  XNOR U3090 ( .A(b[3698]), .B(n2691), .Z(c[3698]) );
  XNOR U3091 ( .A(a[3698]), .B(n2692), .Z(n2691) );
  IV U3092 ( .A(n2689), .Z(n2692) );
  XOR U3093 ( .A(n2693), .B(n2694), .Z(n2689) );
  ANDN U3094 ( .B(n2695), .A(n2696), .Z(n2693) );
  XNOR U3095 ( .A(b[3697]), .B(n2694), .Z(n2695) );
  XNOR U3096 ( .A(b[3697]), .B(n2696), .Z(c[3697]) );
  XNOR U3097 ( .A(a[3697]), .B(n2697), .Z(n2696) );
  IV U3098 ( .A(n2694), .Z(n2697) );
  XOR U3099 ( .A(n2698), .B(n2699), .Z(n2694) );
  ANDN U3100 ( .B(n2700), .A(n2701), .Z(n2698) );
  XNOR U3101 ( .A(b[3696]), .B(n2699), .Z(n2700) );
  XNOR U3102 ( .A(b[3696]), .B(n2701), .Z(c[3696]) );
  XNOR U3103 ( .A(a[3696]), .B(n2702), .Z(n2701) );
  IV U3104 ( .A(n2699), .Z(n2702) );
  XOR U3105 ( .A(n2703), .B(n2704), .Z(n2699) );
  ANDN U3106 ( .B(n2705), .A(n2706), .Z(n2703) );
  XNOR U3107 ( .A(b[3695]), .B(n2704), .Z(n2705) );
  XNOR U3108 ( .A(b[3695]), .B(n2706), .Z(c[3695]) );
  XNOR U3109 ( .A(a[3695]), .B(n2707), .Z(n2706) );
  IV U3110 ( .A(n2704), .Z(n2707) );
  XOR U3111 ( .A(n2708), .B(n2709), .Z(n2704) );
  ANDN U3112 ( .B(n2710), .A(n2711), .Z(n2708) );
  XNOR U3113 ( .A(b[3694]), .B(n2709), .Z(n2710) );
  XNOR U3114 ( .A(b[3694]), .B(n2711), .Z(c[3694]) );
  XNOR U3115 ( .A(a[3694]), .B(n2712), .Z(n2711) );
  IV U3116 ( .A(n2709), .Z(n2712) );
  XOR U3117 ( .A(n2713), .B(n2714), .Z(n2709) );
  ANDN U3118 ( .B(n2715), .A(n2716), .Z(n2713) );
  XNOR U3119 ( .A(b[3693]), .B(n2714), .Z(n2715) );
  XNOR U3120 ( .A(b[3693]), .B(n2716), .Z(c[3693]) );
  XNOR U3121 ( .A(a[3693]), .B(n2717), .Z(n2716) );
  IV U3122 ( .A(n2714), .Z(n2717) );
  XOR U3123 ( .A(n2718), .B(n2719), .Z(n2714) );
  ANDN U3124 ( .B(n2720), .A(n2721), .Z(n2718) );
  XNOR U3125 ( .A(b[3692]), .B(n2719), .Z(n2720) );
  XNOR U3126 ( .A(b[3692]), .B(n2721), .Z(c[3692]) );
  XNOR U3127 ( .A(a[3692]), .B(n2722), .Z(n2721) );
  IV U3128 ( .A(n2719), .Z(n2722) );
  XOR U3129 ( .A(n2723), .B(n2724), .Z(n2719) );
  ANDN U3130 ( .B(n2725), .A(n2726), .Z(n2723) );
  XNOR U3131 ( .A(b[3691]), .B(n2724), .Z(n2725) );
  XNOR U3132 ( .A(b[3691]), .B(n2726), .Z(c[3691]) );
  XNOR U3133 ( .A(a[3691]), .B(n2727), .Z(n2726) );
  IV U3134 ( .A(n2724), .Z(n2727) );
  XOR U3135 ( .A(n2728), .B(n2729), .Z(n2724) );
  ANDN U3136 ( .B(n2730), .A(n2731), .Z(n2728) );
  XNOR U3137 ( .A(b[3690]), .B(n2729), .Z(n2730) );
  XNOR U3138 ( .A(b[3690]), .B(n2731), .Z(c[3690]) );
  XNOR U3139 ( .A(a[3690]), .B(n2732), .Z(n2731) );
  IV U3140 ( .A(n2729), .Z(n2732) );
  XOR U3141 ( .A(n2733), .B(n2734), .Z(n2729) );
  ANDN U3142 ( .B(n2735), .A(n2736), .Z(n2733) );
  XNOR U3143 ( .A(b[3689]), .B(n2734), .Z(n2735) );
  XNOR U3144 ( .A(b[368]), .B(n2737), .Z(c[368]) );
  XNOR U3145 ( .A(b[3689]), .B(n2736), .Z(c[3689]) );
  XNOR U3146 ( .A(a[3689]), .B(n2738), .Z(n2736) );
  IV U3147 ( .A(n2734), .Z(n2738) );
  XOR U3148 ( .A(n2739), .B(n2740), .Z(n2734) );
  ANDN U3149 ( .B(n2741), .A(n2742), .Z(n2739) );
  XNOR U3150 ( .A(b[3688]), .B(n2740), .Z(n2741) );
  XNOR U3151 ( .A(b[3688]), .B(n2742), .Z(c[3688]) );
  XNOR U3152 ( .A(a[3688]), .B(n2743), .Z(n2742) );
  IV U3153 ( .A(n2740), .Z(n2743) );
  XOR U3154 ( .A(n2744), .B(n2745), .Z(n2740) );
  ANDN U3155 ( .B(n2746), .A(n2747), .Z(n2744) );
  XNOR U3156 ( .A(b[3687]), .B(n2745), .Z(n2746) );
  XNOR U3157 ( .A(b[3687]), .B(n2747), .Z(c[3687]) );
  XNOR U3158 ( .A(a[3687]), .B(n2748), .Z(n2747) );
  IV U3159 ( .A(n2745), .Z(n2748) );
  XOR U3160 ( .A(n2749), .B(n2750), .Z(n2745) );
  ANDN U3161 ( .B(n2751), .A(n2752), .Z(n2749) );
  XNOR U3162 ( .A(b[3686]), .B(n2750), .Z(n2751) );
  XNOR U3163 ( .A(b[3686]), .B(n2752), .Z(c[3686]) );
  XNOR U3164 ( .A(a[3686]), .B(n2753), .Z(n2752) );
  IV U3165 ( .A(n2750), .Z(n2753) );
  XOR U3166 ( .A(n2754), .B(n2755), .Z(n2750) );
  ANDN U3167 ( .B(n2756), .A(n2757), .Z(n2754) );
  XNOR U3168 ( .A(b[3685]), .B(n2755), .Z(n2756) );
  XNOR U3169 ( .A(b[3685]), .B(n2757), .Z(c[3685]) );
  XNOR U3170 ( .A(a[3685]), .B(n2758), .Z(n2757) );
  IV U3171 ( .A(n2755), .Z(n2758) );
  XOR U3172 ( .A(n2759), .B(n2760), .Z(n2755) );
  ANDN U3173 ( .B(n2761), .A(n2762), .Z(n2759) );
  XNOR U3174 ( .A(b[3684]), .B(n2760), .Z(n2761) );
  XNOR U3175 ( .A(b[3684]), .B(n2762), .Z(c[3684]) );
  XNOR U3176 ( .A(a[3684]), .B(n2763), .Z(n2762) );
  IV U3177 ( .A(n2760), .Z(n2763) );
  XOR U3178 ( .A(n2764), .B(n2765), .Z(n2760) );
  ANDN U3179 ( .B(n2766), .A(n2767), .Z(n2764) );
  XNOR U3180 ( .A(b[3683]), .B(n2765), .Z(n2766) );
  XNOR U3181 ( .A(b[3683]), .B(n2767), .Z(c[3683]) );
  XNOR U3182 ( .A(a[3683]), .B(n2768), .Z(n2767) );
  IV U3183 ( .A(n2765), .Z(n2768) );
  XOR U3184 ( .A(n2769), .B(n2770), .Z(n2765) );
  ANDN U3185 ( .B(n2771), .A(n2772), .Z(n2769) );
  XNOR U3186 ( .A(b[3682]), .B(n2770), .Z(n2771) );
  XNOR U3187 ( .A(b[3682]), .B(n2772), .Z(c[3682]) );
  XNOR U3188 ( .A(a[3682]), .B(n2773), .Z(n2772) );
  IV U3189 ( .A(n2770), .Z(n2773) );
  XOR U3190 ( .A(n2774), .B(n2775), .Z(n2770) );
  ANDN U3191 ( .B(n2776), .A(n2777), .Z(n2774) );
  XNOR U3192 ( .A(b[3681]), .B(n2775), .Z(n2776) );
  XNOR U3193 ( .A(b[3681]), .B(n2777), .Z(c[3681]) );
  XNOR U3194 ( .A(a[3681]), .B(n2778), .Z(n2777) );
  IV U3195 ( .A(n2775), .Z(n2778) );
  XOR U3196 ( .A(n2779), .B(n2780), .Z(n2775) );
  ANDN U3197 ( .B(n2781), .A(n2782), .Z(n2779) );
  XNOR U3198 ( .A(b[3680]), .B(n2780), .Z(n2781) );
  XNOR U3199 ( .A(b[3680]), .B(n2782), .Z(c[3680]) );
  XNOR U3200 ( .A(a[3680]), .B(n2783), .Z(n2782) );
  IV U3201 ( .A(n2780), .Z(n2783) );
  XOR U3202 ( .A(n2784), .B(n2785), .Z(n2780) );
  ANDN U3203 ( .B(n2786), .A(n2787), .Z(n2784) );
  XNOR U3204 ( .A(b[3679]), .B(n2785), .Z(n2786) );
  XNOR U3205 ( .A(b[367]), .B(n2788), .Z(c[367]) );
  XNOR U3206 ( .A(b[3679]), .B(n2787), .Z(c[3679]) );
  XNOR U3207 ( .A(a[3679]), .B(n2789), .Z(n2787) );
  IV U3208 ( .A(n2785), .Z(n2789) );
  XOR U3209 ( .A(n2790), .B(n2791), .Z(n2785) );
  ANDN U3210 ( .B(n2792), .A(n2793), .Z(n2790) );
  XNOR U3211 ( .A(b[3678]), .B(n2791), .Z(n2792) );
  XNOR U3212 ( .A(b[3678]), .B(n2793), .Z(c[3678]) );
  XNOR U3213 ( .A(a[3678]), .B(n2794), .Z(n2793) );
  IV U3214 ( .A(n2791), .Z(n2794) );
  XOR U3215 ( .A(n2795), .B(n2796), .Z(n2791) );
  ANDN U3216 ( .B(n2797), .A(n2798), .Z(n2795) );
  XNOR U3217 ( .A(b[3677]), .B(n2796), .Z(n2797) );
  XNOR U3218 ( .A(b[3677]), .B(n2798), .Z(c[3677]) );
  XNOR U3219 ( .A(a[3677]), .B(n2799), .Z(n2798) );
  IV U3220 ( .A(n2796), .Z(n2799) );
  XOR U3221 ( .A(n2800), .B(n2801), .Z(n2796) );
  ANDN U3222 ( .B(n2802), .A(n2803), .Z(n2800) );
  XNOR U3223 ( .A(b[3676]), .B(n2801), .Z(n2802) );
  XNOR U3224 ( .A(b[3676]), .B(n2803), .Z(c[3676]) );
  XNOR U3225 ( .A(a[3676]), .B(n2804), .Z(n2803) );
  IV U3226 ( .A(n2801), .Z(n2804) );
  XOR U3227 ( .A(n2805), .B(n2806), .Z(n2801) );
  ANDN U3228 ( .B(n2807), .A(n2808), .Z(n2805) );
  XNOR U3229 ( .A(b[3675]), .B(n2806), .Z(n2807) );
  XNOR U3230 ( .A(b[3675]), .B(n2808), .Z(c[3675]) );
  XNOR U3231 ( .A(a[3675]), .B(n2809), .Z(n2808) );
  IV U3232 ( .A(n2806), .Z(n2809) );
  XOR U3233 ( .A(n2810), .B(n2811), .Z(n2806) );
  ANDN U3234 ( .B(n2812), .A(n2813), .Z(n2810) );
  XNOR U3235 ( .A(b[3674]), .B(n2811), .Z(n2812) );
  XNOR U3236 ( .A(b[3674]), .B(n2813), .Z(c[3674]) );
  XNOR U3237 ( .A(a[3674]), .B(n2814), .Z(n2813) );
  IV U3238 ( .A(n2811), .Z(n2814) );
  XOR U3239 ( .A(n2815), .B(n2816), .Z(n2811) );
  ANDN U3240 ( .B(n2817), .A(n2818), .Z(n2815) );
  XNOR U3241 ( .A(b[3673]), .B(n2816), .Z(n2817) );
  XNOR U3242 ( .A(b[3673]), .B(n2818), .Z(c[3673]) );
  XNOR U3243 ( .A(a[3673]), .B(n2819), .Z(n2818) );
  IV U3244 ( .A(n2816), .Z(n2819) );
  XOR U3245 ( .A(n2820), .B(n2821), .Z(n2816) );
  ANDN U3246 ( .B(n2822), .A(n2823), .Z(n2820) );
  XNOR U3247 ( .A(b[3672]), .B(n2821), .Z(n2822) );
  XNOR U3248 ( .A(b[3672]), .B(n2823), .Z(c[3672]) );
  XNOR U3249 ( .A(a[3672]), .B(n2824), .Z(n2823) );
  IV U3250 ( .A(n2821), .Z(n2824) );
  XOR U3251 ( .A(n2825), .B(n2826), .Z(n2821) );
  ANDN U3252 ( .B(n2827), .A(n2828), .Z(n2825) );
  XNOR U3253 ( .A(b[3671]), .B(n2826), .Z(n2827) );
  XNOR U3254 ( .A(b[3671]), .B(n2828), .Z(c[3671]) );
  XNOR U3255 ( .A(a[3671]), .B(n2829), .Z(n2828) );
  IV U3256 ( .A(n2826), .Z(n2829) );
  XOR U3257 ( .A(n2830), .B(n2831), .Z(n2826) );
  ANDN U3258 ( .B(n2832), .A(n2833), .Z(n2830) );
  XNOR U3259 ( .A(b[3670]), .B(n2831), .Z(n2832) );
  XNOR U3260 ( .A(b[3670]), .B(n2833), .Z(c[3670]) );
  XNOR U3261 ( .A(a[3670]), .B(n2834), .Z(n2833) );
  IV U3262 ( .A(n2831), .Z(n2834) );
  XOR U3263 ( .A(n2835), .B(n2836), .Z(n2831) );
  ANDN U3264 ( .B(n2837), .A(n2838), .Z(n2835) );
  XNOR U3265 ( .A(b[3669]), .B(n2836), .Z(n2837) );
  XNOR U3266 ( .A(b[366]), .B(n2839), .Z(c[366]) );
  XNOR U3267 ( .A(b[3669]), .B(n2838), .Z(c[3669]) );
  XNOR U3268 ( .A(a[3669]), .B(n2840), .Z(n2838) );
  IV U3269 ( .A(n2836), .Z(n2840) );
  XOR U3270 ( .A(n2841), .B(n2842), .Z(n2836) );
  ANDN U3271 ( .B(n2843), .A(n2844), .Z(n2841) );
  XNOR U3272 ( .A(b[3668]), .B(n2842), .Z(n2843) );
  XNOR U3273 ( .A(b[3668]), .B(n2844), .Z(c[3668]) );
  XNOR U3274 ( .A(a[3668]), .B(n2845), .Z(n2844) );
  IV U3275 ( .A(n2842), .Z(n2845) );
  XOR U3276 ( .A(n2846), .B(n2847), .Z(n2842) );
  ANDN U3277 ( .B(n2848), .A(n2849), .Z(n2846) );
  XNOR U3278 ( .A(b[3667]), .B(n2847), .Z(n2848) );
  XNOR U3279 ( .A(b[3667]), .B(n2849), .Z(c[3667]) );
  XNOR U3280 ( .A(a[3667]), .B(n2850), .Z(n2849) );
  IV U3281 ( .A(n2847), .Z(n2850) );
  XOR U3282 ( .A(n2851), .B(n2852), .Z(n2847) );
  ANDN U3283 ( .B(n2853), .A(n2854), .Z(n2851) );
  XNOR U3284 ( .A(b[3666]), .B(n2852), .Z(n2853) );
  XNOR U3285 ( .A(b[3666]), .B(n2854), .Z(c[3666]) );
  XNOR U3286 ( .A(a[3666]), .B(n2855), .Z(n2854) );
  IV U3287 ( .A(n2852), .Z(n2855) );
  XOR U3288 ( .A(n2856), .B(n2857), .Z(n2852) );
  ANDN U3289 ( .B(n2858), .A(n2859), .Z(n2856) );
  XNOR U3290 ( .A(b[3665]), .B(n2857), .Z(n2858) );
  XNOR U3291 ( .A(b[3665]), .B(n2859), .Z(c[3665]) );
  XNOR U3292 ( .A(a[3665]), .B(n2860), .Z(n2859) );
  IV U3293 ( .A(n2857), .Z(n2860) );
  XOR U3294 ( .A(n2861), .B(n2862), .Z(n2857) );
  ANDN U3295 ( .B(n2863), .A(n2864), .Z(n2861) );
  XNOR U3296 ( .A(b[3664]), .B(n2862), .Z(n2863) );
  XNOR U3297 ( .A(b[3664]), .B(n2864), .Z(c[3664]) );
  XNOR U3298 ( .A(a[3664]), .B(n2865), .Z(n2864) );
  IV U3299 ( .A(n2862), .Z(n2865) );
  XOR U3300 ( .A(n2866), .B(n2867), .Z(n2862) );
  ANDN U3301 ( .B(n2868), .A(n2869), .Z(n2866) );
  XNOR U3302 ( .A(b[3663]), .B(n2867), .Z(n2868) );
  XNOR U3303 ( .A(b[3663]), .B(n2869), .Z(c[3663]) );
  XNOR U3304 ( .A(a[3663]), .B(n2870), .Z(n2869) );
  IV U3305 ( .A(n2867), .Z(n2870) );
  XOR U3306 ( .A(n2871), .B(n2872), .Z(n2867) );
  ANDN U3307 ( .B(n2873), .A(n2874), .Z(n2871) );
  XNOR U3308 ( .A(b[3662]), .B(n2872), .Z(n2873) );
  XNOR U3309 ( .A(b[3662]), .B(n2874), .Z(c[3662]) );
  XNOR U3310 ( .A(a[3662]), .B(n2875), .Z(n2874) );
  IV U3311 ( .A(n2872), .Z(n2875) );
  XOR U3312 ( .A(n2876), .B(n2877), .Z(n2872) );
  ANDN U3313 ( .B(n2878), .A(n2879), .Z(n2876) );
  XNOR U3314 ( .A(b[3661]), .B(n2877), .Z(n2878) );
  XNOR U3315 ( .A(b[3661]), .B(n2879), .Z(c[3661]) );
  XNOR U3316 ( .A(a[3661]), .B(n2880), .Z(n2879) );
  IV U3317 ( .A(n2877), .Z(n2880) );
  XOR U3318 ( .A(n2881), .B(n2882), .Z(n2877) );
  ANDN U3319 ( .B(n2883), .A(n2884), .Z(n2881) );
  XNOR U3320 ( .A(b[3660]), .B(n2882), .Z(n2883) );
  XNOR U3321 ( .A(b[3660]), .B(n2884), .Z(c[3660]) );
  XNOR U3322 ( .A(a[3660]), .B(n2885), .Z(n2884) );
  IV U3323 ( .A(n2882), .Z(n2885) );
  XOR U3324 ( .A(n2886), .B(n2887), .Z(n2882) );
  ANDN U3325 ( .B(n2888), .A(n2889), .Z(n2886) );
  XNOR U3326 ( .A(b[3659]), .B(n2887), .Z(n2888) );
  XNOR U3327 ( .A(b[365]), .B(n2890), .Z(c[365]) );
  XNOR U3328 ( .A(b[3659]), .B(n2889), .Z(c[3659]) );
  XNOR U3329 ( .A(a[3659]), .B(n2891), .Z(n2889) );
  IV U3330 ( .A(n2887), .Z(n2891) );
  XOR U3331 ( .A(n2892), .B(n2893), .Z(n2887) );
  ANDN U3332 ( .B(n2894), .A(n2895), .Z(n2892) );
  XNOR U3333 ( .A(b[3658]), .B(n2893), .Z(n2894) );
  XNOR U3334 ( .A(b[3658]), .B(n2895), .Z(c[3658]) );
  XNOR U3335 ( .A(a[3658]), .B(n2896), .Z(n2895) );
  IV U3336 ( .A(n2893), .Z(n2896) );
  XOR U3337 ( .A(n2897), .B(n2898), .Z(n2893) );
  ANDN U3338 ( .B(n2899), .A(n2900), .Z(n2897) );
  XNOR U3339 ( .A(b[3657]), .B(n2898), .Z(n2899) );
  XNOR U3340 ( .A(b[3657]), .B(n2900), .Z(c[3657]) );
  XNOR U3341 ( .A(a[3657]), .B(n2901), .Z(n2900) );
  IV U3342 ( .A(n2898), .Z(n2901) );
  XOR U3343 ( .A(n2902), .B(n2903), .Z(n2898) );
  ANDN U3344 ( .B(n2904), .A(n2905), .Z(n2902) );
  XNOR U3345 ( .A(b[3656]), .B(n2903), .Z(n2904) );
  XNOR U3346 ( .A(b[3656]), .B(n2905), .Z(c[3656]) );
  XNOR U3347 ( .A(a[3656]), .B(n2906), .Z(n2905) );
  IV U3348 ( .A(n2903), .Z(n2906) );
  XOR U3349 ( .A(n2907), .B(n2908), .Z(n2903) );
  ANDN U3350 ( .B(n2909), .A(n2910), .Z(n2907) );
  XNOR U3351 ( .A(b[3655]), .B(n2908), .Z(n2909) );
  XNOR U3352 ( .A(b[3655]), .B(n2910), .Z(c[3655]) );
  XNOR U3353 ( .A(a[3655]), .B(n2911), .Z(n2910) );
  IV U3354 ( .A(n2908), .Z(n2911) );
  XOR U3355 ( .A(n2912), .B(n2913), .Z(n2908) );
  ANDN U3356 ( .B(n2914), .A(n2915), .Z(n2912) );
  XNOR U3357 ( .A(b[3654]), .B(n2913), .Z(n2914) );
  XNOR U3358 ( .A(b[3654]), .B(n2915), .Z(c[3654]) );
  XNOR U3359 ( .A(a[3654]), .B(n2916), .Z(n2915) );
  IV U3360 ( .A(n2913), .Z(n2916) );
  XOR U3361 ( .A(n2917), .B(n2918), .Z(n2913) );
  ANDN U3362 ( .B(n2919), .A(n2920), .Z(n2917) );
  XNOR U3363 ( .A(b[3653]), .B(n2918), .Z(n2919) );
  XNOR U3364 ( .A(b[3653]), .B(n2920), .Z(c[3653]) );
  XNOR U3365 ( .A(a[3653]), .B(n2921), .Z(n2920) );
  IV U3366 ( .A(n2918), .Z(n2921) );
  XOR U3367 ( .A(n2922), .B(n2923), .Z(n2918) );
  ANDN U3368 ( .B(n2924), .A(n2925), .Z(n2922) );
  XNOR U3369 ( .A(b[3652]), .B(n2923), .Z(n2924) );
  XNOR U3370 ( .A(b[3652]), .B(n2925), .Z(c[3652]) );
  XNOR U3371 ( .A(a[3652]), .B(n2926), .Z(n2925) );
  IV U3372 ( .A(n2923), .Z(n2926) );
  XOR U3373 ( .A(n2927), .B(n2928), .Z(n2923) );
  ANDN U3374 ( .B(n2929), .A(n2930), .Z(n2927) );
  XNOR U3375 ( .A(b[3651]), .B(n2928), .Z(n2929) );
  XNOR U3376 ( .A(b[3651]), .B(n2930), .Z(c[3651]) );
  XNOR U3377 ( .A(a[3651]), .B(n2931), .Z(n2930) );
  IV U3378 ( .A(n2928), .Z(n2931) );
  XOR U3379 ( .A(n2932), .B(n2933), .Z(n2928) );
  ANDN U3380 ( .B(n2934), .A(n2935), .Z(n2932) );
  XNOR U3381 ( .A(b[3650]), .B(n2933), .Z(n2934) );
  XNOR U3382 ( .A(b[3650]), .B(n2935), .Z(c[3650]) );
  XNOR U3383 ( .A(a[3650]), .B(n2936), .Z(n2935) );
  IV U3384 ( .A(n2933), .Z(n2936) );
  XOR U3385 ( .A(n2937), .B(n2938), .Z(n2933) );
  ANDN U3386 ( .B(n2939), .A(n2940), .Z(n2937) );
  XNOR U3387 ( .A(b[3649]), .B(n2938), .Z(n2939) );
  XNOR U3388 ( .A(b[364]), .B(n2941), .Z(c[364]) );
  XNOR U3389 ( .A(b[3649]), .B(n2940), .Z(c[3649]) );
  XNOR U3390 ( .A(a[3649]), .B(n2942), .Z(n2940) );
  IV U3391 ( .A(n2938), .Z(n2942) );
  XOR U3392 ( .A(n2943), .B(n2944), .Z(n2938) );
  ANDN U3393 ( .B(n2945), .A(n2946), .Z(n2943) );
  XNOR U3394 ( .A(b[3648]), .B(n2944), .Z(n2945) );
  XNOR U3395 ( .A(b[3648]), .B(n2946), .Z(c[3648]) );
  XNOR U3396 ( .A(a[3648]), .B(n2947), .Z(n2946) );
  IV U3397 ( .A(n2944), .Z(n2947) );
  XOR U3398 ( .A(n2948), .B(n2949), .Z(n2944) );
  ANDN U3399 ( .B(n2950), .A(n2951), .Z(n2948) );
  XNOR U3400 ( .A(b[3647]), .B(n2949), .Z(n2950) );
  XNOR U3401 ( .A(b[3647]), .B(n2951), .Z(c[3647]) );
  XNOR U3402 ( .A(a[3647]), .B(n2952), .Z(n2951) );
  IV U3403 ( .A(n2949), .Z(n2952) );
  XOR U3404 ( .A(n2953), .B(n2954), .Z(n2949) );
  ANDN U3405 ( .B(n2955), .A(n2956), .Z(n2953) );
  XNOR U3406 ( .A(b[3646]), .B(n2954), .Z(n2955) );
  XNOR U3407 ( .A(b[3646]), .B(n2956), .Z(c[3646]) );
  XNOR U3408 ( .A(a[3646]), .B(n2957), .Z(n2956) );
  IV U3409 ( .A(n2954), .Z(n2957) );
  XOR U3410 ( .A(n2958), .B(n2959), .Z(n2954) );
  ANDN U3411 ( .B(n2960), .A(n2961), .Z(n2958) );
  XNOR U3412 ( .A(b[3645]), .B(n2959), .Z(n2960) );
  XNOR U3413 ( .A(b[3645]), .B(n2961), .Z(c[3645]) );
  XNOR U3414 ( .A(a[3645]), .B(n2962), .Z(n2961) );
  IV U3415 ( .A(n2959), .Z(n2962) );
  XOR U3416 ( .A(n2963), .B(n2964), .Z(n2959) );
  ANDN U3417 ( .B(n2965), .A(n2966), .Z(n2963) );
  XNOR U3418 ( .A(b[3644]), .B(n2964), .Z(n2965) );
  XNOR U3419 ( .A(b[3644]), .B(n2966), .Z(c[3644]) );
  XNOR U3420 ( .A(a[3644]), .B(n2967), .Z(n2966) );
  IV U3421 ( .A(n2964), .Z(n2967) );
  XOR U3422 ( .A(n2968), .B(n2969), .Z(n2964) );
  ANDN U3423 ( .B(n2970), .A(n2971), .Z(n2968) );
  XNOR U3424 ( .A(b[3643]), .B(n2969), .Z(n2970) );
  XNOR U3425 ( .A(b[3643]), .B(n2971), .Z(c[3643]) );
  XNOR U3426 ( .A(a[3643]), .B(n2972), .Z(n2971) );
  IV U3427 ( .A(n2969), .Z(n2972) );
  XOR U3428 ( .A(n2973), .B(n2974), .Z(n2969) );
  ANDN U3429 ( .B(n2975), .A(n2976), .Z(n2973) );
  XNOR U3430 ( .A(b[3642]), .B(n2974), .Z(n2975) );
  XNOR U3431 ( .A(b[3642]), .B(n2976), .Z(c[3642]) );
  XNOR U3432 ( .A(a[3642]), .B(n2977), .Z(n2976) );
  IV U3433 ( .A(n2974), .Z(n2977) );
  XOR U3434 ( .A(n2978), .B(n2979), .Z(n2974) );
  ANDN U3435 ( .B(n2980), .A(n2981), .Z(n2978) );
  XNOR U3436 ( .A(b[3641]), .B(n2979), .Z(n2980) );
  XNOR U3437 ( .A(b[3641]), .B(n2981), .Z(c[3641]) );
  XNOR U3438 ( .A(a[3641]), .B(n2982), .Z(n2981) );
  IV U3439 ( .A(n2979), .Z(n2982) );
  XOR U3440 ( .A(n2983), .B(n2984), .Z(n2979) );
  ANDN U3441 ( .B(n2985), .A(n2986), .Z(n2983) );
  XNOR U3442 ( .A(b[3640]), .B(n2984), .Z(n2985) );
  XNOR U3443 ( .A(b[3640]), .B(n2986), .Z(c[3640]) );
  XNOR U3444 ( .A(a[3640]), .B(n2987), .Z(n2986) );
  IV U3445 ( .A(n2984), .Z(n2987) );
  XOR U3446 ( .A(n2988), .B(n2989), .Z(n2984) );
  ANDN U3447 ( .B(n2990), .A(n2991), .Z(n2988) );
  XNOR U3448 ( .A(b[3639]), .B(n2989), .Z(n2990) );
  XNOR U3449 ( .A(b[363]), .B(n2992), .Z(c[363]) );
  XNOR U3450 ( .A(b[3639]), .B(n2991), .Z(c[3639]) );
  XNOR U3451 ( .A(a[3639]), .B(n2993), .Z(n2991) );
  IV U3452 ( .A(n2989), .Z(n2993) );
  XOR U3453 ( .A(n2994), .B(n2995), .Z(n2989) );
  ANDN U3454 ( .B(n2996), .A(n2997), .Z(n2994) );
  XNOR U3455 ( .A(b[3638]), .B(n2995), .Z(n2996) );
  XNOR U3456 ( .A(b[3638]), .B(n2997), .Z(c[3638]) );
  XNOR U3457 ( .A(a[3638]), .B(n2998), .Z(n2997) );
  IV U3458 ( .A(n2995), .Z(n2998) );
  XOR U3459 ( .A(n2999), .B(n3000), .Z(n2995) );
  ANDN U3460 ( .B(n3001), .A(n3002), .Z(n2999) );
  XNOR U3461 ( .A(b[3637]), .B(n3000), .Z(n3001) );
  XNOR U3462 ( .A(b[3637]), .B(n3002), .Z(c[3637]) );
  XNOR U3463 ( .A(a[3637]), .B(n3003), .Z(n3002) );
  IV U3464 ( .A(n3000), .Z(n3003) );
  XOR U3465 ( .A(n3004), .B(n3005), .Z(n3000) );
  ANDN U3466 ( .B(n3006), .A(n3007), .Z(n3004) );
  XNOR U3467 ( .A(b[3636]), .B(n3005), .Z(n3006) );
  XNOR U3468 ( .A(b[3636]), .B(n3007), .Z(c[3636]) );
  XNOR U3469 ( .A(a[3636]), .B(n3008), .Z(n3007) );
  IV U3470 ( .A(n3005), .Z(n3008) );
  XOR U3471 ( .A(n3009), .B(n3010), .Z(n3005) );
  ANDN U3472 ( .B(n3011), .A(n3012), .Z(n3009) );
  XNOR U3473 ( .A(b[3635]), .B(n3010), .Z(n3011) );
  XNOR U3474 ( .A(b[3635]), .B(n3012), .Z(c[3635]) );
  XNOR U3475 ( .A(a[3635]), .B(n3013), .Z(n3012) );
  IV U3476 ( .A(n3010), .Z(n3013) );
  XOR U3477 ( .A(n3014), .B(n3015), .Z(n3010) );
  ANDN U3478 ( .B(n3016), .A(n3017), .Z(n3014) );
  XNOR U3479 ( .A(b[3634]), .B(n3015), .Z(n3016) );
  XNOR U3480 ( .A(b[3634]), .B(n3017), .Z(c[3634]) );
  XNOR U3481 ( .A(a[3634]), .B(n3018), .Z(n3017) );
  IV U3482 ( .A(n3015), .Z(n3018) );
  XOR U3483 ( .A(n3019), .B(n3020), .Z(n3015) );
  ANDN U3484 ( .B(n3021), .A(n3022), .Z(n3019) );
  XNOR U3485 ( .A(b[3633]), .B(n3020), .Z(n3021) );
  XNOR U3486 ( .A(b[3633]), .B(n3022), .Z(c[3633]) );
  XNOR U3487 ( .A(a[3633]), .B(n3023), .Z(n3022) );
  IV U3488 ( .A(n3020), .Z(n3023) );
  XOR U3489 ( .A(n3024), .B(n3025), .Z(n3020) );
  ANDN U3490 ( .B(n3026), .A(n3027), .Z(n3024) );
  XNOR U3491 ( .A(b[3632]), .B(n3025), .Z(n3026) );
  XNOR U3492 ( .A(b[3632]), .B(n3027), .Z(c[3632]) );
  XNOR U3493 ( .A(a[3632]), .B(n3028), .Z(n3027) );
  IV U3494 ( .A(n3025), .Z(n3028) );
  XOR U3495 ( .A(n3029), .B(n3030), .Z(n3025) );
  ANDN U3496 ( .B(n3031), .A(n3032), .Z(n3029) );
  XNOR U3497 ( .A(b[3631]), .B(n3030), .Z(n3031) );
  XNOR U3498 ( .A(b[3631]), .B(n3032), .Z(c[3631]) );
  XNOR U3499 ( .A(a[3631]), .B(n3033), .Z(n3032) );
  IV U3500 ( .A(n3030), .Z(n3033) );
  XOR U3501 ( .A(n3034), .B(n3035), .Z(n3030) );
  ANDN U3502 ( .B(n3036), .A(n3037), .Z(n3034) );
  XNOR U3503 ( .A(b[3630]), .B(n3035), .Z(n3036) );
  XNOR U3504 ( .A(b[3630]), .B(n3037), .Z(c[3630]) );
  XNOR U3505 ( .A(a[3630]), .B(n3038), .Z(n3037) );
  IV U3506 ( .A(n3035), .Z(n3038) );
  XOR U3507 ( .A(n3039), .B(n3040), .Z(n3035) );
  ANDN U3508 ( .B(n3041), .A(n3042), .Z(n3039) );
  XNOR U3509 ( .A(b[3629]), .B(n3040), .Z(n3041) );
  XNOR U3510 ( .A(b[362]), .B(n3043), .Z(c[362]) );
  XNOR U3511 ( .A(b[3629]), .B(n3042), .Z(c[3629]) );
  XNOR U3512 ( .A(a[3629]), .B(n3044), .Z(n3042) );
  IV U3513 ( .A(n3040), .Z(n3044) );
  XOR U3514 ( .A(n3045), .B(n3046), .Z(n3040) );
  ANDN U3515 ( .B(n3047), .A(n3048), .Z(n3045) );
  XNOR U3516 ( .A(b[3628]), .B(n3046), .Z(n3047) );
  XNOR U3517 ( .A(b[3628]), .B(n3048), .Z(c[3628]) );
  XNOR U3518 ( .A(a[3628]), .B(n3049), .Z(n3048) );
  IV U3519 ( .A(n3046), .Z(n3049) );
  XOR U3520 ( .A(n3050), .B(n3051), .Z(n3046) );
  ANDN U3521 ( .B(n3052), .A(n3053), .Z(n3050) );
  XNOR U3522 ( .A(b[3627]), .B(n3051), .Z(n3052) );
  XNOR U3523 ( .A(b[3627]), .B(n3053), .Z(c[3627]) );
  XNOR U3524 ( .A(a[3627]), .B(n3054), .Z(n3053) );
  IV U3525 ( .A(n3051), .Z(n3054) );
  XOR U3526 ( .A(n3055), .B(n3056), .Z(n3051) );
  ANDN U3527 ( .B(n3057), .A(n3058), .Z(n3055) );
  XNOR U3528 ( .A(b[3626]), .B(n3056), .Z(n3057) );
  XNOR U3529 ( .A(b[3626]), .B(n3058), .Z(c[3626]) );
  XNOR U3530 ( .A(a[3626]), .B(n3059), .Z(n3058) );
  IV U3531 ( .A(n3056), .Z(n3059) );
  XOR U3532 ( .A(n3060), .B(n3061), .Z(n3056) );
  ANDN U3533 ( .B(n3062), .A(n3063), .Z(n3060) );
  XNOR U3534 ( .A(b[3625]), .B(n3061), .Z(n3062) );
  XNOR U3535 ( .A(b[3625]), .B(n3063), .Z(c[3625]) );
  XNOR U3536 ( .A(a[3625]), .B(n3064), .Z(n3063) );
  IV U3537 ( .A(n3061), .Z(n3064) );
  XOR U3538 ( .A(n3065), .B(n3066), .Z(n3061) );
  ANDN U3539 ( .B(n3067), .A(n3068), .Z(n3065) );
  XNOR U3540 ( .A(b[3624]), .B(n3066), .Z(n3067) );
  XNOR U3541 ( .A(b[3624]), .B(n3068), .Z(c[3624]) );
  XNOR U3542 ( .A(a[3624]), .B(n3069), .Z(n3068) );
  IV U3543 ( .A(n3066), .Z(n3069) );
  XOR U3544 ( .A(n3070), .B(n3071), .Z(n3066) );
  ANDN U3545 ( .B(n3072), .A(n3073), .Z(n3070) );
  XNOR U3546 ( .A(b[3623]), .B(n3071), .Z(n3072) );
  XNOR U3547 ( .A(b[3623]), .B(n3073), .Z(c[3623]) );
  XNOR U3548 ( .A(a[3623]), .B(n3074), .Z(n3073) );
  IV U3549 ( .A(n3071), .Z(n3074) );
  XOR U3550 ( .A(n3075), .B(n3076), .Z(n3071) );
  ANDN U3551 ( .B(n3077), .A(n3078), .Z(n3075) );
  XNOR U3552 ( .A(b[3622]), .B(n3076), .Z(n3077) );
  XNOR U3553 ( .A(b[3622]), .B(n3078), .Z(c[3622]) );
  XNOR U3554 ( .A(a[3622]), .B(n3079), .Z(n3078) );
  IV U3555 ( .A(n3076), .Z(n3079) );
  XOR U3556 ( .A(n3080), .B(n3081), .Z(n3076) );
  ANDN U3557 ( .B(n3082), .A(n3083), .Z(n3080) );
  XNOR U3558 ( .A(b[3621]), .B(n3081), .Z(n3082) );
  XNOR U3559 ( .A(b[3621]), .B(n3083), .Z(c[3621]) );
  XNOR U3560 ( .A(a[3621]), .B(n3084), .Z(n3083) );
  IV U3561 ( .A(n3081), .Z(n3084) );
  XOR U3562 ( .A(n3085), .B(n3086), .Z(n3081) );
  ANDN U3563 ( .B(n3087), .A(n3088), .Z(n3085) );
  XNOR U3564 ( .A(b[3620]), .B(n3086), .Z(n3087) );
  XNOR U3565 ( .A(b[3620]), .B(n3088), .Z(c[3620]) );
  XNOR U3566 ( .A(a[3620]), .B(n3089), .Z(n3088) );
  IV U3567 ( .A(n3086), .Z(n3089) );
  XOR U3568 ( .A(n3090), .B(n3091), .Z(n3086) );
  ANDN U3569 ( .B(n3092), .A(n3093), .Z(n3090) );
  XNOR U3570 ( .A(b[3619]), .B(n3091), .Z(n3092) );
  XNOR U3571 ( .A(b[361]), .B(n3094), .Z(c[361]) );
  XNOR U3572 ( .A(b[3619]), .B(n3093), .Z(c[3619]) );
  XNOR U3573 ( .A(a[3619]), .B(n3095), .Z(n3093) );
  IV U3574 ( .A(n3091), .Z(n3095) );
  XOR U3575 ( .A(n3096), .B(n3097), .Z(n3091) );
  ANDN U3576 ( .B(n3098), .A(n3099), .Z(n3096) );
  XNOR U3577 ( .A(b[3618]), .B(n3097), .Z(n3098) );
  XNOR U3578 ( .A(b[3618]), .B(n3099), .Z(c[3618]) );
  XNOR U3579 ( .A(a[3618]), .B(n3100), .Z(n3099) );
  IV U3580 ( .A(n3097), .Z(n3100) );
  XOR U3581 ( .A(n3101), .B(n3102), .Z(n3097) );
  ANDN U3582 ( .B(n3103), .A(n3104), .Z(n3101) );
  XNOR U3583 ( .A(b[3617]), .B(n3102), .Z(n3103) );
  XNOR U3584 ( .A(b[3617]), .B(n3104), .Z(c[3617]) );
  XNOR U3585 ( .A(a[3617]), .B(n3105), .Z(n3104) );
  IV U3586 ( .A(n3102), .Z(n3105) );
  XOR U3587 ( .A(n3106), .B(n3107), .Z(n3102) );
  ANDN U3588 ( .B(n3108), .A(n3109), .Z(n3106) );
  XNOR U3589 ( .A(b[3616]), .B(n3107), .Z(n3108) );
  XNOR U3590 ( .A(b[3616]), .B(n3109), .Z(c[3616]) );
  XNOR U3591 ( .A(a[3616]), .B(n3110), .Z(n3109) );
  IV U3592 ( .A(n3107), .Z(n3110) );
  XOR U3593 ( .A(n3111), .B(n3112), .Z(n3107) );
  ANDN U3594 ( .B(n3113), .A(n3114), .Z(n3111) );
  XNOR U3595 ( .A(b[3615]), .B(n3112), .Z(n3113) );
  XNOR U3596 ( .A(b[3615]), .B(n3114), .Z(c[3615]) );
  XNOR U3597 ( .A(a[3615]), .B(n3115), .Z(n3114) );
  IV U3598 ( .A(n3112), .Z(n3115) );
  XOR U3599 ( .A(n3116), .B(n3117), .Z(n3112) );
  ANDN U3600 ( .B(n3118), .A(n3119), .Z(n3116) );
  XNOR U3601 ( .A(b[3614]), .B(n3117), .Z(n3118) );
  XNOR U3602 ( .A(b[3614]), .B(n3119), .Z(c[3614]) );
  XNOR U3603 ( .A(a[3614]), .B(n3120), .Z(n3119) );
  IV U3604 ( .A(n3117), .Z(n3120) );
  XOR U3605 ( .A(n3121), .B(n3122), .Z(n3117) );
  ANDN U3606 ( .B(n3123), .A(n3124), .Z(n3121) );
  XNOR U3607 ( .A(b[3613]), .B(n3122), .Z(n3123) );
  XNOR U3608 ( .A(b[3613]), .B(n3124), .Z(c[3613]) );
  XNOR U3609 ( .A(a[3613]), .B(n3125), .Z(n3124) );
  IV U3610 ( .A(n3122), .Z(n3125) );
  XOR U3611 ( .A(n3126), .B(n3127), .Z(n3122) );
  ANDN U3612 ( .B(n3128), .A(n3129), .Z(n3126) );
  XNOR U3613 ( .A(b[3612]), .B(n3127), .Z(n3128) );
  XNOR U3614 ( .A(b[3612]), .B(n3129), .Z(c[3612]) );
  XNOR U3615 ( .A(a[3612]), .B(n3130), .Z(n3129) );
  IV U3616 ( .A(n3127), .Z(n3130) );
  XOR U3617 ( .A(n3131), .B(n3132), .Z(n3127) );
  ANDN U3618 ( .B(n3133), .A(n3134), .Z(n3131) );
  XNOR U3619 ( .A(b[3611]), .B(n3132), .Z(n3133) );
  XNOR U3620 ( .A(b[3611]), .B(n3134), .Z(c[3611]) );
  XNOR U3621 ( .A(a[3611]), .B(n3135), .Z(n3134) );
  IV U3622 ( .A(n3132), .Z(n3135) );
  XOR U3623 ( .A(n3136), .B(n3137), .Z(n3132) );
  ANDN U3624 ( .B(n3138), .A(n3139), .Z(n3136) );
  XNOR U3625 ( .A(b[3610]), .B(n3137), .Z(n3138) );
  XNOR U3626 ( .A(b[3610]), .B(n3139), .Z(c[3610]) );
  XNOR U3627 ( .A(a[3610]), .B(n3140), .Z(n3139) );
  IV U3628 ( .A(n3137), .Z(n3140) );
  XOR U3629 ( .A(n3141), .B(n3142), .Z(n3137) );
  ANDN U3630 ( .B(n3143), .A(n3144), .Z(n3141) );
  XNOR U3631 ( .A(b[3609]), .B(n3142), .Z(n3143) );
  XNOR U3632 ( .A(b[360]), .B(n3145), .Z(c[360]) );
  XNOR U3633 ( .A(b[3609]), .B(n3144), .Z(c[3609]) );
  XNOR U3634 ( .A(a[3609]), .B(n3146), .Z(n3144) );
  IV U3635 ( .A(n3142), .Z(n3146) );
  XOR U3636 ( .A(n3147), .B(n3148), .Z(n3142) );
  ANDN U3637 ( .B(n3149), .A(n3150), .Z(n3147) );
  XNOR U3638 ( .A(b[3608]), .B(n3148), .Z(n3149) );
  XNOR U3639 ( .A(b[3608]), .B(n3150), .Z(c[3608]) );
  XNOR U3640 ( .A(a[3608]), .B(n3151), .Z(n3150) );
  IV U3641 ( .A(n3148), .Z(n3151) );
  XOR U3642 ( .A(n3152), .B(n3153), .Z(n3148) );
  ANDN U3643 ( .B(n3154), .A(n3155), .Z(n3152) );
  XNOR U3644 ( .A(b[3607]), .B(n3153), .Z(n3154) );
  XNOR U3645 ( .A(b[3607]), .B(n3155), .Z(c[3607]) );
  XNOR U3646 ( .A(a[3607]), .B(n3156), .Z(n3155) );
  IV U3647 ( .A(n3153), .Z(n3156) );
  XOR U3648 ( .A(n3157), .B(n3158), .Z(n3153) );
  ANDN U3649 ( .B(n3159), .A(n3160), .Z(n3157) );
  XNOR U3650 ( .A(b[3606]), .B(n3158), .Z(n3159) );
  XNOR U3651 ( .A(b[3606]), .B(n3160), .Z(c[3606]) );
  XNOR U3652 ( .A(a[3606]), .B(n3161), .Z(n3160) );
  IV U3653 ( .A(n3158), .Z(n3161) );
  XOR U3654 ( .A(n3162), .B(n3163), .Z(n3158) );
  ANDN U3655 ( .B(n3164), .A(n3165), .Z(n3162) );
  XNOR U3656 ( .A(b[3605]), .B(n3163), .Z(n3164) );
  XNOR U3657 ( .A(b[3605]), .B(n3165), .Z(c[3605]) );
  XNOR U3658 ( .A(a[3605]), .B(n3166), .Z(n3165) );
  IV U3659 ( .A(n3163), .Z(n3166) );
  XOR U3660 ( .A(n3167), .B(n3168), .Z(n3163) );
  ANDN U3661 ( .B(n3169), .A(n3170), .Z(n3167) );
  XNOR U3662 ( .A(b[3604]), .B(n3168), .Z(n3169) );
  XNOR U3663 ( .A(b[3604]), .B(n3170), .Z(c[3604]) );
  XNOR U3664 ( .A(a[3604]), .B(n3171), .Z(n3170) );
  IV U3665 ( .A(n3168), .Z(n3171) );
  XOR U3666 ( .A(n3172), .B(n3173), .Z(n3168) );
  ANDN U3667 ( .B(n3174), .A(n3175), .Z(n3172) );
  XNOR U3668 ( .A(b[3603]), .B(n3173), .Z(n3174) );
  XNOR U3669 ( .A(b[3603]), .B(n3175), .Z(c[3603]) );
  XNOR U3670 ( .A(a[3603]), .B(n3176), .Z(n3175) );
  IV U3671 ( .A(n3173), .Z(n3176) );
  XOR U3672 ( .A(n3177), .B(n3178), .Z(n3173) );
  ANDN U3673 ( .B(n3179), .A(n3180), .Z(n3177) );
  XNOR U3674 ( .A(b[3602]), .B(n3178), .Z(n3179) );
  XNOR U3675 ( .A(b[3602]), .B(n3180), .Z(c[3602]) );
  XNOR U3676 ( .A(a[3602]), .B(n3181), .Z(n3180) );
  IV U3677 ( .A(n3178), .Z(n3181) );
  XOR U3678 ( .A(n3182), .B(n3183), .Z(n3178) );
  ANDN U3679 ( .B(n3184), .A(n3185), .Z(n3182) );
  XNOR U3680 ( .A(b[3601]), .B(n3183), .Z(n3184) );
  XNOR U3681 ( .A(b[3601]), .B(n3185), .Z(c[3601]) );
  XNOR U3682 ( .A(a[3601]), .B(n3186), .Z(n3185) );
  IV U3683 ( .A(n3183), .Z(n3186) );
  XOR U3684 ( .A(n3187), .B(n3188), .Z(n3183) );
  ANDN U3685 ( .B(n3189), .A(n3190), .Z(n3187) );
  XNOR U3686 ( .A(b[3600]), .B(n3188), .Z(n3189) );
  XNOR U3687 ( .A(b[3600]), .B(n3190), .Z(c[3600]) );
  XNOR U3688 ( .A(a[3600]), .B(n3191), .Z(n3190) );
  IV U3689 ( .A(n3188), .Z(n3191) );
  XOR U3690 ( .A(n3192), .B(n3193), .Z(n3188) );
  ANDN U3691 ( .B(n3194), .A(n3195), .Z(n3192) );
  XNOR U3692 ( .A(b[3599]), .B(n3193), .Z(n3194) );
  XNOR U3693 ( .A(b[35]), .B(n3196), .Z(c[35]) );
  XNOR U3694 ( .A(b[359]), .B(n3197), .Z(c[359]) );
  XNOR U3695 ( .A(b[3599]), .B(n3195), .Z(c[3599]) );
  XNOR U3696 ( .A(a[3599]), .B(n3198), .Z(n3195) );
  IV U3697 ( .A(n3193), .Z(n3198) );
  XOR U3698 ( .A(n3199), .B(n3200), .Z(n3193) );
  ANDN U3699 ( .B(n3201), .A(n3202), .Z(n3199) );
  XNOR U3700 ( .A(b[3598]), .B(n3200), .Z(n3201) );
  XNOR U3701 ( .A(b[3598]), .B(n3202), .Z(c[3598]) );
  XNOR U3702 ( .A(a[3598]), .B(n3203), .Z(n3202) );
  IV U3703 ( .A(n3200), .Z(n3203) );
  XOR U3704 ( .A(n3204), .B(n3205), .Z(n3200) );
  ANDN U3705 ( .B(n3206), .A(n3207), .Z(n3204) );
  XNOR U3706 ( .A(b[3597]), .B(n3205), .Z(n3206) );
  XNOR U3707 ( .A(b[3597]), .B(n3207), .Z(c[3597]) );
  XNOR U3708 ( .A(a[3597]), .B(n3208), .Z(n3207) );
  IV U3709 ( .A(n3205), .Z(n3208) );
  XOR U3710 ( .A(n3209), .B(n3210), .Z(n3205) );
  ANDN U3711 ( .B(n3211), .A(n3212), .Z(n3209) );
  XNOR U3712 ( .A(b[3596]), .B(n3210), .Z(n3211) );
  XNOR U3713 ( .A(b[3596]), .B(n3212), .Z(c[3596]) );
  XNOR U3714 ( .A(a[3596]), .B(n3213), .Z(n3212) );
  IV U3715 ( .A(n3210), .Z(n3213) );
  XOR U3716 ( .A(n3214), .B(n3215), .Z(n3210) );
  ANDN U3717 ( .B(n3216), .A(n3217), .Z(n3214) );
  XNOR U3718 ( .A(b[3595]), .B(n3215), .Z(n3216) );
  XNOR U3719 ( .A(b[3595]), .B(n3217), .Z(c[3595]) );
  XNOR U3720 ( .A(a[3595]), .B(n3218), .Z(n3217) );
  IV U3721 ( .A(n3215), .Z(n3218) );
  XOR U3722 ( .A(n3219), .B(n3220), .Z(n3215) );
  ANDN U3723 ( .B(n3221), .A(n3222), .Z(n3219) );
  XNOR U3724 ( .A(b[3594]), .B(n3220), .Z(n3221) );
  XNOR U3725 ( .A(b[3594]), .B(n3222), .Z(c[3594]) );
  XNOR U3726 ( .A(a[3594]), .B(n3223), .Z(n3222) );
  IV U3727 ( .A(n3220), .Z(n3223) );
  XOR U3728 ( .A(n3224), .B(n3225), .Z(n3220) );
  ANDN U3729 ( .B(n3226), .A(n3227), .Z(n3224) );
  XNOR U3730 ( .A(b[3593]), .B(n3225), .Z(n3226) );
  XNOR U3731 ( .A(b[3593]), .B(n3227), .Z(c[3593]) );
  XNOR U3732 ( .A(a[3593]), .B(n3228), .Z(n3227) );
  IV U3733 ( .A(n3225), .Z(n3228) );
  XOR U3734 ( .A(n3229), .B(n3230), .Z(n3225) );
  ANDN U3735 ( .B(n3231), .A(n3232), .Z(n3229) );
  XNOR U3736 ( .A(b[3592]), .B(n3230), .Z(n3231) );
  XNOR U3737 ( .A(b[3592]), .B(n3232), .Z(c[3592]) );
  XNOR U3738 ( .A(a[3592]), .B(n3233), .Z(n3232) );
  IV U3739 ( .A(n3230), .Z(n3233) );
  XOR U3740 ( .A(n3234), .B(n3235), .Z(n3230) );
  ANDN U3741 ( .B(n3236), .A(n3237), .Z(n3234) );
  XNOR U3742 ( .A(b[3591]), .B(n3235), .Z(n3236) );
  XNOR U3743 ( .A(b[3591]), .B(n3237), .Z(c[3591]) );
  XNOR U3744 ( .A(a[3591]), .B(n3238), .Z(n3237) );
  IV U3745 ( .A(n3235), .Z(n3238) );
  XOR U3746 ( .A(n3239), .B(n3240), .Z(n3235) );
  ANDN U3747 ( .B(n3241), .A(n3242), .Z(n3239) );
  XNOR U3748 ( .A(b[3590]), .B(n3240), .Z(n3241) );
  XNOR U3749 ( .A(b[3590]), .B(n3242), .Z(c[3590]) );
  XNOR U3750 ( .A(a[3590]), .B(n3243), .Z(n3242) );
  IV U3751 ( .A(n3240), .Z(n3243) );
  XOR U3752 ( .A(n3244), .B(n3245), .Z(n3240) );
  ANDN U3753 ( .B(n3246), .A(n3247), .Z(n3244) );
  XNOR U3754 ( .A(b[3589]), .B(n3245), .Z(n3246) );
  XNOR U3755 ( .A(b[358]), .B(n3248), .Z(c[358]) );
  XNOR U3756 ( .A(b[3589]), .B(n3247), .Z(c[3589]) );
  XNOR U3757 ( .A(a[3589]), .B(n3249), .Z(n3247) );
  IV U3758 ( .A(n3245), .Z(n3249) );
  XOR U3759 ( .A(n3250), .B(n3251), .Z(n3245) );
  ANDN U3760 ( .B(n3252), .A(n3253), .Z(n3250) );
  XNOR U3761 ( .A(b[3588]), .B(n3251), .Z(n3252) );
  XNOR U3762 ( .A(b[3588]), .B(n3253), .Z(c[3588]) );
  XNOR U3763 ( .A(a[3588]), .B(n3254), .Z(n3253) );
  IV U3764 ( .A(n3251), .Z(n3254) );
  XOR U3765 ( .A(n3255), .B(n3256), .Z(n3251) );
  ANDN U3766 ( .B(n3257), .A(n3258), .Z(n3255) );
  XNOR U3767 ( .A(b[3587]), .B(n3256), .Z(n3257) );
  XNOR U3768 ( .A(b[3587]), .B(n3258), .Z(c[3587]) );
  XNOR U3769 ( .A(a[3587]), .B(n3259), .Z(n3258) );
  IV U3770 ( .A(n3256), .Z(n3259) );
  XOR U3771 ( .A(n3260), .B(n3261), .Z(n3256) );
  ANDN U3772 ( .B(n3262), .A(n3263), .Z(n3260) );
  XNOR U3773 ( .A(b[3586]), .B(n3261), .Z(n3262) );
  XNOR U3774 ( .A(b[3586]), .B(n3263), .Z(c[3586]) );
  XNOR U3775 ( .A(a[3586]), .B(n3264), .Z(n3263) );
  IV U3776 ( .A(n3261), .Z(n3264) );
  XOR U3777 ( .A(n3265), .B(n3266), .Z(n3261) );
  ANDN U3778 ( .B(n3267), .A(n3268), .Z(n3265) );
  XNOR U3779 ( .A(b[3585]), .B(n3266), .Z(n3267) );
  XNOR U3780 ( .A(b[3585]), .B(n3268), .Z(c[3585]) );
  XNOR U3781 ( .A(a[3585]), .B(n3269), .Z(n3268) );
  IV U3782 ( .A(n3266), .Z(n3269) );
  XOR U3783 ( .A(n3270), .B(n3271), .Z(n3266) );
  ANDN U3784 ( .B(n3272), .A(n3273), .Z(n3270) );
  XNOR U3785 ( .A(b[3584]), .B(n3271), .Z(n3272) );
  XNOR U3786 ( .A(b[3584]), .B(n3273), .Z(c[3584]) );
  XNOR U3787 ( .A(a[3584]), .B(n3274), .Z(n3273) );
  IV U3788 ( .A(n3271), .Z(n3274) );
  XOR U3789 ( .A(n3275), .B(n3276), .Z(n3271) );
  ANDN U3790 ( .B(n3277), .A(n3278), .Z(n3275) );
  XNOR U3791 ( .A(b[3583]), .B(n3276), .Z(n3277) );
  XNOR U3792 ( .A(b[3583]), .B(n3278), .Z(c[3583]) );
  XNOR U3793 ( .A(a[3583]), .B(n3279), .Z(n3278) );
  IV U3794 ( .A(n3276), .Z(n3279) );
  XOR U3795 ( .A(n3280), .B(n3281), .Z(n3276) );
  ANDN U3796 ( .B(n3282), .A(n3283), .Z(n3280) );
  XNOR U3797 ( .A(b[3582]), .B(n3281), .Z(n3282) );
  XNOR U3798 ( .A(b[3582]), .B(n3283), .Z(c[3582]) );
  XNOR U3799 ( .A(a[3582]), .B(n3284), .Z(n3283) );
  IV U3800 ( .A(n3281), .Z(n3284) );
  XOR U3801 ( .A(n3285), .B(n3286), .Z(n3281) );
  ANDN U3802 ( .B(n3287), .A(n3288), .Z(n3285) );
  XNOR U3803 ( .A(b[3581]), .B(n3286), .Z(n3287) );
  XNOR U3804 ( .A(b[3581]), .B(n3288), .Z(c[3581]) );
  XNOR U3805 ( .A(a[3581]), .B(n3289), .Z(n3288) );
  IV U3806 ( .A(n3286), .Z(n3289) );
  XOR U3807 ( .A(n3290), .B(n3291), .Z(n3286) );
  ANDN U3808 ( .B(n3292), .A(n3293), .Z(n3290) );
  XNOR U3809 ( .A(b[3580]), .B(n3291), .Z(n3292) );
  XNOR U3810 ( .A(b[3580]), .B(n3293), .Z(c[3580]) );
  XNOR U3811 ( .A(a[3580]), .B(n3294), .Z(n3293) );
  IV U3812 ( .A(n3291), .Z(n3294) );
  XOR U3813 ( .A(n3295), .B(n3296), .Z(n3291) );
  ANDN U3814 ( .B(n3297), .A(n3298), .Z(n3295) );
  XNOR U3815 ( .A(b[3579]), .B(n3296), .Z(n3297) );
  XNOR U3816 ( .A(b[357]), .B(n3299), .Z(c[357]) );
  XNOR U3817 ( .A(b[3579]), .B(n3298), .Z(c[3579]) );
  XNOR U3818 ( .A(a[3579]), .B(n3300), .Z(n3298) );
  IV U3819 ( .A(n3296), .Z(n3300) );
  XOR U3820 ( .A(n3301), .B(n3302), .Z(n3296) );
  ANDN U3821 ( .B(n3303), .A(n3304), .Z(n3301) );
  XNOR U3822 ( .A(b[3578]), .B(n3302), .Z(n3303) );
  XNOR U3823 ( .A(b[3578]), .B(n3304), .Z(c[3578]) );
  XNOR U3824 ( .A(a[3578]), .B(n3305), .Z(n3304) );
  IV U3825 ( .A(n3302), .Z(n3305) );
  XOR U3826 ( .A(n3306), .B(n3307), .Z(n3302) );
  ANDN U3827 ( .B(n3308), .A(n3309), .Z(n3306) );
  XNOR U3828 ( .A(b[3577]), .B(n3307), .Z(n3308) );
  XNOR U3829 ( .A(b[3577]), .B(n3309), .Z(c[3577]) );
  XNOR U3830 ( .A(a[3577]), .B(n3310), .Z(n3309) );
  IV U3831 ( .A(n3307), .Z(n3310) );
  XOR U3832 ( .A(n3311), .B(n3312), .Z(n3307) );
  ANDN U3833 ( .B(n3313), .A(n3314), .Z(n3311) );
  XNOR U3834 ( .A(b[3576]), .B(n3312), .Z(n3313) );
  XNOR U3835 ( .A(b[3576]), .B(n3314), .Z(c[3576]) );
  XNOR U3836 ( .A(a[3576]), .B(n3315), .Z(n3314) );
  IV U3837 ( .A(n3312), .Z(n3315) );
  XOR U3838 ( .A(n3316), .B(n3317), .Z(n3312) );
  ANDN U3839 ( .B(n3318), .A(n3319), .Z(n3316) );
  XNOR U3840 ( .A(b[3575]), .B(n3317), .Z(n3318) );
  XNOR U3841 ( .A(b[3575]), .B(n3319), .Z(c[3575]) );
  XNOR U3842 ( .A(a[3575]), .B(n3320), .Z(n3319) );
  IV U3843 ( .A(n3317), .Z(n3320) );
  XOR U3844 ( .A(n3321), .B(n3322), .Z(n3317) );
  ANDN U3845 ( .B(n3323), .A(n3324), .Z(n3321) );
  XNOR U3846 ( .A(b[3574]), .B(n3322), .Z(n3323) );
  XNOR U3847 ( .A(b[3574]), .B(n3324), .Z(c[3574]) );
  XNOR U3848 ( .A(a[3574]), .B(n3325), .Z(n3324) );
  IV U3849 ( .A(n3322), .Z(n3325) );
  XOR U3850 ( .A(n3326), .B(n3327), .Z(n3322) );
  ANDN U3851 ( .B(n3328), .A(n3329), .Z(n3326) );
  XNOR U3852 ( .A(b[3573]), .B(n3327), .Z(n3328) );
  XNOR U3853 ( .A(b[3573]), .B(n3329), .Z(c[3573]) );
  XNOR U3854 ( .A(a[3573]), .B(n3330), .Z(n3329) );
  IV U3855 ( .A(n3327), .Z(n3330) );
  XOR U3856 ( .A(n3331), .B(n3332), .Z(n3327) );
  ANDN U3857 ( .B(n3333), .A(n3334), .Z(n3331) );
  XNOR U3858 ( .A(b[3572]), .B(n3332), .Z(n3333) );
  XNOR U3859 ( .A(b[3572]), .B(n3334), .Z(c[3572]) );
  XNOR U3860 ( .A(a[3572]), .B(n3335), .Z(n3334) );
  IV U3861 ( .A(n3332), .Z(n3335) );
  XOR U3862 ( .A(n3336), .B(n3337), .Z(n3332) );
  ANDN U3863 ( .B(n3338), .A(n3339), .Z(n3336) );
  XNOR U3864 ( .A(b[3571]), .B(n3337), .Z(n3338) );
  XNOR U3865 ( .A(b[3571]), .B(n3339), .Z(c[3571]) );
  XNOR U3866 ( .A(a[3571]), .B(n3340), .Z(n3339) );
  IV U3867 ( .A(n3337), .Z(n3340) );
  XOR U3868 ( .A(n3341), .B(n3342), .Z(n3337) );
  ANDN U3869 ( .B(n3343), .A(n3344), .Z(n3341) );
  XNOR U3870 ( .A(b[3570]), .B(n3342), .Z(n3343) );
  XNOR U3871 ( .A(b[3570]), .B(n3344), .Z(c[3570]) );
  XNOR U3872 ( .A(a[3570]), .B(n3345), .Z(n3344) );
  IV U3873 ( .A(n3342), .Z(n3345) );
  XOR U3874 ( .A(n3346), .B(n3347), .Z(n3342) );
  ANDN U3875 ( .B(n3348), .A(n3349), .Z(n3346) );
  XNOR U3876 ( .A(b[3569]), .B(n3347), .Z(n3348) );
  XNOR U3877 ( .A(b[356]), .B(n3350), .Z(c[356]) );
  XNOR U3878 ( .A(b[3569]), .B(n3349), .Z(c[3569]) );
  XNOR U3879 ( .A(a[3569]), .B(n3351), .Z(n3349) );
  IV U3880 ( .A(n3347), .Z(n3351) );
  XOR U3881 ( .A(n3352), .B(n3353), .Z(n3347) );
  ANDN U3882 ( .B(n3354), .A(n3355), .Z(n3352) );
  XNOR U3883 ( .A(b[3568]), .B(n3353), .Z(n3354) );
  XNOR U3884 ( .A(b[3568]), .B(n3355), .Z(c[3568]) );
  XNOR U3885 ( .A(a[3568]), .B(n3356), .Z(n3355) );
  IV U3886 ( .A(n3353), .Z(n3356) );
  XOR U3887 ( .A(n3357), .B(n3358), .Z(n3353) );
  ANDN U3888 ( .B(n3359), .A(n3360), .Z(n3357) );
  XNOR U3889 ( .A(b[3567]), .B(n3358), .Z(n3359) );
  XNOR U3890 ( .A(b[3567]), .B(n3360), .Z(c[3567]) );
  XNOR U3891 ( .A(a[3567]), .B(n3361), .Z(n3360) );
  IV U3892 ( .A(n3358), .Z(n3361) );
  XOR U3893 ( .A(n3362), .B(n3363), .Z(n3358) );
  ANDN U3894 ( .B(n3364), .A(n3365), .Z(n3362) );
  XNOR U3895 ( .A(b[3566]), .B(n3363), .Z(n3364) );
  XNOR U3896 ( .A(b[3566]), .B(n3365), .Z(c[3566]) );
  XNOR U3897 ( .A(a[3566]), .B(n3366), .Z(n3365) );
  IV U3898 ( .A(n3363), .Z(n3366) );
  XOR U3899 ( .A(n3367), .B(n3368), .Z(n3363) );
  ANDN U3900 ( .B(n3369), .A(n3370), .Z(n3367) );
  XNOR U3901 ( .A(b[3565]), .B(n3368), .Z(n3369) );
  XNOR U3902 ( .A(b[3565]), .B(n3370), .Z(c[3565]) );
  XNOR U3903 ( .A(a[3565]), .B(n3371), .Z(n3370) );
  IV U3904 ( .A(n3368), .Z(n3371) );
  XOR U3905 ( .A(n3372), .B(n3373), .Z(n3368) );
  ANDN U3906 ( .B(n3374), .A(n3375), .Z(n3372) );
  XNOR U3907 ( .A(b[3564]), .B(n3373), .Z(n3374) );
  XNOR U3908 ( .A(b[3564]), .B(n3375), .Z(c[3564]) );
  XNOR U3909 ( .A(a[3564]), .B(n3376), .Z(n3375) );
  IV U3910 ( .A(n3373), .Z(n3376) );
  XOR U3911 ( .A(n3377), .B(n3378), .Z(n3373) );
  ANDN U3912 ( .B(n3379), .A(n3380), .Z(n3377) );
  XNOR U3913 ( .A(b[3563]), .B(n3378), .Z(n3379) );
  XNOR U3914 ( .A(b[3563]), .B(n3380), .Z(c[3563]) );
  XNOR U3915 ( .A(a[3563]), .B(n3381), .Z(n3380) );
  IV U3916 ( .A(n3378), .Z(n3381) );
  XOR U3917 ( .A(n3382), .B(n3383), .Z(n3378) );
  ANDN U3918 ( .B(n3384), .A(n3385), .Z(n3382) );
  XNOR U3919 ( .A(b[3562]), .B(n3383), .Z(n3384) );
  XNOR U3920 ( .A(b[3562]), .B(n3385), .Z(c[3562]) );
  XNOR U3921 ( .A(a[3562]), .B(n3386), .Z(n3385) );
  IV U3922 ( .A(n3383), .Z(n3386) );
  XOR U3923 ( .A(n3387), .B(n3388), .Z(n3383) );
  ANDN U3924 ( .B(n3389), .A(n3390), .Z(n3387) );
  XNOR U3925 ( .A(b[3561]), .B(n3388), .Z(n3389) );
  XNOR U3926 ( .A(b[3561]), .B(n3390), .Z(c[3561]) );
  XNOR U3927 ( .A(a[3561]), .B(n3391), .Z(n3390) );
  IV U3928 ( .A(n3388), .Z(n3391) );
  XOR U3929 ( .A(n3392), .B(n3393), .Z(n3388) );
  ANDN U3930 ( .B(n3394), .A(n3395), .Z(n3392) );
  XNOR U3931 ( .A(b[3560]), .B(n3393), .Z(n3394) );
  XNOR U3932 ( .A(b[3560]), .B(n3395), .Z(c[3560]) );
  XNOR U3933 ( .A(a[3560]), .B(n3396), .Z(n3395) );
  IV U3934 ( .A(n3393), .Z(n3396) );
  XOR U3935 ( .A(n3397), .B(n3398), .Z(n3393) );
  ANDN U3936 ( .B(n3399), .A(n3400), .Z(n3397) );
  XNOR U3937 ( .A(b[3559]), .B(n3398), .Z(n3399) );
  XNOR U3938 ( .A(b[355]), .B(n3401), .Z(c[355]) );
  XNOR U3939 ( .A(b[3559]), .B(n3400), .Z(c[3559]) );
  XNOR U3940 ( .A(a[3559]), .B(n3402), .Z(n3400) );
  IV U3941 ( .A(n3398), .Z(n3402) );
  XOR U3942 ( .A(n3403), .B(n3404), .Z(n3398) );
  ANDN U3943 ( .B(n3405), .A(n3406), .Z(n3403) );
  XNOR U3944 ( .A(b[3558]), .B(n3404), .Z(n3405) );
  XNOR U3945 ( .A(b[3558]), .B(n3406), .Z(c[3558]) );
  XNOR U3946 ( .A(a[3558]), .B(n3407), .Z(n3406) );
  IV U3947 ( .A(n3404), .Z(n3407) );
  XOR U3948 ( .A(n3408), .B(n3409), .Z(n3404) );
  ANDN U3949 ( .B(n3410), .A(n3411), .Z(n3408) );
  XNOR U3950 ( .A(b[3557]), .B(n3409), .Z(n3410) );
  XNOR U3951 ( .A(b[3557]), .B(n3411), .Z(c[3557]) );
  XNOR U3952 ( .A(a[3557]), .B(n3412), .Z(n3411) );
  IV U3953 ( .A(n3409), .Z(n3412) );
  XOR U3954 ( .A(n3413), .B(n3414), .Z(n3409) );
  ANDN U3955 ( .B(n3415), .A(n3416), .Z(n3413) );
  XNOR U3956 ( .A(b[3556]), .B(n3414), .Z(n3415) );
  XNOR U3957 ( .A(b[3556]), .B(n3416), .Z(c[3556]) );
  XNOR U3958 ( .A(a[3556]), .B(n3417), .Z(n3416) );
  IV U3959 ( .A(n3414), .Z(n3417) );
  XOR U3960 ( .A(n3418), .B(n3419), .Z(n3414) );
  ANDN U3961 ( .B(n3420), .A(n3421), .Z(n3418) );
  XNOR U3962 ( .A(b[3555]), .B(n3419), .Z(n3420) );
  XNOR U3963 ( .A(b[3555]), .B(n3421), .Z(c[3555]) );
  XNOR U3964 ( .A(a[3555]), .B(n3422), .Z(n3421) );
  IV U3965 ( .A(n3419), .Z(n3422) );
  XOR U3966 ( .A(n3423), .B(n3424), .Z(n3419) );
  ANDN U3967 ( .B(n3425), .A(n3426), .Z(n3423) );
  XNOR U3968 ( .A(b[3554]), .B(n3424), .Z(n3425) );
  XNOR U3969 ( .A(b[3554]), .B(n3426), .Z(c[3554]) );
  XNOR U3970 ( .A(a[3554]), .B(n3427), .Z(n3426) );
  IV U3971 ( .A(n3424), .Z(n3427) );
  XOR U3972 ( .A(n3428), .B(n3429), .Z(n3424) );
  ANDN U3973 ( .B(n3430), .A(n3431), .Z(n3428) );
  XNOR U3974 ( .A(b[3553]), .B(n3429), .Z(n3430) );
  XNOR U3975 ( .A(b[3553]), .B(n3431), .Z(c[3553]) );
  XNOR U3976 ( .A(a[3553]), .B(n3432), .Z(n3431) );
  IV U3977 ( .A(n3429), .Z(n3432) );
  XOR U3978 ( .A(n3433), .B(n3434), .Z(n3429) );
  ANDN U3979 ( .B(n3435), .A(n3436), .Z(n3433) );
  XNOR U3980 ( .A(b[3552]), .B(n3434), .Z(n3435) );
  XNOR U3981 ( .A(b[3552]), .B(n3436), .Z(c[3552]) );
  XNOR U3982 ( .A(a[3552]), .B(n3437), .Z(n3436) );
  IV U3983 ( .A(n3434), .Z(n3437) );
  XOR U3984 ( .A(n3438), .B(n3439), .Z(n3434) );
  ANDN U3985 ( .B(n3440), .A(n3441), .Z(n3438) );
  XNOR U3986 ( .A(b[3551]), .B(n3439), .Z(n3440) );
  XNOR U3987 ( .A(b[3551]), .B(n3441), .Z(c[3551]) );
  XNOR U3988 ( .A(a[3551]), .B(n3442), .Z(n3441) );
  IV U3989 ( .A(n3439), .Z(n3442) );
  XOR U3990 ( .A(n3443), .B(n3444), .Z(n3439) );
  ANDN U3991 ( .B(n3445), .A(n3446), .Z(n3443) );
  XNOR U3992 ( .A(b[3550]), .B(n3444), .Z(n3445) );
  XNOR U3993 ( .A(b[3550]), .B(n3446), .Z(c[3550]) );
  XNOR U3994 ( .A(a[3550]), .B(n3447), .Z(n3446) );
  IV U3995 ( .A(n3444), .Z(n3447) );
  XOR U3996 ( .A(n3448), .B(n3449), .Z(n3444) );
  ANDN U3997 ( .B(n3450), .A(n3451), .Z(n3448) );
  XNOR U3998 ( .A(b[3549]), .B(n3449), .Z(n3450) );
  XNOR U3999 ( .A(b[354]), .B(n3452), .Z(c[354]) );
  XNOR U4000 ( .A(b[3549]), .B(n3451), .Z(c[3549]) );
  XNOR U4001 ( .A(a[3549]), .B(n3453), .Z(n3451) );
  IV U4002 ( .A(n3449), .Z(n3453) );
  XOR U4003 ( .A(n3454), .B(n3455), .Z(n3449) );
  ANDN U4004 ( .B(n3456), .A(n3457), .Z(n3454) );
  XNOR U4005 ( .A(b[3548]), .B(n3455), .Z(n3456) );
  XNOR U4006 ( .A(b[3548]), .B(n3457), .Z(c[3548]) );
  XNOR U4007 ( .A(a[3548]), .B(n3458), .Z(n3457) );
  IV U4008 ( .A(n3455), .Z(n3458) );
  XOR U4009 ( .A(n3459), .B(n3460), .Z(n3455) );
  ANDN U4010 ( .B(n3461), .A(n3462), .Z(n3459) );
  XNOR U4011 ( .A(b[3547]), .B(n3460), .Z(n3461) );
  XNOR U4012 ( .A(b[3547]), .B(n3462), .Z(c[3547]) );
  XNOR U4013 ( .A(a[3547]), .B(n3463), .Z(n3462) );
  IV U4014 ( .A(n3460), .Z(n3463) );
  XOR U4015 ( .A(n3464), .B(n3465), .Z(n3460) );
  ANDN U4016 ( .B(n3466), .A(n3467), .Z(n3464) );
  XNOR U4017 ( .A(b[3546]), .B(n3465), .Z(n3466) );
  XNOR U4018 ( .A(b[3546]), .B(n3467), .Z(c[3546]) );
  XNOR U4019 ( .A(a[3546]), .B(n3468), .Z(n3467) );
  IV U4020 ( .A(n3465), .Z(n3468) );
  XOR U4021 ( .A(n3469), .B(n3470), .Z(n3465) );
  ANDN U4022 ( .B(n3471), .A(n3472), .Z(n3469) );
  XNOR U4023 ( .A(b[3545]), .B(n3470), .Z(n3471) );
  XNOR U4024 ( .A(b[3545]), .B(n3472), .Z(c[3545]) );
  XNOR U4025 ( .A(a[3545]), .B(n3473), .Z(n3472) );
  IV U4026 ( .A(n3470), .Z(n3473) );
  XOR U4027 ( .A(n3474), .B(n3475), .Z(n3470) );
  ANDN U4028 ( .B(n3476), .A(n3477), .Z(n3474) );
  XNOR U4029 ( .A(b[3544]), .B(n3475), .Z(n3476) );
  XNOR U4030 ( .A(b[3544]), .B(n3477), .Z(c[3544]) );
  XNOR U4031 ( .A(a[3544]), .B(n3478), .Z(n3477) );
  IV U4032 ( .A(n3475), .Z(n3478) );
  XOR U4033 ( .A(n3479), .B(n3480), .Z(n3475) );
  ANDN U4034 ( .B(n3481), .A(n3482), .Z(n3479) );
  XNOR U4035 ( .A(b[3543]), .B(n3480), .Z(n3481) );
  XNOR U4036 ( .A(b[3543]), .B(n3482), .Z(c[3543]) );
  XNOR U4037 ( .A(a[3543]), .B(n3483), .Z(n3482) );
  IV U4038 ( .A(n3480), .Z(n3483) );
  XOR U4039 ( .A(n3484), .B(n3485), .Z(n3480) );
  ANDN U4040 ( .B(n3486), .A(n3487), .Z(n3484) );
  XNOR U4041 ( .A(b[3542]), .B(n3485), .Z(n3486) );
  XNOR U4042 ( .A(b[3542]), .B(n3487), .Z(c[3542]) );
  XNOR U4043 ( .A(a[3542]), .B(n3488), .Z(n3487) );
  IV U4044 ( .A(n3485), .Z(n3488) );
  XOR U4045 ( .A(n3489), .B(n3490), .Z(n3485) );
  ANDN U4046 ( .B(n3491), .A(n3492), .Z(n3489) );
  XNOR U4047 ( .A(b[3541]), .B(n3490), .Z(n3491) );
  XNOR U4048 ( .A(b[3541]), .B(n3492), .Z(c[3541]) );
  XNOR U4049 ( .A(a[3541]), .B(n3493), .Z(n3492) );
  IV U4050 ( .A(n3490), .Z(n3493) );
  XOR U4051 ( .A(n3494), .B(n3495), .Z(n3490) );
  ANDN U4052 ( .B(n3496), .A(n3497), .Z(n3494) );
  XNOR U4053 ( .A(b[3540]), .B(n3495), .Z(n3496) );
  XNOR U4054 ( .A(b[3540]), .B(n3497), .Z(c[3540]) );
  XNOR U4055 ( .A(a[3540]), .B(n3498), .Z(n3497) );
  IV U4056 ( .A(n3495), .Z(n3498) );
  XOR U4057 ( .A(n3499), .B(n3500), .Z(n3495) );
  ANDN U4058 ( .B(n3501), .A(n3502), .Z(n3499) );
  XNOR U4059 ( .A(b[3539]), .B(n3500), .Z(n3501) );
  XNOR U4060 ( .A(b[353]), .B(n3503), .Z(c[353]) );
  XNOR U4061 ( .A(b[3539]), .B(n3502), .Z(c[3539]) );
  XNOR U4062 ( .A(a[3539]), .B(n3504), .Z(n3502) );
  IV U4063 ( .A(n3500), .Z(n3504) );
  XOR U4064 ( .A(n3505), .B(n3506), .Z(n3500) );
  ANDN U4065 ( .B(n3507), .A(n3508), .Z(n3505) );
  XNOR U4066 ( .A(b[3538]), .B(n3506), .Z(n3507) );
  XNOR U4067 ( .A(b[3538]), .B(n3508), .Z(c[3538]) );
  XNOR U4068 ( .A(a[3538]), .B(n3509), .Z(n3508) );
  IV U4069 ( .A(n3506), .Z(n3509) );
  XOR U4070 ( .A(n3510), .B(n3511), .Z(n3506) );
  ANDN U4071 ( .B(n3512), .A(n3513), .Z(n3510) );
  XNOR U4072 ( .A(b[3537]), .B(n3511), .Z(n3512) );
  XNOR U4073 ( .A(b[3537]), .B(n3513), .Z(c[3537]) );
  XNOR U4074 ( .A(a[3537]), .B(n3514), .Z(n3513) );
  IV U4075 ( .A(n3511), .Z(n3514) );
  XOR U4076 ( .A(n3515), .B(n3516), .Z(n3511) );
  ANDN U4077 ( .B(n3517), .A(n3518), .Z(n3515) );
  XNOR U4078 ( .A(b[3536]), .B(n3516), .Z(n3517) );
  XNOR U4079 ( .A(b[3536]), .B(n3518), .Z(c[3536]) );
  XNOR U4080 ( .A(a[3536]), .B(n3519), .Z(n3518) );
  IV U4081 ( .A(n3516), .Z(n3519) );
  XOR U4082 ( .A(n3520), .B(n3521), .Z(n3516) );
  ANDN U4083 ( .B(n3522), .A(n3523), .Z(n3520) );
  XNOR U4084 ( .A(b[3535]), .B(n3521), .Z(n3522) );
  XNOR U4085 ( .A(b[3535]), .B(n3523), .Z(c[3535]) );
  XNOR U4086 ( .A(a[3535]), .B(n3524), .Z(n3523) );
  IV U4087 ( .A(n3521), .Z(n3524) );
  XOR U4088 ( .A(n3525), .B(n3526), .Z(n3521) );
  ANDN U4089 ( .B(n3527), .A(n3528), .Z(n3525) );
  XNOR U4090 ( .A(b[3534]), .B(n3526), .Z(n3527) );
  XNOR U4091 ( .A(b[3534]), .B(n3528), .Z(c[3534]) );
  XNOR U4092 ( .A(a[3534]), .B(n3529), .Z(n3528) );
  IV U4093 ( .A(n3526), .Z(n3529) );
  XOR U4094 ( .A(n3530), .B(n3531), .Z(n3526) );
  ANDN U4095 ( .B(n3532), .A(n3533), .Z(n3530) );
  XNOR U4096 ( .A(b[3533]), .B(n3531), .Z(n3532) );
  XNOR U4097 ( .A(b[3533]), .B(n3533), .Z(c[3533]) );
  XNOR U4098 ( .A(a[3533]), .B(n3534), .Z(n3533) );
  IV U4099 ( .A(n3531), .Z(n3534) );
  XOR U4100 ( .A(n3535), .B(n3536), .Z(n3531) );
  ANDN U4101 ( .B(n3537), .A(n3538), .Z(n3535) );
  XNOR U4102 ( .A(b[3532]), .B(n3536), .Z(n3537) );
  XNOR U4103 ( .A(b[3532]), .B(n3538), .Z(c[3532]) );
  XNOR U4104 ( .A(a[3532]), .B(n3539), .Z(n3538) );
  IV U4105 ( .A(n3536), .Z(n3539) );
  XOR U4106 ( .A(n3540), .B(n3541), .Z(n3536) );
  ANDN U4107 ( .B(n3542), .A(n3543), .Z(n3540) );
  XNOR U4108 ( .A(b[3531]), .B(n3541), .Z(n3542) );
  XNOR U4109 ( .A(b[3531]), .B(n3543), .Z(c[3531]) );
  XNOR U4110 ( .A(a[3531]), .B(n3544), .Z(n3543) );
  IV U4111 ( .A(n3541), .Z(n3544) );
  XOR U4112 ( .A(n3545), .B(n3546), .Z(n3541) );
  ANDN U4113 ( .B(n3547), .A(n3548), .Z(n3545) );
  XNOR U4114 ( .A(b[3530]), .B(n3546), .Z(n3547) );
  XNOR U4115 ( .A(b[3530]), .B(n3548), .Z(c[3530]) );
  XNOR U4116 ( .A(a[3530]), .B(n3549), .Z(n3548) );
  IV U4117 ( .A(n3546), .Z(n3549) );
  XOR U4118 ( .A(n3550), .B(n3551), .Z(n3546) );
  ANDN U4119 ( .B(n3552), .A(n3553), .Z(n3550) );
  XNOR U4120 ( .A(b[3529]), .B(n3551), .Z(n3552) );
  XNOR U4121 ( .A(b[352]), .B(n3554), .Z(c[352]) );
  XNOR U4122 ( .A(b[3529]), .B(n3553), .Z(c[3529]) );
  XNOR U4123 ( .A(a[3529]), .B(n3555), .Z(n3553) );
  IV U4124 ( .A(n3551), .Z(n3555) );
  XOR U4125 ( .A(n3556), .B(n3557), .Z(n3551) );
  ANDN U4126 ( .B(n3558), .A(n3559), .Z(n3556) );
  XNOR U4127 ( .A(b[3528]), .B(n3557), .Z(n3558) );
  XNOR U4128 ( .A(b[3528]), .B(n3559), .Z(c[3528]) );
  XNOR U4129 ( .A(a[3528]), .B(n3560), .Z(n3559) );
  IV U4130 ( .A(n3557), .Z(n3560) );
  XOR U4131 ( .A(n3561), .B(n3562), .Z(n3557) );
  ANDN U4132 ( .B(n3563), .A(n3564), .Z(n3561) );
  XNOR U4133 ( .A(b[3527]), .B(n3562), .Z(n3563) );
  XNOR U4134 ( .A(b[3527]), .B(n3564), .Z(c[3527]) );
  XNOR U4135 ( .A(a[3527]), .B(n3565), .Z(n3564) );
  IV U4136 ( .A(n3562), .Z(n3565) );
  XOR U4137 ( .A(n3566), .B(n3567), .Z(n3562) );
  ANDN U4138 ( .B(n3568), .A(n3569), .Z(n3566) );
  XNOR U4139 ( .A(b[3526]), .B(n3567), .Z(n3568) );
  XNOR U4140 ( .A(b[3526]), .B(n3569), .Z(c[3526]) );
  XNOR U4141 ( .A(a[3526]), .B(n3570), .Z(n3569) );
  IV U4142 ( .A(n3567), .Z(n3570) );
  XOR U4143 ( .A(n3571), .B(n3572), .Z(n3567) );
  ANDN U4144 ( .B(n3573), .A(n3574), .Z(n3571) );
  XNOR U4145 ( .A(b[3525]), .B(n3572), .Z(n3573) );
  XNOR U4146 ( .A(b[3525]), .B(n3574), .Z(c[3525]) );
  XNOR U4147 ( .A(a[3525]), .B(n3575), .Z(n3574) );
  IV U4148 ( .A(n3572), .Z(n3575) );
  XOR U4149 ( .A(n3576), .B(n3577), .Z(n3572) );
  ANDN U4150 ( .B(n3578), .A(n3579), .Z(n3576) );
  XNOR U4151 ( .A(b[3524]), .B(n3577), .Z(n3578) );
  XNOR U4152 ( .A(b[3524]), .B(n3579), .Z(c[3524]) );
  XNOR U4153 ( .A(a[3524]), .B(n3580), .Z(n3579) );
  IV U4154 ( .A(n3577), .Z(n3580) );
  XOR U4155 ( .A(n3581), .B(n3582), .Z(n3577) );
  ANDN U4156 ( .B(n3583), .A(n3584), .Z(n3581) );
  XNOR U4157 ( .A(b[3523]), .B(n3582), .Z(n3583) );
  XNOR U4158 ( .A(b[3523]), .B(n3584), .Z(c[3523]) );
  XNOR U4159 ( .A(a[3523]), .B(n3585), .Z(n3584) );
  IV U4160 ( .A(n3582), .Z(n3585) );
  XOR U4161 ( .A(n3586), .B(n3587), .Z(n3582) );
  ANDN U4162 ( .B(n3588), .A(n3589), .Z(n3586) );
  XNOR U4163 ( .A(b[3522]), .B(n3587), .Z(n3588) );
  XNOR U4164 ( .A(b[3522]), .B(n3589), .Z(c[3522]) );
  XNOR U4165 ( .A(a[3522]), .B(n3590), .Z(n3589) );
  IV U4166 ( .A(n3587), .Z(n3590) );
  XOR U4167 ( .A(n3591), .B(n3592), .Z(n3587) );
  ANDN U4168 ( .B(n3593), .A(n3594), .Z(n3591) );
  XNOR U4169 ( .A(b[3521]), .B(n3592), .Z(n3593) );
  XNOR U4170 ( .A(b[3521]), .B(n3594), .Z(c[3521]) );
  XNOR U4171 ( .A(a[3521]), .B(n3595), .Z(n3594) );
  IV U4172 ( .A(n3592), .Z(n3595) );
  XOR U4173 ( .A(n3596), .B(n3597), .Z(n3592) );
  ANDN U4174 ( .B(n3598), .A(n3599), .Z(n3596) );
  XNOR U4175 ( .A(b[3520]), .B(n3597), .Z(n3598) );
  XNOR U4176 ( .A(b[3520]), .B(n3599), .Z(c[3520]) );
  XNOR U4177 ( .A(a[3520]), .B(n3600), .Z(n3599) );
  IV U4178 ( .A(n3597), .Z(n3600) );
  XOR U4179 ( .A(n3601), .B(n3602), .Z(n3597) );
  ANDN U4180 ( .B(n3603), .A(n3604), .Z(n3601) );
  XNOR U4181 ( .A(b[3519]), .B(n3602), .Z(n3603) );
  XNOR U4182 ( .A(b[351]), .B(n3605), .Z(c[351]) );
  XNOR U4183 ( .A(b[3519]), .B(n3604), .Z(c[3519]) );
  XNOR U4184 ( .A(a[3519]), .B(n3606), .Z(n3604) );
  IV U4185 ( .A(n3602), .Z(n3606) );
  XOR U4186 ( .A(n3607), .B(n3608), .Z(n3602) );
  ANDN U4187 ( .B(n3609), .A(n3610), .Z(n3607) );
  XNOR U4188 ( .A(b[3518]), .B(n3608), .Z(n3609) );
  XNOR U4189 ( .A(b[3518]), .B(n3610), .Z(c[3518]) );
  XNOR U4190 ( .A(a[3518]), .B(n3611), .Z(n3610) );
  IV U4191 ( .A(n3608), .Z(n3611) );
  XOR U4192 ( .A(n3612), .B(n3613), .Z(n3608) );
  ANDN U4193 ( .B(n3614), .A(n3615), .Z(n3612) );
  XNOR U4194 ( .A(b[3517]), .B(n3613), .Z(n3614) );
  XNOR U4195 ( .A(b[3517]), .B(n3615), .Z(c[3517]) );
  XNOR U4196 ( .A(a[3517]), .B(n3616), .Z(n3615) );
  IV U4197 ( .A(n3613), .Z(n3616) );
  XOR U4198 ( .A(n3617), .B(n3618), .Z(n3613) );
  ANDN U4199 ( .B(n3619), .A(n3620), .Z(n3617) );
  XNOR U4200 ( .A(b[3516]), .B(n3618), .Z(n3619) );
  XNOR U4201 ( .A(b[3516]), .B(n3620), .Z(c[3516]) );
  XNOR U4202 ( .A(a[3516]), .B(n3621), .Z(n3620) );
  IV U4203 ( .A(n3618), .Z(n3621) );
  XOR U4204 ( .A(n3622), .B(n3623), .Z(n3618) );
  ANDN U4205 ( .B(n3624), .A(n3625), .Z(n3622) );
  XNOR U4206 ( .A(b[3515]), .B(n3623), .Z(n3624) );
  XNOR U4207 ( .A(b[3515]), .B(n3625), .Z(c[3515]) );
  XNOR U4208 ( .A(a[3515]), .B(n3626), .Z(n3625) );
  IV U4209 ( .A(n3623), .Z(n3626) );
  XOR U4210 ( .A(n3627), .B(n3628), .Z(n3623) );
  ANDN U4211 ( .B(n3629), .A(n3630), .Z(n3627) );
  XNOR U4212 ( .A(b[3514]), .B(n3628), .Z(n3629) );
  XNOR U4213 ( .A(b[3514]), .B(n3630), .Z(c[3514]) );
  XNOR U4214 ( .A(a[3514]), .B(n3631), .Z(n3630) );
  IV U4215 ( .A(n3628), .Z(n3631) );
  XOR U4216 ( .A(n3632), .B(n3633), .Z(n3628) );
  ANDN U4217 ( .B(n3634), .A(n3635), .Z(n3632) );
  XNOR U4218 ( .A(b[3513]), .B(n3633), .Z(n3634) );
  XNOR U4219 ( .A(b[3513]), .B(n3635), .Z(c[3513]) );
  XNOR U4220 ( .A(a[3513]), .B(n3636), .Z(n3635) );
  IV U4221 ( .A(n3633), .Z(n3636) );
  XOR U4222 ( .A(n3637), .B(n3638), .Z(n3633) );
  ANDN U4223 ( .B(n3639), .A(n3640), .Z(n3637) );
  XNOR U4224 ( .A(b[3512]), .B(n3638), .Z(n3639) );
  XNOR U4225 ( .A(b[3512]), .B(n3640), .Z(c[3512]) );
  XNOR U4226 ( .A(a[3512]), .B(n3641), .Z(n3640) );
  IV U4227 ( .A(n3638), .Z(n3641) );
  XOR U4228 ( .A(n3642), .B(n3643), .Z(n3638) );
  ANDN U4229 ( .B(n3644), .A(n3645), .Z(n3642) );
  XNOR U4230 ( .A(b[3511]), .B(n3643), .Z(n3644) );
  XNOR U4231 ( .A(b[3511]), .B(n3645), .Z(c[3511]) );
  XNOR U4232 ( .A(a[3511]), .B(n3646), .Z(n3645) );
  IV U4233 ( .A(n3643), .Z(n3646) );
  XOR U4234 ( .A(n3647), .B(n3648), .Z(n3643) );
  ANDN U4235 ( .B(n3649), .A(n3650), .Z(n3647) );
  XNOR U4236 ( .A(b[3510]), .B(n3648), .Z(n3649) );
  XNOR U4237 ( .A(b[3510]), .B(n3650), .Z(c[3510]) );
  XNOR U4238 ( .A(a[3510]), .B(n3651), .Z(n3650) );
  IV U4239 ( .A(n3648), .Z(n3651) );
  XOR U4240 ( .A(n3652), .B(n3653), .Z(n3648) );
  ANDN U4241 ( .B(n3654), .A(n3655), .Z(n3652) );
  XNOR U4242 ( .A(b[3509]), .B(n3653), .Z(n3654) );
  XNOR U4243 ( .A(b[350]), .B(n3656), .Z(c[350]) );
  XNOR U4244 ( .A(b[3509]), .B(n3655), .Z(c[3509]) );
  XNOR U4245 ( .A(a[3509]), .B(n3657), .Z(n3655) );
  IV U4246 ( .A(n3653), .Z(n3657) );
  XOR U4247 ( .A(n3658), .B(n3659), .Z(n3653) );
  ANDN U4248 ( .B(n3660), .A(n3661), .Z(n3658) );
  XNOR U4249 ( .A(b[3508]), .B(n3659), .Z(n3660) );
  XNOR U4250 ( .A(b[3508]), .B(n3661), .Z(c[3508]) );
  XNOR U4251 ( .A(a[3508]), .B(n3662), .Z(n3661) );
  IV U4252 ( .A(n3659), .Z(n3662) );
  XOR U4253 ( .A(n3663), .B(n3664), .Z(n3659) );
  ANDN U4254 ( .B(n3665), .A(n3666), .Z(n3663) );
  XNOR U4255 ( .A(b[3507]), .B(n3664), .Z(n3665) );
  XNOR U4256 ( .A(b[3507]), .B(n3666), .Z(c[3507]) );
  XNOR U4257 ( .A(a[3507]), .B(n3667), .Z(n3666) );
  IV U4258 ( .A(n3664), .Z(n3667) );
  XOR U4259 ( .A(n3668), .B(n3669), .Z(n3664) );
  ANDN U4260 ( .B(n3670), .A(n3671), .Z(n3668) );
  XNOR U4261 ( .A(b[3506]), .B(n3669), .Z(n3670) );
  XNOR U4262 ( .A(b[3506]), .B(n3671), .Z(c[3506]) );
  XNOR U4263 ( .A(a[3506]), .B(n3672), .Z(n3671) );
  IV U4264 ( .A(n3669), .Z(n3672) );
  XOR U4265 ( .A(n3673), .B(n3674), .Z(n3669) );
  ANDN U4266 ( .B(n3675), .A(n3676), .Z(n3673) );
  XNOR U4267 ( .A(b[3505]), .B(n3674), .Z(n3675) );
  XNOR U4268 ( .A(b[3505]), .B(n3676), .Z(c[3505]) );
  XNOR U4269 ( .A(a[3505]), .B(n3677), .Z(n3676) );
  IV U4270 ( .A(n3674), .Z(n3677) );
  XOR U4271 ( .A(n3678), .B(n3679), .Z(n3674) );
  ANDN U4272 ( .B(n3680), .A(n3681), .Z(n3678) );
  XNOR U4273 ( .A(b[3504]), .B(n3679), .Z(n3680) );
  XNOR U4274 ( .A(b[3504]), .B(n3681), .Z(c[3504]) );
  XNOR U4275 ( .A(a[3504]), .B(n3682), .Z(n3681) );
  IV U4276 ( .A(n3679), .Z(n3682) );
  XOR U4277 ( .A(n3683), .B(n3684), .Z(n3679) );
  ANDN U4278 ( .B(n3685), .A(n3686), .Z(n3683) );
  XNOR U4279 ( .A(b[3503]), .B(n3684), .Z(n3685) );
  XNOR U4280 ( .A(b[3503]), .B(n3686), .Z(c[3503]) );
  XNOR U4281 ( .A(a[3503]), .B(n3687), .Z(n3686) );
  IV U4282 ( .A(n3684), .Z(n3687) );
  XOR U4283 ( .A(n3688), .B(n3689), .Z(n3684) );
  ANDN U4284 ( .B(n3690), .A(n3691), .Z(n3688) );
  XNOR U4285 ( .A(b[3502]), .B(n3689), .Z(n3690) );
  XNOR U4286 ( .A(b[3502]), .B(n3691), .Z(c[3502]) );
  XNOR U4287 ( .A(a[3502]), .B(n3692), .Z(n3691) );
  IV U4288 ( .A(n3689), .Z(n3692) );
  XOR U4289 ( .A(n3693), .B(n3694), .Z(n3689) );
  ANDN U4290 ( .B(n3695), .A(n3696), .Z(n3693) );
  XNOR U4291 ( .A(b[3501]), .B(n3694), .Z(n3695) );
  XNOR U4292 ( .A(b[3501]), .B(n3696), .Z(c[3501]) );
  XNOR U4293 ( .A(a[3501]), .B(n3697), .Z(n3696) );
  IV U4294 ( .A(n3694), .Z(n3697) );
  XOR U4295 ( .A(n3698), .B(n3699), .Z(n3694) );
  ANDN U4296 ( .B(n3700), .A(n3701), .Z(n3698) );
  XNOR U4297 ( .A(b[3500]), .B(n3699), .Z(n3700) );
  XNOR U4298 ( .A(b[3500]), .B(n3701), .Z(c[3500]) );
  XNOR U4299 ( .A(a[3500]), .B(n3702), .Z(n3701) );
  IV U4300 ( .A(n3699), .Z(n3702) );
  XOR U4301 ( .A(n3703), .B(n3704), .Z(n3699) );
  ANDN U4302 ( .B(n3705), .A(n3706), .Z(n3703) );
  XNOR U4303 ( .A(b[3499]), .B(n3704), .Z(n3705) );
  XNOR U4304 ( .A(b[34]), .B(n3707), .Z(c[34]) );
  XNOR U4305 ( .A(b[349]), .B(n3708), .Z(c[349]) );
  XNOR U4306 ( .A(b[3499]), .B(n3706), .Z(c[3499]) );
  XNOR U4307 ( .A(a[3499]), .B(n3709), .Z(n3706) );
  IV U4308 ( .A(n3704), .Z(n3709) );
  XOR U4309 ( .A(n3710), .B(n3711), .Z(n3704) );
  ANDN U4310 ( .B(n3712), .A(n3713), .Z(n3710) );
  XNOR U4311 ( .A(b[3498]), .B(n3711), .Z(n3712) );
  XNOR U4312 ( .A(b[3498]), .B(n3713), .Z(c[3498]) );
  XNOR U4313 ( .A(a[3498]), .B(n3714), .Z(n3713) );
  IV U4314 ( .A(n3711), .Z(n3714) );
  XOR U4315 ( .A(n3715), .B(n3716), .Z(n3711) );
  ANDN U4316 ( .B(n3717), .A(n3718), .Z(n3715) );
  XNOR U4317 ( .A(b[3497]), .B(n3716), .Z(n3717) );
  XNOR U4318 ( .A(b[3497]), .B(n3718), .Z(c[3497]) );
  XNOR U4319 ( .A(a[3497]), .B(n3719), .Z(n3718) );
  IV U4320 ( .A(n3716), .Z(n3719) );
  XOR U4321 ( .A(n3720), .B(n3721), .Z(n3716) );
  ANDN U4322 ( .B(n3722), .A(n3723), .Z(n3720) );
  XNOR U4323 ( .A(b[3496]), .B(n3721), .Z(n3722) );
  XNOR U4324 ( .A(b[3496]), .B(n3723), .Z(c[3496]) );
  XNOR U4325 ( .A(a[3496]), .B(n3724), .Z(n3723) );
  IV U4326 ( .A(n3721), .Z(n3724) );
  XOR U4327 ( .A(n3725), .B(n3726), .Z(n3721) );
  ANDN U4328 ( .B(n3727), .A(n3728), .Z(n3725) );
  XNOR U4329 ( .A(b[3495]), .B(n3726), .Z(n3727) );
  XNOR U4330 ( .A(b[3495]), .B(n3728), .Z(c[3495]) );
  XNOR U4331 ( .A(a[3495]), .B(n3729), .Z(n3728) );
  IV U4332 ( .A(n3726), .Z(n3729) );
  XOR U4333 ( .A(n3730), .B(n3731), .Z(n3726) );
  ANDN U4334 ( .B(n3732), .A(n3733), .Z(n3730) );
  XNOR U4335 ( .A(b[3494]), .B(n3731), .Z(n3732) );
  XNOR U4336 ( .A(b[3494]), .B(n3733), .Z(c[3494]) );
  XNOR U4337 ( .A(a[3494]), .B(n3734), .Z(n3733) );
  IV U4338 ( .A(n3731), .Z(n3734) );
  XOR U4339 ( .A(n3735), .B(n3736), .Z(n3731) );
  ANDN U4340 ( .B(n3737), .A(n3738), .Z(n3735) );
  XNOR U4341 ( .A(b[3493]), .B(n3736), .Z(n3737) );
  XNOR U4342 ( .A(b[3493]), .B(n3738), .Z(c[3493]) );
  XNOR U4343 ( .A(a[3493]), .B(n3739), .Z(n3738) );
  IV U4344 ( .A(n3736), .Z(n3739) );
  XOR U4345 ( .A(n3740), .B(n3741), .Z(n3736) );
  ANDN U4346 ( .B(n3742), .A(n3743), .Z(n3740) );
  XNOR U4347 ( .A(b[3492]), .B(n3741), .Z(n3742) );
  XNOR U4348 ( .A(b[3492]), .B(n3743), .Z(c[3492]) );
  XNOR U4349 ( .A(a[3492]), .B(n3744), .Z(n3743) );
  IV U4350 ( .A(n3741), .Z(n3744) );
  XOR U4351 ( .A(n3745), .B(n3746), .Z(n3741) );
  ANDN U4352 ( .B(n3747), .A(n3748), .Z(n3745) );
  XNOR U4353 ( .A(b[3491]), .B(n3746), .Z(n3747) );
  XNOR U4354 ( .A(b[3491]), .B(n3748), .Z(c[3491]) );
  XNOR U4355 ( .A(a[3491]), .B(n3749), .Z(n3748) );
  IV U4356 ( .A(n3746), .Z(n3749) );
  XOR U4357 ( .A(n3750), .B(n3751), .Z(n3746) );
  ANDN U4358 ( .B(n3752), .A(n3753), .Z(n3750) );
  XNOR U4359 ( .A(b[3490]), .B(n3751), .Z(n3752) );
  XNOR U4360 ( .A(b[3490]), .B(n3753), .Z(c[3490]) );
  XNOR U4361 ( .A(a[3490]), .B(n3754), .Z(n3753) );
  IV U4362 ( .A(n3751), .Z(n3754) );
  XOR U4363 ( .A(n3755), .B(n3756), .Z(n3751) );
  ANDN U4364 ( .B(n3757), .A(n3758), .Z(n3755) );
  XNOR U4365 ( .A(b[3489]), .B(n3756), .Z(n3757) );
  XNOR U4366 ( .A(b[348]), .B(n3759), .Z(c[348]) );
  XNOR U4367 ( .A(b[3489]), .B(n3758), .Z(c[3489]) );
  XNOR U4368 ( .A(a[3489]), .B(n3760), .Z(n3758) );
  IV U4369 ( .A(n3756), .Z(n3760) );
  XOR U4370 ( .A(n3761), .B(n3762), .Z(n3756) );
  ANDN U4371 ( .B(n3763), .A(n3764), .Z(n3761) );
  XNOR U4372 ( .A(b[3488]), .B(n3762), .Z(n3763) );
  XNOR U4373 ( .A(b[3488]), .B(n3764), .Z(c[3488]) );
  XNOR U4374 ( .A(a[3488]), .B(n3765), .Z(n3764) );
  IV U4375 ( .A(n3762), .Z(n3765) );
  XOR U4376 ( .A(n3766), .B(n3767), .Z(n3762) );
  ANDN U4377 ( .B(n3768), .A(n3769), .Z(n3766) );
  XNOR U4378 ( .A(b[3487]), .B(n3767), .Z(n3768) );
  XNOR U4379 ( .A(b[3487]), .B(n3769), .Z(c[3487]) );
  XNOR U4380 ( .A(a[3487]), .B(n3770), .Z(n3769) );
  IV U4381 ( .A(n3767), .Z(n3770) );
  XOR U4382 ( .A(n3771), .B(n3772), .Z(n3767) );
  ANDN U4383 ( .B(n3773), .A(n3774), .Z(n3771) );
  XNOR U4384 ( .A(b[3486]), .B(n3772), .Z(n3773) );
  XNOR U4385 ( .A(b[3486]), .B(n3774), .Z(c[3486]) );
  XNOR U4386 ( .A(a[3486]), .B(n3775), .Z(n3774) );
  IV U4387 ( .A(n3772), .Z(n3775) );
  XOR U4388 ( .A(n3776), .B(n3777), .Z(n3772) );
  ANDN U4389 ( .B(n3778), .A(n3779), .Z(n3776) );
  XNOR U4390 ( .A(b[3485]), .B(n3777), .Z(n3778) );
  XNOR U4391 ( .A(b[3485]), .B(n3779), .Z(c[3485]) );
  XNOR U4392 ( .A(a[3485]), .B(n3780), .Z(n3779) );
  IV U4393 ( .A(n3777), .Z(n3780) );
  XOR U4394 ( .A(n3781), .B(n3782), .Z(n3777) );
  ANDN U4395 ( .B(n3783), .A(n3784), .Z(n3781) );
  XNOR U4396 ( .A(b[3484]), .B(n3782), .Z(n3783) );
  XNOR U4397 ( .A(b[3484]), .B(n3784), .Z(c[3484]) );
  XNOR U4398 ( .A(a[3484]), .B(n3785), .Z(n3784) );
  IV U4399 ( .A(n3782), .Z(n3785) );
  XOR U4400 ( .A(n3786), .B(n3787), .Z(n3782) );
  ANDN U4401 ( .B(n3788), .A(n3789), .Z(n3786) );
  XNOR U4402 ( .A(b[3483]), .B(n3787), .Z(n3788) );
  XNOR U4403 ( .A(b[3483]), .B(n3789), .Z(c[3483]) );
  XNOR U4404 ( .A(a[3483]), .B(n3790), .Z(n3789) );
  IV U4405 ( .A(n3787), .Z(n3790) );
  XOR U4406 ( .A(n3791), .B(n3792), .Z(n3787) );
  ANDN U4407 ( .B(n3793), .A(n3794), .Z(n3791) );
  XNOR U4408 ( .A(b[3482]), .B(n3792), .Z(n3793) );
  XNOR U4409 ( .A(b[3482]), .B(n3794), .Z(c[3482]) );
  XNOR U4410 ( .A(a[3482]), .B(n3795), .Z(n3794) );
  IV U4411 ( .A(n3792), .Z(n3795) );
  XOR U4412 ( .A(n3796), .B(n3797), .Z(n3792) );
  ANDN U4413 ( .B(n3798), .A(n3799), .Z(n3796) );
  XNOR U4414 ( .A(b[3481]), .B(n3797), .Z(n3798) );
  XNOR U4415 ( .A(b[3481]), .B(n3799), .Z(c[3481]) );
  XNOR U4416 ( .A(a[3481]), .B(n3800), .Z(n3799) );
  IV U4417 ( .A(n3797), .Z(n3800) );
  XOR U4418 ( .A(n3801), .B(n3802), .Z(n3797) );
  ANDN U4419 ( .B(n3803), .A(n3804), .Z(n3801) );
  XNOR U4420 ( .A(b[3480]), .B(n3802), .Z(n3803) );
  XNOR U4421 ( .A(b[3480]), .B(n3804), .Z(c[3480]) );
  XNOR U4422 ( .A(a[3480]), .B(n3805), .Z(n3804) );
  IV U4423 ( .A(n3802), .Z(n3805) );
  XOR U4424 ( .A(n3806), .B(n3807), .Z(n3802) );
  ANDN U4425 ( .B(n3808), .A(n3809), .Z(n3806) );
  XNOR U4426 ( .A(b[3479]), .B(n3807), .Z(n3808) );
  XNOR U4427 ( .A(b[347]), .B(n3810), .Z(c[347]) );
  XNOR U4428 ( .A(b[3479]), .B(n3809), .Z(c[3479]) );
  XNOR U4429 ( .A(a[3479]), .B(n3811), .Z(n3809) );
  IV U4430 ( .A(n3807), .Z(n3811) );
  XOR U4431 ( .A(n3812), .B(n3813), .Z(n3807) );
  ANDN U4432 ( .B(n3814), .A(n3815), .Z(n3812) );
  XNOR U4433 ( .A(b[3478]), .B(n3813), .Z(n3814) );
  XNOR U4434 ( .A(b[3478]), .B(n3815), .Z(c[3478]) );
  XNOR U4435 ( .A(a[3478]), .B(n3816), .Z(n3815) );
  IV U4436 ( .A(n3813), .Z(n3816) );
  XOR U4437 ( .A(n3817), .B(n3818), .Z(n3813) );
  ANDN U4438 ( .B(n3819), .A(n3820), .Z(n3817) );
  XNOR U4439 ( .A(b[3477]), .B(n3818), .Z(n3819) );
  XNOR U4440 ( .A(b[3477]), .B(n3820), .Z(c[3477]) );
  XNOR U4441 ( .A(a[3477]), .B(n3821), .Z(n3820) );
  IV U4442 ( .A(n3818), .Z(n3821) );
  XOR U4443 ( .A(n3822), .B(n3823), .Z(n3818) );
  ANDN U4444 ( .B(n3824), .A(n3825), .Z(n3822) );
  XNOR U4445 ( .A(b[3476]), .B(n3823), .Z(n3824) );
  XNOR U4446 ( .A(b[3476]), .B(n3825), .Z(c[3476]) );
  XNOR U4447 ( .A(a[3476]), .B(n3826), .Z(n3825) );
  IV U4448 ( .A(n3823), .Z(n3826) );
  XOR U4449 ( .A(n3827), .B(n3828), .Z(n3823) );
  ANDN U4450 ( .B(n3829), .A(n3830), .Z(n3827) );
  XNOR U4451 ( .A(b[3475]), .B(n3828), .Z(n3829) );
  XNOR U4452 ( .A(b[3475]), .B(n3830), .Z(c[3475]) );
  XNOR U4453 ( .A(a[3475]), .B(n3831), .Z(n3830) );
  IV U4454 ( .A(n3828), .Z(n3831) );
  XOR U4455 ( .A(n3832), .B(n3833), .Z(n3828) );
  ANDN U4456 ( .B(n3834), .A(n3835), .Z(n3832) );
  XNOR U4457 ( .A(b[3474]), .B(n3833), .Z(n3834) );
  XNOR U4458 ( .A(b[3474]), .B(n3835), .Z(c[3474]) );
  XNOR U4459 ( .A(a[3474]), .B(n3836), .Z(n3835) );
  IV U4460 ( .A(n3833), .Z(n3836) );
  XOR U4461 ( .A(n3837), .B(n3838), .Z(n3833) );
  ANDN U4462 ( .B(n3839), .A(n3840), .Z(n3837) );
  XNOR U4463 ( .A(b[3473]), .B(n3838), .Z(n3839) );
  XNOR U4464 ( .A(b[3473]), .B(n3840), .Z(c[3473]) );
  XNOR U4465 ( .A(a[3473]), .B(n3841), .Z(n3840) );
  IV U4466 ( .A(n3838), .Z(n3841) );
  XOR U4467 ( .A(n3842), .B(n3843), .Z(n3838) );
  ANDN U4468 ( .B(n3844), .A(n3845), .Z(n3842) );
  XNOR U4469 ( .A(b[3472]), .B(n3843), .Z(n3844) );
  XNOR U4470 ( .A(b[3472]), .B(n3845), .Z(c[3472]) );
  XNOR U4471 ( .A(a[3472]), .B(n3846), .Z(n3845) );
  IV U4472 ( .A(n3843), .Z(n3846) );
  XOR U4473 ( .A(n3847), .B(n3848), .Z(n3843) );
  ANDN U4474 ( .B(n3849), .A(n3850), .Z(n3847) );
  XNOR U4475 ( .A(b[3471]), .B(n3848), .Z(n3849) );
  XNOR U4476 ( .A(b[3471]), .B(n3850), .Z(c[3471]) );
  XNOR U4477 ( .A(a[3471]), .B(n3851), .Z(n3850) );
  IV U4478 ( .A(n3848), .Z(n3851) );
  XOR U4479 ( .A(n3852), .B(n3853), .Z(n3848) );
  ANDN U4480 ( .B(n3854), .A(n3855), .Z(n3852) );
  XNOR U4481 ( .A(b[3470]), .B(n3853), .Z(n3854) );
  XNOR U4482 ( .A(b[3470]), .B(n3855), .Z(c[3470]) );
  XNOR U4483 ( .A(a[3470]), .B(n3856), .Z(n3855) );
  IV U4484 ( .A(n3853), .Z(n3856) );
  XOR U4485 ( .A(n3857), .B(n3858), .Z(n3853) );
  ANDN U4486 ( .B(n3859), .A(n3860), .Z(n3857) );
  XNOR U4487 ( .A(b[3469]), .B(n3858), .Z(n3859) );
  XNOR U4488 ( .A(b[346]), .B(n3861), .Z(c[346]) );
  XNOR U4489 ( .A(b[3469]), .B(n3860), .Z(c[3469]) );
  XNOR U4490 ( .A(a[3469]), .B(n3862), .Z(n3860) );
  IV U4491 ( .A(n3858), .Z(n3862) );
  XOR U4492 ( .A(n3863), .B(n3864), .Z(n3858) );
  ANDN U4493 ( .B(n3865), .A(n3866), .Z(n3863) );
  XNOR U4494 ( .A(b[3468]), .B(n3864), .Z(n3865) );
  XNOR U4495 ( .A(b[3468]), .B(n3866), .Z(c[3468]) );
  XNOR U4496 ( .A(a[3468]), .B(n3867), .Z(n3866) );
  IV U4497 ( .A(n3864), .Z(n3867) );
  XOR U4498 ( .A(n3868), .B(n3869), .Z(n3864) );
  ANDN U4499 ( .B(n3870), .A(n3871), .Z(n3868) );
  XNOR U4500 ( .A(b[3467]), .B(n3869), .Z(n3870) );
  XNOR U4501 ( .A(b[3467]), .B(n3871), .Z(c[3467]) );
  XNOR U4502 ( .A(a[3467]), .B(n3872), .Z(n3871) );
  IV U4503 ( .A(n3869), .Z(n3872) );
  XOR U4504 ( .A(n3873), .B(n3874), .Z(n3869) );
  ANDN U4505 ( .B(n3875), .A(n3876), .Z(n3873) );
  XNOR U4506 ( .A(b[3466]), .B(n3874), .Z(n3875) );
  XNOR U4507 ( .A(b[3466]), .B(n3876), .Z(c[3466]) );
  XNOR U4508 ( .A(a[3466]), .B(n3877), .Z(n3876) );
  IV U4509 ( .A(n3874), .Z(n3877) );
  XOR U4510 ( .A(n3878), .B(n3879), .Z(n3874) );
  ANDN U4511 ( .B(n3880), .A(n3881), .Z(n3878) );
  XNOR U4512 ( .A(b[3465]), .B(n3879), .Z(n3880) );
  XNOR U4513 ( .A(b[3465]), .B(n3881), .Z(c[3465]) );
  XNOR U4514 ( .A(a[3465]), .B(n3882), .Z(n3881) );
  IV U4515 ( .A(n3879), .Z(n3882) );
  XOR U4516 ( .A(n3883), .B(n3884), .Z(n3879) );
  ANDN U4517 ( .B(n3885), .A(n3886), .Z(n3883) );
  XNOR U4518 ( .A(b[3464]), .B(n3884), .Z(n3885) );
  XNOR U4519 ( .A(b[3464]), .B(n3886), .Z(c[3464]) );
  XNOR U4520 ( .A(a[3464]), .B(n3887), .Z(n3886) );
  IV U4521 ( .A(n3884), .Z(n3887) );
  XOR U4522 ( .A(n3888), .B(n3889), .Z(n3884) );
  ANDN U4523 ( .B(n3890), .A(n3891), .Z(n3888) );
  XNOR U4524 ( .A(b[3463]), .B(n3889), .Z(n3890) );
  XNOR U4525 ( .A(b[3463]), .B(n3891), .Z(c[3463]) );
  XNOR U4526 ( .A(a[3463]), .B(n3892), .Z(n3891) );
  IV U4527 ( .A(n3889), .Z(n3892) );
  XOR U4528 ( .A(n3893), .B(n3894), .Z(n3889) );
  ANDN U4529 ( .B(n3895), .A(n3896), .Z(n3893) );
  XNOR U4530 ( .A(b[3462]), .B(n3894), .Z(n3895) );
  XNOR U4531 ( .A(b[3462]), .B(n3896), .Z(c[3462]) );
  XNOR U4532 ( .A(a[3462]), .B(n3897), .Z(n3896) );
  IV U4533 ( .A(n3894), .Z(n3897) );
  XOR U4534 ( .A(n3898), .B(n3899), .Z(n3894) );
  ANDN U4535 ( .B(n3900), .A(n3901), .Z(n3898) );
  XNOR U4536 ( .A(b[3461]), .B(n3899), .Z(n3900) );
  XNOR U4537 ( .A(b[3461]), .B(n3901), .Z(c[3461]) );
  XNOR U4538 ( .A(a[3461]), .B(n3902), .Z(n3901) );
  IV U4539 ( .A(n3899), .Z(n3902) );
  XOR U4540 ( .A(n3903), .B(n3904), .Z(n3899) );
  ANDN U4541 ( .B(n3905), .A(n3906), .Z(n3903) );
  XNOR U4542 ( .A(b[3460]), .B(n3904), .Z(n3905) );
  XNOR U4543 ( .A(b[3460]), .B(n3906), .Z(c[3460]) );
  XNOR U4544 ( .A(a[3460]), .B(n3907), .Z(n3906) );
  IV U4545 ( .A(n3904), .Z(n3907) );
  XOR U4546 ( .A(n3908), .B(n3909), .Z(n3904) );
  ANDN U4547 ( .B(n3910), .A(n3911), .Z(n3908) );
  XNOR U4548 ( .A(b[3459]), .B(n3909), .Z(n3910) );
  XNOR U4549 ( .A(b[345]), .B(n3912), .Z(c[345]) );
  XNOR U4550 ( .A(b[3459]), .B(n3911), .Z(c[3459]) );
  XNOR U4551 ( .A(a[3459]), .B(n3913), .Z(n3911) );
  IV U4552 ( .A(n3909), .Z(n3913) );
  XOR U4553 ( .A(n3914), .B(n3915), .Z(n3909) );
  ANDN U4554 ( .B(n3916), .A(n3917), .Z(n3914) );
  XNOR U4555 ( .A(b[3458]), .B(n3915), .Z(n3916) );
  XNOR U4556 ( .A(b[3458]), .B(n3917), .Z(c[3458]) );
  XNOR U4557 ( .A(a[3458]), .B(n3918), .Z(n3917) );
  IV U4558 ( .A(n3915), .Z(n3918) );
  XOR U4559 ( .A(n3919), .B(n3920), .Z(n3915) );
  ANDN U4560 ( .B(n3921), .A(n3922), .Z(n3919) );
  XNOR U4561 ( .A(b[3457]), .B(n3920), .Z(n3921) );
  XNOR U4562 ( .A(b[3457]), .B(n3922), .Z(c[3457]) );
  XNOR U4563 ( .A(a[3457]), .B(n3923), .Z(n3922) );
  IV U4564 ( .A(n3920), .Z(n3923) );
  XOR U4565 ( .A(n3924), .B(n3925), .Z(n3920) );
  ANDN U4566 ( .B(n3926), .A(n3927), .Z(n3924) );
  XNOR U4567 ( .A(b[3456]), .B(n3925), .Z(n3926) );
  XNOR U4568 ( .A(b[3456]), .B(n3927), .Z(c[3456]) );
  XNOR U4569 ( .A(a[3456]), .B(n3928), .Z(n3927) );
  IV U4570 ( .A(n3925), .Z(n3928) );
  XOR U4571 ( .A(n3929), .B(n3930), .Z(n3925) );
  ANDN U4572 ( .B(n3931), .A(n3932), .Z(n3929) );
  XNOR U4573 ( .A(b[3455]), .B(n3930), .Z(n3931) );
  XNOR U4574 ( .A(b[3455]), .B(n3932), .Z(c[3455]) );
  XNOR U4575 ( .A(a[3455]), .B(n3933), .Z(n3932) );
  IV U4576 ( .A(n3930), .Z(n3933) );
  XOR U4577 ( .A(n3934), .B(n3935), .Z(n3930) );
  ANDN U4578 ( .B(n3936), .A(n3937), .Z(n3934) );
  XNOR U4579 ( .A(b[3454]), .B(n3935), .Z(n3936) );
  XNOR U4580 ( .A(b[3454]), .B(n3937), .Z(c[3454]) );
  XNOR U4581 ( .A(a[3454]), .B(n3938), .Z(n3937) );
  IV U4582 ( .A(n3935), .Z(n3938) );
  XOR U4583 ( .A(n3939), .B(n3940), .Z(n3935) );
  ANDN U4584 ( .B(n3941), .A(n3942), .Z(n3939) );
  XNOR U4585 ( .A(b[3453]), .B(n3940), .Z(n3941) );
  XNOR U4586 ( .A(b[3453]), .B(n3942), .Z(c[3453]) );
  XNOR U4587 ( .A(a[3453]), .B(n3943), .Z(n3942) );
  IV U4588 ( .A(n3940), .Z(n3943) );
  XOR U4589 ( .A(n3944), .B(n3945), .Z(n3940) );
  ANDN U4590 ( .B(n3946), .A(n3947), .Z(n3944) );
  XNOR U4591 ( .A(b[3452]), .B(n3945), .Z(n3946) );
  XNOR U4592 ( .A(b[3452]), .B(n3947), .Z(c[3452]) );
  XNOR U4593 ( .A(a[3452]), .B(n3948), .Z(n3947) );
  IV U4594 ( .A(n3945), .Z(n3948) );
  XOR U4595 ( .A(n3949), .B(n3950), .Z(n3945) );
  ANDN U4596 ( .B(n3951), .A(n3952), .Z(n3949) );
  XNOR U4597 ( .A(b[3451]), .B(n3950), .Z(n3951) );
  XNOR U4598 ( .A(b[3451]), .B(n3952), .Z(c[3451]) );
  XNOR U4599 ( .A(a[3451]), .B(n3953), .Z(n3952) );
  IV U4600 ( .A(n3950), .Z(n3953) );
  XOR U4601 ( .A(n3954), .B(n3955), .Z(n3950) );
  ANDN U4602 ( .B(n3956), .A(n3957), .Z(n3954) );
  XNOR U4603 ( .A(b[3450]), .B(n3955), .Z(n3956) );
  XNOR U4604 ( .A(b[3450]), .B(n3957), .Z(c[3450]) );
  XNOR U4605 ( .A(a[3450]), .B(n3958), .Z(n3957) );
  IV U4606 ( .A(n3955), .Z(n3958) );
  XOR U4607 ( .A(n3959), .B(n3960), .Z(n3955) );
  ANDN U4608 ( .B(n3961), .A(n3962), .Z(n3959) );
  XNOR U4609 ( .A(b[3449]), .B(n3960), .Z(n3961) );
  XNOR U4610 ( .A(b[344]), .B(n3963), .Z(c[344]) );
  XNOR U4611 ( .A(b[3449]), .B(n3962), .Z(c[3449]) );
  XNOR U4612 ( .A(a[3449]), .B(n3964), .Z(n3962) );
  IV U4613 ( .A(n3960), .Z(n3964) );
  XOR U4614 ( .A(n3965), .B(n3966), .Z(n3960) );
  ANDN U4615 ( .B(n3967), .A(n3968), .Z(n3965) );
  XNOR U4616 ( .A(b[3448]), .B(n3966), .Z(n3967) );
  XNOR U4617 ( .A(b[3448]), .B(n3968), .Z(c[3448]) );
  XNOR U4618 ( .A(a[3448]), .B(n3969), .Z(n3968) );
  IV U4619 ( .A(n3966), .Z(n3969) );
  XOR U4620 ( .A(n3970), .B(n3971), .Z(n3966) );
  ANDN U4621 ( .B(n3972), .A(n3973), .Z(n3970) );
  XNOR U4622 ( .A(b[3447]), .B(n3971), .Z(n3972) );
  XNOR U4623 ( .A(b[3447]), .B(n3973), .Z(c[3447]) );
  XNOR U4624 ( .A(a[3447]), .B(n3974), .Z(n3973) );
  IV U4625 ( .A(n3971), .Z(n3974) );
  XOR U4626 ( .A(n3975), .B(n3976), .Z(n3971) );
  ANDN U4627 ( .B(n3977), .A(n3978), .Z(n3975) );
  XNOR U4628 ( .A(b[3446]), .B(n3976), .Z(n3977) );
  XNOR U4629 ( .A(b[3446]), .B(n3978), .Z(c[3446]) );
  XNOR U4630 ( .A(a[3446]), .B(n3979), .Z(n3978) );
  IV U4631 ( .A(n3976), .Z(n3979) );
  XOR U4632 ( .A(n3980), .B(n3981), .Z(n3976) );
  ANDN U4633 ( .B(n3982), .A(n3983), .Z(n3980) );
  XNOR U4634 ( .A(b[3445]), .B(n3981), .Z(n3982) );
  XNOR U4635 ( .A(b[3445]), .B(n3983), .Z(c[3445]) );
  XNOR U4636 ( .A(a[3445]), .B(n3984), .Z(n3983) );
  IV U4637 ( .A(n3981), .Z(n3984) );
  XOR U4638 ( .A(n3985), .B(n3986), .Z(n3981) );
  ANDN U4639 ( .B(n3987), .A(n3988), .Z(n3985) );
  XNOR U4640 ( .A(b[3444]), .B(n3986), .Z(n3987) );
  XNOR U4641 ( .A(b[3444]), .B(n3988), .Z(c[3444]) );
  XNOR U4642 ( .A(a[3444]), .B(n3989), .Z(n3988) );
  IV U4643 ( .A(n3986), .Z(n3989) );
  XOR U4644 ( .A(n3990), .B(n3991), .Z(n3986) );
  ANDN U4645 ( .B(n3992), .A(n3993), .Z(n3990) );
  XNOR U4646 ( .A(b[3443]), .B(n3991), .Z(n3992) );
  XNOR U4647 ( .A(b[3443]), .B(n3993), .Z(c[3443]) );
  XNOR U4648 ( .A(a[3443]), .B(n3994), .Z(n3993) );
  IV U4649 ( .A(n3991), .Z(n3994) );
  XOR U4650 ( .A(n3995), .B(n3996), .Z(n3991) );
  ANDN U4651 ( .B(n3997), .A(n3998), .Z(n3995) );
  XNOR U4652 ( .A(b[3442]), .B(n3996), .Z(n3997) );
  XNOR U4653 ( .A(b[3442]), .B(n3998), .Z(c[3442]) );
  XNOR U4654 ( .A(a[3442]), .B(n3999), .Z(n3998) );
  IV U4655 ( .A(n3996), .Z(n3999) );
  XOR U4656 ( .A(n4000), .B(n4001), .Z(n3996) );
  ANDN U4657 ( .B(n4002), .A(n4003), .Z(n4000) );
  XNOR U4658 ( .A(b[3441]), .B(n4001), .Z(n4002) );
  XNOR U4659 ( .A(b[3441]), .B(n4003), .Z(c[3441]) );
  XNOR U4660 ( .A(a[3441]), .B(n4004), .Z(n4003) );
  IV U4661 ( .A(n4001), .Z(n4004) );
  XOR U4662 ( .A(n4005), .B(n4006), .Z(n4001) );
  ANDN U4663 ( .B(n4007), .A(n4008), .Z(n4005) );
  XNOR U4664 ( .A(b[3440]), .B(n4006), .Z(n4007) );
  XNOR U4665 ( .A(b[3440]), .B(n4008), .Z(c[3440]) );
  XNOR U4666 ( .A(a[3440]), .B(n4009), .Z(n4008) );
  IV U4667 ( .A(n4006), .Z(n4009) );
  XOR U4668 ( .A(n4010), .B(n4011), .Z(n4006) );
  ANDN U4669 ( .B(n4012), .A(n4013), .Z(n4010) );
  XNOR U4670 ( .A(b[3439]), .B(n4011), .Z(n4012) );
  XNOR U4671 ( .A(b[343]), .B(n4014), .Z(c[343]) );
  XNOR U4672 ( .A(b[3439]), .B(n4013), .Z(c[3439]) );
  XNOR U4673 ( .A(a[3439]), .B(n4015), .Z(n4013) );
  IV U4674 ( .A(n4011), .Z(n4015) );
  XOR U4675 ( .A(n4016), .B(n4017), .Z(n4011) );
  ANDN U4676 ( .B(n4018), .A(n4019), .Z(n4016) );
  XNOR U4677 ( .A(b[3438]), .B(n4017), .Z(n4018) );
  XNOR U4678 ( .A(b[3438]), .B(n4019), .Z(c[3438]) );
  XNOR U4679 ( .A(a[3438]), .B(n4020), .Z(n4019) );
  IV U4680 ( .A(n4017), .Z(n4020) );
  XOR U4681 ( .A(n4021), .B(n4022), .Z(n4017) );
  ANDN U4682 ( .B(n4023), .A(n4024), .Z(n4021) );
  XNOR U4683 ( .A(b[3437]), .B(n4022), .Z(n4023) );
  XNOR U4684 ( .A(b[3437]), .B(n4024), .Z(c[3437]) );
  XNOR U4685 ( .A(a[3437]), .B(n4025), .Z(n4024) );
  IV U4686 ( .A(n4022), .Z(n4025) );
  XOR U4687 ( .A(n4026), .B(n4027), .Z(n4022) );
  ANDN U4688 ( .B(n4028), .A(n4029), .Z(n4026) );
  XNOR U4689 ( .A(b[3436]), .B(n4027), .Z(n4028) );
  XNOR U4690 ( .A(b[3436]), .B(n4029), .Z(c[3436]) );
  XNOR U4691 ( .A(a[3436]), .B(n4030), .Z(n4029) );
  IV U4692 ( .A(n4027), .Z(n4030) );
  XOR U4693 ( .A(n4031), .B(n4032), .Z(n4027) );
  ANDN U4694 ( .B(n4033), .A(n4034), .Z(n4031) );
  XNOR U4695 ( .A(b[3435]), .B(n4032), .Z(n4033) );
  XNOR U4696 ( .A(b[3435]), .B(n4034), .Z(c[3435]) );
  XNOR U4697 ( .A(a[3435]), .B(n4035), .Z(n4034) );
  IV U4698 ( .A(n4032), .Z(n4035) );
  XOR U4699 ( .A(n4036), .B(n4037), .Z(n4032) );
  ANDN U4700 ( .B(n4038), .A(n4039), .Z(n4036) );
  XNOR U4701 ( .A(b[3434]), .B(n4037), .Z(n4038) );
  XNOR U4702 ( .A(b[3434]), .B(n4039), .Z(c[3434]) );
  XNOR U4703 ( .A(a[3434]), .B(n4040), .Z(n4039) );
  IV U4704 ( .A(n4037), .Z(n4040) );
  XOR U4705 ( .A(n4041), .B(n4042), .Z(n4037) );
  ANDN U4706 ( .B(n4043), .A(n4044), .Z(n4041) );
  XNOR U4707 ( .A(b[3433]), .B(n4042), .Z(n4043) );
  XNOR U4708 ( .A(b[3433]), .B(n4044), .Z(c[3433]) );
  XNOR U4709 ( .A(a[3433]), .B(n4045), .Z(n4044) );
  IV U4710 ( .A(n4042), .Z(n4045) );
  XOR U4711 ( .A(n4046), .B(n4047), .Z(n4042) );
  ANDN U4712 ( .B(n4048), .A(n4049), .Z(n4046) );
  XNOR U4713 ( .A(b[3432]), .B(n4047), .Z(n4048) );
  XNOR U4714 ( .A(b[3432]), .B(n4049), .Z(c[3432]) );
  XNOR U4715 ( .A(a[3432]), .B(n4050), .Z(n4049) );
  IV U4716 ( .A(n4047), .Z(n4050) );
  XOR U4717 ( .A(n4051), .B(n4052), .Z(n4047) );
  ANDN U4718 ( .B(n4053), .A(n4054), .Z(n4051) );
  XNOR U4719 ( .A(b[3431]), .B(n4052), .Z(n4053) );
  XNOR U4720 ( .A(b[3431]), .B(n4054), .Z(c[3431]) );
  XNOR U4721 ( .A(a[3431]), .B(n4055), .Z(n4054) );
  IV U4722 ( .A(n4052), .Z(n4055) );
  XOR U4723 ( .A(n4056), .B(n4057), .Z(n4052) );
  ANDN U4724 ( .B(n4058), .A(n4059), .Z(n4056) );
  XNOR U4725 ( .A(b[3430]), .B(n4057), .Z(n4058) );
  XNOR U4726 ( .A(b[3430]), .B(n4059), .Z(c[3430]) );
  XNOR U4727 ( .A(a[3430]), .B(n4060), .Z(n4059) );
  IV U4728 ( .A(n4057), .Z(n4060) );
  XOR U4729 ( .A(n4061), .B(n4062), .Z(n4057) );
  ANDN U4730 ( .B(n4063), .A(n4064), .Z(n4061) );
  XNOR U4731 ( .A(b[3429]), .B(n4062), .Z(n4063) );
  XNOR U4732 ( .A(b[342]), .B(n4065), .Z(c[342]) );
  XNOR U4733 ( .A(b[3429]), .B(n4064), .Z(c[3429]) );
  XNOR U4734 ( .A(a[3429]), .B(n4066), .Z(n4064) );
  IV U4735 ( .A(n4062), .Z(n4066) );
  XOR U4736 ( .A(n4067), .B(n4068), .Z(n4062) );
  ANDN U4737 ( .B(n4069), .A(n4070), .Z(n4067) );
  XNOR U4738 ( .A(b[3428]), .B(n4068), .Z(n4069) );
  XNOR U4739 ( .A(b[3428]), .B(n4070), .Z(c[3428]) );
  XNOR U4740 ( .A(a[3428]), .B(n4071), .Z(n4070) );
  IV U4741 ( .A(n4068), .Z(n4071) );
  XOR U4742 ( .A(n4072), .B(n4073), .Z(n4068) );
  ANDN U4743 ( .B(n4074), .A(n4075), .Z(n4072) );
  XNOR U4744 ( .A(b[3427]), .B(n4073), .Z(n4074) );
  XNOR U4745 ( .A(b[3427]), .B(n4075), .Z(c[3427]) );
  XNOR U4746 ( .A(a[3427]), .B(n4076), .Z(n4075) );
  IV U4747 ( .A(n4073), .Z(n4076) );
  XOR U4748 ( .A(n4077), .B(n4078), .Z(n4073) );
  ANDN U4749 ( .B(n4079), .A(n4080), .Z(n4077) );
  XNOR U4750 ( .A(b[3426]), .B(n4078), .Z(n4079) );
  XNOR U4751 ( .A(b[3426]), .B(n4080), .Z(c[3426]) );
  XNOR U4752 ( .A(a[3426]), .B(n4081), .Z(n4080) );
  IV U4753 ( .A(n4078), .Z(n4081) );
  XOR U4754 ( .A(n4082), .B(n4083), .Z(n4078) );
  ANDN U4755 ( .B(n4084), .A(n4085), .Z(n4082) );
  XNOR U4756 ( .A(b[3425]), .B(n4083), .Z(n4084) );
  XNOR U4757 ( .A(b[3425]), .B(n4085), .Z(c[3425]) );
  XNOR U4758 ( .A(a[3425]), .B(n4086), .Z(n4085) );
  IV U4759 ( .A(n4083), .Z(n4086) );
  XOR U4760 ( .A(n4087), .B(n4088), .Z(n4083) );
  ANDN U4761 ( .B(n4089), .A(n4090), .Z(n4087) );
  XNOR U4762 ( .A(b[3424]), .B(n4088), .Z(n4089) );
  XNOR U4763 ( .A(b[3424]), .B(n4090), .Z(c[3424]) );
  XNOR U4764 ( .A(a[3424]), .B(n4091), .Z(n4090) );
  IV U4765 ( .A(n4088), .Z(n4091) );
  XOR U4766 ( .A(n4092), .B(n4093), .Z(n4088) );
  ANDN U4767 ( .B(n4094), .A(n4095), .Z(n4092) );
  XNOR U4768 ( .A(b[3423]), .B(n4093), .Z(n4094) );
  XNOR U4769 ( .A(b[3423]), .B(n4095), .Z(c[3423]) );
  XNOR U4770 ( .A(a[3423]), .B(n4096), .Z(n4095) );
  IV U4771 ( .A(n4093), .Z(n4096) );
  XOR U4772 ( .A(n4097), .B(n4098), .Z(n4093) );
  ANDN U4773 ( .B(n4099), .A(n4100), .Z(n4097) );
  XNOR U4774 ( .A(b[3422]), .B(n4098), .Z(n4099) );
  XNOR U4775 ( .A(b[3422]), .B(n4100), .Z(c[3422]) );
  XNOR U4776 ( .A(a[3422]), .B(n4101), .Z(n4100) );
  IV U4777 ( .A(n4098), .Z(n4101) );
  XOR U4778 ( .A(n4102), .B(n4103), .Z(n4098) );
  ANDN U4779 ( .B(n4104), .A(n4105), .Z(n4102) );
  XNOR U4780 ( .A(b[3421]), .B(n4103), .Z(n4104) );
  XNOR U4781 ( .A(b[3421]), .B(n4105), .Z(c[3421]) );
  XNOR U4782 ( .A(a[3421]), .B(n4106), .Z(n4105) );
  IV U4783 ( .A(n4103), .Z(n4106) );
  XOR U4784 ( .A(n4107), .B(n4108), .Z(n4103) );
  ANDN U4785 ( .B(n4109), .A(n4110), .Z(n4107) );
  XNOR U4786 ( .A(b[3420]), .B(n4108), .Z(n4109) );
  XNOR U4787 ( .A(b[3420]), .B(n4110), .Z(c[3420]) );
  XNOR U4788 ( .A(a[3420]), .B(n4111), .Z(n4110) );
  IV U4789 ( .A(n4108), .Z(n4111) );
  XOR U4790 ( .A(n4112), .B(n4113), .Z(n4108) );
  ANDN U4791 ( .B(n4114), .A(n4115), .Z(n4112) );
  XNOR U4792 ( .A(b[3419]), .B(n4113), .Z(n4114) );
  XNOR U4793 ( .A(b[341]), .B(n4116), .Z(c[341]) );
  XNOR U4794 ( .A(b[3419]), .B(n4115), .Z(c[3419]) );
  XNOR U4795 ( .A(a[3419]), .B(n4117), .Z(n4115) );
  IV U4796 ( .A(n4113), .Z(n4117) );
  XOR U4797 ( .A(n4118), .B(n4119), .Z(n4113) );
  ANDN U4798 ( .B(n4120), .A(n4121), .Z(n4118) );
  XNOR U4799 ( .A(b[3418]), .B(n4119), .Z(n4120) );
  XNOR U4800 ( .A(b[3418]), .B(n4121), .Z(c[3418]) );
  XNOR U4801 ( .A(a[3418]), .B(n4122), .Z(n4121) );
  IV U4802 ( .A(n4119), .Z(n4122) );
  XOR U4803 ( .A(n4123), .B(n4124), .Z(n4119) );
  ANDN U4804 ( .B(n4125), .A(n4126), .Z(n4123) );
  XNOR U4805 ( .A(b[3417]), .B(n4124), .Z(n4125) );
  XNOR U4806 ( .A(b[3417]), .B(n4126), .Z(c[3417]) );
  XNOR U4807 ( .A(a[3417]), .B(n4127), .Z(n4126) );
  IV U4808 ( .A(n4124), .Z(n4127) );
  XOR U4809 ( .A(n4128), .B(n4129), .Z(n4124) );
  ANDN U4810 ( .B(n4130), .A(n4131), .Z(n4128) );
  XNOR U4811 ( .A(b[3416]), .B(n4129), .Z(n4130) );
  XNOR U4812 ( .A(b[3416]), .B(n4131), .Z(c[3416]) );
  XNOR U4813 ( .A(a[3416]), .B(n4132), .Z(n4131) );
  IV U4814 ( .A(n4129), .Z(n4132) );
  XOR U4815 ( .A(n4133), .B(n4134), .Z(n4129) );
  ANDN U4816 ( .B(n4135), .A(n4136), .Z(n4133) );
  XNOR U4817 ( .A(b[3415]), .B(n4134), .Z(n4135) );
  XNOR U4818 ( .A(b[3415]), .B(n4136), .Z(c[3415]) );
  XNOR U4819 ( .A(a[3415]), .B(n4137), .Z(n4136) );
  IV U4820 ( .A(n4134), .Z(n4137) );
  XOR U4821 ( .A(n4138), .B(n4139), .Z(n4134) );
  ANDN U4822 ( .B(n4140), .A(n4141), .Z(n4138) );
  XNOR U4823 ( .A(b[3414]), .B(n4139), .Z(n4140) );
  XNOR U4824 ( .A(b[3414]), .B(n4141), .Z(c[3414]) );
  XNOR U4825 ( .A(a[3414]), .B(n4142), .Z(n4141) );
  IV U4826 ( .A(n4139), .Z(n4142) );
  XOR U4827 ( .A(n4143), .B(n4144), .Z(n4139) );
  ANDN U4828 ( .B(n4145), .A(n4146), .Z(n4143) );
  XNOR U4829 ( .A(b[3413]), .B(n4144), .Z(n4145) );
  XNOR U4830 ( .A(b[3413]), .B(n4146), .Z(c[3413]) );
  XNOR U4831 ( .A(a[3413]), .B(n4147), .Z(n4146) );
  IV U4832 ( .A(n4144), .Z(n4147) );
  XOR U4833 ( .A(n4148), .B(n4149), .Z(n4144) );
  ANDN U4834 ( .B(n4150), .A(n4151), .Z(n4148) );
  XNOR U4835 ( .A(b[3412]), .B(n4149), .Z(n4150) );
  XNOR U4836 ( .A(b[3412]), .B(n4151), .Z(c[3412]) );
  XNOR U4837 ( .A(a[3412]), .B(n4152), .Z(n4151) );
  IV U4838 ( .A(n4149), .Z(n4152) );
  XOR U4839 ( .A(n4153), .B(n4154), .Z(n4149) );
  ANDN U4840 ( .B(n4155), .A(n4156), .Z(n4153) );
  XNOR U4841 ( .A(b[3411]), .B(n4154), .Z(n4155) );
  XNOR U4842 ( .A(b[3411]), .B(n4156), .Z(c[3411]) );
  XNOR U4843 ( .A(a[3411]), .B(n4157), .Z(n4156) );
  IV U4844 ( .A(n4154), .Z(n4157) );
  XOR U4845 ( .A(n4158), .B(n4159), .Z(n4154) );
  ANDN U4846 ( .B(n4160), .A(n4161), .Z(n4158) );
  XNOR U4847 ( .A(b[3410]), .B(n4159), .Z(n4160) );
  XNOR U4848 ( .A(b[3410]), .B(n4161), .Z(c[3410]) );
  XNOR U4849 ( .A(a[3410]), .B(n4162), .Z(n4161) );
  IV U4850 ( .A(n4159), .Z(n4162) );
  XOR U4851 ( .A(n4163), .B(n4164), .Z(n4159) );
  ANDN U4852 ( .B(n4165), .A(n4166), .Z(n4163) );
  XNOR U4853 ( .A(b[3409]), .B(n4164), .Z(n4165) );
  XNOR U4854 ( .A(b[340]), .B(n4167), .Z(c[340]) );
  XNOR U4855 ( .A(b[3409]), .B(n4166), .Z(c[3409]) );
  XNOR U4856 ( .A(a[3409]), .B(n4168), .Z(n4166) );
  IV U4857 ( .A(n4164), .Z(n4168) );
  XOR U4858 ( .A(n4169), .B(n4170), .Z(n4164) );
  ANDN U4859 ( .B(n4171), .A(n4172), .Z(n4169) );
  XNOR U4860 ( .A(b[3408]), .B(n4170), .Z(n4171) );
  XNOR U4861 ( .A(b[3408]), .B(n4172), .Z(c[3408]) );
  XNOR U4862 ( .A(a[3408]), .B(n4173), .Z(n4172) );
  IV U4863 ( .A(n4170), .Z(n4173) );
  XOR U4864 ( .A(n4174), .B(n4175), .Z(n4170) );
  ANDN U4865 ( .B(n4176), .A(n4177), .Z(n4174) );
  XNOR U4866 ( .A(b[3407]), .B(n4175), .Z(n4176) );
  XNOR U4867 ( .A(b[3407]), .B(n4177), .Z(c[3407]) );
  XNOR U4868 ( .A(a[3407]), .B(n4178), .Z(n4177) );
  IV U4869 ( .A(n4175), .Z(n4178) );
  XOR U4870 ( .A(n4179), .B(n4180), .Z(n4175) );
  ANDN U4871 ( .B(n4181), .A(n4182), .Z(n4179) );
  XNOR U4872 ( .A(b[3406]), .B(n4180), .Z(n4181) );
  XNOR U4873 ( .A(b[3406]), .B(n4182), .Z(c[3406]) );
  XNOR U4874 ( .A(a[3406]), .B(n4183), .Z(n4182) );
  IV U4875 ( .A(n4180), .Z(n4183) );
  XOR U4876 ( .A(n4184), .B(n4185), .Z(n4180) );
  ANDN U4877 ( .B(n4186), .A(n4187), .Z(n4184) );
  XNOR U4878 ( .A(b[3405]), .B(n4185), .Z(n4186) );
  XNOR U4879 ( .A(b[3405]), .B(n4187), .Z(c[3405]) );
  XNOR U4880 ( .A(a[3405]), .B(n4188), .Z(n4187) );
  IV U4881 ( .A(n4185), .Z(n4188) );
  XOR U4882 ( .A(n4189), .B(n4190), .Z(n4185) );
  ANDN U4883 ( .B(n4191), .A(n4192), .Z(n4189) );
  XNOR U4884 ( .A(b[3404]), .B(n4190), .Z(n4191) );
  XNOR U4885 ( .A(b[3404]), .B(n4192), .Z(c[3404]) );
  XNOR U4886 ( .A(a[3404]), .B(n4193), .Z(n4192) );
  IV U4887 ( .A(n4190), .Z(n4193) );
  XOR U4888 ( .A(n4194), .B(n4195), .Z(n4190) );
  ANDN U4889 ( .B(n4196), .A(n4197), .Z(n4194) );
  XNOR U4890 ( .A(b[3403]), .B(n4195), .Z(n4196) );
  XNOR U4891 ( .A(b[3403]), .B(n4197), .Z(c[3403]) );
  XNOR U4892 ( .A(a[3403]), .B(n4198), .Z(n4197) );
  IV U4893 ( .A(n4195), .Z(n4198) );
  XOR U4894 ( .A(n4199), .B(n4200), .Z(n4195) );
  ANDN U4895 ( .B(n4201), .A(n4202), .Z(n4199) );
  XNOR U4896 ( .A(b[3402]), .B(n4200), .Z(n4201) );
  XNOR U4897 ( .A(b[3402]), .B(n4202), .Z(c[3402]) );
  XNOR U4898 ( .A(a[3402]), .B(n4203), .Z(n4202) );
  IV U4899 ( .A(n4200), .Z(n4203) );
  XOR U4900 ( .A(n4204), .B(n4205), .Z(n4200) );
  ANDN U4901 ( .B(n4206), .A(n4207), .Z(n4204) );
  XNOR U4902 ( .A(b[3401]), .B(n4205), .Z(n4206) );
  XNOR U4903 ( .A(b[3401]), .B(n4207), .Z(c[3401]) );
  XNOR U4904 ( .A(a[3401]), .B(n4208), .Z(n4207) );
  IV U4905 ( .A(n4205), .Z(n4208) );
  XOR U4906 ( .A(n4209), .B(n4210), .Z(n4205) );
  ANDN U4907 ( .B(n4211), .A(n4212), .Z(n4209) );
  XNOR U4908 ( .A(b[3400]), .B(n4210), .Z(n4211) );
  XNOR U4909 ( .A(b[3400]), .B(n4212), .Z(c[3400]) );
  XNOR U4910 ( .A(a[3400]), .B(n4213), .Z(n4212) );
  IV U4911 ( .A(n4210), .Z(n4213) );
  XOR U4912 ( .A(n4214), .B(n4215), .Z(n4210) );
  ANDN U4913 ( .B(n4216), .A(n4217), .Z(n4214) );
  XNOR U4914 ( .A(b[3399]), .B(n4215), .Z(n4216) );
  XNOR U4915 ( .A(b[33]), .B(n4218), .Z(c[33]) );
  XNOR U4916 ( .A(b[339]), .B(n4219), .Z(c[339]) );
  XNOR U4917 ( .A(b[3399]), .B(n4217), .Z(c[3399]) );
  XNOR U4918 ( .A(a[3399]), .B(n4220), .Z(n4217) );
  IV U4919 ( .A(n4215), .Z(n4220) );
  XOR U4920 ( .A(n4221), .B(n4222), .Z(n4215) );
  ANDN U4921 ( .B(n4223), .A(n4224), .Z(n4221) );
  XNOR U4922 ( .A(b[3398]), .B(n4222), .Z(n4223) );
  XNOR U4923 ( .A(b[3398]), .B(n4224), .Z(c[3398]) );
  XNOR U4924 ( .A(a[3398]), .B(n4225), .Z(n4224) );
  IV U4925 ( .A(n4222), .Z(n4225) );
  XOR U4926 ( .A(n4226), .B(n4227), .Z(n4222) );
  ANDN U4927 ( .B(n4228), .A(n4229), .Z(n4226) );
  XNOR U4928 ( .A(b[3397]), .B(n4227), .Z(n4228) );
  XNOR U4929 ( .A(b[3397]), .B(n4229), .Z(c[3397]) );
  XNOR U4930 ( .A(a[3397]), .B(n4230), .Z(n4229) );
  IV U4931 ( .A(n4227), .Z(n4230) );
  XOR U4932 ( .A(n4231), .B(n4232), .Z(n4227) );
  ANDN U4933 ( .B(n4233), .A(n4234), .Z(n4231) );
  XNOR U4934 ( .A(b[3396]), .B(n4232), .Z(n4233) );
  XNOR U4935 ( .A(b[3396]), .B(n4234), .Z(c[3396]) );
  XNOR U4936 ( .A(a[3396]), .B(n4235), .Z(n4234) );
  IV U4937 ( .A(n4232), .Z(n4235) );
  XOR U4938 ( .A(n4236), .B(n4237), .Z(n4232) );
  ANDN U4939 ( .B(n4238), .A(n4239), .Z(n4236) );
  XNOR U4940 ( .A(b[3395]), .B(n4237), .Z(n4238) );
  XNOR U4941 ( .A(b[3395]), .B(n4239), .Z(c[3395]) );
  XNOR U4942 ( .A(a[3395]), .B(n4240), .Z(n4239) );
  IV U4943 ( .A(n4237), .Z(n4240) );
  XOR U4944 ( .A(n4241), .B(n4242), .Z(n4237) );
  ANDN U4945 ( .B(n4243), .A(n4244), .Z(n4241) );
  XNOR U4946 ( .A(b[3394]), .B(n4242), .Z(n4243) );
  XNOR U4947 ( .A(b[3394]), .B(n4244), .Z(c[3394]) );
  XNOR U4948 ( .A(a[3394]), .B(n4245), .Z(n4244) );
  IV U4949 ( .A(n4242), .Z(n4245) );
  XOR U4950 ( .A(n4246), .B(n4247), .Z(n4242) );
  ANDN U4951 ( .B(n4248), .A(n4249), .Z(n4246) );
  XNOR U4952 ( .A(b[3393]), .B(n4247), .Z(n4248) );
  XNOR U4953 ( .A(b[3393]), .B(n4249), .Z(c[3393]) );
  XNOR U4954 ( .A(a[3393]), .B(n4250), .Z(n4249) );
  IV U4955 ( .A(n4247), .Z(n4250) );
  XOR U4956 ( .A(n4251), .B(n4252), .Z(n4247) );
  ANDN U4957 ( .B(n4253), .A(n4254), .Z(n4251) );
  XNOR U4958 ( .A(b[3392]), .B(n4252), .Z(n4253) );
  XNOR U4959 ( .A(b[3392]), .B(n4254), .Z(c[3392]) );
  XNOR U4960 ( .A(a[3392]), .B(n4255), .Z(n4254) );
  IV U4961 ( .A(n4252), .Z(n4255) );
  XOR U4962 ( .A(n4256), .B(n4257), .Z(n4252) );
  ANDN U4963 ( .B(n4258), .A(n4259), .Z(n4256) );
  XNOR U4964 ( .A(b[3391]), .B(n4257), .Z(n4258) );
  XNOR U4965 ( .A(b[3391]), .B(n4259), .Z(c[3391]) );
  XNOR U4966 ( .A(a[3391]), .B(n4260), .Z(n4259) );
  IV U4967 ( .A(n4257), .Z(n4260) );
  XOR U4968 ( .A(n4261), .B(n4262), .Z(n4257) );
  ANDN U4969 ( .B(n4263), .A(n4264), .Z(n4261) );
  XNOR U4970 ( .A(b[3390]), .B(n4262), .Z(n4263) );
  XNOR U4971 ( .A(b[3390]), .B(n4264), .Z(c[3390]) );
  XNOR U4972 ( .A(a[3390]), .B(n4265), .Z(n4264) );
  IV U4973 ( .A(n4262), .Z(n4265) );
  XOR U4974 ( .A(n4266), .B(n4267), .Z(n4262) );
  ANDN U4975 ( .B(n4268), .A(n4269), .Z(n4266) );
  XNOR U4976 ( .A(b[3389]), .B(n4267), .Z(n4268) );
  XNOR U4977 ( .A(b[338]), .B(n4270), .Z(c[338]) );
  XNOR U4978 ( .A(b[3389]), .B(n4269), .Z(c[3389]) );
  XNOR U4979 ( .A(a[3389]), .B(n4271), .Z(n4269) );
  IV U4980 ( .A(n4267), .Z(n4271) );
  XOR U4981 ( .A(n4272), .B(n4273), .Z(n4267) );
  ANDN U4982 ( .B(n4274), .A(n4275), .Z(n4272) );
  XNOR U4983 ( .A(b[3388]), .B(n4273), .Z(n4274) );
  XNOR U4984 ( .A(b[3388]), .B(n4275), .Z(c[3388]) );
  XNOR U4985 ( .A(a[3388]), .B(n4276), .Z(n4275) );
  IV U4986 ( .A(n4273), .Z(n4276) );
  XOR U4987 ( .A(n4277), .B(n4278), .Z(n4273) );
  ANDN U4988 ( .B(n4279), .A(n4280), .Z(n4277) );
  XNOR U4989 ( .A(b[3387]), .B(n4278), .Z(n4279) );
  XNOR U4990 ( .A(b[3387]), .B(n4280), .Z(c[3387]) );
  XNOR U4991 ( .A(a[3387]), .B(n4281), .Z(n4280) );
  IV U4992 ( .A(n4278), .Z(n4281) );
  XOR U4993 ( .A(n4282), .B(n4283), .Z(n4278) );
  ANDN U4994 ( .B(n4284), .A(n4285), .Z(n4282) );
  XNOR U4995 ( .A(b[3386]), .B(n4283), .Z(n4284) );
  XNOR U4996 ( .A(b[3386]), .B(n4285), .Z(c[3386]) );
  XNOR U4997 ( .A(a[3386]), .B(n4286), .Z(n4285) );
  IV U4998 ( .A(n4283), .Z(n4286) );
  XOR U4999 ( .A(n4287), .B(n4288), .Z(n4283) );
  ANDN U5000 ( .B(n4289), .A(n4290), .Z(n4287) );
  XNOR U5001 ( .A(b[3385]), .B(n4288), .Z(n4289) );
  XNOR U5002 ( .A(b[3385]), .B(n4290), .Z(c[3385]) );
  XNOR U5003 ( .A(a[3385]), .B(n4291), .Z(n4290) );
  IV U5004 ( .A(n4288), .Z(n4291) );
  XOR U5005 ( .A(n4292), .B(n4293), .Z(n4288) );
  ANDN U5006 ( .B(n4294), .A(n4295), .Z(n4292) );
  XNOR U5007 ( .A(b[3384]), .B(n4293), .Z(n4294) );
  XNOR U5008 ( .A(b[3384]), .B(n4295), .Z(c[3384]) );
  XNOR U5009 ( .A(a[3384]), .B(n4296), .Z(n4295) );
  IV U5010 ( .A(n4293), .Z(n4296) );
  XOR U5011 ( .A(n4297), .B(n4298), .Z(n4293) );
  ANDN U5012 ( .B(n4299), .A(n4300), .Z(n4297) );
  XNOR U5013 ( .A(b[3383]), .B(n4298), .Z(n4299) );
  XNOR U5014 ( .A(b[3383]), .B(n4300), .Z(c[3383]) );
  XNOR U5015 ( .A(a[3383]), .B(n4301), .Z(n4300) );
  IV U5016 ( .A(n4298), .Z(n4301) );
  XOR U5017 ( .A(n4302), .B(n4303), .Z(n4298) );
  ANDN U5018 ( .B(n4304), .A(n4305), .Z(n4302) );
  XNOR U5019 ( .A(b[3382]), .B(n4303), .Z(n4304) );
  XNOR U5020 ( .A(b[3382]), .B(n4305), .Z(c[3382]) );
  XNOR U5021 ( .A(a[3382]), .B(n4306), .Z(n4305) );
  IV U5022 ( .A(n4303), .Z(n4306) );
  XOR U5023 ( .A(n4307), .B(n4308), .Z(n4303) );
  ANDN U5024 ( .B(n4309), .A(n4310), .Z(n4307) );
  XNOR U5025 ( .A(b[3381]), .B(n4308), .Z(n4309) );
  XNOR U5026 ( .A(b[3381]), .B(n4310), .Z(c[3381]) );
  XNOR U5027 ( .A(a[3381]), .B(n4311), .Z(n4310) );
  IV U5028 ( .A(n4308), .Z(n4311) );
  XOR U5029 ( .A(n4312), .B(n4313), .Z(n4308) );
  ANDN U5030 ( .B(n4314), .A(n4315), .Z(n4312) );
  XNOR U5031 ( .A(b[3380]), .B(n4313), .Z(n4314) );
  XNOR U5032 ( .A(b[3380]), .B(n4315), .Z(c[3380]) );
  XNOR U5033 ( .A(a[3380]), .B(n4316), .Z(n4315) );
  IV U5034 ( .A(n4313), .Z(n4316) );
  XOR U5035 ( .A(n4317), .B(n4318), .Z(n4313) );
  ANDN U5036 ( .B(n4319), .A(n4320), .Z(n4317) );
  XNOR U5037 ( .A(b[3379]), .B(n4318), .Z(n4319) );
  XNOR U5038 ( .A(b[337]), .B(n4321), .Z(c[337]) );
  XNOR U5039 ( .A(b[3379]), .B(n4320), .Z(c[3379]) );
  XNOR U5040 ( .A(a[3379]), .B(n4322), .Z(n4320) );
  IV U5041 ( .A(n4318), .Z(n4322) );
  XOR U5042 ( .A(n4323), .B(n4324), .Z(n4318) );
  ANDN U5043 ( .B(n4325), .A(n4326), .Z(n4323) );
  XNOR U5044 ( .A(b[3378]), .B(n4324), .Z(n4325) );
  XNOR U5045 ( .A(b[3378]), .B(n4326), .Z(c[3378]) );
  XNOR U5046 ( .A(a[3378]), .B(n4327), .Z(n4326) );
  IV U5047 ( .A(n4324), .Z(n4327) );
  XOR U5048 ( .A(n4328), .B(n4329), .Z(n4324) );
  ANDN U5049 ( .B(n4330), .A(n4331), .Z(n4328) );
  XNOR U5050 ( .A(b[3377]), .B(n4329), .Z(n4330) );
  XNOR U5051 ( .A(b[3377]), .B(n4331), .Z(c[3377]) );
  XNOR U5052 ( .A(a[3377]), .B(n4332), .Z(n4331) );
  IV U5053 ( .A(n4329), .Z(n4332) );
  XOR U5054 ( .A(n4333), .B(n4334), .Z(n4329) );
  ANDN U5055 ( .B(n4335), .A(n4336), .Z(n4333) );
  XNOR U5056 ( .A(b[3376]), .B(n4334), .Z(n4335) );
  XNOR U5057 ( .A(b[3376]), .B(n4336), .Z(c[3376]) );
  XNOR U5058 ( .A(a[3376]), .B(n4337), .Z(n4336) );
  IV U5059 ( .A(n4334), .Z(n4337) );
  XOR U5060 ( .A(n4338), .B(n4339), .Z(n4334) );
  ANDN U5061 ( .B(n4340), .A(n4341), .Z(n4338) );
  XNOR U5062 ( .A(b[3375]), .B(n4339), .Z(n4340) );
  XNOR U5063 ( .A(b[3375]), .B(n4341), .Z(c[3375]) );
  XNOR U5064 ( .A(a[3375]), .B(n4342), .Z(n4341) );
  IV U5065 ( .A(n4339), .Z(n4342) );
  XOR U5066 ( .A(n4343), .B(n4344), .Z(n4339) );
  ANDN U5067 ( .B(n4345), .A(n4346), .Z(n4343) );
  XNOR U5068 ( .A(b[3374]), .B(n4344), .Z(n4345) );
  XNOR U5069 ( .A(b[3374]), .B(n4346), .Z(c[3374]) );
  XNOR U5070 ( .A(a[3374]), .B(n4347), .Z(n4346) );
  IV U5071 ( .A(n4344), .Z(n4347) );
  XOR U5072 ( .A(n4348), .B(n4349), .Z(n4344) );
  ANDN U5073 ( .B(n4350), .A(n4351), .Z(n4348) );
  XNOR U5074 ( .A(b[3373]), .B(n4349), .Z(n4350) );
  XNOR U5075 ( .A(b[3373]), .B(n4351), .Z(c[3373]) );
  XNOR U5076 ( .A(a[3373]), .B(n4352), .Z(n4351) );
  IV U5077 ( .A(n4349), .Z(n4352) );
  XOR U5078 ( .A(n4353), .B(n4354), .Z(n4349) );
  ANDN U5079 ( .B(n4355), .A(n4356), .Z(n4353) );
  XNOR U5080 ( .A(b[3372]), .B(n4354), .Z(n4355) );
  XNOR U5081 ( .A(b[3372]), .B(n4356), .Z(c[3372]) );
  XNOR U5082 ( .A(a[3372]), .B(n4357), .Z(n4356) );
  IV U5083 ( .A(n4354), .Z(n4357) );
  XOR U5084 ( .A(n4358), .B(n4359), .Z(n4354) );
  ANDN U5085 ( .B(n4360), .A(n4361), .Z(n4358) );
  XNOR U5086 ( .A(b[3371]), .B(n4359), .Z(n4360) );
  XNOR U5087 ( .A(b[3371]), .B(n4361), .Z(c[3371]) );
  XNOR U5088 ( .A(a[3371]), .B(n4362), .Z(n4361) );
  IV U5089 ( .A(n4359), .Z(n4362) );
  XOR U5090 ( .A(n4363), .B(n4364), .Z(n4359) );
  ANDN U5091 ( .B(n4365), .A(n4366), .Z(n4363) );
  XNOR U5092 ( .A(b[3370]), .B(n4364), .Z(n4365) );
  XNOR U5093 ( .A(b[3370]), .B(n4366), .Z(c[3370]) );
  XNOR U5094 ( .A(a[3370]), .B(n4367), .Z(n4366) );
  IV U5095 ( .A(n4364), .Z(n4367) );
  XOR U5096 ( .A(n4368), .B(n4369), .Z(n4364) );
  ANDN U5097 ( .B(n4370), .A(n4371), .Z(n4368) );
  XNOR U5098 ( .A(b[3369]), .B(n4369), .Z(n4370) );
  XNOR U5099 ( .A(b[336]), .B(n4372), .Z(c[336]) );
  XNOR U5100 ( .A(b[3369]), .B(n4371), .Z(c[3369]) );
  XNOR U5101 ( .A(a[3369]), .B(n4373), .Z(n4371) );
  IV U5102 ( .A(n4369), .Z(n4373) );
  XOR U5103 ( .A(n4374), .B(n4375), .Z(n4369) );
  ANDN U5104 ( .B(n4376), .A(n4377), .Z(n4374) );
  XNOR U5105 ( .A(b[3368]), .B(n4375), .Z(n4376) );
  XNOR U5106 ( .A(b[3368]), .B(n4377), .Z(c[3368]) );
  XNOR U5107 ( .A(a[3368]), .B(n4378), .Z(n4377) );
  IV U5108 ( .A(n4375), .Z(n4378) );
  XOR U5109 ( .A(n4379), .B(n4380), .Z(n4375) );
  ANDN U5110 ( .B(n4381), .A(n4382), .Z(n4379) );
  XNOR U5111 ( .A(b[3367]), .B(n4380), .Z(n4381) );
  XNOR U5112 ( .A(b[3367]), .B(n4382), .Z(c[3367]) );
  XNOR U5113 ( .A(a[3367]), .B(n4383), .Z(n4382) );
  IV U5114 ( .A(n4380), .Z(n4383) );
  XOR U5115 ( .A(n4384), .B(n4385), .Z(n4380) );
  ANDN U5116 ( .B(n4386), .A(n4387), .Z(n4384) );
  XNOR U5117 ( .A(b[3366]), .B(n4385), .Z(n4386) );
  XNOR U5118 ( .A(b[3366]), .B(n4387), .Z(c[3366]) );
  XNOR U5119 ( .A(a[3366]), .B(n4388), .Z(n4387) );
  IV U5120 ( .A(n4385), .Z(n4388) );
  XOR U5121 ( .A(n4389), .B(n4390), .Z(n4385) );
  ANDN U5122 ( .B(n4391), .A(n4392), .Z(n4389) );
  XNOR U5123 ( .A(b[3365]), .B(n4390), .Z(n4391) );
  XNOR U5124 ( .A(b[3365]), .B(n4392), .Z(c[3365]) );
  XNOR U5125 ( .A(a[3365]), .B(n4393), .Z(n4392) );
  IV U5126 ( .A(n4390), .Z(n4393) );
  XOR U5127 ( .A(n4394), .B(n4395), .Z(n4390) );
  ANDN U5128 ( .B(n4396), .A(n4397), .Z(n4394) );
  XNOR U5129 ( .A(b[3364]), .B(n4395), .Z(n4396) );
  XNOR U5130 ( .A(b[3364]), .B(n4397), .Z(c[3364]) );
  XNOR U5131 ( .A(a[3364]), .B(n4398), .Z(n4397) );
  IV U5132 ( .A(n4395), .Z(n4398) );
  XOR U5133 ( .A(n4399), .B(n4400), .Z(n4395) );
  ANDN U5134 ( .B(n4401), .A(n4402), .Z(n4399) );
  XNOR U5135 ( .A(b[3363]), .B(n4400), .Z(n4401) );
  XNOR U5136 ( .A(b[3363]), .B(n4402), .Z(c[3363]) );
  XNOR U5137 ( .A(a[3363]), .B(n4403), .Z(n4402) );
  IV U5138 ( .A(n4400), .Z(n4403) );
  XOR U5139 ( .A(n4404), .B(n4405), .Z(n4400) );
  ANDN U5140 ( .B(n4406), .A(n4407), .Z(n4404) );
  XNOR U5141 ( .A(b[3362]), .B(n4405), .Z(n4406) );
  XNOR U5142 ( .A(b[3362]), .B(n4407), .Z(c[3362]) );
  XNOR U5143 ( .A(a[3362]), .B(n4408), .Z(n4407) );
  IV U5144 ( .A(n4405), .Z(n4408) );
  XOR U5145 ( .A(n4409), .B(n4410), .Z(n4405) );
  ANDN U5146 ( .B(n4411), .A(n4412), .Z(n4409) );
  XNOR U5147 ( .A(b[3361]), .B(n4410), .Z(n4411) );
  XNOR U5148 ( .A(b[3361]), .B(n4412), .Z(c[3361]) );
  XNOR U5149 ( .A(a[3361]), .B(n4413), .Z(n4412) );
  IV U5150 ( .A(n4410), .Z(n4413) );
  XOR U5151 ( .A(n4414), .B(n4415), .Z(n4410) );
  ANDN U5152 ( .B(n4416), .A(n4417), .Z(n4414) );
  XNOR U5153 ( .A(b[3360]), .B(n4415), .Z(n4416) );
  XNOR U5154 ( .A(b[3360]), .B(n4417), .Z(c[3360]) );
  XNOR U5155 ( .A(a[3360]), .B(n4418), .Z(n4417) );
  IV U5156 ( .A(n4415), .Z(n4418) );
  XOR U5157 ( .A(n4419), .B(n4420), .Z(n4415) );
  ANDN U5158 ( .B(n4421), .A(n4422), .Z(n4419) );
  XNOR U5159 ( .A(b[3359]), .B(n4420), .Z(n4421) );
  XNOR U5160 ( .A(b[335]), .B(n4423), .Z(c[335]) );
  XNOR U5161 ( .A(b[3359]), .B(n4422), .Z(c[3359]) );
  XNOR U5162 ( .A(a[3359]), .B(n4424), .Z(n4422) );
  IV U5163 ( .A(n4420), .Z(n4424) );
  XOR U5164 ( .A(n4425), .B(n4426), .Z(n4420) );
  ANDN U5165 ( .B(n4427), .A(n4428), .Z(n4425) );
  XNOR U5166 ( .A(b[3358]), .B(n4426), .Z(n4427) );
  XNOR U5167 ( .A(b[3358]), .B(n4428), .Z(c[3358]) );
  XNOR U5168 ( .A(a[3358]), .B(n4429), .Z(n4428) );
  IV U5169 ( .A(n4426), .Z(n4429) );
  XOR U5170 ( .A(n4430), .B(n4431), .Z(n4426) );
  ANDN U5171 ( .B(n4432), .A(n4433), .Z(n4430) );
  XNOR U5172 ( .A(b[3357]), .B(n4431), .Z(n4432) );
  XNOR U5173 ( .A(b[3357]), .B(n4433), .Z(c[3357]) );
  XNOR U5174 ( .A(a[3357]), .B(n4434), .Z(n4433) );
  IV U5175 ( .A(n4431), .Z(n4434) );
  XOR U5176 ( .A(n4435), .B(n4436), .Z(n4431) );
  ANDN U5177 ( .B(n4437), .A(n4438), .Z(n4435) );
  XNOR U5178 ( .A(b[3356]), .B(n4436), .Z(n4437) );
  XNOR U5179 ( .A(b[3356]), .B(n4438), .Z(c[3356]) );
  XNOR U5180 ( .A(a[3356]), .B(n4439), .Z(n4438) );
  IV U5181 ( .A(n4436), .Z(n4439) );
  XOR U5182 ( .A(n4440), .B(n4441), .Z(n4436) );
  ANDN U5183 ( .B(n4442), .A(n4443), .Z(n4440) );
  XNOR U5184 ( .A(b[3355]), .B(n4441), .Z(n4442) );
  XNOR U5185 ( .A(b[3355]), .B(n4443), .Z(c[3355]) );
  XNOR U5186 ( .A(a[3355]), .B(n4444), .Z(n4443) );
  IV U5187 ( .A(n4441), .Z(n4444) );
  XOR U5188 ( .A(n4445), .B(n4446), .Z(n4441) );
  ANDN U5189 ( .B(n4447), .A(n4448), .Z(n4445) );
  XNOR U5190 ( .A(b[3354]), .B(n4446), .Z(n4447) );
  XNOR U5191 ( .A(b[3354]), .B(n4448), .Z(c[3354]) );
  XNOR U5192 ( .A(a[3354]), .B(n4449), .Z(n4448) );
  IV U5193 ( .A(n4446), .Z(n4449) );
  XOR U5194 ( .A(n4450), .B(n4451), .Z(n4446) );
  ANDN U5195 ( .B(n4452), .A(n4453), .Z(n4450) );
  XNOR U5196 ( .A(b[3353]), .B(n4451), .Z(n4452) );
  XNOR U5197 ( .A(b[3353]), .B(n4453), .Z(c[3353]) );
  XNOR U5198 ( .A(a[3353]), .B(n4454), .Z(n4453) );
  IV U5199 ( .A(n4451), .Z(n4454) );
  XOR U5200 ( .A(n4455), .B(n4456), .Z(n4451) );
  ANDN U5201 ( .B(n4457), .A(n4458), .Z(n4455) );
  XNOR U5202 ( .A(b[3352]), .B(n4456), .Z(n4457) );
  XNOR U5203 ( .A(b[3352]), .B(n4458), .Z(c[3352]) );
  XNOR U5204 ( .A(a[3352]), .B(n4459), .Z(n4458) );
  IV U5205 ( .A(n4456), .Z(n4459) );
  XOR U5206 ( .A(n4460), .B(n4461), .Z(n4456) );
  ANDN U5207 ( .B(n4462), .A(n4463), .Z(n4460) );
  XNOR U5208 ( .A(b[3351]), .B(n4461), .Z(n4462) );
  XNOR U5209 ( .A(b[3351]), .B(n4463), .Z(c[3351]) );
  XNOR U5210 ( .A(a[3351]), .B(n4464), .Z(n4463) );
  IV U5211 ( .A(n4461), .Z(n4464) );
  XOR U5212 ( .A(n4465), .B(n4466), .Z(n4461) );
  ANDN U5213 ( .B(n4467), .A(n4468), .Z(n4465) );
  XNOR U5214 ( .A(b[3350]), .B(n4466), .Z(n4467) );
  XNOR U5215 ( .A(b[3350]), .B(n4468), .Z(c[3350]) );
  XNOR U5216 ( .A(a[3350]), .B(n4469), .Z(n4468) );
  IV U5217 ( .A(n4466), .Z(n4469) );
  XOR U5218 ( .A(n4470), .B(n4471), .Z(n4466) );
  ANDN U5219 ( .B(n4472), .A(n4473), .Z(n4470) );
  XNOR U5220 ( .A(b[3349]), .B(n4471), .Z(n4472) );
  XNOR U5221 ( .A(b[334]), .B(n4474), .Z(c[334]) );
  XNOR U5222 ( .A(b[3349]), .B(n4473), .Z(c[3349]) );
  XNOR U5223 ( .A(a[3349]), .B(n4475), .Z(n4473) );
  IV U5224 ( .A(n4471), .Z(n4475) );
  XOR U5225 ( .A(n4476), .B(n4477), .Z(n4471) );
  ANDN U5226 ( .B(n4478), .A(n4479), .Z(n4476) );
  XNOR U5227 ( .A(b[3348]), .B(n4477), .Z(n4478) );
  XNOR U5228 ( .A(b[3348]), .B(n4479), .Z(c[3348]) );
  XNOR U5229 ( .A(a[3348]), .B(n4480), .Z(n4479) );
  IV U5230 ( .A(n4477), .Z(n4480) );
  XOR U5231 ( .A(n4481), .B(n4482), .Z(n4477) );
  ANDN U5232 ( .B(n4483), .A(n4484), .Z(n4481) );
  XNOR U5233 ( .A(b[3347]), .B(n4482), .Z(n4483) );
  XNOR U5234 ( .A(b[3347]), .B(n4484), .Z(c[3347]) );
  XNOR U5235 ( .A(a[3347]), .B(n4485), .Z(n4484) );
  IV U5236 ( .A(n4482), .Z(n4485) );
  XOR U5237 ( .A(n4486), .B(n4487), .Z(n4482) );
  ANDN U5238 ( .B(n4488), .A(n4489), .Z(n4486) );
  XNOR U5239 ( .A(b[3346]), .B(n4487), .Z(n4488) );
  XNOR U5240 ( .A(b[3346]), .B(n4489), .Z(c[3346]) );
  XNOR U5241 ( .A(a[3346]), .B(n4490), .Z(n4489) );
  IV U5242 ( .A(n4487), .Z(n4490) );
  XOR U5243 ( .A(n4491), .B(n4492), .Z(n4487) );
  ANDN U5244 ( .B(n4493), .A(n4494), .Z(n4491) );
  XNOR U5245 ( .A(b[3345]), .B(n4492), .Z(n4493) );
  XNOR U5246 ( .A(b[3345]), .B(n4494), .Z(c[3345]) );
  XNOR U5247 ( .A(a[3345]), .B(n4495), .Z(n4494) );
  IV U5248 ( .A(n4492), .Z(n4495) );
  XOR U5249 ( .A(n4496), .B(n4497), .Z(n4492) );
  ANDN U5250 ( .B(n4498), .A(n4499), .Z(n4496) );
  XNOR U5251 ( .A(b[3344]), .B(n4497), .Z(n4498) );
  XNOR U5252 ( .A(b[3344]), .B(n4499), .Z(c[3344]) );
  XNOR U5253 ( .A(a[3344]), .B(n4500), .Z(n4499) );
  IV U5254 ( .A(n4497), .Z(n4500) );
  XOR U5255 ( .A(n4501), .B(n4502), .Z(n4497) );
  ANDN U5256 ( .B(n4503), .A(n4504), .Z(n4501) );
  XNOR U5257 ( .A(b[3343]), .B(n4502), .Z(n4503) );
  XNOR U5258 ( .A(b[3343]), .B(n4504), .Z(c[3343]) );
  XNOR U5259 ( .A(a[3343]), .B(n4505), .Z(n4504) );
  IV U5260 ( .A(n4502), .Z(n4505) );
  XOR U5261 ( .A(n4506), .B(n4507), .Z(n4502) );
  ANDN U5262 ( .B(n4508), .A(n4509), .Z(n4506) );
  XNOR U5263 ( .A(b[3342]), .B(n4507), .Z(n4508) );
  XNOR U5264 ( .A(b[3342]), .B(n4509), .Z(c[3342]) );
  XNOR U5265 ( .A(a[3342]), .B(n4510), .Z(n4509) );
  IV U5266 ( .A(n4507), .Z(n4510) );
  XOR U5267 ( .A(n4511), .B(n4512), .Z(n4507) );
  ANDN U5268 ( .B(n4513), .A(n4514), .Z(n4511) );
  XNOR U5269 ( .A(b[3341]), .B(n4512), .Z(n4513) );
  XNOR U5270 ( .A(b[3341]), .B(n4514), .Z(c[3341]) );
  XNOR U5271 ( .A(a[3341]), .B(n4515), .Z(n4514) );
  IV U5272 ( .A(n4512), .Z(n4515) );
  XOR U5273 ( .A(n4516), .B(n4517), .Z(n4512) );
  ANDN U5274 ( .B(n4518), .A(n4519), .Z(n4516) );
  XNOR U5275 ( .A(b[3340]), .B(n4517), .Z(n4518) );
  XNOR U5276 ( .A(b[3340]), .B(n4519), .Z(c[3340]) );
  XNOR U5277 ( .A(a[3340]), .B(n4520), .Z(n4519) );
  IV U5278 ( .A(n4517), .Z(n4520) );
  XOR U5279 ( .A(n4521), .B(n4522), .Z(n4517) );
  ANDN U5280 ( .B(n4523), .A(n4524), .Z(n4521) );
  XNOR U5281 ( .A(b[3339]), .B(n4522), .Z(n4523) );
  XNOR U5282 ( .A(b[333]), .B(n4525), .Z(c[333]) );
  XNOR U5283 ( .A(b[3339]), .B(n4524), .Z(c[3339]) );
  XNOR U5284 ( .A(a[3339]), .B(n4526), .Z(n4524) );
  IV U5285 ( .A(n4522), .Z(n4526) );
  XOR U5286 ( .A(n4527), .B(n4528), .Z(n4522) );
  ANDN U5287 ( .B(n4529), .A(n4530), .Z(n4527) );
  XNOR U5288 ( .A(b[3338]), .B(n4528), .Z(n4529) );
  XNOR U5289 ( .A(b[3338]), .B(n4530), .Z(c[3338]) );
  XNOR U5290 ( .A(a[3338]), .B(n4531), .Z(n4530) );
  IV U5291 ( .A(n4528), .Z(n4531) );
  XOR U5292 ( .A(n4532), .B(n4533), .Z(n4528) );
  ANDN U5293 ( .B(n4534), .A(n4535), .Z(n4532) );
  XNOR U5294 ( .A(b[3337]), .B(n4533), .Z(n4534) );
  XNOR U5295 ( .A(b[3337]), .B(n4535), .Z(c[3337]) );
  XNOR U5296 ( .A(a[3337]), .B(n4536), .Z(n4535) );
  IV U5297 ( .A(n4533), .Z(n4536) );
  XOR U5298 ( .A(n4537), .B(n4538), .Z(n4533) );
  ANDN U5299 ( .B(n4539), .A(n4540), .Z(n4537) );
  XNOR U5300 ( .A(b[3336]), .B(n4538), .Z(n4539) );
  XNOR U5301 ( .A(b[3336]), .B(n4540), .Z(c[3336]) );
  XNOR U5302 ( .A(a[3336]), .B(n4541), .Z(n4540) );
  IV U5303 ( .A(n4538), .Z(n4541) );
  XOR U5304 ( .A(n4542), .B(n4543), .Z(n4538) );
  ANDN U5305 ( .B(n4544), .A(n4545), .Z(n4542) );
  XNOR U5306 ( .A(b[3335]), .B(n4543), .Z(n4544) );
  XNOR U5307 ( .A(b[3335]), .B(n4545), .Z(c[3335]) );
  XNOR U5308 ( .A(a[3335]), .B(n4546), .Z(n4545) );
  IV U5309 ( .A(n4543), .Z(n4546) );
  XOR U5310 ( .A(n4547), .B(n4548), .Z(n4543) );
  ANDN U5311 ( .B(n4549), .A(n4550), .Z(n4547) );
  XNOR U5312 ( .A(b[3334]), .B(n4548), .Z(n4549) );
  XNOR U5313 ( .A(b[3334]), .B(n4550), .Z(c[3334]) );
  XNOR U5314 ( .A(a[3334]), .B(n4551), .Z(n4550) );
  IV U5315 ( .A(n4548), .Z(n4551) );
  XOR U5316 ( .A(n4552), .B(n4553), .Z(n4548) );
  ANDN U5317 ( .B(n4554), .A(n4555), .Z(n4552) );
  XNOR U5318 ( .A(b[3333]), .B(n4553), .Z(n4554) );
  XNOR U5319 ( .A(b[3333]), .B(n4555), .Z(c[3333]) );
  XNOR U5320 ( .A(a[3333]), .B(n4556), .Z(n4555) );
  IV U5321 ( .A(n4553), .Z(n4556) );
  XOR U5322 ( .A(n4557), .B(n4558), .Z(n4553) );
  ANDN U5323 ( .B(n4559), .A(n4560), .Z(n4557) );
  XNOR U5324 ( .A(b[3332]), .B(n4558), .Z(n4559) );
  XNOR U5325 ( .A(b[3332]), .B(n4560), .Z(c[3332]) );
  XNOR U5326 ( .A(a[3332]), .B(n4561), .Z(n4560) );
  IV U5327 ( .A(n4558), .Z(n4561) );
  XOR U5328 ( .A(n4562), .B(n4563), .Z(n4558) );
  ANDN U5329 ( .B(n4564), .A(n4565), .Z(n4562) );
  XNOR U5330 ( .A(b[3331]), .B(n4563), .Z(n4564) );
  XNOR U5331 ( .A(b[3331]), .B(n4565), .Z(c[3331]) );
  XNOR U5332 ( .A(a[3331]), .B(n4566), .Z(n4565) );
  IV U5333 ( .A(n4563), .Z(n4566) );
  XOR U5334 ( .A(n4567), .B(n4568), .Z(n4563) );
  ANDN U5335 ( .B(n4569), .A(n4570), .Z(n4567) );
  XNOR U5336 ( .A(b[3330]), .B(n4568), .Z(n4569) );
  XNOR U5337 ( .A(b[3330]), .B(n4570), .Z(c[3330]) );
  XNOR U5338 ( .A(a[3330]), .B(n4571), .Z(n4570) );
  IV U5339 ( .A(n4568), .Z(n4571) );
  XOR U5340 ( .A(n4572), .B(n4573), .Z(n4568) );
  ANDN U5341 ( .B(n4574), .A(n4575), .Z(n4572) );
  XNOR U5342 ( .A(b[3329]), .B(n4573), .Z(n4574) );
  XNOR U5343 ( .A(b[332]), .B(n4576), .Z(c[332]) );
  XNOR U5344 ( .A(b[3329]), .B(n4575), .Z(c[3329]) );
  XNOR U5345 ( .A(a[3329]), .B(n4577), .Z(n4575) );
  IV U5346 ( .A(n4573), .Z(n4577) );
  XOR U5347 ( .A(n4578), .B(n4579), .Z(n4573) );
  ANDN U5348 ( .B(n4580), .A(n4581), .Z(n4578) );
  XNOR U5349 ( .A(b[3328]), .B(n4579), .Z(n4580) );
  XNOR U5350 ( .A(b[3328]), .B(n4581), .Z(c[3328]) );
  XNOR U5351 ( .A(a[3328]), .B(n4582), .Z(n4581) );
  IV U5352 ( .A(n4579), .Z(n4582) );
  XOR U5353 ( .A(n4583), .B(n4584), .Z(n4579) );
  ANDN U5354 ( .B(n4585), .A(n4586), .Z(n4583) );
  XNOR U5355 ( .A(b[3327]), .B(n4584), .Z(n4585) );
  XNOR U5356 ( .A(b[3327]), .B(n4586), .Z(c[3327]) );
  XNOR U5357 ( .A(a[3327]), .B(n4587), .Z(n4586) );
  IV U5358 ( .A(n4584), .Z(n4587) );
  XOR U5359 ( .A(n4588), .B(n4589), .Z(n4584) );
  ANDN U5360 ( .B(n4590), .A(n4591), .Z(n4588) );
  XNOR U5361 ( .A(b[3326]), .B(n4589), .Z(n4590) );
  XNOR U5362 ( .A(b[3326]), .B(n4591), .Z(c[3326]) );
  XNOR U5363 ( .A(a[3326]), .B(n4592), .Z(n4591) );
  IV U5364 ( .A(n4589), .Z(n4592) );
  XOR U5365 ( .A(n4593), .B(n4594), .Z(n4589) );
  ANDN U5366 ( .B(n4595), .A(n4596), .Z(n4593) );
  XNOR U5367 ( .A(b[3325]), .B(n4594), .Z(n4595) );
  XNOR U5368 ( .A(b[3325]), .B(n4596), .Z(c[3325]) );
  XNOR U5369 ( .A(a[3325]), .B(n4597), .Z(n4596) );
  IV U5370 ( .A(n4594), .Z(n4597) );
  XOR U5371 ( .A(n4598), .B(n4599), .Z(n4594) );
  ANDN U5372 ( .B(n4600), .A(n4601), .Z(n4598) );
  XNOR U5373 ( .A(b[3324]), .B(n4599), .Z(n4600) );
  XNOR U5374 ( .A(b[3324]), .B(n4601), .Z(c[3324]) );
  XNOR U5375 ( .A(a[3324]), .B(n4602), .Z(n4601) );
  IV U5376 ( .A(n4599), .Z(n4602) );
  XOR U5377 ( .A(n4603), .B(n4604), .Z(n4599) );
  ANDN U5378 ( .B(n4605), .A(n4606), .Z(n4603) );
  XNOR U5379 ( .A(b[3323]), .B(n4604), .Z(n4605) );
  XNOR U5380 ( .A(b[3323]), .B(n4606), .Z(c[3323]) );
  XNOR U5381 ( .A(a[3323]), .B(n4607), .Z(n4606) );
  IV U5382 ( .A(n4604), .Z(n4607) );
  XOR U5383 ( .A(n4608), .B(n4609), .Z(n4604) );
  ANDN U5384 ( .B(n4610), .A(n4611), .Z(n4608) );
  XNOR U5385 ( .A(b[3322]), .B(n4609), .Z(n4610) );
  XNOR U5386 ( .A(b[3322]), .B(n4611), .Z(c[3322]) );
  XNOR U5387 ( .A(a[3322]), .B(n4612), .Z(n4611) );
  IV U5388 ( .A(n4609), .Z(n4612) );
  XOR U5389 ( .A(n4613), .B(n4614), .Z(n4609) );
  ANDN U5390 ( .B(n4615), .A(n4616), .Z(n4613) );
  XNOR U5391 ( .A(b[3321]), .B(n4614), .Z(n4615) );
  XNOR U5392 ( .A(b[3321]), .B(n4616), .Z(c[3321]) );
  XNOR U5393 ( .A(a[3321]), .B(n4617), .Z(n4616) );
  IV U5394 ( .A(n4614), .Z(n4617) );
  XOR U5395 ( .A(n4618), .B(n4619), .Z(n4614) );
  ANDN U5396 ( .B(n4620), .A(n4621), .Z(n4618) );
  XNOR U5397 ( .A(b[3320]), .B(n4619), .Z(n4620) );
  XNOR U5398 ( .A(b[3320]), .B(n4621), .Z(c[3320]) );
  XNOR U5399 ( .A(a[3320]), .B(n4622), .Z(n4621) );
  IV U5400 ( .A(n4619), .Z(n4622) );
  XOR U5401 ( .A(n4623), .B(n4624), .Z(n4619) );
  ANDN U5402 ( .B(n4625), .A(n4626), .Z(n4623) );
  XNOR U5403 ( .A(b[3319]), .B(n4624), .Z(n4625) );
  XNOR U5404 ( .A(b[331]), .B(n4627), .Z(c[331]) );
  XNOR U5405 ( .A(b[3319]), .B(n4626), .Z(c[3319]) );
  XNOR U5406 ( .A(a[3319]), .B(n4628), .Z(n4626) );
  IV U5407 ( .A(n4624), .Z(n4628) );
  XOR U5408 ( .A(n4629), .B(n4630), .Z(n4624) );
  ANDN U5409 ( .B(n4631), .A(n4632), .Z(n4629) );
  XNOR U5410 ( .A(b[3318]), .B(n4630), .Z(n4631) );
  XNOR U5411 ( .A(b[3318]), .B(n4632), .Z(c[3318]) );
  XNOR U5412 ( .A(a[3318]), .B(n4633), .Z(n4632) );
  IV U5413 ( .A(n4630), .Z(n4633) );
  XOR U5414 ( .A(n4634), .B(n4635), .Z(n4630) );
  ANDN U5415 ( .B(n4636), .A(n4637), .Z(n4634) );
  XNOR U5416 ( .A(b[3317]), .B(n4635), .Z(n4636) );
  XNOR U5417 ( .A(b[3317]), .B(n4637), .Z(c[3317]) );
  XNOR U5418 ( .A(a[3317]), .B(n4638), .Z(n4637) );
  IV U5419 ( .A(n4635), .Z(n4638) );
  XOR U5420 ( .A(n4639), .B(n4640), .Z(n4635) );
  ANDN U5421 ( .B(n4641), .A(n4642), .Z(n4639) );
  XNOR U5422 ( .A(b[3316]), .B(n4640), .Z(n4641) );
  XNOR U5423 ( .A(b[3316]), .B(n4642), .Z(c[3316]) );
  XNOR U5424 ( .A(a[3316]), .B(n4643), .Z(n4642) );
  IV U5425 ( .A(n4640), .Z(n4643) );
  XOR U5426 ( .A(n4644), .B(n4645), .Z(n4640) );
  ANDN U5427 ( .B(n4646), .A(n4647), .Z(n4644) );
  XNOR U5428 ( .A(b[3315]), .B(n4645), .Z(n4646) );
  XNOR U5429 ( .A(b[3315]), .B(n4647), .Z(c[3315]) );
  XNOR U5430 ( .A(a[3315]), .B(n4648), .Z(n4647) );
  IV U5431 ( .A(n4645), .Z(n4648) );
  XOR U5432 ( .A(n4649), .B(n4650), .Z(n4645) );
  ANDN U5433 ( .B(n4651), .A(n4652), .Z(n4649) );
  XNOR U5434 ( .A(b[3314]), .B(n4650), .Z(n4651) );
  XNOR U5435 ( .A(b[3314]), .B(n4652), .Z(c[3314]) );
  XNOR U5436 ( .A(a[3314]), .B(n4653), .Z(n4652) );
  IV U5437 ( .A(n4650), .Z(n4653) );
  XOR U5438 ( .A(n4654), .B(n4655), .Z(n4650) );
  ANDN U5439 ( .B(n4656), .A(n4657), .Z(n4654) );
  XNOR U5440 ( .A(b[3313]), .B(n4655), .Z(n4656) );
  XNOR U5441 ( .A(b[3313]), .B(n4657), .Z(c[3313]) );
  XNOR U5442 ( .A(a[3313]), .B(n4658), .Z(n4657) );
  IV U5443 ( .A(n4655), .Z(n4658) );
  XOR U5444 ( .A(n4659), .B(n4660), .Z(n4655) );
  ANDN U5445 ( .B(n4661), .A(n4662), .Z(n4659) );
  XNOR U5446 ( .A(b[3312]), .B(n4660), .Z(n4661) );
  XNOR U5447 ( .A(b[3312]), .B(n4662), .Z(c[3312]) );
  XNOR U5448 ( .A(a[3312]), .B(n4663), .Z(n4662) );
  IV U5449 ( .A(n4660), .Z(n4663) );
  XOR U5450 ( .A(n4664), .B(n4665), .Z(n4660) );
  ANDN U5451 ( .B(n4666), .A(n4667), .Z(n4664) );
  XNOR U5452 ( .A(b[3311]), .B(n4665), .Z(n4666) );
  XNOR U5453 ( .A(b[3311]), .B(n4667), .Z(c[3311]) );
  XNOR U5454 ( .A(a[3311]), .B(n4668), .Z(n4667) );
  IV U5455 ( .A(n4665), .Z(n4668) );
  XOR U5456 ( .A(n4669), .B(n4670), .Z(n4665) );
  ANDN U5457 ( .B(n4671), .A(n4672), .Z(n4669) );
  XNOR U5458 ( .A(b[3310]), .B(n4670), .Z(n4671) );
  XNOR U5459 ( .A(b[3310]), .B(n4672), .Z(c[3310]) );
  XNOR U5460 ( .A(a[3310]), .B(n4673), .Z(n4672) );
  IV U5461 ( .A(n4670), .Z(n4673) );
  XOR U5462 ( .A(n4674), .B(n4675), .Z(n4670) );
  ANDN U5463 ( .B(n4676), .A(n4677), .Z(n4674) );
  XNOR U5464 ( .A(b[3309]), .B(n4675), .Z(n4676) );
  XNOR U5465 ( .A(b[330]), .B(n4678), .Z(c[330]) );
  XNOR U5466 ( .A(b[3309]), .B(n4677), .Z(c[3309]) );
  XNOR U5467 ( .A(a[3309]), .B(n4679), .Z(n4677) );
  IV U5468 ( .A(n4675), .Z(n4679) );
  XOR U5469 ( .A(n4680), .B(n4681), .Z(n4675) );
  ANDN U5470 ( .B(n4682), .A(n4683), .Z(n4680) );
  XNOR U5471 ( .A(b[3308]), .B(n4681), .Z(n4682) );
  XNOR U5472 ( .A(b[3308]), .B(n4683), .Z(c[3308]) );
  XNOR U5473 ( .A(a[3308]), .B(n4684), .Z(n4683) );
  IV U5474 ( .A(n4681), .Z(n4684) );
  XOR U5475 ( .A(n4685), .B(n4686), .Z(n4681) );
  ANDN U5476 ( .B(n4687), .A(n4688), .Z(n4685) );
  XNOR U5477 ( .A(b[3307]), .B(n4686), .Z(n4687) );
  XNOR U5478 ( .A(b[3307]), .B(n4688), .Z(c[3307]) );
  XNOR U5479 ( .A(a[3307]), .B(n4689), .Z(n4688) );
  IV U5480 ( .A(n4686), .Z(n4689) );
  XOR U5481 ( .A(n4690), .B(n4691), .Z(n4686) );
  ANDN U5482 ( .B(n4692), .A(n4693), .Z(n4690) );
  XNOR U5483 ( .A(b[3306]), .B(n4691), .Z(n4692) );
  XNOR U5484 ( .A(b[3306]), .B(n4693), .Z(c[3306]) );
  XNOR U5485 ( .A(a[3306]), .B(n4694), .Z(n4693) );
  IV U5486 ( .A(n4691), .Z(n4694) );
  XOR U5487 ( .A(n4695), .B(n4696), .Z(n4691) );
  ANDN U5488 ( .B(n4697), .A(n4698), .Z(n4695) );
  XNOR U5489 ( .A(b[3305]), .B(n4696), .Z(n4697) );
  XNOR U5490 ( .A(b[3305]), .B(n4698), .Z(c[3305]) );
  XNOR U5491 ( .A(a[3305]), .B(n4699), .Z(n4698) );
  IV U5492 ( .A(n4696), .Z(n4699) );
  XOR U5493 ( .A(n4700), .B(n4701), .Z(n4696) );
  ANDN U5494 ( .B(n4702), .A(n4703), .Z(n4700) );
  XNOR U5495 ( .A(b[3304]), .B(n4701), .Z(n4702) );
  XNOR U5496 ( .A(b[3304]), .B(n4703), .Z(c[3304]) );
  XNOR U5497 ( .A(a[3304]), .B(n4704), .Z(n4703) );
  IV U5498 ( .A(n4701), .Z(n4704) );
  XOR U5499 ( .A(n4705), .B(n4706), .Z(n4701) );
  ANDN U5500 ( .B(n4707), .A(n4708), .Z(n4705) );
  XNOR U5501 ( .A(b[3303]), .B(n4706), .Z(n4707) );
  XNOR U5502 ( .A(b[3303]), .B(n4708), .Z(c[3303]) );
  XNOR U5503 ( .A(a[3303]), .B(n4709), .Z(n4708) );
  IV U5504 ( .A(n4706), .Z(n4709) );
  XOR U5505 ( .A(n4710), .B(n4711), .Z(n4706) );
  ANDN U5506 ( .B(n4712), .A(n4713), .Z(n4710) );
  XNOR U5507 ( .A(b[3302]), .B(n4711), .Z(n4712) );
  XNOR U5508 ( .A(b[3302]), .B(n4713), .Z(c[3302]) );
  XNOR U5509 ( .A(a[3302]), .B(n4714), .Z(n4713) );
  IV U5510 ( .A(n4711), .Z(n4714) );
  XOR U5511 ( .A(n4715), .B(n4716), .Z(n4711) );
  ANDN U5512 ( .B(n4717), .A(n4718), .Z(n4715) );
  XNOR U5513 ( .A(b[3301]), .B(n4716), .Z(n4717) );
  XNOR U5514 ( .A(b[3301]), .B(n4718), .Z(c[3301]) );
  XNOR U5515 ( .A(a[3301]), .B(n4719), .Z(n4718) );
  IV U5516 ( .A(n4716), .Z(n4719) );
  XOR U5517 ( .A(n4720), .B(n4721), .Z(n4716) );
  ANDN U5518 ( .B(n4722), .A(n4723), .Z(n4720) );
  XNOR U5519 ( .A(b[3300]), .B(n4721), .Z(n4722) );
  XNOR U5520 ( .A(b[3300]), .B(n4723), .Z(c[3300]) );
  XNOR U5521 ( .A(a[3300]), .B(n4724), .Z(n4723) );
  IV U5522 ( .A(n4721), .Z(n4724) );
  XOR U5523 ( .A(n4725), .B(n4726), .Z(n4721) );
  ANDN U5524 ( .B(n4727), .A(n4728), .Z(n4725) );
  XNOR U5525 ( .A(b[3299]), .B(n4726), .Z(n4727) );
  XNOR U5526 ( .A(b[32]), .B(n4729), .Z(c[32]) );
  XNOR U5527 ( .A(b[329]), .B(n4730), .Z(c[329]) );
  XNOR U5528 ( .A(b[3299]), .B(n4728), .Z(c[3299]) );
  XNOR U5529 ( .A(a[3299]), .B(n4731), .Z(n4728) );
  IV U5530 ( .A(n4726), .Z(n4731) );
  XOR U5531 ( .A(n4732), .B(n4733), .Z(n4726) );
  ANDN U5532 ( .B(n4734), .A(n4735), .Z(n4732) );
  XNOR U5533 ( .A(b[3298]), .B(n4733), .Z(n4734) );
  XNOR U5534 ( .A(b[3298]), .B(n4735), .Z(c[3298]) );
  XNOR U5535 ( .A(a[3298]), .B(n4736), .Z(n4735) );
  IV U5536 ( .A(n4733), .Z(n4736) );
  XOR U5537 ( .A(n4737), .B(n4738), .Z(n4733) );
  ANDN U5538 ( .B(n4739), .A(n4740), .Z(n4737) );
  XNOR U5539 ( .A(b[3297]), .B(n4738), .Z(n4739) );
  XNOR U5540 ( .A(b[3297]), .B(n4740), .Z(c[3297]) );
  XNOR U5541 ( .A(a[3297]), .B(n4741), .Z(n4740) );
  IV U5542 ( .A(n4738), .Z(n4741) );
  XOR U5543 ( .A(n4742), .B(n4743), .Z(n4738) );
  ANDN U5544 ( .B(n4744), .A(n4745), .Z(n4742) );
  XNOR U5545 ( .A(b[3296]), .B(n4743), .Z(n4744) );
  XNOR U5546 ( .A(b[3296]), .B(n4745), .Z(c[3296]) );
  XNOR U5547 ( .A(a[3296]), .B(n4746), .Z(n4745) );
  IV U5548 ( .A(n4743), .Z(n4746) );
  XOR U5549 ( .A(n4747), .B(n4748), .Z(n4743) );
  ANDN U5550 ( .B(n4749), .A(n4750), .Z(n4747) );
  XNOR U5551 ( .A(b[3295]), .B(n4748), .Z(n4749) );
  XNOR U5552 ( .A(b[3295]), .B(n4750), .Z(c[3295]) );
  XNOR U5553 ( .A(a[3295]), .B(n4751), .Z(n4750) );
  IV U5554 ( .A(n4748), .Z(n4751) );
  XOR U5555 ( .A(n4752), .B(n4753), .Z(n4748) );
  ANDN U5556 ( .B(n4754), .A(n4755), .Z(n4752) );
  XNOR U5557 ( .A(b[3294]), .B(n4753), .Z(n4754) );
  XNOR U5558 ( .A(b[3294]), .B(n4755), .Z(c[3294]) );
  XNOR U5559 ( .A(a[3294]), .B(n4756), .Z(n4755) );
  IV U5560 ( .A(n4753), .Z(n4756) );
  XOR U5561 ( .A(n4757), .B(n4758), .Z(n4753) );
  ANDN U5562 ( .B(n4759), .A(n4760), .Z(n4757) );
  XNOR U5563 ( .A(b[3293]), .B(n4758), .Z(n4759) );
  XNOR U5564 ( .A(b[3293]), .B(n4760), .Z(c[3293]) );
  XNOR U5565 ( .A(a[3293]), .B(n4761), .Z(n4760) );
  IV U5566 ( .A(n4758), .Z(n4761) );
  XOR U5567 ( .A(n4762), .B(n4763), .Z(n4758) );
  ANDN U5568 ( .B(n4764), .A(n4765), .Z(n4762) );
  XNOR U5569 ( .A(b[3292]), .B(n4763), .Z(n4764) );
  XNOR U5570 ( .A(b[3292]), .B(n4765), .Z(c[3292]) );
  XNOR U5571 ( .A(a[3292]), .B(n4766), .Z(n4765) );
  IV U5572 ( .A(n4763), .Z(n4766) );
  XOR U5573 ( .A(n4767), .B(n4768), .Z(n4763) );
  ANDN U5574 ( .B(n4769), .A(n4770), .Z(n4767) );
  XNOR U5575 ( .A(b[3291]), .B(n4768), .Z(n4769) );
  XNOR U5576 ( .A(b[3291]), .B(n4770), .Z(c[3291]) );
  XNOR U5577 ( .A(a[3291]), .B(n4771), .Z(n4770) );
  IV U5578 ( .A(n4768), .Z(n4771) );
  XOR U5579 ( .A(n4772), .B(n4773), .Z(n4768) );
  ANDN U5580 ( .B(n4774), .A(n4775), .Z(n4772) );
  XNOR U5581 ( .A(b[3290]), .B(n4773), .Z(n4774) );
  XNOR U5582 ( .A(b[3290]), .B(n4775), .Z(c[3290]) );
  XNOR U5583 ( .A(a[3290]), .B(n4776), .Z(n4775) );
  IV U5584 ( .A(n4773), .Z(n4776) );
  XOR U5585 ( .A(n4777), .B(n4778), .Z(n4773) );
  ANDN U5586 ( .B(n4779), .A(n4780), .Z(n4777) );
  XNOR U5587 ( .A(b[3289]), .B(n4778), .Z(n4779) );
  XNOR U5588 ( .A(b[328]), .B(n4781), .Z(c[328]) );
  XNOR U5589 ( .A(b[3289]), .B(n4780), .Z(c[3289]) );
  XNOR U5590 ( .A(a[3289]), .B(n4782), .Z(n4780) );
  IV U5591 ( .A(n4778), .Z(n4782) );
  XOR U5592 ( .A(n4783), .B(n4784), .Z(n4778) );
  ANDN U5593 ( .B(n4785), .A(n4786), .Z(n4783) );
  XNOR U5594 ( .A(b[3288]), .B(n4784), .Z(n4785) );
  XNOR U5595 ( .A(b[3288]), .B(n4786), .Z(c[3288]) );
  XNOR U5596 ( .A(a[3288]), .B(n4787), .Z(n4786) );
  IV U5597 ( .A(n4784), .Z(n4787) );
  XOR U5598 ( .A(n4788), .B(n4789), .Z(n4784) );
  ANDN U5599 ( .B(n4790), .A(n4791), .Z(n4788) );
  XNOR U5600 ( .A(b[3287]), .B(n4789), .Z(n4790) );
  XNOR U5601 ( .A(b[3287]), .B(n4791), .Z(c[3287]) );
  XNOR U5602 ( .A(a[3287]), .B(n4792), .Z(n4791) );
  IV U5603 ( .A(n4789), .Z(n4792) );
  XOR U5604 ( .A(n4793), .B(n4794), .Z(n4789) );
  ANDN U5605 ( .B(n4795), .A(n4796), .Z(n4793) );
  XNOR U5606 ( .A(b[3286]), .B(n4794), .Z(n4795) );
  XNOR U5607 ( .A(b[3286]), .B(n4796), .Z(c[3286]) );
  XNOR U5608 ( .A(a[3286]), .B(n4797), .Z(n4796) );
  IV U5609 ( .A(n4794), .Z(n4797) );
  XOR U5610 ( .A(n4798), .B(n4799), .Z(n4794) );
  ANDN U5611 ( .B(n4800), .A(n4801), .Z(n4798) );
  XNOR U5612 ( .A(b[3285]), .B(n4799), .Z(n4800) );
  XNOR U5613 ( .A(b[3285]), .B(n4801), .Z(c[3285]) );
  XNOR U5614 ( .A(a[3285]), .B(n4802), .Z(n4801) );
  IV U5615 ( .A(n4799), .Z(n4802) );
  XOR U5616 ( .A(n4803), .B(n4804), .Z(n4799) );
  ANDN U5617 ( .B(n4805), .A(n4806), .Z(n4803) );
  XNOR U5618 ( .A(b[3284]), .B(n4804), .Z(n4805) );
  XNOR U5619 ( .A(b[3284]), .B(n4806), .Z(c[3284]) );
  XNOR U5620 ( .A(a[3284]), .B(n4807), .Z(n4806) );
  IV U5621 ( .A(n4804), .Z(n4807) );
  XOR U5622 ( .A(n4808), .B(n4809), .Z(n4804) );
  ANDN U5623 ( .B(n4810), .A(n4811), .Z(n4808) );
  XNOR U5624 ( .A(b[3283]), .B(n4809), .Z(n4810) );
  XNOR U5625 ( .A(b[3283]), .B(n4811), .Z(c[3283]) );
  XNOR U5626 ( .A(a[3283]), .B(n4812), .Z(n4811) );
  IV U5627 ( .A(n4809), .Z(n4812) );
  XOR U5628 ( .A(n4813), .B(n4814), .Z(n4809) );
  ANDN U5629 ( .B(n4815), .A(n4816), .Z(n4813) );
  XNOR U5630 ( .A(b[3282]), .B(n4814), .Z(n4815) );
  XNOR U5631 ( .A(b[3282]), .B(n4816), .Z(c[3282]) );
  XNOR U5632 ( .A(a[3282]), .B(n4817), .Z(n4816) );
  IV U5633 ( .A(n4814), .Z(n4817) );
  XOR U5634 ( .A(n4818), .B(n4819), .Z(n4814) );
  ANDN U5635 ( .B(n4820), .A(n4821), .Z(n4818) );
  XNOR U5636 ( .A(b[3281]), .B(n4819), .Z(n4820) );
  XNOR U5637 ( .A(b[3281]), .B(n4821), .Z(c[3281]) );
  XNOR U5638 ( .A(a[3281]), .B(n4822), .Z(n4821) );
  IV U5639 ( .A(n4819), .Z(n4822) );
  XOR U5640 ( .A(n4823), .B(n4824), .Z(n4819) );
  ANDN U5641 ( .B(n4825), .A(n4826), .Z(n4823) );
  XNOR U5642 ( .A(b[3280]), .B(n4824), .Z(n4825) );
  XNOR U5643 ( .A(b[3280]), .B(n4826), .Z(c[3280]) );
  XNOR U5644 ( .A(a[3280]), .B(n4827), .Z(n4826) );
  IV U5645 ( .A(n4824), .Z(n4827) );
  XOR U5646 ( .A(n4828), .B(n4829), .Z(n4824) );
  ANDN U5647 ( .B(n4830), .A(n4831), .Z(n4828) );
  XNOR U5648 ( .A(b[3279]), .B(n4829), .Z(n4830) );
  XNOR U5649 ( .A(b[327]), .B(n4832), .Z(c[327]) );
  XNOR U5650 ( .A(b[3279]), .B(n4831), .Z(c[3279]) );
  XNOR U5651 ( .A(a[3279]), .B(n4833), .Z(n4831) );
  IV U5652 ( .A(n4829), .Z(n4833) );
  XOR U5653 ( .A(n4834), .B(n4835), .Z(n4829) );
  ANDN U5654 ( .B(n4836), .A(n4837), .Z(n4834) );
  XNOR U5655 ( .A(b[3278]), .B(n4835), .Z(n4836) );
  XNOR U5656 ( .A(b[3278]), .B(n4837), .Z(c[3278]) );
  XNOR U5657 ( .A(a[3278]), .B(n4838), .Z(n4837) );
  IV U5658 ( .A(n4835), .Z(n4838) );
  XOR U5659 ( .A(n4839), .B(n4840), .Z(n4835) );
  ANDN U5660 ( .B(n4841), .A(n4842), .Z(n4839) );
  XNOR U5661 ( .A(b[3277]), .B(n4840), .Z(n4841) );
  XNOR U5662 ( .A(b[3277]), .B(n4842), .Z(c[3277]) );
  XNOR U5663 ( .A(a[3277]), .B(n4843), .Z(n4842) );
  IV U5664 ( .A(n4840), .Z(n4843) );
  XOR U5665 ( .A(n4844), .B(n4845), .Z(n4840) );
  ANDN U5666 ( .B(n4846), .A(n4847), .Z(n4844) );
  XNOR U5667 ( .A(b[3276]), .B(n4845), .Z(n4846) );
  XNOR U5668 ( .A(b[3276]), .B(n4847), .Z(c[3276]) );
  XNOR U5669 ( .A(a[3276]), .B(n4848), .Z(n4847) );
  IV U5670 ( .A(n4845), .Z(n4848) );
  XOR U5671 ( .A(n4849), .B(n4850), .Z(n4845) );
  ANDN U5672 ( .B(n4851), .A(n4852), .Z(n4849) );
  XNOR U5673 ( .A(b[3275]), .B(n4850), .Z(n4851) );
  XNOR U5674 ( .A(b[3275]), .B(n4852), .Z(c[3275]) );
  XNOR U5675 ( .A(a[3275]), .B(n4853), .Z(n4852) );
  IV U5676 ( .A(n4850), .Z(n4853) );
  XOR U5677 ( .A(n4854), .B(n4855), .Z(n4850) );
  ANDN U5678 ( .B(n4856), .A(n4857), .Z(n4854) );
  XNOR U5679 ( .A(b[3274]), .B(n4855), .Z(n4856) );
  XNOR U5680 ( .A(b[3274]), .B(n4857), .Z(c[3274]) );
  XNOR U5681 ( .A(a[3274]), .B(n4858), .Z(n4857) );
  IV U5682 ( .A(n4855), .Z(n4858) );
  XOR U5683 ( .A(n4859), .B(n4860), .Z(n4855) );
  ANDN U5684 ( .B(n4861), .A(n4862), .Z(n4859) );
  XNOR U5685 ( .A(b[3273]), .B(n4860), .Z(n4861) );
  XNOR U5686 ( .A(b[3273]), .B(n4862), .Z(c[3273]) );
  XNOR U5687 ( .A(a[3273]), .B(n4863), .Z(n4862) );
  IV U5688 ( .A(n4860), .Z(n4863) );
  XOR U5689 ( .A(n4864), .B(n4865), .Z(n4860) );
  ANDN U5690 ( .B(n4866), .A(n4867), .Z(n4864) );
  XNOR U5691 ( .A(b[3272]), .B(n4865), .Z(n4866) );
  XNOR U5692 ( .A(b[3272]), .B(n4867), .Z(c[3272]) );
  XNOR U5693 ( .A(a[3272]), .B(n4868), .Z(n4867) );
  IV U5694 ( .A(n4865), .Z(n4868) );
  XOR U5695 ( .A(n4869), .B(n4870), .Z(n4865) );
  ANDN U5696 ( .B(n4871), .A(n4872), .Z(n4869) );
  XNOR U5697 ( .A(b[3271]), .B(n4870), .Z(n4871) );
  XNOR U5698 ( .A(b[3271]), .B(n4872), .Z(c[3271]) );
  XNOR U5699 ( .A(a[3271]), .B(n4873), .Z(n4872) );
  IV U5700 ( .A(n4870), .Z(n4873) );
  XOR U5701 ( .A(n4874), .B(n4875), .Z(n4870) );
  ANDN U5702 ( .B(n4876), .A(n4877), .Z(n4874) );
  XNOR U5703 ( .A(b[3270]), .B(n4875), .Z(n4876) );
  XNOR U5704 ( .A(b[3270]), .B(n4877), .Z(c[3270]) );
  XNOR U5705 ( .A(a[3270]), .B(n4878), .Z(n4877) );
  IV U5706 ( .A(n4875), .Z(n4878) );
  XOR U5707 ( .A(n4879), .B(n4880), .Z(n4875) );
  ANDN U5708 ( .B(n4881), .A(n4882), .Z(n4879) );
  XNOR U5709 ( .A(b[3269]), .B(n4880), .Z(n4881) );
  XNOR U5710 ( .A(b[326]), .B(n4883), .Z(c[326]) );
  XNOR U5711 ( .A(b[3269]), .B(n4882), .Z(c[3269]) );
  XNOR U5712 ( .A(a[3269]), .B(n4884), .Z(n4882) );
  IV U5713 ( .A(n4880), .Z(n4884) );
  XOR U5714 ( .A(n4885), .B(n4886), .Z(n4880) );
  ANDN U5715 ( .B(n4887), .A(n4888), .Z(n4885) );
  XNOR U5716 ( .A(b[3268]), .B(n4886), .Z(n4887) );
  XNOR U5717 ( .A(b[3268]), .B(n4888), .Z(c[3268]) );
  XNOR U5718 ( .A(a[3268]), .B(n4889), .Z(n4888) );
  IV U5719 ( .A(n4886), .Z(n4889) );
  XOR U5720 ( .A(n4890), .B(n4891), .Z(n4886) );
  ANDN U5721 ( .B(n4892), .A(n4893), .Z(n4890) );
  XNOR U5722 ( .A(b[3267]), .B(n4891), .Z(n4892) );
  XNOR U5723 ( .A(b[3267]), .B(n4893), .Z(c[3267]) );
  XNOR U5724 ( .A(a[3267]), .B(n4894), .Z(n4893) );
  IV U5725 ( .A(n4891), .Z(n4894) );
  XOR U5726 ( .A(n4895), .B(n4896), .Z(n4891) );
  ANDN U5727 ( .B(n4897), .A(n4898), .Z(n4895) );
  XNOR U5728 ( .A(b[3266]), .B(n4896), .Z(n4897) );
  XNOR U5729 ( .A(b[3266]), .B(n4898), .Z(c[3266]) );
  XNOR U5730 ( .A(a[3266]), .B(n4899), .Z(n4898) );
  IV U5731 ( .A(n4896), .Z(n4899) );
  XOR U5732 ( .A(n4900), .B(n4901), .Z(n4896) );
  ANDN U5733 ( .B(n4902), .A(n4903), .Z(n4900) );
  XNOR U5734 ( .A(b[3265]), .B(n4901), .Z(n4902) );
  XNOR U5735 ( .A(b[3265]), .B(n4903), .Z(c[3265]) );
  XNOR U5736 ( .A(a[3265]), .B(n4904), .Z(n4903) );
  IV U5737 ( .A(n4901), .Z(n4904) );
  XOR U5738 ( .A(n4905), .B(n4906), .Z(n4901) );
  ANDN U5739 ( .B(n4907), .A(n4908), .Z(n4905) );
  XNOR U5740 ( .A(b[3264]), .B(n4906), .Z(n4907) );
  XNOR U5741 ( .A(b[3264]), .B(n4908), .Z(c[3264]) );
  XNOR U5742 ( .A(a[3264]), .B(n4909), .Z(n4908) );
  IV U5743 ( .A(n4906), .Z(n4909) );
  XOR U5744 ( .A(n4910), .B(n4911), .Z(n4906) );
  ANDN U5745 ( .B(n4912), .A(n4913), .Z(n4910) );
  XNOR U5746 ( .A(b[3263]), .B(n4911), .Z(n4912) );
  XNOR U5747 ( .A(b[3263]), .B(n4913), .Z(c[3263]) );
  XNOR U5748 ( .A(a[3263]), .B(n4914), .Z(n4913) );
  IV U5749 ( .A(n4911), .Z(n4914) );
  XOR U5750 ( .A(n4915), .B(n4916), .Z(n4911) );
  ANDN U5751 ( .B(n4917), .A(n4918), .Z(n4915) );
  XNOR U5752 ( .A(b[3262]), .B(n4916), .Z(n4917) );
  XNOR U5753 ( .A(b[3262]), .B(n4918), .Z(c[3262]) );
  XNOR U5754 ( .A(a[3262]), .B(n4919), .Z(n4918) );
  IV U5755 ( .A(n4916), .Z(n4919) );
  XOR U5756 ( .A(n4920), .B(n4921), .Z(n4916) );
  ANDN U5757 ( .B(n4922), .A(n4923), .Z(n4920) );
  XNOR U5758 ( .A(b[3261]), .B(n4921), .Z(n4922) );
  XNOR U5759 ( .A(b[3261]), .B(n4923), .Z(c[3261]) );
  XNOR U5760 ( .A(a[3261]), .B(n4924), .Z(n4923) );
  IV U5761 ( .A(n4921), .Z(n4924) );
  XOR U5762 ( .A(n4925), .B(n4926), .Z(n4921) );
  ANDN U5763 ( .B(n4927), .A(n4928), .Z(n4925) );
  XNOR U5764 ( .A(b[3260]), .B(n4926), .Z(n4927) );
  XNOR U5765 ( .A(b[3260]), .B(n4928), .Z(c[3260]) );
  XNOR U5766 ( .A(a[3260]), .B(n4929), .Z(n4928) );
  IV U5767 ( .A(n4926), .Z(n4929) );
  XOR U5768 ( .A(n4930), .B(n4931), .Z(n4926) );
  ANDN U5769 ( .B(n4932), .A(n4933), .Z(n4930) );
  XNOR U5770 ( .A(b[3259]), .B(n4931), .Z(n4932) );
  XNOR U5771 ( .A(b[325]), .B(n4934), .Z(c[325]) );
  XNOR U5772 ( .A(b[3259]), .B(n4933), .Z(c[3259]) );
  XNOR U5773 ( .A(a[3259]), .B(n4935), .Z(n4933) );
  IV U5774 ( .A(n4931), .Z(n4935) );
  XOR U5775 ( .A(n4936), .B(n4937), .Z(n4931) );
  ANDN U5776 ( .B(n4938), .A(n4939), .Z(n4936) );
  XNOR U5777 ( .A(b[3258]), .B(n4937), .Z(n4938) );
  XNOR U5778 ( .A(b[3258]), .B(n4939), .Z(c[3258]) );
  XNOR U5779 ( .A(a[3258]), .B(n4940), .Z(n4939) );
  IV U5780 ( .A(n4937), .Z(n4940) );
  XOR U5781 ( .A(n4941), .B(n4942), .Z(n4937) );
  ANDN U5782 ( .B(n4943), .A(n4944), .Z(n4941) );
  XNOR U5783 ( .A(b[3257]), .B(n4942), .Z(n4943) );
  XNOR U5784 ( .A(b[3257]), .B(n4944), .Z(c[3257]) );
  XNOR U5785 ( .A(a[3257]), .B(n4945), .Z(n4944) );
  IV U5786 ( .A(n4942), .Z(n4945) );
  XOR U5787 ( .A(n4946), .B(n4947), .Z(n4942) );
  ANDN U5788 ( .B(n4948), .A(n4949), .Z(n4946) );
  XNOR U5789 ( .A(b[3256]), .B(n4947), .Z(n4948) );
  XNOR U5790 ( .A(b[3256]), .B(n4949), .Z(c[3256]) );
  XNOR U5791 ( .A(a[3256]), .B(n4950), .Z(n4949) );
  IV U5792 ( .A(n4947), .Z(n4950) );
  XOR U5793 ( .A(n4951), .B(n4952), .Z(n4947) );
  ANDN U5794 ( .B(n4953), .A(n4954), .Z(n4951) );
  XNOR U5795 ( .A(b[3255]), .B(n4952), .Z(n4953) );
  XNOR U5796 ( .A(b[3255]), .B(n4954), .Z(c[3255]) );
  XNOR U5797 ( .A(a[3255]), .B(n4955), .Z(n4954) );
  IV U5798 ( .A(n4952), .Z(n4955) );
  XOR U5799 ( .A(n4956), .B(n4957), .Z(n4952) );
  ANDN U5800 ( .B(n4958), .A(n4959), .Z(n4956) );
  XNOR U5801 ( .A(b[3254]), .B(n4957), .Z(n4958) );
  XNOR U5802 ( .A(b[3254]), .B(n4959), .Z(c[3254]) );
  XNOR U5803 ( .A(a[3254]), .B(n4960), .Z(n4959) );
  IV U5804 ( .A(n4957), .Z(n4960) );
  XOR U5805 ( .A(n4961), .B(n4962), .Z(n4957) );
  ANDN U5806 ( .B(n4963), .A(n4964), .Z(n4961) );
  XNOR U5807 ( .A(b[3253]), .B(n4962), .Z(n4963) );
  XNOR U5808 ( .A(b[3253]), .B(n4964), .Z(c[3253]) );
  XNOR U5809 ( .A(a[3253]), .B(n4965), .Z(n4964) );
  IV U5810 ( .A(n4962), .Z(n4965) );
  XOR U5811 ( .A(n4966), .B(n4967), .Z(n4962) );
  ANDN U5812 ( .B(n4968), .A(n4969), .Z(n4966) );
  XNOR U5813 ( .A(b[3252]), .B(n4967), .Z(n4968) );
  XNOR U5814 ( .A(b[3252]), .B(n4969), .Z(c[3252]) );
  XNOR U5815 ( .A(a[3252]), .B(n4970), .Z(n4969) );
  IV U5816 ( .A(n4967), .Z(n4970) );
  XOR U5817 ( .A(n4971), .B(n4972), .Z(n4967) );
  ANDN U5818 ( .B(n4973), .A(n4974), .Z(n4971) );
  XNOR U5819 ( .A(b[3251]), .B(n4972), .Z(n4973) );
  XNOR U5820 ( .A(b[3251]), .B(n4974), .Z(c[3251]) );
  XNOR U5821 ( .A(a[3251]), .B(n4975), .Z(n4974) );
  IV U5822 ( .A(n4972), .Z(n4975) );
  XOR U5823 ( .A(n4976), .B(n4977), .Z(n4972) );
  ANDN U5824 ( .B(n4978), .A(n4979), .Z(n4976) );
  XNOR U5825 ( .A(b[3250]), .B(n4977), .Z(n4978) );
  XNOR U5826 ( .A(b[3250]), .B(n4979), .Z(c[3250]) );
  XNOR U5827 ( .A(a[3250]), .B(n4980), .Z(n4979) );
  IV U5828 ( .A(n4977), .Z(n4980) );
  XOR U5829 ( .A(n4981), .B(n4982), .Z(n4977) );
  ANDN U5830 ( .B(n4983), .A(n4984), .Z(n4981) );
  XNOR U5831 ( .A(b[3249]), .B(n4982), .Z(n4983) );
  XNOR U5832 ( .A(b[324]), .B(n4985), .Z(c[324]) );
  XNOR U5833 ( .A(b[3249]), .B(n4984), .Z(c[3249]) );
  XNOR U5834 ( .A(a[3249]), .B(n4986), .Z(n4984) );
  IV U5835 ( .A(n4982), .Z(n4986) );
  XOR U5836 ( .A(n4987), .B(n4988), .Z(n4982) );
  ANDN U5837 ( .B(n4989), .A(n4990), .Z(n4987) );
  XNOR U5838 ( .A(b[3248]), .B(n4988), .Z(n4989) );
  XNOR U5839 ( .A(b[3248]), .B(n4990), .Z(c[3248]) );
  XNOR U5840 ( .A(a[3248]), .B(n4991), .Z(n4990) );
  IV U5841 ( .A(n4988), .Z(n4991) );
  XOR U5842 ( .A(n4992), .B(n4993), .Z(n4988) );
  ANDN U5843 ( .B(n4994), .A(n4995), .Z(n4992) );
  XNOR U5844 ( .A(b[3247]), .B(n4993), .Z(n4994) );
  XNOR U5845 ( .A(b[3247]), .B(n4995), .Z(c[3247]) );
  XNOR U5846 ( .A(a[3247]), .B(n4996), .Z(n4995) );
  IV U5847 ( .A(n4993), .Z(n4996) );
  XOR U5848 ( .A(n4997), .B(n4998), .Z(n4993) );
  ANDN U5849 ( .B(n4999), .A(n5000), .Z(n4997) );
  XNOR U5850 ( .A(b[3246]), .B(n4998), .Z(n4999) );
  XNOR U5851 ( .A(b[3246]), .B(n5000), .Z(c[3246]) );
  XNOR U5852 ( .A(a[3246]), .B(n5001), .Z(n5000) );
  IV U5853 ( .A(n4998), .Z(n5001) );
  XOR U5854 ( .A(n5002), .B(n5003), .Z(n4998) );
  ANDN U5855 ( .B(n5004), .A(n5005), .Z(n5002) );
  XNOR U5856 ( .A(b[3245]), .B(n5003), .Z(n5004) );
  XNOR U5857 ( .A(b[3245]), .B(n5005), .Z(c[3245]) );
  XNOR U5858 ( .A(a[3245]), .B(n5006), .Z(n5005) );
  IV U5859 ( .A(n5003), .Z(n5006) );
  XOR U5860 ( .A(n5007), .B(n5008), .Z(n5003) );
  ANDN U5861 ( .B(n5009), .A(n5010), .Z(n5007) );
  XNOR U5862 ( .A(b[3244]), .B(n5008), .Z(n5009) );
  XNOR U5863 ( .A(b[3244]), .B(n5010), .Z(c[3244]) );
  XNOR U5864 ( .A(a[3244]), .B(n5011), .Z(n5010) );
  IV U5865 ( .A(n5008), .Z(n5011) );
  XOR U5866 ( .A(n5012), .B(n5013), .Z(n5008) );
  ANDN U5867 ( .B(n5014), .A(n5015), .Z(n5012) );
  XNOR U5868 ( .A(b[3243]), .B(n5013), .Z(n5014) );
  XNOR U5869 ( .A(b[3243]), .B(n5015), .Z(c[3243]) );
  XNOR U5870 ( .A(a[3243]), .B(n5016), .Z(n5015) );
  IV U5871 ( .A(n5013), .Z(n5016) );
  XOR U5872 ( .A(n5017), .B(n5018), .Z(n5013) );
  ANDN U5873 ( .B(n5019), .A(n5020), .Z(n5017) );
  XNOR U5874 ( .A(b[3242]), .B(n5018), .Z(n5019) );
  XNOR U5875 ( .A(b[3242]), .B(n5020), .Z(c[3242]) );
  XNOR U5876 ( .A(a[3242]), .B(n5021), .Z(n5020) );
  IV U5877 ( .A(n5018), .Z(n5021) );
  XOR U5878 ( .A(n5022), .B(n5023), .Z(n5018) );
  ANDN U5879 ( .B(n5024), .A(n5025), .Z(n5022) );
  XNOR U5880 ( .A(b[3241]), .B(n5023), .Z(n5024) );
  XNOR U5881 ( .A(b[3241]), .B(n5025), .Z(c[3241]) );
  XNOR U5882 ( .A(a[3241]), .B(n5026), .Z(n5025) );
  IV U5883 ( .A(n5023), .Z(n5026) );
  XOR U5884 ( .A(n5027), .B(n5028), .Z(n5023) );
  ANDN U5885 ( .B(n5029), .A(n5030), .Z(n5027) );
  XNOR U5886 ( .A(b[3240]), .B(n5028), .Z(n5029) );
  XNOR U5887 ( .A(b[3240]), .B(n5030), .Z(c[3240]) );
  XNOR U5888 ( .A(a[3240]), .B(n5031), .Z(n5030) );
  IV U5889 ( .A(n5028), .Z(n5031) );
  XOR U5890 ( .A(n5032), .B(n5033), .Z(n5028) );
  ANDN U5891 ( .B(n5034), .A(n5035), .Z(n5032) );
  XNOR U5892 ( .A(b[3239]), .B(n5033), .Z(n5034) );
  XNOR U5893 ( .A(b[323]), .B(n5036), .Z(c[323]) );
  XNOR U5894 ( .A(b[3239]), .B(n5035), .Z(c[3239]) );
  XNOR U5895 ( .A(a[3239]), .B(n5037), .Z(n5035) );
  IV U5896 ( .A(n5033), .Z(n5037) );
  XOR U5897 ( .A(n5038), .B(n5039), .Z(n5033) );
  ANDN U5898 ( .B(n5040), .A(n5041), .Z(n5038) );
  XNOR U5899 ( .A(b[3238]), .B(n5039), .Z(n5040) );
  XNOR U5900 ( .A(b[3238]), .B(n5041), .Z(c[3238]) );
  XNOR U5901 ( .A(a[3238]), .B(n5042), .Z(n5041) );
  IV U5902 ( .A(n5039), .Z(n5042) );
  XOR U5903 ( .A(n5043), .B(n5044), .Z(n5039) );
  ANDN U5904 ( .B(n5045), .A(n5046), .Z(n5043) );
  XNOR U5905 ( .A(b[3237]), .B(n5044), .Z(n5045) );
  XNOR U5906 ( .A(b[3237]), .B(n5046), .Z(c[3237]) );
  XNOR U5907 ( .A(a[3237]), .B(n5047), .Z(n5046) );
  IV U5908 ( .A(n5044), .Z(n5047) );
  XOR U5909 ( .A(n5048), .B(n5049), .Z(n5044) );
  ANDN U5910 ( .B(n5050), .A(n5051), .Z(n5048) );
  XNOR U5911 ( .A(b[3236]), .B(n5049), .Z(n5050) );
  XNOR U5912 ( .A(b[3236]), .B(n5051), .Z(c[3236]) );
  XNOR U5913 ( .A(a[3236]), .B(n5052), .Z(n5051) );
  IV U5914 ( .A(n5049), .Z(n5052) );
  XOR U5915 ( .A(n5053), .B(n5054), .Z(n5049) );
  ANDN U5916 ( .B(n5055), .A(n5056), .Z(n5053) );
  XNOR U5917 ( .A(b[3235]), .B(n5054), .Z(n5055) );
  XNOR U5918 ( .A(b[3235]), .B(n5056), .Z(c[3235]) );
  XNOR U5919 ( .A(a[3235]), .B(n5057), .Z(n5056) );
  IV U5920 ( .A(n5054), .Z(n5057) );
  XOR U5921 ( .A(n5058), .B(n5059), .Z(n5054) );
  ANDN U5922 ( .B(n5060), .A(n5061), .Z(n5058) );
  XNOR U5923 ( .A(b[3234]), .B(n5059), .Z(n5060) );
  XNOR U5924 ( .A(b[3234]), .B(n5061), .Z(c[3234]) );
  XNOR U5925 ( .A(a[3234]), .B(n5062), .Z(n5061) );
  IV U5926 ( .A(n5059), .Z(n5062) );
  XOR U5927 ( .A(n5063), .B(n5064), .Z(n5059) );
  ANDN U5928 ( .B(n5065), .A(n5066), .Z(n5063) );
  XNOR U5929 ( .A(b[3233]), .B(n5064), .Z(n5065) );
  XNOR U5930 ( .A(b[3233]), .B(n5066), .Z(c[3233]) );
  XNOR U5931 ( .A(a[3233]), .B(n5067), .Z(n5066) );
  IV U5932 ( .A(n5064), .Z(n5067) );
  XOR U5933 ( .A(n5068), .B(n5069), .Z(n5064) );
  ANDN U5934 ( .B(n5070), .A(n5071), .Z(n5068) );
  XNOR U5935 ( .A(b[3232]), .B(n5069), .Z(n5070) );
  XNOR U5936 ( .A(b[3232]), .B(n5071), .Z(c[3232]) );
  XNOR U5937 ( .A(a[3232]), .B(n5072), .Z(n5071) );
  IV U5938 ( .A(n5069), .Z(n5072) );
  XOR U5939 ( .A(n5073), .B(n5074), .Z(n5069) );
  ANDN U5940 ( .B(n5075), .A(n5076), .Z(n5073) );
  XNOR U5941 ( .A(b[3231]), .B(n5074), .Z(n5075) );
  XNOR U5942 ( .A(b[3231]), .B(n5076), .Z(c[3231]) );
  XNOR U5943 ( .A(a[3231]), .B(n5077), .Z(n5076) );
  IV U5944 ( .A(n5074), .Z(n5077) );
  XOR U5945 ( .A(n5078), .B(n5079), .Z(n5074) );
  ANDN U5946 ( .B(n5080), .A(n5081), .Z(n5078) );
  XNOR U5947 ( .A(b[3230]), .B(n5079), .Z(n5080) );
  XNOR U5948 ( .A(b[3230]), .B(n5081), .Z(c[3230]) );
  XNOR U5949 ( .A(a[3230]), .B(n5082), .Z(n5081) );
  IV U5950 ( .A(n5079), .Z(n5082) );
  XOR U5951 ( .A(n5083), .B(n5084), .Z(n5079) );
  ANDN U5952 ( .B(n5085), .A(n5086), .Z(n5083) );
  XNOR U5953 ( .A(b[3229]), .B(n5084), .Z(n5085) );
  XNOR U5954 ( .A(b[322]), .B(n5087), .Z(c[322]) );
  XNOR U5955 ( .A(b[3229]), .B(n5086), .Z(c[3229]) );
  XNOR U5956 ( .A(a[3229]), .B(n5088), .Z(n5086) );
  IV U5957 ( .A(n5084), .Z(n5088) );
  XOR U5958 ( .A(n5089), .B(n5090), .Z(n5084) );
  ANDN U5959 ( .B(n5091), .A(n5092), .Z(n5089) );
  XNOR U5960 ( .A(b[3228]), .B(n5090), .Z(n5091) );
  XNOR U5961 ( .A(b[3228]), .B(n5092), .Z(c[3228]) );
  XNOR U5962 ( .A(a[3228]), .B(n5093), .Z(n5092) );
  IV U5963 ( .A(n5090), .Z(n5093) );
  XOR U5964 ( .A(n5094), .B(n5095), .Z(n5090) );
  ANDN U5965 ( .B(n5096), .A(n5097), .Z(n5094) );
  XNOR U5966 ( .A(b[3227]), .B(n5095), .Z(n5096) );
  XNOR U5967 ( .A(b[3227]), .B(n5097), .Z(c[3227]) );
  XNOR U5968 ( .A(a[3227]), .B(n5098), .Z(n5097) );
  IV U5969 ( .A(n5095), .Z(n5098) );
  XOR U5970 ( .A(n5099), .B(n5100), .Z(n5095) );
  ANDN U5971 ( .B(n5101), .A(n5102), .Z(n5099) );
  XNOR U5972 ( .A(b[3226]), .B(n5100), .Z(n5101) );
  XNOR U5973 ( .A(b[3226]), .B(n5102), .Z(c[3226]) );
  XNOR U5974 ( .A(a[3226]), .B(n5103), .Z(n5102) );
  IV U5975 ( .A(n5100), .Z(n5103) );
  XOR U5976 ( .A(n5104), .B(n5105), .Z(n5100) );
  ANDN U5977 ( .B(n5106), .A(n5107), .Z(n5104) );
  XNOR U5978 ( .A(b[3225]), .B(n5105), .Z(n5106) );
  XNOR U5979 ( .A(b[3225]), .B(n5107), .Z(c[3225]) );
  XNOR U5980 ( .A(a[3225]), .B(n5108), .Z(n5107) );
  IV U5981 ( .A(n5105), .Z(n5108) );
  XOR U5982 ( .A(n5109), .B(n5110), .Z(n5105) );
  ANDN U5983 ( .B(n5111), .A(n5112), .Z(n5109) );
  XNOR U5984 ( .A(b[3224]), .B(n5110), .Z(n5111) );
  XNOR U5985 ( .A(b[3224]), .B(n5112), .Z(c[3224]) );
  XNOR U5986 ( .A(a[3224]), .B(n5113), .Z(n5112) );
  IV U5987 ( .A(n5110), .Z(n5113) );
  XOR U5988 ( .A(n5114), .B(n5115), .Z(n5110) );
  ANDN U5989 ( .B(n5116), .A(n5117), .Z(n5114) );
  XNOR U5990 ( .A(b[3223]), .B(n5115), .Z(n5116) );
  XNOR U5991 ( .A(b[3223]), .B(n5117), .Z(c[3223]) );
  XNOR U5992 ( .A(a[3223]), .B(n5118), .Z(n5117) );
  IV U5993 ( .A(n5115), .Z(n5118) );
  XOR U5994 ( .A(n5119), .B(n5120), .Z(n5115) );
  ANDN U5995 ( .B(n5121), .A(n5122), .Z(n5119) );
  XNOR U5996 ( .A(b[3222]), .B(n5120), .Z(n5121) );
  XNOR U5997 ( .A(b[3222]), .B(n5122), .Z(c[3222]) );
  XNOR U5998 ( .A(a[3222]), .B(n5123), .Z(n5122) );
  IV U5999 ( .A(n5120), .Z(n5123) );
  XOR U6000 ( .A(n5124), .B(n5125), .Z(n5120) );
  ANDN U6001 ( .B(n5126), .A(n5127), .Z(n5124) );
  XNOR U6002 ( .A(b[3221]), .B(n5125), .Z(n5126) );
  XNOR U6003 ( .A(b[3221]), .B(n5127), .Z(c[3221]) );
  XNOR U6004 ( .A(a[3221]), .B(n5128), .Z(n5127) );
  IV U6005 ( .A(n5125), .Z(n5128) );
  XOR U6006 ( .A(n5129), .B(n5130), .Z(n5125) );
  ANDN U6007 ( .B(n5131), .A(n5132), .Z(n5129) );
  XNOR U6008 ( .A(b[3220]), .B(n5130), .Z(n5131) );
  XNOR U6009 ( .A(b[3220]), .B(n5132), .Z(c[3220]) );
  XNOR U6010 ( .A(a[3220]), .B(n5133), .Z(n5132) );
  IV U6011 ( .A(n5130), .Z(n5133) );
  XOR U6012 ( .A(n5134), .B(n5135), .Z(n5130) );
  ANDN U6013 ( .B(n5136), .A(n5137), .Z(n5134) );
  XNOR U6014 ( .A(b[3219]), .B(n5135), .Z(n5136) );
  XNOR U6015 ( .A(b[321]), .B(n5138), .Z(c[321]) );
  XNOR U6016 ( .A(b[3219]), .B(n5137), .Z(c[3219]) );
  XNOR U6017 ( .A(a[3219]), .B(n5139), .Z(n5137) );
  IV U6018 ( .A(n5135), .Z(n5139) );
  XOR U6019 ( .A(n5140), .B(n5141), .Z(n5135) );
  ANDN U6020 ( .B(n5142), .A(n5143), .Z(n5140) );
  XNOR U6021 ( .A(b[3218]), .B(n5141), .Z(n5142) );
  XNOR U6022 ( .A(b[3218]), .B(n5143), .Z(c[3218]) );
  XNOR U6023 ( .A(a[3218]), .B(n5144), .Z(n5143) );
  IV U6024 ( .A(n5141), .Z(n5144) );
  XOR U6025 ( .A(n5145), .B(n5146), .Z(n5141) );
  ANDN U6026 ( .B(n5147), .A(n5148), .Z(n5145) );
  XNOR U6027 ( .A(b[3217]), .B(n5146), .Z(n5147) );
  XNOR U6028 ( .A(b[3217]), .B(n5148), .Z(c[3217]) );
  XNOR U6029 ( .A(a[3217]), .B(n5149), .Z(n5148) );
  IV U6030 ( .A(n5146), .Z(n5149) );
  XOR U6031 ( .A(n5150), .B(n5151), .Z(n5146) );
  ANDN U6032 ( .B(n5152), .A(n5153), .Z(n5150) );
  XNOR U6033 ( .A(b[3216]), .B(n5151), .Z(n5152) );
  XNOR U6034 ( .A(b[3216]), .B(n5153), .Z(c[3216]) );
  XNOR U6035 ( .A(a[3216]), .B(n5154), .Z(n5153) );
  IV U6036 ( .A(n5151), .Z(n5154) );
  XOR U6037 ( .A(n5155), .B(n5156), .Z(n5151) );
  ANDN U6038 ( .B(n5157), .A(n5158), .Z(n5155) );
  XNOR U6039 ( .A(b[3215]), .B(n5156), .Z(n5157) );
  XNOR U6040 ( .A(b[3215]), .B(n5158), .Z(c[3215]) );
  XNOR U6041 ( .A(a[3215]), .B(n5159), .Z(n5158) );
  IV U6042 ( .A(n5156), .Z(n5159) );
  XOR U6043 ( .A(n5160), .B(n5161), .Z(n5156) );
  ANDN U6044 ( .B(n5162), .A(n5163), .Z(n5160) );
  XNOR U6045 ( .A(b[3214]), .B(n5161), .Z(n5162) );
  XNOR U6046 ( .A(b[3214]), .B(n5163), .Z(c[3214]) );
  XNOR U6047 ( .A(a[3214]), .B(n5164), .Z(n5163) );
  IV U6048 ( .A(n5161), .Z(n5164) );
  XOR U6049 ( .A(n5165), .B(n5166), .Z(n5161) );
  ANDN U6050 ( .B(n5167), .A(n5168), .Z(n5165) );
  XNOR U6051 ( .A(b[3213]), .B(n5166), .Z(n5167) );
  XNOR U6052 ( .A(b[3213]), .B(n5168), .Z(c[3213]) );
  XNOR U6053 ( .A(a[3213]), .B(n5169), .Z(n5168) );
  IV U6054 ( .A(n5166), .Z(n5169) );
  XOR U6055 ( .A(n5170), .B(n5171), .Z(n5166) );
  ANDN U6056 ( .B(n5172), .A(n5173), .Z(n5170) );
  XNOR U6057 ( .A(b[3212]), .B(n5171), .Z(n5172) );
  XNOR U6058 ( .A(b[3212]), .B(n5173), .Z(c[3212]) );
  XNOR U6059 ( .A(a[3212]), .B(n5174), .Z(n5173) );
  IV U6060 ( .A(n5171), .Z(n5174) );
  XOR U6061 ( .A(n5175), .B(n5176), .Z(n5171) );
  ANDN U6062 ( .B(n5177), .A(n5178), .Z(n5175) );
  XNOR U6063 ( .A(b[3211]), .B(n5176), .Z(n5177) );
  XNOR U6064 ( .A(b[3211]), .B(n5178), .Z(c[3211]) );
  XNOR U6065 ( .A(a[3211]), .B(n5179), .Z(n5178) );
  IV U6066 ( .A(n5176), .Z(n5179) );
  XOR U6067 ( .A(n5180), .B(n5181), .Z(n5176) );
  ANDN U6068 ( .B(n5182), .A(n5183), .Z(n5180) );
  XNOR U6069 ( .A(b[3210]), .B(n5181), .Z(n5182) );
  XNOR U6070 ( .A(b[3210]), .B(n5183), .Z(c[3210]) );
  XNOR U6071 ( .A(a[3210]), .B(n5184), .Z(n5183) );
  IV U6072 ( .A(n5181), .Z(n5184) );
  XOR U6073 ( .A(n5185), .B(n5186), .Z(n5181) );
  ANDN U6074 ( .B(n5187), .A(n5188), .Z(n5185) );
  XNOR U6075 ( .A(b[3209]), .B(n5186), .Z(n5187) );
  XNOR U6076 ( .A(b[320]), .B(n5189), .Z(c[320]) );
  XNOR U6077 ( .A(b[3209]), .B(n5188), .Z(c[3209]) );
  XNOR U6078 ( .A(a[3209]), .B(n5190), .Z(n5188) );
  IV U6079 ( .A(n5186), .Z(n5190) );
  XOR U6080 ( .A(n5191), .B(n5192), .Z(n5186) );
  ANDN U6081 ( .B(n5193), .A(n5194), .Z(n5191) );
  XNOR U6082 ( .A(b[3208]), .B(n5192), .Z(n5193) );
  XNOR U6083 ( .A(b[3208]), .B(n5194), .Z(c[3208]) );
  XNOR U6084 ( .A(a[3208]), .B(n5195), .Z(n5194) );
  IV U6085 ( .A(n5192), .Z(n5195) );
  XOR U6086 ( .A(n5196), .B(n5197), .Z(n5192) );
  ANDN U6087 ( .B(n5198), .A(n5199), .Z(n5196) );
  XNOR U6088 ( .A(b[3207]), .B(n5197), .Z(n5198) );
  XNOR U6089 ( .A(b[3207]), .B(n5199), .Z(c[3207]) );
  XNOR U6090 ( .A(a[3207]), .B(n5200), .Z(n5199) );
  IV U6091 ( .A(n5197), .Z(n5200) );
  XOR U6092 ( .A(n5201), .B(n5202), .Z(n5197) );
  ANDN U6093 ( .B(n5203), .A(n5204), .Z(n5201) );
  XNOR U6094 ( .A(b[3206]), .B(n5202), .Z(n5203) );
  XNOR U6095 ( .A(b[3206]), .B(n5204), .Z(c[3206]) );
  XNOR U6096 ( .A(a[3206]), .B(n5205), .Z(n5204) );
  IV U6097 ( .A(n5202), .Z(n5205) );
  XOR U6098 ( .A(n5206), .B(n5207), .Z(n5202) );
  ANDN U6099 ( .B(n5208), .A(n5209), .Z(n5206) );
  XNOR U6100 ( .A(b[3205]), .B(n5207), .Z(n5208) );
  XNOR U6101 ( .A(b[3205]), .B(n5209), .Z(c[3205]) );
  XNOR U6102 ( .A(a[3205]), .B(n5210), .Z(n5209) );
  IV U6103 ( .A(n5207), .Z(n5210) );
  XOR U6104 ( .A(n5211), .B(n5212), .Z(n5207) );
  ANDN U6105 ( .B(n5213), .A(n5214), .Z(n5211) );
  XNOR U6106 ( .A(b[3204]), .B(n5212), .Z(n5213) );
  XNOR U6107 ( .A(b[3204]), .B(n5214), .Z(c[3204]) );
  XNOR U6108 ( .A(a[3204]), .B(n5215), .Z(n5214) );
  IV U6109 ( .A(n5212), .Z(n5215) );
  XOR U6110 ( .A(n5216), .B(n5217), .Z(n5212) );
  ANDN U6111 ( .B(n5218), .A(n5219), .Z(n5216) );
  XNOR U6112 ( .A(b[3203]), .B(n5217), .Z(n5218) );
  XNOR U6113 ( .A(b[3203]), .B(n5219), .Z(c[3203]) );
  XNOR U6114 ( .A(a[3203]), .B(n5220), .Z(n5219) );
  IV U6115 ( .A(n5217), .Z(n5220) );
  XOR U6116 ( .A(n5221), .B(n5222), .Z(n5217) );
  ANDN U6117 ( .B(n5223), .A(n5224), .Z(n5221) );
  XNOR U6118 ( .A(b[3202]), .B(n5222), .Z(n5223) );
  XNOR U6119 ( .A(b[3202]), .B(n5224), .Z(c[3202]) );
  XNOR U6120 ( .A(a[3202]), .B(n5225), .Z(n5224) );
  IV U6121 ( .A(n5222), .Z(n5225) );
  XOR U6122 ( .A(n5226), .B(n5227), .Z(n5222) );
  ANDN U6123 ( .B(n5228), .A(n5229), .Z(n5226) );
  XNOR U6124 ( .A(b[3201]), .B(n5227), .Z(n5228) );
  XNOR U6125 ( .A(b[3201]), .B(n5229), .Z(c[3201]) );
  XNOR U6126 ( .A(a[3201]), .B(n5230), .Z(n5229) );
  IV U6127 ( .A(n5227), .Z(n5230) );
  XOR U6128 ( .A(n5231), .B(n5232), .Z(n5227) );
  ANDN U6129 ( .B(n5233), .A(n5234), .Z(n5231) );
  XNOR U6130 ( .A(b[3200]), .B(n5232), .Z(n5233) );
  XNOR U6131 ( .A(b[3200]), .B(n5234), .Z(c[3200]) );
  XNOR U6132 ( .A(a[3200]), .B(n5235), .Z(n5234) );
  IV U6133 ( .A(n5232), .Z(n5235) );
  XOR U6134 ( .A(n5236), .B(n5237), .Z(n5232) );
  ANDN U6135 ( .B(n5238), .A(n5239), .Z(n5236) );
  XNOR U6136 ( .A(b[3199]), .B(n5237), .Z(n5238) );
  XNOR U6137 ( .A(b[31]), .B(n5240), .Z(c[31]) );
  XNOR U6138 ( .A(b[319]), .B(n5241), .Z(c[319]) );
  XNOR U6139 ( .A(b[3199]), .B(n5239), .Z(c[3199]) );
  XNOR U6140 ( .A(a[3199]), .B(n5242), .Z(n5239) );
  IV U6141 ( .A(n5237), .Z(n5242) );
  XOR U6142 ( .A(n5243), .B(n5244), .Z(n5237) );
  ANDN U6143 ( .B(n5245), .A(n5246), .Z(n5243) );
  XNOR U6144 ( .A(b[3198]), .B(n5244), .Z(n5245) );
  XNOR U6145 ( .A(b[3198]), .B(n5246), .Z(c[3198]) );
  XNOR U6146 ( .A(a[3198]), .B(n5247), .Z(n5246) );
  IV U6147 ( .A(n5244), .Z(n5247) );
  XOR U6148 ( .A(n5248), .B(n5249), .Z(n5244) );
  ANDN U6149 ( .B(n5250), .A(n5251), .Z(n5248) );
  XNOR U6150 ( .A(b[3197]), .B(n5249), .Z(n5250) );
  XNOR U6151 ( .A(b[3197]), .B(n5251), .Z(c[3197]) );
  XNOR U6152 ( .A(a[3197]), .B(n5252), .Z(n5251) );
  IV U6153 ( .A(n5249), .Z(n5252) );
  XOR U6154 ( .A(n5253), .B(n5254), .Z(n5249) );
  ANDN U6155 ( .B(n5255), .A(n5256), .Z(n5253) );
  XNOR U6156 ( .A(b[3196]), .B(n5254), .Z(n5255) );
  XNOR U6157 ( .A(b[3196]), .B(n5256), .Z(c[3196]) );
  XNOR U6158 ( .A(a[3196]), .B(n5257), .Z(n5256) );
  IV U6159 ( .A(n5254), .Z(n5257) );
  XOR U6160 ( .A(n5258), .B(n5259), .Z(n5254) );
  ANDN U6161 ( .B(n5260), .A(n5261), .Z(n5258) );
  XNOR U6162 ( .A(b[3195]), .B(n5259), .Z(n5260) );
  XNOR U6163 ( .A(b[3195]), .B(n5261), .Z(c[3195]) );
  XNOR U6164 ( .A(a[3195]), .B(n5262), .Z(n5261) );
  IV U6165 ( .A(n5259), .Z(n5262) );
  XOR U6166 ( .A(n5263), .B(n5264), .Z(n5259) );
  ANDN U6167 ( .B(n5265), .A(n5266), .Z(n5263) );
  XNOR U6168 ( .A(b[3194]), .B(n5264), .Z(n5265) );
  XNOR U6169 ( .A(b[3194]), .B(n5266), .Z(c[3194]) );
  XNOR U6170 ( .A(a[3194]), .B(n5267), .Z(n5266) );
  IV U6171 ( .A(n5264), .Z(n5267) );
  XOR U6172 ( .A(n5268), .B(n5269), .Z(n5264) );
  ANDN U6173 ( .B(n5270), .A(n5271), .Z(n5268) );
  XNOR U6174 ( .A(b[3193]), .B(n5269), .Z(n5270) );
  XNOR U6175 ( .A(b[3193]), .B(n5271), .Z(c[3193]) );
  XNOR U6176 ( .A(a[3193]), .B(n5272), .Z(n5271) );
  IV U6177 ( .A(n5269), .Z(n5272) );
  XOR U6178 ( .A(n5273), .B(n5274), .Z(n5269) );
  ANDN U6179 ( .B(n5275), .A(n5276), .Z(n5273) );
  XNOR U6180 ( .A(b[3192]), .B(n5274), .Z(n5275) );
  XNOR U6181 ( .A(b[3192]), .B(n5276), .Z(c[3192]) );
  XNOR U6182 ( .A(a[3192]), .B(n5277), .Z(n5276) );
  IV U6183 ( .A(n5274), .Z(n5277) );
  XOR U6184 ( .A(n5278), .B(n5279), .Z(n5274) );
  ANDN U6185 ( .B(n5280), .A(n5281), .Z(n5278) );
  XNOR U6186 ( .A(b[3191]), .B(n5279), .Z(n5280) );
  XNOR U6187 ( .A(b[3191]), .B(n5281), .Z(c[3191]) );
  XNOR U6188 ( .A(a[3191]), .B(n5282), .Z(n5281) );
  IV U6189 ( .A(n5279), .Z(n5282) );
  XOR U6190 ( .A(n5283), .B(n5284), .Z(n5279) );
  ANDN U6191 ( .B(n5285), .A(n5286), .Z(n5283) );
  XNOR U6192 ( .A(b[3190]), .B(n5284), .Z(n5285) );
  XNOR U6193 ( .A(b[3190]), .B(n5286), .Z(c[3190]) );
  XNOR U6194 ( .A(a[3190]), .B(n5287), .Z(n5286) );
  IV U6195 ( .A(n5284), .Z(n5287) );
  XOR U6196 ( .A(n5288), .B(n5289), .Z(n5284) );
  ANDN U6197 ( .B(n5290), .A(n5291), .Z(n5288) );
  XNOR U6198 ( .A(b[3189]), .B(n5289), .Z(n5290) );
  XNOR U6199 ( .A(b[318]), .B(n5292), .Z(c[318]) );
  XNOR U6200 ( .A(b[3189]), .B(n5291), .Z(c[3189]) );
  XNOR U6201 ( .A(a[3189]), .B(n5293), .Z(n5291) );
  IV U6202 ( .A(n5289), .Z(n5293) );
  XOR U6203 ( .A(n5294), .B(n5295), .Z(n5289) );
  ANDN U6204 ( .B(n5296), .A(n5297), .Z(n5294) );
  XNOR U6205 ( .A(b[3188]), .B(n5295), .Z(n5296) );
  XNOR U6206 ( .A(b[3188]), .B(n5297), .Z(c[3188]) );
  XNOR U6207 ( .A(a[3188]), .B(n5298), .Z(n5297) );
  IV U6208 ( .A(n5295), .Z(n5298) );
  XOR U6209 ( .A(n5299), .B(n5300), .Z(n5295) );
  ANDN U6210 ( .B(n5301), .A(n5302), .Z(n5299) );
  XNOR U6211 ( .A(b[3187]), .B(n5300), .Z(n5301) );
  XNOR U6212 ( .A(b[3187]), .B(n5302), .Z(c[3187]) );
  XNOR U6213 ( .A(a[3187]), .B(n5303), .Z(n5302) );
  IV U6214 ( .A(n5300), .Z(n5303) );
  XOR U6215 ( .A(n5304), .B(n5305), .Z(n5300) );
  ANDN U6216 ( .B(n5306), .A(n5307), .Z(n5304) );
  XNOR U6217 ( .A(b[3186]), .B(n5305), .Z(n5306) );
  XNOR U6218 ( .A(b[3186]), .B(n5307), .Z(c[3186]) );
  XNOR U6219 ( .A(a[3186]), .B(n5308), .Z(n5307) );
  IV U6220 ( .A(n5305), .Z(n5308) );
  XOR U6221 ( .A(n5309), .B(n5310), .Z(n5305) );
  ANDN U6222 ( .B(n5311), .A(n5312), .Z(n5309) );
  XNOR U6223 ( .A(b[3185]), .B(n5310), .Z(n5311) );
  XNOR U6224 ( .A(b[3185]), .B(n5312), .Z(c[3185]) );
  XNOR U6225 ( .A(a[3185]), .B(n5313), .Z(n5312) );
  IV U6226 ( .A(n5310), .Z(n5313) );
  XOR U6227 ( .A(n5314), .B(n5315), .Z(n5310) );
  ANDN U6228 ( .B(n5316), .A(n5317), .Z(n5314) );
  XNOR U6229 ( .A(b[3184]), .B(n5315), .Z(n5316) );
  XNOR U6230 ( .A(b[3184]), .B(n5317), .Z(c[3184]) );
  XNOR U6231 ( .A(a[3184]), .B(n5318), .Z(n5317) );
  IV U6232 ( .A(n5315), .Z(n5318) );
  XOR U6233 ( .A(n5319), .B(n5320), .Z(n5315) );
  ANDN U6234 ( .B(n5321), .A(n5322), .Z(n5319) );
  XNOR U6235 ( .A(b[3183]), .B(n5320), .Z(n5321) );
  XNOR U6236 ( .A(b[3183]), .B(n5322), .Z(c[3183]) );
  XNOR U6237 ( .A(a[3183]), .B(n5323), .Z(n5322) );
  IV U6238 ( .A(n5320), .Z(n5323) );
  XOR U6239 ( .A(n5324), .B(n5325), .Z(n5320) );
  ANDN U6240 ( .B(n5326), .A(n5327), .Z(n5324) );
  XNOR U6241 ( .A(b[3182]), .B(n5325), .Z(n5326) );
  XNOR U6242 ( .A(b[3182]), .B(n5327), .Z(c[3182]) );
  XNOR U6243 ( .A(a[3182]), .B(n5328), .Z(n5327) );
  IV U6244 ( .A(n5325), .Z(n5328) );
  XOR U6245 ( .A(n5329), .B(n5330), .Z(n5325) );
  ANDN U6246 ( .B(n5331), .A(n5332), .Z(n5329) );
  XNOR U6247 ( .A(b[3181]), .B(n5330), .Z(n5331) );
  XNOR U6248 ( .A(b[3181]), .B(n5332), .Z(c[3181]) );
  XNOR U6249 ( .A(a[3181]), .B(n5333), .Z(n5332) );
  IV U6250 ( .A(n5330), .Z(n5333) );
  XOR U6251 ( .A(n5334), .B(n5335), .Z(n5330) );
  ANDN U6252 ( .B(n5336), .A(n5337), .Z(n5334) );
  XNOR U6253 ( .A(b[3180]), .B(n5335), .Z(n5336) );
  XNOR U6254 ( .A(b[3180]), .B(n5337), .Z(c[3180]) );
  XNOR U6255 ( .A(a[3180]), .B(n5338), .Z(n5337) );
  IV U6256 ( .A(n5335), .Z(n5338) );
  XOR U6257 ( .A(n5339), .B(n5340), .Z(n5335) );
  ANDN U6258 ( .B(n5341), .A(n5342), .Z(n5339) );
  XNOR U6259 ( .A(b[3179]), .B(n5340), .Z(n5341) );
  XNOR U6260 ( .A(b[317]), .B(n5343), .Z(c[317]) );
  XNOR U6261 ( .A(b[3179]), .B(n5342), .Z(c[3179]) );
  XNOR U6262 ( .A(a[3179]), .B(n5344), .Z(n5342) );
  IV U6263 ( .A(n5340), .Z(n5344) );
  XOR U6264 ( .A(n5345), .B(n5346), .Z(n5340) );
  ANDN U6265 ( .B(n5347), .A(n5348), .Z(n5345) );
  XNOR U6266 ( .A(b[3178]), .B(n5346), .Z(n5347) );
  XNOR U6267 ( .A(b[3178]), .B(n5348), .Z(c[3178]) );
  XNOR U6268 ( .A(a[3178]), .B(n5349), .Z(n5348) );
  IV U6269 ( .A(n5346), .Z(n5349) );
  XOR U6270 ( .A(n5350), .B(n5351), .Z(n5346) );
  ANDN U6271 ( .B(n5352), .A(n5353), .Z(n5350) );
  XNOR U6272 ( .A(b[3177]), .B(n5351), .Z(n5352) );
  XNOR U6273 ( .A(b[3177]), .B(n5353), .Z(c[3177]) );
  XNOR U6274 ( .A(a[3177]), .B(n5354), .Z(n5353) );
  IV U6275 ( .A(n5351), .Z(n5354) );
  XOR U6276 ( .A(n5355), .B(n5356), .Z(n5351) );
  ANDN U6277 ( .B(n5357), .A(n5358), .Z(n5355) );
  XNOR U6278 ( .A(b[3176]), .B(n5356), .Z(n5357) );
  XNOR U6279 ( .A(b[3176]), .B(n5358), .Z(c[3176]) );
  XNOR U6280 ( .A(a[3176]), .B(n5359), .Z(n5358) );
  IV U6281 ( .A(n5356), .Z(n5359) );
  XOR U6282 ( .A(n5360), .B(n5361), .Z(n5356) );
  ANDN U6283 ( .B(n5362), .A(n5363), .Z(n5360) );
  XNOR U6284 ( .A(b[3175]), .B(n5361), .Z(n5362) );
  XNOR U6285 ( .A(b[3175]), .B(n5363), .Z(c[3175]) );
  XNOR U6286 ( .A(a[3175]), .B(n5364), .Z(n5363) );
  IV U6287 ( .A(n5361), .Z(n5364) );
  XOR U6288 ( .A(n5365), .B(n5366), .Z(n5361) );
  ANDN U6289 ( .B(n5367), .A(n5368), .Z(n5365) );
  XNOR U6290 ( .A(b[3174]), .B(n5366), .Z(n5367) );
  XNOR U6291 ( .A(b[3174]), .B(n5368), .Z(c[3174]) );
  XNOR U6292 ( .A(a[3174]), .B(n5369), .Z(n5368) );
  IV U6293 ( .A(n5366), .Z(n5369) );
  XOR U6294 ( .A(n5370), .B(n5371), .Z(n5366) );
  ANDN U6295 ( .B(n5372), .A(n5373), .Z(n5370) );
  XNOR U6296 ( .A(b[3173]), .B(n5371), .Z(n5372) );
  XNOR U6297 ( .A(b[3173]), .B(n5373), .Z(c[3173]) );
  XNOR U6298 ( .A(a[3173]), .B(n5374), .Z(n5373) );
  IV U6299 ( .A(n5371), .Z(n5374) );
  XOR U6300 ( .A(n5375), .B(n5376), .Z(n5371) );
  ANDN U6301 ( .B(n5377), .A(n5378), .Z(n5375) );
  XNOR U6302 ( .A(b[3172]), .B(n5376), .Z(n5377) );
  XNOR U6303 ( .A(b[3172]), .B(n5378), .Z(c[3172]) );
  XNOR U6304 ( .A(a[3172]), .B(n5379), .Z(n5378) );
  IV U6305 ( .A(n5376), .Z(n5379) );
  XOR U6306 ( .A(n5380), .B(n5381), .Z(n5376) );
  ANDN U6307 ( .B(n5382), .A(n5383), .Z(n5380) );
  XNOR U6308 ( .A(b[3171]), .B(n5381), .Z(n5382) );
  XNOR U6309 ( .A(b[3171]), .B(n5383), .Z(c[3171]) );
  XNOR U6310 ( .A(a[3171]), .B(n5384), .Z(n5383) );
  IV U6311 ( .A(n5381), .Z(n5384) );
  XOR U6312 ( .A(n5385), .B(n5386), .Z(n5381) );
  ANDN U6313 ( .B(n5387), .A(n5388), .Z(n5385) );
  XNOR U6314 ( .A(b[3170]), .B(n5386), .Z(n5387) );
  XNOR U6315 ( .A(b[3170]), .B(n5388), .Z(c[3170]) );
  XNOR U6316 ( .A(a[3170]), .B(n5389), .Z(n5388) );
  IV U6317 ( .A(n5386), .Z(n5389) );
  XOR U6318 ( .A(n5390), .B(n5391), .Z(n5386) );
  ANDN U6319 ( .B(n5392), .A(n5393), .Z(n5390) );
  XNOR U6320 ( .A(b[3169]), .B(n5391), .Z(n5392) );
  XNOR U6321 ( .A(b[316]), .B(n5394), .Z(c[316]) );
  XNOR U6322 ( .A(b[3169]), .B(n5393), .Z(c[3169]) );
  XNOR U6323 ( .A(a[3169]), .B(n5395), .Z(n5393) );
  IV U6324 ( .A(n5391), .Z(n5395) );
  XOR U6325 ( .A(n5396), .B(n5397), .Z(n5391) );
  ANDN U6326 ( .B(n5398), .A(n5399), .Z(n5396) );
  XNOR U6327 ( .A(b[3168]), .B(n5397), .Z(n5398) );
  XNOR U6328 ( .A(b[3168]), .B(n5399), .Z(c[3168]) );
  XNOR U6329 ( .A(a[3168]), .B(n5400), .Z(n5399) );
  IV U6330 ( .A(n5397), .Z(n5400) );
  XOR U6331 ( .A(n5401), .B(n5402), .Z(n5397) );
  ANDN U6332 ( .B(n5403), .A(n5404), .Z(n5401) );
  XNOR U6333 ( .A(b[3167]), .B(n5402), .Z(n5403) );
  XNOR U6334 ( .A(b[3167]), .B(n5404), .Z(c[3167]) );
  XNOR U6335 ( .A(a[3167]), .B(n5405), .Z(n5404) );
  IV U6336 ( .A(n5402), .Z(n5405) );
  XOR U6337 ( .A(n5406), .B(n5407), .Z(n5402) );
  ANDN U6338 ( .B(n5408), .A(n5409), .Z(n5406) );
  XNOR U6339 ( .A(b[3166]), .B(n5407), .Z(n5408) );
  XNOR U6340 ( .A(b[3166]), .B(n5409), .Z(c[3166]) );
  XNOR U6341 ( .A(a[3166]), .B(n5410), .Z(n5409) );
  IV U6342 ( .A(n5407), .Z(n5410) );
  XOR U6343 ( .A(n5411), .B(n5412), .Z(n5407) );
  ANDN U6344 ( .B(n5413), .A(n5414), .Z(n5411) );
  XNOR U6345 ( .A(b[3165]), .B(n5412), .Z(n5413) );
  XNOR U6346 ( .A(b[3165]), .B(n5414), .Z(c[3165]) );
  XNOR U6347 ( .A(a[3165]), .B(n5415), .Z(n5414) );
  IV U6348 ( .A(n5412), .Z(n5415) );
  XOR U6349 ( .A(n5416), .B(n5417), .Z(n5412) );
  ANDN U6350 ( .B(n5418), .A(n5419), .Z(n5416) );
  XNOR U6351 ( .A(b[3164]), .B(n5417), .Z(n5418) );
  XNOR U6352 ( .A(b[3164]), .B(n5419), .Z(c[3164]) );
  XNOR U6353 ( .A(a[3164]), .B(n5420), .Z(n5419) );
  IV U6354 ( .A(n5417), .Z(n5420) );
  XOR U6355 ( .A(n5421), .B(n5422), .Z(n5417) );
  ANDN U6356 ( .B(n5423), .A(n5424), .Z(n5421) );
  XNOR U6357 ( .A(b[3163]), .B(n5422), .Z(n5423) );
  XNOR U6358 ( .A(b[3163]), .B(n5424), .Z(c[3163]) );
  XNOR U6359 ( .A(a[3163]), .B(n5425), .Z(n5424) );
  IV U6360 ( .A(n5422), .Z(n5425) );
  XOR U6361 ( .A(n5426), .B(n5427), .Z(n5422) );
  ANDN U6362 ( .B(n5428), .A(n5429), .Z(n5426) );
  XNOR U6363 ( .A(b[3162]), .B(n5427), .Z(n5428) );
  XNOR U6364 ( .A(b[3162]), .B(n5429), .Z(c[3162]) );
  XNOR U6365 ( .A(a[3162]), .B(n5430), .Z(n5429) );
  IV U6366 ( .A(n5427), .Z(n5430) );
  XOR U6367 ( .A(n5431), .B(n5432), .Z(n5427) );
  ANDN U6368 ( .B(n5433), .A(n5434), .Z(n5431) );
  XNOR U6369 ( .A(b[3161]), .B(n5432), .Z(n5433) );
  XNOR U6370 ( .A(b[3161]), .B(n5434), .Z(c[3161]) );
  XNOR U6371 ( .A(a[3161]), .B(n5435), .Z(n5434) );
  IV U6372 ( .A(n5432), .Z(n5435) );
  XOR U6373 ( .A(n5436), .B(n5437), .Z(n5432) );
  ANDN U6374 ( .B(n5438), .A(n5439), .Z(n5436) );
  XNOR U6375 ( .A(b[3160]), .B(n5437), .Z(n5438) );
  XNOR U6376 ( .A(b[3160]), .B(n5439), .Z(c[3160]) );
  XNOR U6377 ( .A(a[3160]), .B(n5440), .Z(n5439) );
  IV U6378 ( .A(n5437), .Z(n5440) );
  XOR U6379 ( .A(n5441), .B(n5442), .Z(n5437) );
  ANDN U6380 ( .B(n5443), .A(n5444), .Z(n5441) );
  XNOR U6381 ( .A(b[3159]), .B(n5442), .Z(n5443) );
  XNOR U6382 ( .A(b[315]), .B(n5445), .Z(c[315]) );
  XNOR U6383 ( .A(b[3159]), .B(n5444), .Z(c[3159]) );
  XNOR U6384 ( .A(a[3159]), .B(n5446), .Z(n5444) );
  IV U6385 ( .A(n5442), .Z(n5446) );
  XOR U6386 ( .A(n5447), .B(n5448), .Z(n5442) );
  ANDN U6387 ( .B(n5449), .A(n5450), .Z(n5447) );
  XNOR U6388 ( .A(b[3158]), .B(n5448), .Z(n5449) );
  XNOR U6389 ( .A(b[3158]), .B(n5450), .Z(c[3158]) );
  XNOR U6390 ( .A(a[3158]), .B(n5451), .Z(n5450) );
  IV U6391 ( .A(n5448), .Z(n5451) );
  XOR U6392 ( .A(n5452), .B(n5453), .Z(n5448) );
  ANDN U6393 ( .B(n5454), .A(n5455), .Z(n5452) );
  XNOR U6394 ( .A(b[3157]), .B(n5453), .Z(n5454) );
  XNOR U6395 ( .A(b[3157]), .B(n5455), .Z(c[3157]) );
  XNOR U6396 ( .A(a[3157]), .B(n5456), .Z(n5455) );
  IV U6397 ( .A(n5453), .Z(n5456) );
  XOR U6398 ( .A(n5457), .B(n5458), .Z(n5453) );
  ANDN U6399 ( .B(n5459), .A(n5460), .Z(n5457) );
  XNOR U6400 ( .A(b[3156]), .B(n5458), .Z(n5459) );
  XNOR U6401 ( .A(b[3156]), .B(n5460), .Z(c[3156]) );
  XNOR U6402 ( .A(a[3156]), .B(n5461), .Z(n5460) );
  IV U6403 ( .A(n5458), .Z(n5461) );
  XOR U6404 ( .A(n5462), .B(n5463), .Z(n5458) );
  ANDN U6405 ( .B(n5464), .A(n5465), .Z(n5462) );
  XNOR U6406 ( .A(b[3155]), .B(n5463), .Z(n5464) );
  XNOR U6407 ( .A(b[3155]), .B(n5465), .Z(c[3155]) );
  XNOR U6408 ( .A(a[3155]), .B(n5466), .Z(n5465) );
  IV U6409 ( .A(n5463), .Z(n5466) );
  XOR U6410 ( .A(n5467), .B(n5468), .Z(n5463) );
  ANDN U6411 ( .B(n5469), .A(n5470), .Z(n5467) );
  XNOR U6412 ( .A(b[3154]), .B(n5468), .Z(n5469) );
  XNOR U6413 ( .A(b[3154]), .B(n5470), .Z(c[3154]) );
  XNOR U6414 ( .A(a[3154]), .B(n5471), .Z(n5470) );
  IV U6415 ( .A(n5468), .Z(n5471) );
  XOR U6416 ( .A(n5472), .B(n5473), .Z(n5468) );
  ANDN U6417 ( .B(n5474), .A(n5475), .Z(n5472) );
  XNOR U6418 ( .A(b[3153]), .B(n5473), .Z(n5474) );
  XNOR U6419 ( .A(b[3153]), .B(n5475), .Z(c[3153]) );
  XNOR U6420 ( .A(a[3153]), .B(n5476), .Z(n5475) );
  IV U6421 ( .A(n5473), .Z(n5476) );
  XOR U6422 ( .A(n5477), .B(n5478), .Z(n5473) );
  ANDN U6423 ( .B(n5479), .A(n5480), .Z(n5477) );
  XNOR U6424 ( .A(b[3152]), .B(n5478), .Z(n5479) );
  XNOR U6425 ( .A(b[3152]), .B(n5480), .Z(c[3152]) );
  XNOR U6426 ( .A(a[3152]), .B(n5481), .Z(n5480) );
  IV U6427 ( .A(n5478), .Z(n5481) );
  XOR U6428 ( .A(n5482), .B(n5483), .Z(n5478) );
  ANDN U6429 ( .B(n5484), .A(n5485), .Z(n5482) );
  XNOR U6430 ( .A(b[3151]), .B(n5483), .Z(n5484) );
  XNOR U6431 ( .A(b[3151]), .B(n5485), .Z(c[3151]) );
  XNOR U6432 ( .A(a[3151]), .B(n5486), .Z(n5485) );
  IV U6433 ( .A(n5483), .Z(n5486) );
  XOR U6434 ( .A(n5487), .B(n5488), .Z(n5483) );
  ANDN U6435 ( .B(n5489), .A(n5490), .Z(n5487) );
  XNOR U6436 ( .A(b[3150]), .B(n5488), .Z(n5489) );
  XNOR U6437 ( .A(b[3150]), .B(n5490), .Z(c[3150]) );
  XNOR U6438 ( .A(a[3150]), .B(n5491), .Z(n5490) );
  IV U6439 ( .A(n5488), .Z(n5491) );
  XOR U6440 ( .A(n5492), .B(n5493), .Z(n5488) );
  ANDN U6441 ( .B(n5494), .A(n5495), .Z(n5492) );
  XNOR U6442 ( .A(b[3149]), .B(n5493), .Z(n5494) );
  XNOR U6443 ( .A(b[314]), .B(n5496), .Z(c[314]) );
  XNOR U6444 ( .A(b[3149]), .B(n5495), .Z(c[3149]) );
  XNOR U6445 ( .A(a[3149]), .B(n5497), .Z(n5495) );
  IV U6446 ( .A(n5493), .Z(n5497) );
  XOR U6447 ( .A(n5498), .B(n5499), .Z(n5493) );
  ANDN U6448 ( .B(n5500), .A(n5501), .Z(n5498) );
  XNOR U6449 ( .A(b[3148]), .B(n5499), .Z(n5500) );
  XNOR U6450 ( .A(b[3148]), .B(n5501), .Z(c[3148]) );
  XNOR U6451 ( .A(a[3148]), .B(n5502), .Z(n5501) );
  IV U6452 ( .A(n5499), .Z(n5502) );
  XOR U6453 ( .A(n5503), .B(n5504), .Z(n5499) );
  ANDN U6454 ( .B(n5505), .A(n5506), .Z(n5503) );
  XNOR U6455 ( .A(b[3147]), .B(n5504), .Z(n5505) );
  XNOR U6456 ( .A(b[3147]), .B(n5506), .Z(c[3147]) );
  XNOR U6457 ( .A(a[3147]), .B(n5507), .Z(n5506) );
  IV U6458 ( .A(n5504), .Z(n5507) );
  XOR U6459 ( .A(n5508), .B(n5509), .Z(n5504) );
  ANDN U6460 ( .B(n5510), .A(n5511), .Z(n5508) );
  XNOR U6461 ( .A(b[3146]), .B(n5509), .Z(n5510) );
  XNOR U6462 ( .A(b[3146]), .B(n5511), .Z(c[3146]) );
  XNOR U6463 ( .A(a[3146]), .B(n5512), .Z(n5511) );
  IV U6464 ( .A(n5509), .Z(n5512) );
  XOR U6465 ( .A(n5513), .B(n5514), .Z(n5509) );
  ANDN U6466 ( .B(n5515), .A(n5516), .Z(n5513) );
  XNOR U6467 ( .A(b[3145]), .B(n5514), .Z(n5515) );
  XNOR U6468 ( .A(b[3145]), .B(n5516), .Z(c[3145]) );
  XNOR U6469 ( .A(a[3145]), .B(n5517), .Z(n5516) );
  IV U6470 ( .A(n5514), .Z(n5517) );
  XOR U6471 ( .A(n5518), .B(n5519), .Z(n5514) );
  ANDN U6472 ( .B(n5520), .A(n5521), .Z(n5518) );
  XNOR U6473 ( .A(b[3144]), .B(n5519), .Z(n5520) );
  XNOR U6474 ( .A(b[3144]), .B(n5521), .Z(c[3144]) );
  XNOR U6475 ( .A(a[3144]), .B(n5522), .Z(n5521) );
  IV U6476 ( .A(n5519), .Z(n5522) );
  XOR U6477 ( .A(n5523), .B(n5524), .Z(n5519) );
  ANDN U6478 ( .B(n5525), .A(n5526), .Z(n5523) );
  XNOR U6479 ( .A(b[3143]), .B(n5524), .Z(n5525) );
  XNOR U6480 ( .A(b[3143]), .B(n5526), .Z(c[3143]) );
  XNOR U6481 ( .A(a[3143]), .B(n5527), .Z(n5526) );
  IV U6482 ( .A(n5524), .Z(n5527) );
  XOR U6483 ( .A(n5528), .B(n5529), .Z(n5524) );
  ANDN U6484 ( .B(n5530), .A(n5531), .Z(n5528) );
  XNOR U6485 ( .A(b[3142]), .B(n5529), .Z(n5530) );
  XNOR U6486 ( .A(b[3142]), .B(n5531), .Z(c[3142]) );
  XNOR U6487 ( .A(a[3142]), .B(n5532), .Z(n5531) );
  IV U6488 ( .A(n5529), .Z(n5532) );
  XOR U6489 ( .A(n5533), .B(n5534), .Z(n5529) );
  ANDN U6490 ( .B(n5535), .A(n5536), .Z(n5533) );
  XNOR U6491 ( .A(b[3141]), .B(n5534), .Z(n5535) );
  XNOR U6492 ( .A(b[3141]), .B(n5536), .Z(c[3141]) );
  XNOR U6493 ( .A(a[3141]), .B(n5537), .Z(n5536) );
  IV U6494 ( .A(n5534), .Z(n5537) );
  XOR U6495 ( .A(n5538), .B(n5539), .Z(n5534) );
  ANDN U6496 ( .B(n5540), .A(n5541), .Z(n5538) );
  XNOR U6497 ( .A(b[3140]), .B(n5539), .Z(n5540) );
  XNOR U6498 ( .A(b[3140]), .B(n5541), .Z(c[3140]) );
  XNOR U6499 ( .A(a[3140]), .B(n5542), .Z(n5541) );
  IV U6500 ( .A(n5539), .Z(n5542) );
  XOR U6501 ( .A(n5543), .B(n5544), .Z(n5539) );
  ANDN U6502 ( .B(n5545), .A(n5546), .Z(n5543) );
  XNOR U6503 ( .A(b[3139]), .B(n5544), .Z(n5545) );
  XNOR U6504 ( .A(b[313]), .B(n5547), .Z(c[313]) );
  XNOR U6505 ( .A(b[3139]), .B(n5546), .Z(c[3139]) );
  XNOR U6506 ( .A(a[3139]), .B(n5548), .Z(n5546) );
  IV U6507 ( .A(n5544), .Z(n5548) );
  XOR U6508 ( .A(n5549), .B(n5550), .Z(n5544) );
  ANDN U6509 ( .B(n5551), .A(n5552), .Z(n5549) );
  XNOR U6510 ( .A(b[3138]), .B(n5550), .Z(n5551) );
  XNOR U6511 ( .A(b[3138]), .B(n5552), .Z(c[3138]) );
  XNOR U6512 ( .A(a[3138]), .B(n5553), .Z(n5552) );
  IV U6513 ( .A(n5550), .Z(n5553) );
  XOR U6514 ( .A(n5554), .B(n5555), .Z(n5550) );
  ANDN U6515 ( .B(n5556), .A(n5557), .Z(n5554) );
  XNOR U6516 ( .A(b[3137]), .B(n5555), .Z(n5556) );
  XNOR U6517 ( .A(b[3137]), .B(n5557), .Z(c[3137]) );
  XNOR U6518 ( .A(a[3137]), .B(n5558), .Z(n5557) );
  IV U6519 ( .A(n5555), .Z(n5558) );
  XOR U6520 ( .A(n5559), .B(n5560), .Z(n5555) );
  ANDN U6521 ( .B(n5561), .A(n5562), .Z(n5559) );
  XNOR U6522 ( .A(b[3136]), .B(n5560), .Z(n5561) );
  XNOR U6523 ( .A(b[3136]), .B(n5562), .Z(c[3136]) );
  XNOR U6524 ( .A(a[3136]), .B(n5563), .Z(n5562) );
  IV U6525 ( .A(n5560), .Z(n5563) );
  XOR U6526 ( .A(n5564), .B(n5565), .Z(n5560) );
  ANDN U6527 ( .B(n5566), .A(n5567), .Z(n5564) );
  XNOR U6528 ( .A(b[3135]), .B(n5565), .Z(n5566) );
  XNOR U6529 ( .A(b[3135]), .B(n5567), .Z(c[3135]) );
  XNOR U6530 ( .A(a[3135]), .B(n5568), .Z(n5567) );
  IV U6531 ( .A(n5565), .Z(n5568) );
  XOR U6532 ( .A(n5569), .B(n5570), .Z(n5565) );
  ANDN U6533 ( .B(n5571), .A(n5572), .Z(n5569) );
  XNOR U6534 ( .A(b[3134]), .B(n5570), .Z(n5571) );
  XNOR U6535 ( .A(b[3134]), .B(n5572), .Z(c[3134]) );
  XNOR U6536 ( .A(a[3134]), .B(n5573), .Z(n5572) );
  IV U6537 ( .A(n5570), .Z(n5573) );
  XOR U6538 ( .A(n5574), .B(n5575), .Z(n5570) );
  ANDN U6539 ( .B(n5576), .A(n5577), .Z(n5574) );
  XNOR U6540 ( .A(b[3133]), .B(n5575), .Z(n5576) );
  XNOR U6541 ( .A(b[3133]), .B(n5577), .Z(c[3133]) );
  XNOR U6542 ( .A(a[3133]), .B(n5578), .Z(n5577) );
  IV U6543 ( .A(n5575), .Z(n5578) );
  XOR U6544 ( .A(n5579), .B(n5580), .Z(n5575) );
  ANDN U6545 ( .B(n5581), .A(n5582), .Z(n5579) );
  XNOR U6546 ( .A(b[3132]), .B(n5580), .Z(n5581) );
  XNOR U6547 ( .A(b[3132]), .B(n5582), .Z(c[3132]) );
  XNOR U6548 ( .A(a[3132]), .B(n5583), .Z(n5582) );
  IV U6549 ( .A(n5580), .Z(n5583) );
  XOR U6550 ( .A(n5584), .B(n5585), .Z(n5580) );
  ANDN U6551 ( .B(n5586), .A(n5587), .Z(n5584) );
  XNOR U6552 ( .A(b[3131]), .B(n5585), .Z(n5586) );
  XNOR U6553 ( .A(b[3131]), .B(n5587), .Z(c[3131]) );
  XNOR U6554 ( .A(a[3131]), .B(n5588), .Z(n5587) );
  IV U6555 ( .A(n5585), .Z(n5588) );
  XOR U6556 ( .A(n5589), .B(n5590), .Z(n5585) );
  ANDN U6557 ( .B(n5591), .A(n5592), .Z(n5589) );
  XNOR U6558 ( .A(b[3130]), .B(n5590), .Z(n5591) );
  XNOR U6559 ( .A(b[3130]), .B(n5592), .Z(c[3130]) );
  XNOR U6560 ( .A(a[3130]), .B(n5593), .Z(n5592) );
  IV U6561 ( .A(n5590), .Z(n5593) );
  XOR U6562 ( .A(n5594), .B(n5595), .Z(n5590) );
  ANDN U6563 ( .B(n5596), .A(n5597), .Z(n5594) );
  XNOR U6564 ( .A(b[3129]), .B(n5595), .Z(n5596) );
  XNOR U6565 ( .A(b[312]), .B(n5598), .Z(c[312]) );
  XNOR U6566 ( .A(b[3129]), .B(n5597), .Z(c[3129]) );
  XNOR U6567 ( .A(a[3129]), .B(n5599), .Z(n5597) );
  IV U6568 ( .A(n5595), .Z(n5599) );
  XOR U6569 ( .A(n5600), .B(n5601), .Z(n5595) );
  ANDN U6570 ( .B(n5602), .A(n5603), .Z(n5600) );
  XNOR U6571 ( .A(b[3128]), .B(n5601), .Z(n5602) );
  XNOR U6572 ( .A(b[3128]), .B(n5603), .Z(c[3128]) );
  XNOR U6573 ( .A(a[3128]), .B(n5604), .Z(n5603) );
  IV U6574 ( .A(n5601), .Z(n5604) );
  XOR U6575 ( .A(n5605), .B(n5606), .Z(n5601) );
  ANDN U6576 ( .B(n5607), .A(n5608), .Z(n5605) );
  XNOR U6577 ( .A(b[3127]), .B(n5606), .Z(n5607) );
  XNOR U6578 ( .A(b[3127]), .B(n5608), .Z(c[3127]) );
  XNOR U6579 ( .A(a[3127]), .B(n5609), .Z(n5608) );
  IV U6580 ( .A(n5606), .Z(n5609) );
  XOR U6581 ( .A(n5610), .B(n5611), .Z(n5606) );
  ANDN U6582 ( .B(n5612), .A(n5613), .Z(n5610) );
  XNOR U6583 ( .A(b[3126]), .B(n5611), .Z(n5612) );
  XNOR U6584 ( .A(b[3126]), .B(n5613), .Z(c[3126]) );
  XNOR U6585 ( .A(a[3126]), .B(n5614), .Z(n5613) );
  IV U6586 ( .A(n5611), .Z(n5614) );
  XOR U6587 ( .A(n5615), .B(n5616), .Z(n5611) );
  ANDN U6588 ( .B(n5617), .A(n5618), .Z(n5615) );
  XNOR U6589 ( .A(b[3125]), .B(n5616), .Z(n5617) );
  XNOR U6590 ( .A(b[3125]), .B(n5618), .Z(c[3125]) );
  XNOR U6591 ( .A(a[3125]), .B(n5619), .Z(n5618) );
  IV U6592 ( .A(n5616), .Z(n5619) );
  XOR U6593 ( .A(n5620), .B(n5621), .Z(n5616) );
  ANDN U6594 ( .B(n5622), .A(n5623), .Z(n5620) );
  XNOR U6595 ( .A(b[3124]), .B(n5621), .Z(n5622) );
  XNOR U6596 ( .A(b[3124]), .B(n5623), .Z(c[3124]) );
  XNOR U6597 ( .A(a[3124]), .B(n5624), .Z(n5623) );
  IV U6598 ( .A(n5621), .Z(n5624) );
  XOR U6599 ( .A(n5625), .B(n5626), .Z(n5621) );
  ANDN U6600 ( .B(n5627), .A(n5628), .Z(n5625) );
  XNOR U6601 ( .A(b[3123]), .B(n5626), .Z(n5627) );
  XNOR U6602 ( .A(b[3123]), .B(n5628), .Z(c[3123]) );
  XNOR U6603 ( .A(a[3123]), .B(n5629), .Z(n5628) );
  IV U6604 ( .A(n5626), .Z(n5629) );
  XOR U6605 ( .A(n5630), .B(n5631), .Z(n5626) );
  ANDN U6606 ( .B(n5632), .A(n5633), .Z(n5630) );
  XNOR U6607 ( .A(b[3122]), .B(n5631), .Z(n5632) );
  XNOR U6608 ( .A(b[3122]), .B(n5633), .Z(c[3122]) );
  XNOR U6609 ( .A(a[3122]), .B(n5634), .Z(n5633) );
  IV U6610 ( .A(n5631), .Z(n5634) );
  XOR U6611 ( .A(n5635), .B(n5636), .Z(n5631) );
  ANDN U6612 ( .B(n5637), .A(n5638), .Z(n5635) );
  XNOR U6613 ( .A(b[3121]), .B(n5636), .Z(n5637) );
  XNOR U6614 ( .A(b[3121]), .B(n5638), .Z(c[3121]) );
  XNOR U6615 ( .A(a[3121]), .B(n5639), .Z(n5638) );
  IV U6616 ( .A(n5636), .Z(n5639) );
  XOR U6617 ( .A(n5640), .B(n5641), .Z(n5636) );
  ANDN U6618 ( .B(n5642), .A(n5643), .Z(n5640) );
  XNOR U6619 ( .A(b[3120]), .B(n5641), .Z(n5642) );
  XNOR U6620 ( .A(b[3120]), .B(n5643), .Z(c[3120]) );
  XNOR U6621 ( .A(a[3120]), .B(n5644), .Z(n5643) );
  IV U6622 ( .A(n5641), .Z(n5644) );
  XOR U6623 ( .A(n5645), .B(n5646), .Z(n5641) );
  ANDN U6624 ( .B(n5647), .A(n5648), .Z(n5645) );
  XNOR U6625 ( .A(b[3119]), .B(n5646), .Z(n5647) );
  XNOR U6626 ( .A(b[311]), .B(n5649), .Z(c[311]) );
  XNOR U6627 ( .A(b[3119]), .B(n5648), .Z(c[3119]) );
  XNOR U6628 ( .A(a[3119]), .B(n5650), .Z(n5648) );
  IV U6629 ( .A(n5646), .Z(n5650) );
  XOR U6630 ( .A(n5651), .B(n5652), .Z(n5646) );
  ANDN U6631 ( .B(n5653), .A(n5654), .Z(n5651) );
  XNOR U6632 ( .A(b[3118]), .B(n5652), .Z(n5653) );
  XNOR U6633 ( .A(b[3118]), .B(n5654), .Z(c[3118]) );
  XNOR U6634 ( .A(a[3118]), .B(n5655), .Z(n5654) );
  IV U6635 ( .A(n5652), .Z(n5655) );
  XOR U6636 ( .A(n5656), .B(n5657), .Z(n5652) );
  ANDN U6637 ( .B(n5658), .A(n5659), .Z(n5656) );
  XNOR U6638 ( .A(b[3117]), .B(n5657), .Z(n5658) );
  XNOR U6639 ( .A(b[3117]), .B(n5659), .Z(c[3117]) );
  XNOR U6640 ( .A(a[3117]), .B(n5660), .Z(n5659) );
  IV U6641 ( .A(n5657), .Z(n5660) );
  XOR U6642 ( .A(n5661), .B(n5662), .Z(n5657) );
  ANDN U6643 ( .B(n5663), .A(n5664), .Z(n5661) );
  XNOR U6644 ( .A(b[3116]), .B(n5662), .Z(n5663) );
  XNOR U6645 ( .A(b[3116]), .B(n5664), .Z(c[3116]) );
  XNOR U6646 ( .A(a[3116]), .B(n5665), .Z(n5664) );
  IV U6647 ( .A(n5662), .Z(n5665) );
  XOR U6648 ( .A(n5666), .B(n5667), .Z(n5662) );
  ANDN U6649 ( .B(n5668), .A(n5669), .Z(n5666) );
  XNOR U6650 ( .A(b[3115]), .B(n5667), .Z(n5668) );
  XNOR U6651 ( .A(b[3115]), .B(n5669), .Z(c[3115]) );
  XNOR U6652 ( .A(a[3115]), .B(n5670), .Z(n5669) );
  IV U6653 ( .A(n5667), .Z(n5670) );
  XOR U6654 ( .A(n5671), .B(n5672), .Z(n5667) );
  ANDN U6655 ( .B(n5673), .A(n5674), .Z(n5671) );
  XNOR U6656 ( .A(b[3114]), .B(n5672), .Z(n5673) );
  XNOR U6657 ( .A(b[3114]), .B(n5674), .Z(c[3114]) );
  XNOR U6658 ( .A(a[3114]), .B(n5675), .Z(n5674) );
  IV U6659 ( .A(n5672), .Z(n5675) );
  XOR U6660 ( .A(n5676), .B(n5677), .Z(n5672) );
  ANDN U6661 ( .B(n5678), .A(n5679), .Z(n5676) );
  XNOR U6662 ( .A(b[3113]), .B(n5677), .Z(n5678) );
  XNOR U6663 ( .A(b[3113]), .B(n5679), .Z(c[3113]) );
  XNOR U6664 ( .A(a[3113]), .B(n5680), .Z(n5679) );
  IV U6665 ( .A(n5677), .Z(n5680) );
  XOR U6666 ( .A(n5681), .B(n5682), .Z(n5677) );
  ANDN U6667 ( .B(n5683), .A(n5684), .Z(n5681) );
  XNOR U6668 ( .A(b[3112]), .B(n5682), .Z(n5683) );
  XNOR U6669 ( .A(b[3112]), .B(n5684), .Z(c[3112]) );
  XNOR U6670 ( .A(a[3112]), .B(n5685), .Z(n5684) );
  IV U6671 ( .A(n5682), .Z(n5685) );
  XOR U6672 ( .A(n5686), .B(n5687), .Z(n5682) );
  ANDN U6673 ( .B(n5688), .A(n5689), .Z(n5686) );
  XNOR U6674 ( .A(b[3111]), .B(n5687), .Z(n5688) );
  XNOR U6675 ( .A(b[3111]), .B(n5689), .Z(c[3111]) );
  XNOR U6676 ( .A(a[3111]), .B(n5690), .Z(n5689) );
  IV U6677 ( .A(n5687), .Z(n5690) );
  XOR U6678 ( .A(n5691), .B(n5692), .Z(n5687) );
  ANDN U6679 ( .B(n5693), .A(n5694), .Z(n5691) );
  XNOR U6680 ( .A(b[3110]), .B(n5692), .Z(n5693) );
  XNOR U6681 ( .A(b[3110]), .B(n5694), .Z(c[3110]) );
  XNOR U6682 ( .A(a[3110]), .B(n5695), .Z(n5694) );
  IV U6683 ( .A(n5692), .Z(n5695) );
  XOR U6684 ( .A(n5696), .B(n5697), .Z(n5692) );
  ANDN U6685 ( .B(n5698), .A(n5699), .Z(n5696) );
  XNOR U6686 ( .A(b[3109]), .B(n5697), .Z(n5698) );
  XNOR U6687 ( .A(b[310]), .B(n5700), .Z(c[310]) );
  XNOR U6688 ( .A(b[3109]), .B(n5699), .Z(c[3109]) );
  XNOR U6689 ( .A(a[3109]), .B(n5701), .Z(n5699) );
  IV U6690 ( .A(n5697), .Z(n5701) );
  XOR U6691 ( .A(n5702), .B(n5703), .Z(n5697) );
  ANDN U6692 ( .B(n5704), .A(n5705), .Z(n5702) );
  XNOR U6693 ( .A(b[3108]), .B(n5703), .Z(n5704) );
  XNOR U6694 ( .A(b[3108]), .B(n5705), .Z(c[3108]) );
  XNOR U6695 ( .A(a[3108]), .B(n5706), .Z(n5705) );
  IV U6696 ( .A(n5703), .Z(n5706) );
  XOR U6697 ( .A(n5707), .B(n5708), .Z(n5703) );
  ANDN U6698 ( .B(n5709), .A(n5710), .Z(n5707) );
  XNOR U6699 ( .A(b[3107]), .B(n5708), .Z(n5709) );
  XNOR U6700 ( .A(b[3107]), .B(n5710), .Z(c[3107]) );
  XNOR U6701 ( .A(a[3107]), .B(n5711), .Z(n5710) );
  IV U6702 ( .A(n5708), .Z(n5711) );
  XOR U6703 ( .A(n5712), .B(n5713), .Z(n5708) );
  ANDN U6704 ( .B(n5714), .A(n5715), .Z(n5712) );
  XNOR U6705 ( .A(b[3106]), .B(n5713), .Z(n5714) );
  XNOR U6706 ( .A(b[3106]), .B(n5715), .Z(c[3106]) );
  XNOR U6707 ( .A(a[3106]), .B(n5716), .Z(n5715) );
  IV U6708 ( .A(n5713), .Z(n5716) );
  XOR U6709 ( .A(n5717), .B(n5718), .Z(n5713) );
  ANDN U6710 ( .B(n5719), .A(n5720), .Z(n5717) );
  XNOR U6711 ( .A(b[3105]), .B(n5718), .Z(n5719) );
  XNOR U6712 ( .A(b[3105]), .B(n5720), .Z(c[3105]) );
  XNOR U6713 ( .A(a[3105]), .B(n5721), .Z(n5720) );
  IV U6714 ( .A(n5718), .Z(n5721) );
  XOR U6715 ( .A(n5722), .B(n5723), .Z(n5718) );
  ANDN U6716 ( .B(n5724), .A(n5725), .Z(n5722) );
  XNOR U6717 ( .A(b[3104]), .B(n5723), .Z(n5724) );
  XNOR U6718 ( .A(b[3104]), .B(n5725), .Z(c[3104]) );
  XNOR U6719 ( .A(a[3104]), .B(n5726), .Z(n5725) );
  IV U6720 ( .A(n5723), .Z(n5726) );
  XOR U6721 ( .A(n5727), .B(n5728), .Z(n5723) );
  ANDN U6722 ( .B(n5729), .A(n5730), .Z(n5727) );
  XNOR U6723 ( .A(b[3103]), .B(n5728), .Z(n5729) );
  XNOR U6724 ( .A(b[3103]), .B(n5730), .Z(c[3103]) );
  XNOR U6725 ( .A(a[3103]), .B(n5731), .Z(n5730) );
  IV U6726 ( .A(n5728), .Z(n5731) );
  XOR U6727 ( .A(n5732), .B(n5733), .Z(n5728) );
  ANDN U6728 ( .B(n5734), .A(n5735), .Z(n5732) );
  XNOR U6729 ( .A(b[3102]), .B(n5733), .Z(n5734) );
  XNOR U6730 ( .A(b[3102]), .B(n5735), .Z(c[3102]) );
  XNOR U6731 ( .A(a[3102]), .B(n5736), .Z(n5735) );
  IV U6732 ( .A(n5733), .Z(n5736) );
  XOR U6733 ( .A(n5737), .B(n5738), .Z(n5733) );
  ANDN U6734 ( .B(n5739), .A(n5740), .Z(n5737) );
  XNOR U6735 ( .A(b[3101]), .B(n5738), .Z(n5739) );
  XNOR U6736 ( .A(b[3101]), .B(n5740), .Z(c[3101]) );
  XNOR U6737 ( .A(a[3101]), .B(n5741), .Z(n5740) );
  IV U6738 ( .A(n5738), .Z(n5741) );
  XOR U6739 ( .A(n5742), .B(n5743), .Z(n5738) );
  ANDN U6740 ( .B(n5744), .A(n5745), .Z(n5742) );
  XNOR U6741 ( .A(b[3100]), .B(n5743), .Z(n5744) );
  XNOR U6742 ( .A(b[3100]), .B(n5745), .Z(c[3100]) );
  XNOR U6743 ( .A(a[3100]), .B(n5746), .Z(n5745) );
  IV U6744 ( .A(n5743), .Z(n5746) );
  XOR U6745 ( .A(n5747), .B(n5748), .Z(n5743) );
  ANDN U6746 ( .B(n5749), .A(n5750), .Z(n5747) );
  XNOR U6747 ( .A(b[3099]), .B(n5748), .Z(n5749) );
  XNOR U6748 ( .A(b[30]), .B(n5751), .Z(c[30]) );
  XNOR U6749 ( .A(b[309]), .B(n5752), .Z(c[309]) );
  XNOR U6750 ( .A(b[3099]), .B(n5750), .Z(c[3099]) );
  XNOR U6751 ( .A(a[3099]), .B(n5753), .Z(n5750) );
  IV U6752 ( .A(n5748), .Z(n5753) );
  XOR U6753 ( .A(n5754), .B(n5755), .Z(n5748) );
  ANDN U6754 ( .B(n5756), .A(n5757), .Z(n5754) );
  XNOR U6755 ( .A(b[3098]), .B(n5755), .Z(n5756) );
  XNOR U6756 ( .A(b[3098]), .B(n5757), .Z(c[3098]) );
  XNOR U6757 ( .A(a[3098]), .B(n5758), .Z(n5757) );
  IV U6758 ( .A(n5755), .Z(n5758) );
  XOR U6759 ( .A(n5759), .B(n5760), .Z(n5755) );
  ANDN U6760 ( .B(n5761), .A(n5762), .Z(n5759) );
  XNOR U6761 ( .A(b[3097]), .B(n5760), .Z(n5761) );
  XNOR U6762 ( .A(b[3097]), .B(n5762), .Z(c[3097]) );
  XNOR U6763 ( .A(a[3097]), .B(n5763), .Z(n5762) );
  IV U6764 ( .A(n5760), .Z(n5763) );
  XOR U6765 ( .A(n5764), .B(n5765), .Z(n5760) );
  ANDN U6766 ( .B(n5766), .A(n5767), .Z(n5764) );
  XNOR U6767 ( .A(b[3096]), .B(n5765), .Z(n5766) );
  XNOR U6768 ( .A(b[3096]), .B(n5767), .Z(c[3096]) );
  XNOR U6769 ( .A(a[3096]), .B(n5768), .Z(n5767) );
  IV U6770 ( .A(n5765), .Z(n5768) );
  XOR U6771 ( .A(n5769), .B(n5770), .Z(n5765) );
  ANDN U6772 ( .B(n5771), .A(n5772), .Z(n5769) );
  XNOR U6773 ( .A(b[3095]), .B(n5770), .Z(n5771) );
  XNOR U6774 ( .A(b[3095]), .B(n5772), .Z(c[3095]) );
  XNOR U6775 ( .A(a[3095]), .B(n5773), .Z(n5772) );
  IV U6776 ( .A(n5770), .Z(n5773) );
  XOR U6777 ( .A(n5774), .B(n5775), .Z(n5770) );
  ANDN U6778 ( .B(n5776), .A(n5777), .Z(n5774) );
  XNOR U6779 ( .A(b[3094]), .B(n5775), .Z(n5776) );
  XNOR U6780 ( .A(b[3094]), .B(n5777), .Z(c[3094]) );
  XNOR U6781 ( .A(a[3094]), .B(n5778), .Z(n5777) );
  IV U6782 ( .A(n5775), .Z(n5778) );
  XOR U6783 ( .A(n5779), .B(n5780), .Z(n5775) );
  ANDN U6784 ( .B(n5781), .A(n5782), .Z(n5779) );
  XNOR U6785 ( .A(b[3093]), .B(n5780), .Z(n5781) );
  XNOR U6786 ( .A(b[3093]), .B(n5782), .Z(c[3093]) );
  XNOR U6787 ( .A(a[3093]), .B(n5783), .Z(n5782) );
  IV U6788 ( .A(n5780), .Z(n5783) );
  XOR U6789 ( .A(n5784), .B(n5785), .Z(n5780) );
  ANDN U6790 ( .B(n5786), .A(n5787), .Z(n5784) );
  XNOR U6791 ( .A(b[3092]), .B(n5785), .Z(n5786) );
  XNOR U6792 ( .A(b[3092]), .B(n5787), .Z(c[3092]) );
  XNOR U6793 ( .A(a[3092]), .B(n5788), .Z(n5787) );
  IV U6794 ( .A(n5785), .Z(n5788) );
  XOR U6795 ( .A(n5789), .B(n5790), .Z(n5785) );
  ANDN U6796 ( .B(n5791), .A(n5792), .Z(n5789) );
  XNOR U6797 ( .A(b[3091]), .B(n5790), .Z(n5791) );
  XNOR U6798 ( .A(b[3091]), .B(n5792), .Z(c[3091]) );
  XNOR U6799 ( .A(a[3091]), .B(n5793), .Z(n5792) );
  IV U6800 ( .A(n5790), .Z(n5793) );
  XOR U6801 ( .A(n5794), .B(n5795), .Z(n5790) );
  ANDN U6802 ( .B(n5796), .A(n5797), .Z(n5794) );
  XNOR U6803 ( .A(b[3090]), .B(n5795), .Z(n5796) );
  XNOR U6804 ( .A(b[3090]), .B(n5797), .Z(c[3090]) );
  XNOR U6805 ( .A(a[3090]), .B(n5798), .Z(n5797) );
  IV U6806 ( .A(n5795), .Z(n5798) );
  XOR U6807 ( .A(n5799), .B(n5800), .Z(n5795) );
  ANDN U6808 ( .B(n5801), .A(n5802), .Z(n5799) );
  XNOR U6809 ( .A(b[3089]), .B(n5800), .Z(n5801) );
  XNOR U6810 ( .A(b[308]), .B(n5803), .Z(c[308]) );
  XNOR U6811 ( .A(b[3089]), .B(n5802), .Z(c[3089]) );
  XNOR U6812 ( .A(a[3089]), .B(n5804), .Z(n5802) );
  IV U6813 ( .A(n5800), .Z(n5804) );
  XOR U6814 ( .A(n5805), .B(n5806), .Z(n5800) );
  ANDN U6815 ( .B(n5807), .A(n5808), .Z(n5805) );
  XNOR U6816 ( .A(b[3088]), .B(n5806), .Z(n5807) );
  XNOR U6817 ( .A(b[3088]), .B(n5808), .Z(c[3088]) );
  XNOR U6818 ( .A(a[3088]), .B(n5809), .Z(n5808) );
  IV U6819 ( .A(n5806), .Z(n5809) );
  XOR U6820 ( .A(n5810), .B(n5811), .Z(n5806) );
  ANDN U6821 ( .B(n5812), .A(n5813), .Z(n5810) );
  XNOR U6822 ( .A(b[3087]), .B(n5811), .Z(n5812) );
  XNOR U6823 ( .A(b[3087]), .B(n5813), .Z(c[3087]) );
  XNOR U6824 ( .A(a[3087]), .B(n5814), .Z(n5813) );
  IV U6825 ( .A(n5811), .Z(n5814) );
  XOR U6826 ( .A(n5815), .B(n5816), .Z(n5811) );
  ANDN U6827 ( .B(n5817), .A(n5818), .Z(n5815) );
  XNOR U6828 ( .A(b[3086]), .B(n5816), .Z(n5817) );
  XNOR U6829 ( .A(b[3086]), .B(n5818), .Z(c[3086]) );
  XNOR U6830 ( .A(a[3086]), .B(n5819), .Z(n5818) );
  IV U6831 ( .A(n5816), .Z(n5819) );
  XOR U6832 ( .A(n5820), .B(n5821), .Z(n5816) );
  ANDN U6833 ( .B(n5822), .A(n5823), .Z(n5820) );
  XNOR U6834 ( .A(b[3085]), .B(n5821), .Z(n5822) );
  XNOR U6835 ( .A(b[3085]), .B(n5823), .Z(c[3085]) );
  XNOR U6836 ( .A(a[3085]), .B(n5824), .Z(n5823) );
  IV U6837 ( .A(n5821), .Z(n5824) );
  XOR U6838 ( .A(n5825), .B(n5826), .Z(n5821) );
  ANDN U6839 ( .B(n5827), .A(n5828), .Z(n5825) );
  XNOR U6840 ( .A(b[3084]), .B(n5826), .Z(n5827) );
  XNOR U6841 ( .A(b[3084]), .B(n5828), .Z(c[3084]) );
  XNOR U6842 ( .A(a[3084]), .B(n5829), .Z(n5828) );
  IV U6843 ( .A(n5826), .Z(n5829) );
  XOR U6844 ( .A(n5830), .B(n5831), .Z(n5826) );
  ANDN U6845 ( .B(n5832), .A(n5833), .Z(n5830) );
  XNOR U6846 ( .A(b[3083]), .B(n5831), .Z(n5832) );
  XNOR U6847 ( .A(b[3083]), .B(n5833), .Z(c[3083]) );
  XNOR U6848 ( .A(a[3083]), .B(n5834), .Z(n5833) );
  IV U6849 ( .A(n5831), .Z(n5834) );
  XOR U6850 ( .A(n5835), .B(n5836), .Z(n5831) );
  ANDN U6851 ( .B(n5837), .A(n5838), .Z(n5835) );
  XNOR U6852 ( .A(b[3082]), .B(n5836), .Z(n5837) );
  XNOR U6853 ( .A(b[3082]), .B(n5838), .Z(c[3082]) );
  XNOR U6854 ( .A(a[3082]), .B(n5839), .Z(n5838) );
  IV U6855 ( .A(n5836), .Z(n5839) );
  XOR U6856 ( .A(n5840), .B(n5841), .Z(n5836) );
  ANDN U6857 ( .B(n5842), .A(n5843), .Z(n5840) );
  XNOR U6858 ( .A(b[3081]), .B(n5841), .Z(n5842) );
  XNOR U6859 ( .A(b[3081]), .B(n5843), .Z(c[3081]) );
  XNOR U6860 ( .A(a[3081]), .B(n5844), .Z(n5843) );
  IV U6861 ( .A(n5841), .Z(n5844) );
  XOR U6862 ( .A(n5845), .B(n5846), .Z(n5841) );
  ANDN U6863 ( .B(n5847), .A(n5848), .Z(n5845) );
  XNOR U6864 ( .A(b[3080]), .B(n5846), .Z(n5847) );
  XNOR U6865 ( .A(b[3080]), .B(n5848), .Z(c[3080]) );
  XNOR U6866 ( .A(a[3080]), .B(n5849), .Z(n5848) );
  IV U6867 ( .A(n5846), .Z(n5849) );
  XOR U6868 ( .A(n5850), .B(n5851), .Z(n5846) );
  ANDN U6869 ( .B(n5852), .A(n5853), .Z(n5850) );
  XNOR U6870 ( .A(b[3079]), .B(n5851), .Z(n5852) );
  XNOR U6871 ( .A(b[307]), .B(n5854), .Z(c[307]) );
  XNOR U6872 ( .A(b[3079]), .B(n5853), .Z(c[3079]) );
  XNOR U6873 ( .A(a[3079]), .B(n5855), .Z(n5853) );
  IV U6874 ( .A(n5851), .Z(n5855) );
  XOR U6875 ( .A(n5856), .B(n5857), .Z(n5851) );
  ANDN U6876 ( .B(n5858), .A(n5859), .Z(n5856) );
  XNOR U6877 ( .A(b[3078]), .B(n5857), .Z(n5858) );
  XNOR U6878 ( .A(b[3078]), .B(n5859), .Z(c[3078]) );
  XNOR U6879 ( .A(a[3078]), .B(n5860), .Z(n5859) );
  IV U6880 ( .A(n5857), .Z(n5860) );
  XOR U6881 ( .A(n5861), .B(n5862), .Z(n5857) );
  ANDN U6882 ( .B(n5863), .A(n5864), .Z(n5861) );
  XNOR U6883 ( .A(b[3077]), .B(n5862), .Z(n5863) );
  XNOR U6884 ( .A(b[3077]), .B(n5864), .Z(c[3077]) );
  XNOR U6885 ( .A(a[3077]), .B(n5865), .Z(n5864) );
  IV U6886 ( .A(n5862), .Z(n5865) );
  XOR U6887 ( .A(n5866), .B(n5867), .Z(n5862) );
  ANDN U6888 ( .B(n5868), .A(n5869), .Z(n5866) );
  XNOR U6889 ( .A(b[3076]), .B(n5867), .Z(n5868) );
  XNOR U6890 ( .A(b[3076]), .B(n5869), .Z(c[3076]) );
  XNOR U6891 ( .A(a[3076]), .B(n5870), .Z(n5869) );
  IV U6892 ( .A(n5867), .Z(n5870) );
  XOR U6893 ( .A(n5871), .B(n5872), .Z(n5867) );
  ANDN U6894 ( .B(n5873), .A(n5874), .Z(n5871) );
  XNOR U6895 ( .A(b[3075]), .B(n5872), .Z(n5873) );
  XNOR U6896 ( .A(b[3075]), .B(n5874), .Z(c[3075]) );
  XNOR U6897 ( .A(a[3075]), .B(n5875), .Z(n5874) );
  IV U6898 ( .A(n5872), .Z(n5875) );
  XOR U6899 ( .A(n5876), .B(n5877), .Z(n5872) );
  ANDN U6900 ( .B(n5878), .A(n5879), .Z(n5876) );
  XNOR U6901 ( .A(b[3074]), .B(n5877), .Z(n5878) );
  XNOR U6902 ( .A(b[3074]), .B(n5879), .Z(c[3074]) );
  XNOR U6903 ( .A(a[3074]), .B(n5880), .Z(n5879) );
  IV U6904 ( .A(n5877), .Z(n5880) );
  XOR U6905 ( .A(n5881), .B(n5882), .Z(n5877) );
  ANDN U6906 ( .B(n5883), .A(n5884), .Z(n5881) );
  XNOR U6907 ( .A(b[3073]), .B(n5882), .Z(n5883) );
  XNOR U6908 ( .A(b[3073]), .B(n5884), .Z(c[3073]) );
  XNOR U6909 ( .A(a[3073]), .B(n5885), .Z(n5884) );
  IV U6910 ( .A(n5882), .Z(n5885) );
  XOR U6911 ( .A(n5886), .B(n5887), .Z(n5882) );
  ANDN U6912 ( .B(n5888), .A(n5889), .Z(n5886) );
  XNOR U6913 ( .A(b[3072]), .B(n5887), .Z(n5888) );
  XNOR U6914 ( .A(b[3072]), .B(n5889), .Z(c[3072]) );
  XNOR U6915 ( .A(a[3072]), .B(n5890), .Z(n5889) );
  IV U6916 ( .A(n5887), .Z(n5890) );
  XOR U6917 ( .A(n5891), .B(n5892), .Z(n5887) );
  ANDN U6918 ( .B(n5893), .A(n5894), .Z(n5891) );
  XNOR U6919 ( .A(b[3071]), .B(n5892), .Z(n5893) );
  XNOR U6920 ( .A(b[3071]), .B(n5894), .Z(c[3071]) );
  XNOR U6921 ( .A(a[3071]), .B(n5895), .Z(n5894) );
  IV U6922 ( .A(n5892), .Z(n5895) );
  XOR U6923 ( .A(n5896), .B(n5897), .Z(n5892) );
  ANDN U6924 ( .B(n5898), .A(n5899), .Z(n5896) );
  XNOR U6925 ( .A(b[3070]), .B(n5897), .Z(n5898) );
  XNOR U6926 ( .A(b[3070]), .B(n5899), .Z(c[3070]) );
  XNOR U6927 ( .A(a[3070]), .B(n5900), .Z(n5899) );
  IV U6928 ( .A(n5897), .Z(n5900) );
  XOR U6929 ( .A(n5901), .B(n5902), .Z(n5897) );
  ANDN U6930 ( .B(n5903), .A(n5904), .Z(n5901) );
  XNOR U6931 ( .A(b[3069]), .B(n5902), .Z(n5903) );
  XNOR U6932 ( .A(b[306]), .B(n5905), .Z(c[306]) );
  XNOR U6933 ( .A(b[3069]), .B(n5904), .Z(c[3069]) );
  XNOR U6934 ( .A(a[3069]), .B(n5906), .Z(n5904) );
  IV U6935 ( .A(n5902), .Z(n5906) );
  XOR U6936 ( .A(n5907), .B(n5908), .Z(n5902) );
  ANDN U6937 ( .B(n5909), .A(n5910), .Z(n5907) );
  XNOR U6938 ( .A(b[3068]), .B(n5908), .Z(n5909) );
  XNOR U6939 ( .A(b[3068]), .B(n5910), .Z(c[3068]) );
  XNOR U6940 ( .A(a[3068]), .B(n5911), .Z(n5910) );
  IV U6941 ( .A(n5908), .Z(n5911) );
  XOR U6942 ( .A(n5912), .B(n5913), .Z(n5908) );
  ANDN U6943 ( .B(n5914), .A(n5915), .Z(n5912) );
  XNOR U6944 ( .A(b[3067]), .B(n5913), .Z(n5914) );
  XNOR U6945 ( .A(b[3067]), .B(n5915), .Z(c[3067]) );
  XNOR U6946 ( .A(a[3067]), .B(n5916), .Z(n5915) );
  IV U6947 ( .A(n5913), .Z(n5916) );
  XOR U6948 ( .A(n5917), .B(n5918), .Z(n5913) );
  ANDN U6949 ( .B(n5919), .A(n5920), .Z(n5917) );
  XNOR U6950 ( .A(b[3066]), .B(n5918), .Z(n5919) );
  XNOR U6951 ( .A(b[3066]), .B(n5920), .Z(c[3066]) );
  XNOR U6952 ( .A(a[3066]), .B(n5921), .Z(n5920) );
  IV U6953 ( .A(n5918), .Z(n5921) );
  XOR U6954 ( .A(n5922), .B(n5923), .Z(n5918) );
  ANDN U6955 ( .B(n5924), .A(n5925), .Z(n5922) );
  XNOR U6956 ( .A(b[3065]), .B(n5923), .Z(n5924) );
  XNOR U6957 ( .A(b[3065]), .B(n5925), .Z(c[3065]) );
  XNOR U6958 ( .A(a[3065]), .B(n5926), .Z(n5925) );
  IV U6959 ( .A(n5923), .Z(n5926) );
  XOR U6960 ( .A(n5927), .B(n5928), .Z(n5923) );
  ANDN U6961 ( .B(n5929), .A(n5930), .Z(n5927) );
  XNOR U6962 ( .A(b[3064]), .B(n5928), .Z(n5929) );
  XNOR U6963 ( .A(b[3064]), .B(n5930), .Z(c[3064]) );
  XNOR U6964 ( .A(a[3064]), .B(n5931), .Z(n5930) );
  IV U6965 ( .A(n5928), .Z(n5931) );
  XOR U6966 ( .A(n5932), .B(n5933), .Z(n5928) );
  ANDN U6967 ( .B(n5934), .A(n5935), .Z(n5932) );
  XNOR U6968 ( .A(b[3063]), .B(n5933), .Z(n5934) );
  XNOR U6969 ( .A(b[3063]), .B(n5935), .Z(c[3063]) );
  XNOR U6970 ( .A(a[3063]), .B(n5936), .Z(n5935) );
  IV U6971 ( .A(n5933), .Z(n5936) );
  XOR U6972 ( .A(n5937), .B(n5938), .Z(n5933) );
  ANDN U6973 ( .B(n5939), .A(n5940), .Z(n5937) );
  XNOR U6974 ( .A(b[3062]), .B(n5938), .Z(n5939) );
  XNOR U6975 ( .A(b[3062]), .B(n5940), .Z(c[3062]) );
  XNOR U6976 ( .A(a[3062]), .B(n5941), .Z(n5940) );
  IV U6977 ( .A(n5938), .Z(n5941) );
  XOR U6978 ( .A(n5942), .B(n5943), .Z(n5938) );
  ANDN U6979 ( .B(n5944), .A(n5945), .Z(n5942) );
  XNOR U6980 ( .A(b[3061]), .B(n5943), .Z(n5944) );
  XNOR U6981 ( .A(b[3061]), .B(n5945), .Z(c[3061]) );
  XNOR U6982 ( .A(a[3061]), .B(n5946), .Z(n5945) );
  IV U6983 ( .A(n5943), .Z(n5946) );
  XOR U6984 ( .A(n5947), .B(n5948), .Z(n5943) );
  ANDN U6985 ( .B(n5949), .A(n5950), .Z(n5947) );
  XNOR U6986 ( .A(b[3060]), .B(n5948), .Z(n5949) );
  XNOR U6987 ( .A(b[3060]), .B(n5950), .Z(c[3060]) );
  XNOR U6988 ( .A(a[3060]), .B(n5951), .Z(n5950) );
  IV U6989 ( .A(n5948), .Z(n5951) );
  XOR U6990 ( .A(n5952), .B(n5953), .Z(n5948) );
  ANDN U6991 ( .B(n5954), .A(n5955), .Z(n5952) );
  XNOR U6992 ( .A(b[3059]), .B(n5953), .Z(n5954) );
  XNOR U6993 ( .A(b[305]), .B(n5956), .Z(c[305]) );
  XNOR U6994 ( .A(b[3059]), .B(n5955), .Z(c[3059]) );
  XNOR U6995 ( .A(a[3059]), .B(n5957), .Z(n5955) );
  IV U6996 ( .A(n5953), .Z(n5957) );
  XOR U6997 ( .A(n5958), .B(n5959), .Z(n5953) );
  ANDN U6998 ( .B(n5960), .A(n5961), .Z(n5958) );
  XNOR U6999 ( .A(b[3058]), .B(n5959), .Z(n5960) );
  XNOR U7000 ( .A(b[3058]), .B(n5961), .Z(c[3058]) );
  XNOR U7001 ( .A(a[3058]), .B(n5962), .Z(n5961) );
  IV U7002 ( .A(n5959), .Z(n5962) );
  XOR U7003 ( .A(n5963), .B(n5964), .Z(n5959) );
  ANDN U7004 ( .B(n5965), .A(n5966), .Z(n5963) );
  XNOR U7005 ( .A(b[3057]), .B(n5964), .Z(n5965) );
  XNOR U7006 ( .A(b[3057]), .B(n5966), .Z(c[3057]) );
  XNOR U7007 ( .A(a[3057]), .B(n5967), .Z(n5966) );
  IV U7008 ( .A(n5964), .Z(n5967) );
  XOR U7009 ( .A(n5968), .B(n5969), .Z(n5964) );
  ANDN U7010 ( .B(n5970), .A(n5971), .Z(n5968) );
  XNOR U7011 ( .A(b[3056]), .B(n5969), .Z(n5970) );
  XNOR U7012 ( .A(b[3056]), .B(n5971), .Z(c[3056]) );
  XNOR U7013 ( .A(a[3056]), .B(n5972), .Z(n5971) );
  IV U7014 ( .A(n5969), .Z(n5972) );
  XOR U7015 ( .A(n5973), .B(n5974), .Z(n5969) );
  ANDN U7016 ( .B(n5975), .A(n5976), .Z(n5973) );
  XNOR U7017 ( .A(b[3055]), .B(n5974), .Z(n5975) );
  XNOR U7018 ( .A(b[3055]), .B(n5976), .Z(c[3055]) );
  XNOR U7019 ( .A(a[3055]), .B(n5977), .Z(n5976) );
  IV U7020 ( .A(n5974), .Z(n5977) );
  XOR U7021 ( .A(n5978), .B(n5979), .Z(n5974) );
  ANDN U7022 ( .B(n5980), .A(n5981), .Z(n5978) );
  XNOR U7023 ( .A(b[3054]), .B(n5979), .Z(n5980) );
  XNOR U7024 ( .A(b[3054]), .B(n5981), .Z(c[3054]) );
  XNOR U7025 ( .A(a[3054]), .B(n5982), .Z(n5981) );
  IV U7026 ( .A(n5979), .Z(n5982) );
  XOR U7027 ( .A(n5983), .B(n5984), .Z(n5979) );
  ANDN U7028 ( .B(n5985), .A(n5986), .Z(n5983) );
  XNOR U7029 ( .A(b[3053]), .B(n5984), .Z(n5985) );
  XNOR U7030 ( .A(b[3053]), .B(n5986), .Z(c[3053]) );
  XNOR U7031 ( .A(a[3053]), .B(n5987), .Z(n5986) );
  IV U7032 ( .A(n5984), .Z(n5987) );
  XOR U7033 ( .A(n5988), .B(n5989), .Z(n5984) );
  ANDN U7034 ( .B(n5990), .A(n5991), .Z(n5988) );
  XNOR U7035 ( .A(b[3052]), .B(n5989), .Z(n5990) );
  XNOR U7036 ( .A(b[3052]), .B(n5991), .Z(c[3052]) );
  XNOR U7037 ( .A(a[3052]), .B(n5992), .Z(n5991) );
  IV U7038 ( .A(n5989), .Z(n5992) );
  XOR U7039 ( .A(n5993), .B(n5994), .Z(n5989) );
  ANDN U7040 ( .B(n5995), .A(n5996), .Z(n5993) );
  XNOR U7041 ( .A(b[3051]), .B(n5994), .Z(n5995) );
  XNOR U7042 ( .A(b[3051]), .B(n5996), .Z(c[3051]) );
  XNOR U7043 ( .A(a[3051]), .B(n5997), .Z(n5996) );
  IV U7044 ( .A(n5994), .Z(n5997) );
  XOR U7045 ( .A(n5998), .B(n5999), .Z(n5994) );
  ANDN U7046 ( .B(n6000), .A(n6001), .Z(n5998) );
  XNOR U7047 ( .A(b[3050]), .B(n5999), .Z(n6000) );
  XNOR U7048 ( .A(b[3050]), .B(n6001), .Z(c[3050]) );
  XNOR U7049 ( .A(a[3050]), .B(n6002), .Z(n6001) );
  IV U7050 ( .A(n5999), .Z(n6002) );
  XOR U7051 ( .A(n6003), .B(n6004), .Z(n5999) );
  ANDN U7052 ( .B(n6005), .A(n6006), .Z(n6003) );
  XNOR U7053 ( .A(b[3049]), .B(n6004), .Z(n6005) );
  XNOR U7054 ( .A(b[304]), .B(n6007), .Z(c[304]) );
  XNOR U7055 ( .A(b[3049]), .B(n6006), .Z(c[3049]) );
  XNOR U7056 ( .A(a[3049]), .B(n6008), .Z(n6006) );
  IV U7057 ( .A(n6004), .Z(n6008) );
  XOR U7058 ( .A(n6009), .B(n6010), .Z(n6004) );
  ANDN U7059 ( .B(n6011), .A(n6012), .Z(n6009) );
  XNOR U7060 ( .A(b[3048]), .B(n6010), .Z(n6011) );
  XNOR U7061 ( .A(b[3048]), .B(n6012), .Z(c[3048]) );
  XNOR U7062 ( .A(a[3048]), .B(n6013), .Z(n6012) );
  IV U7063 ( .A(n6010), .Z(n6013) );
  XOR U7064 ( .A(n6014), .B(n6015), .Z(n6010) );
  ANDN U7065 ( .B(n6016), .A(n6017), .Z(n6014) );
  XNOR U7066 ( .A(b[3047]), .B(n6015), .Z(n6016) );
  XNOR U7067 ( .A(b[3047]), .B(n6017), .Z(c[3047]) );
  XNOR U7068 ( .A(a[3047]), .B(n6018), .Z(n6017) );
  IV U7069 ( .A(n6015), .Z(n6018) );
  XOR U7070 ( .A(n6019), .B(n6020), .Z(n6015) );
  ANDN U7071 ( .B(n6021), .A(n6022), .Z(n6019) );
  XNOR U7072 ( .A(b[3046]), .B(n6020), .Z(n6021) );
  XNOR U7073 ( .A(b[3046]), .B(n6022), .Z(c[3046]) );
  XNOR U7074 ( .A(a[3046]), .B(n6023), .Z(n6022) );
  IV U7075 ( .A(n6020), .Z(n6023) );
  XOR U7076 ( .A(n6024), .B(n6025), .Z(n6020) );
  ANDN U7077 ( .B(n6026), .A(n6027), .Z(n6024) );
  XNOR U7078 ( .A(b[3045]), .B(n6025), .Z(n6026) );
  XNOR U7079 ( .A(b[3045]), .B(n6027), .Z(c[3045]) );
  XNOR U7080 ( .A(a[3045]), .B(n6028), .Z(n6027) );
  IV U7081 ( .A(n6025), .Z(n6028) );
  XOR U7082 ( .A(n6029), .B(n6030), .Z(n6025) );
  ANDN U7083 ( .B(n6031), .A(n6032), .Z(n6029) );
  XNOR U7084 ( .A(b[3044]), .B(n6030), .Z(n6031) );
  XNOR U7085 ( .A(b[3044]), .B(n6032), .Z(c[3044]) );
  XNOR U7086 ( .A(a[3044]), .B(n6033), .Z(n6032) );
  IV U7087 ( .A(n6030), .Z(n6033) );
  XOR U7088 ( .A(n6034), .B(n6035), .Z(n6030) );
  ANDN U7089 ( .B(n6036), .A(n6037), .Z(n6034) );
  XNOR U7090 ( .A(b[3043]), .B(n6035), .Z(n6036) );
  XNOR U7091 ( .A(b[3043]), .B(n6037), .Z(c[3043]) );
  XNOR U7092 ( .A(a[3043]), .B(n6038), .Z(n6037) );
  IV U7093 ( .A(n6035), .Z(n6038) );
  XOR U7094 ( .A(n6039), .B(n6040), .Z(n6035) );
  ANDN U7095 ( .B(n6041), .A(n6042), .Z(n6039) );
  XNOR U7096 ( .A(b[3042]), .B(n6040), .Z(n6041) );
  XNOR U7097 ( .A(b[3042]), .B(n6042), .Z(c[3042]) );
  XNOR U7098 ( .A(a[3042]), .B(n6043), .Z(n6042) );
  IV U7099 ( .A(n6040), .Z(n6043) );
  XOR U7100 ( .A(n6044), .B(n6045), .Z(n6040) );
  ANDN U7101 ( .B(n6046), .A(n6047), .Z(n6044) );
  XNOR U7102 ( .A(b[3041]), .B(n6045), .Z(n6046) );
  XNOR U7103 ( .A(b[3041]), .B(n6047), .Z(c[3041]) );
  XNOR U7104 ( .A(a[3041]), .B(n6048), .Z(n6047) );
  IV U7105 ( .A(n6045), .Z(n6048) );
  XOR U7106 ( .A(n6049), .B(n6050), .Z(n6045) );
  ANDN U7107 ( .B(n6051), .A(n6052), .Z(n6049) );
  XNOR U7108 ( .A(b[3040]), .B(n6050), .Z(n6051) );
  XNOR U7109 ( .A(b[3040]), .B(n6052), .Z(c[3040]) );
  XNOR U7110 ( .A(a[3040]), .B(n6053), .Z(n6052) );
  IV U7111 ( .A(n6050), .Z(n6053) );
  XOR U7112 ( .A(n6054), .B(n6055), .Z(n6050) );
  ANDN U7113 ( .B(n6056), .A(n6057), .Z(n6054) );
  XNOR U7114 ( .A(b[3039]), .B(n6055), .Z(n6056) );
  XNOR U7115 ( .A(b[303]), .B(n6058), .Z(c[303]) );
  XNOR U7116 ( .A(b[3039]), .B(n6057), .Z(c[3039]) );
  XNOR U7117 ( .A(a[3039]), .B(n6059), .Z(n6057) );
  IV U7118 ( .A(n6055), .Z(n6059) );
  XOR U7119 ( .A(n6060), .B(n6061), .Z(n6055) );
  ANDN U7120 ( .B(n6062), .A(n6063), .Z(n6060) );
  XNOR U7121 ( .A(b[3038]), .B(n6061), .Z(n6062) );
  XNOR U7122 ( .A(b[3038]), .B(n6063), .Z(c[3038]) );
  XNOR U7123 ( .A(a[3038]), .B(n6064), .Z(n6063) );
  IV U7124 ( .A(n6061), .Z(n6064) );
  XOR U7125 ( .A(n6065), .B(n6066), .Z(n6061) );
  ANDN U7126 ( .B(n6067), .A(n6068), .Z(n6065) );
  XNOR U7127 ( .A(b[3037]), .B(n6066), .Z(n6067) );
  XNOR U7128 ( .A(b[3037]), .B(n6068), .Z(c[3037]) );
  XNOR U7129 ( .A(a[3037]), .B(n6069), .Z(n6068) );
  IV U7130 ( .A(n6066), .Z(n6069) );
  XOR U7131 ( .A(n6070), .B(n6071), .Z(n6066) );
  ANDN U7132 ( .B(n6072), .A(n6073), .Z(n6070) );
  XNOR U7133 ( .A(b[3036]), .B(n6071), .Z(n6072) );
  XNOR U7134 ( .A(b[3036]), .B(n6073), .Z(c[3036]) );
  XNOR U7135 ( .A(a[3036]), .B(n6074), .Z(n6073) );
  IV U7136 ( .A(n6071), .Z(n6074) );
  XOR U7137 ( .A(n6075), .B(n6076), .Z(n6071) );
  ANDN U7138 ( .B(n6077), .A(n6078), .Z(n6075) );
  XNOR U7139 ( .A(b[3035]), .B(n6076), .Z(n6077) );
  XNOR U7140 ( .A(b[3035]), .B(n6078), .Z(c[3035]) );
  XNOR U7141 ( .A(a[3035]), .B(n6079), .Z(n6078) );
  IV U7142 ( .A(n6076), .Z(n6079) );
  XOR U7143 ( .A(n6080), .B(n6081), .Z(n6076) );
  ANDN U7144 ( .B(n6082), .A(n6083), .Z(n6080) );
  XNOR U7145 ( .A(b[3034]), .B(n6081), .Z(n6082) );
  XNOR U7146 ( .A(b[3034]), .B(n6083), .Z(c[3034]) );
  XNOR U7147 ( .A(a[3034]), .B(n6084), .Z(n6083) );
  IV U7148 ( .A(n6081), .Z(n6084) );
  XOR U7149 ( .A(n6085), .B(n6086), .Z(n6081) );
  ANDN U7150 ( .B(n6087), .A(n6088), .Z(n6085) );
  XNOR U7151 ( .A(b[3033]), .B(n6086), .Z(n6087) );
  XNOR U7152 ( .A(b[3033]), .B(n6088), .Z(c[3033]) );
  XNOR U7153 ( .A(a[3033]), .B(n6089), .Z(n6088) );
  IV U7154 ( .A(n6086), .Z(n6089) );
  XOR U7155 ( .A(n6090), .B(n6091), .Z(n6086) );
  ANDN U7156 ( .B(n6092), .A(n6093), .Z(n6090) );
  XNOR U7157 ( .A(b[3032]), .B(n6091), .Z(n6092) );
  XNOR U7158 ( .A(b[3032]), .B(n6093), .Z(c[3032]) );
  XNOR U7159 ( .A(a[3032]), .B(n6094), .Z(n6093) );
  IV U7160 ( .A(n6091), .Z(n6094) );
  XOR U7161 ( .A(n6095), .B(n6096), .Z(n6091) );
  ANDN U7162 ( .B(n6097), .A(n6098), .Z(n6095) );
  XNOR U7163 ( .A(b[3031]), .B(n6096), .Z(n6097) );
  XNOR U7164 ( .A(b[3031]), .B(n6098), .Z(c[3031]) );
  XNOR U7165 ( .A(a[3031]), .B(n6099), .Z(n6098) );
  IV U7166 ( .A(n6096), .Z(n6099) );
  XOR U7167 ( .A(n6100), .B(n6101), .Z(n6096) );
  ANDN U7168 ( .B(n6102), .A(n6103), .Z(n6100) );
  XNOR U7169 ( .A(b[3030]), .B(n6101), .Z(n6102) );
  XNOR U7170 ( .A(b[3030]), .B(n6103), .Z(c[3030]) );
  XNOR U7171 ( .A(a[3030]), .B(n6104), .Z(n6103) );
  IV U7172 ( .A(n6101), .Z(n6104) );
  XOR U7173 ( .A(n6105), .B(n6106), .Z(n6101) );
  ANDN U7174 ( .B(n6107), .A(n6108), .Z(n6105) );
  XNOR U7175 ( .A(b[3029]), .B(n6106), .Z(n6107) );
  XNOR U7176 ( .A(b[302]), .B(n6109), .Z(c[302]) );
  XNOR U7177 ( .A(b[3029]), .B(n6108), .Z(c[3029]) );
  XNOR U7178 ( .A(a[3029]), .B(n6110), .Z(n6108) );
  IV U7179 ( .A(n6106), .Z(n6110) );
  XOR U7180 ( .A(n6111), .B(n6112), .Z(n6106) );
  ANDN U7181 ( .B(n6113), .A(n6114), .Z(n6111) );
  XNOR U7182 ( .A(b[3028]), .B(n6112), .Z(n6113) );
  XNOR U7183 ( .A(b[3028]), .B(n6114), .Z(c[3028]) );
  XNOR U7184 ( .A(a[3028]), .B(n6115), .Z(n6114) );
  IV U7185 ( .A(n6112), .Z(n6115) );
  XOR U7186 ( .A(n6116), .B(n6117), .Z(n6112) );
  ANDN U7187 ( .B(n6118), .A(n6119), .Z(n6116) );
  XNOR U7188 ( .A(b[3027]), .B(n6117), .Z(n6118) );
  XNOR U7189 ( .A(b[3027]), .B(n6119), .Z(c[3027]) );
  XNOR U7190 ( .A(a[3027]), .B(n6120), .Z(n6119) );
  IV U7191 ( .A(n6117), .Z(n6120) );
  XOR U7192 ( .A(n6121), .B(n6122), .Z(n6117) );
  ANDN U7193 ( .B(n6123), .A(n6124), .Z(n6121) );
  XNOR U7194 ( .A(b[3026]), .B(n6122), .Z(n6123) );
  XNOR U7195 ( .A(b[3026]), .B(n6124), .Z(c[3026]) );
  XNOR U7196 ( .A(a[3026]), .B(n6125), .Z(n6124) );
  IV U7197 ( .A(n6122), .Z(n6125) );
  XOR U7198 ( .A(n6126), .B(n6127), .Z(n6122) );
  ANDN U7199 ( .B(n6128), .A(n6129), .Z(n6126) );
  XNOR U7200 ( .A(b[3025]), .B(n6127), .Z(n6128) );
  XNOR U7201 ( .A(b[3025]), .B(n6129), .Z(c[3025]) );
  XNOR U7202 ( .A(a[3025]), .B(n6130), .Z(n6129) );
  IV U7203 ( .A(n6127), .Z(n6130) );
  XOR U7204 ( .A(n6131), .B(n6132), .Z(n6127) );
  ANDN U7205 ( .B(n6133), .A(n6134), .Z(n6131) );
  XNOR U7206 ( .A(b[3024]), .B(n6132), .Z(n6133) );
  XNOR U7207 ( .A(b[3024]), .B(n6134), .Z(c[3024]) );
  XNOR U7208 ( .A(a[3024]), .B(n6135), .Z(n6134) );
  IV U7209 ( .A(n6132), .Z(n6135) );
  XOR U7210 ( .A(n6136), .B(n6137), .Z(n6132) );
  ANDN U7211 ( .B(n6138), .A(n6139), .Z(n6136) );
  XNOR U7212 ( .A(b[3023]), .B(n6137), .Z(n6138) );
  XNOR U7213 ( .A(b[3023]), .B(n6139), .Z(c[3023]) );
  XNOR U7214 ( .A(a[3023]), .B(n6140), .Z(n6139) );
  IV U7215 ( .A(n6137), .Z(n6140) );
  XOR U7216 ( .A(n6141), .B(n6142), .Z(n6137) );
  ANDN U7217 ( .B(n6143), .A(n6144), .Z(n6141) );
  XNOR U7218 ( .A(b[3022]), .B(n6142), .Z(n6143) );
  XNOR U7219 ( .A(b[3022]), .B(n6144), .Z(c[3022]) );
  XNOR U7220 ( .A(a[3022]), .B(n6145), .Z(n6144) );
  IV U7221 ( .A(n6142), .Z(n6145) );
  XOR U7222 ( .A(n6146), .B(n6147), .Z(n6142) );
  ANDN U7223 ( .B(n6148), .A(n6149), .Z(n6146) );
  XNOR U7224 ( .A(b[3021]), .B(n6147), .Z(n6148) );
  XNOR U7225 ( .A(b[3021]), .B(n6149), .Z(c[3021]) );
  XNOR U7226 ( .A(a[3021]), .B(n6150), .Z(n6149) );
  IV U7227 ( .A(n6147), .Z(n6150) );
  XOR U7228 ( .A(n6151), .B(n6152), .Z(n6147) );
  ANDN U7229 ( .B(n6153), .A(n6154), .Z(n6151) );
  XNOR U7230 ( .A(b[3020]), .B(n6152), .Z(n6153) );
  XNOR U7231 ( .A(b[3020]), .B(n6154), .Z(c[3020]) );
  XNOR U7232 ( .A(a[3020]), .B(n6155), .Z(n6154) );
  IV U7233 ( .A(n6152), .Z(n6155) );
  XOR U7234 ( .A(n6156), .B(n6157), .Z(n6152) );
  ANDN U7235 ( .B(n6158), .A(n6159), .Z(n6156) );
  XNOR U7236 ( .A(b[3019]), .B(n6157), .Z(n6158) );
  XNOR U7237 ( .A(b[301]), .B(n6160), .Z(c[301]) );
  XNOR U7238 ( .A(b[3019]), .B(n6159), .Z(c[3019]) );
  XNOR U7239 ( .A(a[3019]), .B(n6161), .Z(n6159) );
  IV U7240 ( .A(n6157), .Z(n6161) );
  XOR U7241 ( .A(n6162), .B(n6163), .Z(n6157) );
  ANDN U7242 ( .B(n6164), .A(n6165), .Z(n6162) );
  XNOR U7243 ( .A(b[3018]), .B(n6163), .Z(n6164) );
  XNOR U7244 ( .A(b[3018]), .B(n6165), .Z(c[3018]) );
  XNOR U7245 ( .A(a[3018]), .B(n6166), .Z(n6165) );
  IV U7246 ( .A(n6163), .Z(n6166) );
  XOR U7247 ( .A(n6167), .B(n6168), .Z(n6163) );
  ANDN U7248 ( .B(n6169), .A(n6170), .Z(n6167) );
  XNOR U7249 ( .A(b[3017]), .B(n6168), .Z(n6169) );
  XNOR U7250 ( .A(b[3017]), .B(n6170), .Z(c[3017]) );
  XNOR U7251 ( .A(a[3017]), .B(n6171), .Z(n6170) );
  IV U7252 ( .A(n6168), .Z(n6171) );
  XOR U7253 ( .A(n6172), .B(n6173), .Z(n6168) );
  ANDN U7254 ( .B(n6174), .A(n6175), .Z(n6172) );
  XNOR U7255 ( .A(b[3016]), .B(n6173), .Z(n6174) );
  XNOR U7256 ( .A(b[3016]), .B(n6175), .Z(c[3016]) );
  XNOR U7257 ( .A(a[3016]), .B(n6176), .Z(n6175) );
  IV U7258 ( .A(n6173), .Z(n6176) );
  XOR U7259 ( .A(n6177), .B(n6178), .Z(n6173) );
  ANDN U7260 ( .B(n6179), .A(n6180), .Z(n6177) );
  XNOR U7261 ( .A(b[3015]), .B(n6178), .Z(n6179) );
  XNOR U7262 ( .A(b[3015]), .B(n6180), .Z(c[3015]) );
  XNOR U7263 ( .A(a[3015]), .B(n6181), .Z(n6180) );
  IV U7264 ( .A(n6178), .Z(n6181) );
  XOR U7265 ( .A(n6182), .B(n6183), .Z(n6178) );
  ANDN U7266 ( .B(n6184), .A(n6185), .Z(n6182) );
  XNOR U7267 ( .A(b[3014]), .B(n6183), .Z(n6184) );
  XNOR U7268 ( .A(b[3014]), .B(n6185), .Z(c[3014]) );
  XNOR U7269 ( .A(a[3014]), .B(n6186), .Z(n6185) );
  IV U7270 ( .A(n6183), .Z(n6186) );
  XOR U7271 ( .A(n6187), .B(n6188), .Z(n6183) );
  ANDN U7272 ( .B(n6189), .A(n6190), .Z(n6187) );
  XNOR U7273 ( .A(b[3013]), .B(n6188), .Z(n6189) );
  XNOR U7274 ( .A(b[3013]), .B(n6190), .Z(c[3013]) );
  XNOR U7275 ( .A(a[3013]), .B(n6191), .Z(n6190) );
  IV U7276 ( .A(n6188), .Z(n6191) );
  XOR U7277 ( .A(n6192), .B(n6193), .Z(n6188) );
  ANDN U7278 ( .B(n6194), .A(n6195), .Z(n6192) );
  XNOR U7279 ( .A(b[3012]), .B(n6193), .Z(n6194) );
  XNOR U7280 ( .A(b[3012]), .B(n6195), .Z(c[3012]) );
  XNOR U7281 ( .A(a[3012]), .B(n6196), .Z(n6195) );
  IV U7282 ( .A(n6193), .Z(n6196) );
  XOR U7283 ( .A(n6197), .B(n6198), .Z(n6193) );
  ANDN U7284 ( .B(n6199), .A(n6200), .Z(n6197) );
  XNOR U7285 ( .A(b[3011]), .B(n6198), .Z(n6199) );
  XNOR U7286 ( .A(b[3011]), .B(n6200), .Z(c[3011]) );
  XNOR U7287 ( .A(a[3011]), .B(n6201), .Z(n6200) );
  IV U7288 ( .A(n6198), .Z(n6201) );
  XOR U7289 ( .A(n6202), .B(n6203), .Z(n6198) );
  ANDN U7290 ( .B(n6204), .A(n6205), .Z(n6202) );
  XNOR U7291 ( .A(b[3010]), .B(n6203), .Z(n6204) );
  XNOR U7292 ( .A(b[3010]), .B(n6205), .Z(c[3010]) );
  XNOR U7293 ( .A(a[3010]), .B(n6206), .Z(n6205) );
  IV U7294 ( .A(n6203), .Z(n6206) );
  XOR U7295 ( .A(n6207), .B(n6208), .Z(n6203) );
  ANDN U7296 ( .B(n6209), .A(n6210), .Z(n6207) );
  XNOR U7297 ( .A(b[3009]), .B(n6208), .Z(n6209) );
  XNOR U7298 ( .A(b[300]), .B(n6211), .Z(c[300]) );
  XNOR U7299 ( .A(b[3009]), .B(n6210), .Z(c[3009]) );
  XNOR U7300 ( .A(a[3009]), .B(n6212), .Z(n6210) );
  IV U7301 ( .A(n6208), .Z(n6212) );
  XOR U7302 ( .A(n6213), .B(n6214), .Z(n6208) );
  ANDN U7303 ( .B(n6215), .A(n6216), .Z(n6213) );
  XNOR U7304 ( .A(b[3008]), .B(n6214), .Z(n6215) );
  XNOR U7305 ( .A(b[3008]), .B(n6216), .Z(c[3008]) );
  XNOR U7306 ( .A(a[3008]), .B(n6217), .Z(n6216) );
  IV U7307 ( .A(n6214), .Z(n6217) );
  XOR U7308 ( .A(n6218), .B(n6219), .Z(n6214) );
  ANDN U7309 ( .B(n6220), .A(n6221), .Z(n6218) );
  XNOR U7310 ( .A(b[3007]), .B(n6219), .Z(n6220) );
  XNOR U7311 ( .A(b[3007]), .B(n6221), .Z(c[3007]) );
  XNOR U7312 ( .A(a[3007]), .B(n6222), .Z(n6221) );
  IV U7313 ( .A(n6219), .Z(n6222) );
  XOR U7314 ( .A(n6223), .B(n6224), .Z(n6219) );
  ANDN U7315 ( .B(n6225), .A(n6226), .Z(n6223) );
  XNOR U7316 ( .A(b[3006]), .B(n6224), .Z(n6225) );
  XNOR U7317 ( .A(b[3006]), .B(n6226), .Z(c[3006]) );
  XNOR U7318 ( .A(a[3006]), .B(n6227), .Z(n6226) );
  IV U7319 ( .A(n6224), .Z(n6227) );
  XOR U7320 ( .A(n6228), .B(n6229), .Z(n6224) );
  ANDN U7321 ( .B(n6230), .A(n6231), .Z(n6228) );
  XNOR U7322 ( .A(b[3005]), .B(n6229), .Z(n6230) );
  XNOR U7323 ( .A(b[3005]), .B(n6231), .Z(c[3005]) );
  XNOR U7324 ( .A(a[3005]), .B(n6232), .Z(n6231) );
  IV U7325 ( .A(n6229), .Z(n6232) );
  XOR U7326 ( .A(n6233), .B(n6234), .Z(n6229) );
  ANDN U7327 ( .B(n6235), .A(n6236), .Z(n6233) );
  XNOR U7328 ( .A(b[3004]), .B(n6234), .Z(n6235) );
  XNOR U7329 ( .A(b[3004]), .B(n6236), .Z(c[3004]) );
  XNOR U7330 ( .A(a[3004]), .B(n6237), .Z(n6236) );
  IV U7331 ( .A(n6234), .Z(n6237) );
  XOR U7332 ( .A(n6238), .B(n6239), .Z(n6234) );
  ANDN U7333 ( .B(n6240), .A(n6241), .Z(n6238) );
  XNOR U7334 ( .A(b[3003]), .B(n6239), .Z(n6240) );
  XNOR U7335 ( .A(b[3003]), .B(n6241), .Z(c[3003]) );
  XNOR U7336 ( .A(a[3003]), .B(n6242), .Z(n6241) );
  IV U7337 ( .A(n6239), .Z(n6242) );
  XOR U7338 ( .A(n6243), .B(n6244), .Z(n6239) );
  ANDN U7339 ( .B(n6245), .A(n6246), .Z(n6243) );
  XNOR U7340 ( .A(b[3002]), .B(n6244), .Z(n6245) );
  XNOR U7341 ( .A(b[3002]), .B(n6246), .Z(c[3002]) );
  XNOR U7342 ( .A(a[3002]), .B(n6247), .Z(n6246) );
  IV U7343 ( .A(n6244), .Z(n6247) );
  XOR U7344 ( .A(n6248), .B(n6249), .Z(n6244) );
  ANDN U7345 ( .B(n6250), .A(n6251), .Z(n6248) );
  XNOR U7346 ( .A(b[3001]), .B(n6249), .Z(n6250) );
  XNOR U7347 ( .A(b[3001]), .B(n6251), .Z(c[3001]) );
  XNOR U7348 ( .A(a[3001]), .B(n6252), .Z(n6251) );
  IV U7349 ( .A(n6249), .Z(n6252) );
  XOR U7350 ( .A(n6253), .B(n6254), .Z(n6249) );
  ANDN U7351 ( .B(n6255), .A(n6256), .Z(n6253) );
  XNOR U7352 ( .A(b[3000]), .B(n6254), .Z(n6255) );
  XNOR U7353 ( .A(b[3000]), .B(n6256), .Z(c[3000]) );
  XNOR U7354 ( .A(a[3000]), .B(n6257), .Z(n6256) );
  IV U7355 ( .A(n6254), .Z(n6257) );
  XOR U7356 ( .A(n6258), .B(n6259), .Z(n6254) );
  ANDN U7357 ( .B(n6260), .A(n6261), .Z(n6258) );
  XNOR U7358 ( .A(b[2999]), .B(n6259), .Z(n6260) );
  XNOR U7359 ( .A(b[2]), .B(n6262), .Z(c[2]) );
  XNOR U7360 ( .A(b[29]), .B(n6263), .Z(c[29]) );
  XNOR U7361 ( .A(b[299]), .B(n6264), .Z(c[299]) );
  XNOR U7362 ( .A(b[2999]), .B(n6261), .Z(c[2999]) );
  XNOR U7363 ( .A(a[2999]), .B(n6265), .Z(n6261) );
  IV U7364 ( .A(n6259), .Z(n6265) );
  XOR U7365 ( .A(n6266), .B(n6267), .Z(n6259) );
  ANDN U7366 ( .B(n6268), .A(n6269), .Z(n6266) );
  XNOR U7367 ( .A(b[2998]), .B(n6267), .Z(n6268) );
  XNOR U7368 ( .A(b[2998]), .B(n6269), .Z(c[2998]) );
  XNOR U7369 ( .A(a[2998]), .B(n6270), .Z(n6269) );
  IV U7370 ( .A(n6267), .Z(n6270) );
  XOR U7371 ( .A(n6271), .B(n6272), .Z(n6267) );
  ANDN U7372 ( .B(n6273), .A(n6274), .Z(n6271) );
  XNOR U7373 ( .A(b[2997]), .B(n6272), .Z(n6273) );
  XNOR U7374 ( .A(b[2997]), .B(n6274), .Z(c[2997]) );
  XNOR U7375 ( .A(a[2997]), .B(n6275), .Z(n6274) );
  IV U7376 ( .A(n6272), .Z(n6275) );
  XOR U7377 ( .A(n6276), .B(n6277), .Z(n6272) );
  ANDN U7378 ( .B(n6278), .A(n6279), .Z(n6276) );
  XNOR U7379 ( .A(b[2996]), .B(n6277), .Z(n6278) );
  XNOR U7380 ( .A(b[2996]), .B(n6279), .Z(c[2996]) );
  XNOR U7381 ( .A(a[2996]), .B(n6280), .Z(n6279) );
  IV U7382 ( .A(n6277), .Z(n6280) );
  XOR U7383 ( .A(n6281), .B(n6282), .Z(n6277) );
  ANDN U7384 ( .B(n6283), .A(n6284), .Z(n6281) );
  XNOR U7385 ( .A(b[2995]), .B(n6282), .Z(n6283) );
  XNOR U7386 ( .A(b[2995]), .B(n6284), .Z(c[2995]) );
  XNOR U7387 ( .A(a[2995]), .B(n6285), .Z(n6284) );
  IV U7388 ( .A(n6282), .Z(n6285) );
  XOR U7389 ( .A(n6286), .B(n6287), .Z(n6282) );
  ANDN U7390 ( .B(n6288), .A(n6289), .Z(n6286) );
  XNOR U7391 ( .A(b[2994]), .B(n6287), .Z(n6288) );
  XNOR U7392 ( .A(b[2994]), .B(n6289), .Z(c[2994]) );
  XNOR U7393 ( .A(a[2994]), .B(n6290), .Z(n6289) );
  IV U7394 ( .A(n6287), .Z(n6290) );
  XOR U7395 ( .A(n6291), .B(n6292), .Z(n6287) );
  ANDN U7396 ( .B(n6293), .A(n6294), .Z(n6291) );
  XNOR U7397 ( .A(b[2993]), .B(n6292), .Z(n6293) );
  XNOR U7398 ( .A(b[2993]), .B(n6294), .Z(c[2993]) );
  XNOR U7399 ( .A(a[2993]), .B(n6295), .Z(n6294) );
  IV U7400 ( .A(n6292), .Z(n6295) );
  XOR U7401 ( .A(n6296), .B(n6297), .Z(n6292) );
  ANDN U7402 ( .B(n6298), .A(n6299), .Z(n6296) );
  XNOR U7403 ( .A(b[2992]), .B(n6297), .Z(n6298) );
  XNOR U7404 ( .A(b[2992]), .B(n6299), .Z(c[2992]) );
  XNOR U7405 ( .A(a[2992]), .B(n6300), .Z(n6299) );
  IV U7406 ( .A(n6297), .Z(n6300) );
  XOR U7407 ( .A(n6301), .B(n6302), .Z(n6297) );
  ANDN U7408 ( .B(n6303), .A(n6304), .Z(n6301) );
  XNOR U7409 ( .A(b[2991]), .B(n6302), .Z(n6303) );
  XNOR U7410 ( .A(b[2991]), .B(n6304), .Z(c[2991]) );
  XNOR U7411 ( .A(a[2991]), .B(n6305), .Z(n6304) );
  IV U7412 ( .A(n6302), .Z(n6305) );
  XOR U7413 ( .A(n6306), .B(n6307), .Z(n6302) );
  ANDN U7414 ( .B(n6308), .A(n6309), .Z(n6306) );
  XNOR U7415 ( .A(b[2990]), .B(n6307), .Z(n6308) );
  XNOR U7416 ( .A(b[2990]), .B(n6309), .Z(c[2990]) );
  XNOR U7417 ( .A(a[2990]), .B(n6310), .Z(n6309) );
  IV U7418 ( .A(n6307), .Z(n6310) );
  XOR U7419 ( .A(n6311), .B(n6312), .Z(n6307) );
  ANDN U7420 ( .B(n6313), .A(n6314), .Z(n6311) );
  XNOR U7421 ( .A(b[2989]), .B(n6312), .Z(n6313) );
  XNOR U7422 ( .A(b[298]), .B(n6315), .Z(c[298]) );
  XNOR U7423 ( .A(b[2989]), .B(n6314), .Z(c[2989]) );
  XNOR U7424 ( .A(a[2989]), .B(n6316), .Z(n6314) );
  IV U7425 ( .A(n6312), .Z(n6316) );
  XOR U7426 ( .A(n6317), .B(n6318), .Z(n6312) );
  ANDN U7427 ( .B(n6319), .A(n6320), .Z(n6317) );
  XNOR U7428 ( .A(b[2988]), .B(n6318), .Z(n6319) );
  XNOR U7429 ( .A(b[2988]), .B(n6320), .Z(c[2988]) );
  XNOR U7430 ( .A(a[2988]), .B(n6321), .Z(n6320) );
  IV U7431 ( .A(n6318), .Z(n6321) );
  XOR U7432 ( .A(n6322), .B(n6323), .Z(n6318) );
  ANDN U7433 ( .B(n6324), .A(n6325), .Z(n6322) );
  XNOR U7434 ( .A(b[2987]), .B(n6323), .Z(n6324) );
  XNOR U7435 ( .A(b[2987]), .B(n6325), .Z(c[2987]) );
  XNOR U7436 ( .A(a[2987]), .B(n6326), .Z(n6325) );
  IV U7437 ( .A(n6323), .Z(n6326) );
  XOR U7438 ( .A(n6327), .B(n6328), .Z(n6323) );
  ANDN U7439 ( .B(n6329), .A(n6330), .Z(n6327) );
  XNOR U7440 ( .A(b[2986]), .B(n6328), .Z(n6329) );
  XNOR U7441 ( .A(b[2986]), .B(n6330), .Z(c[2986]) );
  XNOR U7442 ( .A(a[2986]), .B(n6331), .Z(n6330) );
  IV U7443 ( .A(n6328), .Z(n6331) );
  XOR U7444 ( .A(n6332), .B(n6333), .Z(n6328) );
  ANDN U7445 ( .B(n6334), .A(n6335), .Z(n6332) );
  XNOR U7446 ( .A(b[2985]), .B(n6333), .Z(n6334) );
  XNOR U7447 ( .A(b[2985]), .B(n6335), .Z(c[2985]) );
  XNOR U7448 ( .A(a[2985]), .B(n6336), .Z(n6335) );
  IV U7449 ( .A(n6333), .Z(n6336) );
  XOR U7450 ( .A(n6337), .B(n6338), .Z(n6333) );
  ANDN U7451 ( .B(n6339), .A(n6340), .Z(n6337) );
  XNOR U7452 ( .A(b[2984]), .B(n6338), .Z(n6339) );
  XNOR U7453 ( .A(b[2984]), .B(n6340), .Z(c[2984]) );
  XNOR U7454 ( .A(a[2984]), .B(n6341), .Z(n6340) );
  IV U7455 ( .A(n6338), .Z(n6341) );
  XOR U7456 ( .A(n6342), .B(n6343), .Z(n6338) );
  ANDN U7457 ( .B(n6344), .A(n6345), .Z(n6342) );
  XNOR U7458 ( .A(b[2983]), .B(n6343), .Z(n6344) );
  XNOR U7459 ( .A(b[2983]), .B(n6345), .Z(c[2983]) );
  XNOR U7460 ( .A(a[2983]), .B(n6346), .Z(n6345) );
  IV U7461 ( .A(n6343), .Z(n6346) );
  XOR U7462 ( .A(n6347), .B(n6348), .Z(n6343) );
  ANDN U7463 ( .B(n6349), .A(n6350), .Z(n6347) );
  XNOR U7464 ( .A(b[2982]), .B(n6348), .Z(n6349) );
  XNOR U7465 ( .A(b[2982]), .B(n6350), .Z(c[2982]) );
  XNOR U7466 ( .A(a[2982]), .B(n6351), .Z(n6350) );
  IV U7467 ( .A(n6348), .Z(n6351) );
  XOR U7468 ( .A(n6352), .B(n6353), .Z(n6348) );
  ANDN U7469 ( .B(n6354), .A(n6355), .Z(n6352) );
  XNOR U7470 ( .A(b[2981]), .B(n6353), .Z(n6354) );
  XNOR U7471 ( .A(b[2981]), .B(n6355), .Z(c[2981]) );
  XNOR U7472 ( .A(a[2981]), .B(n6356), .Z(n6355) );
  IV U7473 ( .A(n6353), .Z(n6356) );
  XOR U7474 ( .A(n6357), .B(n6358), .Z(n6353) );
  ANDN U7475 ( .B(n6359), .A(n6360), .Z(n6357) );
  XNOR U7476 ( .A(b[2980]), .B(n6358), .Z(n6359) );
  XNOR U7477 ( .A(b[2980]), .B(n6360), .Z(c[2980]) );
  XNOR U7478 ( .A(a[2980]), .B(n6361), .Z(n6360) );
  IV U7479 ( .A(n6358), .Z(n6361) );
  XOR U7480 ( .A(n6362), .B(n6363), .Z(n6358) );
  ANDN U7481 ( .B(n6364), .A(n6365), .Z(n6362) );
  XNOR U7482 ( .A(b[2979]), .B(n6363), .Z(n6364) );
  XNOR U7483 ( .A(b[297]), .B(n6366), .Z(c[297]) );
  XNOR U7484 ( .A(b[2979]), .B(n6365), .Z(c[2979]) );
  XNOR U7485 ( .A(a[2979]), .B(n6367), .Z(n6365) );
  IV U7486 ( .A(n6363), .Z(n6367) );
  XOR U7487 ( .A(n6368), .B(n6369), .Z(n6363) );
  ANDN U7488 ( .B(n6370), .A(n6371), .Z(n6368) );
  XNOR U7489 ( .A(b[2978]), .B(n6369), .Z(n6370) );
  XNOR U7490 ( .A(b[2978]), .B(n6371), .Z(c[2978]) );
  XNOR U7491 ( .A(a[2978]), .B(n6372), .Z(n6371) );
  IV U7492 ( .A(n6369), .Z(n6372) );
  XOR U7493 ( .A(n6373), .B(n6374), .Z(n6369) );
  ANDN U7494 ( .B(n6375), .A(n6376), .Z(n6373) );
  XNOR U7495 ( .A(b[2977]), .B(n6374), .Z(n6375) );
  XNOR U7496 ( .A(b[2977]), .B(n6376), .Z(c[2977]) );
  XNOR U7497 ( .A(a[2977]), .B(n6377), .Z(n6376) );
  IV U7498 ( .A(n6374), .Z(n6377) );
  XOR U7499 ( .A(n6378), .B(n6379), .Z(n6374) );
  ANDN U7500 ( .B(n6380), .A(n6381), .Z(n6378) );
  XNOR U7501 ( .A(b[2976]), .B(n6379), .Z(n6380) );
  XNOR U7502 ( .A(b[2976]), .B(n6381), .Z(c[2976]) );
  XNOR U7503 ( .A(a[2976]), .B(n6382), .Z(n6381) );
  IV U7504 ( .A(n6379), .Z(n6382) );
  XOR U7505 ( .A(n6383), .B(n6384), .Z(n6379) );
  ANDN U7506 ( .B(n6385), .A(n6386), .Z(n6383) );
  XNOR U7507 ( .A(b[2975]), .B(n6384), .Z(n6385) );
  XNOR U7508 ( .A(b[2975]), .B(n6386), .Z(c[2975]) );
  XNOR U7509 ( .A(a[2975]), .B(n6387), .Z(n6386) );
  IV U7510 ( .A(n6384), .Z(n6387) );
  XOR U7511 ( .A(n6388), .B(n6389), .Z(n6384) );
  ANDN U7512 ( .B(n6390), .A(n6391), .Z(n6388) );
  XNOR U7513 ( .A(b[2974]), .B(n6389), .Z(n6390) );
  XNOR U7514 ( .A(b[2974]), .B(n6391), .Z(c[2974]) );
  XNOR U7515 ( .A(a[2974]), .B(n6392), .Z(n6391) );
  IV U7516 ( .A(n6389), .Z(n6392) );
  XOR U7517 ( .A(n6393), .B(n6394), .Z(n6389) );
  ANDN U7518 ( .B(n6395), .A(n6396), .Z(n6393) );
  XNOR U7519 ( .A(b[2973]), .B(n6394), .Z(n6395) );
  XNOR U7520 ( .A(b[2973]), .B(n6396), .Z(c[2973]) );
  XNOR U7521 ( .A(a[2973]), .B(n6397), .Z(n6396) );
  IV U7522 ( .A(n6394), .Z(n6397) );
  XOR U7523 ( .A(n6398), .B(n6399), .Z(n6394) );
  ANDN U7524 ( .B(n6400), .A(n6401), .Z(n6398) );
  XNOR U7525 ( .A(b[2972]), .B(n6399), .Z(n6400) );
  XNOR U7526 ( .A(b[2972]), .B(n6401), .Z(c[2972]) );
  XNOR U7527 ( .A(a[2972]), .B(n6402), .Z(n6401) );
  IV U7528 ( .A(n6399), .Z(n6402) );
  XOR U7529 ( .A(n6403), .B(n6404), .Z(n6399) );
  ANDN U7530 ( .B(n6405), .A(n6406), .Z(n6403) );
  XNOR U7531 ( .A(b[2971]), .B(n6404), .Z(n6405) );
  XNOR U7532 ( .A(b[2971]), .B(n6406), .Z(c[2971]) );
  XNOR U7533 ( .A(a[2971]), .B(n6407), .Z(n6406) );
  IV U7534 ( .A(n6404), .Z(n6407) );
  XOR U7535 ( .A(n6408), .B(n6409), .Z(n6404) );
  ANDN U7536 ( .B(n6410), .A(n6411), .Z(n6408) );
  XNOR U7537 ( .A(b[2970]), .B(n6409), .Z(n6410) );
  XNOR U7538 ( .A(b[2970]), .B(n6411), .Z(c[2970]) );
  XNOR U7539 ( .A(a[2970]), .B(n6412), .Z(n6411) );
  IV U7540 ( .A(n6409), .Z(n6412) );
  XOR U7541 ( .A(n6413), .B(n6414), .Z(n6409) );
  ANDN U7542 ( .B(n6415), .A(n6416), .Z(n6413) );
  XNOR U7543 ( .A(b[2969]), .B(n6414), .Z(n6415) );
  XNOR U7544 ( .A(b[296]), .B(n6417), .Z(c[296]) );
  XNOR U7545 ( .A(b[2969]), .B(n6416), .Z(c[2969]) );
  XNOR U7546 ( .A(a[2969]), .B(n6418), .Z(n6416) );
  IV U7547 ( .A(n6414), .Z(n6418) );
  XOR U7548 ( .A(n6419), .B(n6420), .Z(n6414) );
  ANDN U7549 ( .B(n6421), .A(n6422), .Z(n6419) );
  XNOR U7550 ( .A(b[2968]), .B(n6420), .Z(n6421) );
  XNOR U7551 ( .A(b[2968]), .B(n6422), .Z(c[2968]) );
  XNOR U7552 ( .A(a[2968]), .B(n6423), .Z(n6422) );
  IV U7553 ( .A(n6420), .Z(n6423) );
  XOR U7554 ( .A(n6424), .B(n6425), .Z(n6420) );
  ANDN U7555 ( .B(n6426), .A(n6427), .Z(n6424) );
  XNOR U7556 ( .A(b[2967]), .B(n6425), .Z(n6426) );
  XNOR U7557 ( .A(b[2967]), .B(n6427), .Z(c[2967]) );
  XNOR U7558 ( .A(a[2967]), .B(n6428), .Z(n6427) );
  IV U7559 ( .A(n6425), .Z(n6428) );
  XOR U7560 ( .A(n6429), .B(n6430), .Z(n6425) );
  ANDN U7561 ( .B(n6431), .A(n6432), .Z(n6429) );
  XNOR U7562 ( .A(b[2966]), .B(n6430), .Z(n6431) );
  XNOR U7563 ( .A(b[2966]), .B(n6432), .Z(c[2966]) );
  XNOR U7564 ( .A(a[2966]), .B(n6433), .Z(n6432) );
  IV U7565 ( .A(n6430), .Z(n6433) );
  XOR U7566 ( .A(n6434), .B(n6435), .Z(n6430) );
  ANDN U7567 ( .B(n6436), .A(n6437), .Z(n6434) );
  XNOR U7568 ( .A(b[2965]), .B(n6435), .Z(n6436) );
  XNOR U7569 ( .A(b[2965]), .B(n6437), .Z(c[2965]) );
  XNOR U7570 ( .A(a[2965]), .B(n6438), .Z(n6437) );
  IV U7571 ( .A(n6435), .Z(n6438) );
  XOR U7572 ( .A(n6439), .B(n6440), .Z(n6435) );
  ANDN U7573 ( .B(n6441), .A(n6442), .Z(n6439) );
  XNOR U7574 ( .A(b[2964]), .B(n6440), .Z(n6441) );
  XNOR U7575 ( .A(b[2964]), .B(n6442), .Z(c[2964]) );
  XNOR U7576 ( .A(a[2964]), .B(n6443), .Z(n6442) );
  IV U7577 ( .A(n6440), .Z(n6443) );
  XOR U7578 ( .A(n6444), .B(n6445), .Z(n6440) );
  ANDN U7579 ( .B(n6446), .A(n6447), .Z(n6444) );
  XNOR U7580 ( .A(b[2963]), .B(n6445), .Z(n6446) );
  XNOR U7581 ( .A(b[2963]), .B(n6447), .Z(c[2963]) );
  XNOR U7582 ( .A(a[2963]), .B(n6448), .Z(n6447) );
  IV U7583 ( .A(n6445), .Z(n6448) );
  XOR U7584 ( .A(n6449), .B(n6450), .Z(n6445) );
  ANDN U7585 ( .B(n6451), .A(n6452), .Z(n6449) );
  XNOR U7586 ( .A(b[2962]), .B(n6450), .Z(n6451) );
  XNOR U7587 ( .A(b[2962]), .B(n6452), .Z(c[2962]) );
  XNOR U7588 ( .A(a[2962]), .B(n6453), .Z(n6452) );
  IV U7589 ( .A(n6450), .Z(n6453) );
  XOR U7590 ( .A(n6454), .B(n6455), .Z(n6450) );
  ANDN U7591 ( .B(n6456), .A(n6457), .Z(n6454) );
  XNOR U7592 ( .A(b[2961]), .B(n6455), .Z(n6456) );
  XNOR U7593 ( .A(b[2961]), .B(n6457), .Z(c[2961]) );
  XNOR U7594 ( .A(a[2961]), .B(n6458), .Z(n6457) );
  IV U7595 ( .A(n6455), .Z(n6458) );
  XOR U7596 ( .A(n6459), .B(n6460), .Z(n6455) );
  ANDN U7597 ( .B(n6461), .A(n6462), .Z(n6459) );
  XNOR U7598 ( .A(b[2960]), .B(n6460), .Z(n6461) );
  XNOR U7599 ( .A(b[2960]), .B(n6462), .Z(c[2960]) );
  XNOR U7600 ( .A(a[2960]), .B(n6463), .Z(n6462) );
  IV U7601 ( .A(n6460), .Z(n6463) );
  XOR U7602 ( .A(n6464), .B(n6465), .Z(n6460) );
  ANDN U7603 ( .B(n6466), .A(n6467), .Z(n6464) );
  XNOR U7604 ( .A(b[2959]), .B(n6465), .Z(n6466) );
  XNOR U7605 ( .A(b[295]), .B(n6468), .Z(c[295]) );
  XNOR U7606 ( .A(b[2959]), .B(n6467), .Z(c[2959]) );
  XNOR U7607 ( .A(a[2959]), .B(n6469), .Z(n6467) );
  IV U7608 ( .A(n6465), .Z(n6469) );
  XOR U7609 ( .A(n6470), .B(n6471), .Z(n6465) );
  ANDN U7610 ( .B(n6472), .A(n6473), .Z(n6470) );
  XNOR U7611 ( .A(b[2958]), .B(n6471), .Z(n6472) );
  XNOR U7612 ( .A(b[2958]), .B(n6473), .Z(c[2958]) );
  XNOR U7613 ( .A(a[2958]), .B(n6474), .Z(n6473) );
  IV U7614 ( .A(n6471), .Z(n6474) );
  XOR U7615 ( .A(n6475), .B(n6476), .Z(n6471) );
  ANDN U7616 ( .B(n6477), .A(n6478), .Z(n6475) );
  XNOR U7617 ( .A(b[2957]), .B(n6476), .Z(n6477) );
  XNOR U7618 ( .A(b[2957]), .B(n6478), .Z(c[2957]) );
  XNOR U7619 ( .A(a[2957]), .B(n6479), .Z(n6478) );
  IV U7620 ( .A(n6476), .Z(n6479) );
  XOR U7621 ( .A(n6480), .B(n6481), .Z(n6476) );
  ANDN U7622 ( .B(n6482), .A(n6483), .Z(n6480) );
  XNOR U7623 ( .A(b[2956]), .B(n6481), .Z(n6482) );
  XNOR U7624 ( .A(b[2956]), .B(n6483), .Z(c[2956]) );
  XNOR U7625 ( .A(a[2956]), .B(n6484), .Z(n6483) );
  IV U7626 ( .A(n6481), .Z(n6484) );
  XOR U7627 ( .A(n6485), .B(n6486), .Z(n6481) );
  ANDN U7628 ( .B(n6487), .A(n6488), .Z(n6485) );
  XNOR U7629 ( .A(b[2955]), .B(n6486), .Z(n6487) );
  XNOR U7630 ( .A(b[2955]), .B(n6488), .Z(c[2955]) );
  XNOR U7631 ( .A(a[2955]), .B(n6489), .Z(n6488) );
  IV U7632 ( .A(n6486), .Z(n6489) );
  XOR U7633 ( .A(n6490), .B(n6491), .Z(n6486) );
  ANDN U7634 ( .B(n6492), .A(n6493), .Z(n6490) );
  XNOR U7635 ( .A(b[2954]), .B(n6491), .Z(n6492) );
  XNOR U7636 ( .A(b[2954]), .B(n6493), .Z(c[2954]) );
  XNOR U7637 ( .A(a[2954]), .B(n6494), .Z(n6493) );
  IV U7638 ( .A(n6491), .Z(n6494) );
  XOR U7639 ( .A(n6495), .B(n6496), .Z(n6491) );
  ANDN U7640 ( .B(n6497), .A(n6498), .Z(n6495) );
  XNOR U7641 ( .A(b[2953]), .B(n6496), .Z(n6497) );
  XNOR U7642 ( .A(b[2953]), .B(n6498), .Z(c[2953]) );
  XNOR U7643 ( .A(a[2953]), .B(n6499), .Z(n6498) );
  IV U7644 ( .A(n6496), .Z(n6499) );
  XOR U7645 ( .A(n6500), .B(n6501), .Z(n6496) );
  ANDN U7646 ( .B(n6502), .A(n6503), .Z(n6500) );
  XNOR U7647 ( .A(b[2952]), .B(n6501), .Z(n6502) );
  XNOR U7648 ( .A(b[2952]), .B(n6503), .Z(c[2952]) );
  XNOR U7649 ( .A(a[2952]), .B(n6504), .Z(n6503) );
  IV U7650 ( .A(n6501), .Z(n6504) );
  XOR U7651 ( .A(n6505), .B(n6506), .Z(n6501) );
  ANDN U7652 ( .B(n6507), .A(n6508), .Z(n6505) );
  XNOR U7653 ( .A(b[2951]), .B(n6506), .Z(n6507) );
  XNOR U7654 ( .A(b[2951]), .B(n6508), .Z(c[2951]) );
  XNOR U7655 ( .A(a[2951]), .B(n6509), .Z(n6508) );
  IV U7656 ( .A(n6506), .Z(n6509) );
  XOR U7657 ( .A(n6510), .B(n6511), .Z(n6506) );
  ANDN U7658 ( .B(n6512), .A(n6513), .Z(n6510) );
  XNOR U7659 ( .A(b[2950]), .B(n6511), .Z(n6512) );
  XNOR U7660 ( .A(b[2950]), .B(n6513), .Z(c[2950]) );
  XNOR U7661 ( .A(a[2950]), .B(n6514), .Z(n6513) );
  IV U7662 ( .A(n6511), .Z(n6514) );
  XOR U7663 ( .A(n6515), .B(n6516), .Z(n6511) );
  ANDN U7664 ( .B(n6517), .A(n6518), .Z(n6515) );
  XNOR U7665 ( .A(b[2949]), .B(n6516), .Z(n6517) );
  XNOR U7666 ( .A(b[294]), .B(n6519), .Z(c[294]) );
  XNOR U7667 ( .A(b[2949]), .B(n6518), .Z(c[2949]) );
  XNOR U7668 ( .A(a[2949]), .B(n6520), .Z(n6518) );
  IV U7669 ( .A(n6516), .Z(n6520) );
  XOR U7670 ( .A(n6521), .B(n6522), .Z(n6516) );
  ANDN U7671 ( .B(n6523), .A(n6524), .Z(n6521) );
  XNOR U7672 ( .A(b[2948]), .B(n6522), .Z(n6523) );
  XNOR U7673 ( .A(b[2948]), .B(n6524), .Z(c[2948]) );
  XNOR U7674 ( .A(a[2948]), .B(n6525), .Z(n6524) );
  IV U7675 ( .A(n6522), .Z(n6525) );
  XOR U7676 ( .A(n6526), .B(n6527), .Z(n6522) );
  ANDN U7677 ( .B(n6528), .A(n6529), .Z(n6526) );
  XNOR U7678 ( .A(b[2947]), .B(n6527), .Z(n6528) );
  XNOR U7679 ( .A(b[2947]), .B(n6529), .Z(c[2947]) );
  XNOR U7680 ( .A(a[2947]), .B(n6530), .Z(n6529) );
  IV U7681 ( .A(n6527), .Z(n6530) );
  XOR U7682 ( .A(n6531), .B(n6532), .Z(n6527) );
  ANDN U7683 ( .B(n6533), .A(n6534), .Z(n6531) );
  XNOR U7684 ( .A(b[2946]), .B(n6532), .Z(n6533) );
  XNOR U7685 ( .A(b[2946]), .B(n6534), .Z(c[2946]) );
  XNOR U7686 ( .A(a[2946]), .B(n6535), .Z(n6534) );
  IV U7687 ( .A(n6532), .Z(n6535) );
  XOR U7688 ( .A(n6536), .B(n6537), .Z(n6532) );
  ANDN U7689 ( .B(n6538), .A(n6539), .Z(n6536) );
  XNOR U7690 ( .A(b[2945]), .B(n6537), .Z(n6538) );
  XNOR U7691 ( .A(b[2945]), .B(n6539), .Z(c[2945]) );
  XNOR U7692 ( .A(a[2945]), .B(n6540), .Z(n6539) );
  IV U7693 ( .A(n6537), .Z(n6540) );
  XOR U7694 ( .A(n6541), .B(n6542), .Z(n6537) );
  ANDN U7695 ( .B(n6543), .A(n6544), .Z(n6541) );
  XNOR U7696 ( .A(b[2944]), .B(n6542), .Z(n6543) );
  XNOR U7697 ( .A(b[2944]), .B(n6544), .Z(c[2944]) );
  XNOR U7698 ( .A(a[2944]), .B(n6545), .Z(n6544) );
  IV U7699 ( .A(n6542), .Z(n6545) );
  XOR U7700 ( .A(n6546), .B(n6547), .Z(n6542) );
  ANDN U7701 ( .B(n6548), .A(n6549), .Z(n6546) );
  XNOR U7702 ( .A(b[2943]), .B(n6547), .Z(n6548) );
  XNOR U7703 ( .A(b[2943]), .B(n6549), .Z(c[2943]) );
  XNOR U7704 ( .A(a[2943]), .B(n6550), .Z(n6549) );
  IV U7705 ( .A(n6547), .Z(n6550) );
  XOR U7706 ( .A(n6551), .B(n6552), .Z(n6547) );
  ANDN U7707 ( .B(n6553), .A(n6554), .Z(n6551) );
  XNOR U7708 ( .A(b[2942]), .B(n6552), .Z(n6553) );
  XNOR U7709 ( .A(b[2942]), .B(n6554), .Z(c[2942]) );
  XNOR U7710 ( .A(a[2942]), .B(n6555), .Z(n6554) );
  IV U7711 ( .A(n6552), .Z(n6555) );
  XOR U7712 ( .A(n6556), .B(n6557), .Z(n6552) );
  ANDN U7713 ( .B(n6558), .A(n6559), .Z(n6556) );
  XNOR U7714 ( .A(b[2941]), .B(n6557), .Z(n6558) );
  XNOR U7715 ( .A(b[2941]), .B(n6559), .Z(c[2941]) );
  XNOR U7716 ( .A(a[2941]), .B(n6560), .Z(n6559) );
  IV U7717 ( .A(n6557), .Z(n6560) );
  XOR U7718 ( .A(n6561), .B(n6562), .Z(n6557) );
  ANDN U7719 ( .B(n6563), .A(n6564), .Z(n6561) );
  XNOR U7720 ( .A(b[2940]), .B(n6562), .Z(n6563) );
  XNOR U7721 ( .A(b[2940]), .B(n6564), .Z(c[2940]) );
  XNOR U7722 ( .A(a[2940]), .B(n6565), .Z(n6564) );
  IV U7723 ( .A(n6562), .Z(n6565) );
  XOR U7724 ( .A(n6566), .B(n6567), .Z(n6562) );
  ANDN U7725 ( .B(n6568), .A(n6569), .Z(n6566) );
  XNOR U7726 ( .A(b[2939]), .B(n6567), .Z(n6568) );
  XNOR U7727 ( .A(b[293]), .B(n6570), .Z(c[293]) );
  XNOR U7728 ( .A(b[2939]), .B(n6569), .Z(c[2939]) );
  XNOR U7729 ( .A(a[2939]), .B(n6571), .Z(n6569) );
  IV U7730 ( .A(n6567), .Z(n6571) );
  XOR U7731 ( .A(n6572), .B(n6573), .Z(n6567) );
  ANDN U7732 ( .B(n6574), .A(n6575), .Z(n6572) );
  XNOR U7733 ( .A(b[2938]), .B(n6573), .Z(n6574) );
  XNOR U7734 ( .A(b[2938]), .B(n6575), .Z(c[2938]) );
  XNOR U7735 ( .A(a[2938]), .B(n6576), .Z(n6575) );
  IV U7736 ( .A(n6573), .Z(n6576) );
  XOR U7737 ( .A(n6577), .B(n6578), .Z(n6573) );
  ANDN U7738 ( .B(n6579), .A(n6580), .Z(n6577) );
  XNOR U7739 ( .A(b[2937]), .B(n6578), .Z(n6579) );
  XNOR U7740 ( .A(b[2937]), .B(n6580), .Z(c[2937]) );
  XNOR U7741 ( .A(a[2937]), .B(n6581), .Z(n6580) );
  IV U7742 ( .A(n6578), .Z(n6581) );
  XOR U7743 ( .A(n6582), .B(n6583), .Z(n6578) );
  ANDN U7744 ( .B(n6584), .A(n6585), .Z(n6582) );
  XNOR U7745 ( .A(b[2936]), .B(n6583), .Z(n6584) );
  XNOR U7746 ( .A(b[2936]), .B(n6585), .Z(c[2936]) );
  XNOR U7747 ( .A(a[2936]), .B(n6586), .Z(n6585) );
  IV U7748 ( .A(n6583), .Z(n6586) );
  XOR U7749 ( .A(n6587), .B(n6588), .Z(n6583) );
  ANDN U7750 ( .B(n6589), .A(n6590), .Z(n6587) );
  XNOR U7751 ( .A(b[2935]), .B(n6588), .Z(n6589) );
  XNOR U7752 ( .A(b[2935]), .B(n6590), .Z(c[2935]) );
  XNOR U7753 ( .A(a[2935]), .B(n6591), .Z(n6590) );
  IV U7754 ( .A(n6588), .Z(n6591) );
  XOR U7755 ( .A(n6592), .B(n6593), .Z(n6588) );
  ANDN U7756 ( .B(n6594), .A(n6595), .Z(n6592) );
  XNOR U7757 ( .A(b[2934]), .B(n6593), .Z(n6594) );
  XNOR U7758 ( .A(b[2934]), .B(n6595), .Z(c[2934]) );
  XNOR U7759 ( .A(a[2934]), .B(n6596), .Z(n6595) );
  IV U7760 ( .A(n6593), .Z(n6596) );
  XOR U7761 ( .A(n6597), .B(n6598), .Z(n6593) );
  ANDN U7762 ( .B(n6599), .A(n6600), .Z(n6597) );
  XNOR U7763 ( .A(b[2933]), .B(n6598), .Z(n6599) );
  XNOR U7764 ( .A(b[2933]), .B(n6600), .Z(c[2933]) );
  XNOR U7765 ( .A(a[2933]), .B(n6601), .Z(n6600) );
  IV U7766 ( .A(n6598), .Z(n6601) );
  XOR U7767 ( .A(n6602), .B(n6603), .Z(n6598) );
  ANDN U7768 ( .B(n6604), .A(n6605), .Z(n6602) );
  XNOR U7769 ( .A(b[2932]), .B(n6603), .Z(n6604) );
  XNOR U7770 ( .A(b[2932]), .B(n6605), .Z(c[2932]) );
  XNOR U7771 ( .A(a[2932]), .B(n6606), .Z(n6605) );
  IV U7772 ( .A(n6603), .Z(n6606) );
  XOR U7773 ( .A(n6607), .B(n6608), .Z(n6603) );
  ANDN U7774 ( .B(n6609), .A(n6610), .Z(n6607) );
  XNOR U7775 ( .A(b[2931]), .B(n6608), .Z(n6609) );
  XNOR U7776 ( .A(b[2931]), .B(n6610), .Z(c[2931]) );
  XNOR U7777 ( .A(a[2931]), .B(n6611), .Z(n6610) );
  IV U7778 ( .A(n6608), .Z(n6611) );
  XOR U7779 ( .A(n6612), .B(n6613), .Z(n6608) );
  ANDN U7780 ( .B(n6614), .A(n6615), .Z(n6612) );
  XNOR U7781 ( .A(b[2930]), .B(n6613), .Z(n6614) );
  XNOR U7782 ( .A(b[2930]), .B(n6615), .Z(c[2930]) );
  XNOR U7783 ( .A(a[2930]), .B(n6616), .Z(n6615) );
  IV U7784 ( .A(n6613), .Z(n6616) );
  XOR U7785 ( .A(n6617), .B(n6618), .Z(n6613) );
  ANDN U7786 ( .B(n6619), .A(n6620), .Z(n6617) );
  XNOR U7787 ( .A(b[2929]), .B(n6618), .Z(n6619) );
  XNOR U7788 ( .A(b[292]), .B(n6621), .Z(c[292]) );
  XNOR U7789 ( .A(b[2929]), .B(n6620), .Z(c[2929]) );
  XNOR U7790 ( .A(a[2929]), .B(n6622), .Z(n6620) );
  IV U7791 ( .A(n6618), .Z(n6622) );
  XOR U7792 ( .A(n6623), .B(n6624), .Z(n6618) );
  ANDN U7793 ( .B(n6625), .A(n6626), .Z(n6623) );
  XNOR U7794 ( .A(b[2928]), .B(n6624), .Z(n6625) );
  XNOR U7795 ( .A(b[2928]), .B(n6626), .Z(c[2928]) );
  XNOR U7796 ( .A(a[2928]), .B(n6627), .Z(n6626) );
  IV U7797 ( .A(n6624), .Z(n6627) );
  XOR U7798 ( .A(n6628), .B(n6629), .Z(n6624) );
  ANDN U7799 ( .B(n6630), .A(n6631), .Z(n6628) );
  XNOR U7800 ( .A(b[2927]), .B(n6629), .Z(n6630) );
  XNOR U7801 ( .A(b[2927]), .B(n6631), .Z(c[2927]) );
  XNOR U7802 ( .A(a[2927]), .B(n6632), .Z(n6631) );
  IV U7803 ( .A(n6629), .Z(n6632) );
  XOR U7804 ( .A(n6633), .B(n6634), .Z(n6629) );
  ANDN U7805 ( .B(n6635), .A(n6636), .Z(n6633) );
  XNOR U7806 ( .A(b[2926]), .B(n6634), .Z(n6635) );
  XNOR U7807 ( .A(b[2926]), .B(n6636), .Z(c[2926]) );
  XNOR U7808 ( .A(a[2926]), .B(n6637), .Z(n6636) );
  IV U7809 ( .A(n6634), .Z(n6637) );
  XOR U7810 ( .A(n6638), .B(n6639), .Z(n6634) );
  ANDN U7811 ( .B(n6640), .A(n6641), .Z(n6638) );
  XNOR U7812 ( .A(b[2925]), .B(n6639), .Z(n6640) );
  XNOR U7813 ( .A(b[2925]), .B(n6641), .Z(c[2925]) );
  XNOR U7814 ( .A(a[2925]), .B(n6642), .Z(n6641) );
  IV U7815 ( .A(n6639), .Z(n6642) );
  XOR U7816 ( .A(n6643), .B(n6644), .Z(n6639) );
  ANDN U7817 ( .B(n6645), .A(n6646), .Z(n6643) );
  XNOR U7818 ( .A(b[2924]), .B(n6644), .Z(n6645) );
  XNOR U7819 ( .A(b[2924]), .B(n6646), .Z(c[2924]) );
  XNOR U7820 ( .A(a[2924]), .B(n6647), .Z(n6646) );
  IV U7821 ( .A(n6644), .Z(n6647) );
  XOR U7822 ( .A(n6648), .B(n6649), .Z(n6644) );
  ANDN U7823 ( .B(n6650), .A(n6651), .Z(n6648) );
  XNOR U7824 ( .A(b[2923]), .B(n6649), .Z(n6650) );
  XNOR U7825 ( .A(b[2923]), .B(n6651), .Z(c[2923]) );
  XNOR U7826 ( .A(a[2923]), .B(n6652), .Z(n6651) );
  IV U7827 ( .A(n6649), .Z(n6652) );
  XOR U7828 ( .A(n6653), .B(n6654), .Z(n6649) );
  ANDN U7829 ( .B(n6655), .A(n6656), .Z(n6653) );
  XNOR U7830 ( .A(b[2922]), .B(n6654), .Z(n6655) );
  XNOR U7831 ( .A(b[2922]), .B(n6656), .Z(c[2922]) );
  XNOR U7832 ( .A(a[2922]), .B(n6657), .Z(n6656) );
  IV U7833 ( .A(n6654), .Z(n6657) );
  XOR U7834 ( .A(n6658), .B(n6659), .Z(n6654) );
  ANDN U7835 ( .B(n6660), .A(n6661), .Z(n6658) );
  XNOR U7836 ( .A(b[2921]), .B(n6659), .Z(n6660) );
  XNOR U7837 ( .A(b[2921]), .B(n6661), .Z(c[2921]) );
  XNOR U7838 ( .A(a[2921]), .B(n6662), .Z(n6661) );
  IV U7839 ( .A(n6659), .Z(n6662) );
  XOR U7840 ( .A(n6663), .B(n6664), .Z(n6659) );
  ANDN U7841 ( .B(n6665), .A(n6666), .Z(n6663) );
  XNOR U7842 ( .A(b[2920]), .B(n6664), .Z(n6665) );
  XNOR U7843 ( .A(b[2920]), .B(n6666), .Z(c[2920]) );
  XNOR U7844 ( .A(a[2920]), .B(n6667), .Z(n6666) );
  IV U7845 ( .A(n6664), .Z(n6667) );
  XOR U7846 ( .A(n6668), .B(n6669), .Z(n6664) );
  ANDN U7847 ( .B(n6670), .A(n6671), .Z(n6668) );
  XNOR U7848 ( .A(b[2919]), .B(n6669), .Z(n6670) );
  XNOR U7849 ( .A(b[291]), .B(n6672), .Z(c[291]) );
  XNOR U7850 ( .A(b[2919]), .B(n6671), .Z(c[2919]) );
  XNOR U7851 ( .A(a[2919]), .B(n6673), .Z(n6671) );
  IV U7852 ( .A(n6669), .Z(n6673) );
  XOR U7853 ( .A(n6674), .B(n6675), .Z(n6669) );
  ANDN U7854 ( .B(n6676), .A(n6677), .Z(n6674) );
  XNOR U7855 ( .A(b[2918]), .B(n6675), .Z(n6676) );
  XNOR U7856 ( .A(b[2918]), .B(n6677), .Z(c[2918]) );
  XNOR U7857 ( .A(a[2918]), .B(n6678), .Z(n6677) );
  IV U7858 ( .A(n6675), .Z(n6678) );
  XOR U7859 ( .A(n6679), .B(n6680), .Z(n6675) );
  ANDN U7860 ( .B(n6681), .A(n6682), .Z(n6679) );
  XNOR U7861 ( .A(b[2917]), .B(n6680), .Z(n6681) );
  XNOR U7862 ( .A(b[2917]), .B(n6682), .Z(c[2917]) );
  XNOR U7863 ( .A(a[2917]), .B(n6683), .Z(n6682) );
  IV U7864 ( .A(n6680), .Z(n6683) );
  XOR U7865 ( .A(n6684), .B(n6685), .Z(n6680) );
  ANDN U7866 ( .B(n6686), .A(n6687), .Z(n6684) );
  XNOR U7867 ( .A(b[2916]), .B(n6685), .Z(n6686) );
  XNOR U7868 ( .A(b[2916]), .B(n6687), .Z(c[2916]) );
  XNOR U7869 ( .A(a[2916]), .B(n6688), .Z(n6687) );
  IV U7870 ( .A(n6685), .Z(n6688) );
  XOR U7871 ( .A(n6689), .B(n6690), .Z(n6685) );
  ANDN U7872 ( .B(n6691), .A(n6692), .Z(n6689) );
  XNOR U7873 ( .A(b[2915]), .B(n6690), .Z(n6691) );
  XNOR U7874 ( .A(b[2915]), .B(n6692), .Z(c[2915]) );
  XNOR U7875 ( .A(a[2915]), .B(n6693), .Z(n6692) );
  IV U7876 ( .A(n6690), .Z(n6693) );
  XOR U7877 ( .A(n6694), .B(n6695), .Z(n6690) );
  ANDN U7878 ( .B(n6696), .A(n6697), .Z(n6694) );
  XNOR U7879 ( .A(b[2914]), .B(n6695), .Z(n6696) );
  XNOR U7880 ( .A(b[2914]), .B(n6697), .Z(c[2914]) );
  XNOR U7881 ( .A(a[2914]), .B(n6698), .Z(n6697) );
  IV U7882 ( .A(n6695), .Z(n6698) );
  XOR U7883 ( .A(n6699), .B(n6700), .Z(n6695) );
  ANDN U7884 ( .B(n6701), .A(n6702), .Z(n6699) );
  XNOR U7885 ( .A(b[2913]), .B(n6700), .Z(n6701) );
  XNOR U7886 ( .A(b[2913]), .B(n6702), .Z(c[2913]) );
  XNOR U7887 ( .A(a[2913]), .B(n6703), .Z(n6702) );
  IV U7888 ( .A(n6700), .Z(n6703) );
  XOR U7889 ( .A(n6704), .B(n6705), .Z(n6700) );
  ANDN U7890 ( .B(n6706), .A(n6707), .Z(n6704) );
  XNOR U7891 ( .A(b[2912]), .B(n6705), .Z(n6706) );
  XNOR U7892 ( .A(b[2912]), .B(n6707), .Z(c[2912]) );
  XNOR U7893 ( .A(a[2912]), .B(n6708), .Z(n6707) );
  IV U7894 ( .A(n6705), .Z(n6708) );
  XOR U7895 ( .A(n6709), .B(n6710), .Z(n6705) );
  ANDN U7896 ( .B(n6711), .A(n6712), .Z(n6709) );
  XNOR U7897 ( .A(b[2911]), .B(n6710), .Z(n6711) );
  XNOR U7898 ( .A(b[2911]), .B(n6712), .Z(c[2911]) );
  XNOR U7899 ( .A(a[2911]), .B(n6713), .Z(n6712) );
  IV U7900 ( .A(n6710), .Z(n6713) );
  XOR U7901 ( .A(n6714), .B(n6715), .Z(n6710) );
  ANDN U7902 ( .B(n6716), .A(n6717), .Z(n6714) );
  XNOR U7903 ( .A(b[2910]), .B(n6715), .Z(n6716) );
  XNOR U7904 ( .A(b[2910]), .B(n6717), .Z(c[2910]) );
  XNOR U7905 ( .A(a[2910]), .B(n6718), .Z(n6717) );
  IV U7906 ( .A(n6715), .Z(n6718) );
  XOR U7907 ( .A(n6719), .B(n6720), .Z(n6715) );
  ANDN U7908 ( .B(n6721), .A(n6722), .Z(n6719) );
  XNOR U7909 ( .A(b[2909]), .B(n6720), .Z(n6721) );
  XNOR U7910 ( .A(b[290]), .B(n6723), .Z(c[290]) );
  XNOR U7911 ( .A(b[2909]), .B(n6722), .Z(c[2909]) );
  XNOR U7912 ( .A(a[2909]), .B(n6724), .Z(n6722) );
  IV U7913 ( .A(n6720), .Z(n6724) );
  XOR U7914 ( .A(n6725), .B(n6726), .Z(n6720) );
  ANDN U7915 ( .B(n6727), .A(n6728), .Z(n6725) );
  XNOR U7916 ( .A(b[2908]), .B(n6726), .Z(n6727) );
  XNOR U7917 ( .A(b[2908]), .B(n6728), .Z(c[2908]) );
  XNOR U7918 ( .A(a[2908]), .B(n6729), .Z(n6728) );
  IV U7919 ( .A(n6726), .Z(n6729) );
  XOR U7920 ( .A(n6730), .B(n6731), .Z(n6726) );
  ANDN U7921 ( .B(n6732), .A(n6733), .Z(n6730) );
  XNOR U7922 ( .A(b[2907]), .B(n6731), .Z(n6732) );
  XNOR U7923 ( .A(b[2907]), .B(n6733), .Z(c[2907]) );
  XNOR U7924 ( .A(a[2907]), .B(n6734), .Z(n6733) );
  IV U7925 ( .A(n6731), .Z(n6734) );
  XOR U7926 ( .A(n6735), .B(n6736), .Z(n6731) );
  ANDN U7927 ( .B(n6737), .A(n6738), .Z(n6735) );
  XNOR U7928 ( .A(b[2906]), .B(n6736), .Z(n6737) );
  XNOR U7929 ( .A(b[2906]), .B(n6738), .Z(c[2906]) );
  XNOR U7930 ( .A(a[2906]), .B(n6739), .Z(n6738) );
  IV U7931 ( .A(n6736), .Z(n6739) );
  XOR U7932 ( .A(n6740), .B(n6741), .Z(n6736) );
  ANDN U7933 ( .B(n6742), .A(n6743), .Z(n6740) );
  XNOR U7934 ( .A(b[2905]), .B(n6741), .Z(n6742) );
  XNOR U7935 ( .A(b[2905]), .B(n6743), .Z(c[2905]) );
  XNOR U7936 ( .A(a[2905]), .B(n6744), .Z(n6743) );
  IV U7937 ( .A(n6741), .Z(n6744) );
  XOR U7938 ( .A(n6745), .B(n6746), .Z(n6741) );
  ANDN U7939 ( .B(n6747), .A(n6748), .Z(n6745) );
  XNOR U7940 ( .A(b[2904]), .B(n6746), .Z(n6747) );
  XNOR U7941 ( .A(b[2904]), .B(n6748), .Z(c[2904]) );
  XNOR U7942 ( .A(a[2904]), .B(n6749), .Z(n6748) );
  IV U7943 ( .A(n6746), .Z(n6749) );
  XOR U7944 ( .A(n6750), .B(n6751), .Z(n6746) );
  ANDN U7945 ( .B(n6752), .A(n6753), .Z(n6750) );
  XNOR U7946 ( .A(b[2903]), .B(n6751), .Z(n6752) );
  XNOR U7947 ( .A(b[2903]), .B(n6753), .Z(c[2903]) );
  XNOR U7948 ( .A(a[2903]), .B(n6754), .Z(n6753) );
  IV U7949 ( .A(n6751), .Z(n6754) );
  XOR U7950 ( .A(n6755), .B(n6756), .Z(n6751) );
  ANDN U7951 ( .B(n6757), .A(n6758), .Z(n6755) );
  XNOR U7952 ( .A(b[2902]), .B(n6756), .Z(n6757) );
  XNOR U7953 ( .A(b[2902]), .B(n6758), .Z(c[2902]) );
  XNOR U7954 ( .A(a[2902]), .B(n6759), .Z(n6758) );
  IV U7955 ( .A(n6756), .Z(n6759) );
  XOR U7956 ( .A(n6760), .B(n6761), .Z(n6756) );
  ANDN U7957 ( .B(n6762), .A(n6763), .Z(n6760) );
  XNOR U7958 ( .A(b[2901]), .B(n6761), .Z(n6762) );
  XNOR U7959 ( .A(b[2901]), .B(n6763), .Z(c[2901]) );
  XNOR U7960 ( .A(a[2901]), .B(n6764), .Z(n6763) );
  IV U7961 ( .A(n6761), .Z(n6764) );
  XOR U7962 ( .A(n6765), .B(n6766), .Z(n6761) );
  ANDN U7963 ( .B(n6767), .A(n6768), .Z(n6765) );
  XNOR U7964 ( .A(b[2900]), .B(n6766), .Z(n6767) );
  XNOR U7965 ( .A(b[2900]), .B(n6768), .Z(c[2900]) );
  XNOR U7966 ( .A(a[2900]), .B(n6769), .Z(n6768) );
  IV U7967 ( .A(n6766), .Z(n6769) );
  XOR U7968 ( .A(n6770), .B(n6771), .Z(n6766) );
  ANDN U7969 ( .B(n6772), .A(n6773), .Z(n6770) );
  XNOR U7970 ( .A(b[2899]), .B(n6771), .Z(n6772) );
  XNOR U7971 ( .A(b[28]), .B(n6774), .Z(c[28]) );
  XNOR U7972 ( .A(b[289]), .B(n6775), .Z(c[289]) );
  XNOR U7973 ( .A(b[2899]), .B(n6773), .Z(c[2899]) );
  XNOR U7974 ( .A(a[2899]), .B(n6776), .Z(n6773) );
  IV U7975 ( .A(n6771), .Z(n6776) );
  XOR U7976 ( .A(n6777), .B(n6778), .Z(n6771) );
  ANDN U7977 ( .B(n6779), .A(n6780), .Z(n6777) );
  XNOR U7978 ( .A(b[2898]), .B(n6778), .Z(n6779) );
  XNOR U7979 ( .A(b[2898]), .B(n6780), .Z(c[2898]) );
  XNOR U7980 ( .A(a[2898]), .B(n6781), .Z(n6780) );
  IV U7981 ( .A(n6778), .Z(n6781) );
  XOR U7982 ( .A(n6782), .B(n6783), .Z(n6778) );
  ANDN U7983 ( .B(n6784), .A(n6785), .Z(n6782) );
  XNOR U7984 ( .A(b[2897]), .B(n6783), .Z(n6784) );
  XNOR U7985 ( .A(b[2897]), .B(n6785), .Z(c[2897]) );
  XNOR U7986 ( .A(a[2897]), .B(n6786), .Z(n6785) );
  IV U7987 ( .A(n6783), .Z(n6786) );
  XOR U7988 ( .A(n6787), .B(n6788), .Z(n6783) );
  ANDN U7989 ( .B(n6789), .A(n6790), .Z(n6787) );
  XNOR U7990 ( .A(b[2896]), .B(n6788), .Z(n6789) );
  XNOR U7991 ( .A(b[2896]), .B(n6790), .Z(c[2896]) );
  XNOR U7992 ( .A(a[2896]), .B(n6791), .Z(n6790) );
  IV U7993 ( .A(n6788), .Z(n6791) );
  XOR U7994 ( .A(n6792), .B(n6793), .Z(n6788) );
  ANDN U7995 ( .B(n6794), .A(n6795), .Z(n6792) );
  XNOR U7996 ( .A(b[2895]), .B(n6793), .Z(n6794) );
  XNOR U7997 ( .A(b[2895]), .B(n6795), .Z(c[2895]) );
  XNOR U7998 ( .A(a[2895]), .B(n6796), .Z(n6795) );
  IV U7999 ( .A(n6793), .Z(n6796) );
  XOR U8000 ( .A(n6797), .B(n6798), .Z(n6793) );
  ANDN U8001 ( .B(n6799), .A(n6800), .Z(n6797) );
  XNOR U8002 ( .A(b[2894]), .B(n6798), .Z(n6799) );
  XNOR U8003 ( .A(b[2894]), .B(n6800), .Z(c[2894]) );
  XNOR U8004 ( .A(a[2894]), .B(n6801), .Z(n6800) );
  IV U8005 ( .A(n6798), .Z(n6801) );
  XOR U8006 ( .A(n6802), .B(n6803), .Z(n6798) );
  ANDN U8007 ( .B(n6804), .A(n6805), .Z(n6802) );
  XNOR U8008 ( .A(b[2893]), .B(n6803), .Z(n6804) );
  XNOR U8009 ( .A(b[2893]), .B(n6805), .Z(c[2893]) );
  XNOR U8010 ( .A(a[2893]), .B(n6806), .Z(n6805) );
  IV U8011 ( .A(n6803), .Z(n6806) );
  XOR U8012 ( .A(n6807), .B(n6808), .Z(n6803) );
  ANDN U8013 ( .B(n6809), .A(n6810), .Z(n6807) );
  XNOR U8014 ( .A(b[2892]), .B(n6808), .Z(n6809) );
  XNOR U8015 ( .A(b[2892]), .B(n6810), .Z(c[2892]) );
  XNOR U8016 ( .A(a[2892]), .B(n6811), .Z(n6810) );
  IV U8017 ( .A(n6808), .Z(n6811) );
  XOR U8018 ( .A(n6812), .B(n6813), .Z(n6808) );
  ANDN U8019 ( .B(n6814), .A(n6815), .Z(n6812) );
  XNOR U8020 ( .A(b[2891]), .B(n6813), .Z(n6814) );
  XNOR U8021 ( .A(b[2891]), .B(n6815), .Z(c[2891]) );
  XNOR U8022 ( .A(a[2891]), .B(n6816), .Z(n6815) );
  IV U8023 ( .A(n6813), .Z(n6816) );
  XOR U8024 ( .A(n6817), .B(n6818), .Z(n6813) );
  ANDN U8025 ( .B(n6819), .A(n6820), .Z(n6817) );
  XNOR U8026 ( .A(b[2890]), .B(n6818), .Z(n6819) );
  XNOR U8027 ( .A(b[2890]), .B(n6820), .Z(c[2890]) );
  XNOR U8028 ( .A(a[2890]), .B(n6821), .Z(n6820) );
  IV U8029 ( .A(n6818), .Z(n6821) );
  XOR U8030 ( .A(n6822), .B(n6823), .Z(n6818) );
  ANDN U8031 ( .B(n6824), .A(n6825), .Z(n6822) );
  XNOR U8032 ( .A(b[2889]), .B(n6823), .Z(n6824) );
  XNOR U8033 ( .A(b[288]), .B(n6826), .Z(c[288]) );
  XNOR U8034 ( .A(b[2889]), .B(n6825), .Z(c[2889]) );
  XNOR U8035 ( .A(a[2889]), .B(n6827), .Z(n6825) );
  IV U8036 ( .A(n6823), .Z(n6827) );
  XOR U8037 ( .A(n6828), .B(n6829), .Z(n6823) );
  ANDN U8038 ( .B(n6830), .A(n6831), .Z(n6828) );
  XNOR U8039 ( .A(b[2888]), .B(n6829), .Z(n6830) );
  XNOR U8040 ( .A(b[2888]), .B(n6831), .Z(c[2888]) );
  XNOR U8041 ( .A(a[2888]), .B(n6832), .Z(n6831) );
  IV U8042 ( .A(n6829), .Z(n6832) );
  XOR U8043 ( .A(n6833), .B(n6834), .Z(n6829) );
  ANDN U8044 ( .B(n6835), .A(n6836), .Z(n6833) );
  XNOR U8045 ( .A(b[2887]), .B(n6834), .Z(n6835) );
  XNOR U8046 ( .A(b[2887]), .B(n6836), .Z(c[2887]) );
  XNOR U8047 ( .A(a[2887]), .B(n6837), .Z(n6836) );
  IV U8048 ( .A(n6834), .Z(n6837) );
  XOR U8049 ( .A(n6838), .B(n6839), .Z(n6834) );
  ANDN U8050 ( .B(n6840), .A(n6841), .Z(n6838) );
  XNOR U8051 ( .A(b[2886]), .B(n6839), .Z(n6840) );
  XNOR U8052 ( .A(b[2886]), .B(n6841), .Z(c[2886]) );
  XNOR U8053 ( .A(a[2886]), .B(n6842), .Z(n6841) );
  IV U8054 ( .A(n6839), .Z(n6842) );
  XOR U8055 ( .A(n6843), .B(n6844), .Z(n6839) );
  ANDN U8056 ( .B(n6845), .A(n6846), .Z(n6843) );
  XNOR U8057 ( .A(b[2885]), .B(n6844), .Z(n6845) );
  XNOR U8058 ( .A(b[2885]), .B(n6846), .Z(c[2885]) );
  XNOR U8059 ( .A(a[2885]), .B(n6847), .Z(n6846) );
  IV U8060 ( .A(n6844), .Z(n6847) );
  XOR U8061 ( .A(n6848), .B(n6849), .Z(n6844) );
  ANDN U8062 ( .B(n6850), .A(n6851), .Z(n6848) );
  XNOR U8063 ( .A(b[2884]), .B(n6849), .Z(n6850) );
  XNOR U8064 ( .A(b[2884]), .B(n6851), .Z(c[2884]) );
  XNOR U8065 ( .A(a[2884]), .B(n6852), .Z(n6851) );
  IV U8066 ( .A(n6849), .Z(n6852) );
  XOR U8067 ( .A(n6853), .B(n6854), .Z(n6849) );
  ANDN U8068 ( .B(n6855), .A(n6856), .Z(n6853) );
  XNOR U8069 ( .A(b[2883]), .B(n6854), .Z(n6855) );
  XNOR U8070 ( .A(b[2883]), .B(n6856), .Z(c[2883]) );
  XNOR U8071 ( .A(a[2883]), .B(n6857), .Z(n6856) );
  IV U8072 ( .A(n6854), .Z(n6857) );
  XOR U8073 ( .A(n6858), .B(n6859), .Z(n6854) );
  ANDN U8074 ( .B(n6860), .A(n6861), .Z(n6858) );
  XNOR U8075 ( .A(b[2882]), .B(n6859), .Z(n6860) );
  XNOR U8076 ( .A(b[2882]), .B(n6861), .Z(c[2882]) );
  XNOR U8077 ( .A(a[2882]), .B(n6862), .Z(n6861) );
  IV U8078 ( .A(n6859), .Z(n6862) );
  XOR U8079 ( .A(n6863), .B(n6864), .Z(n6859) );
  ANDN U8080 ( .B(n6865), .A(n6866), .Z(n6863) );
  XNOR U8081 ( .A(b[2881]), .B(n6864), .Z(n6865) );
  XNOR U8082 ( .A(b[2881]), .B(n6866), .Z(c[2881]) );
  XNOR U8083 ( .A(a[2881]), .B(n6867), .Z(n6866) );
  IV U8084 ( .A(n6864), .Z(n6867) );
  XOR U8085 ( .A(n6868), .B(n6869), .Z(n6864) );
  ANDN U8086 ( .B(n6870), .A(n6871), .Z(n6868) );
  XNOR U8087 ( .A(b[2880]), .B(n6869), .Z(n6870) );
  XNOR U8088 ( .A(b[2880]), .B(n6871), .Z(c[2880]) );
  XNOR U8089 ( .A(a[2880]), .B(n6872), .Z(n6871) );
  IV U8090 ( .A(n6869), .Z(n6872) );
  XOR U8091 ( .A(n6873), .B(n6874), .Z(n6869) );
  ANDN U8092 ( .B(n6875), .A(n6876), .Z(n6873) );
  XNOR U8093 ( .A(b[2879]), .B(n6874), .Z(n6875) );
  XNOR U8094 ( .A(b[287]), .B(n6877), .Z(c[287]) );
  XNOR U8095 ( .A(b[2879]), .B(n6876), .Z(c[2879]) );
  XNOR U8096 ( .A(a[2879]), .B(n6878), .Z(n6876) );
  IV U8097 ( .A(n6874), .Z(n6878) );
  XOR U8098 ( .A(n6879), .B(n6880), .Z(n6874) );
  ANDN U8099 ( .B(n6881), .A(n6882), .Z(n6879) );
  XNOR U8100 ( .A(b[2878]), .B(n6880), .Z(n6881) );
  XNOR U8101 ( .A(b[2878]), .B(n6882), .Z(c[2878]) );
  XNOR U8102 ( .A(a[2878]), .B(n6883), .Z(n6882) );
  IV U8103 ( .A(n6880), .Z(n6883) );
  XOR U8104 ( .A(n6884), .B(n6885), .Z(n6880) );
  ANDN U8105 ( .B(n6886), .A(n6887), .Z(n6884) );
  XNOR U8106 ( .A(b[2877]), .B(n6885), .Z(n6886) );
  XNOR U8107 ( .A(b[2877]), .B(n6887), .Z(c[2877]) );
  XNOR U8108 ( .A(a[2877]), .B(n6888), .Z(n6887) );
  IV U8109 ( .A(n6885), .Z(n6888) );
  XOR U8110 ( .A(n6889), .B(n6890), .Z(n6885) );
  ANDN U8111 ( .B(n6891), .A(n6892), .Z(n6889) );
  XNOR U8112 ( .A(b[2876]), .B(n6890), .Z(n6891) );
  XNOR U8113 ( .A(b[2876]), .B(n6892), .Z(c[2876]) );
  XNOR U8114 ( .A(a[2876]), .B(n6893), .Z(n6892) );
  IV U8115 ( .A(n6890), .Z(n6893) );
  XOR U8116 ( .A(n6894), .B(n6895), .Z(n6890) );
  ANDN U8117 ( .B(n6896), .A(n6897), .Z(n6894) );
  XNOR U8118 ( .A(b[2875]), .B(n6895), .Z(n6896) );
  XNOR U8119 ( .A(b[2875]), .B(n6897), .Z(c[2875]) );
  XNOR U8120 ( .A(a[2875]), .B(n6898), .Z(n6897) );
  IV U8121 ( .A(n6895), .Z(n6898) );
  XOR U8122 ( .A(n6899), .B(n6900), .Z(n6895) );
  ANDN U8123 ( .B(n6901), .A(n6902), .Z(n6899) );
  XNOR U8124 ( .A(b[2874]), .B(n6900), .Z(n6901) );
  XNOR U8125 ( .A(b[2874]), .B(n6902), .Z(c[2874]) );
  XNOR U8126 ( .A(a[2874]), .B(n6903), .Z(n6902) );
  IV U8127 ( .A(n6900), .Z(n6903) );
  XOR U8128 ( .A(n6904), .B(n6905), .Z(n6900) );
  ANDN U8129 ( .B(n6906), .A(n6907), .Z(n6904) );
  XNOR U8130 ( .A(b[2873]), .B(n6905), .Z(n6906) );
  XNOR U8131 ( .A(b[2873]), .B(n6907), .Z(c[2873]) );
  XNOR U8132 ( .A(a[2873]), .B(n6908), .Z(n6907) );
  IV U8133 ( .A(n6905), .Z(n6908) );
  XOR U8134 ( .A(n6909), .B(n6910), .Z(n6905) );
  ANDN U8135 ( .B(n6911), .A(n6912), .Z(n6909) );
  XNOR U8136 ( .A(b[2872]), .B(n6910), .Z(n6911) );
  XNOR U8137 ( .A(b[2872]), .B(n6912), .Z(c[2872]) );
  XNOR U8138 ( .A(a[2872]), .B(n6913), .Z(n6912) );
  IV U8139 ( .A(n6910), .Z(n6913) );
  XOR U8140 ( .A(n6914), .B(n6915), .Z(n6910) );
  ANDN U8141 ( .B(n6916), .A(n6917), .Z(n6914) );
  XNOR U8142 ( .A(b[2871]), .B(n6915), .Z(n6916) );
  XNOR U8143 ( .A(b[2871]), .B(n6917), .Z(c[2871]) );
  XNOR U8144 ( .A(a[2871]), .B(n6918), .Z(n6917) );
  IV U8145 ( .A(n6915), .Z(n6918) );
  XOR U8146 ( .A(n6919), .B(n6920), .Z(n6915) );
  ANDN U8147 ( .B(n6921), .A(n6922), .Z(n6919) );
  XNOR U8148 ( .A(b[2870]), .B(n6920), .Z(n6921) );
  XNOR U8149 ( .A(b[2870]), .B(n6922), .Z(c[2870]) );
  XNOR U8150 ( .A(a[2870]), .B(n6923), .Z(n6922) );
  IV U8151 ( .A(n6920), .Z(n6923) );
  XOR U8152 ( .A(n6924), .B(n6925), .Z(n6920) );
  ANDN U8153 ( .B(n6926), .A(n6927), .Z(n6924) );
  XNOR U8154 ( .A(b[2869]), .B(n6925), .Z(n6926) );
  XNOR U8155 ( .A(b[286]), .B(n6928), .Z(c[286]) );
  XNOR U8156 ( .A(b[2869]), .B(n6927), .Z(c[2869]) );
  XNOR U8157 ( .A(a[2869]), .B(n6929), .Z(n6927) );
  IV U8158 ( .A(n6925), .Z(n6929) );
  XOR U8159 ( .A(n6930), .B(n6931), .Z(n6925) );
  ANDN U8160 ( .B(n6932), .A(n6933), .Z(n6930) );
  XNOR U8161 ( .A(b[2868]), .B(n6931), .Z(n6932) );
  XNOR U8162 ( .A(b[2868]), .B(n6933), .Z(c[2868]) );
  XNOR U8163 ( .A(a[2868]), .B(n6934), .Z(n6933) );
  IV U8164 ( .A(n6931), .Z(n6934) );
  XOR U8165 ( .A(n6935), .B(n6936), .Z(n6931) );
  ANDN U8166 ( .B(n6937), .A(n6938), .Z(n6935) );
  XNOR U8167 ( .A(b[2867]), .B(n6936), .Z(n6937) );
  XNOR U8168 ( .A(b[2867]), .B(n6938), .Z(c[2867]) );
  XNOR U8169 ( .A(a[2867]), .B(n6939), .Z(n6938) );
  IV U8170 ( .A(n6936), .Z(n6939) );
  XOR U8171 ( .A(n6940), .B(n6941), .Z(n6936) );
  ANDN U8172 ( .B(n6942), .A(n6943), .Z(n6940) );
  XNOR U8173 ( .A(b[2866]), .B(n6941), .Z(n6942) );
  XNOR U8174 ( .A(b[2866]), .B(n6943), .Z(c[2866]) );
  XNOR U8175 ( .A(a[2866]), .B(n6944), .Z(n6943) );
  IV U8176 ( .A(n6941), .Z(n6944) );
  XOR U8177 ( .A(n6945), .B(n6946), .Z(n6941) );
  ANDN U8178 ( .B(n6947), .A(n6948), .Z(n6945) );
  XNOR U8179 ( .A(b[2865]), .B(n6946), .Z(n6947) );
  XNOR U8180 ( .A(b[2865]), .B(n6948), .Z(c[2865]) );
  XNOR U8181 ( .A(a[2865]), .B(n6949), .Z(n6948) );
  IV U8182 ( .A(n6946), .Z(n6949) );
  XOR U8183 ( .A(n6950), .B(n6951), .Z(n6946) );
  ANDN U8184 ( .B(n6952), .A(n6953), .Z(n6950) );
  XNOR U8185 ( .A(b[2864]), .B(n6951), .Z(n6952) );
  XNOR U8186 ( .A(b[2864]), .B(n6953), .Z(c[2864]) );
  XNOR U8187 ( .A(a[2864]), .B(n6954), .Z(n6953) );
  IV U8188 ( .A(n6951), .Z(n6954) );
  XOR U8189 ( .A(n6955), .B(n6956), .Z(n6951) );
  ANDN U8190 ( .B(n6957), .A(n6958), .Z(n6955) );
  XNOR U8191 ( .A(b[2863]), .B(n6956), .Z(n6957) );
  XNOR U8192 ( .A(b[2863]), .B(n6958), .Z(c[2863]) );
  XNOR U8193 ( .A(a[2863]), .B(n6959), .Z(n6958) );
  IV U8194 ( .A(n6956), .Z(n6959) );
  XOR U8195 ( .A(n6960), .B(n6961), .Z(n6956) );
  ANDN U8196 ( .B(n6962), .A(n6963), .Z(n6960) );
  XNOR U8197 ( .A(b[2862]), .B(n6961), .Z(n6962) );
  XNOR U8198 ( .A(b[2862]), .B(n6963), .Z(c[2862]) );
  XNOR U8199 ( .A(a[2862]), .B(n6964), .Z(n6963) );
  IV U8200 ( .A(n6961), .Z(n6964) );
  XOR U8201 ( .A(n6965), .B(n6966), .Z(n6961) );
  ANDN U8202 ( .B(n6967), .A(n6968), .Z(n6965) );
  XNOR U8203 ( .A(b[2861]), .B(n6966), .Z(n6967) );
  XNOR U8204 ( .A(b[2861]), .B(n6968), .Z(c[2861]) );
  XNOR U8205 ( .A(a[2861]), .B(n6969), .Z(n6968) );
  IV U8206 ( .A(n6966), .Z(n6969) );
  XOR U8207 ( .A(n6970), .B(n6971), .Z(n6966) );
  ANDN U8208 ( .B(n6972), .A(n6973), .Z(n6970) );
  XNOR U8209 ( .A(b[2860]), .B(n6971), .Z(n6972) );
  XNOR U8210 ( .A(b[2860]), .B(n6973), .Z(c[2860]) );
  XNOR U8211 ( .A(a[2860]), .B(n6974), .Z(n6973) );
  IV U8212 ( .A(n6971), .Z(n6974) );
  XOR U8213 ( .A(n6975), .B(n6976), .Z(n6971) );
  ANDN U8214 ( .B(n6977), .A(n6978), .Z(n6975) );
  XNOR U8215 ( .A(b[2859]), .B(n6976), .Z(n6977) );
  XNOR U8216 ( .A(b[285]), .B(n6979), .Z(c[285]) );
  XNOR U8217 ( .A(b[2859]), .B(n6978), .Z(c[2859]) );
  XNOR U8218 ( .A(a[2859]), .B(n6980), .Z(n6978) );
  IV U8219 ( .A(n6976), .Z(n6980) );
  XOR U8220 ( .A(n6981), .B(n6982), .Z(n6976) );
  ANDN U8221 ( .B(n6983), .A(n6984), .Z(n6981) );
  XNOR U8222 ( .A(b[2858]), .B(n6982), .Z(n6983) );
  XNOR U8223 ( .A(b[2858]), .B(n6984), .Z(c[2858]) );
  XNOR U8224 ( .A(a[2858]), .B(n6985), .Z(n6984) );
  IV U8225 ( .A(n6982), .Z(n6985) );
  XOR U8226 ( .A(n6986), .B(n6987), .Z(n6982) );
  ANDN U8227 ( .B(n6988), .A(n6989), .Z(n6986) );
  XNOR U8228 ( .A(b[2857]), .B(n6987), .Z(n6988) );
  XNOR U8229 ( .A(b[2857]), .B(n6989), .Z(c[2857]) );
  XNOR U8230 ( .A(a[2857]), .B(n6990), .Z(n6989) );
  IV U8231 ( .A(n6987), .Z(n6990) );
  XOR U8232 ( .A(n6991), .B(n6992), .Z(n6987) );
  ANDN U8233 ( .B(n6993), .A(n6994), .Z(n6991) );
  XNOR U8234 ( .A(b[2856]), .B(n6992), .Z(n6993) );
  XNOR U8235 ( .A(b[2856]), .B(n6994), .Z(c[2856]) );
  XNOR U8236 ( .A(a[2856]), .B(n6995), .Z(n6994) );
  IV U8237 ( .A(n6992), .Z(n6995) );
  XOR U8238 ( .A(n6996), .B(n6997), .Z(n6992) );
  ANDN U8239 ( .B(n6998), .A(n6999), .Z(n6996) );
  XNOR U8240 ( .A(b[2855]), .B(n6997), .Z(n6998) );
  XNOR U8241 ( .A(b[2855]), .B(n6999), .Z(c[2855]) );
  XNOR U8242 ( .A(a[2855]), .B(n7000), .Z(n6999) );
  IV U8243 ( .A(n6997), .Z(n7000) );
  XOR U8244 ( .A(n7001), .B(n7002), .Z(n6997) );
  ANDN U8245 ( .B(n7003), .A(n7004), .Z(n7001) );
  XNOR U8246 ( .A(b[2854]), .B(n7002), .Z(n7003) );
  XNOR U8247 ( .A(b[2854]), .B(n7004), .Z(c[2854]) );
  XNOR U8248 ( .A(a[2854]), .B(n7005), .Z(n7004) );
  IV U8249 ( .A(n7002), .Z(n7005) );
  XOR U8250 ( .A(n7006), .B(n7007), .Z(n7002) );
  ANDN U8251 ( .B(n7008), .A(n7009), .Z(n7006) );
  XNOR U8252 ( .A(b[2853]), .B(n7007), .Z(n7008) );
  XNOR U8253 ( .A(b[2853]), .B(n7009), .Z(c[2853]) );
  XNOR U8254 ( .A(a[2853]), .B(n7010), .Z(n7009) );
  IV U8255 ( .A(n7007), .Z(n7010) );
  XOR U8256 ( .A(n7011), .B(n7012), .Z(n7007) );
  ANDN U8257 ( .B(n7013), .A(n7014), .Z(n7011) );
  XNOR U8258 ( .A(b[2852]), .B(n7012), .Z(n7013) );
  XNOR U8259 ( .A(b[2852]), .B(n7014), .Z(c[2852]) );
  XNOR U8260 ( .A(a[2852]), .B(n7015), .Z(n7014) );
  IV U8261 ( .A(n7012), .Z(n7015) );
  XOR U8262 ( .A(n7016), .B(n7017), .Z(n7012) );
  ANDN U8263 ( .B(n7018), .A(n7019), .Z(n7016) );
  XNOR U8264 ( .A(b[2851]), .B(n7017), .Z(n7018) );
  XNOR U8265 ( .A(b[2851]), .B(n7019), .Z(c[2851]) );
  XNOR U8266 ( .A(a[2851]), .B(n7020), .Z(n7019) );
  IV U8267 ( .A(n7017), .Z(n7020) );
  XOR U8268 ( .A(n7021), .B(n7022), .Z(n7017) );
  ANDN U8269 ( .B(n7023), .A(n7024), .Z(n7021) );
  XNOR U8270 ( .A(b[2850]), .B(n7022), .Z(n7023) );
  XNOR U8271 ( .A(b[2850]), .B(n7024), .Z(c[2850]) );
  XNOR U8272 ( .A(a[2850]), .B(n7025), .Z(n7024) );
  IV U8273 ( .A(n7022), .Z(n7025) );
  XOR U8274 ( .A(n7026), .B(n7027), .Z(n7022) );
  ANDN U8275 ( .B(n7028), .A(n7029), .Z(n7026) );
  XNOR U8276 ( .A(b[2849]), .B(n7027), .Z(n7028) );
  XNOR U8277 ( .A(b[284]), .B(n7030), .Z(c[284]) );
  XNOR U8278 ( .A(b[2849]), .B(n7029), .Z(c[2849]) );
  XNOR U8279 ( .A(a[2849]), .B(n7031), .Z(n7029) );
  IV U8280 ( .A(n7027), .Z(n7031) );
  XOR U8281 ( .A(n7032), .B(n7033), .Z(n7027) );
  ANDN U8282 ( .B(n7034), .A(n7035), .Z(n7032) );
  XNOR U8283 ( .A(b[2848]), .B(n7033), .Z(n7034) );
  XNOR U8284 ( .A(b[2848]), .B(n7035), .Z(c[2848]) );
  XNOR U8285 ( .A(a[2848]), .B(n7036), .Z(n7035) );
  IV U8286 ( .A(n7033), .Z(n7036) );
  XOR U8287 ( .A(n7037), .B(n7038), .Z(n7033) );
  ANDN U8288 ( .B(n7039), .A(n7040), .Z(n7037) );
  XNOR U8289 ( .A(b[2847]), .B(n7038), .Z(n7039) );
  XNOR U8290 ( .A(b[2847]), .B(n7040), .Z(c[2847]) );
  XNOR U8291 ( .A(a[2847]), .B(n7041), .Z(n7040) );
  IV U8292 ( .A(n7038), .Z(n7041) );
  XOR U8293 ( .A(n7042), .B(n7043), .Z(n7038) );
  ANDN U8294 ( .B(n7044), .A(n7045), .Z(n7042) );
  XNOR U8295 ( .A(b[2846]), .B(n7043), .Z(n7044) );
  XNOR U8296 ( .A(b[2846]), .B(n7045), .Z(c[2846]) );
  XNOR U8297 ( .A(a[2846]), .B(n7046), .Z(n7045) );
  IV U8298 ( .A(n7043), .Z(n7046) );
  XOR U8299 ( .A(n7047), .B(n7048), .Z(n7043) );
  ANDN U8300 ( .B(n7049), .A(n7050), .Z(n7047) );
  XNOR U8301 ( .A(b[2845]), .B(n7048), .Z(n7049) );
  XNOR U8302 ( .A(b[2845]), .B(n7050), .Z(c[2845]) );
  XNOR U8303 ( .A(a[2845]), .B(n7051), .Z(n7050) );
  IV U8304 ( .A(n7048), .Z(n7051) );
  XOR U8305 ( .A(n7052), .B(n7053), .Z(n7048) );
  ANDN U8306 ( .B(n7054), .A(n7055), .Z(n7052) );
  XNOR U8307 ( .A(b[2844]), .B(n7053), .Z(n7054) );
  XNOR U8308 ( .A(b[2844]), .B(n7055), .Z(c[2844]) );
  XNOR U8309 ( .A(a[2844]), .B(n7056), .Z(n7055) );
  IV U8310 ( .A(n7053), .Z(n7056) );
  XOR U8311 ( .A(n7057), .B(n7058), .Z(n7053) );
  ANDN U8312 ( .B(n7059), .A(n7060), .Z(n7057) );
  XNOR U8313 ( .A(b[2843]), .B(n7058), .Z(n7059) );
  XNOR U8314 ( .A(b[2843]), .B(n7060), .Z(c[2843]) );
  XNOR U8315 ( .A(a[2843]), .B(n7061), .Z(n7060) );
  IV U8316 ( .A(n7058), .Z(n7061) );
  XOR U8317 ( .A(n7062), .B(n7063), .Z(n7058) );
  ANDN U8318 ( .B(n7064), .A(n7065), .Z(n7062) );
  XNOR U8319 ( .A(b[2842]), .B(n7063), .Z(n7064) );
  XNOR U8320 ( .A(b[2842]), .B(n7065), .Z(c[2842]) );
  XNOR U8321 ( .A(a[2842]), .B(n7066), .Z(n7065) );
  IV U8322 ( .A(n7063), .Z(n7066) );
  XOR U8323 ( .A(n7067), .B(n7068), .Z(n7063) );
  ANDN U8324 ( .B(n7069), .A(n7070), .Z(n7067) );
  XNOR U8325 ( .A(b[2841]), .B(n7068), .Z(n7069) );
  XNOR U8326 ( .A(b[2841]), .B(n7070), .Z(c[2841]) );
  XNOR U8327 ( .A(a[2841]), .B(n7071), .Z(n7070) );
  IV U8328 ( .A(n7068), .Z(n7071) );
  XOR U8329 ( .A(n7072), .B(n7073), .Z(n7068) );
  ANDN U8330 ( .B(n7074), .A(n7075), .Z(n7072) );
  XNOR U8331 ( .A(b[2840]), .B(n7073), .Z(n7074) );
  XNOR U8332 ( .A(b[2840]), .B(n7075), .Z(c[2840]) );
  XNOR U8333 ( .A(a[2840]), .B(n7076), .Z(n7075) );
  IV U8334 ( .A(n7073), .Z(n7076) );
  XOR U8335 ( .A(n7077), .B(n7078), .Z(n7073) );
  ANDN U8336 ( .B(n7079), .A(n7080), .Z(n7077) );
  XNOR U8337 ( .A(b[2839]), .B(n7078), .Z(n7079) );
  XNOR U8338 ( .A(b[283]), .B(n7081), .Z(c[283]) );
  XNOR U8339 ( .A(b[2839]), .B(n7080), .Z(c[2839]) );
  XNOR U8340 ( .A(a[2839]), .B(n7082), .Z(n7080) );
  IV U8341 ( .A(n7078), .Z(n7082) );
  XOR U8342 ( .A(n7083), .B(n7084), .Z(n7078) );
  ANDN U8343 ( .B(n7085), .A(n7086), .Z(n7083) );
  XNOR U8344 ( .A(b[2838]), .B(n7084), .Z(n7085) );
  XNOR U8345 ( .A(b[2838]), .B(n7086), .Z(c[2838]) );
  XNOR U8346 ( .A(a[2838]), .B(n7087), .Z(n7086) );
  IV U8347 ( .A(n7084), .Z(n7087) );
  XOR U8348 ( .A(n7088), .B(n7089), .Z(n7084) );
  ANDN U8349 ( .B(n7090), .A(n7091), .Z(n7088) );
  XNOR U8350 ( .A(b[2837]), .B(n7089), .Z(n7090) );
  XNOR U8351 ( .A(b[2837]), .B(n7091), .Z(c[2837]) );
  XNOR U8352 ( .A(a[2837]), .B(n7092), .Z(n7091) );
  IV U8353 ( .A(n7089), .Z(n7092) );
  XOR U8354 ( .A(n7093), .B(n7094), .Z(n7089) );
  ANDN U8355 ( .B(n7095), .A(n7096), .Z(n7093) );
  XNOR U8356 ( .A(b[2836]), .B(n7094), .Z(n7095) );
  XNOR U8357 ( .A(b[2836]), .B(n7096), .Z(c[2836]) );
  XNOR U8358 ( .A(a[2836]), .B(n7097), .Z(n7096) );
  IV U8359 ( .A(n7094), .Z(n7097) );
  XOR U8360 ( .A(n7098), .B(n7099), .Z(n7094) );
  ANDN U8361 ( .B(n7100), .A(n7101), .Z(n7098) );
  XNOR U8362 ( .A(b[2835]), .B(n7099), .Z(n7100) );
  XNOR U8363 ( .A(b[2835]), .B(n7101), .Z(c[2835]) );
  XNOR U8364 ( .A(a[2835]), .B(n7102), .Z(n7101) );
  IV U8365 ( .A(n7099), .Z(n7102) );
  XOR U8366 ( .A(n7103), .B(n7104), .Z(n7099) );
  ANDN U8367 ( .B(n7105), .A(n7106), .Z(n7103) );
  XNOR U8368 ( .A(b[2834]), .B(n7104), .Z(n7105) );
  XNOR U8369 ( .A(b[2834]), .B(n7106), .Z(c[2834]) );
  XNOR U8370 ( .A(a[2834]), .B(n7107), .Z(n7106) );
  IV U8371 ( .A(n7104), .Z(n7107) );
  XOR U8372 ( .A(n7108), .B(n7109), .Z(n7104) );
  ANDN U8373 ( .B(n7110), .A(n7111), .Z(n7108) );
  XNOR U8374 ( .A(b[2833]), .B(n7109), .Z(n7110) );
  XNOR U8375 ( .A(b[2833]), .B(n7111), .Z(c[2833]) );
  XNOR U8376 ( .A(a[2833]), .B(n7112), .Z(n7111) );
  IV U8377 ( .A(n7109), .Z(n7112) );
  XOR U8378 ( .A(n7113), .B(n7114), .Z(n7109) );
  ANDN U8379 ( .B(n7115), .A(n7116), .Z(n7113) );
  XNOR U8380 ( .A(b[2832]), .B(n7114), .Z(n7115) );
  XNOR U8381 ( .A(b[2832]), .B(n7116), .Z(c[2832]) );
  XNOR U8382 ( .A(a[2832]), .B(n7117), .Z(n7116) );
  IV U8383 ( .A(n7114), .Z(n7117) );
  XOR U8384 ( .A(n7118), .B(n7119), .Z(n7114) );
  ANDN U8385 ( .B(n7120), .A(n7121), .Z(n7118) );
  XNOR U8386 ( .A(b[2831]), .B(n7119), .Z(n7120) );
  XNOR U8387 ( .A(b[2831]), .B(n7121), .Z(c[2831]) );
  XNOR U8388 ( .A(a[2831]), .B(n7122), .Z(n7121) );
  IV U8389 ( .A(n7119), .Z(n7122) );
  XOR U8390 ( .A(n7123), .B(n7124), .Z(n7119) );
  ANDN U8391 ( .B(n7125), .A(n7126), .Z(n7123) );
  XNOR U8392 ( .A(b[2830]), .B(n7124), .Z(n7125) );
  XNOR U8393 ( .A(b[2830]), .B(n7126), .Z(c[2830]) );
  XNOR U8394 ( .A(a[2830]), .B(n7127), .Z(n7126) );
  IV U8395 ( .A(n7124), .Z(n7127) );
  XOR U8396 ( .A(n7128), .B(n7129), .Z(n7124) );
  ANDN U8397 ( .B(n7130), .A(n7131), .Z(n7128) );
  XNOR U8398 ( .A(b[2829]), .B(n7129), .Z(n7130) );
  XNOR U8399 ( .A(b[282]), .B(n7132), .Z(c[282]) );
  XNOR U8400 ( .A(b[2829]), .B(n7131), .Z(c[2829]) );
  XNOR U8401 ( .A(a[2829]), .B(n7133), .Z(n7131) );
  IV U8402 ( .A(n7129), .Z(n7133) );
  XOR U8403 ( .A(n7134), .B(n7135), .Z(n7129) );
  ANDN U8404 ( .B(n7136), .A(n7137), .Z(n7134) );
  XNOR U8405 ( .A(b[2828]), .B(n7135), .Z(n7136) );
  XNOR U8406 ( .A(b[2828]), .B(n7137), .Z(c[2828]) );
  XNOR U8407 ( .A(a[2828]), .B(n7138), .Z(n7137) );
  IV U8408 ( .A(n7135), .Z(n7138) );
  XOR U8409 ( .A(n7139), .B(n7140), .Z(n7135) );
  ANDN U8410 ( .B(n7141), .A(n7142), .Z(n7139) );
  XNOR U8411 ( .A(b[2827]), .B(n7140), .Z(n7141) );
  XNOR U8412 ( .A(b[2827]), .B(n7142), .Z(c[2827]) );
  XNOR U8413 ( .A(a[2827]), .B(n7143), .Z(n7142) );
  IV U8414 ( .A(n7140), .Z(n7143) );
  XOR U8415 ( .A(n7144), .B(n7145), .Z(n7140) );
  ANDN U8416 ( .B(n7146), .A(n7147), .Z(n7144) );
  XNOR U8417 ( .A(b[2826]), .B(n7145), .Z(n7146) );
  XNOR U8418 ( .A(b[2826]), .B(n7147), .Z(c[2826]) );
  XNOR U8419 ( .A(a[2826]), .B(n7148), .Z(n7147) );
  IV U8420 ( .A(n7145), .Z(n7148) );
  XOR U8421 ( .A(n7149), .B(n7150), .Z(n7145) );
  ANDN U8422 ( .B(n7151), .A(n7152), .Z(n7149) );
  XNOR U8423 ( .A(b[2825]), .B(n7150), .Z(n7151) );
  XNOR U8424 ( .A(b[2825]), .B(n7152), .Z(c[2825]) );
  XNOR U8425 ( .A(a[2825]), .B(n7153), .Z(n7152) );
  IV U8426 ( .A(n7150), .Z(n7153) );
  XOR U8427 ( .A(n7154), .B(n7155), .Z(n7150) );
  ANDN U8428 ( .B(n7156), .A(n7157), .Z(n7154) );
  XNOR U8429 ( .A(b[2824]), .B(n7155), .Z(n7156) );
  XNOR U8430 ( .A(b[2824]), .B(n7157), .Z(c[2824]) );
  XNOR U8431 ( .A(a[2824]), .B(n7158), .Z(n7157) );
  IV U8432 ( .A(n7155), .Z(n7158) );
  XOR U8433 ( .A(n7159), .B(n7160), .Z(n7155) );
  ANDN U8434 ( .B(n7161), .A(n7162), .Z(n7159) );
  XNOR U8435 ( .A(b[2823]), .B(n7160), .Z(n7161) );
  XNOR U8436 ( .A(b[2823]), .B(n7162), .Z(c[2823]) );
  XNOR U8437 ( .A(a[2823]), .B(n7163), .Z(n7162) );
  IV U8438 ( .A(n7160), .Z(n7163) );
  XOR U8439 ( .A(n7164), .B(n7165), .Z(n7160) );
  ANDN U8440 ( .B(n7166), .A(n7167), .Z(n7164) );
  XNOR U8441 ( .A(b[2822]), .B(n7165), .Z(n7166) );
  XNOR U8442 ( .A(b[2822]), .B(n7167), .Z(c[2822]) );
  XNOR U8443 ( .A(a[2822]), .B(n7168), .Z(n7167) );
  IV U8444 ( .A(n7165), .Z(n7168) );
  XOR U8445 ( .A(n7169), .B(n7170), .Z(n7165) );
  ANDN U8446 ( .B(n7171), .A(n7172), .Z(n7169) );
  XNOR U8447 ( .A(b[2821]), .B(n7170), .Z(n7171) );
  XNOR U8448 ( .A(b[2821]), .B(n7172), .Z(c[2821]) );
  XNOR U8449 ( .A(a[2821]), .B(n7173), .Z(n7172) );
  IV U8450 ( .A(n7170), .Z(n7173) );
  XOR U8451 ( .A(n7174), .B(n7175), .Z(n7170) );
  ANDN U8452 ( .B(n7176), .A(n7177), .Z(n7174) );
  XNOR U8453 ( .A(b[2820]), .B(n7175), .Z(n7176) );
  XNOR U8454 ( .A(b[2820]), .B(n7177), .Z(c[2820]) );
  XNOR U8455 ( .A(a[2820]), .B(n7178), .Z(n7177) );
  IV U8456 ( .A(n7175), .Z(n7178) );
  XOR U8457 ( .A(n7179), .B(n7180), .Z(n7175) );
  ANDN U8458 ( .B(n7181), .A(n7182), .Z(n7179) );
  XNOR U8459 ( .A(b[2819]), .B(n7180), .Z(n7181) );
  XNOR U8460 ( .A(b[281]), .B(n7183), .Z(c[281]) );
  XNOR U8461 ( .A(b[2819]), .B(n7182), .Z(c[2819]) );
  XNOR U8462 ( .A(a[2819]), .B(n7184), .Z(n7182) );
  IV U8463 ( .A(n7180), .Z(n7184) );
  XOR U8464 ( .A(n7185), .B(n7186), .Z(n7180) );
  ANDN U8465 ( .B(n7187), .A(n7188), .Z(n7185) );
  XNOR U8466 ( .A(b[2818]), .B(n7186), .Z(n7187) );
  XNOR U8467 ( .A(b[2818]), .B(n7188), .Z(c[2818]) );
  XNOR U8468 ( .A(a[2818]), .B(n7189), .Z(n7188) );
  IV U8469 ( .A(n7186), .Z(n7189) );
  XOR U8470 ( .A(n7190), .B(n7191), .Z(n7186) );
  ANDN U8471 ( .B(n7192), .A(n7193), .Z(n7190) );
  XNOR U8472 ( .A(b[2817]), .B(n7191), .Z(n7192) );
  XNOR U8473 ( .A(b[2817]), .B(n7193), .Z(c[2817]) );
  XNOR U8474 ( .A(a[2817]), .B(n7194), .Z(n7193) );
  IV U8475 ( .A(n7191), .Z(n7194) );
  XOR U8476 ( .A(n7195), .B(n7196), .Z(n7191) );
  ANDN U8477 ( .B(n7197), .A(n7198), .Z(n7195) );
  XNOR U8478 ( .A(b[2816]), .B(n7196), .Z(n7197) );
  XNOR U8479 ( .A(b[2816]), .B(n7198), .Z(c[2816]) );
  XNOR U8480 ( .A(a[2816]), .B(n7199), .Z(n7198) );
  IV U8481 ( .A(n7196), .Z(n7199) );
  XOR U8482 ( .A(n7200), .B(n7201), .Z(n7196) );
  ANDN U8483 ( .B(n7202), .A(n7203), .Z(n7200) );
  XNOR U8484 ( .A(b[2815]), .B(n7201), .Z(n7202) );
  XNOR U8485 ( .A(b[2815]), .B(n7203), .Z(c[2815]) );
  XNOR U8486 ( .A(a[2815]), .B(n7204), .Z(n7203) );
  IV U8487 ( .A(n7201), .Z(n7204) );
  XOR U8488 ( .A(n7205), .B(n7206), .Z(n7201) );
  ANDN U8489 ( .B(n7207), .A(n7208), .Z(n7205) );
  XNOR U8490 ( .A(b[2814]), .B(n7206), .Z(n7207) );
  XNOR U8491 ( .A(b[2814]), .B(n7208), .Z(c[2814]) );
  XNOR U8492 ( .A(a[2814]), .B(n7209), .Z(n7208) );
  IV U8493 ( .A(n7206), .Z(n7209) );
  XOR U8494 ( .A(n7210), .B(n7211), .Z(n7206) );
  ANDN U8495 ( .B(n7212), .A(n7213), .Z(n7210) );
  XNOR U8496 ( .A(b[2813]), .B(n7211), .Z(n7212) );
  XNOR U8497 ( .A(b[2813]), .B(n7213), .Z(c[2813]) );
  XNOR U8498 ( .A(a[2813]), .B(n7214), .Z(n7213) );
  IV U8499 ( .A(n7211), .Z(n7214) );
  XOR U8500 ( .A(n7215), .B(n7216), .Z(n7211) );
  ANDN U8501 ( .B(n7217), .A(n7218), .Z(n7215) );
  XNOR U8502 ( .A(b[2812]), .B(n7216), .Z(n7217) );
  XNOR U8503 ( .A(b[2812]), .B(n7218), .Z(c[2812]) );
  XNOR U8504 ( .A(a[2812]), .B(n7219), .Z(n7218) );
  IV U8505 ( .A(n7216), .Z(n7219) );
  XOR U8506 ( .A(n7220), .B(n7221), .Z(n7216) );
  ANDN U8507 ( .B(n7222), .A(n7223), .Z(n7220) );
  XNOR U8508 ( .A(b[2811]), .B(n7221), .Z(n7222) );
  XNOR U8509 ( .A(b[2811]), .B(n7223), .Z(c[2811]) );
  XNOR U8510 ( .A(a[2811]), .B(n7224), .Z(n7223) );
  IV U8511 ( .A(n7221), .Z(n7224) );
  XOR U8512 ( .A(n7225), .B(n7226), .Z(n7221) );
  ANDN U8513 ( .B(n7227), .A(n7228), .Z(n7225) );
  XNOR U8514 ( .A(b[2810]), .B(n7226), .Z(n7227) );
  XNOR U8515 ( .A(b[2810]), .B(n7228), .Z(c[2810]) );
  XNOR U8516 ( .A(a[2810]), .B(n7229), .Z(n7228) );
  IV U8517 ( .A(n7226), .Z(n7229) );
  XOR U8518 ( .A(n7230), .B(n7231), .Z(n7226) );
  ANDN U8519 ( .B(n7232), .A(n7233), .Z(n7230) );
  XNOR U8520 ( .A(b[2809]), .B(n7231), .Z(n7232) );
  XNOR U8521 ( .A(b[280]), .B(n7234), .Z(c[280]) );
  XNOR U8522 ( .A(b[2809]), .B(n7233), .Z(c[2809]) );
  XNOR U8523 ( .A(a[2809]), .B(n7235), .Z(n7233) );
  IV U8524 ( .A(n7231), .Z(n7235) );
  XOR U8525 ( .A(n7236), .B(n7237), .Z(n7231) );
  ANDN U8526 ( .B(n7238), .A(n7239), .Z(n7236) );
  XNOR U8527 ( .A(b[2808]), .B(n7237), .Z(n7238) );
  XNOR U8528 ( .A(b[2808]), .B(n7239), .Z(c[2808]) );
  XNOR U8529 ( .A(a[2808]), .B(n7240), .Z(n7239) );
  IV U8530 ( .A(n7237), .Z(n7240) );
  XOR U8531 ( .A(n7241), .B(n7242), .Z(n7237) );
  ANDN U8532 ( .B(n7243), .A(n7244), .Z(n7241) );
  XNOR U8533 ( .A(b[2807]), .B(n7242), .Z(n7243) );
  XNOR U8534 ( .A(b[2807]), .B(n7244), .Z(c[2807]) );
  XNOR U8535 ( .A(a[2807]), .B(n7245), .Z(n7244) );
  IV U8536 ( .A(n7242), .Z(n7245) );
  XOR U8537 ( .A(n7246), .B(n7247), .Z(n7242) );
  ANDN U8538 ( .B(n7248), .A(n7249), .Z(n7246) );
  XNOR U8539 ( .A(b[2806]), .B(n7247), .Z(n7248) );
  XNOR U8540 ( .A(b[2806]), .B(n7249), .Z(c[2806]) );
  XNOR U8541 ( .A(a[2806]), .B(n7250), .Z(n7249) );
  IV U8542 ( .A(n7247), .Z(n7250) );
  XOR U8543 ( .A(n7251), .B(n7252), .Z(n7247) );
  ANDN U8544 ( .B(n7253), .A(n7254), .Z(n7251) );
  XNOR U8545 ( .A(b[2805]), .B(n7252), .Z(n7253) );
  XNOR U8546 ( .A(b[2805]), .B(n7254), .Z(c[2805]) );
  XNOR U8547 ( .A(a[2805]), .B(n7255), .Z(n7254) );
  IV U8548 ( .A(n7252), .Z(n7255) );
  XOR U8549 ( .A(n7256), .B(n7257), .Z(n7252) );
  ANDN U8550 ( .B(n7258), .A(n7259), .Z(n7256) );
  XNOR U8551 ( .A(b[2804]), .B(n7257), .Z(n7258) );
  XNOR U8552 ( .A(b[2804]), .B(n7259), .Z(c[2804]) );
  XNOR U8553 ( .A(a[2804]), .B(n7260), .Z(n7259) );
  IV U8554 ( .A(n7257), .Z(n7260) );
  XOR U8555 ( .A(n7261), .B(n7262), .Z(n7257) );
  ANDN U8556 ( .B(n7263), .A(n7264), .Z(n7261) );
  XNOR U8557 ( .A(b[2803]), .B(n7262), .Z(n7263) );
  XNOR U8558 ( .A(b[2803]), .B(n7264), .Z(c[2803]) );
  XNOR U8559 ( .A(a[2803]), .B(n7265), .Z(n7264) );
  IV U8560 ( .A(n7262), .Z(n7265) );
  XOR U8561 ( .A(n7266), .B(n7267), .Z(n7262) );
  ANDN U8562 ( .B(n7268), .A(n7269), .Z(n7266) );
  XNOR U8563 ( .A(b[2802]), .B(n7267), .Z(n7268) );
  XNOR U8564 ( .A(b[2802]), .B(n7269), .Z(c[2802]) );
  XNOR U8565 ( .A(a[2802]), .B(n7270), .Z(n7269) );
  IV U8566 ( .A(n7267), .Z(n7270) );
  XOR U8567 ( .A(n7271), .B(n7272), .Z(n7267) );
  ANDN U8568 ( .B(n7273), .A(n7274), .Z(n7271) );
  XNOR U8569 ( .A(b[2801]), .B(n7272), .Z(n7273) );
  XNOR U8570 ( .A(b[2801]), .B(n7274), .Z(c[2801]) );
  XNOR U8571 ( .A(a[2801]), .B(n7275), .Z(n7274) );
  IV U8572 ( .A(n7272), .Z(n7275) );
  XOR U8573 ( .A(n7276), .B(n7277), .Z(n7272) );
  ANDN U8574 ( .B(n7278), .A(n7279), .Z(n7276) );
  XNOR U8575 ( .A(b[2800]), .B(n7277), .Z(n7278) );
  XNOR U8576 ( .A(b[2800]), .B(n7279), .Z(c[2800]) );
  XNOR U8577 ( .A(a[2800]), .B(n7280), .Z(n7279) );
  IV U8578 ( .A(n7277), .Z(n7280) );
  XOR U8579 ( .A(n7281), .B(n7282), .Z(n7277) );
  ANDN U8580 ( .B(n7283), .A(n7284), .Z(n7281) );
  XNOR U8581 ( .A(b[2799]), .B(n7282), .Z(n7283) );
  XNOR U8582 ( .A(b[27]), .B(n7285), .Z(c[27]) );
  XNOR U8583 ( .A(b[279]), .B(n7286), .Z(c[279]) );
  XNOR U8584 ( .A(b[2799]), .B(n7284), .Z(c[2799]) );
  XNOR U8585 ( .A(a[2799]), .B(n7287), .Z(n7284) );
  IV U8586 ( .A(n7282), .Z(n7287) );
  XOR U8587 ( .A(n7288), .B(n7289), .Z(n7282) );
  ANDN U8588 ( .B(n7290), .A(n7291), .Z(n7288) );
  XNOR U8589 ( .A(b[2798]), .B(n7289), .Z(n7290) );
  XNOR U8590 ( .A(b[2798]), .B(n7291), .Z(c[2798]) );
  XNOR U8591 ( .A(a[2798]), .B(n7292), .Z(n7291) );
  IV U8592 ( .A(n7289), .Z(n7292) );
  XOR U8593 ( .A(n7293), .B(n7294), .Z(n7289) );
  ANDN U8594 ( .B(n7295), .A(n7296), .Z(n7293) );
  XNOR U8595 ( .A(b[2797]), .B(n7294), .Z(n7295) );
  XNOR U8596 ( .A(b[2797]), .B(n7296), .Z(c[2797]) );
  XNOR U8597 ( .A(a[2797]), .B(n7297), .Z(n7296) );
  IV U8598 ( .A(n7294), .Z(n7297) );
  XOR U8599 ( .A(n7298), .B(n7299), .Z(n7294) );
  ANDN U8600 ( .B(n7300), .A(n7301), .Z(n7298) );
  XNOR U8601 ( .A(b[2796]), .B(n7299), .Z(n7300) );
  XNOR U8602 ( .A(b[2796]), .B(n7301), .Z(c[2796]) );
  XNOR U8603 ( .A(a[2796]), .B(n7302), .Z(n7301) );
  IV U8604 ( .A(n7299), .Z(n7302) );
  XOR U8605 ( .A(n7303), .B(n7304), .Z(n7299) );
  ANDN U8606 ( .B(n7305), .A(n7306), .Z(n7303) );
  XNOR U8607 ( .A(b[2795]), .B(n7304), .Z(n7305) );
  XNOR U8608 ( .A(b[2795]), .B(n7306), .Z(c[2795]) );
  XNOR U8609 ( .A(a[2795]), .B(n7307), .Z(n7306) );
  IV U8610 ( .A(n7304), .Z(n7307) );
  XOR U8611 ( .A(n7308), .B(n7309), .Z(n7304) );
  ANDN U8612 ( .B(n7310), .A(n7311), .Z(n7308) );
  XNOR U8613 ( .A(b[2794]), .B(n7309), .Z(n7310) );
  XNOR U8614 ( .A(b[2794]), .B(n7311), .Z(c[2794]) );
  XNOR U8615 ( .A(a[2794]), .B(n7312), .Z(n7311) );
  IV U8616 ( .A(n7309), .Z(n7312) );
  XOR U8617 ( .A(n7313), .B(n7314), .Z(n7309) );
  ANDN U8618 ( .B(n7315), .A(n7316), .Z(n7313) );
  XNOR U8619 ( .A(b[2793]), .B(n7314), .Z(n7315) );
  XNOR U8620 ( .A(b[2793]), .B(n7316), .Z(c[2793]) );
  XNOR U8621 ( .A(a[2793]), .B(n7317), .Z(n7316) );
  IV U8622 ( .A(n7314), .Z(n7317) );
  XOR U8623 ( .A(n7318), .B(n7319), .Z(n7314) );
  ANDN U8624 ( .B(n7320), .A(n7321), .Z(n7318) );
  XNOR U8625 ( .A(b[2792]), .B(n7319), .Z(n7320) );
  XNOR U8626 ( .A(b[2792]), .B(n7321), .Z(c[2792]) );
  XNOR U8627 ( .A(a[2792]), .B(n7322), .Z(n7321) );
  IV U8628 ( .A(n7319), .Z(n7322) );
  XOR U8629 ( .A(n7323), .B(n7324), .Z(n7319) );
  ANDN U8630 ( .B(n7325), .A(n7326), .Z(n7323) );
  XNOR U8631 ( .A(b[2791]), .B(n7324), .Z(n7325) );
  XNOR U8632 ( .A(b[2791]), .B(n7326), .Z(c[2791]) );
  XNOR U8633 ( .A(a[2791]), .B(n7327), .Z(n7326) );
  IV U8634 ( .A(n7324), .Z(n7327) );
  XOR U8635 ( .A(n7328), .B(n7329), .Z(n7324) );
  ANDN U8636 ( .B(n7330), .A(n7331), .Z(n7328) );
  XNOR U8637 ( .A(b[2790]), .B(n7329), .Z(n7330) );
  XNOR U8638 ( .A(b[2790]), .B(n7331), .Z(c[2790]) );
  XNOR U8639 ( .A(a[2790]), .B(n7332), .Z(n7331) );
  IV U8640 ( .A(n7329), .Z(n7332) );
  XOR U8641 ( .A(n7333), .B(n7334), .Z(n7329) );
  ANDN U8642 ( .B(n7335), .A(n7336), .Z(n7333) );
  XNOR U8643 ( .A(b[2789]), .B(n7334), .Z(n7335) );
  XNOR U8644 ( .A(b[278]), .B(n7337), .Z(c[278]) );
  XNOR U8645 ( .A(b[2789]), .B(n7336), .Z(c[2789]) );
  XNOR U8646 ( .A(a[2789]), .B(n7338), .Z(n7336) );
  IV U8647 ( .A(n7334), .Z(n7338) );
  XOR U8648 ( .A(n7339), .B(n7340), .Z(n7334) );
  ANDN U8649 ( .B(n7341), .A(n7342), .Z(n7339) );
  XNOR U8650 ( .A(b[2788]), .B(n7340), .Z(n7341) );
  XNOR U8651 ( .A(b[2788]), .B(n7342), .Z(c[2788]) );
  XNOR U8652 ( .A(a[2788]), .B(n7343), .Z(n7342) );
  IV U8653 ( .A(n7340), .Z(n7343) );
  XOR U8654 ( .A(n7344), .B(n7345), .Z(n7340) );
  ANDN U8655 ( .B(n7346), .A(n7347), .Z(n7344) );
  XNOR U8656 ( .A(b[2787]), .B(n7345), .Z(n7346) );
  XNOR U8657 ( .A(b[2787]), .B(n7347), .Z(c[2787]) );
  XNOR U8658 ( .A(a[2787]), .B(n7348), .Z(n7347) );
  IV U8659 ( .A(n7345), .Z(n7348) );
  XOR U8660 ( .A(n7349), .B(n7350), .Z(n7345) );
  ANDN U8661 ( .B(n7351), .A(n7352), .Z(n7349) );
  XNOR U8662 ( .A(b[2786]), .B(n7350), .Z(n7351) );
  XNOR U8663 ( .A(b[2786]), .B(n7352), .Z(c[2786]) );
  XNOR U8664 ( .A(a[2786]), .B(n7353), .Z(n7352) );
  IV U8665 ( .A(n7350), .Z(n7353) );
  XOR U8666 ( .A(n7354), .B(n7355), .Z(n7350) );
  ANDN U8667 ( .B(n7356), .A(n7357), .Z(n7354) );
  XNOR U8668 ( .A(b[2785]), .B(n7355), .Z(n7356) );
  XNOR U8669 ( .A(b[2785]), .B(n7357), .Z(c[2785]) );
  XNOR U8670 ( .A(a[2785]), .B(n7358), .Z(n7357) );
  IV U8671 ( .A(n7355), .Z(n7358) );
  XOR U8672 ( .A(n7359), .B(n7360), .Z(n7355) );
  ANDN U8673 ( .B(n7361), .A(n7362), .Z(n7359) );
  XNOR U8674 ( .A(b[2784]), .B(n7360), .Z(n7361) );
  XNOR U8675 ( .A(b[2784]), .B(n7362), .Z(c[2784]) );
  XNOR U8676 ( .A(a[2784]), .B(n7363), .Z(n7362) );
  IV U8677 ( .A(n7360), .Z(n7363) );
  XOR U8678 ( .A(n7364), .B(n7365), .Z(n7360) );
  ANDN U8679 ( .B(n7366), .A(n7367), .Z(n7364) );
  XNOR U8680 ( .A(b[2783]), .B(n7365), .Z(n7366) );
  XNOR U8681 ( .A(b[2783]), .B(n7367), .Z(c[2783]) );
  XNOR U8682 ( .A(a[2783]), .B(n7368), .Z(n7367) );
  IV U8683 ( .A(n7365), .Z(n7368) );
  XOR U8684 ( .A(n7369), .B(n7370), .Z(n7365) );
  ANDN U8685 ( .B(n7371), .A(n7372), .Z(n7369) );
  XNOR U8686 ( .A(b[2782]), .B(n7370), .Z(n7371) );
  XNOR U8687 ( .A(b[2782]), .B(n7372), .Z(c[2782]) );
  XNOR U8688 ( .A(a[2782]), .B(n7373), .Z(n7372) );
  IV U8689 ( .A(n7370), .Z(n7373) );
  XOR U8690 ( .A(n7374), .B(n7375), .Z(n7370) );
  ANDN U8691 ( .B(n7376), .A(n7377), .Z(n7374) );
  XNOR U8692 ( .A(b[2781]), .B(n7375), .Z(n7376) );
  XNOR U8693 ( .A(b[2781]), .B(n7377), .Z(c[2781]) );
  XNOR U8694 ( .A(a[2781]), .B(n7378), .Z(n7377) );
  IV U8695 ( .A(n7375), .Z(n7378) );
  XOR U8696 ( .A(n7379), .B(n7380), .Z(n7375) );
  ANDN U8697 ( .B(n7381), .A(n7382), .Z(n7379) );
  XNOR U8698 ( .A(b[2780]), .B(n7380), .Z(n7381) );
  XNOR U8699 ( .A(b[2780]), .B(n7382), .Z(c[2780]) );
  XNOR U8700 ( .A(a[2780]), .B(n7383), .Z(n7382) );
  IV U8701 ( .A(n7380), .Z(n7383) );
  XOR U8702 ( .A(n7384), .B(n7385), .Z(n7380) );
  ANDN U8703 ( .B(n7386), .A(n7387), .Z(n7384) );
  XNOR U8704 ( .A(b[2779]), .B(n7385), .Z(n7386) );
  XNOR U8705 ( .A(b[277]), .B(n7388), .Z(c[277]) );
  XNOR U8706 ( .A(b[2779]), .B(n7387), .Z(c[2779]) );
  XNOR U8707 ( .A(a[2779]), .B(n7389), .Z(n7387) );
  IV U8708 ( .A(n7385), .Z(n7389) );
  XOR U8709 ( .A(n7390), .B(n7391), .Z(n7385) );
  ANDN U8710 ( .B(n7392), .A(n7393), .Z(n7390) );
  XNOR U8711 ( .A(b[2778]), .B(n7391), .Z(n7392) );
  XNOR U8712 ( .A(b[2778]), .B(n7393), .Z(c[2778]) );
  XNOR U8713 ( .A(a[2778]), .B(n7394), .Z(n7393) );
  IV U8714 ( .A(n7391), .Z(n7394) );
  XOR U8715 ( .A(n7395), .B(n7396), .Z(n7391) );
  ANDN U8716 ( .B(n7397), .A(n7398), .Z(n7395) );
  XNOR U8717 ( .A(b[2777]), .B(n7396), .Z(n7397) );
  XNOR U8718 ( .A(b[2777]), .B(n7398), .Z(c[2777]) );
  XNOR U8719 ( .A(a[2777]), .B(n7399), .Z(n7398) );
  IV U8720 ( .A(n7396), .Z(n7399) );
  XOR U8721 ( .A(n7400), .B(n7401), .Z(n7396) );
  ANDN U8722 ( .B(n7402), .A(n7403), .Z(n7400) );
  XNOR U8723 ( .A(b[2776]), .B(n7401), .Z(n7402) );
  XNOR U8724 ( .A(b[2776]), .B(n7403), .Z(c[2776]) );
  XNOR U8725 ( .A(a[2776]), .B(n7404), .Z(n7403) );
  IV U8726 ( .A(n7401), .Z(n7404) );
  XOR U8727 ( .A(n7405), .B(n7406), .Z(n7401) );
  ANDN U8728 ( .B(n7407), .A(n7408), .Z(n7405) );
  XNOR U8729 ( .A(b[2775]), .B(n7406), .Z(n7407) );
  XNOR U8730 ( .A(b[2775]), .B(n7408), .Z(c[2775]) );
  XNOR U8731 ( .A(a[2775]), .B(n7409), .Z(n7408) );
  IV U8732 ( .A(n7406), .Z(n7409) );
  XOR U8733 ( .A(n7410), .B(n7411), .Z(n7406) );
  ANDN U8734 ( .B(n7412), .A(n7413), .Z(n7410) );
  XNOR U8735 ( .A(b[2774]), .B(n7411), .Z(n7412) );
  XNOR U8736 ( .A(b[2774]), .B(n7413), .Z(c[2774]) );
  XNOR U8737 ( .A(a[2774]), .B(n7414), .Z(n7413) );
  IV U8738 ( .A(n7411), .Z(n7414) );
  XOR U8739 ( .A(n7415), .B(n7416), .Z(n7411) );
  ANDN U8740 ( .B(n7417), .A(n7418), .Z(n7415) );
  XNOR U8741 ( .A(b[2773]), .B(n7416), .Z(n7417) );
  XNOR U8742 ( .A(b[2773]), .B(n7418), .Z(c[2773]) );
  XNOR U8743 ( .A(a[2773]), .B(n7419), .Z(n7418) );
  IV U8744 ( .A(n7416), .Z(n7419) );
  XOR U8745 ( .A(n7420), .B(n7421), .Z(n7416) );
  ANDN U8746 ( .B(n7422), .A(n7423), .Z(n7420) );
  XNOR U8747 ( .A(b[2772]), .B(n7421), .Z(n7422) );
  XNOR U8748 ( .A(b[2772]), .B(n7423), .Z(c[2772]) );
  XNOR U8749 ( .A(a[2772]), .B(n7424), .Z(n7423) );
  IV U8750 ( .A(n7421), .Z(n7424) );
  XOR U8751 ( .A(n7425), .B(n7426), .Z(n7421) );
  ANDN U8752 ( .B(n7427), .A(n7428), .Z(n7425) );
  XNOR U8753 ( .A(b[2771]), .B(n7426), .Z(n7427) );
  XNOR U8754 ( .A(b[2771]), .B(n7428), .Z(c[2771]) );
  XNOR U8755 ( .A(a[2771]), .B(n7429), .Z(n7428) );
  IV U8756 ( .A(n7426), .Z(n7429) );
  XOR U8757 ( .A(n7430), .B(n7431), .Z(n7426) );
  ANDN U8758 ( .B(n7432), .A(n7433), .Z(n7430) );
  XNOR U8759 ( .A(b[2770]), .B(n7431), .Z(n7432) );
  XNOR U8760 ( .A(b[2770]), .B(n7433), .Z(c[2770]) );
  XNOR U8761 ( .A(a[2770]), .B(n7434), .Z(n7433) );
  IV U8762 ( .A(n7431), .Z(n7434) );
  XOR U8763 ( .A(n7435), .B(n7436), .Z(n7431) );
  ANDN U8764 ( .B(n7437), .A(n7438), .Z(n7435) );
  XNOR U8765 ( .A(b[2769]), .B(n7436), .Z(n7437) );
  XNOR U8766 ( .A(b[276]), .B(n7439), .Z(c[276]) );
  XNOR U8767 ( .A(b[2769]), .B(n7438), .Z(c[2769]) );
  XNOR U8768 ( .A(a[2769]), .B(n7440), .Z(n7438) );
  IV U8769 ( .A(n7436), .Z(n7440) );
  XOR U8770 ( .A(n7441), .B(n7442), .Z(n7436) );
  ANDN U8771 ( .B(n7443), .A(n7444), .Z(n7441) );
  XNOR U8772 ( .A(b[2768]), .B(n7442), .Z(n7443) );
  XNOR U8773 ( .A(b[2768]), .B(n7444), .Z(c[2768]) );
  XNOR U8774 ( .A(a[2768]), .B(n7445), .Z(n7444) );
  IV U8775 ( .A(n7442), .Z(n7445) );
  XOR U8776 ( .A(n7446), .B(n7447), .Z(n7442) );
  ANDN U8777 ( .B(n7448), .A(n7449), .Z(n7446) );
  XNOR U8778 ( .A(b[2767]), .B(n7447), .Z(n7448) );
  XNOR U8779 ( .A(b[2767]), .B(n7449), .Z(c[2767]) );
  XNOR U8780 ( .A(a[2767]), .B(n7450), .Z(n7449) );
  IV U8781 ( .A(n7447), .Z(n7450) );
  XOR U8782 ( .A(n7451), .B(n7452), .Z(n7447) );
  ANDN U8783 ( .B(n7453), .A(n7454), .Z(n7451) );
  XNOR U8784 ( .A(b[2766]), .B(n7452), .Z(n7453) );
  XNOR U8785 ( .A(b[2766]), .B(n7454), .Z(c[2766]) );
  XNOR U8786 ( .A(a[2766]), .B(n7455), .Z(n7454) );
  IV U8787 ( .A(n7452), .Z(n7455) );
  XOR U8788 ( .A(n7456), .B(n7457), .Z(n7452) );
  ANDN U8789 ( .B(n7458), .A(n7459), .Z(n7456) );
  XNOR U8790 ( .A(b[2765]), .B(n7457), .Z(n7458) );
  XNOR U8791 ( .A(b[2765]), .B(n7459), .Z(c[2765]) );
  XNOR U8792 ( .A(a[2765]), .B(n7460), .Z(n7459) );
  IV U8793 ( .A(n7457), .Z(n7460) );
  XOR U8794 ( .A(n7461), .B(n7462), .Z(n7457) );
  ANDN U8795 ( .B(n7463), .A(n7464), .Z(n7461) );
  XNOR U8796 ( .A(b[2764]), .B(n7462), .Z(n7463) );
  XNOR U8797 ( .A(b[2764]), .B(n7464), .Z(c[2764]) );
  XNOR U8798 ( .A(a[2764]), .B(n7465), .Z(n7464) );
  IV U8799 ( .A(n7462), .Z(n7465) );
  XOR U8800 ( .A(n7466), .B(n7467), .Z(n7462) );
  ANDN U8801 ( .B(n7468), .A(n7469), .Z(n7466) );
  XNOR U8802 ( .A(b[2763]), .B(n7467), .Z(n7468) );
  XNOR U8803 ( .A(b[2763]), .B(n7469), .Z(c[2763]) );
  XNOR U8804 ( .A(a[2763]), .B(n7470), .Z(n7469) );
  IV U8805 ( .A(n7467), .Z(n7470) );
  XOR U8806 ( .A(n7471), .B(n7472), .Z(n7467) );
  ANDN U8807 ( .B(n7473), .A(n7474), .Z(n7471) );
  XNOR U8808 ( .A(b[2762]), .B(n7472), .Z(n7473) );
  XNOR U8809 ( .A(b[2762]), .B(n7474), .Z(c[2762]) );
  XNOR U8810 ( .A(a[2762]), .B(n7475), .Z(n7474) );
  IV U8811 ( .A(n7472), .Z(n7475) );
  XOR U8812 ( .A(n7476), .B(n7477), .Z(n7472) );
  ANDN U8813 ( .B(n7478), .A(n7479), .Z(n7476) );
  XNOR U8814 ( .A(b[2761]), .B(n7477), .Z(n7478) );
  XNOR U8815 ( .A(b[2761]), .B(n7479), .Z(c[2761]) );
  XNOR U8816 ( .A(a[2761]), .B(n7480), .Z(n7479) );
  IV U8817 ( .A(n7477), .Z(n7480) );
  XOR U8818 ( .A(n7481), .B(n7482), .Z(n7477) );
  ANDN U8819 ( .B(n7483), .A(n7484), .Z(n7481) );
  XNOR U8820 ( .A(b[2760]), .B(n7482), .Z(n7483) );
  XNOR U8821 ( .A(b[2760]), .B(n7484), .Z(c[2760]) );
  XNOR U8822 ( .A(a[2760]), .B(n7485), .Z(n7484) );
  IV U8823 ( .A(n7482), .Z(n7485) );
  XOR U8824 ( .A(n7486), .B(n7487), .Z(n7482) );
  ANDN U8825 ( .B(n7488), .A(n7489), .Z(n7486) );
  XNOR U8826 ( .A(b[2759]), .B(n7487), .Z(n7488) );
  XNOR U8827 ( .A(b[275]), .B(n7490), .Z(c[275]) );
  XNOR U8828 ( .A(b[2759]), .B(n7489), .Z(c[2759]) );
  XNOR U8829 ( .A(a[2759]), .B(n7491), .Z(n7489) );
  IV U8830 ( .A(n7487), .Z(n7491) );
  XOR U8831 ( .A(n7492), .B(n7493), .Z(n7487) );
  ANDN U8832 ( .B(n7494), .A(n7495), .Z(n7492) );
  XNOR U8833 ( .A(b[2758]), .B(n7493), .Z(n7494) );
  XNOR U8834 ( .A(b[2758]), .B(n7495), .Z(c[2758]) );
  XNOR U8835 ( .A(a[2758]), .B(n7496), .Z(n7495) );
  IV U8836 ( .A(n7493), .Z(n7496) );
  XOR U8837 ( .A(n7497), .B(n7498), .Z(n7493) );
  ANDN U8838 ( .B(n7499), .A(n7500), .Z(n7497) );
  XNOR U8839 ( .A(b[2757]), .B(n7498), .Z(n7499) );
  XNOR U8840 ( .A(b[2757]), .B(n7500), .Z(c[2757]) );
  XNOR U8841 ( .A(a[2757]), .B(n7501), .Z(n7500) );
  IV U8842 ( .A(n7498), .Z(n7501) );
  XOR U8843 ( .A(n7502), .B(n7503), .Z(n7498) );
  ANDN U8844 ( .B(n7504), .A(n7505), .Z(n7502) );
  XNOR U8845 ( .A(b[2756]), .B(n7503), .Z(n7504) );
  XNOR U8846 ( .A(b[2756]), .B(n7505), .Z(c[2756]) );
  XNOR U8847 ( .A(a[2756]), .B(n7506), .Z(n7505) );
  IV U8848 ( .A(n7503), .Z(n7506) );
  XOR U8849 ( .A(n7507), .B(n7508), .Z(n7503) );
  ANDN U8850 ( .B(n7509), .A(n7510), .Z(n7507) );
  XNOR U8851 ( .A(b[2755]), .B(n7508), .Z(n7509) );
  XNOR U8852 ( .A(b[2755]), .B(n7510), .Z(c[2755]) );
  XNOR U8853 ( .A(a[2755]), .B(n7511), .Z(n7510) );
  IV U8854 ( .A(n7508), .Z(n7511) );
  XOR U8855 ( .A(n7512), .B(n7513), .Z(n7508) );
  ANDN U8856 ( .B(n7514), .A(n7515), .Z(n7512) );
  XNOR U8857 ( .A(b[2754]), .B(n7513), .Z(n7514) );
  XNOR U8858 ( .A(b[2754]), .B(n7515), .Z(c[2754]) );
  XNOR U8859 ( .A(a[2754]), .B(n7516), .Z(n7515) );
  IV U8860 ( .A(n7513), .Z(n7516) );
  XOR U8861 ( .A(n7517), .B(n7518), .Z(n7513) );
  ANDN U8862 ( .B(n7519), .A(n7520), .Z(n7517) );
  XNOR U8863 ( .A(b[2753]), .B(n7518), .Z(n7519) );
  XNOR U8864 ( .A(b[2753]), .B(n7520), .Z(c[2753]) );
  XNOR U8865 ( .A(a[2753]), .B(n7521), .Z(n7520) );
  IV U8866 ( .A(n7518), .Z(n7521) );
  XOR U8867 ( .A(n7522), .B(n7523), .Z(n7518) );
  ANDN U8868 ( .B(n7524), .A(n7525), .Z(n7522) );
  XNOR U8869 ( .A(b[2752]), .B(n7523), .Z(n7524) );
  XNOR U8870 ( .A(b[2752]), .B(n7525), .Z(c[2752]) );
  XNOR U8871 ( .A(a[2752]), .B(n7526), .Z(n7525) );
  IV U8872 ( .A(n7523), .Z(n7526) );
  XOR U8873 ( .A(n7527), .B(n7528), .Z(n7523) );
  ANDN U8874 ( .B(n7529), .A(n7530), .Z(n7527) );
  XNOR U8875 ( .A(b[2751]), .B(n7528), .Z(n7529) );
  XNOR U8876 ( .A(b[2751]), .B(n7530), .Z(c[2751]) );
  XNOR U8877 ( .A(a[2751]), .B(n7531), .Z(n7530) );
  IV U8878 ( .A(n7528), .Z(n7531) );
  XOR U8879 ( .A(n7532), .B(n7533), .Z(n7528) );
  ANDN U8880 ( .B(n7534), .A(n7535), .Z(n7532) );
  XNOR U8881 ( .A(b[2750]), .B(n7533), .Z(n7534) );
  XNOR U8882 ( .A(b[2750]), .B(n7535), .Z(c[2750]) );
  XNOR U8883 ( .A(a[2750]), .B(n7536), .Z(n7535) );
  IV U8884 ( .A(n7533), .Z(n7536) );
  XOR U8885 ( .A(n7537), .B(n7538), .Z(n7533) );
  ANDN U8886 ( .B(n7539), .A(n7540), .Z(n7537) );
  XNOR U8887 ( .A(b[2749]), .B(n7538), .Z(n7539) );
  XNOR U8888 ( .A(b[274]), .B(n7541), .Z(c[274]) );
  XNOR U8889 ( .A(b[2749]), .B(n7540), .Z(c[2749]) );
  XNOR U8890 ( .A(a[2749]), .B(n7542), .Z(n7540) );
  IV U8891 ( .A(n7538), .Z(n7542) );
  XOR U8892 ( .A(n7543), .B(n7544), .Z(n7538) );
  ANDN U8893 ( .B(n7545), .A(n7546), .Z(n7543) );
  XNOR U8894 ( .A(b[2748]), .B(n7544), .Z(n7545) );
  XNOR U8895 ( .A(b[2748]), .B(n7546), .Z(c[2748]) );
  XNOR U8896 ( .A(a[2748]), .B(n7547), .Z(n7546) );
  IV U8897 ( .A(n7544), .Z(n7547) );
  XOR U8898 ( .A(n7548), .B(n7549), .Z(n7544) );
  ANDN U8899 ( .B(n7550), .A(n7551), .Z(n7548) );
  XNOR U8900 ( .A(b[2747]), .B(n7549), .Z(n7550) );
  XNOR U8901 ( .A(b[2747]), .B(n7551), .Z(c[2747]) );
  XNOR U8902 ( .A(a[2747]), .B(n7552), .Z(n7551) );
  IV U8903 ( .A(n7549), .Z(n7552) );
  XOR U8904 ( .A(n7553), .B(n7554), .Z(n7549) );
  ANDN U8905 ( .B(n7555), .A(n7556), .Z(n7553) );
  XNOR U8906 ( .A(b[2746]), .B(n7554), .Z(n7555) );
  XNOR U8907 ( .A(b[2746]), .B(n7556), .Z(c[2746]) );
  XNOR U8908 ( .A(a[2746]), .B(n7557), .Z(n7556) );
  IV U8909 ( .A(n7554), .Z(n7557) );
  XOR U8910 ( .A(n7558), .B(n7559), .Z(n7554) );
  ANDN U8911 ( .B(n7560), .A(n7561), .Z(n7558) );
  XNOR U8912 ( .A(b[2745]), .B(n7559), .Z(n7560) );
  XNOR U8913 ( .A(b[2745]), .B(n7561), .Z(c[2745]) );
  XNOR U8914 ( .A(a[2745]), .B(n7562), .Z(n7561) );
  IV U8915 ( .A(n7559), .Z(n7562) );
  XOR U8916 ( .A(n7563), .B(n7564), .Z(n7559) );
  ANDN U8917 ( .B(n7565), .A(n7566), .Z(n7563) );
  XNOR U8918 ( .A(b[2744]), .B(n7564), .Z(n7565) );
  XNOR U8919 ( .A(b[2744]), .B(n7566), .Z(c[2744]) );
  XNOR U8920 ( .A(a[2744]), .B(n7567), .Z(n7566) );
  IV U8921 ( .A(n7564), .Z(n7567) );
  XOR U8922 ( .A(n7568), .B(n7569), .Z(n7564) );
  ANDN U8923 ( .B(n7570), .A(n7571), .Z(n7568) );
  XNOR U8924 ( .A(b[2743]), .B(n7569), .Z(n7570) );
  XNOR U8925 ( .A(b[2743]), .B(n7571), .Z(c[2743]) );
  XNOR U8926 ( .A(a[2743]), .B(n7572), .Z(n7571) );
  IV U8927 ( .A(n7569), .Z(n7572) );
  XOR U8928 ( .A(n7573), .B(n7574), .Z(n7569) );
  ANDN U8929 ( .B(n7575), .A(n7576), .Z(n7573) );
  XNOR U8930 ( .A(b[2742]), .B(n7574), .Z(n7575) );
  XNOR U8931 ( .A(b[2742]), .B(n7576), .Z(c[2742]) );
  XNOR U8932 ( .A(a[2742]), .B(n7577), .Z(n7576) );
  IV U8933 ( .A(n7574), .Z(n7577) );
  XOR U8934 ( .A(n7578), .B(n7579), .Z(n7574) );
  ANDN U8935 ( .B(n7580), .A(n7581), .Z(n7578) );
  XNOR U8936 ( .A(b[2741]), .B(n7579), .Z(n7580) );
  XNOR U8937 ( .A(b[2741]), .B(n7581), .Z(c[2741]) );
  XNOR U8938 ( .A(a[2741]), .B(n7582), .Z(n7581) );
  IV U8939 ( .A(n7579), .Z(n7582) );
  XOR U8940 ( .A(n7583), .B(n7584), .Z(n7579) );
  ANDN U8941 ( .B(n7585), .A(n7586), .Z(n7583) );
  XNOR U8942 ( .A(b[2740]), .B(n7584), .Z(n7585) );
  XNOR U8943 ( .A(b[2740]), .B(n7586), .Z(c[2740]) );
  XNOR U8944 ( .A(a[2740]), .B(n7587), .Z(n7586) );
  IV U8945 ( .A(n7584), .Z(n7587) );
  XOR U8946 ( .A(n7588), .B(n7589), .Z(n7584) );
  ANDN U8947 ( .B(n7590), .A(n7591), .Z(n7588) );
  XNOR U8948 ( .A(b[2739]), .B(n7589), .Z(n7590) );
  XNOR U8949 ( .A(b[273]), .B(n7592), .Z(c[273]) );
  XNOR U8950 ( .A(b[2739]), .B(n7591), .Z(c[2739]) );
  XNOR U8951 ( .A(a[2739]), .B(n7593), .Z(n7591) );
  IV U8952 ( .A(n7589), .Z(n7593) );
  XOR U8953 ( .A(n7594), .B(n7595), .Z(n7589) );
  ANDN U8954 ( .B(n7596), .A(n7597), .Z(n7594) );
  XNOR U8955 ( .A(b[2738]), .B(n7595), .Z(n7596) );
  XNOR U8956 ( .A(b[2738]), .B(n7597), .Z(c[2738]) );
  XNOR U8957 ( .A(a[2738]), .B(n7598), .Z(n7597) );
  IV U8958 ( .A(n7595), .Z(n7598) );
  XOR U8959 ( .A(n7599), .B(n7600), .Z(n7595) );
  ANDN U8960 ( .B(n7601), .A(n7602), .Z(n7599) );
  XNOR U8961 ( .A(b[2737]), .B(n7600), .Z(n7601) );
  XNOR U8962 ( .A(b[2737]), .B(n7602), .Z(c[2737]) );
  XNOR U8963 ( .A(a[2737]), .B(n7603), .Z(n7602) );
  IV U8964 ( .A(n7600), .Z(n7603) );
  XOR U8965 ( .A(n7604), .B(n7605), .Z(n7600) );
  ANDN U8966 ( .B(n7606), .A(n7607), .Z(n7604) );
  XNOR U8967 ( .A(b[2736]), .B(n7605), .Z(n7606) );
  XNOR U8968 ( .A(b[2736]), .B(n7607), .Z(c[2736]) );
  XNOR U8969 ( .A(a[2736]), .B(n7608), .Z(n7607) );
  IV U8970 ( .A(n7605), .Z(n7608) );
  XOR U8971 ( .A(n7609), .B(n7610), .Z(n7605) );
  ANDN U8972 ( .B(n7611), .A(n7612), .Z(n7609) );
  XNOR U8973 ( .A(b[2735]), .B(n7610), .Z(n7611) );
  XNOR U8974 ( .A(b[2735]), .B(n7612), .Z(c[2735]) );
  XNOR U8975 ( .A(a[2735]), .B(n7613), .Z(n7612) );
  IV U8976 ( .A(n7610), .Z(n7613) );
  XOR U8977 ( .A(n7614), .B(n7615), .Z(n7610) );
  ANDN U8978 ( .B(n7616), .A(n7617), .Z(n7614) );
  XNOR U8979 ( .A(b[2734]), .B(n7615), .Z(n7616) );
  XNOR U8980 ( .A(b[2734]), .B(n7617), .Z(c[2734]) );
  XNOR U8981 ( .A(a[2734]), .B(n7618), .Z(n7617) );
  IV U8982 ( .A(n7615), .Z(n7618) );
  XOR U8983 ( .A(n7619), .B(n7620), .Z(n7615) );
  ANDN U8984 ( .B(n7621), .A(n7622), .Z(n7619) );
  XNOR U8985 ( .A(b[2733]), .B(n7620), .Z(n7621) );
  XNOR U8986 ( .A(b[2733]), .B(n7622), .Z(c[2733]) );
  XNOR U8987 ( .A(a[2733]), .B(n7623), .Z(n7622) );
  IV U8988 ( .A(n7620), .Z(n7623) );
  XOR U8989 ( .A(n7624), .B(n7625), .Z(n7620) );
  ANDN U8990 ( .B(n7626), .A(n7627), .Z(n7624) );
  XNOR U8991 ( .A(b[2732]), .B(n7625), .Z(n7626) );
  XNOR U8992 ( .A(b[2732]), .B(n7627), .Z(c[2732]) );
  XNOR U8993 ( .A(a[2732]), .B(n7628), .Z(n7627) );
  IV U8994 ( .A(n7625), .Z(n7628) );
  XOR U8995 ( .A(n7629), .B(n7630), .Z(n7625) );
  ANDN U8996 ( .B(n7631), .A(n7632), .Z(n7629) );
  XNOR U8997 ( .A(b[2731]), .B(n7630), .Z(n7631) );
  XNOR U8998 ( .A(b[2731]), .B(n7632), .Z(c[2731]) );
  XNOR U8999 ( .A(a[2731]), .B(n7633), .Z(n7632) );
  IV U9000 ( .A(n7630), .Z(n7633) );
  XOR U9001 ( .A(n7634), .B(n7635), .Z(n7630) );
  ANDN U9002 ( .B(n7636), .A(n7637), .Z(n7634) );
  XNOR U9003 ( .A(b[2730]), .B(n7635), .Z(n7636) );
  XNOR U9004 ( .A(b[2730]), .B(n7637), .Z(c[2730]) );
  XNOR U9005 ( .A(a[2730]), .B(n7638), .Z(n7637) );
  IV U9006 ( .A(n7635), .Z(n7638) );
  XOR U9007 ( .A(n7639), .B(n7640), .Z(n7635) );
  ANDN U9008 ( .B(n7641), .A(n7642), .Z(n7639) );
  XNOR U9009 ( .A(b[2729]), .B(n7640), .Z(n7641) );
  XNOR U9010 ( .A(b[272]), .B(n7643), .Z(c[272]) );
  XNOR U9011 ( .A(b[2729]), .B(n7642), .Z(c[2729]) );
  XNOR U9012 ( .A(a[2729]), .B(n7644), .Z(n7642) );
  IV U9013 ( .A(n7640), .Z(n7644) );
  XOR U9014 ( .A(n7645), .B(n7646), .Z(n7640) );
  ANDN U9015 ( .B(n7647), .A(n7648), .Z(n7645) );
  XNOR U9016 ( .A(b[2728]), .B(n7646), .Z(n7647) );
  XNOR U9017 ( .A(b[2728]), .B(n7648), .Z(c[2728]) );
  XNOR U9018 ( .A(a[2728]), .B(n7649), .Z(n7648) );
  IV U9019 ( .A(n7646), .Z(n7649) );
  XOR U9020 ( .A(n7650), .B(n7651), .Z(n7646) );
  ANDN U9021 ( .B(n7652), .A(n7653), .Z(n7650) );
  XNOR U9022 ( .A(b[2727]), .B(n7651), .Z(n7652) );
  XNOR U9023 ( .A(b[2727]), .B(n7653), .Z(c[2727]) );
  XNOR U9024 ( .A(a[2727]), .B(n7654), .Z(n7653) );
  IV U9025 ( .A(n7651), .Z(n7654) );
  XOR U9026 ( .A(n7655), .B(n7656), .Z(n7651) );
  ANDN U9027 ( .B(n7657), .A(n7658), .Z(n7655) );
  XNOR U9028 ( .A(b[2726]), .B(n7656), .Z(n7657) );
  XNOR U9029 ( .A(b[2726]), .B(n7658), .Z(c[2726]) );
  XNOR U9030 ( .A(a[2726]), .B(n7659), .Z(n7658) );
  IV U9031 ( .A(n7656), .Z(n7659) );
  XOR U9032 ( .A(n7660), .B(n7661), .Z(n7656) );
  ANDN U9033 ( .B(n7662), .A(n7663), .Z(n7660) );
  XNOR U9034 ( .A(b[2725]), .B(n7661), .Z(n7662) );
  XNOR U9035 ( .A(b[2725]), .B(n7663), .Z(c[2725]) );
  XNOR U9036 ( .A(a[2725]), .B(n7664), .Z(n7663) );
  IV U9037 ( .A(n7661), .Z(n7664) );
  XOR U9038 ( .A(n7665), .B(n7666), .Z(n7661) );
  ANDN U9039 ( .B(n7667), .A(n7668), .Z(n7665) );
  XNOR U9040 ( .A(b[2724]), .B(n7666), .Z(n7667) );
  XNOR U9041 ( .A(b[2724]), .B(n7668), .Z(c[2724]) );
  XNOR U9042 ( .A(a[2724]), .B(n7669), .Z(n7668) );
  IV U9043 ( .A(n7666), .Z(n7669) );
  XOR U9044 ( .A(n7670), .B(n7671), .Z(n7666) );
  ANDN U9045 ( .B(n7672), .A(n7673), .Z(n7670) );
  XNOR U9046 ( .A(b[2723]), .B(n7671), .Z(n7672) );
  XNOR U9047 ( .A(b[2723]), .B(n7673), .Z(c[2723]) );
  XNOR U9048 ( .A(a[2723]), .B(n7674), .Z(n7673) );
  IV U9049 ( .A(n7671), .Z(n7674) );
  XOR U9050 ( .A(n7675), .B(n7676), .Z(n7671) );
  ANDN U9051 ( .B(n7677), .A(n7678), .Z(n7675) );
  XNOR U9052 ( .A(b[2722]), .B(n7676), .Z(n7677) );
  XNOR U9053 ( .A(b[2722]), .B(n7678), .Z(c[2722]) );
  XNOR U9054 ( .A(a[2722]), .B(n7679), .Z(n7678) );
  IV U9055 ( .A(n7676), .Z(n7679) );
  XOR U9056 ( .A(n7680), .B(n7681), .Z(n7676) );
  ANDN U9057 ( .B(n7682), .A(n7683), .Z(n7680) );
  XNOR U9058 ( .A(b[2721]), .B(n7681), .Z(n7682) );
  XNOR U9059 ( .A(b[2721]), .B(n7683), .Z(c[2721]) );
  XNOR U9060 ( .A(a[2721]), .B(n7684), .Z(n7683) );
  IV U9061 ( .A(n7681), .Z(n7684) );
  XOR U9062 ( .A(n7685), .B(n7686), .Z(n7681) );
  ANDN U9063 ( .B(n7687), .A(n7688), .Z(n7685) );
  XNOR U9064 ( .A(b[2720]), .B(n7686), .Z(n7687) );
  XNOR U9065 ( .A(b[2720]), .B(n7688), .Z(c[2720]) );
  XNOR U9066 ( .A(a[2720]), .B(n7689), .Z(n7688) );
  IV U9067 ( .A(n7686), .Z(n7689) );
  XOR U9068 ( .A(n7690), .B(n7691), .Z(n7686) );
  ANDN U9069 ( .B(n7692), .A(n7693), .Z(n7690) );
  XNOR U9070 ( .A(b[2719]), .B(n7691), .Z(n7692) );
  XNOR U9071 ( .A(b[271]), .B(n7694), .Z(c[271]) );
  XNOR U9072 ( .A(b[2719]), .B(n7693), .Z(c[2719]) );
  XNOR U9073 ( .A(a[2719]), .B(n7695), .Z(n7693) );
  IV U9074 ( .A(n7691), .Z(n7695) );
  XOR U9075 ( .A(n7696), .B(n7697), .Z(n7691) );
  ANDN U9076 ( .B(n7698), .A(n7699), .Z(n7696) );
  XNOR U9077 ( .A(b[2718]), .B(n7697), .Z(n7698) );
  XNOR U9078 ( .A(b[2718]), .B(n7699), .Z(c[2718]) );
  XNOR U9079 ( .A(a[2718]), .B(n7700), .Z(n7699) );
  IV U9080 ( .A(n7697), .Z(n7700) );
  XOR U9081 ( .A(n7701), .B(n7702), .Z(n7697) );
  ANDN U9082 ( .B(n7703), .A(n7704), .Z(n7701) );
  XNOR U9083 ( .A(b[2717]), .B(n7702), .Z(n7703) );
  XNOR U9084 ( .A(b[2717]), .B(n7704), .Z(c[2717]) );
  XNOR U9085 ( .A(a[2717]), .B(n7705), .Z(n7704) );
  IV U9086 ( .A(n7702), .Z(n7705) );
  XOR U9087 ( .A(n7706), .B(n7707), .Z(n7702) );
  ANDN U9088 ( .B(n7708), .A(n7709), .Z(n7706) );
  XNOR U9089 ( .A(b[2716]), .B(n7707), .Z(n7708) );
  XNOR U9090 ( .A(b[2716]), .B(n7709), .Z(c[2716]) );
  XNOR U9091 ( .A(a[2716]), .B(n7710), .Z(n7709) );
  IV U9092 ( .A(n7707), .Z(n7710) );
  XOR U9093 ( .A(n7711), .B(n7712), .Z(n7707) );
  ANDN U9094 ( .B(n7713), .A(n7714), .Z(n7711) );
  XNOR U9095 ( .A(b[2715]), .B(n7712), .Z(n7713) );
  XNOR U9096 ( .A(b[2715]), .B(n7714), .Z(c[2715]) );
  XNOR U9097 ( .A(a[2715]), .B(n7715), .Z(n7714) );
  IV U9098 ( .A(n7712), .Z(n7715) );
  XOR U9099 ( .A(n7716), .B(n7717), .Z(n7712) );
  ANDN U9100 ( .B(n7718), .A(n7719), .Z(n7716) );
  XNOR U9101 ( .A(b[2714]), .B(n7717), .Z(n7718) );
  XNOR U9102 ( .A(b[2714]), .B(n7719), .Z(c[2714]) );
  XNOR U9103 ( .A(a[2714]), .B(n7720), .Z(n7719) );
  IV U9104 ( .A(n7717), .Z(n7720) );
  XOR U9105 ( .A(n7721), .B(n7722), .Z(n7717) );
  ANDN U9106 ( .B(n7723), .A(n7724), .Z(n7721) );
  XNOR U9107 ( .A(b[2713]), .B(n7722), .Z(n7723) );
  XNOR U9108 ( .A(b[2713]), .B(n7724), .Z(c[2713]) );
  XNOR U9109 ( .A(a[2713]), .B(n7725), .Z(n7724) );
  IV U9110 ( .A(n7722), .Z(n7725) );
  XOR U9111 ( .A(n7726), .B(n7727), .Z(n7722) );
  ANDN U9112 ( .B(n7728), .A(n7729), .Z(n7726) );
  XNOR U9113 ( .A(b[2712]), .B(n7727), .Z(n7728) );
  XNOR U9114 ( .A(b[2712]), .B(n7729), .Z(c[2712]) );
  XNOR U9115 ( .A(a[2712]), .B(n7730), .Z(n7729) );
  IV U9116 ( .A(n7727), .Z(n7730) );
  XOR U9117 ( .A(n7731), .B(n7732), .Z(n7727) );
  ANDN U9118 ( .B(n7733), .A(n7734), .Z(n7731) );
  XNOR U9119 ( .A(b[2711]), .B(n7732), .Z(n7733) );
  XNOR U9120 ( .A(b[2711]), .B(n7734), .Z(c[2711]) );
  XNOR U9121 ( .A(a[2711]), .B(n7735), .Z(n7734) );
  IV U9122 ( .A(n7732), .Z(n7735) );
  XOR U9123 ( .A(n7736), .B(n7737), .Z(n7732) );
  ANDN U9124 ( .B(n7738), .A(n7739), .Z(n7736) );
  XNOR U9125 ( .A(b[2710]), .B(n7737), .Z(n7738) );
  XNOR U9126 ( .A(b[2710]), .B(n7739), .Z(c[2710]) );
  XNOR U9127 ( .A(a[2710]), .B(n7740), .Z(n7739) );
  IV U9128 ( .A(n7737), .Z(n7740) );
  XOR U9129 ( .A(n7741), .B(n7742), .Z(n7737) );
  ANDN U9130 ( .B(n7743), .A(n7744), .Z(n7741) );
  XNOR U9131 ( .A(b[2709]), .B(n7742), .Z(n7743) );
  XNOR U9132 ( .A(b[270]), .B(n7745), .Z(c[270]) );
  XNOR U9133 ( .A(b[2709]), .B(n7744), .Z(c[2709]) );
  XNOR U9134 ( .A(a[2709]), .B(n7746), .Z(n7744) );
  IV U9135 ( .A(n7742), .Z(n7746) );
  XOR U9136 ( .A(n7747), .B(n7748), .Z(n7742) );
  ANDN U9137 ( .B(n7749), .A(n7750), .Z(n7747) );
  XNOR U9138 ( .A(b[2708]), .B(n7748), .Z(n7749) );
  XNOR U9139 ( .A(b[2708]), .B(n7750), .Z(c[2708]) );
  XNOR U9140 ( .A(a[2708]), .B(n7751), .Z(n7750) );
  IV U9141 ( .A(n7748), .Z(n7751) );
  XOR U9142 ( .A(n7752), .B(n7753), .Z(n7748) );
  ANDN U9143 ( .B(n7754), .A(n7755), .Z(n7752) );
  XNOR U9144 ( .A(b[2707]), .B(n7753), .Z(n7754) );
  XNOR U9145 ( .A(b[2707]), .B(n7755), .Z(c[2707]) );
  XNOR U9146 ( .A(a[2707]), .B(n7756), .Z(n7755) );
  IV U9147 ( .A(n7753), .Z(n7756) );
  XOR U9148 ( .A(n7757), .B(n7758), .Z(n7753) );
  ANDN U9149 ( .B(n7759), .A(n7760), .Z(n7757) );
  XNOR U9150 ( .A(b[2706]), .B(n7758), .Z(n7759) );
  XNOR U9151 ( .A(b[2706]), .B(n7760), .Z(c[2706]) );
  XNOR U9152 ( .A(a[2706]), .B(n7761), .Z(n7760) );
  IV U9153 ( .A(n7758), .Z(n7761) );
  XOR U9154 ( .A(n7762), .B(n7763), .Z(n7758) );
  ANDN U9155 ( .B(n7764), .A(n7765), .Z(n7762) );
  XNOR U9156 ( .A(b[2705]), .B(n7763), .Z(n7764) );
  XNOR U9157 ( .A(b[2705]), .B(n7765), .Z(c[2705]) );
  XNOR U9158 ( .A(a[2705]), .B(n7766), .Z(n7765) );
  IV U9159 ( .A(n7763), .Z(n7766) );
  XOR U9160 ( .A(n7767), .B(n7768), .Z(n7763) );
  ANDN U9161 ( .B(n7769), .A(n7770), .Z(n7767) );
  XNOR U9162 ( .A(b[2704]), .B(n7768), .Z(n7769) );
  XNOR U9163 ( .A(b[2704]), .B(n7770), .Z(c[2704]) );
  XNOR U9164 ( .A(a[2704]), .B(n7771), .Z(n7770) );
  IV U9165 ( .A(n7768), .Z(n7771) );
  XOR U9166 ( .A(n7772), .B(n7773), .Z(n7768) );
  ANDN U9167 ( .B(n7774), .A(n7775), .Z(n7772) );
  XNOR U9168 ( .A(b[2703]), .B(n7773), .Z(n7774) );
  XNOR U9169 ( .A(b[2703]), .B(n7775), .Z(c[2703]) );
  XNOR U9170 ( .A(a[2703]), .B(n7776), .Z(n7775) );
  IV U9171 ( .A(n7773), .Z(n7776) );
  XOR U9172 ( .A(n7777), .B(n7778), .Z(n7773) );
  ANDN U9173 ( .B(n7779), .A(n7780), .Z(n7777) );
  XNOR U9174 ( .A(b[2702]), .B(n7778), .Z(n7779) );
  XNOR U9175 ( .A(b[2702]), .B(n7780), .Z(c[2702]) );
  XNOR U9176 ( .A(a[2702]), .B(n7781), .Z(n7780) );
  IV U9177 ( .A(n7778), .Z(n7781) );
  XOR U9178 ( .A(n7782), .B(n7783), .Z(n7778) );
  ANDN U9179 ( .B(n7784), .A(n7785), .Z(n7782) );
  XNOR U9180 ( .A(b[2701]), .B(n7783), .Z(n7784) );
  XNOR U9181 ( .A(b[2701]), .B(n7785), .Z(c[2701]) );
  XNOR U9182 ( .A(a[2701]), .B(n7786), .Z(n7785) );
  IV U9183 ( .A(n7783), .Z(n7786) );
  XOR U9184 ( .A(n7787), .B(n7788), .Z(n7783) );
  ANDN U9185 ( .B(n7789), .A(n7790), .Z(n7787) );
  XNOR U9186 ( .A(b[2700]), .B(n7788), .Z(n7789) );
  XNOR U9187 ( .A(b[2700]), .B(n7790), .Z(c[2700]) );
  XNOR U9188 ( .A(a[2700]), .B(n7791), .Z(n7790) );
  IV U9189 ( .A(n7788), .Z(n7791) );
  XOR U9190 ( .A(n7792), .B(n7793), .Z(n7788) );
  ANDN U9191 ( .B(n7794), .A(n7795), .Z(n7792) );
  XNOR U9192 ( .A(b[2699]), .B(n7793), .Z(n7794) );
  XNOR U9193 ( .A(b[26]), .B(n7796), .Z(c[26]) );
  XNOR U9194 ( .A(b[269]), .B(n7797), .Z(c[269]) );
  XNOR U9195 ( .A(b[2699]), .B(n7795), .Z(c[2699]) );
  XNOR U9196 ( .A(a[2699]), .B(n7798), .Z(n7795) );
  IV U9197 ( .A(n7793), .Z(n7798) );
  XOR U9198 ( .A(n7799), .B(n7800), .Z(n7793) );
  ANDN U9199 ( .B(n7801), .A(n7802), .Z(n7799) );
  XNOR U9200 ( .A(b[2698]), .B(n7800), .Z(n7801) );
  XNOR U9201 ( .A(b[2698]), .B(n7802), .Z(c[2698]) );
  XNOR U9202 ( .A(a[2698]), .B(n7803), .Z(n7802) );
  IV U9203 ( .A(n7800), .Z(n7803) );
  XOR U9204 ( .A(n7804), .B(n7805), .Z(n7800) );
  ANDN U9205 ( .B(n7806), .A(n7807), .Z(n7804) );
  XNOR U9206 ( .A(b[2697]), .B(n7805), .Z(n7806) );
  XNOR U9207 ( .A(b[2697]), .B(n7807), .Z(c[2697]) );
  XNOR U9208 ( .A(a[2697]), .B(n7808), .Z(n7807) );
  IV U9209 ( .A(n7805), .Z(n7808) );
  XOR U9210 ( .A(n7809), .B(n7810), .Z(n7805) );
  ANDN U9211 ( .B(n7811), .A(n7812), .Z(n7809) );
  XNOR U9212 ( .A(b[2696]), .B(n7810), .Z(n7811) );
  XNOR U9213 ( .A(b[2696]), .B(n7812), .Z(c[2696]) );
  XNOR U9214 ( .A(a[2696]), .B(n7813), .Z(n7812) );
  IV U9215 ( .A(n7810), .Z(n7813) );
  XOR U9216 ( .A(n7814), .B(n7815), .Z(n7810) );
  ANDN U9217 ( .B(n7816), .A(n7817), .Z(n7814) );
  XNOR U9218 ( .A(b[2695]), .B(n7815), .Z(n7816) );
  XNOR U9219 ( .A(b[2695]), .B(n7817), .Z(c[2695]) );
  XNOR U9220 ( .A(a[2695]), .B(n7818), .Z(n7817) );
  IV U9221 ( .A(n7815), .Z(n7818) );
  XOR U9222 ( .A(n7819), .B(n7820), .Z(n7815) );
  ANDN U9223 ( .B(n7821), .A(n7822), .Z(n7819) );
  XNOR U9224 ( .A(b[2694]), .B(n7820), .Z(n7821) );
  XNOR U9225 ( .A(b[2694]), .B(n7822), .Z(c[2694]) );
  XNOR U9226 ( .A(a[2694]), .B(n7823), .Z(n7822) );
  IV U9227 ( .A(n7820), .Z(n7823) );
  XOR U9228 ( .A(n7824), .B(n7825), .Z(n7820) );
  ANDN U9229 ( .B(n7826), .A(n7827), .Z(n7824) );
  XNOR U9230 ( .A(b[2693]), .B(n7825), .Z(n7826) );
  XNOR U9231 ( .A(b[2693]), .B(n7827), .Z(c[2693]) );
  XNOR U9232 ( .A(a[2693]), .B(n7828), .Z(n7827) );
  IV U9233 ( .A(n7825), .Z(n7828) );
  XOR U9234 ( .A(n7829), .B(n7830), .Z(n7825) );
  ANDN U9235 ( .B(n7831), .A(n7832), .Z(n7829) );
  XNOR U9236 ( .A(b[2692]), .B(n7830), .Z(n7831) );
  XNOR U9237 ( .A(b[2692]), .B(n7832), .Z(c[2692]) );
  XNOR U9238 ( .A(a[2692]), .B(n7833), .Z(n7832) );
  IV U9239 ( .A(n7830), .Z(n7833) );
  XOR U9240 ( .A(n7834), .B(n7835), .Z(n7830) );
  ANDN U9241 ( .B(n7836), .A(n7837), .Z(n7834) );
  XNOR U9242 ( .A(b[2691]), .B(n7835), .Z(n7836) );
  XNOR U9243 ( .A(b[2691]), .B(n7837), .Z(c[2691]) );
  XNOR U9244 ( .A(a[2691]), .B(n7838), .Z(n7837) );
  IV U9245 ( .A(n7835), .Z(n7838) );
  XOR U9246 ( .A(n7839), .B(n7840), .Z(n7835) );
  ANDN U9247 ( .B(n7841), .A(n7842), .Z(n7839) );
  XNOR U9248 ( .A(b[2690]), .B(n7840), .Z(n7841) );
  XNOR U9249 ( .A(b[2690]), .B(n7842), .Z(c[2690]) );
  XNOR U9250 ( .A(a[2690]), .B(n7843), .Z(n7842) );
  IV U9251 ( .A(n7840), .Z(n7843) );
  XOR U9252 ( .A(n7844), .B(n7845), .Z(n7840) );
  ANDN U9253 ( .B(n7846), .A(n7847), .Z(n7844) );
  XNOR U9254 ( .A(b[2689]), .B(n7845), .Z(n7846) );
  XNOR U9255 ( .A(b[268]), .B(n7848), .Z(c[268]) );
  XNOR U9256 ( .A(b[2689]), .B(n7847), .Z(c[2689]) );
  XNOR U9257 ( .A(a[2689]), .B(n7849), .Z(n7847) );
  IV U9258 ( .A(n7845), .Z(n7849) );
  XOR U9259 ( .A(n7850), .B(n7851), .Z(n7845) );
  ANDN U9260 ( .B(n7852), .A(n7853), .Z(n7850) );
  XNOR U9261 ( .A(b[2688]), .B(n7851), .Z(n7852) );
  XNOR U9262 ( .A(b[2688]), .B(n7853), .Z(c[2688]) );
  XNOR U9263 ( .A(a[2688]), .B(n7854), .Z(n7853) );
  IV U9264 ( .A(n7851), .Z(n7854) );
  XOR U9265 ( .A(n7855), .B(n7856), .Z(n7851) );
  ANDN U9266 ( .B(n7857), .A(n7858), .Z(n7855) );
  XNOR U9267 ( .A(b[2687]), .B(n7856), .Z(n7857) );
  XNOR U9268 ( .A(b[2687]), .B(n7858), .Z(c[2687]) );
  XNOR U9269 ( .A(a[2687]), .B(n7859), .Z(n7858) );
  IV U9270 ( .A(n7856), .Z(n7859) );
  XOR U9271 ( .A(n7860), .B(n7861), .Z(n7856) );
  ANDN U9272 ( .B(n7862), .A(n7863), .Z(n7860) );
  XNOR U9273 ( .A(b[2686]), .B(n7861), .Z(n7862) );
  XNOR U9274 ( .A(b[2686]), .B(n7863), .Z(c[2686]) );
  XNOR U9275 ( .A(a[2686]), .B(n7864), .Z(n7863) );
  IV U9276 ( .A(n7861), .Z(n7864) );
  XOR U9277 ( .A(n7865), .B(n7866), .Z(n7861) );
  ANDN U9278 ( .B(n7867), .A(n7868), .Z(n7865) );
  XNOR U9279 ( .A(b[2685]), .B(n7866), .Z(n7867) );
  XNOR U9280 ( .A(b[2685]), .B(n7868), .Z(c[2685]) );
  XNOR U9281 ( .A(a[2685]), .B(n7869), .Z(n7868) );
  IV U9282 ( .A(n7866), .Z(n7869) );
  XOR U9283 ( .A(n7870), .B(n7871), .Z(n7866) );
  ANDN U9284 ( .B(n7872), .A(n7873), .Z(n7870) );
  XNOR U9285 ( .A(b[2684]), .B(n7871), .Z(n7872) );
  XNOR U9286 ( .A(b[2684]), .B(n7873), .Z(c[2684]) );
  XNOR U9287 ( .A(a[2684]), .B(n7874), .Z(n7873) );
  IV U9288 ( .A(n7871), .Z(n7874) );
  XOR U9289 ( .A(n7875), .B(n7876), .Z(n7871) );
  ANDN U9290 ( .B(n7877), .A(n7878), .Z(n7875) );
  XNOR U9291 ( .A(b[2683]), .B(n7876), .Z(n7877) );
  XNOR U9292 ( .A(b[2683]), .B(n7878), .Z(c[2683]) );
  XNOR U9293 ( .A(a[2683]), .B(n7879), .Z(n7878) );
  IV U9294 ( .A(n7876), .Z(n7879) );
  XOR U9295 ( .A(n7880), .B(n7881), .Z(n7876) );
  ANDN U9296 ( .B(n7882), .A(n7883), .Z(n7880) );
  XNOR U9297 ( .A(b[2682]), .B(n7881), .Z(n7882) );
  XNOR U9298 ( .A(b[2682]), .B(n7883), .Z(c[2682]) );
  XNOR U9299 ( .A(a[2682]), .B(n7884), .Z(n7883) );
  IV U9300 ( .A(n7881), .Z(n7884) );
  XOR U9301 ( .A(n7885), .B(n7886), .Z(n7881) );
  ANDN U9302 ( .B(n7887), .A(n7888), .Z(n7885) );
  XNOR U9303 ( .A(b[2681]), .B(n7886), .Z(n7887) );
  XNOR U9304 ( .A(b[2681]), .B(n7888), .Z(c[2681]) );
  XNOR U9305 ( .A(a[2681]), .B(n7889), .Z(n7888) );
  IV U9306 ( .A(n7886), .Z(n7889) );
  XOR U9307 ( .A(n7890), .B(n7891), .Z(n7886) );
  ANDN U9308 ( .B(n7892), .A(n7893), .Z(n7890) );
  XNOR U9309 ( .A(b[2680]), .B(n7891), .Z(n7892) );
  XNOR U9310 ( .A(b[2680]), .B(n7893), .Z(c[2680]) );
  XNOR U9311 ( .A(a[2680]), .B(n7894), .Z(n7893) );
  IV U9312 ( .A(n7891), .Z(n7894) );
  XOR U9313 ( .A(n7895), .B(n7896), .Z(n7891) );
  ANDN U9314 ( .B(n7897), .A(n7898), .Z(n7895) );
  XNOR U9315 ( .A(b[2679]), .B(n7896), .Z(n7897) );
  XNOR U9316 ( .A(b[267]), .B(n7899), .Z(c[267]) );
  XNOR U9317 ( .A(b[2679]), .B(n7898), .Z(c[2679]) );
  XNOR U9318 ( .A(a[2679]), .B(n7900), .Z(n7898) );
  IV U9319 ( .A(n7896), .Z(n7900) );
  XOR U9320 ( .A(n7901), .B(n7902), .Z(n7896) );
  ANDN U9321 ( .B(n7903), .A(n7904), .Z(n7901) );
  XNOR U9322 ( .A(b[2678]), .B(n7902), .Z(n7903) );
  XNOR U9323 ( .A(b[2678]), .B(n7904), .Z(c[2678]) );
  XNOR U9324 ( .A(a[2678]), .B(n7905), .Z(n7904) );
  IV U9325 ( .A(n7902), .Z(n7905) );
  XOR U9326 ( .A(n7906), .B(n7907), .Z(n7902) );
  ANDN U9327 ( .B(n7908), .A(n7909), .Z(n7906) );
  XNOR U9328 ( .A(b[2677]), .B(n7907), .Z(n7908) );
  XNOR U9329 ( .A(b[2677]), .B(n7909), .Z(c[2677]) );
  XNOR U9330 ( .A(a[2677]), .B(n7910), .Z(n7909) );
  IV U9331 ( .A(n7907), .Z(n7910) );
  XOR U9332 ( .A(n7911), .B(n7912), .Z(n7907) );
  ANDN U9333 ( .B(n7913), .A(n7914), .Z(n7911) );
  XNOR U9334 ( .A(b[2676]), .B(n7912), .Z(n7913) );
  XNOR U9335 ( .A(b[2676]), .B(n7914), .Z(c[2676]) );
  XNOR U9336 ( .A(a[2676]), .B(n7915), .Z(n7914) );
  IV U9337 ( .A(n7912), .Z(n7915) );
  XOR U9338 ( .A(n7916), .B(n7917), .Z(n7912) );
  ANDN U9339 ( .B(n7918), .A(n7919), .Z(n7916) );
  XNOR U9340 ( .A(b[2675]), .B(n7917), .Z(n7918) );
  XNOR U9341 ( .A(b[2675]), .B(n7919), .Z(c[2675]) );
  XNOR U9342 ( .A(a[2675]), .B(n7920), .Z(n7919) );
  IV U9343 ( .A(n7917), .Z(n7920) );
  XOR U9344 ( .A(n7921), .B(n7922), .Z(n7917) );
  ANDN U9345 ( .B(n7923), .A(n7924), .Z(n7921) );
  XNOR U9346 ( .A(b[2674]), .B(n7922), .Z(n7923) );
  XNOR U9347 ( .A(b[2674]), .B(n7924), .Z(c[2674]) );
  XNOR U9348 ( .A(a[2674]), .B(n7925), .Z(n7924) );
  IV U9349 ( .A(n7922), .Z(n7925) );
  XOR U9350 ( .A(n7926), .B(n7927), .Z(n7922) );
  ANDN U9351 ( .B(n7928), .A(n7929), .Z(n7926) );
  XNOR U9352 ( .A(b[2673]), .B(n7927), .Z(n7928) );
  XNOR U9353 ( .A(b[2673]), .B(n7929), .Z(c[2673]) );
  XNOR U9354 ( .A(a[2673]), .B(n7930), .Z(n7929) );
  IV U9355 ( .A(n7927), .Z(n7930) );
  XOR U9356 ( .A(n7931), .B(n7932), .Z(n7927) );
  ANDN U9357 ( .B(n7933), .A(n7934), .Z(n7931) );
  XNOR U9358 ( .A(b[2672]), .B(n7932), .Z(n7933) );
  XNOR U9359 ( .A(b[2672]), .B(n7934), .Z(c[2672]) );
  XNOR U9360 ( .A(a[2672]), .B(n7935), .Z(n7934) );
  IV U9361 ( .A(n7932), .Z(n7935) );
  XOR U9362 ( .A(n7936), .B(n7937), .Z(n7932) );
  ANDN U9363 ( .B(n7938), .A(n7939), .Z(n7936) );
  XNOR U9364 ( .A(b[2671]), .B(n7937), .Z(n7938) );
  XNOR U9365 ( .A(b[2671]), .B(n7939), .Z(c[2671]) );
  XNOR U9366 ( .A(a[2671]), .B(n7940), .Z(n7939) );
  IV U9367 ( .A(n7937), .Z(n7940) );
  XOR U9368 ( .A(n7941), .B(n7942), .Z(n7937) );
  ANDN U9369 ( .B(n7943), .A(n7944), .Z(n7941) );
  XNOR U9370 ( .A(b[2670]), .B(n7942), .Z(n7943) );
  XNOR U9371 ( .A(b[2670]), .B(n7944), .Z(c[2670]) );
  XNOR U9372 ( .A(a[2670]), .B(n7945), .Z(n7944) );
  IV U9373 ( .A(n7942), .Z(n7945) );
  XOR U9374 ( .A(n7946), .B(n7947), .Z(n7942) );
  ANDN U9375 ( .B(n7948), .A(n7949), .Z(n7946) );
  XNOR U9376 ( .A(b[2669]), .B(n7947), .Z(n7948) );
  XNOR U9377 ( .A(b[266]), .B(n7950), .Z(c[266]) );
  XNOR U9378 ( .A(b[2669]), .B(n7949), .Z(c[2669]) );
  XNOR U9379 ( .A(a[2669]), .B(n7951), .Z(n7949) );
  IV U9380 ( .A(n7947), .Z(n7951) );
  XOR U9381 ( .A(n7952), .B(n7953), .Z(n7947) );
  ANDN U9382 ( .B(n7954), .A(n7955), .Z(n7952) );
  XNOR U9383 ( .A(b[2668]), .B(n7953), .Z(n7954) );
  XNOR U9384 ( .A(b[2668]), .B(n7955), .Z(c[2668]) );
  XNOR U9385 ( .A(a[2668]), .B(n7956), .Z(n7955) );
  IV U9386 ( .A(n7953), .Z(n7956) );
  XOR U9387 ( .A(n7957), .B(n7958), .Z(n7953) );
  ANDN U9388 ( .B(n7959), .A(n7960), .Z(n7957) );
  XNOR U9389 ( .A(b[2667]), .B(n7958), .Z(n7959) );
  XNOR U9390 ( .A(b[2667]), .B(n7960), .Z(c[2667]) );
  XNOR U9391 ( .A(a[2667]), .B(n7961), .Z(n7960) );
  IV U9392 ( .A(n7958), .Z(n7961) );
  XOR U9393 ( .A(n7962), .B(n7963), .Z(n7958) );
  ANDN U9394 ( .B(n7964), .A(n7965), .Z(n7962) );
  XNOR U9395 ( .A(b[2666]), .B(n7963), .Z(n7964) );
  XNOR U9396 ( .A(b[2666]), .B(n7965), .Z(c[2666]) );
  XNOR U9397 ( .A(a[2666]), .B(n7966), .Z(n7965) );
  IV U9398 ( .A(n7963), .Z(n7966) );
  XOR U9399 ( .A(n7967), .B(n7968), .Z(n7963) );
  ANDN U9400 ( .B(n7969), .A(n7970), .Z(n7967) );
  XNOR U9401 ( .A(b[2665]), .B(n7968), .Z(n7969) );
  XNOR U9402 ( .A(b[2665]), .B(n7970), .Z(c[2665]) );
  XNOR U9403 ( .A(a[2665]), .B(n7971), .Z(n7970) );
  IV U9404 ( .A(n7968), .Z(n7971) );
  XOR U9405 ( .A(n7972), .B(n7973), .Z(n7968) );
  ANDN U9406 ( .B(n7974), .A(n7975), .Z(n7972) );
  XNOR U9407 ( .A(b[2664]), .B(n7973), .Z(n7974) );
  XNOR U9408 ( .A(b[2664]), .B(n7975), .Z(c[2664]) );
  XNOR U9409 ( .A(a[2664]), .B(n7976), .Z(n7975) );
  IV U9410 ( .A(n7973), .Z(n7976) );
  XOR U9411 ( .A(n7977), .B(n7978), .Z(n7973) );
  ANDN U9412 ( .B(n7979), .A(n7980), .Z(n7977) );
  XNOR U9413 ( .A(b[2663]), .B(n7978), .Z(n7979) );
  XNOR U9414 ( .A(b[2663]), .B(n7980), .Z(c[2663]) );
  XNOR U9415 ( .A(a[2663]), .B(n7981), .Z(n7980) );
  IV U9416 ( .A(n7978), .Z(n7981) );
  XOR U9417 ( .A(n7982), .B(n7983), .Z(n7978) );
  ANDN U9418 ( .B(n7984), .A(n7985), .Z(n7982) );
  XNOR U9419 ( .A(b[2662]), .B(n7983), .Z(n7984) );
  XNOR U9420 ( .A(b[2662]), .B(n7985), .Z(c[2662]) );
  XNOR U9421 ( .A(a[2662]), .B(n7986), .Z(n7985) );
  IV U9422 ( .A(n7983), .Z(n7986) );
  XOR U9423 ( .A(n7987), .B(n7988), .Z(n7983) );
  ANDN U9424 ( .B(n7989), .A(n7990), .Z(n7987) );
  XNOR U9425 ( .A(b[2661]), .B(n7988), .Z(n7989) );
  XNOR U9426 ( .A(b[2661]), .B(n7990), .Z(c[2661]) );
  XNOR U9427 ( .A(a[2661]), .B(n7991), .Z(n7990) );
  IV U9428 ( .A(n7988), .Z(n7991) );
  XOR U9429 ( .A(n7992), .B(n7993), .Z(n7988) );
  ANDN U9430 ( .B(n7994), .A(n7995), .Z(n7992) );
  XNOR U9431 ( .A(b[2660]), .B(n7993), .Z(n7994) );
  XNOR U9432 ( .A(b[2660]), .B(n7995), .Z(c[2660]) );
  XNOR U9433 ( .A(a[2660]), .B(n7996), .Z(n7995) );
  IV U9434 ( .A(n7993), .Z(n7996) );
  XOR U9435 ( .A(n7997), .B(n7998), .Z(n7993) );
  ANDN U9436 ( .B(n7999), .A(n8000), .Z(n7997) );
  XNOR U9437 ( .A(b[2659]), .B(n7998), .Z(n7999) );
  XNOR U9438 ( .A(b[265]), .B(n8001), .Z(c[265]) );
  XNOR U9439 ( .A(b[2659]), .B(n8000), .Z(c[2659]) );
  XNOR U9440 ( .A(a[2659]), .B(n8002), .Z(n8000) );
  IV U9441 ( .A(n7998), .Z(n8002) );
  XOR U9442 ( .A(n8003), .B(n8004), .Z(n7998) );
  ANDN U9443 ( .B(n8005), .A(n8006), .Z(n8003) );
  XNOR U9444 ( .A(b[2658]), .B(n8004), .Z(n8005) );
  XNOR U9445 ( .A(b[2658]), .B(n8006), .Z(c[2658]) );
  XNOR U9446 ( .A(a[2658]), .B(n8007), .Z(n8006) );
  IV U9447 ( .A(n8004), .Z(n8007) );
  XOR U9448 ( .A(n8008), .B(n8009), .Z(n8004) );
  ANDN U9449 ( .B(n8010), .A(n8011), .Z(n8008) );
  XNOR U9450 ( .A(b[2657]), .B(n8009), .Z(n8010) );
  XNOR U9451 ( .A(b[2657]), .B(n8011), .Z(c[2657]) );
  XNOR U9452 ( .A(a[2657]), .B(n8012), .Z(n8011) );
  IV U9453 ( .A(n8009), .Z(n8012) );
  XOR U9454 ( .A(n8013), .B(n8014), .Z(n8009) );
  ANDN U9455 ( .B(n8015), .A(n8016), .Z(n8013) );
  XNOR U9456 ( .A(b[2656]), .B(n8014), .Z(n8015) );
  XNOR U9457 ( .A(b[2656]), .B(n8016), .Z(c[2656]) );
  XNOR U9458 ( .A(a[2656]), .B(n8017), .Z(n8016) );
  IV U9459 ( .A(n8014), .Z(n8017) );
  XOR U9460 ( .A(n8018), .B(n8019), .Z(n8014) );
  ANDN U9461 ( .B(n8020), .A(n8021), .Z(n8018) );
  XNOR U9462 ( .A(b[2655]), .B(n8019), .Z(n8020) );
  XNOR U9463 ( .A(b[2655]), .B(n8021), .Z(c[2655]) );
  XNOR U9464 ( .A(a[2655]), .B(n8022), .Z(n8021) );
  IV U9465 ( .A(n8019), .Z(n8022) );
  XOR U9466 ( .A(n8023), .B(n8024), .Z(n8019) );
  ANDN U9467 ( .B(n8025), .A(n8026), .Z(n8023) );
  XNOR U9468 ( .A(b[2654]), .B(n8024), .Z(n8025) );
  XNOR U9469 ( .A(b[2654]), .B(n8026), .Z(c[2654]) );
  XNOR U9470 ( .A(a[2654]), .B(n8027), .Z(n8026) );
  IV U9471 ( .A(n8024), .Z(n8027) );
  XOR U9472 ( .A(n8028), .B(n8029), .Z(n8024) );
  ANDN U9473 ( .B(n8030), .A(n8031), .Z(n8028) );
  XNOR U9474 ( .A(b[2653]), .B(n8029), .Z(n8030) );
  XNOR U9475 ( .A(b[2653]), .B(n8031), .Z(c[2653]) );
  XNOR U9476 ( .A(a[2653]), .B(n8032), .Z(n8031) );
  IV U9477 ( .A(n8029), .Z(n8032) );
  XOR U9478 ( .A(n8033), .B(n8034), .Z(n8029) );
  ANDN U9479 ( .B(n8035), .A(n8036), .Z(n8033) );
  XNOR U9480 ( .A(b[2652]), .B(n8034), .Z(n8035) );
  XNOR U9481 ( .A(b[2652]), .B(n8036), .Z(c[2652]) );
  XNOR U9482 ( .A(a[2652]), .B(n8037), .Z(n8036) );
  IV U9483 ( .A(n8034), .Z(n8037) );
  XOR U9484 ( .A(n8038), .B(n8039), .Z(n8034) );
  ANDN U9485 ( .B(n8040), .A(n8041), .Z(n8038) );
  XNOR U9486 ( .A(b[2651]), .B(n8039), .Z(n8040) );
  XNOR U9487 ( .A(b[2651]), .B(n8041), .Z(c[2651]) );
  XNOR U9488 ( .A(a[2651]), .B(n8042), .Z(n8041) );
  IV U9489 ( .A(n8039), .Z(n8042) );
  XOR U9490 ( .A(n8043), .B(n8044), .Z(n8039) );
  ANDN U9491 ( .B(n8045), .A(n8046), .Z(n8043) );
  XNOR U9492 ( .A(b[2650]), .B(n8044), .Z(n8045) );
  XNOR U9493 ( .A(b[2650]), .B(n8046), .Z(c[2650]) );
  XNOR U9494 ( .A(a[2650]), .B(n8047), .Z(n8046) );
  IV U9495 ( .A(n8044), .Z(n8047) );
  XOR U9496 ( .A(n8048), .B(n8049), .Z(n8044) );
  ANDN U9497 ( .B(n8050), .A(n8051), .Z(n8048) );
  XNOR U9498 ( .A(b[2649]), .B(n8049), .Z(n8050) );
  XNOR U9499 ( .A(b[264]), .B(n8052), .Z(c[264]) );
  XNOR U9500 ( .A(b[2649]), .B(n8051), .Z(c[2649]) );
  XNOR U9501 ( .A(a[2649]), .B(n8053), .Z(n8051) );
  IV U9502 ( .A(n8049), .Z(n8053) );
  XOR U9503 ( .A(n8054), .B(n8055), .Z(n8049) );
  ANDN U9504 ( .B(n8056), .A(n8057), .Z(n8054) );
  XNOR U9505 ( .A(b[2648]), .B(n8055), .Z(n8056) );
  XNOR U9506 ( .A(b[2648]), .B(n8057), .Z(c[2648]) );
  XNOR U9507 ( .A(a[2648]), .B(n8058), .Z(n8057) );
  IV U9508 ( .A(n8055), .Z(n8058) );
  XOR U9509 ( .A(n8059), .B(n8060), .Z(n8055) );
  ANDN U9510 ( .B(n8061), .A(n8062), .Z(n8059) );
  XNOR U9511 ( .A(b[2647]), .B(n8060), .Z(n8061) );
  XNOR U9512 ( .A(b[2647]), .B(n8062), .Z(c[2647]) );
  XNOR U9513 ( .A(a[2647]), .B(n8063), .Z(n8062) );
  IV U9514 ( .A(n8060), .Z(n8063) );
  XOR U9515 ( .A(n8064), .B(n8065), .Z(n8060) );
  ANDN U9516 ( .B(n8066), .A(n8067), .Z(n8064) );
  XNOR U9517 ( .A(b[2646]), .B(n8065), .Z(n8066) );
  XNOR U9518 ( .A(b[2646]), .B(n8067), .Z(c[2646]) );
  XNOR U9519 ( .A(a[2646]), .B(n8068), .Z(n8067) );
  IV U9520 ( .A(n8065), .Z(n8068) );
  XOR U9521 ( .A(n8069), .B(n8070), .Z(n8065) );
  ANDN U9522 ( .B(n8071), .A(n8072), .Z(n8069) );
  XNOR U9523 ( .A(b[2645]), .B(n8070), .Z(n8071) );
  XNOR U9524 ( .A(b[2645]), .B(n8072), .Z(c[2645]) );
  XNOR U9525 ( .A(a[2645]), .B(n8073), .Z(n8072) );
  IV U9526 ( .A(n8070), .Z(n8073) );
  XOR U9527 ( .A(n8074), .B(n8075), .Z(n8070) );
  ANDN U9528 ( .B(n8076), .A(n8077), .Z(n8074) );
  XNOR U9529 ( .A(b[2644]), .B(n8075), .Z(n8076) );
  XNOR U9530 ( .A(b[2644]), .B(n8077), .Z(c[2644]) );
  XNOR U9531 ( .A(a[2644]), .B(n8078), .Z(n8077) );
  IV U9532 ( .A(n8075), .Z(n8078) );
  XOR U9533 ( .A(n8079), .B(n8080), .Z(n8075) );
  ANDN U9534 ( .B(n8081), .A(n8082), .Z(n8079) );
  XNOR U9535 ( .A(b[2643]), .B(n8080), .Z(n8081) );
  XNOR U9536 ( .A(b[2643]), .B(n8082), .Z(c[2643]) );
  XNOR U9537 ( .A(a[2643]), .B(n8083), .Z(n8082) );
  IV U9538 ( .A(n8080), .Z(n8083) );
  XOR U9539 ( .A(n8084), .B(n8085), .Z(n8080) );
  ANDN U9540 ( .B(n8086), .A(n8087), .Z(n8084) );
  XNOR U9541 ( .A(b[2642]), .B(n8085), .Z(n8086) );
  XNOR U9542 ( .A(b[2642]), .B(n8087), .Z(c[2642]) );
  XNOR U9543 ( .A(a[2642]), .B(n8088), .Z(n8087) );
  IV U9544 ( .A(n8085), .Z(n8088) );
  XOR U9545 ( .A(n8089), .B(n8090), .Z(n8085) );
  ANDN U9546 ( .B(n8091), .A(n8092), .Z(n8089) );
  XNOR U9547 ( .A(b[2641]), .B(n8090), .Z(n8091) );
  XNOR U9548 ( .A(b[2641]), .B(n8092), .Z(c[2641]) );
  XNOR U9549 ( .A(a[2641]), .B(n8093), .Z(n8092) );
  IV U9550 ( .A(n8090), .Z(n8093) );
  XOR U9551 ( .A(n8094), .B(n8095), .Z(n8090) );
  ANDN U9552 ( .B(n8096), .A(n8097), .Z(n8094) );
  XNOR U9553 ( .A(b[2640]), .B(n8095), .Z(n8096) );
  XNOR U9554 ( .A(b[2640]), .B(n8097), .Z(c[2640]) );
  XNOR U9555 ( .A(a[2640]), .B(n8098), .Z(n8097) );
  IV U9556 ( .A(n8095), .Z(n8098) );
  XOR U9557 ( .A(n8099), .B(n8100), .Z(n8095) );
  ANDN U9558 ( .B(n8101), .A(n8102), .Z(n8099) );
  XNOR U9559 ( .A(b[2639]), .B(n8100), .Z(n8101) );
  XNOR U9560 ( .A(b[263]), .B(n8103), .Z(c[263]) );
  XNOR U9561 ( .A(b[2639]), .B(n8102), .Z(c[2639]) );
  XNOR U9562 ( .A(a[2639]), .B(n8104), .Z(n8102) );
  IV U9563 ( .A(n8100), .Z(n8104) );
  XOR U9564 ( .A(n8105), .B(n8106), .Z(n8100) );
  ANDN U9565 ( .B(n8107), .A(n8108), .Z(n8105) );
  XNOR U9566 ( .A(b[2638]), .B(n8106), .Z(n8107) );
  XNOR U9567 ( .A(b[2638]), .B(n8108), .Z(c[2638]) );
  XNOR U9568 ( .A(a[2638]), .B(n8109), .Z(n8108) );
  IV U9569 ( .A(n8106), .Z(n8109) );
  XOR U9570 ( .A(n8110), .B(n8111), .Z(n8106) );
  ANDN U9571 ( .B(n8112), .A(n8113), .Z(n8110) );
  XNOR U9572 ( .A(b[2637]), .B(n8111), .Z(n8112) );
  XNOR U9573 ( .A(b[2637]), .B(n8113), .Z(c[2637]) );
  XNOR U9574 ( .A(a[2637]), .B(n8114), .Z(n8113) );
  IV U9575 ( .A(n8111), .Z(n8114) );
  XOR U9576 ( .A(n8115), .B(n8116), .Z(n8111) );
  ANDN U9577 ( .B(n8117), .A(n8118), .Z(n8115) );
  XNOR U9578 ( .A(b[2636]), .B(n8116), .Z(n8117) );
  XNOR U9579 ( .A(b[2636]), .B(n8118), .Z(c[2636]) );
  XNOR U9580 ( .A(a[2636]), .B(n8119), .Z(n8118) );
  IV U9581 ( .A(n8116), .Z(n8119) );
  XOR U9582 ( .A(n8120), .B(n8121), .Z(n8116) );
  ANDN U9583 ( .B(n8122), .A(n8123), .Z(n8120) );
  XNOR U9584 ( .A(b[2635]), .B(n8121), .Z(n8122) );
  XNOR U9585 ( .A(b[2635]), .B(n8123), .Z(c[2635]) );
  XNOR U9586 ( .A(a[2635]), .B(n8124), .Z(n8123) );
  IV U9587 ( .A(n8121), .Z(n8124) );
  XOR U9588 ( .A(n8125), .B(n8126), .Z(n8121) );
  ANDN U9589 ( .B(n8127), .A(n8128), .Z(n8125) );
  XNOR U9590 ( .A(b[2634]), .B(n8126), .Z(n8127) );
  XNOR U9591 ( .A(b[2634]), .B(n8128), .Z(c[2634]) );
  XNOR U9592 ( .A(a[2634]), .B(n8129), .Z(n8128) );
  IV U9593 ( .A(n8126), .Z(n8129) );
  XOR U9594 ( .A(n8130), .B(n8131), .Z(n8126) );
  ANDN U9595 ( .B(n8132), .A(n8133), .Z(n8130) );
  XNOR U9596 ( .A(b[2633]), .B(n8131), .Z(n8132) );
  XNOR U9597 ( .A(b[2633]), .B(n8133), .Z(c[2633]) );
  XNOR U9598 ( .A(a[2633]), .B(n8134), .Z(n8133) );
  IV U9599 ( .A(n8131), .Z(n8134) );
  XOR U9600 ( .A(n8135), .B(n8136), .Z(n8131) );
  ANDN U9601 ( .B(n8137), .A(n8138), .Z(n8135) );
  XNOR U9602 ( .A(b[2632]), .B(n8136), .Z(n8137) );
  XNOR U9603 ( .A(b[2632]), .B(n8138), .Z(c[2632]) );
  XNOR U9604 ( .A(a[2632]), .B(n8139), .Z(n8138) );
  IV U9605 ( .A(n8136), .Z(n8139) );
  XOR U9606 ( .A(n8140), .B(n8141), .Z(n8136) );
  ANDN U9607 ( .B(n8142), .A(n8143), .Z(n8140) );
  XNOR U9608 ( .A(b[2631]), .B(n8141), .Z(n8142) );
  XNOR U9609 ( .A(b[2631]), .B(n8143), .Z(c[2631]) );
  XNOR U9610 ( .A(a[2631]), .B(n8144), .Z(n8143) );
  IV U9611 ( .A(n8141), .Z(n8144) );
  XOR U9612 ( .A(n8145), .B(n8146), .Z(n8141) );
  ANDN U9613 ( .B(n8147), .A(n8148), .Z(n8145) );
  XNOR U9614 ( .A(b[2630]), .B(n8146), .Z(n8147) );
  XNOR U9615 ( .A(b[2630]), .B(n8148), .Z(c[2630]) );
  XNOR U9616 ( .A(a[2630]), .B(n8149), .Z(n8148) );
  IV U9617 ( .A(n8146), .Z(n8149) );
  XOR U9618 ( .A(n8150), .B(n8151), .Z(n8146) );
  ANDN U9619 ( .B(n8152), .A(n8153), .Z(n8150) );
  XNOR U9620 ( .A(b[2629]), .B(n8151), .Z(n8152) );
  XNOR U9621 ( .A(b[262]), .B(n8154), .Z(c[262]) );
  XNOR U9622 ( .A(b[2629]), .B(n8153), .Z(c[2629]) );
  XNOR U9623 ( .A(a[2629]), .B(n8155), .Z(n8153) );
  IV U9624 ( .A(n8151), .Z(n8155) );
  XOR U9625 ( .A(n8156), .B(n8157), .Z(n8151) );
  ANDN U9626 ( .B(n8158), .A(n8159), .Z(n8156) );
  XNOR U9627 ( .A(b[2628]), .B(n8157), .Z(n8158) );
  XNOR U9628 ( .A(b[2628]), .B(n8159), .Z(c[2628]) );
  XNOR U9629 ( .A(a[2628]), .B(n8160), .Z(n8159) );
  IV U9630 ( .A(n8157), .Z(n8160) );
  XOR U9631 ( .A(n8161), .B(n8162), .Z(n8157) );
  ANDN U9632 ( .B(n8163), .A(n8164), .Z(n8161) );
  XNOR U9633 ( .A(b[2627]), .B(n8162), .Z(n8163) );
  XNOR U9634 ( .A(b[2627]), .B(n8164), .Z(c[2627]) );
  XNOR U9635 ( .A(a[2627]), .B(n8165), .Z(n8164) );
  IV U9636 ( .A(n8162), .Z(n8165) );
  XOR U9637 ( .A(n8166), .B(n8167), .Z(n8162) );
  ANDN U9638 ( .B(n8168), .A(n8169), .Z(n8166) );
  XNOR U9639 ( .A(b[2626]), .B(n8167), .Z(n8168) );
  XNOR U9640 ( .A(b[2626]), .B(n8169), .Z(c[2626]) );
  XNOR U9641 ( .A(a[2626]), .B(n8170), .Z(n8169) );
  IV U9642 ( .A(n8167), .Z(n8170) );
  XOR U9643 ( .A(n8171), .B(n8172), .Z(n8167) );
  ANDN U9644 ( .B(n8173), .A(n8174), .Z(n8171) );
  XNOR U9645 ( .A(b[2625]), .B(n8172), .Z(n8173) );
  XNOR U9646 ( .A(b[2625]), .B(n8174), .Z(c[2625]) );
  XNOR U9647 ( .A(a[2625]), .B(n8175), .Z(n8174) );
  IV U9648 ( .A(n8172), .Z(n8175) );
  XOR U9649 ( .A(n8176), .B(n8177), .Z(n8172) );
  ANDN U9650 ( .B(n8178), .A(n8179), .Z(n8176) );
  XNOR U9651 ( .A(b[2624]), .B(n8177), .Z(n8178) );
  XNOR U9652 ( .A(b[2624]), .B(n8179), .Z(c[2624]) );
  XNOR U9653 ( .A(a[2624]), .B(n8180), .Z(n8179) );
  IV U9654 ( .A(n8177), .Z(n8180) );
  XOR U9655 ( .A(n8181), .B(n8182), .Z(n8177) );
  ANDN U9656 ( .B(n8183), .A(n8184), .Z(n8181) );
  XNOR U9657 ( .A(b[2623]), .B(n8182), .Z(n8183) );
  XNOR U9658 ( .A(b[2623]), .B(n8184), .Z(c[2623]) );
  XNOR U9659 ( .A(a[2623]), .B(n8185), .Z(n8184) );
  IV U9660 ( .A(n8182), .Z(n8185) );
  XOR U9661 ( .A(n8186), .B(n8187), .Z(n8182) );
  ANDN U9662 ( .B(n8188), .A(n8189), .Z(n8186) );
  XNOR U9663 ( .A(b[2622]), .B(n8187), .Z(n8188) );
  XNOR U9664 ( .A(b[2622]), .B(n8189), .Z(c[2622]) );
  XNOR U9665 ( .A(a[2622]), .B(n8190), .Z(n8189) );
  IV U9666 ( .A(n8187), .Z(n8190) );
  XOR U9667 ( .A(n8191), .B(n8192), .Z(n8187) );
  ANDN U9668 ( .B(n8193), .A(n8194), .Z(n8191) );
  XNOR U9669 ( .A(b[2621]), .B(n8192), .Z(n8193) );
  XNOR U9670 ( .A(b[2621]), .B(n8194), .Z(c[2621]) );
  XNOR U9671 ( .A(a[2621]), .B(n8195), .Z(n8194) );
  IV U9672 ( .A(n8192), .Z(n8195) );
  XOR U9673 ( .A(n8196), .B(n8197), .Z(n8192) );
  ANDN U9674 ( .B(n8198), .A(n8199), .Z(n8196) );
  XNOR U9675 ( .A(b[2620]), .B(n8197), .Z(n8198) );
  XNOR U9676 ( .A(b[2620]), .B(n8199), .Z(c[2620]) );
  XNOR U9677 ( .A(a[2620]), .B(n8200), .Z(n8199) );
  IV U9678 ( .A(n8197), .Z(n8200) );
  XOR U9679 ( .A(n8201), .B(n8202), .Z(n8197) );
  ANDN U9680 ( .B(n8203), .A(n8204), .Z(n8201) );
  XNOR U9681 ( .A(b[2619]), .B(n8202), .Z(n8203) );
  XNOR U9682 ( .A(b[261]), .B(n8205), .Z(c[261]) );
  XNOR U9683 ( .A(b[2619]), .B(n8204), .Z(c[2619]) );
  XNOR U9684 ( .A(a[2619]), .B(n8206), .Z(n8204) );
  IV U9685 ( .A(n8202), .Z(n8206) );
  XOR U9686 ( .A(n8207), .B(n8208), .Z(n8202) );
  ANDN U9687 ( .B(n8209), .A(n8210), .Z(n8207) );
  XNOR U9688 ( .A(b[2618]), .B(n8208), .Z(n8209) );
  XNOR U9689 ( .A(b[2618]), .B(n8210), .Z(c[2618]) );
  XNOR U9690 ( .A(a[2618]), .B(n8211), .Z(n8210) );
  IV U9691 ( .A(n8208), .Z(n8211) );
  XOR U9692 ( .A(n8212), .B(n8213), .Z(n8208) );
  ANDN U9693 ( .B(n8214), .A(n8215), .Z(n8212) );
  XNOR U9694 ( .A(b[2617]), .B(n8213), .Z(n8214) );
  XNOR U9695 ( .A(b[2617]), .B(n8215), .Z(c[2617]) );
  XNOR U9696 ( .A(a[2617]), .B(n8216), .Z(n8215) );
  IV U9697 ( .A(n8213), .Z(n8216) );
  XOR U9698 ( .A(n8217), .B(n8218), .Z(n8213) );
  ANDN U9699 ( .B(n8219), .A(n8220), .Z(n8217) );
  XNOR U9700 ( .A(b[2616]), .B(n8218), .Z(n8219) );
  XNOR U9701 ( .A(b[2616]), .B(n8220), .Z(c[2616]) );
  XNOR U9702 ( .A(a[2616]), .B(n8221), .Z(n8220) );
  IV U9703 ( .A(n8218), .Z(n8221) );
  XOR U9704 ( .A(n8222), .B(n8223), .Z(n8218) );
  ANDN U9705 ( .B(n8224), .A(n8225), .Z(n8222) );
  XNOR U9706 ( .A(b[2615]), .B(n8223), .Z(n8224) );
  XNOR U9707 ( .A(b[2615]), .B(n8225), .Z(c[2615]) );
  XNOR U9708 ( .A(a[2615]), .B(n8226), .Z(n8225) );
  IV U9709 ( .A(n8223), .Z(n8226) );
  XOR U9710 ( .A(n8227), .B(n8228), .Z(n8223) );
  ANDN U9711 ( .B(n8229), .A(n8230), .Z(n8227) );
  XNOR U9712 ( .A(b[2614]), .B(n8228), .Z(n8229) );
  XNOR U9713 ( .A(b[2614]), .B(n8230), .Z(c[2614]) );
  XNOR U9714 ( .A(a[2614]), .B(n8231), .Z(n8230) );
  IV U9715 ( .A(n8228), .Z(n8231) );
  XOR U9716 ( .A(n8232), .B(n8233), .Z(n8228) );
  ANDN U9717 ( .B(n8234), .A(n8235), .Z(n8232) );
  XNOR U9718 ( .A(b[2613]), .B(n8233), .Z(n8234) );
  XNOR U9719 ( .A(b[2613]), .B(n8235), .Z(c[2613]) );
  XNOR U9720 ( .A(a[2613]), .B(n8236), .Z(n8235) );
  IV U9721 ( .A(n8233), .Z(n8236) );
  XOR U9722 ( .A(n8237), .B(n8238), .Z(n8233) );
  ANDN U9723 ( .B(n8239), .A(n8240), .Z(n8237) );
  XNOR U9724 ( .A(b[2612]), .B(n8238), .Z(n8239) );
  XNOR U9725 ( .A(b[2612]), .B(n8240), .Z(c[2612]) );
  XNOR U9726 ( .A(a[2612]), .B(n8241), .Z(n8240) );
  IV U9727 ( .A(n8238), .Z(n8241) );
  XOR U9728 ( .A(n8242), .B(n8243), .Z(n8238) );
  ANDN U9729 ( .B(n8244), .A(n8245), .Z(n8242) );
  XNOR U9730 ( .A(b[2611]), .B(n8243), .Z(n8244) );
  XNOR U9731 ( .A(b[2611]), .B(n8245), .Z(c[2611]) );
  XNOR U9732 ( .A(a[2611]), .B(n8246), .Z(n8245) );
  IV U9733 ( .A(n8243), .Z(n8246) );
  XOR U9734 ( .A(n8247), .B(n8248), .Z(n8243) );
  ANDN U9735 ( .B(n8249), .A(n8250), .Z(n8247) );
  XNOR U9736 ( .A(b[2610]), .B(n8248), .Z(n8249) );
  XNOR U9737 ( .A(b[2610]), .B(n8250), .Z(c[2610]) );
  XNOR U9738 ( .A(a[2610]), .B(n8251), .Z(n8250) );
  IV U9739 ( .A(n8248), .Z(n8251) );
  XOR U9740 ( .A(n8252), .B(n8253), .Z(n8248) );
  ANDN U9741 ( .B(n8254), .A(n8255), .Z(n8252) );
  XNOR U9742 ( .A(b[2609]), .B(n8253), .Z(n8254) );
  XNOR U9743 ( .A(b[260]), .B(n8256), .Z(c[260]) );
  XNOR U9744 ( .A(b[2609]), .B(n8255), .Z(c[2609]) );
  XNOR U9745 ( .A(a[2609]), .B(n8257), .Z(n8255) );
  IV U9746 ( .A(n8253), .Z(n8257) );
  XOR U9747 ( .A(n8258), .B(n8259), .Z(n8253) );
  ANDN U9748 ( .B(n8260), .A(n8261), .Z(n8258) );
  XNOR U9749 ( .A(b[2608]), .B(n8259), .Z(n8260) );
  XNOR U9750 ( .A(b[2608]), .B(n8261), .Z(c[2608]) );
  XNOR U9751 ( .A(a[2608]), .B(n8262), .Z(n8261) );
  IV U9752 ( .A(n8259), .Z(n8262) );
  XOR U9753 ( .A(n8263), .B(n8264), .Z(n8259) );
  ANDN U9754 ( .B(n8265), .A(n8266), .Z(n8263) );
  XNOR U9755 ( .A(b[2607]), .B(n8264), .Z(n8265) );
  XNOR U9756 ( .A(b[2607]), .B(n8266), .Z(c[2607]) );
  XNOR U9757 ( .A(a[2607]), .B(n8267), .Z(n8266) );
  IV U9758 ( .A(n8264), .Z(n8267) );
  XOR U9759 ( .A(n8268), .B(n8269), .Z(n8264) );
  ANDN U9760 ( .B(n8270), .A(n8271), .Z(n8268) );
  XNOR U9761 ( .A(b[2606]), .B(n8269), .Z(n8270) );
  XNOR U9762 ( .A(b[2606]), .B(n8271), .Z(c[2606]) );
  XNOR U9763 ( .A(a[2606]), .B(n8272), .Z(n8271) );
  IV U9764 ( .A(n8269), .Z(n8272) );
  XOR U9765 ( .A(n8273), .B(n8274), .Z(n8269) );
  ANDN U9766 ( .B(n8275), .A(n8276), .Z(n8273) );
  XNOR U9767 ( .A(b[2605]), .B(n8274), .Z(n8275) );
  XNOR U9768 ( .A(b[2605]), .B(n8276), .Z(c[2605]) );
  XNOR U9769 ( .A(a[2605]), .B(n8277), .Z(n8276) );
  IV U9770 ( .A(n8274), .Z(n8277) );
  XOR U9771 ( .A(n8278), .B(n8279), .Z(n8274) );
  ANDN U9772 ( .B(n8280), .A(n8281), .Z(n8278) );
  XNOR U9773 ( .A(b[2604]), .B(n8279), .Z(n8280) );
  XNOR U9774 ( .A(b[2604]), .B(n8281), .Z(c[2604]) );
  XNOR U9775 ( .A(a[2604]), .B(n8282), .Z(n8281) );
  IV U9776 ( .A(n8279), .Z(n8282) );
  XOR U9777 ( .A(n8283), .B(n8284), .Z(n8279) );
  ANDN U9778 ( .B(n8285), .A(n8286), .Z(n8283) );
  XNOR U9779 ( .A(b[2603]), .B(n8284), .Z(n8285) );
  XNOR U9780 ( .A(b[2603]), .B(n8286), .Z(c[2603]) );
  XNOR U9781 ( .A(a[2603]), .B(n8287), .Z(n8286) );
  IV U9782 ( .A(n8284), .Z(n8287) );
  XOR U9783 ( .A(n8288), .B(n8289), .Z(n8284) );
  ANDN U9784 ( .B(n8290), .A(n8291), .Z(n8288) );
  XNOR U9785 ( .A(b[2602]), .B(n8289), .Z(n8290) );
  XNOR U9786 ( .A(b[2602]), .B(n8291), .Z(c[2602]) );
  XNOR U9787 ( .A(a[2602]), .B(n8292), .Z(n8291) );
  IV U9788 ( .A(n8289), .Z(n8292) );
  XOR U9789 ( .A(n8293), .B(n8294), .Z(n8289) );
  ANDN U9790 ( .B(n8295), .A(n8296), .Z(n8293) );
  XNOR U9791 ( .A(b[2601]), .B(n8294), .Z(n8295) );
  XNOR U9792 ( .A(b[2601]), .B(n8296), .Z(c[2601]) );
  XNOR U9793 ( .A(a[2601]), .B(n8297), .Z(n8296) );
  IV U9794 ( .A(n8294), .Z(n8297) );
  XOR U9795 ( .A(n8298), .B(n8299), .Z(n8294) );
  ANDN U9796 ( .B(n8300), .A(n8301), .Z(n8298) );
  XNOR U9797 ( .A(b[2600]), .B(n8299), .Z(n8300) );
  XNOR U9798 ( .A(b[2600]), .B(n8301), .Z(c[2600]) );
  XNOR U9799 ( .A(a[2600]), .B(n8302), .Z(n8301) );
  IV U9800 ( .A(n8299), .Z(n8302) );
  XOR U9801 ( .A(n8303), .B(n8304), .Z(n8299) );
  ANDN U9802 ( .B(n8305), .A(n8306), .Z(n8303) );
  XNOR U9803 ( .A(b[2599]), .B(n8304), .Z(n8305) );
  XNOR U9804 ( .A(b[25]), .B(n8307), .Z(c[25]) );
  XNOR U9805 ( .A(b[259]), .B(n8308), .Z(c[259]) );
  XNOR U9806 ( .A(b[2599]), .B(n8306), .Z(c[2599]) );
  XNOR U9807 ( .A(a[2599]), .B(n8309), .Z(n8306) );
  IV U9808 ( .A(n8304), .Z(n8309) );
  XOR U9809 ( .A(n8310), .B(n8311), .Z(n8304) );
  ANDN U9810 ( .B(n8312), .A(n8313), .Z(n8310) );
  XNOR U9811 ( .A(b[2598]), .B(n8311), .Z(n8312) );
  XNOR U9812 ( .A(b[2598]), .B(n8313), .Z(c[2598]) );
  XNOR U9813 ( .A(a[2598]), .B(n8314), .Z(n8313) );
  IV U9814 ( .A(n8311), .Z(n8314) );
  XOR U9815 ( .A(n8315), .B(n8316), .Z(n8311) );
  ANDN U9816 ( .B(n8317), .A(n8318), .Z(n8315) );
  XNOR U9817 ( .A(b[2597]), .B(n8316), .Z(n8317) );
  XNOR U9818 ( .A(b[2597]), .B(n8318), .Z(c[2597]) );
  XNOR U9819 ( .A(a[2597]), .B(n8319), .Z(n8318) );
  IV U9820 ( .A(n8316), .Z(n8319) );
  XOR U9821 ( .A(n8320), .B(n8321), .Z(n8316) );
  ANDN U9822 ( .B(n8322), .A(n8323), .Z(n8320) );
  XNOR U9823 ( .A(b[2596]), .B(n8321), .Z(n8322) );
  XNOR U9824 ( .A(b[2596]), .B(n8323), .Z(c[2596]) );
  XNOR U9825 ( .A(a[2596]), .B(n8324), .Z(n8323) );
  IV U9826 ( .A(n8321), .Z(n8324) );
  XOR U9827 ( .A(n8325), .B(n8326), .Z(n8321) );
  ANDN U9828 ( .B(n8327), .A(n8328), .Z(n8325) );
  XNOR U9829 ( .A(b[2595]), .B(n8326), .Z(n8327) );
  XNOR U9830 ( .A(b[2595]), .B(n8328), .Z(c[2595]) );
  XNOR U9831 ( .A(a[2595]), .B(n8329), .Z(n8328) );
  IV U9832 ( .A(n8326), .Z(n8329) );
  XOR U9833 ( .A(n8330), .B(n8331), .Z(n8326) );
  ANDN U9834 ( .B(n8332), .A(n8333), .Z(n8330) );
  XNOR U9835 ( .A(b[2594]), .B(n8331), .Z(n8332) );
  XNOR U9836 ( .A(b[2594]), .B(n8333), .Z(c[2594]) );
  XNOR U9837 ( .A(a[2594]), .B(n8334), .Z(n8333) );
  IV U9838 ( .A(n8331), .Z(n8334) );
  XOR U9839 ( .A(n8335), .B(n8336), .Z(n8331) );
  ANDN U9840 ( .B(n8337), .A(n8338), .Z(n8335) );
  XNOR U9841 ( .A(b[2593]), .B(n8336), .Z(n8337) );
  XNOR U9842 ( .A(b[2593]), .B(n8338), .Z(c[2593]) );
  XNOR U9843 ( .A(a[2593]), .B(n8339), .Z(n8338) );
  IV U9844 ( .A(n8336), .Z(n8339) );
  XOR U9845 ( .A(n8340), .B(n8341), .Z(n8336) );
  ANDN U9846 ( .B(n8342), .A(n8343), .Z(n8340) );
  XNOR U9847 ( .A(b[2592]), .B(n8341), .Z(n8342) );
  XNOR U9848 ( .A(b[2592]), .B(n8343), .Z(c[2592]) );
  XNOR U9849 ( .A(a[2592]), .B(n8344), .Z(n8343) );
  IV U9850 ( .A(n8341), .Z(n8344) );
  XOR U9851 ( .A(n8345), .B(n8346), .Z(n8341) );
  ANDN U9852 ( .B(n8347), .A(n8348), .Z(n8345) );
  XNOR U9853 ( .A(b[2591]), .B(n8346), .Z(n8347) );
  XNOR U9854 ( .A(b[2591]), .B(n8348), .Z(c[2591]) );
  XNOR U9855 ( .A(a[2591]), .B(n8349), .Z(n8348) );
  IV U9856 ( .A(n8346), .Z(n8349) );
  XOR U9857 ( .A(n8350), .B(n8351), .Z(n8346) );
  ANDN U9858 ( .B(n8352), .A(n8353), .Z(n8350) );
  XNOR U9859 ( .A(b[2590]), .B(n8351), .Z(n8352) );
  XNOR U9860 ( .A(b[2590]), .B(n8353), .Z(c[2590]) );
  XNOR U9861 ( .A(a[2590]), .B(n8354), .Z(n8353) );
  IV U9862 ( .A(n8351), .Z(n8354) );
  XOR U9863 ( .A(n8355), .B(n8356), .Z(n8351) );
  ANDN U9864 ( .B(n8357), .A(n8358), .Z(n8355) );
  XNOR U9865 ( .A(b[2589]), .B(n8356), .Z(n8357) );
  XNOR U9866 ( .A(b[258]), .B(n8359), .Z(c[258]) );
  XNOR U9867 ( .A(b[2589]), .B(n8358), .Z(c[2589]) );
  XNOR U9868 ( .A(a[2589]), .B(n8360), .Z(n8358) );
  IV U9869 ( .A(n8356), .Z(n8360) );
  XOR U9870 ( .A(n8361), .B(n8362), .Z(n8356) );
  ANDN U9871 ( .B(n8363), .A(n8364), .Z(n8361) );
  XNOR U9872 ( .A(b[2588]), .B(n8362), .Z(n8363) );
  XNOR U9873 ( .A(b[2588]), .B(n8364), .Z(c[2588]) );
  XNOR U9874 ( .A(a[2588]), .B(n8365), .Z(n8364) );
  IV U9875 ( .A(n8362), .Z(n8365) );
  XOR U9876 ( .A(n8366), .B(n8367), .Z(n8362) );
  ANDN U9877 ( .B(n8368), .A(n8369), .Z(n8366) );
  XNOR U9878 ( .A(b[2587]), .B(n8367), .Z(n8368) );
  XNOR U9879 ( .A(b[2587]), .B(n8369), .Z(c[2587]) );
  XNOR U9880 ( .A(a[2587]), .B(n8370), .Z(n8369) );
  IV U9881 ( .A(n8367), .Z(n8370) );
  XOR U9882 ( .A(n8371), .B(n8372), .Z(n8367) );
  ANDN U9883 ( .B(n8373), .A(n8374), .Z(n8371) );
  XNOR U9884 ( .A(b[2586]), .B(n8372), .Z(n8373) );
  XNOR U9885 ( .A(b[2586]), .B(n8374), .Z(c[2586]) );
  XNOR U9886 ( .A(a[2586]), .B(n8375), .Z(n8374) );
  IV U9887 ( .A(n8372), .Z(n8375) );
  XOR U9888 ( .A(n8376), .B(n8377), .Z(n8372) );
  ANDN U9889 ( .B(n8378), .A(n8379), .Z(n8376) );
  XNOR U9890 ( .A(b[2585]), .B(n8377), .Z(n8378) );
  XNOR U9891 ( .A(b[2585]), .B(n8379), .Z(c[2585]) );
  XNOR U9892 ( .A(a[2585]), .B(n8380), .Z(n8379) );
  IV U9893 ( .A(n8377), .Z(n8380) );
  XOR U9894 ( .A(n8381), .B(n8382), .Z(n8377) );
  ANDN U9895 ( .B(n8383), .A(n8384), .Z(n8381) );
  XNOR U9896 ( .A(b[2584]), .B(n8382), .Z(n8383) );
  XNOR U9897 ( .A(b[2584]), .B(n8384), .Z(c[2584]) );
  XNOR U9898 ( .A(a[2584]), .B(n8385), .Z(n8384) );
  IV U9899 ( .A(n8382), .Z(n8385) );
  XOR U9900 ( .A(n8386), .B(n8387), .Z(n8382) );
  ANDN U9901 ( .B(n8388), .A(n8389), .Z(n8386) );
  XNOR U9902 ( .A(b[2583]), .B(n8387), .Z(n8388) );
  XNOR U9903 ( .A(b[2583]), .B(n8389), .Z(c[2583]) );
  XNOR U9904 ( .A(a[2583]), .B(n8390), .Z(n8389) );
  IV U9905 ( .A(n8387), .Z(n8390) );
  XOR U9906 ( .A(n8391), .B(n8392), .Z(n8387) );
  ANDN U9907 ( .B(n8393), .A(n8394), .Z(n8391) );
  XNOR U9908 ( .A(b[2582]), .B(n8392), .Z(n8393) );
  XNOR U9909 ( .A(b[2582]), .B(n8394), .Z(c[2582]) );
  XNOR U9910 ( .A(a[2582]), .B(n8395), .Z(n8394) );
  IV U9911 ( .A(n8392), .Z(n8395) );
  XOR U9912 ( .A(n8396), .B(n8397), .Z(n8392) );
  ANDN U9913 ( .B(n8398), .A(n8399), .Z(n8396) );
  XNOR U9914 ( .A(b[2581]), .B(n8397), .Z(n8398) );
  XNOR U9915 ( .A(b[2581]), .B(n8399), .Z(c[2581]) );
  XNOR U9916 ( .A(a[2581]), .B(n8400), .Z(n8399) );
  IV U9917 ( .A(n8397), .Z(n8400) );
  XOR U9918 ( .A(n8401), .B(n8402), .Z(n8397) );
  ANDN U9919 ( .B(n8403), .A(n8404), .Z(n8401) );
  XNOR U9920 ( .A(b[2580]), .B(n8402), .Z(n8403) );
  XNOR U9921 ( .A(b[2580]), .B(n8404), .Z(c[2580]) );
  XNOR U9922 ( .A(a[2580]), .B(n8405), .Z(n8404) );
  IV U9923 ( .A(n8402), .Z(n8405) );
  XOR U9924 ( .A(n8406), .B(n8407), .Z(n8402) );
  ANDN U9925 ( .B(n8408), .A(n8409), .Z(n8406) );
  XNOR U9926 ( .A(b[2579]), .B(n8407), .Z(n8408) );
  XNOR U9927 ( .A(b[257]), .B(n8410), .Z(c[257]) );
  XNOR U9928 ( .A(b[2579]), .B(n8409), .Z(c[2579]) );
  XNOR U9929 ( .A(a[2579]), .B(n8411), .Z(n8409) );
  IV U9930 ( .A(n8407), .Z(n8411) );
  XOR U9931 ( .A(n8412), .B(n8413), .Z(n8407) );
  ANDN U9932 ( .B(n8414), .A(n8415), .Z(n8412) );
  XNOR U9933 ( .A(b[2578]), .B(n8413), .Z(n8414) );
  XNOR U9934 ( .A(b[2578]), .B(n8415), .Z(c[2578]) );
  XNOR U9935 ( .A(a[2578]), .B(n8416), .Z(n8415) );
  IV U9936 ( .A(n8413), .Z(n8416) );
  XOR U9937 ( .A(n8417), .B(n8418), .Z(n8413) );
  ANDN U9938 ( .B(n8419), .A(n8420), .Z(n8417) );
  XNOR U9939 ( .A(b[2577]), .B(n8418), .Z(n8419) );
  XNOR U9940 ( .A(b[2577]), .B(n8420), .Z(c[2577]) );
  XNOR U9941 ( .A(a[2577]), .B(n8421), .Z(n8420) );
  IV U9942 ( .A(n8418), .Z(n8421) );
  XOR U9943 ( .A(n8422), .B(n8423), .Z(n8418) );
  ANDN U9944 ( .B(n8424), .A(n8425), .Z(n8422) );
  XNOR U9945 ( .A(b[2576]), .B(n8423), .Z(n8424) );
  XNOR U9946 ( .A(b[2576]), .B(n8425), .Z(c[2576]) );
  XNOR U9947 ( .A(a[2576]), .B(n8426), .Z(n8425) );
  IV U9948 ( .A(n8423), .Z(n8426) );
  XOR U9949 ( .A(n8427), .B(n8428), .Z(n8423) );
  ANDN U9950 ( .B(n8429), .A(n8430), .Z(n8427) );
  XNOR U9951 ( .A(b[2575]), .B(n8428), .Z(n8429) );
  XNOR U9952 ( .A(b[2575]), .B(n8430), .Z(c[2575]) );
  XNOR U9953 ( .A(a[2575]), .B(n8431), .Z(n8430) );
  IV U9954 ( .A(n8428), .Z(n8431) );
  XOR U9955 ( .A(n8432), .B(n8433), .Z(n8428) );
  ANDN U9956 ( .B(n8434), .A(n8435), .Z(n8432) );
  XNOR U9957 ( .A(b[2574]), .B(n8433), .Z(n8434) );
  XNOR U9958 ( .A(b[2574]), .B(n8435), .Z(c[2574]) );
  XNOR U9959 ( .A(a[2574]), .B(n8436), .Z(n8435) );
  IV U9960 ( .A(n8433), .Z(n8436) );
  XOR U9961 ( .A(n8437), .B(n8438), .Z(n8433) );
  ANDN U9962 ( .B(n8439), .A(n8440), .Z(n8437) );
  XNOR U9963 ( .A(b[2573]), .B(n8438), .Z(n8439) );
  XNOR U9964 ( .A(b[2573]), .B(n8440), .Z(c[2573]) );
  XNOR U9965 ( .A(a[2573]), .B(n8441), .Z(n8440) );
  IV U9966 ( .A(n8438), .Z(n8441) );
  XOR U9967 ( .A(n8442), .B(n8443), .Z(n8438) );
  ANDN U9968 ( .B(n8444), .A(n8445), .Z(n8442) );
  XNOR U9969 ( .A(b[2572]), .B(n8443), .Z(n8444) );
  XNOR U9970 ( .A(b[2572]), .B(n8445), .Z(c[2572]) );
  XNOR U9971 ( .A(a[2572]), .B(n8446), .Z(n8445) );
  IV U9972 ( .A(n8443), .Z(n8446) );
  XOR U9973 ( .A(n8447), .B(n8448), .Z(n8443) );
  ANDN U9974 ( .B(n8449), .A(n8450), .Z(n8447) );
  XNOR U9975 ( .A(b[2571]), .B(n8448), .Z(n8449) );
  XNOR U9976 ( .A(b[2571]), .B(n8450), .Z(c[2571]) );
  XNOR U9977 ( .A(a[2571]), .B(n8451), .Z(n8450) );
  IV U9978 ( .A(n8448), .Z(n8451) );
  XOR U9979 ( .A(n8452), .B(n8453), .Z(n8448) );
  ANDN U9980 ( .B(n8454), .A(n8455), .Z(n8452) );
  XNOR U9981 ( .A(b[2570]), .B(n8453), .Z(n8454) );
  XNOR U9982 ( .A(b[2570]), .B(n8455), .Z(c[2570]) );
  XNOR U9983 ( .A(a[2570]), .B(n8456), .Z(n8455) );
  IV U9984 ( .A(n8453), .Z(n8456) );
  XOR U9985 ( .A(n8457), .B(n8458), .Z(n8453) );
  ANDN U9986 ( .B(n8459), .A(n8460), .Z(n8457) );
  XNOR U9987 ( .A(b[2569]), .B(n8458), .Z(n8459) );
  XNOR U9988 ( .A(b[256]), .B(n8461), .Z(c[256]) );
  XNOR U9989 ( .A(b[2569]), .B(n8460), .Z(c[2569]) );
  XNOR U9990 ( .A(a[2569]), .B(n8462), .Z(n8460) );
  IV U9991 ( .A(n8458), .Z(n8462) );
  XOR U9992 ( .A(n8463), .B(n8464), .Z(n8458) );
  ANDN U9993 ( .B(n8465), .A(n8466), .Z(n8463) );
  XNOR U9994 ( .A(b[2568]), .B(n8464), .Z(n8465) );
  XNOR U9995 ( .A(b[2568]), .B(n8466), .Z(c[2568]) );
  XNOR U9996 ( .A(a[2568]), .B(n8467), .Z(n8466) );
  IV U9997 ( .A(n8464), .Z(n8467) );
  XOR U9998 ( .A(n8468), .B(n8469), .Z(n8464) );
  ANDN U9999 ( .B(n8470), .A(n8471), .Z(n8468) );
  XNOR U10000 ( .A(b[2567]), .B(n8469), .Z(n8470) );
  XNOR U10001 ( .A(b[2567]), .B(n8471), .Z(c[2567]) );
  XNOR U10002 ( .A(a[2567]), .B(n8472), .Z(n8471) );
  IV U10003 ( .A(n8469), .Z(n8472) );
  XOR U10004 ( .A(n8473), .B(n8474), .Z(n8469) );
  ANDN U10005 ( .B(n8475), .A(n8476), .Z(n8473) );
  XNOR U10006 ( .A(b[2566]), .B(n8474), .Z(n8475) );
  XNOR U10007 ( .A(b[2566]), .B(n8476), .Z(c[2566]) );
  XNOR U10008 ( .A(a[2566]), .B(n8477), .Z(n8476) );
  IV U10009 ( .A(n8474), .Z(n8477) );
  XOR U10010 ( .A(n8478), .B(n8479), .Z(n8474) );
  ANDN U10011 ( .B(n8480), .A(n8481), .Z(n8478) );
  XNOR U10012 ( .A(b[2565]), .B(n8479), .Z(n8480) );
  XNOR U10013 ( .A(b[2565]), .B(n8481), .Z(c[2565]) );
  XNOR U10014 ( .A(a[2565]), .B(n8482), .Z(n8481) );
  IV U10015 ( .A(n8479), .Z(n8482) );
  XOR U10016 ( .A(n8483), .B(n8484), .Z(n8479) );
  ANDN U10017 ( .B(n8485), .A(n8486), .Z(n8483) );
  XNOR U10018 ( .A(b[2564]), .B(n8484), .Z(n8485) );
  XNOR U10019 ( .A(b[2564]), .B(n8486), .Z(c[2564]) );
  XNOR U10020 ( .A(a[2564]), .B(n8487), .Z(n8486) );
  IV U10021 ( .A(n8484), .Z(n8487) );
  XOR U10022 ( .A(n8488), .B(n8489), .Z(n8484) );
  ANDN U10023 ( .B(n8490), .A(n8491), .Z(n8488) );
  XNOR U10024 ( .A(b[2563]), .B(n8489), .Z(n8490) );
  XNOR U10025 ( .A(b[2563]), .B(n8491), .Z(c[2563]) );
  XNOR U10026 ( .A(a[2563]), .B(n8492), .Z(n8491) );
  IV U10027 ( .A(n8489), .Z(n8492) );
  XOR U10028 ( .A(n8493), .B(n8494), .Z(n8489) );
  ANDN U10029 ( .B(n8495), .A(n8496), .Z(n8493) );
  XNOR U10030 ( .A(b[2562]), .B(n8494), .Z(n8495) );
  XNOR U10031 ( .A(b[2562]), .B(n8496), .Z(c[2562]) );
  XNOR U10032 ( .A(a[2562]), .B(n8497), .Z(n8496) );
  IV U10033 ( .A(n8494), .Z(n8497) );
  XOR U10034 ( .A(n8498), .B(n8499), .Z(n8494) );
  ANDN U10035 ( .B(n8500), .A(n8501), .Z(n8498) );
  XNOR U10036 ( .A(b[2561]), .B(n8499), .Z(n8500) );
  XNOR U10037 ( .A(b[2561]), .B(n8501), .Z(c[2561]) );
  XNOR U10038 ( .A(a[2561]), .B(n8502), .Z(n8501) );
  IV U10039 ( .A(n8499), .Z(n8502) );
  XOR U10040 ( .A(n8503), .B(n8504), .Z(n8499) );
  ANDN U10041 ( .B(n8505), .A(n8506), .Z(n8503) );
  XNOR U10042 ( .A(b[2560]), .B(n8504), .Z(n8505) );
  XNOR U10043 ( .A(b[2560]), .B(n8506), .Z(c[2560]) );
  XNOR U10044 ( .A(a[2560]), .B(n8507), .Z(n8506) );
  IV U10045 ( .A(n8504), .Z(n8507) );
  XOR U10046 ( .A(n8508), .B(n8509), .Z(n8504) );
  ANDN U10047 ( .B(n8510), .A(n8511), .Z(n8508) );
  XNOR U10048 ( .A(b[2559]), .B(n8509), .Z(n8510) );
  XNOR U10049 ( .A(b[255]), .B(n8512), .Z(c[255]) );
  XNOR U10050 ( .A(b[2559]), .B(n8511), .Z(c[2559]) );
  XNOR U10051 ( .A(a[2559]), .B(n8513), .Z(n8511) );
  IV U10052 ( .A(n8509), .Z(n8513) );
  XOR U10053 ( .A(n8514), .B(n8515), .Z(n8509) );
  ANDN U10054 ( .B(n8516), .A(n8517), .Z(n8514) );
  XNOR U10055 ( .A(b[2558]), .B(n8515), .Z(n8516) );
  XNOR U10056 ( .A(b[2558]), .B(n8517), .Z(c[2558]) );
  XNOR U10057 ( .A(a[2558]), .B(n8518), .Z(n8517) );
  IV U10058 ( .A(n8515), .Z(n8518) );
  XOR U10059 ( .A(n8519), .B(n8520), .Z(n8515) );
  ANDN U10060 ( .B(n8521), .A(n8522), .Z(n8519) );
  XNOR U10061 ( .A(b[2557]), .B(n8520), .Z(n8521) );
  XNOR U10062 ( .A(b[2557]), .B(n8522), .Z(c[2557]) );
  XNOR U10063 ( .A(a[2557]), .B(n8523), .Z(n8522) );
  IV U10064 ( .A(n8520), .Z(n8523) );
  XOR U10065 ( .A(n8524), .B(n8525), .Z(n8520) );
  ANDN U10066 ( .B(n8526), .A(n8527), .Z(n8524) );
  XNOR U10067 ( .A(b[2556]), .B(n8525), .Z(n8526) );
  XNOR U10068 ( .A(b[2556]), .B(n8527), .Z(c[2556]) );
  XNOR U10069 ( .A(a[2556]), .B(n8528), .Z(n8527) );
  IV U10070 ( .A(n8525), .Z(n8528) );
  XOR U10071 ( .A(n8529), .B(n8530), .Z(n8525) );
  ANDN U10072 ( .B(n8531), .A(n8532), .Z(n8529) );
  XNOR U10073 ( .A(b[2555]), .B(n8530), .Z(n8531) );
  XNOR U10074 ( .A(b[2555]), .B(n8532), .Z(c[2555]) );
  XNOR U10075 ( .A(a[2555]), .B(n8533), .Z(n8532) );
  IV U10076 ( .A(n8530), .Z(n8533) );
  XOR U10077 ( .A(n8534), .B(n8535), .Z(n8530) );
  ANDN U10078 ( .B(n8536), .A(n8537), .Z(n8534) );
  XNOR U10079 ( .A(b[2554]), .B(n8535), .Z(n8536) );
  XNOR U10080 ( .A(b[2554]), .B(n8537), .Z(c[2554]) );
  XNOR U10081 ( .A(a[2554]), .B(n8538), .Z(n8537) );
  IV U10082 ( .A(n8535), .Z(n8538) );
  XOR U10083 ( .A(n8539), .B(n8540), .Z(n8535) );
  ANDN U10084 ( .B(n8541), .A(n8542), .Z(n8539) );
  XNOR U10085 ( .A(b[2553]), .B(n8540), .Z(n8541) );
  XNOR U10086 ( .A(b[2553]), .B(n8542), .Z(c[2553]) );
  XNOR U10087 ( .A(a[2553]), .B(n8543), .Z(n8542) );
  IV U10088 ( .A(n8540), .Z(n8543) );
  XOR U10089 ( .A(n8544), .B(n8545), .Z(n8540) );
  ANDN U10090 ( .B(n8546), .A(n8547), .Z(n8544) );
  XNOR U10091 ( .A(b[2552]), .B(n8545), .Z(n8546) );
  XNOR U10092 ( .A(b[2552]), .B(n8547), .Z(c[2552]) );
  XNOR U10093 ( .A(a[2552]), .B(n8548), .Z(n8547) );
  IV U10094 ( .A(n8545), .Z(n8548) );
  XOR U10095 ( .A(n8549), .B(n8550), .Z(n8545) );
  ANDN U10096 ( .B(n8551), .A(n8552), .Z(n8549) );
  XNOR U10097 ( .A(b[2551]), .B(n8550), .Z(n8551) );
  XNOR U10098 ( .A(b[2551]), .B(n8552), .Z(c[2551]) );
  XNOR U10099 ( .A(a[2551]), .B(n8553), .Z(n8552) );
  IV U10100 ( .A(n8550), .Z(n8553) );
  XOR U10101 ( .A(n8554), .B(n8555), .Z(n8550) );
  ANDN U10102 ( .B(n8556), .A(n8557), .Z(n8554) );
  XNOR U10103 ( .A(b[2550]), .B(n8555), .Z(n8556) );
  XNOR U10104 ( .A(b[2550]), .B(n8557), .Z(c[2550]) );
  XNOR U10105 ( .A(a[2550]), .B(n8558), .Z(n8557) );
  IV U10106 ( .A(n8555), .Z(n8558) );
  XOR U10107 ( .A(n8559), .B(n8560), .Z(n8555) );
  ANDN U10108 ( .B(n8561), .A(n8562), .Z(n8559) );
  XNOR U10109 ( .A(b[2549]), .B(n8560), .Z(n8561) );
  XNOR U10110 ( .A(b[254]), .B(n8563), .Z(c[254]) );
  XNOR U10111 ( .A(b[2549]), .B(n8562), .Z(c[2549]) );
  XNOR U10112 ( .A(a[2549]), .B(n8564), .Z(n8562) );
  IV U10113 ( .A(n8560), .Z(n8564) );
  XOR U10114 ( .A(n8565), .B(n8566), .Z(n8560) );
  ANDN U10115 ( .B(n8567), .A(n8568), .Z(n8565) );
  XNOR U10116 ( .A(b[2548]), .B(n8566), .Z(n8567) );
  XNOR U10117 ( .A(b[2548]), .B(n8568), .Z(c[2548]) );
  XNOR U10118 ( .A(a[2548]), .B(n8569), .Z(n8568) );
  IV U10119 ( .A(n8566), .Z(n8569) );
  XOR U10120 ( .A(n8570), .B(n8571), .Z(n8566) );
  ANDN U10121 ( .B(n8572), .A(n8573), .Z(n8570) );
  XNOR U10122 ( .A(b[2547]), .B(n8571), .Z(n8572) );
  XNOR U10123 ( .A(b[2547]), .B(n8573), .Z(c[2547]) );
  XNOR U10124 ( .A(a[2547]), .B(n8574), .Z(n8573) );
  IV U10125 ( .A(n8571), .Z(n8574) );
  XOR U10126 ( .A(n8575), .B(n8576), .Z(n8571) );
  ANDN U10127 ( .B(n8577), .A(n8578), .Z(n8575) );
  XNOR U10128 ( .A(b[2546]), .B(n8576), .Z(n8577) );
  XNOR U10129 ( .A(b[2546]), .B(n8578), .Z(c[2546]) );
  XNOR U10130 ( .A(a[2546]), .B(n8579), .Z(n8578) );
  IV U10131 ( .A(n8576), .Z(n8579) );
  XOR U10132 ( .A(n8580), .B(n8581), .Z(n8576) );
  ANDN U10133 ( .B(n8582), .A(n8583), .Z(n8580) );
  XNOR U10134 ( .A(b[2545]), .B(n8581), .Z(n8582) );
  XNOR U10135 ( .A(b[2545]), .B(n8583), .Z(c[2545]) );
  XNOR U10136 ( .A(a[2545]), .B(n8584), .Z(n8583) );
  IV U10137 ( .A(n8581), .Z(n8584) );
  XOR U10138 ( .A(n8585), .B(n8586), .Z(n8581) );
  ANDN U10139 ( .B(n8587), .A(n8588), .Z(n8585) );
  XNOR U10140 ( .A(b[2544]), .B(n8586), .Z(n8587) );
  XNOR U10141 ( .A(b[2544]), .B(n8588), .Z(c[2544]) );
  XNOR U10142 ( .A(a[2544]), .B(n8589), .Z(n8588) );
  IV U10143 ( .A(n8586), .Z(n8589) );
  XOR U10144 ( .A(n8590), .B(n8591), .Z(n8586) );
  ANDN U10145 ( .B(n8592), .A(n8593), .Z(n8590) );
  XNOR U10146 ( .A(b[2543]), .B(n8591), .Z(n8592) );
  XNOR U10147 ( .A(b[2543]), .B(n8593), .Z(c[2543]) );
  XNOR U10148 ( .A(a[2543]), .B(n8594), .Z(n8593) );
  IV U10149 ( .A(n8591), .Z(n8594) );
  XOR U10150 ( .A(n8595), .B(n8596), .Z(n8591) );
  ANDN U10151 ( .B(n8597), .A(n8598), .Z(n8595) );
  XNOR U10152 ( .A(b[2542]), .B(n8596), .Z(n8597) );
  XNOR U10153 ( .A(b[2542]), .B(n8598), .Z(c[2542]) );
  XNOR U10154 ( .A(a[2542]), .B(n8599), .Z(n8598) );
  IV U10155 ( .A(n8596), .Z(n8599) );
  XOR U10156 ( .A(n8600), .B(n8601), .Z(n8596) );
  ANDN U10157 ( .B(n8602), .A(n8603), .Z(n8600) );
  XNOR U10158 ( .A(b[2541]), .B(n8601), .Z(n8602) );
  XNOR U10159 ( .A(b[2541]), .B(n8603), .Z(c[2541]) );
  XNOR U10160 ( .A(a[2541]), .B(n8604), .Z(n8603) );
  IV U10161 ( .A(n8601), .Z(n8604) );
  XOR U10162 ( .A(n8605), .B(n8606), .Z(n8601) );
  ANDN U10163 ( .B(n8607), .A(n8608), .Z(n8605) );
  XNOR U10164 ( .A(b[2540]), .B(n8606), .Z(n8607) );
  XNOR U10165 ( .A(b[2540]), .B(n8608), .Z(c[2540]) );
  XNOR U10166 ( .A(a[2540]), .B(n8609), .Z(n8608) );
  IV U10167 ( .A(n8606), .Z(n8609) );
  XOR U10168 ( .A(n8610), .B(n8611), .Z(n8606) );
  ANDN U10169 ( .B(n8612), .A(n8613), .Z(n8610) );
  XNOR U10170 ( .A(b[2539]), .B(n8611), .Z(n8612) );
  XNOR U10171 ( .A(b[253]), .B(n8614), .Z(c[253]) );
  XNOR U10172 ( .A(b[2539]), .B(n8613), .Z(c[2539]) );
  XNOR U10173 ( .A(a[2539]), .B(n8615), .Z(n8613) );
  IV U10174 ( .A(n8611), .Z(n8615) );
  XOR U10175 ( .A(n8616), .B(n8617), .Z(n8611) );
  ANDN U10176 ( .B(n8618), .A(n8619), .Z(n8616) );
  XNOR U10177 ( .A(b[2538]), .B(n8617), .Z(n8618) );
  XNOR U10178 ( .A(b[2538]), .B(n8619), .Z(c[2538]) );
  XNOR U10179 ( .A(a[2538]), .B(n8620), .Z(n8619) );
  IV U10180 ( .A(n8617), .Z(n8620) );
  XOR U10181 ( .A(n8621), .B(n8622), .Z(n8617) );
  ANDN U10182 ( .B(n8623), .A(n8624), .Z(n8621) );
  XNOR U10183 ( .A(b[2537]), .B(n8622), .Z(n8623) );
  XNOR U10184 ( .A(b[2537]), .B(n8624), .Z(c[2537]) );
  XNOR U10185 ( .A(a[2537]), .B(n8625), .Z(n8624) );
  IV U10186 ( .A(n8622), .Z(n8625) );
  XOR U10187 ( .A(n8626), .B(n8627), .Z(n8622) );
  ANDN U10188 ( .B(n8628), .A(n8629), .Z(n8626) );
  XNOR U10189 ( .A(b[2536]), .B(n8627), .Z(n8628) );
  XNOR U10190 ( .A(b[2536]), .B(n8629), .Z(c[2536]) );
  XNOR U10191 ( .A(a[2536]), .B(n8630), .Z(n8629) );
  IV U10192 ( .A(n8627), .Z(n8630) );
  XOR U10193 ( .A(n8631), .B(n8632), .Z(n8627) );
  ANDN U10194 ( .B(n8633), .A(n8634), .Z(n8631) );
  XNOR U10195 ( .A(b[2535]), .B(n8632), .Z(n8633) );
  XNOR U10196 ( .A(b[2535]), .B(n8634), .Z(c[2535]) );
  XNOR U10197 ( .A(a[2535]), .B(n8635), .Z(n8634) );
  IV U10198 ( .A(n8632), .Z(n8635) );
  XOR U10199 ( .A(n8636), .B(n8637), .Z(n8632) );
  ANDN U10200 ( .B(n8638), .A(n8639), .Z(n8636) );
  XNOR U10201 ( .A(b[2534]), .B(n8637), .Z(n8638) );
  XNOR U10202 ( .A(b[2534]), .B(n8639), .Z(c[2534]) );
  XNOR U10203 ( .A(a[2534]), .B(n8640), .Z(n8639) );
  IV U10204 ( .A(n8637), .Z(n8640) );
  XOR U10205 ( .A(n8641), .B(n8642), .Z(n8637) );
  ANDN U10206 ( .B(n8643), .A(n8644), .Z(n8641) );
  XNOR U10207 ( .A(b[2533]), .B(n8642), .Z(n8643) );
  XNOR U10208 ( .A(b[2533]), .B(n8644), .Z(c[2533]) );
  XNOR U10209 ( .A(a[2533]), .B(n8645), .Z(n8644) );
  IV U10210 ( .A(n8642), .Z(n8645) );
  XOR U10211 ( .A(n8646), .B(n8647), .Z(n8642) );
  ANDN U10212 ( .B(n8648), .A(n8649), .Z(n8646) );
  XNOR U10213 ( .A(b[2532]), .B(n8647), .Z(n8648) );
  XNOR U10214 ( .A(b[2532]), .B(n8649), .Z(c[2532]) );
  XNOR U10215 ( .A(a[2532]), .B(n8650), .Z(n8649) );
  IV U10216 ( .A(n8647), .Z(n8650) );
  XOR U10217 ( .A(n8651), .B(n8652), .Z(n8647) );
  ANDN U10218 ( .B(n8653), .A(n8654), .Z(n8651) );
  XNOR U10219 ( .A(b[2531]), .B(n8652), .Z(n8653) );
  XNOR U10220 ( .A(b[2531]), .B(n8654), .Z(c[2531]) );
  XNOR U10221 ( .A(a[2531]), .B(n8655), .Z(n8654) );
  IV U10222 ( .A(n8652), .Z(n8655) );
  XOR U10223 ( .A(n8656), .B(n8657), .Z(n8652) );
  ANDN U10224 ( .B(n8658), .A(n8659), .Z(n8656) );
  XNOR U10225 ( .A(b[2530]), .B(n8657), .Z(n8658) );
  XNOR U10226 ( .A(b[2530]), .B(n8659), .Z(c[2530]) );
  XNOR U10227 ( .A(a[2530]), .B(n8660), .Z(n8659) );
  IV U10228 ( .A(n8657), .Z(n8660) );
  XOR U10229 ( .A(n8661), .B(n8662), .Z(n8657) );
  ANDN U10230 ( .B(n8663), .A(n8664), .Z(n8661) );
  XNOR U10231 ( .A(b[2529]), .B(n8662), .Z(n8663) );
  XNOR U10232 ( .A(b[252]), .B(n8665), .Z(c[252]) );
  XNOR U10233 ( .A(b[2529]), .B(n8664), .Z(c[2529]) );
  XNOR U10234 ( .A(a[2529]), .B(n8666), .Z(n8664) );
  IV U10235 ( .A(n8662), .Z(n8666) );
  XOR U10236 ( .A(n8667), .B(n8668), .Z(n8662) );
  ANDN U10237 ( .B(n8669), .A(n8670), .Z(n8667) );
  XNOR U10238 ( .A(b[2528]), .B(n8668), .Z(n8669) );
  XNOR U10239 ( .A(b[2528]), .B(n8670), .Z(c[2528]) );
  XNOR U10240 ( .A(a[2528]), .B(n8671), .Z(n8670) );
  IV U10241 ( .A(n8668), .Z(n8671) );
  XOR U10242 ( .A(n8672), .B(n8673), .Z(n8668) );
  ANDN U10243 ( .B(n8674), .A(n8675), .Z(n8672) );
  XNOR U10244 ( .A(b[2527]), .B(n8673), .Z(n8674) );
  XNOR U10245 ( .A(b[2527]), .B(n8675), .Z(c[2527]) );
  XNOR U10246 ( .A(a[2527]), .B(n8676), .Z(n8675) );
  IV U10247 ( .A(n8673), .Z(n8676) );
  XOR U10248 ( .A(n8677), .B(n8678), .Z(n8673) );
  ANDN U10249 ( .B(n8679), .A(n8680), .Z(n8677) );
  XNOR U10250 ( .A(b[2526]), .B(n8678), .Z(n8679) );
  XNOR U10251 ( .A(b[2526]), .B(n8680), .Z(c[2526]) );
  XNOR U10252 ( .A(a[2526]), .B(n8681), .Z(n8680) );
  IV U10253 ( .A(n8678), .Z(n8681) );
  XOR U10254 ( .A(n8682), .B(n8683), .Z(n8678) );
  ANDN U10255 ( .B(n8684), .A(n8685), .Z(n8682) );
  XNOR U10256 ( .A(b[2525]), .B(n8683), .Z(n8684) );
  XNOR U10257 ( .A(b[2525]), .B(n8685), .Z(c[2525]) );
  XNOR U10258 ( .A(a[2525]), .B(n8686), .Z(n8685) );
  IV U10259 ( .A(n8683), .Z(n8686) );
  XOR U10260 ( .A(n8687), .B(n8688), .Z(n8683) );
  ANDN U10261 ( .B(n8689), .A(n8690), .Z(n8687) );
  XNOR U10262 ( .A(b[2524]), .B(n8688), .Z(n8689) );
  XNOR U10263 ( .A(b[2524]), .B(n8690), .Z(c[2524]) );
  XNOR U10264 ( .A(a[2524]), .B(n8691), .Z(n8690) );
  IV U10265 ( .A(n8688), .Z(n8691) );
  XOR U10266 ( .A(n8692), .B(n8693), .Z(n8688) );
  ANDN U10267 ( .B(n8694), .A(n8695), .Z(n8692) );
  XNOR U10268 ( .A(b[2523]), .B(n8693), .Z(n8694) );
  XNOR U10269 ( .A(b[2523]), .B(n8695), .Z(c[2523]) );
  XNOR U10270 ( .A(a[2523]), .B(n8696), .Z(n8695) );
  IV U10271 ( .A(n8693), .Z(n8696) );
  XOR U10272 ( .A(n8697), .B(n8698), .Z(n8693) );
  ANDN U10273 ( .B(n8699), .A(n8700), .Z(n8697) );
  XNOR U10274 ( .A(b[2522]), .B(n8698), .Z(n8699) );
  XNOR U10275 ( .A(b[2522]), .B(n8700), .Z(c[2522]) );
  XNOR U10276 ( .A(a[2522]), .B(n8701), .Z(n8700) );
  IV U10277 ( .A(n8698), .Z(n8701) );
  XOR U10278 ( .A(n8702), .B(n8703), .Z(n8698) );
  ANDN U10279 ( .B(n8704), .A(n8705), .Z(n8702) );
  XNOR U10280 ( .A(b[2521]), .B(n8703), .Z(n8704) );
  XNOR U10281 ( .A(b[2521]), .B(n8705), .Z(c[2521]) );
  XNOR U10282 ( .A(a[2521]), .B(n8706), .Z(n8705) );
  IV U10283 ( .A(n8703), .Z(n8706) );
  XOR U10284 ( .A(n8707), .B(n8708), .Z(n8703) );
  ANDN U10285 ( .B(n8709), .A(n8710), .Z(n8707) );
  XNOR U10286 ( .A(b[2520]), .B(n8708), .Z(n8709) );
  XNOR U10287 ( .A(b[2520]), .B(n8710), .Z(c[2520]) );
  XNOR U10288 ( .A(a[2520]), .B(n8711), .Z(n8710) );
  IV U10289 ( .A(n8708), .Z(n8711) );
  XOR U10290 ( .A(n8712), .B(n8713), .Z(n8708) );
  ANDN U10291 ( .B(n8714), .A(n8715), .Z(n8712) );
  XNOR U10292 ( .A(b[2519]), .B(n8713), .Z(n8714) );
  XNOR U10293 ( .A(b[251]), .B(n8716), .Z(c[251]) );
  XNOR U10294 ( .A(b[2519]), .B(n8715), .Z(c[2519]) );
  XNOR U10295 ( .A(a[2519]), .B(n8717), .Z(n8715) );
  IV U10296 ( .A(n8713), .Z(n8717) );
  XOR U10297 ( .A(n8718), .B(n8719), .Z(n8713) );
  ANDN U10298 ( .B(n8720), .A(n8721), .Z(n8718) );
  XNOR U10299 ( .A(b[2518]), .B(n8719), .Z(n8720) );
  XNOR U10300 ( .A(b[2518]), .B(n8721), .Z(c[2518]) );
  XNOR U10301 ( .A(a[2518]), .B(n8722), .Z(n8721) );
  IV U10302 ( .A(n8719), .Z(n8722) );
  XOR U10303 ( .A(n8723), .B(n8724), .Z(n8719) );
  ANDN U10304 ( .B(n8725), .A(n8726), .Z(n8723) );
  XNOR U10305 ( .A(b[2517]), .B(n8724), .Z(n8725) );
  XNOR U10306 ( .A(b[2517]), .B(n8726), .Z(c[2517]) );
  XNOR U10307 ( .A(a[2517]), .B(n8727), .Z(n8726) );
  IV U10308 ( .A(n8724), .Z(n8727) );
  XOR U10309 ( .A(n8728), .B(n8729), .Z(n8724) );
  ANDN U10310 ( .B(n8730), .A(n8731), .Z(n8728) );
  XNOR U10311 ( .A(b[2516]), .B(n8729), .Z(n8730) );
  XNOR U10312 ( .A(b[2516]), .B(n8731), .Z(c[2516]) );
  XNOR U10313 ( .A(a[2516]), .B(n8732), .Z(n8731) );
  IV U10314 ( .A(n8729), .Z(n8732) );
  XOR U10315 ( .A(n8733), .B(n8734), .Z(n8729) );
  ANDN U10316 ( .B(n8735), .A(n8736), .Z(n8733) );
  XNOR U10317 ( .A(b[2515]), .B(n8734), .Z(n8735) );
  XNOR U10318 ( .A(b[2515]), .B(n8736), .Z(c[2515]) );
  XNOR U10319 ( .A(a[2515]), .B(n8737), .Z(n8736) );
  IV U10320 ( .A(n8734), .Z(n8737) );
  XOR U10321 ( .A(n8738), .B(n8739), .Z(n8734) );
  ANDN U10322 ( .B(n8740), .A(n8741), .Z(n8738) );
  XNOR U10323 ( .A(b[2514]), .B(n8739), .Z(n8740) );
  XNOR U10324 ( .A(b[2514]), .B(n8741), .Z(c[2514]) );
  XNOR U10325 ( .A(a[2514]), .B(n8742), .Z(n8741) );
  IV U10326 ( .A(n8739), .Z(n8742) );
  XOR U10327 ( .A(n8743), .B(n8744), .Z(n8739) );
  ANDN U10328 ( .B(n8745), .A(n8746), .Z(n8743) );
  XNOR U10329 ( .A(b[2513]), .B(n8744), .Z(n8745) );
  XNOR U10330 ( .A(b[2513]), .B(n8746), .Z(c[2513]) );
  XNOR U10331 ( .A(a[2513]), .B(n8747), .Z(n8746) );
  IV U10332 ( .A(n8744), .Z(n8747) );
  XOR U10333 ( .A(n8748), .B(n8749), .Z(n8744) );
  ANDN U10334 ( .B(n8750), .A(n8751), .Z(n8748) );
  XNOR U10335 ( .A(b[2512]), .B(n8749), .Z(n8750) );
  XNOR U10336 ( .A(b[2512]), .B(n8751), .Z(c[2512]) );
  XNOR U10337 ( .A(a[2512]), .B(n8752), .Z(n8751) );
  IV U10338 ( .A(n8749), .Z(n8752) );
  XOR U10339 ( .A(n8753), .B(n8754), .Z(n8749) );
  ANDN U10340 ( .B(n8755), .A(n8756), .Z(n8753) );
  XNOR U10341 ( .A(b[2511]), .B(n8754), .Z(n8755) );
  XNOR U10342 ( .A(b[2511]), .B(n8756), .Z(c[2511]) );
  XNOR U10343 ( .A(a[2511]), .B(n8757), .Z(n8756) );
  IV U10344 ( .A(n8754), .Z(n8757) );
  XOR U10345 ( .A(n8758), .B(n8759), .Z(n8754) );
  ANDN U10346 ( .B(n8760), .A(n8761), .Z(n8758) );
  XNOR U10347 ( .A(b[2510]), .B(n8759), .Z(n8760) );
  XNOR U10348 ( .A(b[2510]), .B(n8761), .Z(c[2510]) );
  XNOR U10349 ( .A(a[2510]), .B(n8762), .Z(n8761) );
  IV U10350 ( .A(n8759), .Z(n8762) );
  XOR U10351 ( .A(n8763), .B(n8764), .Z(n8759) );
  ANDN U10352 ( .B(n8765), .A(n8766), .Z(n8763) );
  XNOR U10353 ( .A(b[2509]), .B(n8764), .Z(n8765) );
  XNOR U10354 ( .A(b[250]), .B(n8767), .Z(c[250]) );
  XNOR U10355 ( .A(b[2509]), .B(n8766), .Z(c[2509]) );
  XNOR U10356 ( .A(a[2509]), .B(n8768), .Z(n8766) );
  IV U10357 ( .A(n8764), .Z(n8768) );
  XOR U10358 ( .A(n8769), .B(n8770), .Z(n8764) );
  ANDN U10359 ( .B(n8771), .A(n8772), .Z(n8769) );
  XNOR U10360 ( .A(b[2508]), .B(n8770), .Z(n8771) );
  XNOR U10361 ( .A(b[2508]), .B(n8772), .Z(c[2508]) );
  XNOR U10362 ( .A(a[2508]), .B(n8773), .Z(n8772) );
  IV U10363 ( .A(n8770), .Z(n8773) );
  XOR U10364 ( .A(n8774), .B(n8775), .Z(n8770) );
  ANDN U10365 ( .B(n8776), .A(n8777), .Z(n8774) );
  XNOR U10366 ( .A(b[2507]), .B(n8775), .Z(n8776) );
  XNOR U10367 ( .A(b[2507]), .B(n8777), .Z(c[2507]) );
  XNOR U10368 ( .A(a[2507]), .B(n8778), .Z(n8777) );
  IV U10369 ( .A(n8775), .Z(n8778) );
  XOR U10370 ( .A(n8779), .B(n8780), .Z(n8775) );
  ANDN U10371 ( .B(n8781), .A(n8782), .Z(n8779) );
  XNOR U10372 ( .A(b[2506]), .B(n8780), .Z(n8781) );
  XNOR U10373 ( .A(b[2506]), .B(n8782), .Z(c[2506]) );
  XNOR U10374 ( .A(a[2506]), .B(n8783), .Z(n8782) );
  IV U10375 ( .A(n8780), .Z(n8783) );
  XOR U10376 ( .A(n8784), .B(n8785), .Z(n8780) );
  ANDN U10377 ( .B(n8786), .A(n8787), .Z(n8784) );
  XNOR U10378 ( .A(b[2505]), .B(n8785), .Z(n8786) );
  XNOR U10379 ( .A(b[2505]), .B(n8787), .Z(c[2505]) );
  XNOR U10380 ( .A(a[2505]), .B(n8788), .Z(n8787) );
  IV U10381 ( .A(n8785), .Z(n8788) );
  XOR U10382 ( .A(n8789), .B(n8790), .Z(n8785) );
  ANDN U10383 ( .B(n8791), .A(n8792), .Z(n8789) );
  XNOR U10384 ( .A(b[2504]), .B(n8790), .Z(n8791) );
  XNOR U10385 ( .A(b[2504]), .B(n8792), .Z(c[2504]) );
  XNOR U10386 ( .A(a[2504]), .B(n8793), .Z(n8792) );
  IV U10387 ( .A(n8790), .Z(n8793) );
  XOR U10388 ( .A(n8794), .B(n8795), .Z(n8790) );
  ANDN U10389 ( .B(n8796), .A(n8797), .Z(n8794) );
  XNOR U10390 ( .A(b[2503]), .B(n8795), .Z(n8796) );
  XNOR U10391 ( .A(b[2503]), .B(n8797), .Z(c[2503]) );
  XNOR U10392 ( .A(a[2503]), .B(n8798), .Z(n8797) );
  IV U10393 ( .A(n8795), .Z(n8798) );
  XOR U10394 ( .A(n8799), .B(n8800), .Z(n8795) );
  ANDN U10395 ( .B(n8801), .A(n8802), .Z(n8799) );
  XNOR U10396 ( .A(b[2502]), .B(n8800), .Z(n8801) );
  XNOR U10397 ( .A(b[2502]), .B(n8802), .Z(c[2502]) );
  XNOR U10398 ( .A(a[2502]), .B(n8803), .Z(n8802) );
  IV U10399 ( .A(n8800), .Z(n8803) );
  XOR U10400 ( .A(n8804), .B(n8805), .Z(n8800) );
  ANDN U10401 ( .B(n8806), .A(n8807), .Z(n8804) );
  XNOR U10402 ( .A(b[2501]), .B(n8805), .Z(n8806) );
  XNOR U10403 ( .A(b[2501]), .B(n8807), .Z(c[2501]) );
  XNOR U10404 ( .A(a[2501]), .B(n8808), .Z(n8807) );
  IV U10405 ( .A(n8805), .Z(n8808) );
  XOR U10406 ( .A(n8809), .B(n8810), .Z(n8805) );
  ANDN U10407 ( .B(n8811), .A(n8812), .Z(n8809) );
  XNOR U10408 ( .A(b[2500]), .B(n8810), .Z(n8811) );
  XNOR U10409 ( .A(b[2500]), .B(n8812), .Z(c[2500]) );
  XNOR U10410 ( .A(a[2500]), .B(n8813), .Z(n8812) );
  IV U10411 ( .A(n8810), .Z(n8813) );
  XOR U10412 ( .A(n8814), .B(n8815), .Z(n8810) );
  ANDN U10413 ( .B(n8816), .A(n8817), .Z(n8814) );
  XNOR U10414 ( .A(b[2499]), .B(n8815), .Z(n8816) );
  XNOR U10415 ( .A(b[24]), .B(n8818), .Z(c[24]) );
  XNOR U10416 ( .A(b[249]), .B(n8819), .Z(c[249]) );
  XNOR U10417 ( .A(b[2499]), .B(n8817), .Z(c[2499]) );
  XNOR U10418 ( .A(a[2499]), .B(n8820), .Z(n8817) );
  IV U10419 ( .A(n8815), .Z(n8820) );
  XOR U10420 ( .A(n8821), .B(n8822), .Z(n8815) );
  ANDN U10421 ( .B(n8823), .A(n8824), .Z(n8821) );
  XNOR U10422 ( .A(b[2498]), .B(n8822), .Z(n8823) );
  XNOR U10423 ( .A(b[2498]), .B(n8824), .Z(c[2498]) );
  XNOR U10424 ( .A(a[2498]), .B(n8825), .Z(n8824) );
  IV U10425 ( .A(n8822), .Z(n8825) );
  XOR U10426 ( .A(n8826), .B(n8827), .Z(n8822) );
  ANDN U10427 ( .B(n8828), .A(n8829), .Z(n8826) );
  XNOR U10428 ( .A(b[2497]), .B(n8827), .Z(n8828) );
  XNOR U10429 ( .A(b[2497]), .B(n8829), .Z(c[2497]) );
  XNOR U10430 ( .A(a[2497]), .B(n8830), .Z(n8829) );
  IV U10431 ( .A(n8827), .Z(n8830) );
  XOR U10432 ( .A(n8831), .B(n8832), .Z(n8827) );
  ANDN U10433 ( .B(n8833), .A(n8834), .Z(n8831) );
  XNOR U10434 ( .A(b[2496]), .B(n8832), .Z(n8833) );
  XNOR U10435 ( .A(b[2496]), .B(n8834), .Z(c[2496]) );
  XNOR U10436 ( .A(a[2496]), .B(n8835), .Z(n8834) );
  IV U10437 ( .A(n8832), .Z(n8835) );
  XOR U10438 ( .A(n8836), .B(n8837), .Z(n8832) );
  ANDN U10439 ( .B(n8838), .A(n8839), .Z(n8836) );
  XNOR U10440 ( .A(b[2495]), .B(n8837), .Z(n8838) );
  XNOR U10441 ( .A(b[2495]), .B(n8839), .Z(c[2495]) );
  XNOR U10442 ( .A(a[2495]), .B(n8840), .Z(n8839) );
  IV U10443 ( .A(n8837), .Z(n8840) );
  XOR U10444 ( .A(n8841), .B(n8842), .Z(n8837) );
  ANDN U10445 ( .B(n8843), .A(n8844), .Z(n8841) );
  XNOR U10446 ( .A(b[2494]), .B(n8842), .Z(n8843) );
  XNOR U10447 ( .A(b[2494]), .B(n8844), .Z(c[2494]) );
  XNOR U10448 ( .A(a[2494]), .B(n8845), .Z(n8844) );
  IV U10449 ( .A(n8842), .Z(n8845) );
  XOR U10450 ( .A(n8846), .B(n8847), .Z(n8842) );
  ANDN U10451 ( .B(n8848), .A(n8849), .Z(n8846) );
  XNOR U10452 ( .A(b[2493]), .B(n8847), .Z(n8848) );
  XNOR U10453 ( .A(b[2493]), .B(n8849), .Z(c[2493]) );
  XNOR U10454 ( .A(a[2493]), .B(n8850), .Z(n8849) );
  IV U10455 ( .A(n8847), .Z(n8850) );
  XOR U10456 ( .A(n8851), .B(n8852), .Z(n8847) );
  ANDN U10457 ( .B(n8853), .A(n8854), .Z(n8851) );
  XNOR U10458 ( .A(b[2492]), .B(n8852), .Z(n8853) );
  XNOR U10459 ( .A(b[2492]), .B(n8854), .Z(c[2492]) );
  XNOR U10460 ( .A(a[2492]), .B(n8855), .Z(n8854) );
  IV U10461 ( .A(n8852), .Z(n8855) );
  XOR U10462 ( .A(n8856), .B(n8857), .Z(n8852) );
  ANDN U10463 ( .B(n8858), .A(n8859), .Z(n8856) );
  XNOR U10464 ( .A(b[2491]), .B(n8857), .Z(n8858) );
  XNOR U10465 ( .A(b[2491]), .B(n8859), .Z(c[2491]) );
  XNOR U10466 ( .A(a[2491]), .B(n8860), .Z(n8859) );
  IV U10467 ( .A(n8857), .Z(n8860) );
  XOR U10468 ( .A(n8861), .B(n8862), .Z(n8857) );
  ANDN U10469 ( .B(n8863), .A(n8864), .Z(n8861) );
  XNOR U10470 ( .A(b[2490]), .B(n8862), .Z(n8863) );
  XNOR U10471 ( .A(b[2490]), .B(n8864), .Z(c[2490]) );
  XNOR U10472 ( .A(a[2490]), .B(n8865), .Z(n8864) );
  IV U10473 ( .A(n8862), .Z(n8865) );
  XOR U10474 ( .A(n8866), .B(n8867), .Z(n8862) );
  ANDN U10475 ( .B(n8868), .A(n8869), .Z(n8866) );
  XNOR U10476 ( .A(b[2489]), .B(n8867), .Z(n8868) );
  XNOR U10477 ( .A(b[248]), .B(n8870), .Z(c[248]) );
  XNOR U10478 ( .A(b[2489]), .B(n8869), .Z(c[2489]) );
  XNOR U10479 ( .A(a[2489]), .B(n8871), .Z(n8869) );
  IV U10480 ( .A(n8867), .Z(n8871) );
  XOR U10481 ( .A(n8872), .B(n8873), .Z(n8867) );
  ANDN U10482 ( .B(n8874), .A(n8875), .Z(n8872) );
  XNOR U10483 ( .A(b[2488]), .B(n8873), .Z(n8874) );
  XNOR U10484 ( .A(b[2488]), .B(n8875), .Z(c[2488]) );
  XNOR U10485 ( .A(a[2488]), .B(n8876), .Z(n8875) );
  IV U10486 ( .A(n8873), .Z(n8876) );
  XOR U10487 ( .A(n8877), .B(n8878), .Z(n8873) );
  ANDN U10488 ( .B(n8879), .A(n8880), .Z(n8877) );
  XNOR U10489 ( .A(b[2487]), .B(n8878), .Z(n8879) );
  XNOR U10490 ( .A(b[2487]), .B(n8880), .Z(c[2487]) );
  XNOR U10491 ( .A(a[2487]), .B(n8881), .Z(n8880) );
  IV U10492 ( .A(n8878), .Z(n8881) );
  XOR U10493 ( .A(n8882), .B(n8883), .Z(n8878) );
  ANDN U10494 ( .B(n8884), .A(n8885), .Z(n8882) );
  XNOR U10495 ( .A(b[2486]), .B(n8883), .Z(n8884) );
  XNOR U10496 ( .A(b[2486]), .B(n8885), .Z(c[2486]) );
  XNOR U10497 ( .A(a[2486]), .B(n8886), .Z(n8885) );
  IV U10498 ( .A(n8883), .Z(n8886) );
  XOR U10499 ( .A(n8887), .B(n8888), .Z(n8883) );
  ANDN U10500 ( .B(n8889), .A(n8890), .Z(n8887) );
  XNOR U10501 ( .A(b[2485]), .B(n8888), .Z(n8889) );
  XNOR U10502 ( .A(b[2485]), .B(n8890), .Z(c[2485]) );
  XNOR U10503 ( .A(a[2485]), .B(n8891), .Z(n8890) );
  IV U10504 ( .A(n8888), .Z(n8891) );
  XOR U10505 ( .A(n8892), .B(n8893), .Z(n8888) );
  ANDN U10506 ( .B(n8894), .A(n8895), .Z(n8892) );
  XNOR U10507 ( .A(b[2484]), .B(n8893), .Z(n8894) );
  XNOR U10508 ( .A(b[2484]), .B(n8895), .Z(c[2484]) );
  XNOR U10509 ( .A(a[2484]), .B(n8896), .Z(n8895) );
  IV U10510 ( .A(n8893), .Z(n8896) );
  XOR U10511 ( .A(n8897), .B(n8898), .Z(n8893) );
  ANDN U10512 ( .B(n8899), .A(n8900), .Z(n8897) );
  XNOR U10513 ( .A(b[2483]), .B(n8898), .Z(n8899) );
  XNOR U10514 ( .A(b[2483]), .B(n8900), .Z(c[2483]) );
  XNOR U10515 ( .A(a[2483]), .B(n8901), .Z(n8900) );
  IV U10516 ( .A(n8898), .Z(n8901) );
  XOR U10517 ( .A(n8902), .B(n8903), .Z(n8898) );
  ANDN U10518 ( .B(n8904), .A(n8905), .Z(n8902) );
  XNOR U10519 ( .A(b[2482]), .B(n8903), .Z(n8904) );
  XNOR U10520 ( .A(b[2482]), .B(n8905), .Z(c[2482]) );
  XNOR U10521 ( .A(a[2482]), .B(n8906), .Z(n8905) );
  IV U10522 ( .A(n8903), .Z(n8906) );
  XOR U10523 ( .A(n8907), .B(n8908), .Z(n8903) );
  ANDN U10524 ( .B(n8909), .A(n8910), .Z(n8907) );
  XNOR U10525 ( .A(b[2481]), .B(n8908), .Z(n8909) );
  XNOR U10526 ( .A(b[2481]), .B(n8910), .Z(c[2481]) );
  XNOR U10527 ( .A(a[2481]), .B(n8911), .Z(n8910) );
  IV U10528 ( .A(n8908), .Z(n8911) );
  XOR U10529 ( .A(n8912), .B(n8913), .Z(n8908) );
  ANDN U10530 ( .B(n8914), .A(n8915), .Z(n8912) );
  XNOR U10531 ( .A(b[2480]), .B(n8913), .Z(n8914) );
  XNOR U10532 ( .A(b[2480]), .B(n8915), .Z(c[2480]) );
  XNOR U10533 ( .A(a[2480]), .B(n8916), .Z(n8915) );
  IV U10534 ( .A(n8913), .Z(n8916) );
  XOR U10535 ( .A(n8917), .B(n8918), .Z(n8913) );
  ANDN U10536 ( .B(n8919), .A(n8920), .Z(n8917) );
  XNOR U10537 ( .A(b[2479]), .B(n8918), .Z(n8919) );
  XNOR U10538 ( .A(b[247]), .B(n8921), .Z(c[247]) );
  XNOR U10539 ( .A(b[2479]), .B(n8920), .Z(c[2479]) );
  XNOR U10540 ( .A(a[2479]), .B(n8922), .Z(n8920) );
  IV U10541 ( .A(n8918), .Z(n8922) );
  XOR U10542 ( .A(n8923), .B(n8924), .Z(n8918) );
  ANDN U10543 ( .B(n8925), .A(n8926), .Z(n8923) );
  XNOR U10544 ( .A(b[2478]), .B(n8924), .Z(n8925) );
  XNOR U10545 ( .A(b[2478]), .B(n8926), .Z(c[2478]) );
  XNOR U10546 ( .A(a[2478]), .B(n8927), .Z(n8926) );
  IV U10547 ( .A(n8924), .Z(n8927) );
  XOR U10548 ( .A(n8928), .B(n8929), .Z(n8924) );
  ANDN U10549 ( .B(n8930), .A(n8931), .Z(n8928) );
  XNOR U10550 ( .A(b[2477]), .B(n8929), .Z(n8930) );
  XNOR U10551 ( .A(b[2477]), .B(n8931), .Z(c[2477]) );
  XNOR U10552 ( .A(a[2477]), .B(n8932), .Z(n8931) );
  IV U10553 ( .A(n8929), .Z(n8932) );
  XOR U10554 ( .A(n8933), .B(n8934), .Z(n8929) );
  ANDN U10555 ( .B(n8935), .A(n8936), .Z(n8933) );
  XNOR U10556 ( .A(b[2476]), .B(n8934), .Z(n8935) );
  XNOR U10557 ( .A(b[2476]), .B(n8936), .Z(c[2476]) );
  XNOR U10558 ( .A(a[2476]), .B(n8937), .Z(n8936) );
  IV U10559 ( .A(n8934), .Z(n8937) );
  XOR U10560 ( .A(n8938), .B(n8939), .Z(n8934) );
  ANDN U10561 ( .B(n8940), .A(n8941), .Z(n8938) );
  XNOR U10562 ( .A(b[2475]), .B(n8939), .Z(n8940) );
  XNOR U10563 ( .A(b[2475]), .B(n8941), .Z(c[2475]) );
  XNOR U10564 ( .A(a[2475]), .B(n8942), .Z(n8941) );
  IV U10565 ( .A(n8939), .Z(n8942) );
  XOR U10566 ( .A(n8943), .B(n8944), .Z(n8939) );
  ANDN U10567 ( .B(n8945), .A(n8946), .Z(n8943) );
  XNOR U10568 ( .A(b[2474]), .B(n8944), .Z(n8945) );
  XNOR U10569 ( .A(b[2474]), .B(n8946), .Z(c[2474]) );
  XNOR U10570 ( .A(a[2474]), .B(n8947), .Z(n8946) );
  IV U10571 ( .A(n8944), .Z(n8947) );
  XOR U10572 ( .A(n8948), .B(n8949), .Z(n8944) );
  ANDN U10573 ( .B(n8950), .A(n8951), .Z(n8948) );
  XNOR U10574 ( .A(b[2473]), .B(n8949), .Z(n8950) );
  XNOR U10575 ( .A(b[2473]), .B(n8951), .Z(c[2473]) );
  XNOR U10576 ( .A(a[2473]), .B(n8952), .Z(n8951) );
  IV U10577 ( .A(n8949), .Z(n8952) );
  XOR U10578 ( .A(n8953), .B(n8954), .Z(n8949) );
  ANDN U10579 ( .B(n8955), .A(n8956), .Z(n8953) );
  XNOR U10580 ( .A(b[2472]), .B(n8954), .Z(n8955) );
  XNOR U10581 ( .A(b[2472]), .B(n8956), .Z(c[2472]) );
  XNOR U10582 ( .A(a[2472]), .B(n8957), .Z(n8956) );
  IV U10583 ( .A(n8954), .Z(n8957) );
  XOR U10584 ( .A(n8958), .B(n8959), .Z(n8954) );
  ANDN U10585 ( .B(n8960), .A(n8961), .Z(n8958) );
  XNOR U10586 ( .A(b[2471]), .B(n8959), .Z(n8960) );
  XNOR U10587 ( .A(b[2471]), .B(n8961), .Z(c[2471]) );
  XNOR U10588 ( .A(a[2471]), .B(n8962), .Z(n8961) );
  IV U10589 ( .A(n8959), .Z(n8962) );
  XOR U10590 ( .A(n8963), .B(n8964), .Z(n8959) );
  ANDN U10591 ( .B(n8965), .A(n8966), .Z(n8963) );
  XNOR U10592 ( .A(b[2470]), .B(n8964), .Z(n8965) );
  XNOR U10593 ( .A(b[2470]), .B(n8966), .Z(c[2470]) );
  XNOR U10594 ( .A(a[2470]), .B(n8967), .Z(n8966) );
  IV U10595 ( .A(n8964), .Z(n8967) );
  XOR U10596 ( .A(n8968), .B(n8969), .Z(n8964) );
  ANDN U10597 ( .B(n8970), .A(n8971), .Z(n8968) );
  XNOR U10598 ( .A(b[2469]), .B(n8969), .Z(n8970) );
  XNOR U10599 ( .A(b[246]), .B(n8972), .Z(c[246]) );
  XNOR U10600 ( .A(b[2469]), .B(n8971), .Z(c[2469]) );
  XNOR U10601 ( .A(a[2469]), .B(n8973), .Z(n8971) );
  IV U10602 ( .A(n8969), .Z(n8973) );
  XOR U10603 ( .A(n8974), .B(n8975), .Z(n8969) );
  ANDN U10604 ( .B(n8976), .A(n8977), .Z(n8974) );
  XNOR U10605 ( .A(b[2468]), .B(n8975), .Z(n8976) );
  XNOR U10606 ( .A(b[2468]), .B(n8977), .Z(c[2468]) );
  XNOR U10607 ( .A(a[2468]), .B(n8978), .Z(n8977) );
  IV U10608 ( .A(n8975), .Z(n8978) );
  XOR U10609 ( .A(n8979), .B(n8980), .Z(n8975) );
  ANDN U10610 ( .B(n8981), .A(n8982), .Z(n8979) );
  XNOR U10611 ( .A(b[2467]), .B(n8980), .Z(n8981) );
  XNOR U10612 ( .A(b[2467]), .B(n8982), .Z(c[2467]) );
  XNOR U10613 ( .A(a[2467]), .B(n8983), .Z(n8982) );
  IV U10614 ( .A(n8980), .Z(n8983) );
  XOR U10615 ( .A(n8984), .B(n8985), .Z(n8980) );
  ANDN U10616 ( .B(n8986), .A(n8987), .Z(n8984) );
  XNOR U10617 ( .A(b[2466]), .B(n8985), .Z(n8986) );
  XNOR U10618 ( .A(b[2466]), .B(n8987), .Z(c[2466]) );
  XNOR U10619 ( .A(a[2466]), .B(n8988), .Z(n8987) );
  IV U10620 ( .A(n8985), .Z(n8988) );
  XOR U10621 ( .A(n8989), .B(n8990), .Z(n8985) );
  ANDN U10622 ( .B(n8991), .A(n8992), .Z(n8989) );
  XNOR U10623 ( .A(b[2465]), .B(n8990), .Z(n8991) );
  XNOR U10624 ( .A(b[2465]), .B(n8992), .Z(c[2465]) );
  XNOR U10625 ( .A(a[2465]), .B(n8993), .Z(n8992) );
  IV U10626 ( .A(n8990), .Z(n8993) );
  XOR U10627 ( .A(n8994), .B(n8995), .Z(n8990) );
  ANDN U10628 ( .B(n8996), .A(n8997), .Z(n8994) );
  XNOR U10629 ( .A(b[2464]), .B(n8995), .Z(n8996) );
  XNOR U10630 ( .A(b[2464]), .B(n8997), .Z(c[2464]) );
  XNOR U10631 ( .A(a[2464]), .B(n8998), .Z(n8997) );
  IV U10632 ( .A(n8995), .Z(n8998) );
  XOR U10633 ( .A(n8999), .B(n9000), .Z(n8995) );
  ANDN U10634 ( .B(n9001), .A(n9002), .Z(n8999) );
  XNOR U10635 ( .A(b[2463]), .B(n9000), .Z(n9001) );
  XNOR U10636 ( .A(b[2463]), .B(n9002), .Z(c[2463]) );
  XNOR U10637 ( .A(a[2463]), .B(n9003), .Z(n9002) );
  IV U10638 ( .A(n9000), .Z(n9003) );
  XOR U10639 ( .A(n9004), .B(n9005), .Z(n9000) );
  ANDN U10640 ( .B(n9006), .A(n9007), .Z(n9004) );
  XNOR U10641 ( .A(b[2462]), .B(n9005), .Z(n9006) );
  XNOR U10642 ( .A(b[2462]), .B(n9007), .Z(c[2462]) );
  XNOR U10643 ( .A(a[2462]), .B(n9008), .Z(n9007) );
  IV U10644 ( .A(n9005), .Z(n9008) );
  XOR U10645 ( .A(n9009), .B(n9010), .Z(n9005) );
  ANDN U10646 ( .B(n9011), .A(n9012), .Z(n9009) );
  XNOR U10647 ( .A(b[2461]), .B(n9010), .Z(n9011) );
  XNOR U10648 ( .A(b[2461]), .B(n9012), .Z(c[2461]) );
  XNOR U10649 ( .A(a[2461]), .B(n9013), .Z(n9012) );
  IV U10650 ( .A(n9010), .Z(n9013) );
  XOR U10651 ( .A(n9014), .B(n9015), .Z(n9010) );
  ANDN U10652 ( .B(n9016), .A(n9017), .Z(n9014) );
  XNOR U10653 ( .A(b[2460]), .B(n9015), .Z(n9016) );
  XNOR U10654 ( .A(b[2460]), .B(n9017), .Z(c[2460]) );
  XNOR U10655 ( .A(a[2460]), .B(n9018), .Z(n9017) );
  IV U10656 ( .A(n9015), .Z(n9018) );
  XOR U10657 ( .A(n9019), .B(n9020), .Z(n9015) );
  ANDN U10658 ( .B(n9021), .A(n9022), .Z(n9019) );
  XNOR U10659 ( .A(b[2459]), .B(n9020), .Z(n9021) );
  XNOR U10660 ( .A(b[245]), .B(n9023), .Z(c[245]) );
  XNOR U10661 ( .A(b[2459]), .B(n9022), .Z(c[2459]) );
  XNOR U10662 ( .A(a[2459]), .B(n9024), .Z(n9022) );
  IV U10663 ( .A(n9020), .Z(n9024) );
  XOR U10664 ( .A(n9025), .B(n9026), .Z(n9020) );
  ANDN U10665 ( .B(n9027), .A(n9028), .Z(n9025) );
  XNOR U10666 ( .A(b[2458]), .B(n9026), .Z(n9027) );
  XNOR U10667 ( .A(b[2458]), .B(n9028), .Z(c[2458]) );
  XNOR U10668 ( .A(a[2458]), .B(n9029), .Z(n9028) );
  IV U10669 ( .A(n9026), .Z(n9029) );
  XOR U10670 ( .A(n9030), .B(n9031), .Z(n9026) );
  ANDN U10671 ( .B(n9032), .A(n9033), .Z(n9030) );
  XNOR U10672 ( .A(b[2457]), .B(n9031), .Z(n9032) );
  XNOR U10673 ( .A(b[2457]), .B(n9033), .Z(c[2457]) );
  XNOR U10674 ( .A(a[2457]), .B(n9034), .Z(n9033) );
  IV U10675 ( .A(n9031), .Z(n9034) );
  XOR U10676 ( .A(n9035), .B(n9036), .Z(n9031) );
  ANDN U10677 ( .B(n9037), .A(n9038), .Z(n9035) );
  XNOR U10678 ( .A(b[2456]), .B(n9036), .Z(n9037) );
  XNOR U10679 ( .A(b[2456]), .B(n9038), .Z(c[2456]) );
  XNOR U10680 ( .A(a[2456]), .B(n9039), .Z(n9038) );
  IV U10681 ( .A(n9036), .Z(n9039) );
  XOR U10682 ( .A(n9040), .B(n9041), .Z(n9036) );
  ANDN U10683 ( .B(n9042), .A(n9043), .Z(n9040) );
  XNOR U10684 ( .A(b[2455]), .B(n9041), .Z(n9042) );
  XNOR U10685 ( .A(b[2455]), .B(n9043), .Z(c[2455]) );
  XNOR U10686 ( .A(a[2455]), .B(n9044), .Z(n9043) );
  IV U10687 ( .A(n9041), .Z(n9044) );
  XOR U10688 ( .A(n9045), .B(n9046), .Z(n9041) );
  ANDN U10689 ( .B(n9047), .A(n9048), .Z(n9045) );
  XNOR U10690 ( .A(b[2454]), .B(n9046), .Z(n9047) );
  XNOR U10691 ( .A(b[2454]), .B(n9048), .Z(c[2454]) );
  XNOR U10692 ( .A(a[2454]), .B(n9049), .Z(n9048) );
  IV U10693 ( .A(n9046), .Z(n9049) );
  XOR U10694 ( .A(n9050), .B(n9051), .Z(n9046) );
  ANDN U10695 ( .B(n9052), .A(n9053), .Z(n9050) );
  XNOR U10696 ( .A(b[2453]), .B(n9051), .Z(n9052) );
  XNOR U10697 ( .A(b[2453]), .B(n9053), .Z(c[2453]) );
  XNOR U10698 ( .A(a[2453]), .B(n9054), .Z(n9053) );
  IV U10699 ( .A(n9051), .Z(n9054) );
  XOR U10700 ( .A(n9055), .B(n9056), .Z(n9051) );
  ANDN U10701 ( .B(n9057), .A(n9058), .Z(n9055) );
  XNOR U10702 ( .A(b[2452]), .B(n9056), .Z(n9057) );
  XNOR U10703 ( .A(b[2452]), .B(n9058), .Z(c[2452]) );
  XNOR U10704 ( .A(a[2452]), .B(n9059), .Z(n9058) );
  IV U10705 ( .A(n9056), .Z(n9059) );
  XOR U10706 ( .A(n9060), .B(n9061), .Z(n9056) );
  ANDN U10707 ( .B(n9062), .A(n9063), .Z(n9060) );
  XNOR U10708 ( .A(b[2451]), .B(n9061), .Z(n9062) );
  XNOR U10709 ( .A(b[2451]), .B(n9063), .Z(c[2451]) );
  XNOR U10710 ( .A(a[2451]), .B(n9064), .Z(n9063) );
  IV U10711 ( .A(n9061), .Z(n9064) );
  XOR U10712 ( .A(n9065), .B(n9066), .Z(n9061) );
  ANDN U10713 ( .B(n9067), .A(n9068), .Z(n9065) );
  XNOR U10714 ( .A(b[2450]), .B(n9066), .Z(n9067) );
  XNOR U10715 ( .A(b[2450]), .B(n9068), .Z(c[2450]) );
  XNOR U10716 ( .A(a[2450]), .B(n9069), .Z(n9068) );
  IV U10717 ( .A(n9066), .Z(n9069) );
  XOR U10718 ( .A(n9070), .B(n9071), .Z(n9066) );
  ANDN U10719 ( .B(n9072), .A(n9073), .Z(n9070) );
  XNOR U10720 ( .A(b[2449]), .B(n9071), .Z(n9072) );
  XNOR U10721 ( .A(b[244]), .B(n9074), .Z(c[244]) );
  XNOR U10722 ( .A(b[2449]), .B(n9073), .Z(c[2449]) );
  XNOR U10723 ( .A(a[2449]), .B(n9075), .Z(n9073) );
  IV U10724 ( .A(n9071), .Z(n9075) );
  XOR U10725 ( .A(n9076), .B(n9077), .Z(n9071) );
  ANDN U10726 ( .B(n9078), .A(n9079), .Z(n9076) );
  XNOR U10727 ( .A(b[2448]), .B(n9077), .Z(n9078) );
  XNOR U10728 ( .A(b[2448]), .B(n9079), .Z(c[2448]) );
  XNOR U10729 ( .A(a[2448]), .B(n9080), .Z(n9079) );
  IV U10730 ( .A(n9077), .Z(n9080) );
  XOR U10731 ( .A(n9081), .B(n9082), .Z(n9077) );
  ANDN U10732 ( .B(n9083), .A(n9084), .Z(n9081) );
  XNOR U10733 ( .A(b[2447]), .B(n9082), .Z(n9083) );
  XNOR U10734 ( .A(b[2447]), .B(n9084), .Z(c[2447]) );
  XNOR U10735 ( .A(a[2447]), .B(n9085), .Z(n9084) );
  IV U10736 ( .A(n9082), .Z(n9085) );
  XOR U10737 ( .A(n9086), .B(n9087), .Z(n9082) );
  ANDN U10738 ( .B(n9088), .A(n9089), .Z(n9086) );
  XNOR U10739 ( .A(b[2446]), .B(n9087), .Z(n9088) );
  XNOR U10740 ( .A(b[2446]), .B(n9089), .Z(c[2446]) );
  XNOR U10741 ( .A(a[2446]), .B(n9090), .Z(n9089) );
  IV U10742 ( .A(n9087), .Z(n9090) );
  XOR U10743 ( .A(n9091), .B(n9092), .Z(n9087) );
  ANDN U10744 ( .B(n9093), .A(n9094), .Z(n9091) );
  XNOR U10745 ( .A(b[2445]), .B(n9092), .Z(n9093) );
  XNOR U10746 ( .A(b[2445]), .B(n9094), .Z(c[2445]) );
  XNOR U10747 ( .A(a[2445]), .B(n9095), .Z(n9094) );
  IV U10748 ( .A(n9092), .Z(n9095) );
  XOR U10749 ( .A(n9096), .B(n9097), .Z(n9092) );
  ANDN U10750 ( .B(n9098), .A(n9099), .Z(n9096) );
  XNOR U10751 ( .A(b[2444]), .B(n9097), .Z(n9098) );
  XNOR U10752 ( .A(b[2444]), .B(n9099), .Z(c[2444]) );
  XNOR U10753 ( .A(a[2444]), .B(n9100), .Z(n9099) );
  IV U10754 ( .A(n9097), .Z(n9100) );
  XOR U10755 ( .A(n9101), .B(n9102), .Z(n9097) );
  ANDN U10756 ( .B(n9103), .A(n9104), .Z(n9101) );
  XNOR U10757 ( .A(b[2443]), .B(n9102), .Z(n9103) );
  XNOR U10758 ( .A(b[2443]), .B(n9104), .Z(c[2443]) );
  XNOR U10759 ( .A(a[2443]), .B(n9105), .Z(n9104) );
  IV U10760 ( .A(n9102), .Z(n9105) );
  XOR U10761 ( .A(n9106), .B(n9107), .Z(n9102) );
  ANDN U10762 ( .B(n9108), .A(n9109), .Z(n9106) );
  XNOR U10763 ( .A(b[2442]), .B(n9107), .Z(n9108) );
  XNOR U10764 ( .A(b[2442]), .B(n9109), .Z(c[2442]) );
  XNOR U10765 ( .A(a[2442]), .B(n9110), .Z(n9109) );
  IV U10766 ( .A(n9107), .Z(n9110) );
  XOR U10767 ( .A(n9111), .B(n9112), .Z(n9107) );
  ANDN U10768 ( .B(n9113), .A(n9114), .Z(n9111) );
  XNOR U10769 ( .A(b[2441]), .B(n9112), .Z(n9113) );
  XNOR U10770 ( .A(b[2441]), .B(n9114), .Z(c[2441]) );
  XNOR U10771 ( .A(a[2441]), .B(n9115), .Z(n9114) );
  IV U10772 ( .A(n9112), .Z(n9115) );
  XOR U10773 ( .A(n9116), .B(n9117), .Z(n9112) );
  ANDN U10774 ( .B(n9118), .A(n9119), .Z(n9116) );
  XNOR U10775 ( .A(b[2440]), .B(n9117), .Z(n9118) );
  XNOR U10776 ( .A(b[2440]), .B(n9119), .Z(c[2440]) );
  XNOR U10777 ( .A(a[2440]), .B(n9120), .Z(n9119) );
  IV U10778 ( .A(n9117), .Z(n9120) );
  XOR U10779 ( .A(n9121), .B(n9122), .Z(n9117) );
  ANDN U10780 ( .B(n9123), .A(n9124), .Z(n9121) );
  XNOR U10781 ( .A(b[2439]), .B(n9122), .Z(n9123) );
  XNOR U10782 ( .A(b[243]), .B(n9125), .Z(c[243]) );
  XNOR U10783 ( .A(b[2439]), .B(n9124), .Z(c[2439]) );
  XNOR U10784 ( .A(a[2439]), .B(n9126), .Z(n9124) );
  IV U10785 ( .A(n9122), .Z(n9126) );
  XOR U10786 ( .A(n9127), .B(n9128), .Z(n9122) );
  ANDN U10787 ( .B(n9129), .A(n9130), .Z(n9127) );
  XNOR U10788 ( .A(b[2438]), .B(n9128), .Z(n9129) );
  XNOR U10789 ( .A(b[2438]), .B(n9130), .Z(c[2438]) );
  XNOR U10790 ( .A(a[2438]), .B(n9131), .Z(n9130) );
  IV U10791 ( .A(n9128), .Z(n9131) );
  XOR U10792 ( .A(n9132), .B(n9133), .Z(n9128) );
  ANDN U10793 ( .B(n9134), .A(n9135), .Z(n9132) );
  XNOR U10794 ( .A(b[2437]), .B(n9133), .Z(n9134) );
  XNOR U10795 ( .A(b[2437]), .B(n9135), .Z(c[2437]) );
  XNOR U10796 ( .A(a[2437]), .B(n9136), .Z(n9135) );
  IV U10797 ( .A(n9133), .Z(n9136) );
  XOR U10798 ( .A(n9137), .B(n9138), .Z(n9133) );
  ANDN U10799 ( .B(n9139), .A(n9140), .Z(n9137) );
  XNOR U10800 ( .A(b[2436]), .B(n9138), .Z(n9139) );
  XNOR U10801 ( .A(b[2436]), .B(n9140), .Z(c[2436]) );
  XNOR U10802 ( .A(a[2436]), .B(n9141), .Z(n9140) );
  IV U10803 ( .A(n9138), .Z(n9141) );
  XOR U10804 ( .A(n9142), .B(n9143), .Z(n9138) );
  ANDN U10805 ( .B(n9144), .A(n9145), .Z(n9142) );
  XNOR U10806 ( .A(b[2435]), .B(n9143), .Z(n9144) );
  XNOR U10807 ( .A(b[2435]), .B(n9145), .Z(c[2435]) );
  XNOR U10808 ( .A(a[2435]), .B(n9146), .Z(n9145) );
  IV U10809 ( .A(n9143), .Z(n9146) );
  XOR U10810 ( .A(n9147), .B(n9148), .Z(n9143) );
  ANDN U10811 ( .B(n9149), .A(n9150), .Z(n9147) );
  XNOR U10812 ( .A(b[2434]), .B(n9148), .Z(n9149) );
  XNOR U10813 ( .A(b[2434]), .B(n9150), .Z(c[2434]) );
  XNOR U10814 ( .A(a[2434]), .B(n9151), .Z(n9150) );
  IV U10815 ( .A(n9148), .Z(n9151) );
  XOR U10816 ( .A(n9152), .B(n9153), .Z(n9148) );
  ANDN U10817 ( .B(n9154), .A(n9155), .Z(n9152) );
  XNOR U10818 ( .A(b[2433]), .B(n9153), .Z(n9154) );
  XNOR U10819 ( .A(b[2433]), .B(n9155), .Z(c[2433]) );
  XNOR U10820 ( .A(a[2433]), .B(n9156), .Z(n9155) );
  IV U10821 ( .A(n9153), .Z(n9156) );
  XOR U10822 ( .A(n9157), .B(n9158), .Z(n9153) );
  ANDN U10823 ( .B(n9159), .A(n9160), .Z(n9157) );
  XNOR U10824 ( .A(b[2432]), .B(n9158), .Z(n9159) );
  XNOR U10825 ( .A(b[2432]), .B(n9160), .Z(c[2432]) );
  XNOR U10826 ( .A(a[2432]), .B(n9161), .Z(n9160) );
  IV U10827 ( .A(n9158), .Z(n9161) );
  XOR U10828 ( .A(n9162), .B(n9163), .Z(n9158) );
  ANDN U10829 ( .B(n9164), .A(n9165), .Z(n9162) );
  XNOR U10830 ( .A(b[2431]), .B(n9163), .Z(n9164) );
  XNOR U10831 ( .A(b[2431]), .B(n9165), .Z(c[2431]) );
  XNOR U10832 ( .A(a[2431]), .B(n9166), .Z(n9165) );
  IV U10833 ( .A(n9163), .Z(n9166) );
  XOR U10834 ( .A(n9167), .B(n9168), .Z(n9163) );
  ANDN U10835 ( .B(n9169), .A(n9170), .Z(n9167) );
  XNOR U10836 ( .A(b[2430]), .B(n9168), .Z(n9169) );
  XNOR U10837 ( .A(b[2430]), .B(n9170), .Z(c[2430]) );
  XNOR U10838 ( .A(a[2430]), .B(n9171), .Z(n9170) );
  IV U10839 ( .A(n9168), .Z(n9171) );
  XOR U10840 ( .A(n9172), .B(n9173), .Z(n9168) );
  ANDN U10841 ( .B(n9174), .A(n9175), .Z(n9172) );
  XNOR U10842 ( .A(b[2429]), .B(n9173), .Z(n9174) );
  XNOR U10843 ( .A(b[242]), .B(n9176), .Z(c[242]) );
  XNOR U10844 ( .A(b[2429]), .B(n9175), .Z(c[2429]) );
  XNOR U10845 ( .A(a[2429]), .B(n9177), .Z(n9175) );
  IV U10846 ( .A(n9173), .Z(n9177) );
  XOR U10847 ( .A(n9178), .B(n9179), .Z(n9173) );
  ANDN U10848 ( .B(n9180), .A(n9181), .Z(n9178) );
  XNOR U10849 ( .A(b[2428]), .B(n9179), .Z(n9180) );
  XNOR U10850 ( .A(b[2428]), .B(n9181), .Z(c[2428]) );
  XNOR U10851 ( .A(a[2428]), .B(n9182), .Z(n9181) );
  IV U10852 ( .A(n9179), .Z(n9182) );
  XOR U10853 ( .A(n9183), .B(n9184), .Z(n9179) );
  ANDN U10854 ( .B(n9185), .A(n9186), .Z(n9183) );
  XNOR U10855 ( .A(b[2427]), .B(n9184), .Z(n9185) );
  XNOR U10856 ( .A(b[2427]), .B(n9186), .Z(c[2427]) );
  XNOR U10857 ( .A(a[2427]), .B(n9187), .Z(n9186) );
  IV U10858 ( .A(n9184), .Z(n9187) );
  XOR U10859 ( .A(n9188), .B(n9189), .Z(n9184) );
  ANDN U10860 ( .B(n9190), .A(n9191), .Z(n9188) );
  XNOR U10861 ( .A(b[2426]), .B(n9189), .Z(n9190) );
  XNOR U10862 ( .A(b[2426]), .B(n9191), .Z(c[2426]) );
  XNOR U10863 ( .A(a[2426]), .B(n9192), .Z(n9191) );
  IV U10864 ( .A(n9189), .Z(n9192) );
  XOR U10865 ( .A(n9193), .B(n9194), .Z(n9189) );
  ANDN U10866 ( .B(n9195), .A(n9196), .Z(n9193) );
  XNOR U10867 ( .A(b[2425]), .B(n9194), .Z(n9195) );
  XNOR U10868 ( .A(b[2425]), .B(n9196), .Z(c[2425]) );
  XNOR U10869 ( .A(a[2425]), .B(n9197), .Z(n9196) );
  IV U10870 ( .A(n9194), .Z(n9197) );
  XOR U10871 ( .A(n9198), .B(n9199), .Z(n9194) );
  ANDN U10872 ( .B(n9200), .A(n9201), .Z(n9198) );
  XNOR U10873 ( .A(b[2424]), .B(n9199), .Z(n9200) );
  XNOR U10874 ( .A(b[2424]), .B(n9201), .Z(c[2424]) );
  XNOR U10875 ( .A(a[2424]), .B(n9202), .Z(n9201) );
  IV U10876 ( .A(n9199), .Z(n9202) );
  XOR U10877 ( .A(n9203), .B(n9204), .Z(n9199) );
  ANDN U10878 ( .B(n9205), .A(n9206), .Z(n9203) );
  XNOR U10879 ( .A(b[2423]), .B(n9204), .Z(n9205) );
  XNOR U10880 ( .A(b[2423]), .B(n9206), .Z(c[2423]) );
  XNOR U10881 ( .A(a[2423]), .B(n9207), .Z(n9206) );
  IV U10882 ( .A(n9204), .Z(n9207) );
  XOR U10883 ( .A(n9208), .B(n9209), .Z(n9204) );
  ANDN U10884 ( .B(n9210), .A(n9211), .Z(n9208) );
  XNOR U10885 ( .A(b[2422]), .B(n9209), .Z(n9210) );
  XNOR U10886 ( .A(b[2422]), .B(n9211), .Z(c[2422]) );
  XNOR U10887 ( .A(a[2422]), .B(n9212), .Z(n9211) );
  IV U10888 ( .A(n9209), .Z(n9212) );
  XOR U10889 ( .A(n9213), .B(n9214), .Z(n9209) );
  ANDN U10890 ( .B(n9215), .A(n9216), .Z(n9213) );
  XNOR U10891 ( .A(b[2421]), .B(n9214), .Z(n9215) );
  XNOR U10892 ( .A(b[2421]), .B(n9216), .Z(c[2421]) );
  XNOR U10893 ( .A(a[2421]), .B(n9217), .Z(n9216) );
  IV U10894 ( .A(n9214), .Z(n9217) );
  XOR U10895 ( .A(n9218), .B(n9219), .Z(n9214) );
  ANDN U10896 ( .B(n9220), .A(n9221), .Z(n9218) );
  XNOR U10897 ( .A(b[2420]), .B(n9219), .Z(n9220) );
  XNOR U10898 ( .A(b[2420]), .B(n9221), .Z(c[2420]) );
  XNOR U10899 ( .A(a[2420]), .B(n9222), .Z(n9221) );
  IV U10900 ( .A(n9219), .Z(n9222) );
  XOR U10901 ( .A(n9223), .B(n9224), .Z(n9219) );
  ANDN U10902 ( .B(n9225), .A(n9226), .Z(n9223) );
  XNOR U10903 ( .A(b[2419]), .B(n9224), .Z(n9225) );
  XNOR U10904 ( .A(b[241]), .B(n9227), .Z(c[241]) );
  XNOR U10905 ( .A(b[2419]), .B(n9226), .Z(c[2419]) );
  XNOR U10906 ( .A(a[2419]), .B(n9228), .Z(n9226) );
  IV U10907 ( .A(n9224), .Z(n9228) );
  XOR U10908 ( .A(n9229), .B(n9230), .Z(n9224) );
  ANDN U10909 ( .B(n9231), .A(n9232), .Z(n9229) );
  XNOR U10910 ( .A(b[2418]), .B(n9230), .Z(n9231) );
  XNOR U10911 ( .A(b[2418]), .B(n9232), .Z(c[2418]) );
  XNOR U10912 ( .A(a[2418]), .B(n9233), .Z(n9232) );
  IV U10913 ( .A(n9230), .Z(n9233) );
  XOR U10914 ( .A(n9234), .B(n9235), .Z(n9230) );
  ANDN U10915 ( .B(n9236), .A(n9237), .Z(n9234) );
  XNOR U10916 ( .A(b[2417]), .B(n9235), .Z(n9236) );
  XNOR U10917 ( .A(b[2417]), .B(n9237), .Z(c[2417]) );
  XNOR U10918 ( .A(a[2417]), .B(n9238), .Z(n9237) );
  IV U10919 ( .A(n9235), .Z(n9238) );
  XOR U10920 ( .A(n9239), .B(n9240), .Z(n9235) );
  ANDN U10921 ( .B(n9241), .A(n9242), .Z(n9239) );
  XNOR U10922 ( .A(b[2416]), .B(n9240), .Z(n9241) );
  XNOR U10923 ( .A(b[2416]), .B(n9242), .Z(c[2416]) );
  XNOR U10924 ( .A(a[2416]), .B(n9243), .Z(n9242) );
  IV U10925 ( .A(n9240), .Z(n9243) );
  XOR U10926 ( .A(n9244), .B(n9245), .Z(n9240) );
  ANDN U10927 ( .B(n9246), .A(n9247), .Z(n9244) );
  XNOR U10928 ( .A(b[2415]), .B(n9245), .Z(n9246) );
  XNOR U10929 ( .A(b[2415]), .B(n9247), .Z(c[2415]) );
  XNOR U10930 ( .A(a[2415]), .B(n9248), .Z(n9247) );
  IV U10931 ( .A(n9245), .Z(n9248) );
  XOR U10932 ( .A(n9249), .B(n9250), .Z(n9245) );
  ANDN U10933 ( .B(n9251), .A(n9252), .Z(n9249) );
  XNOR U10934 ( .A(b[2414]), .B(n9250), .Z(n9251) );
  XNOR U10935 ( .A(b[2414]), .B(n9252), .Z(c[2414]) );
  XNOR U10936 ( .A(a[2414]), .B(n9253), .Z(n9252) );
  IV U10937 ( .A(n9250), .Z(n9253) );
  XOR U10938 ( .A(n9254), .B(n9255), .Z(n9250) );
  ANDN U10939 ( .B(n9256), .A(n9257), .Z(n9254) );
  XNOR U10940 ( .A(b[2413]), .B(n9255), .Z(n9256) );
  XNOR U10941 ( .A(b[2413]), .B(n9257), .Z(c[2413]) );
  XNOR U10942 ( .A(a[2413]), .B(n9258), .Z(n9257) );
  IV U10943 ( .A(n9255), .Z(n9258) );
  XOR U10944 ( .A(n9259), .B(n9260), .Z(n9255) );
  ANDN U10945 ( .B(n9261), .A(n9262), .Z(n9259) );
  XNOR U10946 ( .A(b[2412]), .B(n9260), .Z(n9261) );
  XNOR U10947 ( .A(b[2412]), .B(n9262), .Z(c[2412]) );
  XNOR U10948 ( .A(a[2412]), .B(n9263), .Z(n9262) );
  IV U10949 ( .A(n9260), .Z(n9263) );
  XOR U10950 ( .A(n9264), .B(n9265), .Z(n9260) );
  ANDN U10951 ( .B(n9266), .A(n9267), .Z(n9264) );
  XNOR U10952 ( .A(b[2411]), .B(n9265), .Z(n9266) );
  XNOR U10953 ( .A(b[2411]), .B(n9267), .Z(c[2411]) );
  XNOR U10954 ( .A(a[2411]), .B(n9268), .Z(n9267) );
  IV U10955 ( .A(n9265), .Z(n9268) );
  XOR U10956 ( .A(n9269), .B(n9270), .Z(n9265) );
  ANDN U10957 ( .B(n9271), .A(n9272), .Z(n9269) );
  XNOR U10958 ( .A(b[2410]), .B(n9270), .Z(n9271) );
  XNOR U10959 ( .A(b[2410]), .B(n9272), .Z(c[2410]) );
  XNOR U10960 ( .A(a[2410]), .B(n9273), .Z(n9272) );
  IV U10961 ( .A(n9270), .Z(n9273) );
  XOR U10962 ( .A(n9274), .B(n9275), .Z(n9270) );
  ANDN U10963 ( .B(n9276), .A(n9277), .Z(n9274) );
  XNOR U10964 ( .A(b[2409]), .B(n9275), .Z(n9276) );
  XNOR U10965 ( .A(b[240]), .B(n9278), .Z(c[240]) );
  XNOR U10966 ( .A(b[2409]), .B(n9277), .Z(c[2409]) );
  XNOR U10967 ( .A(a[2409]), .B(n9279), .Z(n9277) );
  IV U10968 ( .A(n9275), .Z(n9279) );
  XOR U10969 ( .A(n9280), .B(n9281), .Z(n9275) );
  ANDN U10970 ( .B(n9282), .A(n9283), .Z(n9280) );
  XNOR U10971 ( .A(b[2408]), .B(n9281), .Z(n9282) );
  XNOR U10972 ( .A(b[2408]), .B(n9283), .Z(c[2408]) );
  XNOR U10973 ( .A(a[2408]), .B(n9284), .Z(n9283) );
  IV U10974 ( .A(n9281), .Z(n9284) );
  XOR U10975 ( .A(n9285), .B(n9286), .Z(n9281) );
  ANDN U10976 ( .B(n9287), .A(n9288), .Z(n9285) );
  XNOR U10977 ( .A(b[2407]), .B(n9286), .Z(n9287) );
  XNOR U10978 ( .A(b[2407]), .B(n9288), .Z(c[2407]) );
  XNOR U10979 ( .A(a[2407]), .B(n9289), .Z(n9288) );
  IV U10980 ( .A(n9286), .Z(n9289) );
  XOR U10981 ( .A(n9290), .B(n9291), .Z(n9286) );
  ANDN U10982 ( .B(n9292), .A(n9293), .Z(n9290) );
  XNOR U10983 ( .A(b[2406]), .B(n9291), .Z(n9292) );
  XNOR U10984 ( .A(b[2406]), .B(n9293), .Z(c[2406]) );
  XNOR U10985 ( .A(a[2406]), .B(n9294), .Z(n9293) );
  IV U10986 ( .A(n9291), .Z(n9294) );
  XOR U10987 ( .A(n9295), .B(n9296), .Z(n9291) );
  ANDN U10988 ( .B(n9297), .A(n9298), .Z(n9295) );
  XNOR U10989 ( .A(b[2405]), .B(n9296), .Z(n9297) );
  XNOR U10990 ( .A(b[2405]), .B(n9298), .Z(c[2405]) );
  XNOR U10991 ( .A(a[2405]), .B(n9299), .Z(n9298) );
  IV U10992 ( .A(n9296), .Z(n9299) );
  XOR U10993 ( .A(n9300), .B(n9301), .Z(n9296) );
  ANDN U10994 ( .B(n9302), .A(n9303), .Z(n9300) );
  XNOR U10995 ( .A(b[2404]), .B(n9301), .Z(n9302) );
  XNOR U10996 ( .A(b[2404]), .B(n9303), .Z(c[2404]) );
  XNOR U10997 ( .A(a[2404]), .B(n9304), .Z(n9303) );
  IV U10998 ( .A(n9301), .Z(n9304) );
  XOR U10999 ( .A(n9305), .B(n9306), .Z(n9301) );
  ANDN U11000 ( .B(n9307), .A(n9308), .Z(n9305) );
  XNOR U11001 ( .A(b[2403]), .B(n9306), .Z(n9307) );
  XNOR U11002 ( .A(b[2403]), .B(n9308), .Z(c[2403]) );
  XNOR U11003 ( .A(a[2403]), .B(n9309), .Z(n9308) );
  IV U11004 ( .A(n9306), .Z(n9309) );
  XOR U11005 ( .A(n9310), .B(n9311), .Z(n9306) );
  ANDN U11006 ( .B(n9312), .A(n9313), .Z(n9310) );
  XNOR U11007 ( .A(b[2402]), .B(n9311), .Z(n9312) );
  XNOR U11008 ( .A(b[2402]), .B(n9313), .Z(c[2402]) );
  XNOR U11009 ( .A(a[2402]), .B(n9314), .Z(n9313) );
  IV U11010 ( .A(n9311), .Z(n9314) );
  XOR U11011 ( .A(n9315), .B(n9316), .Z(n9311) );
  ANDN U11012 ( .B(n9317), .A(n9318), .Z(n9315) );
  XNOR U11013 ( .A(b[2401]), .B(n9316), .Z(n9317) );
  XNOR U11014 ( .A(b[2401]), .B(n9318), .Z(c[2401]) );
  XNOR U11015 ( .A(a[2401]), .B(n9319), .Z(n9318) );
  IV U11016 ( .A(n9316), .Z(n9319) );
  XOR U11017 ( .A(n9320), .B(n9321), .Z(n9316) );
  ANDN U11018 ( .B(n9322), .A(n9323), .Z(n9320) );
  XNOR U11019 ( .A(b[2400]), .B(n9321), .Z(n9322) );
  XNOR U11020 ( .A(b[2400]), .B(n9323), .Z(c[2400]) );
  XNOR U11021 ( .A(a[2400]), .B(n9324), .Z(n9323) );
  IV U11022 ( .A(n9321), .Z(n9324) );
  XOR U11023 ( .A(n9325), .B(n9326), .Z(n9321) );
  ANDN U11024 ( .B(n9327), .A(n9328), .Z(n9325) );
  XNOR U11025 ( .A(b[2399]), .B(n9326), .Z(n9327) );
  XNOR U11026 ( .A(b[23]), .B(n9329), .Z(c[23]) );
  XNOR U11027 ( .A(b[239]), .B(n9330), .Z(c[239]) );
  XNOR U11028 ( .A(b[2399]), .B(n9328), .Z(c[2399]) );
  XNOR U11029 ( .A(a[2399]), .B(n9331), .Z(n9328) );
  IV U11030 ( .A(n9326), .Z(n9331) );
  XOR U11031 ( .A(n9332), .B(n9333), .Z(n9326) );
  ANDN U11032 ( .B(n9334), .A(n9335), .Z(n9332) );
  XNOR U11033 ( .A(b[2398]), .B(n9333), .Z(n9334) );
  XNOR U11034 ( .A(b[2398]), .B(n9335), .Z(c[2398]) );
  XNOR U11035 ( .A(a[2398]), .B(n9336), .Z(n9335) );
  IV U11036 ( .A(n9333), .Z(n9336) );
  XOR U11037 ( .A(n9337), .B(n9338), .Z(n9333) );
  ANDN U11038 ( .B(n9339), .A(n9340), .Z(n9337) );
  XNOR U11039 ( .A(b[2397]), .B(n9338), .Z(n9339) );
  XNOR U11040 ( .A(b[2397]), .B(n9340), .Z(c[2397]) );
  XNOR U11041 ( .A(a[2397]), .B(n9341), .Z(n9340) );
  IV U11042 ( .A(n9338), .Z(n9341) );
  XOR U11043 ( .A(n9342), .B(n9343), .Z(n9338) );
  ANDN U11044 ( .B(n9344), .A(n9345), .Z(n9342) );
  XNOR U11045 ( .A(b[2396]), .B(n9343), .Z(n9344) );
  XNOR U11046 ( .A(b[2396]), .B(n9345), .Z(c[2396]) );
  XNOR U11047 ( .A(a[2396]), .B(n9346), .Z(n9345) );
  IV U11048 ( .A(n9343), .Z(n9346) );
  XOR U11049 ( .A(n9347), .B(n9348), .Z(n9343) );
  ANDN U11050 ( .B(n9349), .A(n9350), .Z(n9347) );
  XNOR U11051 ( .A(b[2395]), .B(n9348), .Z(n9349) );
  XNOR U11052 ( .A(b[2395]), .B(n9350), .Z(c[2395]) );
  XNOR U11053 ( .A(a[2395]), .B(n9351), .Z(n9350) );
  IV U11054 ( .A(n9348), .Z(n9351) );
  XOR U11055 ( .A(n9352), .B(n9353), .Z(n9348) );
  ANDN U11056 ( .B(n9354), .A(n9355), .Z(n9352) );
  XNOR U11057 ( .A(b[2394]), .B(n9353), .Z(n9354) );
  XNOR U11058 ( .A(b[2394]), .B(n9355), .Z(c[2394]) );
  XNOR U11059 ( .A(a[2394]), .B(n9356), .Z(n9355) );
  IV U11060 ( .A(n9353), .Z(n9356) );
  XOR U11061 ( .A(n9357), .B(n9358), .Z(n9353) );
  ANDN U11062 ( .B(n9359), .A(n9360), .Z(n9357) );
  XNOR U11063 ( .A(b[2393]), .B(n9358), .Z(n9359) );
  XNOR U11064 ( .A(b[2393]), .B(n9360), .Z(c[2393]) );
  XNOR U11065 ( .A(a[2393]), .B(n9361), .Z(n9360) );
  IV U11066 ( .A(n9358), .Z(n9361) );
  XOR U11067 ( .A(n9362), .B(n9363), .Z(n9358) );
  ANDN U11068 ( .B(n9364), .A(n9365), .Z(n9362) );
  XNOR U11069 ( .A(b[2392]), .B(n9363), .Z(n9364) );
  XNOR U11070 ( .A(b[2392]), .B(n9365), .Z(c[2392]) );
  XNOR U11071 ( .A(a[2392]), .B(n9366), .Z(n9365) );
  IV U11072 ( .A(n9363), .Z(n9366) );
  XOR U11073 ( .A(n9367), .B(n9368), .Z(n9363) );
  ANDN U11074 ( .B(n9369), .A(n9370), .Z(n9367) );
  XNOR U11075 ( .A(b[2391]), .B(n9368), .Z(n9369) );
  XNOR U11076 ( .A(b[2391]), .B(n9370), .Z(c[2391]) );
  XNOR U11077 ( .A(a[2391]), .B(n9371), .Z(n9370) );
  IV U11078 ( .A(n9368), .Z(n9371) );
  XOR U11079 ( .A(n9372), .B(n9373), .Z(n9368) );
  ANDN U11080 ( .B(n9374), .A(n9375), .Z(n9372) );
  XNOR U11081 ( .A(b[2390]), .B(n9373), .Z(n9374) );
  XNOR U11082 ( .A(b[2390]), .B(n9375), .Z(c[2390]) );
  XNOR U11083 ( .A(a[2390]), .B(n9376), .Z(n9375) );
  IV U11084 ( .A(n9373), .Z(n9376) );
  XOR U11085 ( .A(n9377), .B(n9378), .Z(n9373) );
  ANDN U11086 ( .B(n9379), .A(n9380), .Z(n9377) );
  XNOR U11087 ( .A(b[2389]), .B(n9378), .Z(n9379) );
  XNOR U11088 ( .A(b[238]), .B(n9381), .Z(c[238]) );
  XNOR U11089 ( .A(b[2389]), .B(n9380), .Z(c[2389]) );
  XNOR U11090 ( .A(a[2389]), .B(n9382), .Z(n9380) );
  IV U11091 ( .A(n9378), .Z(n9382) );
  XOR U11092 ( .A(n9383), .B(n9384), .Z(n9378) );
  ANDN U11093 ( .B(n9385), .A(n9386), .Z(n9383) );
  XNOR U11094 ( .A(b[2388]), .B(n9384), .Z(n9385) );
  XNOR U11095 ( .A(b[2388]), .B(n9386), .Z(c[2388]) );
  XNOR U11096 ( .A(a[2388]), .B(n9387), .Z(n9386) );
  IV U11097 ( .A(n9384), .Z(n9387) );
  XOR U11098 ( .A(n9388), .B(n9389), .Z(n9384) );
  ANDN U11099 ( .B(n9390), .A(n9391), .Z(n9388) );
  XNOR U11100 ( .A(b[2387]), .B(n9389), .Z(n9390) );
  XNOR U11101 ( .A(b[2387]), .B(n9391), .Z(c[2387]) );
  XNOR U11102 ( .A(a[2387]), .B(n9392), .Z(n9391) );
  IV U11103 ( .A(n9389), .Z(n9392) );
  XOR U11104 ( .A(n9393), .B(n9394), .Z(n9389) );
  ANDN U11105 ( .B(n9395), .A(n9396), .Z(n9393) );
  XNOR U11106 ( .A(b[2386]), .B(n9394), .Z(n9395) );
  XNOR U11107 ( .A(b[2386]), .B(n9396), .Z(c[2386]) );
  XNOR U11108 ( .A(a[2386]), .B(n9397), .Z(n9396) );
  IV U11109 ( .A(n9394), .Z(n9397) );
  XOR U11110 ( .A(n9398), .B(n9399), .Z(n9394) );
  ANDN U11111 ( .B(n9400), .A(n9401), .Z(n9398) );
  XNOR U11112 ( .A(b[2385]), .B(n9399), .Z(n9400) );
  XNOR U11113 ( .A(b[2385]), .B(n9401), .Z(c[2385]) );
  XNOR U11114 ( .A(a[2385]), .B(n9402), .Z(n9401) );
  IV U11115 ( .A(n9399), .Z(n9402) );
  XOR U11116 ( .A(n9403), .B(n9404), .Z(n9399) );
  ANDN U11117 ( .B(n9405), .A(n9406), .Z(n9403) );
  XNOR U11118 ( .A(b[2384]), .B(n9404), .Z(n9405) );
  XNOR U11119 ( .A(b[2384]), .B(n9406), .Z(c[2384]) );
  XNOR U11120 ( .A(a[2384]), .B(n9407), .Z(n9406) );
  IV U11121 ( .A(n9404), .Z(n9407) );
  XOR U11122 ( .A(n9408), .B(n9409), .Z(n9404) );
  ANDN U11123 ( .B(n9410), .A(n9411), .Z(n9408) );
  XNOR U11124 ( .A(b[2383]), .B(n9409), .Z(n9410) );
  XNOR U11125 ( .A(b[2383]), .B(n9411), .Z(c[2383]) );
  XNOR U11126 ( .A(a[2383]), .B(n9412), .Z(n9411) );
  IV U11127 ( .A(n9409), .Z(n9412) );
  XOR U11128 ( .A(n9413), .B(n9414), .Z(n9409) );
  ANDN U11129 ( .B(n9415), .A(n9416), .Z(n9413) );
  XNOR U11130 ( .A(b[2382]), .B(n9414), .Z(n9415) );
  XNOR U11131 ( .A(b[2382]), .B(n9416), .Z(c[2382]) );
  XNOR U11132 ( .A(a[2382]), .B(n9417), .Z(n9416) );
  IV U11133 ( .A(n9414), .Z(n9417) );
  XOR U11134 ( .A(n9418), .B(n9419), .Z(n9414) );
  ANDN U11135 ( .B(n9420), .A(n9421), .Z(n9418) );
  XNOR U11136 ( .A(b[2381]), .B(n9419), .Z(n9420) );
  XNOR U11137 ( .A(b[2381]), .B(n9421), .Z(c[2381]) );
  XNOR U11138 ( .A(a[2381]), .B(n9422), .Z(n9421) );
  IV U11139 ( .A(n9419), .Z(n9422) );
  XOR U11140 ( .A(n9423), .B(n9424), .Z(n9419) );
  ANDN U11141 ( .B(n9425), .A(n9426), .Z(n9423) );
  XNOR U11142 ( .A(b[2380]), .B(n9424), .Z(n9425) );
  XNOR U11143 ( .A(b[2380]), .B(n9426), .Z(c[2380]) );
  XNOR U11144 ( .A(a[2380]), .B(n9427), .Z(n9426) );
  IV U11145 ( .A(n9424), .Z(n9427) );
  XOR U11146 ( .A(n9428), .B(n9429), .Z(n9424) );
  ANDN U11147 ( .B(n9430), .A(n9431), .Z(n9428) );
  XNOR U11148 ( .A(b[2379]), .B(n9429), .Z(n9430) );
  XNOR U11149 ( .A(b[237]), .B(n9432), .Z(c[237]) );
  XNOR U11150 ( .A(b[2379]), .B(n9431), .Z(c[2379]) );
  XNOR U11151 ( .A(a[2379]), .B(n9433), .Z(n9431) );
  IV U11152 ( .A(n9429), .Z(n9433) );
  XOR U11153 ( .A(n9434), .B(n9435), .Z(n9429) );
  ANDN U11154 ( .B(n9436), .A(n9437), .Z(n9434) );
  XNOR U11155 ( .A(b[2378]), .B(n9435), .Z(n9436) );
  XNOR U11156 ( .A(b[2378]), .B(n9437), .Z(c[2378]) );
  XNOR U11157 ( .A(a[2378]), .B(n9438), .Z(n9437) );
  IV U11158 ( .A(n9435), .Z(n9438) );
  XOR U11159 ( .A(n9439), .B(n9440), .Z(n9435) );
  ANDN U11160 ( .B(n9441), .A(n9442), .Z(n9439) );
  XNOR U11161 ( .A(b[2377]), .B(n9440), .Z(n9441) );
  XNOR U11162 ( .A(b[2377]), .B(n9442), .Z(c[2377]) );
  XNOR U11163 ( .A(a[2377]), .B(n9443), .Z(n9442) );
  IV U11164 ( .A(n9440), .Z(n9443) );
  XOR U11165 ( .A(n9444), .B(n9445), .Z(n9440) );
  ANDN U11166 ( .B(n9446), .A(n9447), .Z(n9444) );
  XNOR U11167 ( .A(b[2376]), .B(n9445), .Z(n9446) );
  XNOR U11168 ( .A(b[2376]), .B(n9447), .Z(c[2376]) );
  XNOR U11169 ( .A(a[2376]), .B(n9448), .Z(n9447) );
  IV U11170 ( .A(n9445), .Z(n9448) );
  XOR U11171 ( .A(n9449), .B(n9450), .Z(n9445) );
  ANDN U11172 ( .B(n9451), .A(n9452), .Z(n9449) );
  XNOR U11173 ( .A(b[2375]), .B(n9450), .Z(n9451) );
  XNOR U11174 ( .A(b[2375]), .B(n9452), .Z(c[2375]) );
  XNOR U11175 ( .A(a[2375]), .B(n9453), .Z(n9452) );
  IV U11176 ( .A(n9450), .Z(n9453) );
  XOR U11177 ( .A(n9454), .B(n9455), .Z(n9450) );
  ANDN U11178 ( .B(n9456), .A(n9457), .Z(n9454) );
  XNOR U11179 ( .A(b[2374]), .B(n9455), .Z(n9456) );
  XNOR U11180 ( .A(b[2374]), .B(n9457), .Z(c[2374]) );
  XNOR U11181 ( .A(a[2374]), .B(n9458), .Z(n9457) );
  IV U11182 ( .A(n9455), .Z(n9458) );
  XOR U11183 ( .A(n9459), .B(n9460), .Z(n9455) );
  ANDN U11184 ( .B(n9461), .A(n9462), .Z(n9459) );
  XNOR U11185 ( .A(b[2373]), .B(n9460), .Z(n9461) );
  XNOR U11186 ( .A(b[2373]), .B(n9462), .Z(c[2373]) );
  XNOR U11187 ( .A(a[2373]), .B(n9463), .Z(n9462) );
  IV U11188 ( .A(n9460), .Z(n9463) );
  XOR U11189 ( .A(n9464), .B(n9465), .Z(n9460) );
  ANDN U11190 ( .B(n9466), .A(n9467), .Z(n9464) );
  XNOR U11191 ( .A(b[2372]), .B(n9465), .Z(n9466) );
  XNOR U11192 ( .A(b[2372]), .B(n9467), .Z(c[2372]) );
  XNOR U11193 ( .A(a[2372]), .B(n9468), .Z(n9467) );
  IV U11194 ( .A(n9465), .Z(n9468) );
  XOR U11195 ( .A(n9469), .B(n9470), .Z(n9465) );
  ANDN U11196 ( .B(n9471), .A(n9472), .Z(n9469) );
  XNOR U11197 ( .A(b[2371]), .B(n9470), .Z(n9471) );
  XNOR U11198 ( .A(b[2371]), .B(n9472), .Z(c[2371]) );
  XNOR U11199 ( .A(a[2371]), .B(n9473), .Z(n9472) );
  IV U11200 ( .A(n9470), .Z(n9473) );
  XOR U11201 ( .A(n9474), .B(n9475), .Z(n9470) );
  ANDN U11202 ( .B(n9476), .A(n9477), .Z(n9474) );
  XNOR U11203 ( .A(b[2370]), .B(n9475), .Z(n9476) );
  XNOR U11204 ( .A(b[2370]), .B(n9477), .Z(c[2370]) );
  XNOR U11205 ( .A(a[2370]), .B(n9478), .Z(n9477) );
  IV U11206 ( .A(n9475), .Z(n9478) );
  XOR U11207 ( .A(n9479), .B(n9480), .Z(n9475) );
  ANDN U11208 ( .B(n9481), .A(n9482), .Z(n9479) );
  XNOR U11209 ( .A(b[2369]), .B(n9480), .Z(n9481) );
  XNOR U11210 ( .A(b[236]), .B(n9483), .Z(c[236]) );
  XNOR U11211 ( .A(b[2369]), .B(n9482), .Z(c[2369]) );
  XNOR U11212 ( .A(a[2369]), .B(n9484), .Z(n9482) );
  IV U11213 ( .A(n9480), .Z(n9484) );
  XOR U11214 ( .A(n9485), .B(n9486), .Z(n9480) );
  ANDN U11215 ( .B(n9487), .A(n9488), .Z(n9485) );
  XNOR U11216 ( .A(b[2368]), .B(n9486), .Z(n9487) );
  XNOR U11217 ( .A(b[2368]), .B(n9488), .Z(c[2368]) );
  XNOR U11218 ( .A(a[2368]), .B(n9489), .Z(n9488) );
  IV U11219 ( .A(n9486), .Z(n9489) );
  XOR U11220 ( .A(n9490), .B(n9491), .Z(n9486) );
  ANDN U11221 ( .B(n9492), .A(n9493), .Z(n9490) );
  XNOR U11222 ( .A(b[2367]), .B(n9491), .Z(n9492) );
  XNOR U11223 ( .A(b[2367]), .B(n9493), .Z(c[2367]) );
  XNOR U11224 ( .A(a[2367]), .B(n9494), .Z(n9493) );
  IV U11225 ( .A(n9491), .Z(n9494) );
  XOR U11226 ( .A(n9495), .B(n9496), .Z(n9491) );
  ANDN U11227 ( .B(n9497), .A(n9498), .Z(n9495) );
  XNOR U11228 ( .A(b[2366]), .B(n9496), .Z(n9497) );
  XNOR U11229 ( .A(b[2366]), .B(n9498), .Z(c[2366]) );
  XNOR U11230 ( .A(a[2366]), .B(n9499), .Z(n9498) );
  IV U11231 ( .A(n9496), .Z(n9499) );
  XOR U11232 ( .A(n9500), .B(n9501), .Z(n9496) );
  ANDN U11233 ( .B(n9502), .A(n9503), .Z(n9500) );
  XNOR U11234 ( .A(b[2365]), .B(n9501), .Z(n9502) );
  XNOR U11235 ( .A(b[2365]), .B(n9503), .Z(c[2365]) );
  XNOR U11236 ( .A(a[2365]), .B(n9504), .Z(n9503) );
  IV U11237 ( .A(n9501), .Z(n9504) );
  XOR U11238 ( .A(n9505), .B(n9506), .Z(n9501) );
  ANDN U11239 ( .B(n9507), .A(n9508), .Z(n9505) );
  XNOR U11240 ( .A(b[2364]), .B(n9506), .Z(n9507) );
  XNOR U11241 ( .A(b[2364]), .B(n9508), .Z(c[2364]) );
  XNOR U11242 ( .A(a[2364]), .B(n9509), .Z(n9508) );
  IV U11243 ( .A(n9506), .Z(n9509) );
  XOR U11244 ( .A(n9510), .B(n9511), .Z(n9506) );
  ANDN U11245 ( .B(n9512), .A(n9513), .Z(n9510) );
  XNOR U11246 ( .A(b[2363]), .B(n9511), .Z(n9512) );
  XNOR U11247 ( .A(b[2363]), .B(n9513), .Z(c[2363]) );
  XNOR U11248 ( .A(a[2363]), .B(n9514), .Z(n9513) );
  IV U11249 ( .A(n9511), .Z(n9514) );
  XOR U11250 ( .A(n9515), .B(n9516), .Z(n9511) );
  ANDN U11251 ( .B(n9517), .A(n9518), .Z(n9515) );
  XNOR U11252 ( .A(b[2362]), .B(n9516), .Z(n9517) );
  XNOR U11253 ( .A(b[2362]), .B(n9518), .Z(c[2362]) );
  XNOR U11254 ( .A(a[2362]), .B(n9519), .Z(n9518) );
  IV U11255 ( .A(n9516), .Z(n9519) );
  XOR U11256 ( .A(n9520), .B(n9521), .Z(n9516) );
  ANDN U11257 ( .B(n9522), .A(n9523), .Z(n9520) );
  XNOR U11258 ( .A(b[2361]), .B(n9521), .Z(n9522) );
  XNOR U11259 ( .A(b[2361]), .B(n9523), .Z(c[2361]) );
  XNOR U11260 ( .A(a[2361]), .B(n9524), .Z(n9523) );
  IV U11261 ( .A(n9521), .Z(n9524) );
  XOR U11262 ( .A(n9525), .B(n9526), .Z(n9521) );
  ANDN U11263 ( .B(n9527), .A(n9528), .Z(n9525) );
  XNOR U11264 ( .A(b[2360]), .B(n9526), .Z(n9527) );
  XNOR U11265 ( .A(b[2360]), .B(n9528), .Z(c[2360]) );
  XNOR U11266 ( .A(a[2360]), .B(n9529), .Z(n9528) );
  IV U11267 ( .A(n9526), .Z(n9529) );
  XOR U11268 ( .A(n9530), .B(n9531), .Z(n9526) );
  ANDN U11269 ( .B(n9532), .A(n9533), .Z(n9530) );
  XNOR U11270 ( .A(b[2359]), .B(n9531), .Z(n9532) );
  XNOR U11271 ( .A(b[235]), .B(n9534), .Z(c[235]) );
  XNOR U11272 ( .A(b[2359]), .B(n9533), .Z(c[2359]) );
  XNOR U11273 ( .A(a[2359]), .B(n9535), .Z(n9533) );
  IV U11274 ( .A(n9531), .Z(n9535) );
  XOR U11275 ( .A(n9536), .B(n9537), .Z(n9531) );
  ANDN U11276 ( .B(n9538), .A(n9539), .Z(n9536) );
  XNOR U11277 ( .A(b[2358]), .B(n9537), .Z(n9538) );
  XNOR U11278 ( .A(b[2358]), .B(n9539), .Z(c[2358]) );
  XNOR U11279 ( .A(a[2358]), .B(n9540), .Z(n9539) );
  IV U11280 ( .A(n9537), .Z(n9540) );
  XOR U11281 ( .A(n9541), .B(n9542), .Z(n9537) );
  ANDN U11282 ( .B(n9543), .A(n9544), .Z(n9541) );
  XNOR U11283 ( .A(b[2357]), .B(n9542), .Z(n9543) );
  XNOR U11284 ( .A(b[2357]), .B(n9544), .Z(c[2357]) );
  XNOR U11285 ( .A(a[2357]), .B(n9545), .Z(n9544) );
  IV U11286 ( .A(n9542), .Z(n9545) );
  XOR U11287 ( .A(n9546), .B(n9547), .Z(n9542) );
  ANDN U11288 ( .B(n9548), .A(n9549), .Z(n9546) );
  XNOR U11289 ( .A(b[2356]), .B(n9547), .Z(n9548) );
  XNOR U11290 ( .A(b[2356]), .B(n9549), .Z(c[2356]) );
  XNOR U11291 ( .A(a[2356]), .B(n9550), .Z(n9549) );
  IV U11292 ( .A(n9547), .Z(n9550) );
  XOR U11293 ( .A(n9551), .B(n9552), .Z(n9547) );
  ANDN U11294 ( .B(n9553), .A(n9554), .Z(n9551) );
  XNOR U11295 ( .A(b[2355]), .B(n9552), .Z(n9553) );
  XNOR U11296 ( .A(b[2355]), .B(n9554), .Z(c[2355]) );
  XNOR U11297 ( .A(a[2355]), .B(n9555), .Z(n9554) );
  IV U11298 ( .A(n9552), .Z(n9555) );
  XOR U11299 ( .A(n9556), .B(n9557), .Z(n9552) );
  ANDN U11300 ( .B(n9558), .A(n9559), .Z(n9556) );
  XNOR U11301 ( .A(b[2354]), .B(n9557), .Z(n9558) );
  XNOR U11302 ( .A(b[2354]), .B(n9559), .Z(c[2354]) );
  XNOR U11303 ( .A(a[2354]), .B(n9560), .Z(n9559) );
  IV U11304 ( .A(n9557), .Z(n9560) );
  XOR U11305 ( .A(n9561), .B(n9562), .Z(n9557) );
  ANDN U11306 ( .B(n9563), .A(n9564), .Z(n9561) );
  XNOR U11307 ( .A(b[2353]), .B(n9562), .Z(n9563) );
  XNOR U11308 ( .A(b[2353]), .B(n9564), .Z(c[2353]) );
  XNOR U11309 ( .A(a[2353]), .B(n9565), .Z(n9564) );
  IV U11310 ( .A(n9562), .Z(n9565) );
  XOR U11311 ( .A(n9566), .B(n9567), .Z(n9562) );
  ANDN U11312 ( .B(n9568), .A(n9569), .Z(n9566) );
  XNOR U11313 ( .A(b[2352]), .B(n9567), .Z(n9568) );
  XNOR U11314 ( .A(b[2352]), .B(n9569), .Z(c[2352]) );
  XNOR U11315 ( .A(a[2352]), .B(n9570), .Z(n9569) );
  IV U11316 ( .A(n9567), .Z(n9570) );
  XOR U11317 ( .A(n9571), .B(n9572), .Z(n9567) );
  ANDN U11318 ( .B(n9573), .A(n9574), .Z(n9571) );
  XNOR U11319 ( .A(b[2351]), .B(n9572), .Z(n9573) );
  XNOR U11320 ( .A(b[2351]), .B(n9574), .Z(c[2351]) );
  XNOR U11321 ( .A(a[2351]), .B(n9575), .Z(n9574) );
  IV U11322 ( .A(n9572), .Z(n9575) );
  XOR U11323 ( .A(n9576), .B(n9577), .Z(n9572) );
  ANDN U11324 ( .B(n9578), .A(n9579), .Z(n9576) );
  XNOR U11325 ( .A(b[2350]), .B(n9577), .Z(n9578) );
  XNOR U11326 ( .A(b[2350]), .B(n9579), .Z(c[2350]) );
  XNOR U11327 ( .A(a[2350]), .B(n9580), .Z(n9579) );
  IV U11328 ( .A(n9577), .Z(n9580) );
  XOR U11329 ( .A(n9581), .B(n9582), .Z(n9577) );
  ANDN U11330 ( .B(n9583), .A(n9584), .Z(n9581) );
  XNOR U11331 ( .A(b[2349]), .B(n9582), .Z(n9583) );
  XNOR U11332 ( .A(b[234]), .B(n9585), .Z(c[234]) );
  XNOR U11333 ( .A(b[2349]), .B(n9584), .Z(c[2349]) );
  XNOR U11334 ( .A(a[2349]), .B(n9586), .Z(n9584) );
  IV U11335 ( .A(n9582), .Z(n9586) );
  XOR U11336 ( .A(n9587), .B(n9588), .Z(n9582) );
  ANDN U11337 ( .B(n9589), .A(n9590), .Z(n9587) );
  XNOR U11338 ( .A(b[2348]), .B(n9588), .Z(n9589) );
  XNOR U11339 ( .A(b[2348]), .B(n9590), .Z(c[2348]) );
  XNOR U11340 ( .A(a[2348]), .B(n9591), .Z(n9590) );
  IV U11341 ( .A(n9588), .Z(n9591) );
  XOR U11342 ( .A(n9592), .B(n9593), .Z(n9588) );
  ANDN U11343 ( .B(n9594), .A(n9595), .Z(n9592) );
  XNOR U11344 ( .A(b[2347]), .B(n9593), .Z(n9594) );
  XNOR U11345 ( .A(b[2347]), .B(n9595), .Z(c[2347]) );
  XNOR U11346 ( .A(a[2347]), .B(n9596), .Z(n9595) );
  IV U11347 ( .A(n9593), .Z(n9596) );
  XOR U11348 ( .A(n9597), .B(n9598), .Z(n9593) );
  ANDN U11349 ( .B(n9599), .A(n9600), .Z(n9597) );
  XNOR U11350 ( .A(b[2346]), .B(n9598), .Z(n9599) );
  XNOR U11351 ( .A(b[2346]), .B(n9600), .Z(c[2346]) );
  XNOR U11352 ( .A(a[2346]), .B(n9601), .Z(n9600) );
  IV U11353 ( .A(n9598), .Z(n9601) );
  XOR U11354 ( .A(n9602), .B(n9603), .Z(n9598) );
  ANDN U11355 ( .B(n9604), .A(n9605), .Z(n9602) );
  XNOR U11356 ( .A(b[2345]), .B(n9603), .Z(n9604) );
  XNOR U11357 ( .A(b[2345]), .B(n9605), .Z(c[2345]) );
  XNOR U11358 ( .A(a[2345]), .B(n9606), .Z(n9605) );
  IV U11359 ( .A(n9603), .Z(n9606) );
  XOR U11360 ( .A(n9607), .B(n9608), .Z(n9603) );
  ANDN U11361 ( .B(n9609), .A(n9610), .Z(n9607) );
  XNOR U11362 ( .A(b[2344]), .B(n9608), .Z(n9609) );
  XNOR U11363 ( .A(b[2344]), .B(n9610), .Z(c[2344]) );
  XNOR U11364 ( .A(a[2344]), .B(n9611), .Z(n9610) );
  IV U11365 ( .A(n9608), .Z(n9611) );
  XOR U11366 ( .A(n9612), .B(n9613), .Z(n9608) );
  ANDN U11367 ( .B(n9614), .A(n9615), .Z(n9612) );
  XNOR U11368 ( .A(b[2343]), .B(n9613), .Z(n9614) );
  XNOR U11369 ( .A(b[2343]), .B(n9615), .Z(c[2343]) );
  XNOR U11370 ( .A(a[2343]), .B(n9616), .Z(n9615) );
  IV U11371 ( .A(n9613), .Z(n9616) );
  XOR U11372 ( .A(n9617), .B(n9618), .Z(n9613) );
  ANDN U11373 ( .B(n9619), .A(n9620), .Z(n9617) );
  XNOR U11374 ( .A(b[2342]), .B(n9618), .Z(n9619) );
  XNOR U11375 ( .A(b[2342]), .B(n9620), .Z(c[2342]) );
  XNOR U11376 ( .A(a[2342]), .B(n9621), .Z(n9620) );
  IV U11377 ( .A(n9618), .Z(n9621) );
  XOR U11378 ( .A(n9622), .B(n9623), .Z(n9618) );
  ANDN U11379 ( .B(n9624), .A(n9625), .Z(n9622) );
  XNOR U11380 ( .A(b[2341]), .B(n9623), .Z(n9624) );
  XNOR U11381 ( .A(b[2341]), .B(n9625), .Z(c[2341]) );
  XNOR U11382 ( .A(a[2341]), .B(n9626), .Z(n9625) );
  IV U11383 ( .A(n9623), .Z(n9626) );
  XOR U11384 ( .A(n9627), .B(n9628), .Z(n9623) );
  ANDN U11385 ( .B(n9629), .A(n9630), .Z(n9627) );
  XNOR U11386 ( .A(b[2340]), .B(n9628), .Z(n9629) );
  XNOR U11387 ( .A(b[2340]), .B(n9630), .Z(c[2340]) );
  XNOR U11388 ( .A(a[2340]), .B(n9631), .Z(n9630) );
  IV U11389 ( .A(n9628), .Z(n9631) );
  XOR U11390 ( .A(n9632), .B(n9633), .Z(n9628) );
  ANDN U11391 ( .B(n9634), .A(n9635), .Z(n9632) );
  XNOR U11392 ( .A(b[2339]), .B(n9633), .Z(n9634) );
  XNOR U11393 ( .A(b[233]), .B(n9636), .Z(c[233]) );
  XNOR U11394 ( .A(b[2339]), .B(n9635), .Z(c[2339]) );
  XNOR U11395 ( .A(a[2339]), .B(n9637), .Z(n9635) );
  IV U11396 ( .A(n9633), .Z(n9637) );
  XOR U11397 ( .A(n9638), .B(n9639), .Z(n9633) );
  ANDN U11398 ( .B(n9640), .A(n9641), .Z(n9638) );
  XNOR U11399 ( .A(b[2338]), .B(n9639), .Z(n9640) );
  XNOR U11400 ( .A(b[2338]), .B(n9641), .Z(c[2338]) );
  XNOR U11401 ( .A(a[2338]), .B(n9642), .Z(n9641) );
  IV U11402 ( .A(n9639), .Z(n9642) );
  XOR U11403 ( .A(n9643), .B(n9644), .Z(n9639) );
  ANDN U11404 ( .B(n9645), .A(n9646), .Z(n9643) );
  XNOR U11405 ( .A(b[2337]), .B(n9644), .Z(n9645) );
  XNOR U11406 ( .A(b[2337]), .B(n9646), .Z(c[2337]) );
  XNOR U11407 ( .A(a[2337]), .B(n9647), .Z(n9646) );
  IV U11408 ( .A(n9644), .Z(n9647) );
  XOR U11409 ( .A(n9648), .B(n9649), .Z(n9644) );
  ANDN U11410 ( .B(n9650), .A(n9651), .Z(n9648) );
  XNOR U11411 ( .A(b[2336]), .B(n9649), .Z(n9650) );
  XNOR U11412 ( .A(b[2336]), .B(n9651), .Z(c[2336]) );
  XNOR U11413 ( .A(a[2336]), .B(n9652), .Z(n9651) );
  IV U11414 ( .A(n9649), .Z(n9652) );
  XOR U11415 ( .A(n9653), .B(n9654), .Z(n9649) );
  ANDN U11416 ( .B(n9655), .A(n9656), .Z(n9653) );
  XNOR U11417 ( .A(b[2335]), .B(n9654), .Z(n9655) );
  XNOR U11418 ( .A(b[2335]), .B(n9656), .Z(c[2335]) );
  XNOR U11419 ( .A(a[2335]), .B(n9657), .Z(n9656) );
  IV U11420 ( .A(n9654), .Z(n9657) );
  XOR U11421 ( .A(n9658), .B(n9659), .Z(n9654) );
  ANDN U11422 ( .B(n9660), .A(n9661), .Z(n9658) );
  XNOR U11423 ( .A(b[2334]), .B(n9659), .Z(n9660) );
  XNOR U11424 ( .A(b[2334]), .B(n9661), .Z(c[2334]) );
  XNOR U11425 ( .A(a[2334]), .B(n9662), .Z(n9661) );
  IV U11426 ( .A(n9659), .Z(n9662) );
  XOR U11427 ( .A(n9663), .B(n9664), .Z(n9659) );
  ANDN U11428 ( .B(n9665), .A(n9666), .Z(n9663) );
  XNOR U11429 ( .A(b[2333]), .B(n9664), .Z(n9665) );
  XNOR U11430 ( .A(b[2333]), .B(n9666), .Z(c[2333]) );
  XNOR U11431 ( .A(a[2333]), .B(n9667), .Z(n9666) );
  IV U11432 ( .A(n9664), .Z(n9667) );
  XOR U11433 ( .A(n9668), .B(n9669), .Z(n9664) );
  ANDN U11434 ( .B(n9670), .A(n9671), .Z(n9668) );
  XNOR U11435 ( .A(b[2332]), .B(n9669), .Z(n9670) );
  XNOR U11436 ( .A(b[2332]), .B(n9671), .Z(c[2332]) );
  XNOR U11437 ( .A(a[2332]), .B(n9672), .Z(n9671) );
  IV U11438 ( .A(n9669), .Z(n9672) );
  XOR U11439 ( .A(n9673), .B(n9674), .Z(n9669) );
  ANDN U11440 ( .B(n9675), .A(n9676), .Z(n9673) );
  XNOR U11441 ( .A(b[2331]), .B(n9674), .Z(n9675) );
  XNOR U11442 ( .A(b[2331]), .B(n9676), .Z(c[2331]) );
  XNOR U11443 ( .A(a[2331]), .B(n9677), .Z(n9676) );
  IV U11444 ( .A(n9674), .Z(n9677) );
  XOR U11445 ( .A(n9678), .B(n9679), .Z(n9674) );
  ANDN U11446 ( .B(n9680), .A(n9681), .Z(n9678) );
  XNOR U11447 ( .A(b[2330]), .B(n9679), .Z(n9680) );
  XNOR U11448 ( .A(b[2330]), .B(n9681), .Z(c[2330]) );
  XNOR U11449 ( .A(a[2330]), .B(n9682), .Z(n9681) );
  IV U11450 ( .A(n9679), .Z(n9682) );
  XOR U11451 ( .A(n9683), .B(n9684), .Z(n9679) );
  ANDN U11452 ( .B(n9685), .A(n9686), .Z(n9683) );
  XNOR U11453 ( .A(b[2329]), .B(n9684), .Z(n9685) );
  XNOR U11454 ( .A(b[232]), .B(n9687), .Z(c[232]) );
  XNOR U11455 ( .A(b[2329]), .B(n9686), .Z(c[2329]) );
  XNOR U11456 ( .A(a[2329]), .B(n9688), .Z(n9686) );
  IV U11457 ( .A(n9684), .Z(n9688) );
  XOR U11458 ( .A(n9689), .B(n9690), .Z(n9684) );
  ANDN U11459 ( .B(n9691), .A(n9692), .Z(n9689) );
  XNOR U11460 ( .A(b[2328]), .B(n9690), .Z(n9691) );
  XNOR U11461 ( .A(b[2328]), .B(n9692), .Z(c[2328]) );
  XNOR U11462 ( .A(a[2328]), .B(n9693), .Z(n9692) );
  IV U11463 ( .A(n9690), .Z(n9693) );
  XOR U11464 ( .A(n9694), .B(n9695), .Z(n9690) );
  ANDN U11465 ( .B(n9696), .A(n9697), .Z(n9694) );
  XNOR U11466 ( .A(b[2327]), .B(n9695), .Z(n9696) );
  XNOR U11467 ( .A(b[2327]), .B(n9697), .Z(c[2327]) );
  XNOR U11468 ( .A(a[2327]), .B(n9698), .Z(n9697) );
  IV U11469 ( .A(n9695), .Z(n9698) );
  XOR U11470 ( .A(n9699), .B(n9700), .Z(n9695) );
  ANDN U11471 ( .B(n9701), .A(n9702), .Z(n9699) );
  XNOR U11472 ( .A(b[2326]), .B(n9700), .Z(n9701) );
  XNOR U11473 ( .A(b[2326]), .B(n9702), .Z(c[2326]) );
  XNOR U11474 ( .A(a[2326]), .B(n9703), .Z(n9702) );
  IV U11475 ( .A(n9700), .Z(n9703) );
  XOR U11476 ( .A(n9704), .B(n9705), .Z(n9700) );
  ANDN U11477 ( .B(n9706), .A(n9707), .Z(n9704) );
  XNOR U11478 ( .A(b[2325]), .B(n9705), .Z(n9706) );
  XNOR U11479 ( .A(b[2325]), .B(n9707), .Z(c[2325]) );
  XNOR U11480 ( .A(a[2325]), .B(n9708), .Z(n9707) );
  IV U11481 ( .A(n9705), .Z(n9708) );
  XOR U11482 ( .A(n9709), .B(n9710), .Z(n9705) );
  ANDN U11483 ( .B(n9711), .A(n9712), .Z(n9709) );
  XNOR U11484 ( .A(b[2324]), .B(n9710), .Z(n9711) );
  XNOR U11485 ( .A(b[2324]), .B(n9712), .Z(c[2324]) );
  XNOR U11486 ( .A(a[2324]), .B(n9713), .Z(n9712) );
  IV U11487 ( .A(n9710), .Z(n9713) );
  XOR U11488 ( .A(n9714), .B(n9715), .Z(n9710) );
  ANDN U11489 ( .B(n9716), .A(n9717), .Z(n9714) );
  XNOR U11490 ( .A(b[2323]), .B(n9715), .Z(n9716) );
  XNOR U11491 ( .A(b[2323]), .B(n9717), .Z(c[2323]) );
  XNOR U11492 ( .A(a[2323]), .B(n9718), .Z(n9717) );
  IV U11493 ( .A(n9715), .Z(n9718) );
  XOR U11494 ( .A(n9719), .B(n9720), .Z(n9715) );
  ANDN U11495 ( .B(n9721), .A(n9722), .Z(n9719) );
  XNOR U11496 ( .A(b[2322]), .B(n9720), .Z(n9721) );
  XNOR U11497 ( .A(b[2322]), .B(n9722), .Z(c[2322]) );
  XNOR U11498 ( .A(a[2322]), .B(n9723), .Z(n9722) );
  IV U11499 ( .A(n9720), .Z(n9723) );
  XOR U11500 ( .A(n9724), .B(n9725), .Z(n9720) );
  ANDN U11501 ( .B(n9726), .A(n9727), .Z(n9724) );
  XNOR U11502 ( .A(b[2321]), .B(n9725), .Z(n9726) );
  XNOR U11503 ( .A(b[2321]), .B(n9727), .Z(c[2321]) );
  XNOR U11504 ( .A(a[2321]), .B(n9728), .Z(n9727) );
  IV U11505 ( .A(n9725), .Z(n9728) );
  XOR U11506 ( .A(n9729), .B(n9730), .Z(n9725) );
  ANDN U11507 ( .B(n9731), .A(n9732), .Z(n9729) );
  XNOR U11508 ( .A(b[2320]), .B(n9730), .Z(n9731) );
  XNOR U11509 ( .A(b[2320]), .B(n9732), .Z(c[2320]) );
  XNOR U11510 ( .A(a[2320]), .B(n9733), .Z(n9732) );
  IV U11511 ( .A(n9730), .Z(n9733) );
  XOR U11512 ( .A(n9734), .B(n9735), .Z(n9730) );
  ANDN U11513 ( .B(n9736), .A(n9737), .Z(n9734) );
  XNOR U11514 ( .A(b[2319]), .B(n9735), .Z(n9736) );
  XNOR U11515 ( .A(b[231]), .B(n9738), .Z(c[231]) );
  XNOR U11516 ( .A(b[2319]), .B(n9737), .Z(c[2319]) );
  XNOR U11517 ( .A(a[2319]), .B(n9739), .Z(n9737) );
  IV U11518 ( .A(n9735), .Z(n9739) );
  XOR U11519 ( .A(n9740), .B(n9741), .Z(n9735) );
  ANDN U11520 ( .B(n9742), .A(n9743), .Z(n9740) );
  XNOR U11521 ( .A(b[2318]), .B(n9741), .Z(n9742) );
  XNOR U11522 ( .A(b[2318]), .B(n9743), .Z(c[2318]) );
  XNOR U11523 ( .A(a[2318]), .B(n9744), .Z(n9743) );
  IV U11524 ( .A(n9741), .Z(n9744) );
  XOR U11525 ( .A(n9745), .B(n9746), .Z(n9741) );
  ANDN U11526 ( .B(n9747), .A(n9748), .Z(n9745) );
  XNOR U11527 ( .A(b[2317]), .B(n9746), .Z(n9747) );
  XNOR U11528 ( .A(b[2317]), .B(n9748), .Z(c[2317]) );
  XNOR U11529 ( .A(a[2317]), .B(n9749), .Z(n9748) );
  IV U11530 ( .A(n9746), .Z(n9749) );
  XOR U11531 ( .A(n9750), .B(n9751), .Z(n9746) );
  ANDN U11532 ( .B(n9752), .A(n9753), .Z(n9750) );
  XNOR U11533 ( .A(b[2316]), .B(n9751), .Z(n9752) );
  XNOR U11534 ( .A(b[2316]), .B(n9753), .Z(c[2316]) );
  XNOR U11535 ( .A(a[2316]), .B(n9754), .Z(n9753) );
  IV U11536 ( .A(n9751), .Z(n9754) );
  XOR U11537 ( .A(n9755), .B(n9756), .Z(n9751) );
  ANDN U11538 ( .B(n9757), .A(n9758), .Z(n9755) );
  XNOR U11539 ( .A(b[2315]), .B(n9756), .Z(n9757) );
  XNOR U11540 ( .A(b[2315]), .B(n9758), .Z(c[2315]) );
  XNOR U11541 ( .A(a[2315]), .B(n9759), .Z(n9758) );
  IV U11542 ( .A(n9756), .Z(n9759) );
  XOR U11543 ( .A(n9760), .B(n9761), .Z(n9756) );
  ANDN U11544 ( .B(n9762), .A(n9763), .Z(n9760) );
  XNOR U11545 ( .A(b[2314]), .B(n9761), .Z(n9762) );
  XNOR U11546 ( .A(b[2314]), .B(n9763), .Z(c[2314]) );
  XNOR U11547 ( .A(a[2314]), .B(n9764), .Z(n9763) );
  IV U11548 ( .A(n9761), .Z(n9764) );
  XOR U11549 ( .A(n9765), .B(n9766), .Z(n9761) );
  ANDN U11550 ( .B(n9767), .A(n9768), .Z(n9765) );
  XNOR U11551 ( .A(b[2313]), .B(n9766), .Z(n9767) );
  XNOR U11552 ( .A(b[2313]), .B(n9768), .Z(c[2313]) );
  XNOR U11553 ( .A(a[2313]), .B(n9769), .Z(n9768) );
  IV U11554 ( .A(n9766), .Z(n9769) );
  XOR U11555 ( .A(n9770), .B(n9771), .Z(n9766) );
  ANDN U11556 ( .B(n9772), .A(n9773), .Z(n9770) );
  XNOR U11557 ( .A(b[2312]), .B(n9771), .Z(n9772) );
  XNOR U11558 ( .A(b[2312]), .B(n9773), .Z(c[2312]) );
  XNOR U11559 ( .A(a[2312]), .B(n9774), .Z(n9773) );
  IV U11560 ( .A(n9771), .Z(n9774) );
  XOR U11561 ( .A(n9775), .B(n9776), .Z(n9771) );
  ANDN U11562 ( .B(n9777), .A(n9778), .Z(n9775) );
  XNOR U11563 ( .A(b[2311]), .B(n9776), .Z(n9777) );
  XNOR U11564 ( .A(b[2311]), .B(n9778), .Z(c[2311]) );
  XNOR U11565 ( .A(a[2311]), .B(n9779), .Z(n9778) );
  IV U11566 ( .A(n9776), .Z(n9779) );
  XOR U11567 ( .A(n9780), .B(n9781), .Z(n9776) );
  ANDN U11568 ( .B(n9782), .A(n9783), .Z(n9780) );
  XNOR U11569 ( .A(b[2310]), .B(n9781), .Z(n9782) );
  XNOR U11570 ( .A(b[2310]), .B(n9783), .Z(c[2310]) );
  XNOR U11571 ( .A(a[2310]), .B(n9784), .Z(n9783) );
  IV U11572 ( .A(n9781), .Z(n9784) );
  XOR U11573 ( .A(n9785), .B(n9786), .Z(n9781) );
  ANDN U11574 ( .B(n9787), .A(n9788), .Z(n9785) );
  XNOR U11575 ( .A(b[2309]), .B(n9786), .Z(n9787) );
  XNOR U11576 ( .A(b[230]), .B(n9789), .Z(c[230]) );
  XNOR U11577 ( .A(b[2309]), .B(n9788), .Z(c[2309]) );
  XNOR U11578 ( .A(a[2309]), .B(n9790), .Z(n9788) );
  IV U11579 ( .A(n9786), .Z(n9790) );
  XOR U11580 ( .A(n9791), .B(n9792), .Z(n9786) );
  ANDN U11581 ( .B(n9793), .A(n9794), .Z(n9791) );
  XNOR U11582 ( .A(b[2308]), .B(n9792), .Z(n9793) );
  XNOR U11583 ( .A(b[2308]), .B(n9794), .Z(c[2308]) );
  XNOR U11584 ( .A(a[2308]), .B(n9795), .Z(n9794) );
  IV U11585 ( .A(n9792), .Z(n9795) );
  XOR U11586 ( .A(n9796), .B(n9797), .Z(n9792) );
  ANDN U11587 ( .B(n9798), .A(n9799), .Z(n9796) );
  XNOR U11588 ( .A(b[2307]), .B(n9797), .Z(n9798) );
  XNOR U11589 ( .A(b[2307]), .B(n9799), .Z(c[2307]) );
  XNOR U11590 ( .A(a[2307]), .B(n9800), .Z(n9799) );
  IV U11591 ( .A(n9797), .Z(n9800) );
  XOR U11592 ( .A(n9801), .B(n9802), .Z(n9797) );
  ANDN U11593 ( .B(n9803), .A(n9804), .Z(n9801) );
  XNOR U11594 ( .A(b[2306]), .B(n9802), .Z(n9803) );
  XNOR U11595 ( .A(b[2306]), .B(n9804), .Z(c[2306]) );
  XNOR U11596 ( .A(a[2306]), .B(n9805), .Z(n9804) );
  IV U11597 ( .A(n9802), .Z(n9805) );
  XOR U11598 ( .A(n9806), .B(n9807), .Z(n9802) );
  ANDN U11599 ( .B(n9808), .A(n9809), .Z(n9806) );
  XNOR U11600 ( .A(b[2305]), .B(n9807), .Z(n9808) );
  XNOR U11601 ( .A(b[2305]), .B(n9809), .Z(c[2305]) );
  XNOR U11602 ( .A(a[2305]), .B(n9810), .Z(n9809) );
  IV U11603 ( .A(n9807), .Z(n9810) );
  XOR U11604 ( .A(n9811), .B(n9812), .Z(n9807) );
  ANDN U11605 ( .B(n9813), .A(n9814), .Z(n9811) );
  XNOR U11606 ( .A(b[2304]), .B(n9812), .Z(n9813) );
  XNOR U11607 ( .A(b[2304]), .B(n9814), .Z(c[2304]) );
  XNOR U11608 ( .A(a[2304]), .B(n9815), .Z(n9814) );
  IV U11609 ( .A(n9812), .Z(n9815) );
  XOR U11610 ( .A(n9816), .B(n9817), .Z(n9812) );
  ANDN U11611 ( .B(n9818), .A(n9819), .Z(n9816) );
  XNOR U11612 ( .A(b[2303]), .B(n9817), .Z(n9818) );
  XNOR U11613 ( .A(b[2303]), .B(n9819), .Z(c[2303]) );
  XNOR U11614 ( .A(a[2303]), .B(n9820), .Z(n9819) );
  IV U11615 ( .A(n9817), .Z(n9820) );
  XOR U11616 ( .A(n9821), .B(n9822), .Z(n9817) );
  ANDN U11617 ( .B(n9823), .A(n9824), .Z(n9821) );
  XNOR U11618 ( .A(b[2302]), .B(n9822), .Z(n9823) );
  XNOR U11619 ( .A(b[2302]), .B(n9824), .Z(c[2302]) );
  XNOR U11620 ( .A(a[2302]), .B(n9825), .Z(n9824) );
  IV U11621 ( .A(n9822), .Z(n9825) );
  XOR U11622 ( .A(n9826), .B(n9827), .Z(n9822) );
  ANDN U11623 ( .B(n9828), .A(n9829), .Z(n9826) );
  XNOR U11624 ( .A(b[2301]), .B(n9827), .Z(n9828) );
  XNOR U11625 ( .A(b[2301]), .B(n9829), .Z(c[2301]) );
  XNOR U11626 ( .A(a[2301]), .B(n9830), .Z(n9829) );
  IV U11627 ( .A(n9827), .Z(n9830) );
  XOR U11628 ( .A(n9831), .B(n9832), .Z(n9827) );
  ANDN U11629 ( .B(n9833), .A(n9834), .Z(n9831) );
  XNOR U11630 ( .A(b[2300]), .B(n9832), .Z(n9833) );
  XNOR U11631 ( .A(b[2300]), .B(n9834), .Z(c[2300]) );
  XNOR U11632 ( .A(a[2300]), .B(n9835), .Z(n9834) );
  IV U11633 ( .A(n9832), .Z(n9835) );
  XOR U11634 ( .A(n9836), .B(n9837), .Z(n9832) );
  ANDN U11635 ( .B(n9838), .A(n9839), .Z(n9836) );
  XNOR U11636 ( .A(b[2299]), .B(n9837), .Z(n9838) );
  XNOR U11637 ( .A(b[22]), .B(n9840), .Z(c[22]) );
  XNOR U11638 ( .A(b[229]), .B(n9841), .Z(c[229]) );
  XNOR U11639 ( .A(b[2299]), .B(n9839), .Z(c[2299]) );
  XNOR U11640 ( .A(a[2299]), .B(n9842), .Z(n9839) );
  IV U11641 ( .A(n9837), .Z(n9842) );
  XOR U11642 ( .A(n9843), .B(n9844), .Z(n9837) );
  ANDN U11643 ( .B(n9845), .A(n9846), .Z(n9843) );
  XNOR U11644 ( .A(b[2298]), .B(n9844), .Z(n9845) );
  XNOR U11645 ( .A(b[2298]), .B(n9846), .Z(c[2298]) );
  XNOR U11646 ( .A(a[2298]), .B(n9847), .Z(n9846) );
  IV U11647 ( .A(n9844), .Z(n9847) );
  XOR U11648 ( .A(n9848), .B(n9849), .Z(n9844) );
  ANDN U11649 ( .B(n9850), .A(n9851), .Z(n9848) );
  XNOR U11650 ( .A(b[2297]), .B(n9849), .Z(n9850) );
  XNOR U11651 ( .A(b[2297]), .B(n9851), .Z(c[2297]) );
  XNOR U11652 ( .A(a[2297]), .B(n9852), .Z(n9851) );
  IV U11653 ( .A(n9849), .Z(n9852) );
  XOR U11654 ( .A(n9853), .B(n9854), .Z(n9849) );
  ANDN U11655 ( .B(n9855), .A(n9856), .Z(n9853) );
  XNOR U11656 ( .A(b[2296]), .B(n9854), .Z(n9855) );
  XNOR U11657 ( .A(b[2296]), .B(n9856), .Z(c[2296]) );
  XNOR U11658 ( .A(a[2296]), .B(n9857), .Z(n9856) );
  IV U11659 ( .A(n9854), .Z(n9857) );
  XOR U11660 ( .A(n9858), .B(n9859), .Z(n9854) );
  ANDN U11661 ( .B(n9860), .A(n9861), .Z(n9858) );
  XNOR U11662 ( .A(b[2295]), .B(n9859), .Z(n9860) );
  XNOR U11663 ( .A(b[2295]), .B(n9861), .Z(c[2295]) );
  XNOR U11664 ( .A(a[2295]), .B(n9862), .Z(n9861) );
  IV U11665 ( .A(n9859), .Z(n9862) );
  XOR U11666 ( .A(n9863), .B(n9864), .Z(n9859) );
  ANDN U11667 ( .B(n9865), .A(n9866), .Z(n9863) );
  XNOR U11668 ( .A(b[2294]), .B(n9864), .Z(n9865) );
  XNOR U11669 ( .A(b[2294]), .B(n9866), .Z(c[2294]) );
  XNOR U11670 ( .A(a[2294]), .B(n9867), .Z(n9866) );
  IV U11671 ( .A(n9864), .Z(n9867) );
  XOR U11672 ( .A(n9868), .B(n9869), .Z(n9864) );
  ANDN U11673 ( .B(n9870), .A(n9871), .Z(n9868) );
  XNOR U11674 ( .A(b[2293]), .B(n9869), .Z(n9870) );
  XNOR U11675 ( .A(b[2293]), .B(n9871), .Z(c[2293]) );
  XNOR U11676 ( .A(a[2293]), .B(n9872), .Z(n9871) );
  IV U11677 ( .A(n9869), .Z(n9872) );
  XOR U11678 ( .A(n9873), .B(n9874), .Z(n9869) );
  ANDN U11679 ( .B(n9875), .A(n9876), .Z(n9873) );
  XNOR U11680 ( .A(b[2292]), .B(n9874), .Z(n9875) );
  XNOR U11681 ( .A(b[2292]), .B(n9876), .Z(c[2292]) );
  XNOR U11682 ( .A(a[2292]), .B(n9877), .Z(n9876) );
  IV U11683 ( .A(n9874), .Z(n9877) );
  XOR U11684 ( .A(n9878), .B(n9879), .Z(n9874) );
  ANDN U11685 ( .B(n9880), .A(n9881), .Z(n9878) );
  XNOR U11686 ( .A(b[2291]), .B(n9879), .Z(n9880) );
  XNOR U11687 ( .A(b[2291]), .B(n9881), .Z(c[2291]) );
  XNOR U11688 ( .A(a[2291]), .B(n9882), .Z(n9881) );
  IV U11689 ( .A(n9879), .Z(n9882) );
  XOR U11690 ( .A(n9883), .B(n9884), .Z(n9879) );
  ANDN U11691 ( .B(n9885), .A(n9886), .Z(n9883) );
  XNOR U11692 ( .A(b[2290]), .B(n9884), .Z(n9885) );
  XNOR U11693 ( .A(b[2290]), .B(n9886), .Z(c[2290]) );
  XNOR U11694 ( .A(a[2290]), .B(n9887), .Z(n9886) );
  IV U11695 ( .A(n9884), .Z(n9887) );
  XOR U11696 ( .A(n9888), .B(n9889), .Z(n9884) );
  ANDN U11697 ( .B(n9890), .A(n9891), .Z(n9888) );
  XNOR U11698 ( .A(b[2289]), .B(n9889), .Z(n9890) );
  XNOR U11699 ( .A(b[228]), .B(n9892), .Z(c[228]) );
  XNOR U11700 ( .A(b[2289]), .B(n9891), .Z(c[2289]) );
  XNOR U11701 ( .A(a[2289]), .B(n9893), .Z(n9891) );
  IV U11702 ( .A(n9889), .Z(n9893) );
  XOR U11703 ( .A(n9894), .B(n9895), .Z(n9889) );
  ANDN U11704 ( .B(n9896), .A(n9897), .Z(n9894) );
  XNOR U11705 ( .A(b[2288]), .B(n9895), .Z(n9896) );
  XNOR U11706 ( .A(b[2288]), .B(n9897), .Z(c[2288]) );
  XNOR U11707 ( .A(a[2288]), .B(n9898), .Z(n9897) );
  IV U11708 ( .A(n9895), .Z(n9898) );
  XOR U11709 ( .A(n9899), .B(n9900), .Z(n9895) );
  ANDN U11710 ( .B(n9901), .A(n9902), .Z(n9899) );
  XNOR U11711 ( .A(b[2287]), .B(n9900), .Z(n9901) );
  XNOR U11712 ( .A(b[2287]), .B(n9902), .Z(c[2287]) );
  XNOR U11713 ( .A(a[2287]), .B(n9903), .Z(n9902) );
  IV U11714 ( .A(n9900), .Z(n9903) );
  XOR U11715 ( .A(n9904), .B(n9905), .Z(n9900) );
  ANDN U11716 ( .B(n9906), .A(n9907), .Z(n9904) );
  XNOR U11717 ( .A(b[2286]), .B(n9905), .Z(n9906) );
  XNOR U11718 ( .A(b[2286]), .B(n9907), .Z(c[2286]) );
  XNOR U11719 ( .A(a[2286]), .B(n9908), .Z(n9907) );
  IV U11720 ( .A(n9905), .Z(n9908) );
  XOR U11721 ( .A(n9909), .B(n9910), .Z(n9905) );
  ANDN U11722 ( .B(n9911), .A(n9912), .Z(n9909) );
  XNOR U11723 ( .A(b[2285]), .B(n9910), .Z(n9911) );
  XNOR U11724 ( .A(b[2285]), .B(n9912), .Z(c[2285]) );
  XNOR U11725 ( .A(a[2285]), .B(n9913), .Z(n9912) );
  IV U11726 ( .A(n9910), .Z(n9913) );
  XOR U11727 ( .A(n9914), .B(n9915), .Z(n9910) );
  ANDN U11728 ( .B(n9916), .A(n9917), .Z(n9914) );
  XNOR U11729 ( .A(b[2284]), .B(n9915), .Z(n9916) );
  XNOR U11730 ( .A(b[2284]), .B(n9917), .Z(c[2284]) );
  XNOR U11731 ( .A(a[2284]), .B(n9918), .Z(n9917) );
  IV U11732 ( .A(n9915), .Z(n9918) );
  XOR U11733 ( .A(n9919), .B(n9920), .Z(n9915) );
  ANDN U11734 ( .B(n9921), .A(n9922), .Z(n9919) );
  XNOR U11735 ( .A(b[2283]), .B(n9920), .Z(n9921) );
  XNOR U11736 ( .A(b[2283]), .B(n9922), .Z(c[2283]) );
  XNOR U11737 ( .A(a[2283]), .B(n9923), .Z(n9922) );
  IV U11738 ( .A(n9920), .Z(n9923) );
  XOR U11739 ( .A(n9924), .B(n9925), .Z(n9920) );
  ANDN U11740 ( .B(n9926), .A(n9927), .Z(n9924) );
  XNOR U11741 ( .A(b[2282]), .B(n9925), .Z(n9926) );
  XNOR U11742 ( .A(b[2282]), .B(n9927), .Z(c[2282]) );
  XNOR U11743 ( .A(a[2282]), .B(n9928), .Z(n9927) );
  IV U11744 ( .A(n9925), .Z(n9928) );
  XOR U11745 ( .A(n9929), .B(n9930), .Z(n9925) );
  ANDN U11746 ( .B(n9931), .A(n9932), .Z(n9929) );
  XNOR U11747 ( .A(b[2281]), .B(n9930), .Z(n9931) );
  XNOR U11748 ( .A(b[2281]), .B(n9932), .Z(c[2281]) );
  XNOR U11749 ( .A(a[2281]), .B(n9933), .Z(n9932) );
  IV U11750 ( .A(n9930), .Z(n9933) );
  XOR U11751 ( .A(n9934), .B(n9935), .Z(n9930) );
  ANDN U11752 ( .B(n9936), .A(n9937), .Z(n9934) );
  XNOR U11753 ( .A(b[2280]), .B(n9935), .Z(n9936) );
  XNOR U11754 ( .A(b[2280]), .B(n9937), .Z(c[2280]) );
  XNOR U11755 ( .A(a[2280]), .B(n9938), .Z(n9937) );
  IV U11756 ( .A(n9935), .Z(n9938) );
  XOR U11757 ( .A(n9939), .B(n9940), .Z(n9935) );
  ANDN U11758 ( .B(n9941), .A(n9942), .Z(n9939) );
  XNOR U11759 ( .A(b[2279]), .B(n9940), .Z(n9941) );
  XNOR U11760 ( .A(b[227]), .B(n9943), .Z(c[227]) );
  XNOR U11761 ( .A(b[2279]), .B(n9942), .Z(c[2279]) );
  XNOR U11762 ( .A(a[2279]), .B(n9944), .Z(n9942) );
  IV U11763 ( .A(n9940), .Z(n9944) );
  XOR U11764 ( .A(n9945), .B(n9946), .Z(n9940) );
  ANDN U11765 ( .B(n9947), .A(n9948), .Z(n9945) );
  XNOR U11766 ( .A(b[2278]), .B(n9946), .Z(n9947) );
  XNOR U11767 ( .A(b[2278]), .B(n9948), .Z(c[2278]) );
  XNOR U11768 ( .A(a[2278]), .B(n9949), .Z(n9948) );
  IV U11769 ( .A(n9946), .Z(n9949) );
  XOR U11770 ( .A(n9950), .B(n9951), .Z(n9946) );
  ANDN U11771 ( .B(n9952), .A(n9953), .Z(n9950) );
  XNOR U11772 ( .A(b[2277]), .B(n9951), .Z(n9952) );
  XNOR U11773 ( .A(b[2277]), .B(n9953), .Z(c[2277]) );
  XNOR U11774 ( .A(a[2277]), .B(n9954), .Z(n9953) );
  IV U11775 ( .A(n9951), .Z(n9954) );
  XOR U11776 ( .A(n9955), .B(n9956), .Z(n9951) );
  ANDN U11777 ( .B(n9957), .A(n9958), .Z(n9955) );
  XNOR U11778 ( .A(b[2276]), .B(n9956), .Z(n9957) );
  XNOR U11779 ( .A(b[2276]), .B(n9958), .Z(c[2276]) );
  XNOR U11780 ( .A(a[2276]), .B(n9959), .Z(n9958) );
  IV U11781 ( .A(n9956), .Z(n9959) );
  XOR U11782 ( .A(n9960), .B(n9961), .Z(n9956) );
  ANDN U11783 ( .B(n9962), .A(n9963), .Z(n9960) );
  XNOR U11784 ( .A(b[2275]), .B(n9961), .Z(n9962) );
  XNOR U11785 ( .A(b[2275]), .B(n9963), .Z(c[2275]) );
  XNOR U11786 ( .A(a[2275]), .B(n9964), .Z(n9963) );
  IV U11787 ( .A(n9961), .Z(n9964) );
  XOR U11788 ( .A(n9965), .B(n9966), .Z(n9961) );
  ANDN U11789 ( .B(n9967), .A(n9968), .Z(n9965) );
  XNOR U11790 ( .A(b[2274]), .B(n9966), .Z(n9967) );
  XNOR U11791 ( .A(b[2274]), .B(n9968), .Z(c[2274]) );
  XNOR U11792 ( .A(a[2274]), .B(n9969), .Z(n9968) );
  IV U11793 ( .A(n9966), .Z(n9969) );
  XOR U11794 ( .A(n9970), .B(n9971), .Z(n9966) );
  ANDN U11795 ( .B(n9972), .A(n9973), .Z(n9970) );
  XNOR U11796 ( .A(b[2273]), .B(n9971), .Z(n9972) );
  XNOR U11797 ( .A(b[2273]), .B(n9973), .Z(c[2273]) );
  XNOR U11798 ( .A(a[2273]), .B(n9974), .Z(n9973) );
  IV U11799 ( .A(n9971), .Z(n9974) );
  XOR U11800 ( .A(n9975), .B(n9976), .Z(n9971) );
  ANDN U11801 ( .B(n9977), .A(n9978), .Z(n9975) );
  XNOR U11802 ( .A(b[2272]), .B(n9976), .Z(n9977) );
  XNOR U11803 ( .A(b[2272]), .B(n9978), .Z(c[2272]) );
  XNOR U11804 ( .A(a[2272]), .B(n9979), .Z(n9978) );
  IV U11805 ( .A(n9976), .Z(n9979) );
  XOR U11806 ( .A(n9980), .B(n9981), .Z(n9976) );
  ANDN U11807 ( .B(n9982), .A(n9983), .Z(n9980) );
  XNOR U11808 ( .A(b[2271]), .B(n9981), .Z(n9982) );
  XNOR U11809 ( .A(b[2271]), .B(n9983), .Z(c[2271]) );
  XNOR U11810 ( .A(a[2271]), .B(n9984), .Z(n9983) );
  IV U11811 ( .A(n9981), .Z(n9984) );
  XOR U11812 ( .A(n9985), .B(n9986), .Z(n9981) );
  ANDN U11813 ( .B(n9987), .A(n9988), .Z(n9985) );
  XNOR U11814 ( .A(b[2270]), .B(n9986), .Z(n9987) );
  XNOR U11815 ( .A(b[2270]), .B(n9988), .Z(c[2270]) );
  XNOR U11816 ( .A(a[2270]), .B(n9989), .Z(n9988) );
  IV U11817 ( .A(n9986), .Z(n9989) );
  XOR U11818 ( .A(n9990), .B(n9991), .Z(n9986) );
  ANDN U11819 ( .B(n9992), .A(n9993), .Z(n9990) );
  XNOR U11820 ( .A(b[2269]), .B(n9991), .Z(n9992) );
  XNOR U11821 ( .A(b[226]), .B(n9994), .Z(c[226]) );
  XNOR U11822 ( .A(b[2269]), .B(n9993), .Z(c[2269]) );
  XNOR U11823 ( .A(a[2269]), .B(n9995), .Z(n9993) );
  IV U11824 ( .A(n9991), .Z(n9995) );
  XOR U11825 ( .A(n9996), .B(n9997), .Z(n9991) );
  ANDN U11826 ( .B(n9998), .A(n9999), .Z(n9996) );
  XNOR U11827 ( .A(b[2268]), .B(n9997), .Z(n9998) );
  XNOR U11828 ( .A(b[2268]), .B(n9999), .Z(c[2268]) );
  XNOR U11829 ( .A(a[2268]), .B(n10000), .Z(n9999) );
  IV U11830 ( .A(n9997), .Z(n10000) );
  XOR U11831 ( .A(n10001), .B(n10002), .Z(n9997) );
  ANDN U11832 ( .B(n10003), .A(n10004), .Z(n10001) );
  XNOR U11833 ( .A(b[2267]), .B(n10002), .Z(n10003) );
  XNOR U11834 ( .A(b[2267]), .B(n10004), .Z(c[2267]) );
  XNOR U11835 ( .A(a[2267]), .B(n10005), .Z(n10004) );
  IV U11836 ( .A(n10002), .Z(n10005) );
  XOR U11837 ( .A(n10006), .B(n10007), .Z(n10002) );
  ANDN U11838 ( .B(n10008), .A(n10009), .Z(n10006) );
  XNOR U11839 ( .A(b[2266]), .B(n10007), .Z(n10008) );
  XNOR U11840 ( .A(b[2266]), .B(n10009), .Z(c[2266]) );
  XNOR U11841 ( .A(a[2266]), .B(n10010), .Z(n10009) );
  IV U11842 ( .A(n10007), .Z(n10010) );
  XOR U11843 ( .A(n10011), .B(n10012), .Z(n10007) );
  ANDN U11844 ( .B(n10013), .A(n10014), .Z(n10011) );
  XNOR U11845 ( .A(b[2265]), .B(n10012), .Z(n10013) );
  XNOR U11846 ( .A(b[2265]), .B(n10014), .Z(c[2265]) );
  XNOR U11847 ( .A(a[2265]), .B(n10015), .Z(n10014) );
  IV U11848 ( .A(n10012), .Z(n10015) );
  XOR U11849 ( .A(n10016), .B(n10017), .Z(n10012) );
  ANDN U11850 ( .B(n10018), .A(n10019), .Z(n10016) );
  XNOR U11851 ( .A(b[2264]), .B(n10017), .Z(n10018) );
  XNOR U11852 ( .A(b[2264]), .B(n10019), .Z(c[2264]) );
  XNOR U11853 ( .A(a[2264]), .B(n10020), .Z(n10019) );
  IV U11854 ( .A(n10017), .Z(n10020) );
  XOR U11855 ( .A(n10021), .B(n10022), .Z(n10017) );
  ANDN U11856 ( .B(n10023), .A(n10024), .Z(n10021) );
  XNOR U11857 ( .A(b[2263]), .B(n10022), .Z(n10023) );
  XNOR U11858 ( .A(b[2263]), .B(n10024), .Z(c[2263]) );
  XNOR U11859 ( .A(a[2263]), .B(n10025), .Z(n10024) );
  IV U11860 ( .A(n10022), .Z(n10025) );
  XOR U11861 ( .A(n10026), .B(n10027), .Z(n10022) );
  ANDN U11862 ( .B(n10028), .A(n10029), .Z(n10026) );
  XNOR U11863 ( .A(b[2262]), .B(n10027), .Z(n10028) );
  XNOR U11864 ( .A(b[2262]), .B(n10029), .Z(c[2262]) );
  XNOR U11865 ( .A(a[2262]), .B(n10030), .Z(n10029) );
  IV U11866 ( .A(n10027), .Z(n10030) );
  XOR U11867 ( .A(n10031), .B(n10032), .Z(n10027) );
  ANDN U11868 ( .B(n10033), .A(n10034), .Z(n10031) );
  XNOR U11869 ( .A(b[2261]), .B(n10032), .Z(n10033) );
  XNOR U11870 ( .A(b[2261]), .B(n10034), .Z(c[2261]) );
  XNOR U11871 ( .A(a[2261]), .B(n10035), .Z(n10034) );
  IV U11872 ( .A(n10032), .Z(n10035) );
  XOR U11873 ( .A(n10036), .B(n10037), .Z(n10032) );
  ANDN U11874 ( .B(n10038), .A(n10039), .Z(n10036) );
  XNOR U11875 ( .A(b[2260]), .B(n10037), .Z(n10038) );
  XNOR U11876 ( .A(b[2260]), .B(n10039), .Z(c[2260]) );
  XNOR U11877 ( .A(a[2260]), .B(n10040), .Z(n10039) );
  IV U11878 ( .A(n10037), .Z(n10040) );
  XOR U11879 ( .A(n10041), .B(n10042), .Z(n10037) );
  ANDN U11880 ( .B(n10043), .A(n10044), .Z(n10041) );
  XNOR U11881 ( .A(b[2259]), .B(n10042), .Z(n10043) );
  XNOR U11882 ( .A(b[225]), .B(n10045), .Z(c[225]) );
  XNOR U11883 ( .A(b[2259]), .B(n10044), .Z(c[2259]) );
  XNOR U11884 ( .A(a[2259]), .B(n10046), .Z(n10044) );
  IV U11885 ( .A(n10042), .Z(n10046) );
  XOR U11886 ( .A(n10047), .B(n10048), .Z(n10042) );
  ANDN U11887 ( .B(n10049), .A(n10050), .Z(n10047) );
  XNOR U11888 ( .A(b[2258]), .B(n10048), .Z(n10049) );
  XNOR U11889 ( .A(b[2258]), .B(n10050), .Z(c[2258]) );
  XNOR U11890 ( .A(a[2258]), .B(n10051), .Z(n10050) );
  IV U11891 ( .A(n10048), .Z(n10051) );
  XOR U11892 ( .A(n10052), .B(n10053), .Z(n10048) );
  ANDN U11893 ( .B(n10054), .A(n10055), .Z(n10052) );
  XNOR U11894 ( .A(b[2257]), .B(n10053), .Z(n10054) );
  XNOR U11895 ( .A(b[2257]), .B(n10055), .Z(c[2257]) );
  XNOR U11896 ( .A(a[2257]), .B(n10056), .Z(n10055) );
  IV U11897 ( .A(n10053), .Z(n10056) );
  XOR U11898 ( .A(n10057), .B(n10058), .Z(n10053) );
  ANDN U11899 ( .B(n10059), .A(n10060), .Z(n10057) );
  XNOR U11900 ( .A(b[2256]), .B(n10058), .Z(n10059) );
  XNOR U11901 ( .A(b[2256]), .B(n10060), .Z(c[2256]) );
  XNOR U11902 ( .A(a[2256]), .B(n10061), .Z(n10060) );
  IV U11903 ( .A(n10058), .Z(n10061) );
  XOR U11904 ( .A(n10062), .B(n10063), .Z(n10058) );
  ANDN U11905 ( .B(n10064), .A(n10065), .Z(n10062) );
  XNOR U11906 ( .A(b[2255]), .B(n10063), .Z(n10064) );
  XNOR U11907 ( .A(b[2255]), .B(n10065), .Z(c[2255]) );
  XNOR U11908 ( .A(a[2255]), .B(n10066), .Z(n10065) );
  IV U11909 ( .A(n10063), .Z(n10066) );
  XOR U11910 ( .A(n10067), .B(n10068), .Z(n10063) );
  ANDN U11911 ( .B(n10069), .A(n10070), .Z(n10067) );
  XNOR U11912 ( .A(b[2254]), .B(n10068), .Z(n10069) );
  XNOR U11913 ( .A(b[2254]), .B(n10070), .Z(c[2254]) );
  XNOR U11914 ( .A(a[2254]), .B(n10071), .Z(n10070) );
  IV U11915 ( .A(n10068), .Z(n10071) );
  XOR U11916 ( .A(n10072), .B(n10073), .Z(n10068) );
  ANDN U11917 ( .B(n10074), .A(n10075), .Z(n10072) );
  XNOR U11918 ( .A(b[2253]), .B(n10073), .Z(n10074) );
  XNOR U11919 ( .A(b[2253]), .B(n10075), .Z(c[2253]) );
  XNOR U11920 ( .A(a[2253]), .B(n10076), .Z(n10075) );
  IV U11921 ( .A(n10073), .Z(n10076) );
  XOR U11922 ( .A(n10077), .B(n10078), .Z(n10073) );
  ANDN U11923 ( .B(n10079), .A(n10080), .Z(n10077) );
  XNOR U11924 ( .A(b[2252]), .B(n10078), .Z(n10079) );
  XNOR U11925 ( .A(b[2252]), .B(n10080), .Z(c[2252]) );
  XNOR U11926 ( .A(a[2252]), .B(n10081), .Z(n10080) );
  IV U11927 ( .A(n10078), .Z(n10081) );
  XOR U11928 ( .A(n10082), .B(n10083), .Z(n10078) );
  ANDN U11929 ( .B(n10084), .A(n10085), .Z(n10082) );
  XNOR U11930 ( .A(b[2251]), .B(n10083), .Z(n10084) );
  XNOR U11931 ( .A(b[2251]), .B(n10085), .Z(c[2251]) );
  XNOR U11932 ( .A(a[2251]), .B(n10086), .Z(n10085) );
  IV U11933 ( .A(n10083), .Z(n10086) );
  XOR U11934 ( .A(n10087), .B(n10088), .Z(n10083) );
  ANDN U11935 ( .B(n10089), .A(n10090), .Z(n10087) );
  XNOR U11936 ( .A(b[2250]), .B(n10088), .Z(n10089) );
  XNOR U11937 ( .A(b[2250]), .B(n10090), .Z(c[2250]) );
  XNOR U11938 ( .A(a[2250]), .B(n10091), .Z(n10090) );
  IV U11939 ( .A(n10088), .Z(n10091) );
  XOR U11940 ( .A(n10092), .B(n10093), .Z(n10088) );
  ANDN U11941 ( .B(n10094), .A(n10095), .Z(n10092) );
  XNOR U11942 ( .A(b[2249]), .B(n10093), .Z(n10094) );
  XNOR U11943 ( .A(b[224]), .B(n10096), .Z(c[224]) );
  XNOR U11944 ( .A(b[2249]), .B(n10095), .Z(c[2249]) );
  XNOR U11945 ( .A(a[2249]), .B(n10097), .Z(n10095) );
  IV U11946 ( .A(n10093), .Z(n10097) );
  XOR U11947 ( .A(n10098), .B(n10099), .Z(n10093) );
  ANDN U11948 ( .B(n10100), .A(n10101), .Z(n10098) );
  XNOR U11949 ( .A(b[2248]), .B(n10099), .Z(n10100) );
  XNOR U11950 ( .A(b[2248]), .B(n10101), .Z(c[2248]) );
  XNOR U11951 ( .A(a[2248]), .B(n10102), .Z(n10101) );
  IV U11952 ( .A(n10099), .Z(n10102) );
  XOR U11953 ( .A(n10103), .B(n10104), .Z(n10099) );
  ANDN U11954 ( .B(n10105), .A(n10106), .Z(n10103) );
  XNOR U11955 ( .A(b[2247]), .B(n10104), .Z(n10105) );
  XNOR U11956 ( .A(b[2247]), .B(n10106), .Z(c[2247]) );
  XNOR U11957 ( .A(a[2247]), .B(n10107), .Z(n10106) );
  IV U11958 ( .A(n10104), .Z(n10107) );
  XOR U11959 ( .A(n10108), .B(n10109), .Z(n10104) );
  ANDN U11960 ( .B(n10110), .A(n10111), .Z(n10108) );
  XNOR U11961 ( .A(b[2246]), .B(n10109), .Z(n10110) );
  XNOR U11962 ( .A(b[2246]), .B(n10111), .Z(c[2246]) );
  XNOR U11963 ( .A(a[2246]), .B(n10112), .Z(n10111) );
  IV U11964 ( .A(n10109), .Z(n10112) );
  XOR U11965 ( .A(n10113), .B(n10114), .Z(n10109) );
  ANDN U11966 ( .B(n10115), .A(n10116), .Z(n10113) );
  XNOR U11967 ( .A(b[2245]), .B(n10114), .Z(n10115) );
  XNOR U11968 ( .A(b[2245]), .B(n10116), .Z(c[2245]) );
  XNOR U11969 ( .A(a[2245]), .B(n10117), .Z(n10116) );
  IV U11970 ( .A(n10114), .Z(n10117) );
  XOR U11971 ( .A(n10118), .B(n10119), .Z(n10114) );
  ANDN U11972 ( .B(n10120), .A(n10121), .Z(n10118) );
  XNOR U11973 ( .A(b[2244]), .B(n10119), .Z(n10120) );
  XNOR U11974 ( .A(b[2244]), .B(n10121), .Z(c[2244]) );
  XNOR U11975 ( .A(a[2244]), .B(n10122), .Z(n10121) );
  IV U11976 ( .A(n10119), .Z(n10122) );
  XOR U11977 ( .A(n10123), .B(n10124), .Z(n10119) );
  ANDN U11978 ( .B(n10125), .A(n10126), .Z(n10123) );
  XNOR U11979 ( .A(b[2243]), .B(n10124), .Z(n10125) );
  XNOR U11980 ( .A(b[2243]), .B(n10126), .Z(c[2243]) );
  XNOR U11981 ( .A(a[2243]), .B(n10127), .Z(n10126) );
  IV U11982 ( .A(n10124), .Z(n10127) );
  XOR U11983 ( .A(n10128), .B(n10129), .Z(n10124) );
  ANDN U11984 ( .B(n10130), .A(n10131), .Z(n10128) );
  XNOR U11985 ( .A(b[2242]), .B(n10129), .Z(n10130) );
  XNOR U11986 ( .A(b[2242]), .B(n10131), .Z(c[2242]) );
  XNOR U11987 ( .A(a[2242]), .B(n10132), .Z(n10131) );
  IV U11988 ( .A(n10129), .Z(n10132) );
  XOR U11989 ( .A(n10133), .B(n10134), .Z(n10129) );
  ANDN U11990 ( .B(n10135), .A(n10136), .Z(n10133) );
  XNOR U11991 ( .A(b[2241]), .B(n10134), .Z(n10135) );
  XNOR U11992 ( .A(b[2241]), .B(n10136), .Z(c[2241]) );
  XNOR U11993 ( .A(a[2241]), .B(n10137), .Z(n10136) );
  IV U11994 ( .A(n10134), .Z(n10137) );
  XOR U11995 ( .A(n10138), .B(n10139), .Z(n10134) );
  ANDN U11996 ( .B(n10140), .A(n10141), .Z(n10138) );
  XNOR U11997 ( .A(b[2240]), .B(n10139), .Z(n10140) );
  XNOR U11998 ( .A(b[2240]), .B(n10141), .Z(c[2240]) );
  XNOR U11999 ( .A(a[2240]), .B(n10142), .Z(n10141) );
  IV U12000 ( .A(n10139), .Z(n10142) );
  XOR U12001 ( .A(n10143), .B(n10144), .Z(n10139) );
  ANDN U12002 ( .B(n10145), .A(n10146), .Z(n10143) );
  XNOR U12003 ( .A(b[2239]), .B(n10144), .Z(n10145) );
  XNOR U12004 ( .A(b[223]), .B(n10147), .Z(c[223]) );
  XNOR U12005 ( .A(b[2239]), .B(n10146), .Z(c[2239]) );
  XNOR U12006 ( .A(a[2239]), .B(n10148), .Z(n10146) );
  IV U12007 ( .A(n10144), .Z(n10148) );
  XOR U12008 ( .A(n10149), .B(n10150), .Z(n10144) );
  ANDN U12009 ( .B(n10151), .A(n10152), .Z(n10149) );
  XNOR U12010 ( .A(b[2238]), .B(n10150), .Z(n10151) );
  XNOR U12011 ( .A(b[2238]), .B(n10152), .Z(c[2238]) );
  XNOR U12012 ( .A(a[2238]), .B(n10153), .Z(n10152) );
  IV U12013 ( .A(n10150), .Z(n10153) );
  XOR U12014 ( .A(n10154), .B(n10155), .Z(n10150) );
  ANDN U12015 ( .B(n10156), .A(n10157), .Z(n10154) );
  XNOR U12016 ( .A(b[2237]), .B(n10155), .Z(n10156) );
  XNOR U12017 ( .A(b[2237]), .B(n10157), .Z(c[2237]) );
  XNOR U12018 ( .A(a[2237]), .B(n10158), .Z(n10157) );
  IV U12019 ( .A(n10155), .Z(n10158) );
  XOR U12020 ( .A(n10159), .B(n10160), .Z(n10155) );
  ANDN U12021 ( .B(n10161), .A(n10162), .Z(n10159) );
  XNOR U12022 ( .A(b[2236]), .B(n10160), .Z(n10161) );
  XNOR U12023 ( .A(b[2236]), .B(n10162), .Z(c[2236]) );
  XNOR U12024 ( .A(a[2236]), .B(n10163), .Z(n10162) );
  IV U12025 ( .A(n10160), .Z(n10163) );
  XOR U12026 ( .A(n10164), .B(n10165), .Z(n10160) );
  ANDN U12027 ( .B(n10166), .A(n10167), .Z(n10164) );
  XNOR U12028 ( .A(b[2235]), .B(n10165), .Z(n10166) );
  XNOR U12029 ( .A(b[2235]), .B(n10167), .Z(c[2235]) );
  XNOR U12030 ( .A(a[2235]), .B(n10168), .Z(n10167) );
  IV U12031 ( .A(n10165), .Z(n10168) );
  XOR U12032 ( .A(n10169), .B(n10170), .Z(n10165) );
  ANDN U12033 ( .B(n10171), .A(n10172), .Z(n10169) );
  XNOR U12034 ( .A(b[2234]), .B(n10170), .Z(n10171) );
  XNOR U12035 ( .A(b[2234]), .B(n10172), .Z(c[2234]) );
  XNOR U12036 ( .A(a[2234]), .B(n10173), .Z(n10172) );
  IV U12037 ( .A(n10170), .Z(n10173) );
  XOR U12038 ( .A(n10174), .B(n10175), .Z(n10170) );
  ANDN U12039 ( .B(n10176), .A(n10177), .Z(n10174) );
  XNOR U12040 ( .A(b[2233]), .B(n10175), .Z(n10176) );
  XNOR U12041 ( .A(b[2233]), .B(n10177), .Z(c[2233]) );
  XNOR U12042 ( .A(a[2233]), .B(n10178), .Z(n10177) );
  IV U12043 ( .A(n10175), .Z(n10178) );
  XOR U12044 ( .A(n10179), .B(n10180), .Z(n10175) );
  ANDN U12045 ( .B(n10181), .A(n10182), .Z(n10179) );
  XNOR U12046 ( .A(b[2232]), .B(n10180), .Z(n10181) );
  XNOR U12047 ( .A(b[2232]), .B(n10182), .Z(c[2232]) );
  XNOR U12048 ( .A(a[2232]), .B(n10183), .Z(n10182) );
  IV U12049 ( .A(n10180), .Z(n10183) );
  XOR U12050 ( .A(n10184), .B(n10185), .Z(n10180) );
  ANDN U12051 ( .B(n10186), .A(n10187), .Z(n10184) );
  XNOR U12052 ( .A(b[2231]), .B(n10185), .Z(n10186) );
  XNOR U12053 ( .A(b[2231]), .B(n10187), .Z(c[2231]) );
  XNOR U12054 ( .A(a[2231]), .B(n10188), .Z(n10187) );
  IV U12055 ( .A(n10185), .Z(n10188) );
  XOR U12056 ( .A(n10189), .B(n10190), .Z(n10185) );
  ANDN U12057 ( .B(n10191), .A(n10192), .Z(n10189) );
  XNOR U12058 ( .A(b[2230]), .B(n10190), .Z(n10191) );
  XNOR U12059 ( .A(b[2230]), .B(n10192), .Z(c[2230]) );
  XNOR U12060 ( .A(a[2230]), .B(n10193), .Z(n10192) );
  IV U12061 ( .A(n10190), .Z(n10193) );
  XOR U12062 ( .A(n10194), .B(n10195), .Z(n10190) );
  ANDN U12063 ( .B(n10196), .A(n10197), .Z(n10194) );
  XNOR U12064 ( .A(b[2229]), .B(n10195), .Z(n10196) );
  XNOR U12065 ( .A(b[222]), .B(n10198), .Z(c[222]) );
  XNOR U12066 ( .A(b[2229]), .B(n10197), .Z(c[2229]) );
  XNOR U12067 ( .A(a[2229]), .B(n10199), .Z(n10197) );
  IV U12068 ( .A(n10195), .Z(n10199) );
  XOR U12069 ( .A(n10200), .B(n10201), .Z(n10195) );
  ANDN U12070 ( .B(n10202), .A(n10203), .Z(n10200) );
  XNOR U12071 ( .A(b[2228]), .B(n10201), .Z(n10202) );
  XNOR U12072 ( .A(b[2228]), .B(n10203), .Z(c[2228]) );
  XNOR U12073 ( .A(a[2228]), .B(n10204), .Z(n10203) );
  IV U12074 ( .A(n10201), .Z(n10204) );
  XOR U12075 ( .A(n10205), .B(n10206), .Z(n10201) );
  ANDN U12076 ( .B(n10207), .A(n10208), .Z(n10205) );
  XNOR U12077 ( .A(b[2227]), .B(n10206), .Z(n10207) );
  XNOR U12078 ( .A(b[2227]), .B(n10208), .Z(c[2227]) );
  XNOR U12079 ( .A(a[2227]), .B(n10209), .Z(n10208) );
  IV U12080 ( .A(n10206), .Z(n10209) );
  XOR U12081 ( .A(n10210), .B(n10211), .Z(n10206) );
  ANDN U12082 ( .B(n10212), .A(n10213), .Z(n10210) );
  XNOR U12083 ( .A(b[2226]), .B(n10211), .Z(n10212) );
  XNOR U12084 ( .A(b[2226]), .B(n10213), .Z(c[2226]) );
  XNOR U12085 ( .A(a[2226]), .B(n10214), .Z(n10213) );
  IV U12086 ( .A(n10211), .Z(n10214) );
  XOR U12087 ( .A(n10215), .B(n10216), .Z(n10211) );
  ANDN U12088 ( .B(n10217), .A(n10218), .Z(n10215) );
  XNOR U12089 ( .A(b[2225]), .B(n10216), .Z(n10217) );
  XNOR U12090 ( .A(b[2225]), .B(n10218), .Z(c[2225]) );
  XNOR U12091 ( .A(a[2225]), .B(n10219), .Z(n10218) );
  IV U12092 ( .A(n10216), .Z(n10219) );
  XOR U12093 ( .A(n10220), .B(n10221), .Z(n10216) );
  ANDN U12094 ( .B(n10222), .A(n10223), .Z(n10220) );
  XNOR U12095 ( .A(b[2224]), .B(n10221), .Z(n10222) );
  XNOR U12096 ( .A(b[2224]), .B(n10223), .Z(c[2224]) );
  XNOR U12097 ( .A(a[2224]), .B(n10224), .Z(n10223) );
  IV U12098 ( .A(n10221), .Z(n10224) );
  XOR U12099 ( .A(n10225), .B(n10226), .Z(n10221) );
  ANDN U12100 ( .B(n10227), .A(n10228), .Z(n10225) );
  XNOR U12101 ( .A(b[2223]), .B(n10226), .Z(n10227) );
  XNOR U12102 ( .A(b[2223]), .B(n10228), .Z(c[2223]) );
  XNOR U12103 ( .A(a[2223]), .B(n10229), .Z(n10228) );
  IV U12104 ( .A(n10226), .Z(n10229) );
  XOR U12105 ( .A(n10230), .B(n10231), .Z(n10226) );
  ANDN U12106 ( .B(n10232), .A(n10233), .Z(n10230) );
  XNOR U12107 ( .A(b[2222]), .B(n10231), .Z(n10232) );
  XNOR U12108 ( .A(b[2222]), .B(n10233), .Z(c[2222]) );
  XNOR U12109 ( .A(a[2222]), .B(n10234), .Z(n10233) );
  IV U12110 ( .A(n10231), .Z(n10234) );
  XOR U12111 ( .A(n10235), .B(n10236), .Z(n10231) );
  ANDN U12112 ( .B(n10237), .A(n10238), .Z(n10235) );
  XNOR U12113 ( .A(b[2221]), .B(n10236), .Z(n10237) );
  XNOR U12114 ( .A(b[2221]), .B(n10238), .Z(c[2221]) );
  XNOR U12115 ( .A(a[2221]), .B(n10239), .Z(n10238) );
  IV U12116 ( .A(n10236), .Z(n10239) );
  XOR U12117 ( .A(n10240), .B(n10241), .Z(n10236) );
  ANDN U12118 ( .B(n10242), .A(n10243), .Z(n10240) );
  XNOR U12119 ( .A(b[2220]), .B(n10241), .Z(n10242) );
  XNOR U12120 ( .A(b[2220]), .B(n10243), .Z(c[2220]) );
  XNOR U12121 ( .A(a[2220]), .B(n10244), .Z(n10243) );
  IV U12122 ( .A(n10241), .Z(n10244) );
  XOR U12123 ( .A(n10245), .B(n10246), .Z(n10241) );
  ANDN U12124 ( .B(n10247), .A(n10248), .Z(n10245) );
  XNOR U12125 ( .A(b[2219]), .B(n10246), .Z(n10247) );
  XNOR U12126 ( .A(b[221]), .B(n10249), .Z(c[221]) );
  XNOR U12127 ( .A(b[2219]), .B(n10248), .Z(c[2219]) );
  XNOR U12128 ( .A(a[2219]), .B(n10250), .Z(n10248) );
  IV U12129 ( .A(n10246), .Z(n10250) );
  XOR U12130 ( .A(n10251), .B(n10252), .Z(n10246) );
  ANDN U12131 ( .B(n10253), .A(n10254), .Z(n10251) );
  XNOR U12132 ( .A(b[2218]), .B(n10252), .Z(n10253) );
  XNOR U12133 ( .A(b[2218]), .B(n10254), .Z(c[2218]) );
  XNOR U12134 ( .A(a[2218]), .B(n10255), .Z(n10254) );
  IV U12135 ( .A(n10252), .Z(n10255) );
  XOR U12136 ( .A(n10256), .B(n10257), .Z(n10252) );
  ANDN U12137 ( .B(n10258), .A(n10259), .Z(n10256) );
  XNOR U12138 ( .A(b[2217]), .B(n10257), .Z(n10258) );
  XNOR U12139 ( .A(b[2217]), .B(n10259), .Z(c[2217]) );
  XNOR U12140 ( .A(a[2217]), .B(n10260), .Z(n10259) );
  IV U12141 ( .A(n10257), .Z(n10260) );
  XOR U12142 ( .A(n10261), .B(n10262), .Z(n10257) );
  ANDN U12143 ( .B(n10263), .A(n10264), .Z(n10261) );
  XNOR U12144 ( .A(b[2216]), .B(n10262), .Z(n10263) );
  XNOR U12145 ( .A(b[2216]), .B(n10264), .Z(c[2216]) );
  XNOR U12146 ( .A(a[2216]), .B(n10265), .Z(n10264) );
  IV U12147 ( .A(n10262), .Z(n10265) );
  XOR U12148 ( .A(n10266), .B(n10267), .Z(n10262) );
  ANDN U12149 ( .B(n10268), .A(n10269), .Z(n10266) );
  XNOR U12150 ( .A(b[2215]), .B(n10267), .Z(n10268) );
  XNOR U12151 ( .A(b[2215]), .B(n10269), .Z(c[2215]) );
  XNOR U12152 ( .A(a[2215]), .B(n10270), .Z(n10269) );
  IV U12153 ( .A(n10267), .Z(n10270) );
  XOR U12154 ( .A(n10271), .B(n10272), .Z(n10267) );
  ANDN U12155 ( .B(n10273), .A(n10274), .Z(n10271) );
  XNOR U12156 ( .A(b[2214]), .B(n10272), .Z(n10273) );
  XNOR U12157 ( .A(b[2214]), .B(n10274), .Z(c[2214]) );
  XNOR U12158 ( .A(a[2214]), .B(n10275), .Z(n10274) );
  IV U12159 ( .A(n10272), .Z(n10275) );
  XOR U12160 ( .A(n10276), .B(n10277), .Z(n10272) );
  ANDN U12161 ( .B(n10278), .A(n10279), .Z(n10276) );
  XNOR U12162 ( .A(b[2213]), .B(n10277), .Z(n10278) );
  XNOR U12163 ( .A(b[2213]), .B(n10279), .Z(c[2213]) );
  XNOR U12164 ( .A(a[2213]), .B(n10280), .Z(n10279) );
  IV U12165 ( .A(n10277), .Z(n10280) );
  XOR U12166 ( .A(n10281), .B(n10282), .Z(n10277) );
  ANDN U12167 ( .B(n10283), .A(n10284), .Z(n10281) );
  XNOR U12168 ( .A(b[2212]), .B(n10282), .Z(n10283) );
  XNOR U12169 ( .A(b[2212]), .B(n10284), .Z(c[2212]) );
  XNOR U12170 ( .A(a[2212]), .B(n10285), .Z(n10284) );
  IV U12171 ( .A(n10282), .Z(n10285) );
  XOR U12172 ( .A(n10286), .B(n10287), .Z(n10282) );
  ANDN U12173 ( .B(n10288), .A(n10289), .Z(n10286) );
  XNOR U12174 ( .A(b[2211]), .B(n10287), .Z(n10288) );
  XNOR U12175 ( .A(b[2211]), .B(n10289), .Z(c[2211]) );
  XNOR U12176 ( .A(a[2211]), .B(n10290), .Z(n10289) );
  IV U12177 ( .A(n10287), .Z(n10290) );
  XOR U12178 ( .A(n10291), .B(n10292), .Z(n10287) );
  ANDN U12179 ( .B(n10293), .A(n10294), .Z(n10291) );
  XNOR U12180 ( .A(b[2210]), .B(n10292), .Z(n10293) );
  XNOR U12181 ( .A(b[2210]), .B(n10294), .Z(c[2210]) );
  XNOR U12182 ( .A(a[2210]), .B(n10295), .Z(n10294) );
  IV U12183 ( .A(n10292), .Z(n10295) );
  XOR U12184 ( .A(n10296), .B(n10297), .Z(n10292) );
  ANDN U12185 ( .B(n10298), .A(n10299), .Z(n10296) );
  XNOR U12186 ( .A(b[2209]), .B(n10297), .Z(n10298) );
  XNOR U12187 ( .A(b[220]), .B(n10300), .Z(c[220]) );
  XNOR U12188 ( .A(b[2209]), .B(n10299), .Z(c[2209]) );
  XNOR U12189 ( .A(a[2209]), .B(n10301), .Z(n10299) );
  IV U12190 ( .A(n10297), .Z(n10301) );
  XOR U12191 ( .A(n10302), .B(n10303), .Z(n10297) );
  ANDN U12192 ( .B(n10304), .A(n10305), .Z(n10302) );
  XNOR U12193 ( .A(b[2208]), .B(n10303), .Z(n10304) );
  XNOR U12194 ( .A(b[2208]), .B(n10305), .Z(c[2208]) );
  XNOR U12195 ( .A(a[2208]), .B(n10306), .Z(n10305) );
  IV U12196 ( .A(n10303), .Z(n10306) );
  XOR U12197 ( .A(n10307), .B(n10308), .Z(n10303) );
  ANDN U12198 ( .B(n10309), .A(n10310), .Z(n10307) );
  XNOR U12199 ( .A(b[2207]), .B(n10308), .Z(n10309) );
  XNOR U12200 ( .A(b[2207]), .B(n10310), .Z(c[2207]) );
  XNOR U12201 ( .A(a[2207]), .B(n10311), .Z(n10310) );
  IV U12202 ( .A(n10308), .Z(n10311) );
  XOR U12203 ( .A(n10312), .B(n10313), .Z(n10308) );
  ANDN U12204 ( .B(n10314), .A(n10315), .Z(n10312) );
  XNOR U12205 ( .A(b[2206]), .B(n10313), .Z(n10314) );
  XNOR U12206 ( .A(b[2206]), .B(n10315), .Z(c[2206]) );
  XNOR U12207 ( .A(a[2206]), .B(n10316), .Z(n10315) );
  IV U12208 ( .A(n10313), .Z(n10316) );
  XOR U12209 ( .A(n10317), .B(n10318), .Z(n10313) );
  ANDN U12210 ( .B(n10319), .A(n10320), .Z(n10317) );
  XNOR U12211 ( .A(b[2205]), .B(n10318), .Z(n10319) );
  XNOR U12212 ( .A(b[2205]), .B(n10320), .Z(c[2205]) );
  XNOR U12213 ( .A(a[2205]), .B(n10321), .Z(n10320) );
  IV U12214 ( .A(n10318), .Z(n10321) );
  XOR U12215 ( .A(n10322), .B(n10323), .Z(n10318) );
  ANDN U12216 ( .B(n10324), .A(n10325), .Z(n10322) );
  XNOR U12217 ( .A(b[2204]), .B(n10323), .Z(n10324) );
  XNOR U12218 ( .A(b[2204]), .B(n10325), .Z(c[2204]) );
  XNOR U12219 ( .A(a[2204]), .B(n10326), .Z(n10325) );
  IV U12220 ( .A(n10323), .Z(n10326) );
  XOR U12221 ( .A(n10327), .B(n10328), .Z(n10323) );
  ANDN U12222 ( .B(n10329), .A(n10330), .Z(n10327) );
  XNOR U12223 ( .A(b[2203]), .B(n10328), .Z(n10329) );
  XNOR U12224 ( .A(b[2203]), .B(n10330), .Z(c[2203]) );
  XNOR U12225 ( .A(a[2203]), .B(n10331), .Z(n10330) );
  IV U12226 ( .A(n10328), .Z(n10331) );
  XOR U12227 ( .A(n10332), .B(n10333), .Z(n10328) );
  ANDN U12228 ( .B(n10334), .A(n10335), .Z(n10332) );
  XNOR U12229 ( .A(b[2202]), .B(n10333), .Z(n10334) );
  XNOR U12230 ( .A(b[2202]), .B(n10335), .Z(c[2202]) );
  XNOR U12231 ( .A(a[2202]), .B(n10336), .Z(n10335) );
  IV U12232 ( .A(n10333), .Z(n10336) );
  XOR U12233 ( .A(n10337), .B(n10338), .Z(n10333) );
  ANDN U12234 ( .B(n10339), .A(n10340), .Z(n10337) );
  XNOR U12235 ( .A(b[2201]), .B(n10338), .Z(n10339) );
  XNOR U12236 ( .A(b[2201]), .B(n10340), .Z(c[2201]) );
  XNOR U12237 ( .A(a[2201]), .B(n10341), .Z(n10340) );
  IV U12238 ( .A(n10338), .Z(n10341) );
  XOR U12239 ( .A(n10342), .B(n10343), .Z(n10338) );
  ANDN U12240 ( .B(n10344), .A(n10345), .Z(n10342) );
  XNOR U12241 ( .A(b[2200]), .B(n10343), .Z(n10344) );
  XNOR U12242 ( .A(b[2200]), .B(n10345), .Z(c[2200]) );
  XNOR U12243 ( .A(a[2200]), .B(n10346), .Z(n10345) );
  IV U12244 ( .A(n10343), .Z(n10346) );
  XOR U12245 ( .A(n10347), .B(n10348), .Z(n10343) );
  ANDN U12246 ( .B(n10349), .A(n10350), .Z(n10347) );
  XNOR U12247 ( .A(b[2199]), .B(n10348), .Z(n10349) );
  XNOR U12248 ( .A(b[21]), .B(n10351), .Z(c[21]) );
  XNOR U12249 ( .A(b[219]), .B(n10352), .Z(c[219]) );
  XNOR U12250 ( .A(b[2199]), .B(n10350), .Z(c[2199]) );
  XNOR U12251 ( .A(a[2199]), .B(n10353), .Z(n10350) );
  IV U12252 ( .A(n10348), .Z(n10353) );
  XOR U12253 ( .A(n10354), .B(n10355), .Z(n10348) );
  ANDN U12254 ( .B(n10356), .A(n10357), .Z(n10354) );
  XNOR U12255 ( .A(b[2198]), .B(n10355), .Z(n10356) );
  XNOR U12256 ( .A(b[2198]), .B(n10357), .Z(c[2198]) );
  XNOR U12257 ( .A(a[2198]), .B(n10358), .Z(n10357) );
  IV U12258 ( .A(n10355), .Z(n10358) );
  XOR U12259 ( .A(n10359), .B(n10360), .Z(n10355) );
  ANDN U12260 ( .B(n10361), .A(n10362), .Z(n10359) );
  XNOR U12261 ( .A(b[2197]), .B(n10360), .Z(n10361) );
  XNOR U12262 ( .A(b[2197]), .B(n10362), .Z(c[2197]) );
  XNOR U12263 ( .A(a[2197]), .B(n10363), .Z(n10362) );
  IV U12264 ( .A(n10360), .Z(n10363) );
  XOR U12265 ( .A(n10364), .B(n10365), .Z(n10360) );
  ANDN U12266 ( .B(n10366), .A(n10367), .Z(n10364) );
  XNOR U12267 ( .A(b[2196]), .B(n10365), .Z(n10366) );
  XNOR U12268 ( .A(b[2196]), .B(n10367), .Z(c[2196]) );
  XNOR U12269 ( .A(a[2196]), .B(n10368), .Z(n10367) );
  IV U12270 ( .A(n10365), .Z(n10368) );
  XOR U12271 ( .A(n10369), .B(n10370), .Z(n10365) );
  ANDN U12272 ( .B(n10371), .A(n10372), .Z(n10369) );
  XNOR U12273 ( .A(b[2195]), .B(n10370), .Z(n10371) );
  XNOR U12274 ( .A(b[2195]), .B(n10372), .Z(c[2195]) );
  XNOR U12275 ( .A(a[2195]), .B(n10373), .Z(n10372) );
  IV U12276 ( .A(n10370), .Z(n10373) );
  XOR U12277 ( .A(n10374), .B(n10375), .Z(n10370) );
  ANDN U12278 ( .B(n10376), .A(n10377), .Z(n10374) );
  XNOR U12279 ( .A(b[2194]), .B(n10375), .Z(n10376) );
  XNOR U12280 ( .A(b[2194]), .B(n10377), .Z(c[2194]) );
  XNOR U12281 ( .A(a[2194]), .B(n10378), .Z(n10377) );
  IV U12282 ( .A(n10375), .Z(n10378) );
  XOR U12283 ( .A(n10379), .B(n10380), .Z(n10375) );
  ANDN U12284 ( .B(n10381), .A(n10382), .Z(n10379) );
  XNOR U12285 ( .A(b[2193]), .B(n10380), .Z(n10381) );
  XNOR U12286 ( .A(b[2193]), .B(n10382), .Z(c[2193]) );
  XNOR U12287 ( .A(a[2193]), .B(n10383), .Z(n10382) );
  IV U12288 ( .A(n10380), .Z(n10383) );
  XOR U12289 ( .A(n10384), .B(n10385), .Z(n10380) );
  ANDN U12290 ( .B(n10386), .A(n10387), .Z(n10384) );
  XNOR U12291 ( .A(b[2192]), .B(n10385), .Z(n10386) );
  XNOR U12292 ( .A(b[2192]), .B(n10387), .Z(c[2192]) );
  XNOR U12293 ( .A(a[2192]), .B(n10388), .Z(n10387) );
  IV U12294 ( .A(n10385), .Z(n10388) );
  XOR U12295 ( .A(n10389), .B(n10390), .Z(n10385) );
  ANDN U12296 ( .B(n10391), .A(n10392), .Z(n10389) );
  XNOR U12297 ( .A(b[2191]), .B(n10390), .Z(n10391) );
  XNOR U12298 ( .A(b[2191]), .B(n10392), .Z(c[2191]) );
  XNOR U12299 ( .A(a[2191]), .B(n10393), .Z(n10392) );
  IV U12300 ( .A(n10390), .Z(n10393) );
  XOR U12301 ( .A(n10394), .B(n10395), .Z(n10390) );
  ANDN U12302 ( .B(n10396), .A(n10397), .Z(n10394) );
  XNOR U12303 ( .A(b[2190]), .B(n10395), .Z(n10396) );
  XNOR U12304 ( .A(b[2190]), .B(n10397), .Z(c[2190]) );
  XNOR U12305 ( .A(a[2190]), .B(n10398), .Z(n10397) );
  IV U12306 ( .A(n10395), .Z(n10398) );
  XOR U12307 ( .A(n10399), .B(n10400), .Z(n10395) );
  ANDN U12308 ( .B(n10401), .A(n10402), .Z(n10399) );
  XNOR U12309 ( .A(b[2189]), .B(n10400), .Z(n10401) );
  XNOR U12310 ( .A(b[218]), .B(n10403), .Z(c[218]) );
  XNOR U12311 ( .A(b[2189]), .B(n10402), .Z(c[2189]) );
  XNOR U12312 ( .A(a[2189]), .B(n10404), .Z(n10402) );
  IV U12313 ( .A(n10400), .Z(n10404) );
  XOR U12314 ( .A(n10405), .B(n10406), .Z(n10400) );
  ANDN U12315 ( .B(n10407), .A(n10408), .Z(n10405) );
  XNOR U12316 ( .A(b[2188]), .B(n10406), .Z(n10407) );
  XNOR U12317 ( .A(b[2188]), .B(n10408), .Z(c[2188]) );
  XNOR U12318 ( .A(a[2188]), .B(n10409), .Z(n10408) );
  IV U12319 ( .A(n10406), .Z(n10409) );
  XOR U12320 ( .A(n10410), .B(n10411), .Z(n10406) );
  ANDN U12321 ( .B(n10412), .A(n10413), .Z(n10410) );
  XNOR U12322 ( .A(b[2187]), .B(n10411), .Z(n10412) );
  XNOR U12323 ( .A(b[2187]), .B(n10413), .Z(c[2187]) );
  XNOR U12324 ( .A(a[2187]), .B(n10414), .Z(n10413) );
  IV U12325 ( .A(n10411), .Z(n10414) );
  XOR U12326 ( .A(n10415), .B(n10416), .Z(n10411) );
  ANDN U12327 ( .B(n10417), .A(n10418), .Z(n10415) );
  XNOR U12328 ( .A(b[2186]), .B(n10416), .Z(n10417) );
  XNOR U12329 ( .A(b[2186]), .B(n10418), .Z(c[2186]) );
  XNOR U12330 ( .A(a[2186]), .B(n10419), .Z(n10418) );
  IV U12331 ( .A(n10416), .Z(n10419) );
  XOR U12332 ( .A(n10420), .B(n10421), .Z(n10416) );
  ANDN U12333 ( .B(n10422), .A(n10423), .Z(n10420) );
  XNOR U12334 ( .A(b[2185]), .B(n10421), .Z(n10422) );
  XNOR U12335 ( .A(b[2185]), .B(n10423), .Z(c[2185]) );
  XNOR U12336 ( .A(a[2185]), .B(n10424), .Z(n10423) );
  IV U12337 ( .A(n10421), .Z(n10424) );
  XOR U12338 ( .A(n10425), .B(n10426), .Z(n10421) );
  ANDN U12339 ( .B(n10427), .A(n10428), .Z(n10425) );
  XNOR U12340 ( .A(b[2184]), .B(n10426), .Z(n10427) );
  XNOR U12341 ( .A(b[2184]), .B(n10428), .Z(c[2184]) );
  XNOR U12342 ( .A(a[2184]), .B(n10429), .Z(n10428) );
  IV U12343 ( .A(n10426), .Z(n10429) );
  XOR U12344 ( .A(n10430), .B(n10431), .Z(n10426) );
  ANDN U12345 ( .B(n10432), .A(n10433), .Z(n10430) );
  XNOR U12346 ( .A(b[2183]), .B(n10431), .Z(n10432) );
  XNOR U12347 ( .A(b[2183]), .B(n10433), .Z(c[2183]) );
  XNOR U12348 ( .A(a[2183]), .B(n10434), .Z(n10433) );
  IV U12349 ( .A(n10431), .Z(n10434) );
  XOR U12350 ( .A(n10435), .B(n10436), .Z(n10431) );
  ANDN U12351 ( .B(n10437), .A(n10438), .Z(n10435) );
  XNOR U12352 ( .A(b[2182]), .B(n10436), .Z(n10437) );
  XNOR U12353 ( .A(b[2182]), .B(n10438), .Z(c[2182]) );
  XNOR U12354 ( .A(a[2182]), .B(n10439), .Z(n10438) );
  IV U12355 ( .A(n10436), .Z(n10439) );
  XOR U12356 ( .A(n10440), .B(n10441), .Z(n10436) );
  ANDN U12357 ( .B(n10442), .A(n10443), .Z(n10440) );
  XNOR U12358 ( .A(b[2181]), .B(n10441), .Z(n10442) );
  XNOR U12359 ( .A(b[2181]), .B(n10443), .Z(c[2181]) );
  XNOR U12360 ( .A(a[2181]), .B(n10444), .Z(n10443) );
  IV U12361 ( .A(n10441), .Z(n10444) );
  XOR U12362 ( .A(n10445), .B(n10446), .Z(n10441) );
  ANDN U12363 ( .B(n10447), .A(n10448), .Z(n10445) );
  XNOR U12364 ( .A(b[2180]), .B(n10446), .Z(n10447) );
  XNOR U12365 ( .A(b[2180]), .B(n10448), .Z(c[2180]) );
  XNOR U12366 ( .A(a[2180]), .B(n10449), .Z(n10448) );
  IV U12367 ( .A(n10446), .Z(n10449) );
  XOR U12368 ( .A(n10450), .B(n10451), .Z(n10446) );
  ANDN U12369 ( .B(n10452), .A(n10453), .Z(n10450) );
  XNOR U12370 ( .A(b[2179]), .B(n10451), .Z(n10452) );
  XNOR U12371 ( .A(b[217]), .B(n10454), .Z(c[217]) );
  XNOR U12372 ( .A(b[2179]), .B(n10453), .Z(c[2179]) );
  XNOR U12373 ( .A(a[2179]), .B(n10455), .Z(n10453) );
  IV U12374 ( .A(n10451), .Z(n10455) );
  XOR U12375 ( .A(n10456), .B(n10457), .Z(n10451) );
  ANDN U12376 ( .B(n10458), .A(n10459), .Z(n10456) );
  XNOR U12377 ( .A(b[2178]), .B(n10457), .Z(n10458) );
  XNOR U12378 ( .A(b[2178]), .B(n10459), .Z(c[2178]) );
  XNOR U12379 ( .A(a[2178]), .B(n10460), .Z(n10459) );
  IV U12380 ( .A(n10457), .Z(n10460) );
  XOR U12381 ( .A(n10461), .B(n10462), .Z(n10457) );
  ANDN U12382 ( .B(n10463), .A(n10464), .Z(n10461) );
  XNOR U12383 ( .A(b[2177]), .B(n10462), .Z(n10463) );
  XNOR U12384 ( .A(b[2177]), .B(n10464), .Z(c[2177]) );
  XNOR U12385 ( .A(a[2177]), .B(n10465), .Z(n10464) );
  IV U12386 ( .A(n10462), .Z(n10465) );
  XOR U12387 ( .A(n10466), .B(n10467), .Z(n10462) );
  ANDN U12388 ( .B(n10468), .A(n10469), .Z(n10466) );
  XNOR U12389 ( .A(b[2176]), .B(n10467), .Z(n10468) );
  XNOR U12390 ( .A(b[2176]), .B(n10469), .Z(c[2176]) );
  XNOR U12391 ( .A(a[2176]), .B(n10470), .Z(n10469) );
  IV U12392 ( .A(n10467), .Z(n10470) );
  XOR U12393 ( .A(n10471), .B(n10472), .Z(n10467) );
  ANDN U12394 ( .B(n10473), .A(n10474), .Z(n10471) );
  XNOR U12395 ( .A(b[2175]), .B(n10472), .Z(n10473) );
  XNOR U12396 ( .A(b[2175]), .B(n10474), .Z(c[2175]) );
  XNOR U12397 ( .A(a[2175]), .B(n10475), .Z(n10474) );
  IV U12398 ( .A(n10472), .Z(n10475) );
  XOR U12399 ( .A(n10476), .B(n10477), .Z(n10472) );
  ANDN U12400 ( .B(n10478), .A(n10479), .Z(n10476) );
  XNOR U12401 ( .A(b[2174]), .B(n10477), .Z(n10478) );
  XNOR U12402 ( .A(b[2174]), .B(n10479), .Z(c[2174]) );
  XNOR U12403 ( .A(a[2174]), .B(n10480), .Z(n10479) );
  IV U12404 ( .A(n10477), .Z(n10480) );
  XOR U12405 ( .A(n10481), .B(n10482), .Z(n10477) );
  ANDN U12406 ( .B(n10483), .A(n10484), .Z(n10481) );
  XNOR U12407 ( .A(b[2173]), .B(n10482), .Z(n10483) );
  XNOR U12408 ( .A(b[2173]), .B(n10484), .Z(c[2173]) );
  XNOR U12409 ( .A(a[2173]), .B(n10485), .Z(n10484) );
  IV U12410 ( .A(n10482), .Z(n10485) );
  XOR U12411 ( .A(n10486), .B(n10487), .Z(n10482) );
  ANDN U12412 ( .B(n10488), .A(n10489), .Z(n10486) );
  XNOR U12413 ( .A(b[2172]), .B(n10487), .Z(n10488) );
  XNOR U12414 ( .A(b[2172]), .B(n10489), .Z(c[2172]) );
  XNOR U12415 ( .A(a[2172]), .B(n10490), .Z(n10489) );
  IV U12416 ( .A(n10487), .Z(n10490) );
  XOR U12417 ( .A(n10491), .B(n10492), .Z(n10487) );
  ANDN U12418 ( .B(n10493), .A(n10494), .Z(n10491) );
  XNOR U12419 ( .A(b[2171]), .B(n10492), .Z(n10493) );
  XNOR U12420 ( .A(b[2171]), .B(n10494), .Z(c[2171]) );
  XNOR U12421 ( .A(a[2171]), .B(n10495), .Z(n10494) );
  IV U12422 ( .A(n10492), .Z(n10495) );
  XOR U12423 ( .A(n10496), .B(n10497), .Z(n10492) );
  ANDN U12424 ( .B(n10498), .A(n10499), .Z(n10496) );
  XNOR U12425 ( .A(b[2170]), .B(n10497), .Z(n10498) );
  XNOR U12426 ( .A(b[2170]), .B(n10499), .Z(c[2170]) );
  XNOR U12427 ( .A(a[2170]), .B(n10500), .Z(n10499) );
  IV U12428 ( .A(n10497), .Z(n10500) );
  XOR U12429 ( .A(n10501), .B(n10502), .Z(n10497) );
  ANDN U12430 ( .B(n10503), .A(n10504), .Z(n10501) );
  XNOR U12431 ( .A(b[2169]), .B(n10502), .Z(n10503) );
  XNOR U12432 ( .A(b[216]), .B(n10505), .Z(c[216]) );
  XNOR U12433 ( .A(b[2169]), .B(n10504), .Z(c[2169]) );
  XNOR U12434 ( .A(a[2169]), .B(n10506), .Z(n10504) );
  IV U12435 ( .A(n10502), .Z(n10506) );
  XOR U12436 ( .A(n10507), .B(n10508), .Z(n10502) );
  ANDN U12437 ( .B(n10509), .A(n10510), .Z(n10507) );
  XNOR U12438 ( .A(b[2168]), .B(n10508), .Z(n10509) );
  XNOR U12439 ( .A(b[2168]), .B(n10510), .Z(c[2168]) );
  XNOR U12440 ( .A(a[2168]), .B(n10511), .Z(n10510) );
  IV U12441 ( .A(n10508), .Z(n10511) );
  XOR U12442 ( .A(n10512), .B(n10513), .Z(n10508) );
  ANDN U12443 ( .B(n10514), .A(n10515), .Z(n10512) );
  XNOR U12444 ( .A(b[2167]), .B(n10513), .Z(n10514) );
  XNOR U12445 ( .A(b[2167]), .B(n10515), .Z(c[2167]) );
  XNOR U12446 ( .A(a[2167]), .B(n10516), .Z(n10515) );
  IV U12447 ( .A(n10513), .Z(n10516) );
  XOR U12448 ( .A(n10517), .B(n10518), .Z(n10513) );
  ANDN U12449 ( .B(n10519), .A(n10520), .Z(n10517) );
  XNOR U12450 ( .A(b[2166]), .B(n10518), .Z(n10519) );
  XNOR U12451 ( .A(b[2166]), .B(n10520), .Z(c[2166]) );
  XNOR U12452 ( .A(a[2166]), .B(n10521), .Z(n10520) );
  IV U12453 ( .A(n10518), .Z(n10521) );
  XOR U12454 ( .A(n10522), .B(n10523), .Z(n10518) );
  ANDN U12455 ( .B(n10524), .A(n10525), .Z(n10522) );
  XNOR U12456 ( .A(b[2165]), .B(n10523), .Z(n10524) );
  XNOR U12457 ( .A(b[2165]), .B(n10525), .Z(c[2165]) );
  XNOR U12458 ( .A(a[2165]), .B(n10526), .Z(n10525) );
  IV U12459 ( .A(n10523), .Z(n10526) );
  XOR U12460 ( .A(n10527), .B(n10528), .Z(n10523) );
  ANDN U12461 ( .B(n10529), .A(n10530), .Z(n10527) );
  XNOR U12462 ( .A(b[2164]), .B(n10528), .Z(n10529) );
  XNOR U12463 ( .A(b[2164]), .B(n10530), .Z(c[2164]) );
  XNOR U12464 ( .A(a[2164]), .B(n10531), .Z(n10530) );
  IV U12465 ( .A(n10528), .Z(n10531) );
  XOR U12466 ( .A(n10532), .B(n10533), .Z(n10528) );
  ANDN U12467 ( .B(n10534), .A(n10535), .Z(n10532) );
  XNOR U12468 ( .A(b[2163]), .B(n10533), .Z(n10534) );
  XNOR U12469 ( .A(b[2163]), .B(n10535), .Z(c[2163]) );
  XNOR U12470 ( .A(a[2163]), .B(n10536), .Z(n10535) );
  IV U12471 ( .A(n10533), .Z(n10536) );
  XOR U12472 ( .A(n10537), .B(n10538), .Z(n10533) );
  ANDN U12473 ( .B(n10539), .A(n10540), .Z(n10537) );
  XNOR U12474 ( .A(b[2162]), .B(n10538), .Z(n10539) );
  XNOR U12475 ( .A(b[2162]), .B(n10540), .Z(c[2162]) );
  XNOR U12476 ( .A(a[2162]), .B(n10541), .Z(n10540) );
  IV U12477 ( .A(n10538), .Z(n10541) );
  XOR U12478 ( .A(n10542), .B(n10543), .Z(n10538) );
  ANDN U12479 ( .B(n10544), .A(n10545), .Z(n10542) );
  XNOR U12480 ( .A(b[2161]), .B(n10543), .Z(n10544) );
  XNOR U12481 ( .A(b[2161]), .B(n10545), .Z(c[2161]) );
  XNOR U12482 ( .A(a[2161]), .B(n10546), .Z(n10545) );
  IV U12483 ( .A(n10543), .Z(n10546) );
  XOR U12484 ( .A(n10547), .B(n10548), .Z(n10543) );
  ANDN U12485 ( .B(n10549), .A(n10550), .Z(n10547) );
  XNOR U12486 ( .A(b[2160]), .B(n10548), .Z(n10549) );
  XNOR U12487 ( .A(b[2160]), .B(n10550), .Z(c[2160]) );
  XNOR U12488 ( .A(a[2160]), .B(n10551), .Z(n10550) );
  IV U12489 ( .A(n10548), .Z(n10551) );
  XOR U12490 ( .A(n10552), .B(n10553), .Z(n10548) );
  ANDN U12491 ( .B(n10554), .A(n10555), .Z(n10552) );
  XNOR U12492 ( .A(b[2159]), .B(n10553), .Z(n10554) );
  XNOR U12493 ( .A(b[215]), .B(n10556), .Z(c[215]) );
  XNOR U12494 ( .A(b[2159]), .B(n10555), .Z(c[2159]) );
  XNOR U12495 ( .A(a[2159]), .B(n10557), .Z(n10555) );
  IV U12496 ( .A(n10553), .Z(n10557) );
  XOR U12497 ( .A(n10558), .B(n10559), .Z(n10553) );
  ANDN U12498 ( .B(n10560), .A(n10561), .Z(n10558) );
  XNOR U12499 ( .A(b[2158]), .B(n10559), .Z(n10560) );
  XNOR U12500 ( .A(b[2158]), .B(n10561), .Z(c[2158]) );
  XNOR U12501 ( .A(a[2158]), .B(n10562), .Z(n10561) );
  IV U12502 ( .A(n10559), .Z(n10562) );
  XOR U12503 ( .A(n10563), .B(n10564), .Z(n10559) );
  ANDN U12504 ( .B(n10565), .A(n10566), .Z(n10563) );
  XNOR U12505 ( .A(b[2157]), .B(n10564), .Z(n10565) );
  XNOR U12506 ( .A(b[2157]), .B(n10566), .Z(c[2157]) );
  XNOR U12507 ( .A(a[2157]), .B(n10567), .Z(n10566) );
  IV U12508 ( .A(n10564), .Z(n10567) );
  XOR U12509 ( .A(n10568), .B(n10569), .Z(n10564) );
  ANDN U12510 ( .B(n10570), .A(n10571), .Z(n10568) );
  XNOR U12511 ( .A(b[2156]), .B(n10569), .Z(n10570) );
  XNOR U12512 ( .A(b[2156]), .B(n10571), .Z(c[2156]) );
  XNOR U12513 ( .A(a[2156]), .B(n10572), .Z(n10571) );
  IV U12514 ( .A(n10569), .Z(n10572) );
  XOR U12515 ( .A(n10573), .B(n10574), .Z(n10569) );
  ANDN U12516 ( .B(n10575), .A(n10576), .Z(n10573) );
  XNOR U12517 ( .A(b[2155]), .B(n10574), .Z(n10575) );
  XNOR U12518 ( .A(b[2155]), .B(n10576), .Z(c[2155]) );
  XNOR U12519 ( .A(a[2155]), .B(n10577), .Z(n10576) );
  IV U12520 ( .A(n10574), .Z(n10577) );
  XOR U12521 ( .A(n10578), .B(n10579), .Z(n10574) );
  ANDN U12522 ( .B(n10580), .A(n10581), .Z(n10578) );
  XNOR U12523 ( .A(b[2154]), .B(n10579), .Z(n10580) );
  XNOR U12524 ( .A(b[2154]), .B(n10581), .Z(c[2154]) );
  XNOR U12525 ( .A(a[2154]), .B(n10582), .Z(n10581) );
  IV U12526 ( .A(n10579), .Z(n10582) );
  XOR U12527 ( .A(n10583), .B(n10584), .Z(n10579) );
  ANDN U12528 ( .B(n10585), .A(n10586), .Z(n10583) );
  XNOR U12529 ( .A(b[2153]), .B(n10584), .Z(n10585) );
  XNOR U12530 ( .A(b[2153]), .B(n10586), .Z(c[2153]) );
  XNOR U12531 ( .A(a[2153]), .B(n10587), .Z(n10586) );
  IV U12532 ( .A(n10584), .Z(n10587) );
  XOR U12533 ( .A(n10588), .B(n10589), .Z(n10584) );
  ANDN U12534 ( .B(n10590), .A(n10591), .Z(n10588) );
  XNOR U12535 ( .A(b[2152]), .B(n10589), .Z(n10590) );
  XNOR U12536 ( .A(b[2152]), .B(n10591), .Z(c[2152]) );
  XNOR U12537 ( .A(a[2152]), .B(n10592), .Z(n10591) );
  IV U12538 ( .A(n10589), .Z(n10592) );
  XOR U12539 ( .A(n10593), .B(n10594), .Z(n10589) );
  ANDN U12540 ( .B(n10595), .A(n10596), .Z(n10593) );
  XNOR U12541 ( .A(b[2151]), .B(n10594), .Z(n10595) );
  XNOR U12542 ( .A(b[2151]), .B(n10596), .Z(c[2151]) );
  XNOR U12543 ( .A(a[2151]), .B(n10597), .Z(n10596) );
  IV U12544 ( .A(n10594), .Z(n10597) );
  XOR U12545 ( .A(n10598), .B(n10599), .Z(n10594) );
  ANDN U12546 ( .B(n10600), .A(n10601), .Z(n10598) );
  XNOR U12547 ( .A(b[2150]), .B(n10599), .Z(n10600) );
  XNOR U12548 ( .A(b[2150]), .B(n10601), .Z(c[2150]) );
  XNOR U12549 ( .A(a[2150]), .B(n10602), .Z(n10601) );
  IV U12550 ( .A(n10599), .Z(n10602) );
  XOR U12551 ( .A(n10603), .B(n10604), .Z(n10599) );
  ANDN U12552 ( .B(n10605), .A(n10606), .Z(n10603) );
  XNOR U12553 ( .A(b[2149]), .B(n10604), .Z(n10605) );
  XNOR U12554 ( .A(b[214]), .B(n10607), .Z(c[214]) );
  XNOR U12555 ( .A(b[2149]), .B(n10606), .Z(c[2149]) );
  XNOR U12556 ( .A(a[2149]), .B(n10608), .Z(n10606) );
  IV U12557 ( .A(n10604), .Z(n10608) );
  XOR U12558 ( .A(n10609), .B(n10610), .Z(n10604) );
  ANDN U12559 ( .B(n10611), .A(n10612), .Z(n10609) );
  XNOR U12560 ( .A(b[2148]), .B(n10610), .Z(n10611) );
  XNOR U12561 ( .A(b[2148]), .B(n10612), .Z(c[2148]) );
  XNOR U12562 ( .A(a[2148]), .B(n10613), .Z(n10612) );
  IV U12563 ( .A(n10610), .Z(n10613) );
  XOR U12564 ( .A(n10614), .B(n10615), .Z(n10610) );
  ANDN U12565 ( .B(n10616), .A(n10617), .Z(n10614) );
  XNOR U12566 ( .A(b[2147]), .B(n10615), .Z(n10616) );
  XNOR U12567 ( .A(b[2147]), .B(n10617), .Z(c[2147]) );
  XNOR U12568 ( .A(a[2147]), .B(n10618), .Z(n10617) );
  IV U12569 ( .A(n10615), .Z(n10618) );
  XOR U12570 ( .A(n10619), .B(n10620), .Z(n10615) );
  ANDN U12571 ( .B(n10621), .A(n10622), .Z(n10619) );
  XNOR U12572 ( .A(b[2146]), .B(n10620), .Z(n10621) );
  XNOR U12573 ( .A(b[2146]), .B(n10622), .Z(c[2146]) );
  XNOR U12574 ( .A(a[2146]), .B(n10623), .Z(n10622) );
  IV U12575 ( .A(n10620), .Z(n10623) );
  XOR U12576 ( .A(n10624), .B(n10625), .Z(n10620) );
  ANDN U12577 ( .B(n10626), .A(n10627), .Z(n10624) );
  XNOR U12578 ( .A(b[2145]), .B(n10625), .Z(n10626) );
  XNOR U12579 ( .A(b[2145]), .B(n10627), .Z(c[2145]) );
  XNOR U12580 ( .A(a[2145]), .B(n10628), .Z(n10627) );
  IV U12581 ( .A(n10625), .Z(n10628) );
  XOR U12582 ( .A(n10629), .B(n10630), .Z(n10625) );
  ANDN U12583 ( .B(n10631), .A(n10632), .Z(n10629) );
  XNOR U12584 ( .A(b[2144]), .B(n10630), .Z(n10631) );
  XNOR U12585 ( .A(b[2144]), .B(n10632), .Z(c[2144]) );
  XNOR U12586 ( .A(a[2144]), .B(n10633), .Z(n10632) );
  IV U12587 ( .A(n10630), .Z(n10633) );
  XOR U12588 ( .A(n10634), .B(n10635), .Z(n10630) );
  ANDN U12589 ( .B(n10636), .A(n10637), .Z(n10634) );
  XNOR U12590 ( .A(b[2143]), .B(n10635), .Z(n10636) );
  XNOR U12591 ( .A(b[2143]), .B(n10637), .Z(c[2143]) );
  XNOR U12592 ( .A(a[2143]), .B(n10638), .Z(n10637) );
  IV U12593 ( .A(n10635), .Z(n10638) );
  XOR U12594 ( .A(n10639), .B(n10640), .Z(n10635) );
  ANDN U12595 ( .B(n10641), .A(n10642), .Z(n10639) );
  XNOR U12596 ( .A(b[2142]), .B(n10640), .Z(n10641) );
  XNOR U12597 ( .A(b[2142]), .B(n10642), .Z(c[2142]) );
  XNOR U12598 ( .A(a[2142]), .B(n10643), .Z(n10642) );
  IV U12599 ( .A(n10640), .Z(n10643) );
  XOR U12600 ( .A(n10644), .B(n10645), .Z(n10640) );
  ANDN U12601 ( .B(n10646), .A(n10647), .Z(n10644) );
  XNOR U12602 ( .A(b[2141]), .B(n10645), .Z(n10646) );
  XNOR U12603 ( .A(b[2141]), .B(n10647), .Z(c[2141]) );
  XNOR U12604 ( .A(a[2141]), .B(n10648), .Z(n10647) );
  IV U12605 ( .A(n10645), .Z(n10648) );
  XOR U12606 ( .A(n10649), .B(n10650), .Z(n10645) );
  ANDN U12607 ( .B(n10651), .A(n10652), .Z(n10649) );
  XNOR U12608 ( .A(b[2140]), .B(n10650), .Z(n10651) );
  XNOR U12609 ( .A(b[2140]), .B(n10652), .Z(c[2140]) );
  XNOR U12610 ( .A(a[2140]), .B(n10653), .Z(n10652) );
  IV U12611 ( .A(n10650), .Z(n10653) );
  XOR U12612 ( .A(n10654), .B(n10655), .Z(n10650) );
  ANDN U12613 ( .B(n10656), .A(n10657), .Z(n10654) );
  XNOR U12614 ( .A(b[2139]), .B(n10655), .Z(n10656) );
  XNOR U12615 ( .A(b[213]), .B(n10658), .Z(c[213]) );
  XNOR U12616 ( .A(b[2139]), .B(n10657), .Z(c[2139]) );
  XNOR U12617 ( .A(a[2139]), .B(n10659), .Z(n10657) );
  IV U12618 ( .A(n10655), .Z(n10659) );
  XOR U12619 ( .A(n10660), .B(n10661), .Z(n10655) );
  ANDN U12620 ( .B(n10662), .A(n10663), .Z(n10660) );
  XNOR U12621 ( .A(b[2138]), .B(n10661), .Z(n10662) );
  XNOR U12622 ( .A(b[2138]), .B(n10663), .Z(c[2138]) );
  XNOR U12623 ( .A(a[2138]), .B(n10664), .Z(n10663) );
  IV U12624 ( .A(n10661), .Z(n10664) );
  XOR U12625 ( .A(n10665), .B(n10666), .Z(n10661) );
  ANDN U12626 ( .B(n10667), .A(n10668), .Z(n10665) );
  XNOR U12627 ( .A(b[2137]), .B(n10666), .Z(n10667) );
  XNOR U12628 ( .A(b[2137]), .B(n10668), .Z(c[2137]) );
  XNOR U12629 ( .A(a[2137]), .B(n10669), .Z(n10668) );
  IV U12630 ( .A(n10666), .Z(n10669) );
  XOR U12631 ( .A(n10670), .B(n10671), .Z(n10666) );
  ANDN U12632 ( .B(n10672), .A(n10673), .Z(n10670) );
  XNOR U12633 ( .A(b[2136]), .B(n10671), .Z(n10672) );
  XNOR U12634 ( .A(b[2136]), .B(n10673), .Z(c[2136]) );
  XNOR U12635 ( .A(a[2136]), .B(n10674), .Z(n10673) );
  IV U12636 ( .A(n10671), .Z(n10674) );
  XOR U12637 ( .A(n10675), .B(n10676), .Z(n10671) );
  ANDN U12638 ( .B(n10677), .A(n10678), .Z(n10675) );
  XNOR U12639 ( .A(b[2135]), .B(n10676), .Z(n10677) );
  XNOR U12640 ( .A(b[2135]), .B(n10678), .Z(c[2135]) );
  XNOR U12641 ( .A(a[2135]), .B(n10679), .Z(n10678) );
  IV U12642 ( .A(n10676), .Z(n10679) );
  XOR U12643 ( .A(n10680), .B(n10681), .Z(n10676) );
  ANDN U12644 ( .B(n10682), .A(n10683), .Z(n10680) );
  XNOR U12645 ( .A(b[2134]), .B(n10681), .Z(n10682) );
  XNOR U12646 ( .A(b[2134]), .B(n10683), .Z(c[2134]) );
  XNOR U12647 ( .A(a[2134]), .B(n10684), .Z(n10683) );
  IV U12648 ( .A(n10681), .Z(n10684) );
  XOR U12649 ( .A(n10685), .B(n10686), .Z(n10681) );
  ANDN U12650 ( .B(n10687), .A(n10688), .Z(n10685) );
  XNOR U12651 ( .A(b[2133]), .B(n10686), .Z(n10687) );
  XNOR U12652 ( .A(b[2133]), .B(n10688), .Z(c[2133]) );
  XNOR U12653 ( .A(a[2133]), .B(n10689), .Z(n10688) );
  IV U12654 ( .A(n10686), .Z(n10689) );
  XOR U12655 ( .A(n10690), .B(n10691), .Z(n10686) );
  ANDN U12656 ( .B(n10692), .A(n10693), .Z(n10690) );
  XNOR U12657 ( .A(b[2132]), .B(n10691), .Z(n10692) );
  XNOR U12658 ( .A(b[2132]), .B(n10693), .Z(c[2132]) );
  XNOR U12659 ( .A(a[2132]), .B(n10694), .Z(n10693) );
  IV U12660 ( .A(n10691), .Z(n10694) );
  XOR U12661 ( .A(n10695), .B(n10696), .Z(n10691) );
  ANDN U12662 ( .B(n10697), .A(n10698), .Z(n10695) );
  XNOR U12663 ( .A(b[2131]), .B(n10696), .Z(n10697) );
  XNOR U12664 ( .A(b[2131]), .B(n10698), .Z(c[2131]) );
  XNOR U12665 ( .A(a[2131]), .B(n10699), .Z(n10698) );
  IV U12666 ( .A(n10696), .Z(n10699) );
  XOR U12667 ( .A(n10700), .B(n10701), .Z(n10696) );
  ANDN U12668 ( .B(n10702), .A(n10703), .Z(n10700) );
  XNOR U12669 ( .A(b[2130]), .B(n10701), .Z(n10702) );
  XNOR U12670 ( .A(b[2130]), .B(n10703), .Z(c[2130]) );
  XNOR U12671 ( .A(a[2130]), .B(n10704), .Z(n10703) );
  IV U12672 ( .A(n10701), .Z(n10704) );
  XOR U12673 ( .A(n10705), .B(n10706), .Z(n10701) );
  ANDN U12674 ( .B(n10707), .A(n10708), .Z(n10705) );
  XNOR U12675 ( .A(b[2129]), .B(n10706), .Z(n10707) );
  XNOR U12676 ( .A(b[212]), .B(n10709), .Z(c[212]) );
  XNOR U12677 ( .A(b[2129]), .B(n10708), .Z(c[2129]) );
  XNOR U12678 ( .A(a[2129]), .B(n10710), .Z(n10708) );
  IV U12679 ( .A(n10706), .Z(n10710) );
  XOR U12680 ( .A(n10711), .B(n10712), .Z(n10706) );
  ANDN U12681 ( .B(n10713), .A(n10714), .Z(n10711) );
  XNOR U12682 ( .A(b[2128]), .B(n10712), .Z(n10713) );
  XNOR U12683 ( .A(b[2128]), .B(n10714), .Z(c[2128]) );
  XNOR U12684 ( .A(a[2128]), .B(n10715), .Z(n10714) );
  IV U12685 ( .A(n10712), .Z(n10715) );
  XOR U12686 ( .A(n10716), .B(n10717), .Z(n10712) );
  ANDN U12687 ( .B(n10718), .A(n10719), .Z(n10716) );
  XNOR U12688 ( .A(b[2127]), .B(n10717), .Z(n10718) );
  XNOR U12689 ( .A(b[2127]), .B(n10719), .Z(c[2127]) );
  XNOR U12690 ( .A(a[2127]), .B(n10720), .Z(n10719) );
  IV U12691 ( .A(n10717), .Z(n10720) );
  XOR U12692 ( .A(n10721), .B(n10722), .Z(n10717) );
  ANDN U12693 ( .B(n10723), .A(n10724), .Z(n10721) );
  XNOR U12694 ( .A(b[2126]), .B(n10722), .Z(n10723) );
  XNOR U12695 ( .A(b[2126]), .B(n10724), .Z(c[2126]) );
  XNOR U12696 ( .A(a[2126]), .B(n10725), .Z(n10724) );
  IV U12697 ( .A(n10722), .Z(n10725) );
  XOR U12698 ( .A(n10726), .B(n10727), .Z(n10722) );
  ANDN U12699 ( .B(n10728), .A(n10729), .Z(n10726) );
  XNOR U12700 ( .A(b[2125]), .B(n10727), .Z(n10728) );
  XNOR U12701 ( .A(b[2125]), .B(n10729), .Z(c[2125]) );
  XNOR U12702 ( .A(a[2125]), .B(n10730), .Z(n10729) );
  IV U12703 ( .A(n10727), .Z(n10730) );
  XOR U12704 ( .A(n10731), .B(n10732), .Z(n10727) );
  ANDN U12705 ( .B(n10733), .A(n10734), .Z(n10731) );
  XNOR U12706 ( .A(b[2124]), .B(n10732), .Z(n10733) );
  XNOR U12707 ( .A(b[2124]), .B(n10734), .Z(c[2124]) );
  XNOR U12708 ( .A(a[2124]), .B(n10735), .Z(n10734) );
  IV U12709 ( .A(n10732), .Z(n10735) );
  XOR U12710 ( .A(n10736), .B(n10737), .Z(n10732) );
  ANDN U12711 ( .B(n10738), .A(n10739), .Z(n10736) );
  XNOR U12712 ( .A(b[2123]), .B(n10737), .Z(n10738) );
  XNOR U12713 ( .A(b[2123]), .B(n10739), .Z(c[2123]) );
  XNOR U12714 ( .A(a[2123]), .B(n10740), .Z(n10739) );
  IV U12715 ( .A(n10737), .Z(n10740) );
  XOR U12716 ( .A(n10741), .B(n10742), .Z(n10737) );
  ANDN U12717 ( .B(n10743), .A(n10744), .Z(n10741) );
  XNOR U12718 ( .A(b[2122]), .B(n10742), .Z(n10743) );
  XNOR U12719 ( .A(b[2122]), .B(n10744), .Z(c[2122]) );
  XNOR U12720 ( .A(a[2122]), .B(n10745), .Z(n10744) );
  IV U12721 ( .A(n10742), .Z(n10745) );
  XOR U12722 ( .A(n10746), .B(n10747), .Z(n10742) );
  ANDN U12723 ( .B(n10748), .A(n10749), .Z(n10746) );
  XNOR U12724 ( .A(b[2121]), .B(n10747), .Z(n10748) );
  XNOR U12725 ( .A(b[2121]), .B(n10749), .Z(c[2121]) );
  XNOR U12726 ( .A(a[2121]), .B(n10750), .Z(n10749) );
  IV U12727 ( .A(n10747), .Z(n10750) );
  XOR U12728 ( .A(n10751), .B(n10752), .Z(n10747) );
  ANDN U12729 ( .B(n10753), .A(n10754), .Z(n10751) );
  XNOR U12730 ( .A(b[2120]), .B(n10752), .Z(n10753) );
  XNOR U12731 ( .A(b[2120]), .B(n10754), .Z(c[2120]) );
  XNOR U12732 ( .A(a[2120]), .B(n10755), .Z(n10754) );
  IV U12733 ( .A(n10752), .Z(n10755) );
  XOR U12734 ( .A(n10756), .B(n10757), .Z(n10752) );
  ANDN U12735 ( .B(n10758), .A(n10759), .Z(n10756) );
  XNOR U12736 ( .A(b[2119]), .B(n10757), .Z(n10758) );
  XNOR U12737 ( .A(b[211]), .B(n10760), .Z(c[211]) );
  XNOR U12738 ( .A(b[2119]), .B(n10759), .Z(c[2119]) );
  XNOR U12739 ( .A(a[2119]), .B(n10761), .Z(n10759) );
  IV U12740 ( .A(n10757), .Z(n10761) );
  XOR U12741 ( .A(n10762), .B(n10763), .Z(n10757) );
  ANDN U12742 ( .B(n10764), .A(n10765), .Z(n10762) );
  XNOR U12743 ( .A(b[2118]), .B(n10763), .Z(n10764) );
  XNOR U12744 ( .A(b[2118]), .B(n10765), .Z(c[2118]) );
  XNOR U12745 ( .A(a[2118]), .B(n10766), .Z(n10765) );
  IV U12746 ( .A(n10763), .Z(n10766) );
  XOR U12747 ( .A(n10767), .B(n10768), .Z(n10763) );
  ANDN U12748 ( .B(n10769), .A(n10770), .Z(n10767) );
  XNOR U12749 ( .A(b[2117]), .B(n10768), .Z(n10769) );
  XNOR U12750 ( .A(b[2117]), .B(n10770), .Z(c[2117]) );
  XNOR U12751 ( .A(a[2117]), .B(n10771), .Z(n10770) );
  IV U12752 ( .A(n10768), .Z(n10771) );
  XOR U12753 ( .A(n10772), .B(n10773), .Z(n10768) );
  ANDN U12754 ( .B(n10774), .A(n10775), .Z(n10772) );
  XNOR U12755 ( .A(b[2116]), .B(n10773), .Z(n10774) );
  XNOR U12756 ( .A(b[2116]), .B(n10775), .Z(c[2116]) );
  XNOR U12757 ( .A(a[2116]), .B(n10776), .Z(n10775) );
  IV U12758 ( .A(n10773), .Z(n10776) );
  XOR U12759 ( .A(n10777), .B(n10778), .Z(n10773) );
  ANDN U12760 ( .B(n10779), .A(n10780), .Z(n10777) );
  XNOR U12761 ( .A(b[2115]), .B(n10778), .Z(n10779) );
  XNOR U12762 ( .A(b[2115]), .B(n10780), .Z(c[2115]) );
  XNOR U12763 ( .A(a[2115]), .B(n10781), .Z(n10780) );
  IV U12764 ( .A(n10778), .Z(n10781) );
  XOR U12765 ( .A(n10782), .B(n10783), .Z(n10778) );
  ANDN U12766 ( .B(n10784), .A(n10785), .Z(n10782) );
  XNOR U12767 ( .A(b[2114]), .B(n10783), .Z(n10784) );
  XNOR U12768 ( .A(b[2114]), .B(n10785), .Z(c[2114]) );
  XNOR U12769 ( .A(a[2114]), .B(n10786), .Z(n10785) );
  IV U12770 ( .A(n10783), .Z(n10786) );
  XOR U12771 ( .A(n10787), .B(n10788), .Z(n10783) );
  ANDN U12772 ( .B(n10789), .A(n10790), .Z(n10787) );
  XNOR U12773 ( .A(b[2113]), .B(n10788), .Z(n10789) );
  XNOR U12774 ( .A(b[2113]), .B(n10790), .Z(c[2113]) );
  XNOR U12775 ( .A(a[2113]), .B(n10791), .Z(n10790) );
  IV U12776 ( .A(n10788), .Z(n10791) );
  XOR U12777 ( .A(n10792), .B(n10793), .Z(n10788) );
  ANDN U12778 ( .B(n10794), .A(n10795), .Z(n10792) );
  XNOR U12779 ( .A(b[2112]), .B(n10793), .Z(n10794) );
  XNOR U12780 ( .A(b[2112]), .B(n10795), .Z(c[2112]) );
  XNOR U12781 ( .A(a[2112]), .B(n10796), .Z(n10795) );
  IV U12782 ( .A(n10793), .Z(n10796) );
  XOR U12783 ( .A(n10797), .B(n10798), .Z(n10793) );
  ANDN U12784 ( .B(n10799), .A(n10800), .Z(n10797) );
  XNOR U12785 ( .A(b[2111]), .B(n10798), .Z(n10799) );
  XNOR U12786 ( .A(b[2111]), .B(n10800), .Z(c[2111]) );
  XNOR U12787 ( .A(a[2111]), .B(n10801), .Z(n10800) );
  IV U12788 ( .A(n10798), .Z(n10801) );
  XOR U12789 ( .A(n10802), .B(n10803), .Z(n10798) );
  ANDN U12790 ( .B(n10804), .A(n10805), .Z(n10802) );
  XNOR U12791 ( .A(b[2110]), .B(n10803), .Z(n10804) );
  XNOR U12792 ( .A(b[2110]), .B(n10805), .Z(c[2110]) );
  XNOR U12793 ( .A(a[2110]), .B(n10806), .Z(n10805) );
  IV U12794 ( .A(n10803), .Z(n10806) );
  XOR U12795 ( .A(n10807), .B(n10808), .Z(n10803) );
  ANDN U12796 ( .B(n10809), .A(n10810), .Z(n10807) );
  XNOR U12797 ( .A(b[2109]), .B(n10808), .Z(n10809) );
  XNOR U12798 ( .A(b[210]), .B(n10811), .Z(c[210]) );
  XNOR U12799 ( .A(b[2109]), .B(n10810), .Z(c[2109]) );
  XNOR U12800 ( .A(a[2109]), .B(n10812), .Z(n10810) );
  IV U12801 ( .A(n10808), .Z(n10812) );
  XOR U12802 ( .A(n10813), .B(n10814), .Z(n10808) );
  ANDN U12803 ( .B(n10815), .A(n10816), .Z(n10813) );
  XNOR U12804 ( .A(b[2108]), .B(n10814), .Z(n10815) );
  XNOR U12805 ( .A(b[2108]), .B(n10816), .Z(c[2108]) );
  XNOR U12806 ( .A(a[2108]), .B(n10817), .Z(n10816) );
  IV U12807 ( .A(n10814), .Z(n10817) );
  XOR U12808 ( .A(n10818), .B(n10819), .Z(n10814) );
  ANDN U12809 ( .B(n10820), .A(n10821), .Z(n10818) );
  XNOR U12810 ( .A(b[2107]), .B(n10819), .Z(n10820) );
  XNOR U12811 ( .A(b[2107]), .B(n10821), .Z(c[2107]) );
  XNOR U12812 ( .A(a[2107]), .B(n10822), .Z(n10821) );
  IV U12813 ( .A(n10819), .Z(n10822) );
  XOR U12814 ( .A(n10823), .B(n10824), .Z(n10819) );
  ANDN U12815 ( .B(n10825), .A(n10826), .Z(n10823) );
  XNOR U12816 ( .A(b[2106]), .B(n10824), .Z(n10825) );
  XNOR U12817 ( .A(b[2106]), .B(n10826), .Z(c[2106]) );
  XNOR U12818 ( .A(a[2106]), .B(n10827), .Z(n10826) );
  IV U12819 ( .A(n10824), .Z(n10827) );
  XOR U12820 ( .A(n10828), .B(n10829), .Z(n10824) );
  ANDN U12821 ( .B(n10830), .A(n10831), .Z(n10828) );
  XNOR U12822 ( .A(b[2105]), .B(n10829), .Z(n10830) );
  XNOR U12823 ( .A(b[2105]), .B(n10831), .Z(c[2105]) );
  XNOR U12824 ( .A(a[2105]), .B(n10832), .Z(n10831) );
  IV U12825 ( .A(n10829), .Z(n10832) );
  XOR U12826 ( .A(n10833), .B(n10834), .Z(n10829) );
  ANDN U12827 ( .B(n10835), .A(n10836), .Z(n10833) );
  XNOR U12828 ( .A(b[2104]), .B(n10834), .Z(n10835) );
  XNOR U12829 ( .A(b[2104]), .B(n10836), .Z(c[2104]) );
  XNOR U12830 ( .A(a[2104]), .B(n10837), .Z(n10836) );
  IV U12831 ( .A(n10834), .Z(n10837) );
  XOR U12832 ( .A(n10838), .B(n10839), .Z(n10834) );
  ANDN U12833 ( .B(n10840), .A(n10841), .Z(n10838) );
  XNOR U12834 ( .A(b[2103]), .B(n10839), .Z(n10840) );
  XNOR U12835 ( .A(b[2103]), .B(n10841), .Z(c[2103]) );
  XNOR U12836 ( .A(a[2103]), .B(n10842), .Z(n10841) );
  IV U12837 ( .A(n10839), .Z(n10842) );
  XOR U12838 ( .A(n10843), .B(n10844), .Z(n10839) );
  ANDN U12839 ( .B(n10845), .A(n10846), .Z(n10843) );
  XNOR U12840 ( .A(b[2102]), .B(n10844), .Z(n10845) );
  XNOR U12841 ( .A(b[2102]), .B(n10846), .Z(c[2102]) );
  XNOR U12842 ( .A(a[2102]), .B(n10847), .Z(n10846) );
  IV U12843 ( .A(n10844), .Z(n10847) );
  XOR U12844 ( .A(n10848), .B(n10849), .Z(n10844) );
  ANDN U12845 ( .B(n10850), .A(n10851), .Z(n10848) );
  XNOR U12846 ( .A(b[2101]), .B(n10849), .Z(n10850) );
  XNOR U12847 ( .A(b[2101]), .B(n10851), .Z(c[2101]) );
  XNOR U12848 ( .A(a[2101]), .B(n10852), .Z(n10851) );
  IV U12849 ( .A(n10849), .Z(n10852) );
  XOR U12850 ( .A(n10853), .B(n10854), .Z(n10849) );
  ANDN U12851 ( .B(n10855), .A(n10856), .Z(n10853) );
  XNOR U12852 ( .A(b[2100]), .B(n10854), .Z(n10855) );
  XNOR U12853 ( .A(b[2100]), .B(n10856), .Z(c[2100]) );
  XNOR U12854 ( .A(a[2100]), .B(n10857), .Z(n10856) );
  IV U12855 ( .A(n10854), .Z(n10857) );
  XOR U12856 ( .A(n10858), .B(n10859), .Z(n10854) );
  ANDN U12857 ( .B(n10860), .A(n10861), .Z(n10858) );
  XNOR U12858 ( .A(b[2099]), .B(n10859), .Z(n10860) );
  XNOR U12859 ( .A(b[20]), .B(n10862), .Z(c[20]) );
  XNOR U12860 ( .A(b[209]), .B(n10863), .Z(c[209]) );
  XNOR U12861 ( .A(b[2099]), .B(n10861), .Z(c[2099]) );
  XNOR U12862 ( .A(a[2099]), .B(n10864), .Z(n10861) );
  IV U12863 ( .A(n10859), .Z(n10864) );
  XOR U12864 ( .A(n10865), .B(n10866), .Z(n10859) );
  ANDN U12865 ( .B(n10867), .A(n10868), .Z(n10865) );
  XNOR U12866 ( .A(b[2098]), .B(n10866), .Z(n10867) );
  XNOR U12867 ( .A(b[2098]), .B(n10868), .Z(c[2098]) );
  XNOR U12868 ( .A(a[2098]), .B(n10869), .Z(n10868) );
  IV U12869 ( .A(n10866), .Z(n10869) );
  XOR U12870 ( .A(n10870), .B(n10871), .Z(n10866) );
  ANDN U12871 ( .B(n10872), .A(n10873), .Z(n10870) );
  XNOR U12872 ( .A(b[2097]), .B(n10871), .Z(n10872) );
  XNOR U12873 ( .A(b[2097]), .B(n10873), .Z(c[2097]) );
  XNOR U12874 ( .A(a[2097]), .B(n10874), .Z(n10873) );
  IV U12875 ( .A(n10871), .Z(n10874) );
  XOR U12876 ( .A(n10875), .B(n10876), .Z(n10871) );
  ANDN U12877 ( .B(n10877), .A(n10878), .Z(n10875) );
  XNOR U12878 ( .A(b[2096]), .B(n10876), .Z(n10877) );
  XNOR U12879 ( .A(b[2096]), .B(n10878), .Z(c[2096]) );
  XNOR U12880 ( .A(a[2096]), .B(n10879), .Z(n10878) );
  IV U12881 ( .A(n10876), .Z(n10879) );
  XOR U12882 ( .A(n10880), .B(n10881), .Z(n10876) );
  ANDN U12883 ( .B(n10882), .A(n10883), .Z(n10880) );
  XNOR U12884 ( .A(b[2095]), .B(n10881), .Z(n10882) );
  XNOR U12885 ( .A(b[2095]), .B(n10883), .Z(c[2095]) );
  XNOR U12886 ( .A(a[2095]), .B(n10884), .Z(n10883) );
  IV U12887 ( .A(n10881), .Z(n10884) );
  XOR U12888 ( .A(n10885), .B(n10886), .Z(n10881) );
  ANDN U12889 ( .B(n10887), .A(n10888), .Z(n10885) );
  XNOR U12890 ( .A(b[2094]), .B(n10886), .Z(n10887) );
  XNOR U12891 ( .A(b[2094]), .B(n10888), .Z(c[2094]) );
  XNOR U12892 ( .A(a[2094]), .B(n10889), .Z(n10888) );
  IV U12893 ( .A(n10886), .Z(n10889) );
  XOR U12894 ( .A(n10890), .B(n10891), .Z(n10886) );
  ANDN U12895 ( .B(n10892), .A(n10893), .Z(n10890) );
  XNOR U12896 ( .A(b[2093]), .B(n10891), .Z(n10892) );
  XNOR U12897 ( .A(b[2093]), .B(n10893), .Z(c[2093]) );
  XNOR U12898 ( .A(a[2093]), .B(n10894), .Z(n10893) );
  IV U12899 ( .A(n10891), .Z(n10894) );
  XOR U12900 ( .A(n10895), .B(n10896), .Z(n10891) );
  ANDN U12901 ( .B(n10897), .A(n10898), .Z(n10895) );
  XNOR U12902 ( .A(b[2092]), .B(n10896), .Z(n10897) );
  XNOR U12903 ( .A(b[2092]), .B(n10898), .Z(c[2092]) );
  XNOR U12904 ( .A(a[2092]), .B(n10899), .Z(n10898) );
  IV U12905 ( .A(n10896), .Z(n10899) );
  XOR U12906 ( .A(n10900), .B(n10901), .Z(n10896) );
  ANDN U12907 ( .B(n10902), .A(n10903), .Z(n10900) );
  XNOR U12908 ( .A(b[2091]), .B(n10901), .Z(n10902) );
  XNOR U12909 ( .A(b[2091]), .B(n10903), .Z(c[2091]) );
  XNOR U12910 ( .A(a[2091]), .B(n10904), .Z(n10903) );
  IV U12911 ( .A(n10901), .Z(n10904) );
  XOR U12912 ( .A(n10905), .B(n10906), .Z(n10901) );
  ANDN U12913 ( .B(n10907), .A(n10908), .Z(n10905) );
  XNOR U12914 ( .A(b[2090]), .B(n10906), .Z(n10907) );
  XNOR U12915 ( .A(b[2090]), .B(n10908), .Z(c[2090]) );
  XNOR U12916 ( .A(a[2090]), .B(n10909), .Z(n10908) );
  IV U12917 ( .A(n10906), .Z(n10909) );
  XOR U12918 ( .A(n10910), .B(n10911), .Z(n10906) );
  ANDN U12919 ( .B(n10912), .A(n10913), .Z(n10910) );
  XNOR U12920 ( .A(b[2089]), .B(n10911), .Z(n10912) );
  XNOR U12921 ( .A(b[208]), .B(n10914), .Z(c[208]) );
  XNOR U12922 ( .A(b[2089]), .B(n10913), .Z(c[2089]) );
  XNOR U12923 ( .A(a[2089]), .B(n10915), .Z(n10913) );
  IV U12924 ( .A(n10911), .Z(n10915) );
  XOR U12925 ( .A(n10916), .B(n10917), .Z(n10911) );
  ANDN U12926 ( .B(n10918), .A(n10919), .Z(n10916) );
  XNOR U12927 ( .A(b[2088]), .B(n10917), .Z(n10918) );
  XNOR U12928 ( .A(b[2088]), .B(n10919), .Z(c[2088]) );
  XNOR U12929 ( .A(a[2088]), .B(n10920), .Z(n10919) );
  IV U12930 ( .A(n10917), .Z(n10920) );
  XOR U12931 ( .A(n10921), .B(n10922), .Z(n10917) );
  ANDN U12932 ( .B(n10923), .A(n10924), .Z(n10921) );
  XNOR U12933 ( .A(b[2087]), .B(n10922), .Z(n10923) );
  XNOR U12934 ( .A(b[2087]), .B(n10924), .Z(c[2087]) );
  XNOR U12935 ( .A(a[2087]), .B(n10925), .Z(n10924) );
  IV U12936 ( .A(n10922), .Z(n10925) );
  XOR U12937 ( .A(n10926), .B(n10927), .Z(n10922) );
  ANDN U12938 ( .B(n10928), .A(n10929), .Z(n10926) );
  XNOR U12939 ( .A(b[2086]), .B(n10927), .Z(n10928) );
  XNOR U12940 ( .A(b[2086]), .B(n10929), .Z(c[2086]) );
  XNOR U12941 ( .A(a[2086]), .B(n10930), .Z(n10929) );
  IV U12942 ( .A(n10927), .Z(n10930) );
  XOR U12943 ( .A(n10931), .B(n10932), .Z(n10927) );
  ANDN U12944 ( .B(n10933), .A(n10934), .Z(n10931) );
  XNOR U12945 ( .A(b[2085]), .B(n10932), .Z(n10933) );
  XNOR U12946 ( .A(b[2085]), .B(n10934), .Z(c[2085]) );
  XNOR U12947 ( .A(a[2085]), .B(n10935), .Z(n10934) );
  IV U12948 ( .A(n10932), .Z(n10935) );
  XOR U12949 ( .A(n10936), .B(n10937), .Z(n10932) );
  ANDN U12950 ( .B(n10938), .A(n10939), .Z(n10936) );
  XNOR U12951 ( .A(b[2084]), .B(n10937), .Z(n10938) );
  XNOR U12952 ( .A(b[2084]), .B(n10939), .Z(c[2084]) );
  XNOR U12953 ( .A(a[2084]), .B(n10940), .Z(n10939) );
  IV U12954 ( .A(n10937), .Z(n10940) );
  XOR U12955 ( .A(n10941), .B(n10942), .Z(n10937) );
  ANDN U12956 ( .B(n10943), .A(n10944), .Z(n10941) );
  XNOR U12957 ( .A(b[2083]), .B(n10942), .Z(n10943) );
  XNOR U12958 ( .A(b[2083]), .B(n10944), .Z(c[2083]) );
  XNOR U12959 ( .A(a[2083]), .B(n10945), .Z(n10944) );
  IV U12960 ( .A(n10942), .Z(n10945) );
  XOR U12961 ( .A(n10946), .B(n10947), .Z(n10942) );
  ANDN U12962 ( .B(n10948), .A(n10949), .Z(n10946) );
  XNOR U12963 ( .A(b[2082]), .B(n10947), .Z(n10948) );
  XNOR U12964 ( .A(b[2082]), .B(n10949), .Z(c[2082]) );
  XNOR U12965 ( .A(a[2082]), .B(n10950), .Z(n10949) );
  IV U12966 ( .A(n10947), .Z(n10950) );
  XOR U12967 ( .A(n10951), .B(n10952), .Z(n10947) );
  ANDN U12968 ( .B(n10953), .A(n10954), .Z(n10951) );
  XNOR U12969 ( .A(b[2081]), .B(n10952), .Z(n10953) );
  XNOR U12970 ( .A(b[2081]), .B(n10954), .Z(c[2081]) );
  XNOR U12971 ( .A(a[2081]), .B(n10955), .Z(n10954) );
  IV U12972 ( .A(n10952), .Z(n10955) );
  XOR U12973 ( .A(n10956), .B(n10957), .Z(n10952) );
  ANDN U12974 ( .B(n10958), .A(n10959), .Z(n10956) );
  XNOR U12975 ( .A(b[2080]), .B(n10957), .Z(n10958) );
  XNOR U12976 ( .A(b[2080]), .B(n10959), .Z(c[2080]) );
  XNOR U12977 ( .A(a[2080]), .B(n10960), .Z(n10959) );
  IV U12978 ( .A(n10957), .Z(n10960) );
  XOR U12979 ( .A(n10961), .B(n10962), .Z(n10957) );
  ANDN U12980 ( .B(n10963), .A(n10964), .Z(n10961) );
  XNOR U12981 ( .A(b[2079]), .B(n10962), .Z(n10963) );
  XNOR U12982 ( .A(b[207]), .B(n10965), .Z(c[207]) );
  XNOR U12983 ( .A(b[2079]), .B(n10964), .Z(c[2079]) );
  XNOR U12984 ( .A(a[2079]), .B(n10966), .Z(n10964) );
  IV U12985 ( .A(n10962), .Z(n10966) );
  XOR U12986 ( .A(n10967), .B(n10968), .Z(n10962) );
  ANDN U12987 ( .B(n10969), .A(n10970), .Z(n10967) );
  XNOR U12988 ( .A(b[2078]), .B(n10968), .Z(n10969) );
  XNOR U12989 ( .A(b[2078]), .B(n10970), .Z(c[2078]) );
  XNOR U12990 ( .A(a[2078]), .B(n10971), .Z(n10970) );
  IV U12991 ( .A(n10968), .Z(n10971) );
  XOR U12992 ( .A(n10972), .B(n10973), .Z(n10968) );
  ANDN U12993 ( .B(n10974), .A(n10975), .Z(n10972) );
  XNOR U12994 ( .A(b[2077]), .B(n10973), .Z(n10974) );
  XNOR U12995 ( .A(b[2077]), .B(n10975), .Z(c[2077]) );
  XNOR U12996 ( .A(a[2077]), .B(n10976), .Z(n10975) );
  IV U12997 ( .A(n10973), .Z(n10976) );
  XOR U12998 ( .A(n10977), .B(n10978), .Z(n10973) );
  ANDN U12999 ( .B(n10979), .A(n10980), .Z(n10977) );
  XNOR U13000 ( .A(b[2076]), .B(n10978), .Z(n10979) );
  XNOR U13001 ( .A(b[2076]), .B(n10980), .Z(c[2076]) );
  XNOR U13002 ( .A(a[2076]), .B(n10981), .Z(n10980) );
  IV U13003 ( .A(n10978), .Z(n10981) );
  XOR U13004 ( .A(n10982), .B(n10983), .Z(n10978) );
  ANDN U13005 ( .B(n10984), .A(n10985), .Z(n10982) );
  XNOR U13006 ( .A(b[2075]), .B(n10983), .Z(n10984) );
  XNOR U13007 ( .A(b[2075]), .B(n10985), .Z(c[2075]) );
  XNOR U13008 ( .A(a[2075]), .B(n10986), .Z(n10985) );
  IV U13009 ( .A(n10983), .Z(n10986) );
  XOR U13010 ( .A(n10987), .B(n10988), .Z(n10983) );
  ANDN U13011 ( .B(n10989), .A(n10990), .Z(n10987) );
  XNOR U13012 ( .A(b[2074]), .B(n10988), .Z(n10989) );
  XNOR U13013 ( .A(b[2074]), .B(n10990), .Z(c[2074]) );
  XNOR U13014 ( .A(a[2074]), .B(n10991), .Z(n10990) );
  IV U13015 ( .A(n10988), .Z(n10991) );
  XOR U13016 ( .A(n10992), .B(n10993), .Z(n10988) );
  ANDN U13017 ( .B(n10994), .A(n10995), .Z(n10992) );
  XNOR U13018 ( .A(b[2073]), .B(n10993), .Z(n10994) );
  XNOR U13019 ( .A(b[2073]), .B(n10995), .Z(c[2073]) );
  XNOR U13020 ( .A(a[2073]), .B(n10996), .Z(n10995) );
  IV U13021 ( .A(n10993), .Z(n10996) );
  XOR U13022 ( .A(n10997), .B(n10998), .Z(n10993) );
  ANDN U13023 ( .B(n10999), .A(n11000), .Z(n10997) );
  XNOR U13024 ( .A(b[2072]), .B(n10998), .Z(n10999) );
  XNOR U13025 ( .A(b[2072]), .B(n11000), .Z(c[2072]) );
  XNOR U13026 ( .A(a[2072]), .B(n11001), .Z(n11000) );
  IV U13027 ( .A(n10998), .Z(n11001) );
  XOR U13028 ( .A(n11002), .B(n11003), .Z(n10998) );
  ANDN U13029 ( .B(n11004), .A(n11005), .Z(n11002) );
  XNOR U13030 ( .A(b[2071]), .B(n11003), .Z(n11004) );
  XNOR U13031 ( .A(b[2071]), .B(n11005), .Z(c[2071]) );
  XNOR U13032 ( .A(a[2071]), .B(n11006), .Z(n11005) );
  IV U13033 ( .A(n11003), .Z(n11006) );
  XOR U13034 ( .A(n11007), .B(n11008), .Z(n11003) );
  ANDN U13035 ( .B(n11009), .A(n11010), .Z(n11007) );
  XNOR U13036 ( .A(b[2070]), .B(n11008), .Z(n11009) );
  XNOR U13037 ( .A(b[2070]), .B(n11010), .Z(c[2070]) );
  XNOR U13038 ( .A(a[2070]), .B(n11011), .Z(n11010) );
  IV U13039 ( .A(n11008), .Z(n11011) );
  XOR U13040 ( .A(n11012), .B(n11013), .Z(n11008) );
  ANDN U13041 ( .B(n11014), .A(n11015), .Z(n11012) );
  XNOR U13042 ( .A(b[2069]), .B(n11013), .Z(n11014) );
  XNOR U13043 ( .A(b[206]), .B(n11016), .Z(c[206]) );
  XNOR U13044 ( .A(b[2069]), .B(n11015), .Z(c[2069]) );
  XNOR U13045 ( .A(a[2069]), .B(n11017), .Z(n11015) );
  IV U13046 ( .A(n11013), .Z(n11017) );
  XOR U13047 ( .A(n11018), .B(n11019), .Z(n11013) );
  ANDN U13048 ( .B(n11020), .A(n11021), .Z(n11018) );
  XNOR U13049 ( .A(b[2068]), .B(n11019), .Z(n11020) );
  XNOR U13050 ( .A(b[2068]), .B(n11021), .Z(c[2068]) );
  XNOR U13051 ( .A(a[2068]), .B(n11022), .Z(n11021) );
  IV U13052 ( .A(n11019), .Z(n11022) );
  XOR U13053 ( .A(n11023), .B(n11024), .Z(n11019) );
  ANDN U13054 ( .B(n11025), .A(n11026), .Z(n11023) );
  XNOR U13055 ( .A(b[2067]), .B(n11024), .Z(n11025) );
  XNOR U13056 ( .A(b[2067]), .B(n11026), .Z(c[2067]) );
  XNOR U13057 ( .A(a[2067]), .B(n11027), .Z(n11026) );
  IV U13058 ( .A(n11024), .Z(n11027) );
  XOR U13059 ( .A(n11028), .B(n11029), .Z(n11024) );
  ANDN U13060 ( .B(n11030), .A(n11031), .Z(n11028) );
  XNOR U13061 ( .A(b[2066]), .B(n11029), .Z(n11030) );
  XNOR U13062 ( .A(b[2066]), .B(n11031), .Z(c[2066]) );
  XNOR U13063 ( .A(a[2066]), .B(n11032), .Z(n11031) );
  IV U13064 ( .A(n11029), .Z(n11032) );
  XOR U13065 ( .A(n11033), .B(n11034), .Z(n11029) );
  ANDN U13066 ( .B(n11035), .A(n11036), .Z(n11033) );
  XNOR U13067 ( .A(b[2065]), .B(n11034), .Z(n11035) );
  XNOR U13068 ( .A(b[2065]), .B(n11036), .Z(c[2065]) );
  XNOR U13069 ( .A(a[2065]), .B(n11037), .Z(n11036) );
  IV U13070 ( .A(n11034), .Z(n11037) );
  XOR U13071 ( .A(n11038), .B(n11039), .Z(n11034) );
  ANDN U13072 ( .B(n11040), .A(n11041), .Z(n11038) );
  XNOR U13073 ( .A(b[2064]), .B(n11039), .Z(n11040) );
  XNOR U13074 ( .A(b[2064]), .B(n11041), .Z(c[2064]) );
  XNOR U13075 ( .A(a[2064]), .B(n11042), .Z(n11041) );
  IV U13076 ( .A(n11039), .Z(n11042) );
  XOR U13077 ( .A(n11043), .B(n11044), .Z(n11039) );
  ANDN U13078 ( .B(n11045), .A(n11046), .Z(n11043) );
  XNOR U13079 ( .A(b[2063]), .B(n11044), .Z(n11045) );
  XNOR U13080 ( .A(b[2063]), .B(n11046), .Z(c[2063]) );
  XNOR U13081 ( .A(a[2063]), .B(n11047), .Z(n11046) );
  IV U13082 ( .A(n11044), .Z(n11047) );
  XOR U13083 ( .A(n11048), .B(n11049), .Z(n11044) );
  ANDN U13084 ( .B(n11050), .A(n11051), .Z(n11048) );
  XNOR U13085 ( .A(b[2062]), .B(n11049), .Z(n11050) );
  XNOR U13086 ( .A(b[2062]), .B(n11051), .Z(c[2062]) );
  XNOR U13087 ( .A(a[2062]), .B(n11052), .Z(n11051) );
  IV U13088 ( .A(n11049), .Z(n11052) );
  XOR U13089 ( .A(n11053), .B(n11054), .Z(n11049) );
  ANDN U13090 ( .B(n11055), .A(n11056), .Z(n11053) );
  XNOR U13091 ( .A(b[2061]), .B(n11054), .Z(n11055) );
  XNOR U13092 ( .A(b[2061]), .B(n11056), .Z(c[2061]) );
  XNOR U13093 ( .A(a[2061]), .B(n11057), .Z(n11056) );
  IV U13094 ( .A(n11054), .Z(n11057) );
  XOR U13095 ( .A(n11058), .B(n11059), .Z(n11054) );
  ANDN U13096 ( .B(n11060), .A(n11061), .Z(n11058) );
  XNOR U13097 ( .A(b[2060]), .B(n11059), .Z(n11060) );
  XNOR U13098 ( .A(b[2060]), .B(n11061), .Z(c[2060]) );
  XNOR U13099 ( .A(a[2060]), .B(n11062), .Z(n11061) );
  IV U13100 ( .A(n11059), .Z(n11062) );
  XOR U13101 ( .A(n11063), .B(n11064), .Z(n11059) );
  ANDN U13102 ( .B(n11065), .A(n11066), .Z(n11063) );
  XNOR U13103 ( .A(b[2059]), .B(n11064), .Z(n11065) );
  XNOR U13104 ( .A(b[205]), .B(n11067), .Z(c[205]) );
  XNOR U13105 ( .A(b[2059]), .B(n11066), .Z(c[2059]) );
  XNOR U13106 ( .A(a[2059]), .B(n11068), .Z(n11066) );
  IV U13107 ( .A(n11064), .Z(n11068) );
  XOR U13108 ( .A(n11069), .B(n11070), .Z(n11064) );
  ANDN U13109 ( .B(n11071), .A(n11072), .Z(n11069) );
  XNOR U13110 ( .A(b[2058]), .B(n11070), .Z(n11071) );
  XNOR U13111 ( .A(b[2058]), .B(n11072), .Z(c[2058]) );
  XNOR U13112 ( .A(a[2058]), .B(n11073), .Z(n11072) );
  IV U13113 ( .A(n11070), .Z(n11073) );
  XOR U13114 ( .A(n11074), .B(n11075), .Z(n11070) );
  ANDN U13115 ( .B(n11076), .A(n11077), .Z(n11074) );
  XNOR U13116 ( .A(b[2057]), .B(n11075), .Z(n11076) );
  XNOR U13117 ( .A(b[2057]), .B(n11077), .Z(c[2057]) );
  XNOR U13118 ( .A(a[2057]), .B(n11078), .Z(n11077) );
  IV U13119 ( .A(n11075), .Z(n11078) );
  XOR U13120 ( .A(n11079), .B(n11080), .Z(n11075) );
  ANDN U13121 ( .B(n11081), .A(n11082), .Z(n11079) );
  XNOR U13122 ( .A(b[2056]), .B(n11080), .Z(n11081) );
  XNOR U13123 ( .A(b[2056]), .B(n11082), .Z(c[2056]) );
  XNOR U13124 ( .A(a[2056]), .B(n11083), .Z(n11082) );
  IV U13125 ( .A(n11080), .Z(n11083) );
  XOR U13126 ( .A(n11084), .B(n11085), .Z(n11080) );
  ANDN U13127 ( .B(n11086), .A(n11087), .Z(n11084) );
  XNOR U13128 ( .A(b[2055]), .B(n11085), .Z(n11086) );
  XNOR U13129 ( .A(b[2055]), .B(n11087), .Z(c[2055]) );
  XNOR U13130 ( .A(a[2055]), .B(n11088), .Z(n11087) );
  IV U13131 ( .A(n11085), .Z(n11088) );
  XOR U13132 ( .A(n11089), .B(n11090), .Z(n11085) );
  ANDN U13133 ( .B(n11091), .A(n11092), .Z(n11089) );
  XNOR U13134 ( .A(b[2054]), .B(n11090), .Z(n11091) );
  XNOR U13135 ( .A(b[2054]), .B(n11092), .Z(c[2054]) );
  XNOR U13136 ( .A(a[2054]), .B(n11093), .Z(n11092) );
  IV U13137 ( .A(n11090), .Z(n11093) );
  XOR U13138 ( .A(n11094), .B(n11095), .Z(n11090) );
  ANDN U13139 ( .B(n11096), .A(n11097), .Z(n11094) );
  XNOR U13140 ( .A(b[2053]), .B(n11095), .Z(n11096) );
  XNOR U13141 ( .A(b[2053]), .B(n11097), .Z(c[2053]) );
  XNOR U13142 ( .A(a[2053]), .B(n11098), .Z(n11097) );
  IV U13143 ( .A(n11095), .Z(n11098) );
  XOR U13144 ( .A(n11099), .B(n11100), .Z(n11095) );
  ANDN U13145 ( .B(n11101), .A(n11102), .Z(n11099) );
  XNOR U13146 ( .A(b[2052]), .B(n11100), .Z(n11101) );
  XNOR U13147 ( .A(b[2052]), .B(n11102), .Z(c[2052]) );
  XNOR U13148 ( .A(a[2052]), .B(n11103), .Z(n11102) );
  IV U13149 ( .A(n11100), .Z(n11103) );
  XOR U13150 ( .A(n11104), .B(n11105), .Z(n11100) );
  ANDN U13151 ( .B(n11106), .A(n11107), .Z(n11104) );
  XNOR U13152 ( .A(b[2051]), .B(n11105), .Z(n11106) );
  XNOR U13153 ( .A(b[2051]), .B(n11107), .Z(c[2051]) );
  XNOR U13154 ( .A(a[2051]), .B(n11108), .Z(n11107) );
  IV U13155 ( .A(n11105), .Z(n11108) );
  XOR U13156 ( .A(n11109), .B(n11110), .Z(n11105) );
  ANDN U13157 ( .B(n11111), .A(n11112), .Z(n11109) );
  XNOR U13158 ( .A(b[2050]), .B(n11110), .Z(n11111) );
  XNOR U13159 ( .A(b[2050]), .B(n11112), .Z(c[2050]) );
  XNOR U13160 ( .A(a[2050]), .B(n11113), .Z(n11112) );
  IV U13161 ( .A(n11110), .Z(n11113) );
  XOR U13162 ( .A(n11114), .B(n11115), .Z(n11110) );
  ANDN U13163 ( .B(n11116), .A(n11117), .Z(n11114) );
  XNOR U13164 ( .A(b[2049]), .B(n11115), .Z(n11116) );
  XNOR U13165 ( .A(b[204]), .B(n11118), .Z(c[204]) );
  XNOR U13166 ( .A(b[2049]), .B(n11117), .Z(c[2049]) );
  XNOR U13167 ( .A(a[2049]), .B(n11119), .Z(n11117) );
  IV U13168 ( .A(n11115), .Z(n11119) );
  XOR U13169 ( .A(n11120), .B(n11121), .Z(n11115) );
  ANDN U13170 ( .B(n11122), .A(n11123), .Z(n11120) );
  XNOR U13171 ( .A(b[2048]), .B(n11121), .Z(n11122) );
  XNOR U13172 ( .A(b[2048]), .B(n11123), .Z(c[2048]) );
  XNOR U13173 ( .A(a[2048]), .B(n11124), .Z(n11123) );
  IV U13174 ( .A(n11121), .Z(n11124) );
  XOR U13175 ( .A(n11125), .B(n11126), .Z(n11121) );
  ANDN U13176 ( .B(n11127), .A(n11128), .Z(n11125) );
  XNOR U13177 ( .A(b[2047]), .B(n11126), .Z(n11127) );
  XNOR U13178 ( .A(b[2047]), .B(n11128), .Z(c[2047]) );
  XNOR U13179 ( .A(a[2047]), .B(n11129), .Z(n11128) );
  IV U13180 ( .A(n11126), .Z(n11129) );
  XOR U13181 ( .A(n11130), .B(n11131), .Z(n11126) );
  ANDN U13182 ( .B(n11132), .A(n11133), .Z(n11130) );
  XNOR U13183 ( .A(b[2046]), .B(n11131), .Z(n11132) );
  XNOR U13184 ( .A(b[2046]), .B(n11133), .Z(c[2046]) );
  XNOR U13185 ( .A(a[2046]), .B(n11134), .Z(n11133) );
  IV U13186 ( .A(n11131), .Z(n11134) );
  XOR U13187 ( .A(n11135), .B(n11136), .Z(n11131) );
  ANDN U13188 ( .B(n11137), .A(n11138), .Z(n11135) );
  XNOR U13189 ( .A(b[2045]), .B(n11136), .Z(n11137) );
  XNOR U13190 ( .A(b[2045]), .B(n11138), .Z(c[2045]) );
  XNOR U13191 ( .A(a[2045]), .B(n11139), .Z(n11138) );
  IV U13192 ( .A(n11136), .Z(n11139) );
  XOR U13193 ( .A(n11140), .B(n11141), .Z(n11136) );
  ANDN U13194 ( .B(n11142), .A(n11143), .Z(n11140) );
  XNOR U13195 ( .A(b[2044]), .B(n11141), .Z(n11142) );
  XNOR U13196 ( .A(b[2044]), .B(n11143), .Z(c[2044]) );
  XNOR U13197 ( .A(a[2044]), .B(n11144), .Z(n11143) );
  IV U13198 ( .A(n11141), .Z(n11144) );
  XOR U13199 ( .A(n11145), .B(n11146), .Z(n11141) );
  ANDN U13200 ( .B(n11147), .A(n11148), .Z(n11145) );
  XNOR U13201 ( .A(b[2043]), .B(n11146), .Z(n11147) );
  XNOR U13202 ( .A(b[2043]), .B(n11148), .Z(c[2043]) );
  XNOR U13203 ( .A(a[2043]), .B(n11149), .Z(n11148) );
  IV U13204 ( .A(n11146), .Z(n11149) );
  XOR U13205 ( .A(n11150), .B(n11151), .Z(n11146) );
  ANDN U13206 ( .B(n11152), .A(n11153), .Z(n11150) );
  XNOR U13207 ( .A(b[2042]), .B(n11151), .Z(n11152) );
  XNOR U13208 ( .A(b[2042]), .B(n11153), .Z(c[2042]) );
  XNOR U13209 ( .A(a[2042]), .B(n11154), .Z(n11153) );
  IV U13210 ( .A(n11151), .Z(n11154) );
  XOR U13211 ( .A(n11155), .B(n11156), .Z(n11151) );
  ANDN U13212 ( .B(n11157), .A(n11158), .Z(n11155) );
  XNOR U13213 ( .A(b[2041]), .B(n11156), .Z(n11157) );
  XNOR U13214 ( .A(b[2041]), .B(n11158), .Z(c[2041]) );
  XNOR U13215 ( .A(a[2041]), .B(n11159), .Z(n11158) );
  IV U13216 ( .A(n11156), .Z(n11159) );
  XOR U13217 ( .A(n11160), .B(n11161), .Z(n11156) );
  ANDN U13218 ( .B(n11162), .A(n11163), .Z(n11160) );
  XNOR U13219 ( .A(b[2040]), .B(n11161), .Z(n11162) );
  XNOR U13220 ( .A(b[2040]), .B(n11163), .Z(c[2040]) );
  XNOR U13221 ( .A(a[2040]), .B(n11164), .Z(n11163) );
  IV U13222 ( .A(n11161), .Z(n11164) );
  XOR U13223 ( .A(n11165), .B(n11166), .Z(n11161) );
  ANDN U13224 ( .B(n11167), .A(n11168), .Z(n11165) );
  XNOR U13225 ( .A(b[2039]), .B(n11166), .Z(n11167) );
  XNOR U13226 ( .A(b[203]), .B(n11169), .Z(c[203]) );
  XNOR U13227 ( .A(b[2039]), .B(n11168), .Z(c[2039]) );
  XNOR U13228 ( .A(a[2039]), .B(n11170), .Z(n11168) );
  IV U13229 ( .A(n11166), .Z(n11170) );
  XOR U13230 ( .A(n11171), .B(n11172), .Z(n11166) );
  ANDN U13231 ( .B(n11173), .A(n11174), .Z(n11171) );
  XNOR U13232 ( .A(b[2038]), .B(n11172), .Z(n11173) );
  XNOR U13233 ( .A(b[2038]), .B(n11174), .Z(c[2038]) );
  XNOR U13234 ( .A(a[2038]), .B(n11175), .Z(n11174) );
  IV U13235 ( .A(n11172), .Z(n11175) );
  XOR U13236 ( .A(n11176), .B(n11177), .Z(n11172) );
  ANDN U13237 ( .B(n11178), .A(n11179), .Z(n11176) );
  XNOR U13238 ( .A(b[2037]), .B(n11177), .Z(n11178) );
  XNOR U13239 ( .A(b[2037]), .B(n11179), .Z(c[2037]) );
  XNOR U13240 ( .A(a[2037]), .B(n11180), .Z(n11179) );
  IV U13241 ( .A(n11177), .Z(n11180) );
  XOR U13242 ( .A(n11181), .B(n11182), .Z(n11177) );
  ANDN U13243 ( .B(n11183), .A(n11184), .Z(n11181) );
  XNOR U13244 ( .A(b[2036]), .B(n11182), .Z(n11183) );
  XNOR U13245 ( .A(b[2036]), .B(n11184), .Z(c[2036]) );
  XNOR U13246 ( .A(a[2036]), .B(n11185), .Z(n11184) );
  IV U13247 ( .A(n11182), .Z(n11185) );
  XOR U13248 ( .A(n11186), .B(n11187), .Z(n11182) );
  ANDN U13249 ( .B(n11188), .A(n11189), .Z(n11186) );
  XNOR U13250 ( .A(b[2035]), .B(n11187), .Z(n11188) );
  XNOR U13251 ( .A(b[2035]), .B(n11189), .Z(c[2035]) );
  XNOR U13252 ( .A(a[2035]), .B(n11190), .Z(n11189) );
  IV U13253 ( .A(n11187), .Z(n11190) );
  XOR U13254 ( .A(n11191), .B(n11192), .Z(n11187) );
  ANDN U13255 ( .B(n11193), .A(n11194), .Z(n11191) );
  XNOR U13256 ( .A(b[2034]), .B(n11192), .Z(n11193) );
  XNOR U13257 ( .A(b[2034]), .B(n11194), .Z(c[2034]) );
  XNOR U13258 ( .A(a[2034]), .B(n11195), .Z(n11194) );
  IV U13259 ( .A(n11192), .Z(n11195) );
  XOR U13260 ( .A(n11196), .B(n11197), .Z(n11192) );
  ANDN U13261 ( .B(n11198), .A(n11199), .Z(n11196) );
  XNOR U13262 ( .A(b[2033]), .B(n11197), .Z(n11198) );
  XNOR U13263 ( .A(b[2033]), .B(n11199), .Z(c[2033]) );
  XNOR U13264 ( .A(a[2033]), .B(n11200), .Z(n11199) );
  IV U13265 ( .A(n11197), .Z(n11200) );
  XOR U13266 ( .A(n11201), .B(n11202), .Z(n11197) );
  ANDN U13267 ( .B(n11203), .A(n11204), .Z(n11201) );
  XNOR U13268 ( .A(b[2032]), .B(n11202), .Z(n11203) );
  XNOR U13269 ( .A(b[2032]), .B(n11204), .Z(c[2032]) );
  XNOR U13270 ( .A(a[2032]), .B(n11205), .Z(n11204) );
  IV U13271 ( .A(n11202), .Z(n11205) );
  XOR U13272 ( .A(n11206), .B(n11207), .Z(n11202) );
  ANDN U13273 ( .B(n11208), .A(n11209), .Z(n11206) );
  XNOR U13274 ( .A(b[2031]), .B(n11207), .Z(n11208) );
  XNOR U13275 ( .A(b[2031]), .B(n11209), .Z(c[2031]) );
  XNOR U13276 ( .A(a[2031]), .B(n11210), .Z(n11209) );
  IV U13277 ( .A(n11207), .Z(n11210) );
  XOR U13278 ( .A(n11211), .B(n11212), .Z(n11207) );
  ANDN U13279 ( .B(n11213), .A(n11214), .Z(n11211) );
  XNOR U13280 ( .A(b[2030]), .B(n11212), .Z(n11213) );
  XNOR U13281 ( .A(b[2030]), .B(n11214), .Z(c[2030]) );
  XNOR U13282 ( .A(a[2030]), .B(n11215), .Z(n11214) );
  IV U13283 ( .A(n11212), .Z(n11215) );
  XOR U13284 ( .A(n11216), .B(n11217), .Z(n11212) );
  ANDN U13285 ( .B(n11218), .A(n11219), .Z(n11216) );
  XNOR U13286 ( .A(b[2029]), .B(n11217), .Z(n11218) );
  XNOR U13287 ( .A(b[202]), .B(n11220), .Z(c[202]) );
  XNOR U13288 ( .A(b[2029]), .B(n11219), .Z(c[2029]) );
  XNOR U13289 ( .A(a[2029]), .B(n11221), .Z(n11219) );
  IV U13290 ( .A(n11217), .Z(n11221) );
  XOR U13291 ( .A(n11222), .B(n11223), .Z(n11217) );
  ANDN U13292 ( .B(n11224), .A(n11225), .Z(n11222) );
  XNOR U13293 ( .A(b[2028]), .B(n11223), .Z(n11224) );
  XNOR U13294 ( .A(b[2028]), .B(n11225), .Z(c[2028]) );
  XNOR U13295 ( .A(a[2028]), .B(n11226), .Z(n11225) );
  IV U13296 ( .A(n11223), .Z(n11226) );
  XOR U13297 ( .A(n11227), .B(n11228), .Z(n11223) );
  ANDN U13298 ( .B(n11229), .A(n11230), .Z(n11227) );
  XNOR U13299 ( .A(b[2027]), .B(n11228), .Z(n11229) );
  XNOR U13300 ( .A(b[2027]), .B(n11230), .Z(c[2027]) );
  XNOR U13301 ( .A(a[2027]), .B(n11231), .Z(n11230) );
  IV U13302 ( .A(n11228), .Z(n11231) );
  XOR U13303 ( .A(n11232), .B(n11233), .Z(n11228) );
  ANDN U13304 ( .B(n11234), .A(n11235), .Z(n11232) );
  XNOR U13305 ( .A(b[2026]), .B(n11233), .Z(n11234) );
  XNOR U13306 ( .A(b[2026]), .B(n11235), .Z(c[2026]) );
  XNOR U13307 ( .A(a[2026]), .B(n11236), .Z(n11235) );
  IV U13308 ( .A(n11233), .Z(n11236) );
  XOR U13309 ( .A(n11237), .B(n11238), .Z(n11233) );
  ANDN U13310 ( .B(n11239), .A(n11240), .Z(n11237) );
  XNOR U13311 ( .A(b[2025]), .B(n11238), .Z(n11239) );
  XNOR U13312 ( .A(b[2025]), .B(n11240), .Z(c[2025]) );
  XNOR U13313 ( .A(a[2025]), .B(n11241), .Z(n11240) );
  IV U13314 ( .A(n11238), .Z(n11241) );
  XOR U13315 ( .A(n11242), .B(n11243), .Z(n11238) );
  ANDN U13316 ( .B(n11244), .A(n11245), .Z(n11242) );
  XNOR U13317 ( .A(b[2024]), .B(n11243), .Z(n11244) );
  XNOR U13318 ( .A(b[2024]), .B(n11245), .Z(c[2024]) );
  XNOR U13319 ( .A(a[2024]), .B(n11246), .Z(n11245) );
  IV U13320 ( .A(n11243), .Z(n11246) );
  XOR U13321 ( .A(n11247), .B(n11248), .Z(n11243) );
  ANDN U13322 ( .B(n11249), .A(n11250), .Z(n11247) );
  XNOR U13323 ( .A(b[2023]), .B(n11248), .Z(n11249) );
  XNOR U13324 ( .A(b[2023]), .B(n11250), .Z(c[2023]) );
  XNOR U13325 ( .A(a[2023]), .B(n11251), .Z(n11250) );
  IV U13326 ( .A(n11248), .Z(n11251) );
  XOR U13327 ( .A(n11252), .B(n11253), .Z(n11248) );
  ANDN U13328 ( .B(n11254), .A(n11255), .Z(n11252) );
  XNOR U13329 ( .A(b[2022]), .B(n11253), .Z(n11254) );
  XNOR U13330 ( .A(b[2022]), .B(n11255), .Z(c[2022]) );
  XNOR U13331 ( .A(a[2022]), .B(n11256), .Z(n11255) );
  IV U13332 ( .A(n11253), .Z(n11256) );
  XOR U13333 ( .A(n11257), .B(n11258), .Z(n11253) );
  ANDN U13334 ( .B(n11259), .A(n11260), .Z(n11257) );
  XNOR U13335 ( .A(b[2021]), .B(n11258), .Z(n11259) );
  XNOR U13336 ( .A(b[2021]), .B(n11260), .Z(c[2021]) );
  XNOR U13337 ( .A(a[2021]), .B(n11261), .Z(n11260) );
  IV U13338 ( .A(n11258), .Z(n11261) );
  XOR U13339 ( .A(n11262), .B(n11263), .Z(n11258) );
  ANDN U13340 ( .B(n11264), .A(n11265), .Z(n11262) );
  XNOR U13341 ( .A(b[2020]), .B(n11263), .Z(n11264) );
  XNOR U13342 ( .A(b[2020]), .B(n11265), .Z(c[2020]) );
  XNOR U13343 ( .A(a[2020]), .B(n11266), .Z(n11265) );
  IV U13344 ( .A(n11263), .Z(n11266) );
  XOR U13345 ( .A(n11267), .B(n11268), .Z(n11263) );
  ANDN U13346 ( .B(n11269), .A(n11270), .Z(n11267) );
  XNOR U13347 ( .A(b[2019]), .B(n11268), .Z(n11269) );
  XNOR U13348 ( .A(b[201]), .B(n11271), .Z(c[201]) );
  XNOR U13349 ( .A(b[2019]), .B(n11270), .Z(c[2019]) );
  XNOR U13350 ( .A(a[2019]), .B(n11272), .Z(n11270) );
  IV U13351 ( .A(n11268), .Z(n11272) );
  XOR U13352 ( .A(n11273), .B(n11274), .Z(n11268) );
  ANDN U13353 ( .B(n11275), .A(n11276), .Z(n11273) );
  XNOR U13354 ( .A(b[2018]), .B(n11274), .Z(n11275) );
  XNOR U13355 ( .A(b[2018]), .B(n11276), .Z(c[2018]) );
  XNOR U13356 ( .A(a[2018]), .B(n11277), .Z(n11276) );
  IV U13357 ( .A(n11274), .Z(n11277) );
  XOR U13358 ( .A(n11278), .B(n11279), .Z(n11274) );
  ANDN U13359 ( .B(n11280), .A(n11281), .Z(n11278) );
  XNOR U13360 ( .A(b[2017]), .B(n11279), .Z(n11280) );
  XNOR U13361 ( .A(b[2017]), .B(n11281), .Z(c[2017]) );
  XNOR U13362 ( .A(a[2017]), .B(n11282), .Z(n11281) );
  IV U13363 ( .A(n11279), .Z(n11282) );
  XOR U13364 ( .A(n11283), .B(n11284), .Z(n11279) );
  ANDN U13365 ( .B(n11285), .A(n11286), .Z(n11283) );
  XNOR U13366 ( .A(b[2016]), .B(n11284), .Z(n11285) );
  XNOR U13367 ( .A(b[2016]), .B(n11286), .Z(c[2016]) );
  XNOR U13368 ( .A(a[2016]), .B(n11287), .Z(n11286) );
  IV U13369 ( .A(n11284), .Z(n11287) );
  XOR U13370 ( .A(n11288), .B(n11289), .Z(n11284) );
  ANDN U13371 ( .B(n11290), .A(n11291), .Z(n11288) );
  XNOR U13372 ( .A(b[2015]), .B(n11289), .Z(n11290) );
  XNOR U13373 ( .A(b[2015]), .B(n11291), .Z(c[2015]) );
  XNOR U13374 ( .A(a[2015]), .B(n11292), .Z(n11291) );
  IV U13375 ( .A(n11289), .Z(n11292) );
  XOR U13376 ( .A(n11293), .B(n11294), .Z(n11289) );
  ANDN U13377 ( .B(n11295), .A(n11296), .Z(n11293) );
  XNOR U13378 ( .A(b[2014]), .B(n11294), .Z(n11295) );
  XNOR U13379 ( .A(b[2014]), .B(n11296), .Z(c[2014]) );
  XNOR U13380 ( .A(a[2014]), .B(n11297), .Z(n11296) );
  IV U13381 ( .A(n11294), .Z(n11297) );
  XOR U13382 ( .A(n11298), .B(n11299), .Z(n11294) );
  ANDN U13383 ( .B(n11300), .A(n11301), .Z(n11298) );
  XNOR U13384 ( .A(b[2013]), .B(n11299), .Z(n11300) );
  XNOR U13385 ( .A(b[2013]), .B(n11301), .Z(c[2013]) );
  XNOR U13386 ( .A(a[2013]), .B(n11302), .Z(n11301) );
  IV U13387 ( .A(n11299), .Z(n11302) );
  XOR U13388 ( .A(n11303), .B(n11304), .Z(n11299) );
  ANDN U13389 ( .B(n11305), .A(n11306), .Z(n11303) );
  XNOR U13390 ( .A(b[2012]), .B(n11304), .Z(n11305) );
  XNOR U13391 ( .A(b[2012]), .B(n11306), .Z(c[2012]) );
  XNOR U13392 ( .A(a[2012]), .B(n11307), .Z(n11306) );
  IV U13393 ( .A(n11304), .Z(n11307) );
  XOR U13394 ( .A(n11308), .B(n11309), .Z(n11304) );
  ANDN U13395 ( .B(n11310), .A(n11311), .Z(n11308) );
  XNOR U13396 ( .A(b[2011]), .B(n11309), .Z(n11310) );
  XNOR U13397 ( .A(b[2011]), .B(n11311), .Z(c[2011]) );
  XNOR U13398 ( .A(a[2011]), .B(n11312), .Z(n11311) );
  IV U13399 ( .A(n11309), .Z(n11312) );
  XOR U13400 ( .A(n11313), .B(n11314), .Z(n11309) );
  ANDN U13401 ( .B(n11315), .A(n11316), .Z(n11313) );
  XNOR U13402 ( .A(b[2010]), .B(n11314), .Z(n11315) );
  XNOR U13403 ( .A(b[2010]), .B(n11316), .Z(c[2010]) );
  XNOR U13404 ( .A(a[2010]), .B(n11317), .Z(n11316) );
  IV U13405 ( .A(n11314), .Z(n11317) );
  XOR U13406 ( .A(n11318), .B(n11319), .Z(n11314) );
  ANDN U13407 ( .B(n11320), .A(n11321), .Z(n11318) );
  XNOR U13408 ( .A(b[2009]), .B(n11319), .Z(n11320) );
  XNOR U13409 ( .A(b[200]), .B(n11322), .Z(c[200]) );
  XNOR U13410 ( .A(b[2009]), .B(n11321), .Z(c[2009]) );
  XNOR U13411 ( .A(a[2009]), .B(n11323), .Z(n11321) );
  IV U13412 ( .A(n11319), .Z(n11323) );
  XOR U13413 ( .A(n11324), .B(n11325), .Z(n11319) );
  ANDN U13414 ( .B(n11326), .A(n11327), .Z(n11324) );
  XNOR U13415 ( .A(b[2008]), .B(n11325), .Z(n11326) );
  XNOR U13416 ( .A(b[2008]), .B(n11327), .Z(c[2008]) );
  XNOR U13417 ( .A(a[2008]), .B(n11328), .Z(n11327) );
  IV U13418 ( .A(n11325), .Z(n11328) );
  XOR U13419 ( .A(n11329), .B(n11330), .Z(n11325) );
  ANDN U13420 ( .B(n11331), .A(n11332), .Z(n11329) );
  XNOR U13421 ( .A(b[2007]), .B(n11330), .Z(n11331) );
  XNOR U13422 ( .A(b[2007]), .B(n11332), .Z(c[2007]) );
  XNOR U13423 ( .A(a[2007]), .B(n11333), .Z(n11332) );
  IV U13424 ( .A(n11330), .Z(n11333) );
  XOR U13425 ( .A(n11334), .B(n11335), .Z(n11330) );
  ANDN U13426 ( .B(n11336), .A(n11337), .Z(n11334) );
  XNOR U13427 ( .A(b[2006]), .B(n11335), .Z(n11336) );
  XNOR U13428 ( .A(b[2006]), .B(n11337), .Z(c[2006]) );
  XNOR U13429 ( .A(a[2006]), .B(n11338), .Z(n11337) );
  IV U13430 ( .A(n11335), .Z(n11338) );
  XOR U13431 ( .A(n11339), .B(n11340), .Z(n11335) );
  ANDN U13432 ( .B(n11341), .A(n11342), .Z(n11339) );
  XNOR U13433 ( .A(b[2005]), .B(n11340), .Z(n11341) );
  XNOR U13434 ( .A(b[2005]), .B(n11342), .Z(c[2005]) );
  XNOR U13435 ( .A(a[2005]), .B(n11343), .Z(n11342) );
  IV U13436 ( .A(n11340), .Z(n11343) );
  XOR U13437 ( .A(n11344), .B(n11345), .Z(n11340) );
  ANDN U13438 ( .B(n11346), .A(n11347), .Z(n11344) );
  XNOR U13439 ( .A(b[2004]), .B(n11345), .Z(n11346) );
  XNOR U13440 ( .A(b[2004]), .B(n11347), .Z(c[2004]) );
  XNOR U13441 ( .A(a[2004]), .B(n11348), .Z(n11347) );
  IV U13442 ( .A(n11345), .Z(n11348) );
  XOR U13443 ( .A(n11349), .B(n11350), .Z(n11345) );
  ANDN U13444 ( .B(n11351), .A(n11352), .Z(n11349) );
  XNOR U13445 ( .A(b[2003]), .B(n11350), .Z(n11351) );
  XNOR U13446 ( .A(b[2003]), .B(n11352), .Z(c[2003]) );
  XNOR U13447 ( .A(a[2003]), .B(n11353), .Z(n11352) );
  IV U13448 ( .A(n11350), .Z(n11353) );
  XOR U13449 ( .A(n11354), .B(n11355), .Z(n11350) );
  ANDN U13450 ( .B(n11356), .A(n11357), .Z(n11354) );
  XNOR U13451 ( .A(b[2002]), .B(n11355), .Z(n11356) );
  XNOR U13452 ( .A(b[2002]), .B(n11357), .Z(c[2002]) );
  XNOR U13453 ( .A(a[2002]), .B(n11358), .Z(n11357) );
  IV U13454 ( .A(n11355), .Z(n11358) );
  XOR U13455 ( .A(n11359), .B(n11360), .Z(n11355) );
  ANDN U13456 ( .B(n11361), .A(n11362), .Z(n11359) );
  XNOR U13457 ( .A(b[2001]), .B(n11360), .Z(n11361) );
  XNOR U13458 ( .A(b[2001]), .B(n11362), .Z(c[2001]) );
  XNOR U13459 ( .A(a[2001]), .B(n11363), .Z(n11362) );
  IV U13460 ( .A(n11360), .Z(n11363) );
  XOR U13461 ( .A(n11364), .B(n11365), .Z(n11360) );
  ANDN U13462 ( .B(n11366), .A(n11367), .Z(n11364) );
  XNOR U13463 ( .A(b[2000]), .B(n11365), .Z(n11366) );
  XNOR U13464 ( .A(b[2000]), .B(n11367), .Z(c[2000]) );
  XNOR U13465 ( .A(a[2000]), .B(n11368), .Z(n11367) );
  IV U13466 ( .A(n11365), .Z(n11368) );
  XOR U13467 ( .A(n11369), .B(n11370), .Z(n11365) );
  ANDN U13468 ( .B(n11371), .A(n11372), .Z(n11369) );
  XNOR U13469 ( .A(b[1999]), .B(n11370), .Z(n11371) );
  XNOR U13470 ( .A(b[1]), .B(n11373), .Z(c[1]) );
  XNOR U13471 ( .A(b[19]), .B(n11374), .Z(c[19]) );
  XNOR U13472 ( .A(b[199]), .B(n11375), .Z(c[199]) );
  XNOR U13473 ( .A(b[1999]), .B(n11372), .Z(c[1999]) );
  XNOR U13474 ( .A(a[1999]), .B(n11376), .Z(n11372) );
  IV U13475 ( .A(n11370), .Z(n11376) );
  XOR U13476 ( .A(n11377), .B(n11378), .Z(n11370) );
  ANDN U13477 ( .B(n11379), .A(n11380), .Z(n11377) );
  XNOR U13478 ( .A(b[1998]), .B(n11378), .Z(n11379) );
  XNOR U13479 ( .A(b[1998]), .B(n11380), .Z(c[1998]) );
  XNOR U13480 ( .A(a[1998]), .B(n11381), .Z(n11380) );
  IV U13481 ( .A(n11378), .Z(n11381) );
  XOR U13482 ( .A(n11382), .B(n11383), .Z(n11378) );
  ANDN U13483 ( .B(n11384), .A(n11385), .Z(n11382) );
  XNOR U13484 ( .A(b[1997]), .B(n11383), .Z(n11384) );
  XNOR U13485 ( .A(b[1997]), .B(n11385), .Z(c[1997]) );
  XNOR U13486 ( .A(a[1997]), .B(n11386), .Z(n11385) );
  IV U13487 ( .A(n11383), .Z(n11386) );
  XOR U13488 ( .A(n11387), .B(n11388), .Z(n11383) );
  ANDN U13489 ( .B(n11389), .A(n11390), .Z(n11387) );
  XNOR U13490 ( .A(b[1996]), .B(n11388), .Z(n11389) );
  XNOR U13491 ( .A(b[1996]), .B(n11390), .Z(c[1996]) );
  XNOR U13492 ( .A(a[1996]), .B(n11391), .Z(n11390) );
  IV U13493 ( .A(n11388), .Z(n11391) );
  XOR U13494 ( .A(n11392), .B(n11393), .Z(n11388) );
  ANDN U13495 ( .B(n11394), .A(n11395), .Z(n11392) );
  XNOR U13496 ( .A(b[1995]), .B(n11393), .Z(n11394) );
  XNOR U13497 ( .A(b[1995]), .B(n11395), .Z(c[1995]) );
  XNOR U13498 ( .A(a[1995]), .B(n11396), .Z(n11395) );
  IV U13499 ( .A(n11393), .Z(n11396) );
  XOR U13500 ( .A(n11397), .B(n11398), .Z(n11393) );
  ANDN U13501 ( .B(n11399), .A(n11400), .Z(n11397) );
  XNOR U13502 ( .A(b[1994]), .B(n11398), .Z(n11399) );
  XNOR U13503 ( .A(b[1994]), .B(n11400), .Z(c[1994]) );
  XNOR U13504 ( .A(a[1994]), .B(n11401), .Z(n11400) );
  IV U13505 ( .A(n11398), .Z(n11401) );
  XOR U13506 ( .A(n11402), .B(n11403), .Z(n11398) );
  ANDN U13507 ( .B(n11404), .A(n11405), .Z(n11402) );
  XNOR U13508 ( .A(b[1993]), .B(n11403), .Z(n11404) );
  XNOR U13509 ( .A(b[1993]), .B(n11405), .Z(c[1993]) );
  XNOR U13510 ( .A(a[1993]), .B(n11406), .Z(n11405) );
  IV U13511 ( .A(n11403), .Z(n11406) );
  XOR U13512 ( .A(n11407), .B(n11408), .Z(n11403) );
  ANDN U13513 ( .B(n11409), .A(n11410), .Z(n11407) );
  XNOR U13514 ( .A(b[1992]), .B(n11408), .Z(n11409) );
  XNOR U13515 ( .A(b[1992]), .B(n11410), .Z(c[1992]) );
  XNOR U13516 ( .A(a[1992]), .B(n11411), .Z(n11410) );
  IV U13517 ( .A(n11408), .Z(n11411) );
  XOR U13518 ( .A(n11412), .B(n11413), .Z(n11408) );
  ANDN U13519 ( .B(n11414), .A(n11415), .Z(n11412) );
  XNOR U13520 ( .A(b[1991]), .B(n11413), .Z(n11414) );
  XNOR U13521 ( .A(b[1991]), .B(n11415), .Z(c[1991]) );
  XNOR U13522 ( .A(a[1991]), .B(n11416), .Z(n11415) );
  IV U13523 ( .A(n11413), .Z(n11416) );
  XOR U13524 ( .A(n11417), .B(n11418), .Z(n11413) );
  ANDN U13525 ( .B(n11419), .A(n11420), .Z(n11417) );
  XNOR U13526 ( .A(b[1990]), .B(n11418), .Z(n11419) );
  XNOR U13527 ( .A(b[1990]), .B(n11420), .Z(c[1990]) );
  XNOR U13528 ( .A(a[1990]), .B(n11421), .Z(n11420) );
  IV U13529 ( .A(n11418), .Z(n11421) );
  XOR U13530 ( .A(n11422), .B(n11423), .Z(n11418) );
  ANDN U13531 ( .B(n11424), .A(n11425), .Z(n11422) );
  XNOR U13532 ( .A(b[1989]), .B(n11423), .Z(n11424) );
  XNOR U13533 ( .A(b[198]), .B(n11426), .Z(c[198]) );
  XNOR U13534 ( .A(b[1989]), .B(n11425), .Z(c[1989]) );
  XNOR U13535 ( .A(a[1989]), .B(n11427), .Z(n11425) );
  IV U13536 ( .A(n11423), .Z(n11427) );
  XOR U13537 ( .A(n11428), .B(n11429), .Z(n11423) );
  ANDN U13538 ( .B(n11430), .A(n11431), .Z(n11428) );
  XNOR U13539 ( .A(b[1988]), .B(n11429), .Z(n11430) );
  XNOR U13540 ( .A(b[1988]), .B(n11431), .Z(c[1988]) );
  XNOR U13541 ( .A(a[1988]), .B(n11432), .Z(n11431) );
  IV U13542 ( .A(n11429), .Z(n11432) );
  XOR U13543 ( .A(n11433), .B(n11434), .Z(n11429) );
  ANDN U13544 ( .B(n11435), .A(n11436), .Z(n11433) );
  XNOR U13545 ( .A(b[1987]), .B(n11434), .Z(n11435) );
  XNOR U13546 ( .A(b[1987]), .B(n11436), .Z(c[1987]) );
  XNOR U13547 ( .A(a[1987]), .B(n11437), .Z(n11436) );
  IV U13548 ( .A(n11434), .Z(n11437) );
  XOR U13549 ( .A(n11438), .B(n11439), .Z(n11434) );
  ANDN U13550 ( .B(n11440), .A(n11441), .Z(n11438) );
  XNOR U13551 ( .A(b[1986]), .B(n11439), .Z(n11440) );
  XNOR U13552 ( .A(b[1986]), .B(n11441), .Z(c[1986]) );
  XNOR U13553 ( .A(a[1986]), .B(n11442), .Z(n11441) );
  IV U13554 ( .A(n11439), .Z(n11442) );
  XOR U13555 ( .A(n11443), .B(n11444), .Z(n11439) );
  ANDN U13556 ( .B(n11445), .A(n11446), .Z(n11443) );
  XNOR U13557 ( .A(b[1985]), .B(n11444), .Z(n11445) );
  XNOR U13558 ( .A(b[1985]), .B(n11446), .Z(c[1985]) );
  XNOR U13559 ( .A(a[1985]), .B(n11447), .Z(n11446) );
  IV U13560 ( .A(n11444), .Z(n11447) );
  XOR U13561 ( .A(n11448), .B(n11449), .Z(n11444) );
  ANDN U13562 ( .B(n11450), .A(n11451), .Z(n11448) );
  XNOR U13563 ( .A(b[1984]), .B(n11449), .Z(n11450) );
  XNOR U13564 ( .A(b[1984]), .B(n11451), .Z(c[1984]) );
  XNOR U13565 ( .A(a[1984]), .B(n11452), .Z(n11451) );
  IV U13566 ( .A(n11449), .Z(n11452) );
  XOR U13567 ( .A(n11453), .B(n11454), .Z(n11449) );
  ANDN U13568 ( .B(n11455), .A(n11456), .Z(n11453) );
  XNOR U13569 ( .A(b[1983]), .B(n11454), .Z(n11455) );
  XNOR U13570 ( .A(b[1983]), .B(n11456), .Z(c[1983]) );
  XNOR U13571 ( .A(a[1983]), .B(n11457), .Z(n11456) );
  IV U13572 ( .A(n11454), .Z(n11457) );
  XOR U13573 ( .A(n11458), .B(n11459), .Z(n11454) );
  ANDN U13574 ( .B(n11460), .A(n11461), .Z(n11458) );
  XNOR U13575 ( .A(b[1982]), .B(n11459), .Z(n11460) );
  XNOR U13576 ( .A(b[1982]), .B(n11461), .Z(c[1982]) );
  XNOR U13577 ( .A(a[1982]), .B(n11462), .Z(n11461) );
  IV U13578 ( .A(n11459), .Z(n11462) );
  XOR U13579 ( .A(n11463), .B(n11464), .Z(n11459) );
  ANDN U13580 ( .B(n11465), .A(n11466), .Z(n11463) );
  XNOR U13581 ( .A(b[1981]), .B(n11464), .Z(n11465) );
  XNOR U13582 ( .A(b[1981]), .B(n11466), .Z(c[1981]) );
  XNOR U13583 ( .A(a[1981]), .B(n11467), .Z(n11466) );
  IV U13584 ( .A(n11464), .Z(n11467) );
  XOR U13585 ( .A(n11468), .B(n11469), .Z(n11464) );
  ANDN U13586 ( .B(n11470), .A(n11471), .Z(n11468) );
  XNOR U13587 ( .A(b[1980]), .B(n11469), .Z(n11470) );
  XNOR U13588 ( .A(b[1980]), .B(n11471), .Z(c[1980]) );
  XNOR U13589 ( .A(a[1980]), .B(n11472), .Z(n11471) );
  IV U13590 ( .A(n11469), .Z(n11472) );
  XOR U13591 ( .A(n11473), .B(n11474), .Z(n11469) );
  ANDN U13592 ( .B(n11475), .A(n11476), .Z(n11473) );
  XNOR U13593 ( .A(b[1979]), .B(n11474), .Z(n11475) );
  XNOR U13594 ( .A(b[197]), .B(n11477), .Z(c[197]) );
  XNOR U13595 ( .A(b[1979]), .B(n11476), .Z(c[1979]) );
  XNOR U13596 ( .A(a[1979]), .B(n11478), .Z(n11476) );
  IV U13597 ( .A(n11474), .Z(n11478) );
  XOR U13598 ( .A(n11479), .B(n11480), .Z(n11474) );
  ANDN U13599 ( .B(n11481), .A(n11482), .Z(n11479) );
  XNOR U13600 ( .A(b[1978]), .B(n11480), .Z(n11481) );
  XNOR U13601 ( .A(b[1978]), .B(n11482), .Z(c[1978]) );
  XNOR U13602 ( .A(a[1978]), .B(n11483), .Z(n11482) );
  IV U13603 ( .A(n11480), .Z(n11483) );
  XOR U13604 ( .A(n11484), .B(n11485), .Z(n11480) );
  ANDN U13605 ( .B(n11486), .A(n11487), .Z(n11484) );
  XNOR U13606 ( .A(b[1977]), .B(n11485), .Z(n11486) );
  XNOR U13607 ( .A(b[1977]), .B(n11487), .Z(c[1977]) );
  XNOR U13608 ( .A(a[1977]), .B(n11488), .Z(n11487) );
  IV U13609 ( .A(n11485), .Z(n11488) );
  XOR U13610 ( .A(n11489), .B(n11490), .Z(n11485) );
  ANDN U13611 ( .B(n11491), .A(n11492), .Z(n11489) );
  XNOR U13612 ( .A(b[1976]), .B(n11490), .Z(n11491) );
  XNOR U13613 ( .A(b[1976]), .B(n11492), .Z(c[1976]) );
  XNOR U13614 ( .A(a[1976]), .B(n11493), .Z(n11492) );
  IV U13615 ( .A(n11490), .Z(n11493) );
  XOR U13616 ( .A(n11494), .B(n11495), .Z(n11490) );
  ANDN U13617 ( .B(n11496), .A(n11497), .Z(n11494) );
  XNOR U13618 ( .A(b[1975]), .B(n11495), .Z(n11496) );
  XNOR U13619 ( .A(b[1975]), .B(n11497), .Z(c[1975]) );
  XNOR U13620 ( .A(a[1975]), .B(n11498), .Z(n11497) );
  IV U13621 ( .A(n11495), .Z(n11498) );
  XOR U13622 ( .A(n11499), .B(n11500), .Z(n11495) );
  ANDN U13623 ( .B(n11501), .A(n11502), .Z(n11499) );
  XNOR U13624 ( .A(b[1974]), .B(n11500), .Z(n11501) );
  XNOR U13625 ( .A(b[1974]), .B(n11502), .Z(c[1974]) );
  XNOR U13626 ( .A(a[1974]), .B(n11503), .Z(n11502) );
  IV U13627 ( .A(n11500), .Z(n11503) );
  XOR U13628 ( .A(n11504), .B(n11505), .Z(n11500) );
  ANDN U13629 ( .B(n11506), .A(n11507), .Z(n11504) );
  XNOR U13630 ( .A(b[1973]), .B(n11505), .Z(n11506) );
  XNOR U13631 ( .A(b[1973]), .B(n11507), .Z(c[1973]) );
  XNOR U13632 ( .A(a[1973]), .B(n11508), .Z(n11507) );
  IV U13633 ( .A(n11505), .Z(n11508) );
  XOR U13634 ( .A(n11509), .B(n11510), .Z(n11505) );
  ANDN U13635 ( .B(n11511), .A(n11512), .Z(n11509) );
  XNOR U13636 ( .A(b[1972]), .B(n11510), .Z(n11511) );
  XNOR U13637 ( .A(b[1972]), .B(n11512), .Z(c[1972]) );
  XNOR U13638 ( .A(a[1972]), .B(n11513), .Z(n11512) );
  IV U13639 ( .A(n11510), .Z(n11513) );
  XOR U13640 ( .A(n11514), .B(n11515), .Z(n11510) );
  ANDN U13641 ( .B(n11516), .A(n11517), .Z(n11514) );
  XNOR U13642 ( .A(b[1971]), .B(n11515), .Z(n11516) );
  XNOR U13643 ( .A(b[1971]), .B(n11517), .Z(c[1971]) );
  XNOR U13644 ( .A(a[1971]), .B(n11518), .Z(n11517) );
  IV U13645 ( .A(n11515), .Z(n11518) );
  XOR U13646 ( .A(n11519), .B(n11520), .Z(n11515) );
  ANDN U13647 ( .B(n11521), .A(n11522), .Z(n11519) );
  XNOR U13648 ( .A(b[1970]), .B(n11520), .Z(n11521) );
  XNOR U13649 ( .A(b[1970]), .B(n11522), .Z(c[1970]) );
  XNOR U13650 ( .A(a[1970]), .B(n11523), .Z(n11522) );
  IV U13651 ( .A(n11520), .Z(n11523) );
  XOR U13652 ( .A(n11524), .B(n11525), .Z(n11520) );
  ANDN U13653 ( .B(n11526), .A(n11527), .Z(n11524) );
  XNOR U13654 ( .A(b[1969]), .B(n11525), .Z(n11526) );
  XNOR U13655 ( .A(b[196]), .B(n11528), .Z(c[196]) );
  XNOR U13656 ( .A(b[1969]), .B(n11527), .Z(c[1969]) );
  XNOR U13657 ( .A(a[1969]), .B(n11529), .Z(n11527) );
  IV U13658 ( .A(n11525), .Z(n11529) );
  XOR U13659 ( .A(n11530), .B(n11531), .Z(n11525) );
  ANDN U13660 ( .B(n11532), .A(n11533), .Z(n11530) );
  XNOR U13661 ( .A(b[1968]), .B(n11531), .Z(n11532) );
  XNOR U13662 ( .A(b[1968]), .B(n11533), .Z(c[1968]) );
  XNOR U13663 ( .A(a[1968]), .B(n11534), .Z(n11533) );
  IV U13664 ( .A(n11531), .Z(n11534) );
  XOR U13665 ( .A(n11535), .B(n11536), .Z(n11531) );
  ANDN U13666 ( .B(n11537), .A(n11538), .Z(n11535) );
  XNOR U13667 ( .A(b[1967]), .B(n11536), .Z(n11537) );
  XNOR U13668 ( .A(b[1967]), .B(n11538), .Z(c[1967]) );
  XNOR U13669 ( .A(a[1967]), .B(n11539), .Z(n11538) );
  IV U13670 ( .A(n11536), .Z(n11539) );
  XOR U13671 ( .A(n11540), .B(n11541), .Z(n11536) );
  ANDN U13672 ( .B(n11542), .A(n11543), .Z(n11540) );
  XNOR U13673 ( .A(b[1966]), .B(n11541), .Z(n11542) );
  XNOR U13674 ( .A(b[1966]), .B(n11543), .Z(c[1966]) );
  XNOR U13675 ( .A(a[1966]), .B(n11544), .Z(n11543) );
  IV U13676 ( .A(n11541), .Z(n11544) );
  XOR U13677 ( .A(n11545), .B(n11546), .Z(n11541) );
  ANDN U13678 ( .B(n11547), .A(n11548), .Z(n11545) );
  XNOR U13679 ( .A(b[1965]), .B(n11546), .Z(n11547) );
  XNOR U13680 ( .A(b[1965]), .B(n11548), .Z(c[1965]) );
  XNOR U13681 ( .A(a[1965]), .B(n11549), .Z(n11548) );
  IV U13682 ( .A(n11546), .Z(n11549) );
  XOR U13683 ( .A(n11550), .B(n11551), .Z(n11546) );
  ANDN U13684 ( .B(n11552), .A(n11553), .Z(n11550) );
  XNOR U13685 ( .A(b[1964]), .B(n11551), .Z(n11552) );
  XNOR U13686 ( .A(b[1964]), .B(n11553), .Z(c[1964]) );
  XNOR U13687 ( .A(a[1964]), .B(n11554), .Z(n11553) );
  IV U13688 ( .A(n11551), .Z(n11554) );
  XOR U13689 ( .A(n11555), .B(n11556), .Z(n11551) );
  ANDN U13690 ( .B(n11557), .A(n11558), .Z(n11555) );
  XNOR U13691 ( .A(b[1963]), .B(n11556), .Z(n11557) );
  XNOR U13692 ( .A(b[1963]), .B(n11558), .Z(c[1963]) );
  XNOR U13693 ( .A(a[1963]), .B(n11559), .Z(n11558) );
  IV U13694 ( .A(n11556), .Z(n11559) );
  XOR U13695 ( .A(n11560), .B(n11561), .Z(n11556) );
  ANDN U13696 ( .B(n11562), .A(n11563), .Z(n11560) );
  XNOR U13697 ( .A(b[1962]), .B(n11561), .Z(n11562) );
  XNOR U13698 ( .A(b[1962]), .B(n11563), .Z(c[1962]) );
  XNOR U13699 ( .A(a[1962]), .B(n11564), .Z(n11563) );
  IV U13700 ( .A(n11561), .Z(n11564) );
  XOR U13701 ( .A(n11565), .B(n11566), .Z(n11561) );
  ANDN U13702 ( .B(n11567), .A(n11568), .Z(n11565) );
  XNOR U13703 ( .A(b[1961]), .B(n11566), .Z(n11567) );
  XNOR U13704 ( .A(b[1961]), .B(n11568), .Z(c[1961]) );
  XNOR U13705 ( .A(a[1961]), .B(n11569), .Z(n11568) );
  IV U13706 ( .A(n11566), .Z(n11569) );
  XOR U13707 ( .A(n11570), .B(n11571), .Z(n11566) );
  ANDN U13708 ( .B(n11572), .A(n11573), .Z(n11570) );
  XNOR U13709 ( .A(b[1960]), .B(n11571), .Z(n11572) );
  XNOR U13710 ( .A(b[1960]), .B(n11573), .Z(c[1960]) );
  XNOR U13711 ( .A(a[1960]), .B(n11574), .Z(n11573) );
  IV U13712 ( .A(n11571), .Z(n11574) );
  XOR U13713 ( .A(n11575), .B(n11576), .Z(n11571) );
  ANDN U13714 ( .B(n11577), .A(n11578), .Z(n11575) );
  XNOR U13715 ( .A(b[1959]), .B(n11576), .Z(n11577) );
  XNOR U13716 ( .A(b[195]), .B(n11579), .Z(c[195]) );
  XNOR U13717 ( .A(b[1959]), .B(n11578), .Z(c[1959]) );
  XNOR U13718 ( .A(a[1959]), .B(n11580), .Z(n11578) );
  IV U13719 ( .A(n11576), .Z(n11580) );
  XOR U13720 ( .A(n11581), .B(n11582), .Z(n11576) );
  ANDN U13721 ( .B(n11583), .A(n11584), .Z(n11581) );
  XNOR U13722 ( .A(b[1958]), .B(n11582), .Z(n11583) );
  XNOR U13723 ( .A(b[1958]), .B(n11584), .Z(c[1958]) );
  XNOR U13724 ( .A(a[1958]), .B(n11585), .Z(n11584) );
  IV U13725 ( .A(n11582), .Z(n11585) );
  XOR U13726 ( .A(n11586), .B(n11587), .Z(n11582) );
  ANDN U13727 ( .B(n11588), .A(n11589), .Z(n11586) );
  XNOR U13728 ( .A(b[1957]), .B(n11587), .Z(n11588) );
  XNOR U13729 ( .A(b[1957]), .B(n11589), .Z(c[1957]) );
  XNOR U13730 ( .A(a[1957]), .B(n11590), .Z(n11589) );
  IV U13731 ( .A(n11587), .Z(n11590) );
  XOR U13732 ( .A(n11591), .B(n11592), .Z(n11587) );
  ANDN U13733 ( .B(n11593), .A(n11594), .Z(n11591) );
  XNOR U13734 ( .A(b[1956]), .B(n11592), .Z(n11593) );
  XNOR U13735 ( .A(b[1956]), .B(n11594), .Z(c[1956]) );
  XNOR U13736 ( .A(a[1956]), .B(n11595), .Z(n11594) );
  IV U13737 ( .A(n11592), .Z(n11595) );
  XOR U13738 ( .A(n11596), .B(n11597), .Z(n11592) );
  ANDN U13739 ( .B(n11598), .A(n11599), .Z(n11596) );
  XNOR U13740 ( .A(b[1955]), .B(n11597), .Z(n11598) );
  XNOR U13741 ( .A(b[1955]), .B(n11599), .Z(c[1955]) );
  XNOR U13742 ( .A(a[1955]), .B(n11600), .Z(n11599) );
  IV U13743 ( .A(n11597), .Z(n11600) );
  XOR U13744 ( .A(n11601), .B(n11602), .Z(n11597) );
  ANDN U13745 ( .B(n11603), .A(n11604), .Z(n11601) );
  XNOR U13746 ( .A(b[1954]), .B(n11602), .Z(n11603) );
  XNOR U13747 ( .A(b[1954]), .B(n11604), .Z(c[1954]) );
  XNOR U13748 ( .A(a[1954]), .B(n11605), .Z(n11604) );
  IV U13749 ( .A(n11602), .Z(n11605) );
  XOR U13750 ( .A(n11606), .B(n11607), .Z(n11602) );
  ANDN U13751 ( .B(n11608), .A(n11609), .Z(n11606) );
  XNOR U13752 ( .A(b[1953]), .B(n11607), .Z(n11608) );
  XNOR U13753 ( .A(b[1953]), .B(n11609), .Z(c[1953]) );
  XNOR U13754 ( .A(a[1953]), .B(n11610), .Z(n11609) );
  IV U13755 ( .A(n11607), .Z(n11610) );
  XOR U13756 ( .A(n11611), .B(n11612), .Z(n11607) );
  ANDN U13757 ( .B(n11613), .A(n11614), .Z(n11611) );
  XNOR U13758 ( .A(b[1952]), .B(n11612), .Z(n11613) );
  XNOR U13759 ( .A(b[1952]), .B(n11614), .Z(c[1952]) );
  XNOR U13760 ( .A(a[1952]), .B(n11615), .Z(n11614) );
  IV U13761 ( .A(n11612), .Z(n11615) );
  XOR U13762 ( .A(n11616), .B(n11617), .Z(n11612) );
  ANDN U13763 ( .B(n11618), .A(n11619), .Z(n11616) );
  XNOR U13764 ( .A(b[1951]), .B(n11617), .Z(n11618) );
  XNOR U13765 ( .A(b[1951]), .B(n11619), .Z(c[1951]) );
  XNOR U13766 ( .A(a[1951]), .B(n11620), .Z(n11619) );
  IV U13767 ( .A(n11617), .Z(n11620) );
  XOR U13768 ( .A(n11621), .B(n11622), .Z(n11617) );
  ANDN U13769 ( .B(n11623), .A(n11624), .Z(n11621) );
  XNOR U13770 ( .A(b[1950]), .B(n11622), .Z(n11623) );
  XNOR U13771 ( .A(b[1950]), .B(n11624), .Z(c[1950]) );
  XNOR U13772 ( .A(a[1950]), .B(n11625), .Z(n11624) );
  IV U13773 ( .A(n11622), .Z(n11625) );
  XOR U13774 ( .A(n11626), .B(n11627), .Z(n11622) );
  ANDN U13775 ( .B(n11628), .A(n11629), .Z(n11626) );
  XNOR U13776 ( .A(b[1949]), .B(n11627), .Z(n11628) );
  XNOR U13777 ( .A(b[194]), .B(n11630), .Z(c[194]) );
  XNOR U13778 ( .A(b[1949]), .B(n11629), .Z(c[1949]) );
  XNOR U13779 ( .A(a[1949]), .B(n11631), .Z(n11629) );
  IV U13780 ( .A(n11627), .Z(n11631) );
  XOR U13781 ( .A(n11632), .B(n11633), .Z(n11627) );
  ANDN U13782 ( .B(n11634), .A(n11635), .Z(n11632) );
  XNOR U13783 ( .A(b[1948]), .B(n11633), .Z(n11634) );
  XNOR U13784 ( .A(b[1948]), .B(n11635), .Z(c[1948]) );
  XNOR U13785 ( .A(a[1948]), .B(n11636), .Z(n11635) );
  IV U13786 ( .A(n11633), .Z(n11636) );
  XOR U13787 ( .A(n11637), .B(n11638), .Z(n11633) );
  ANDN U13788 ( .B(n11639), .A(n11640), .Z(n11637) );
  XNOR U13789 ( .A(b[1947]), .B(n11638), .Z(n11639) );
  XNOR U13790 ( .A(b[1947]), .B(n11640), .Z(c[1947]) );
  XNOR U13791 ( .A(a[1947]), .B(n11641), .Z(n11640) );
  IV U13792 ( .A(n11638), .Z(n11641) );
  XOR U13793 ( .A(n11642), .B(n11643), .Z(n11638) );
  ANDN U13794 ( .B(n11644), .A(n11645), .Z(n11642) );
  XNOR U13795 ( .A(b[1946]), .B(n11643), .Z(n11644) );
  XNOR U13796 ( .A(b[1946]), .B(n11645), .Z(c[1946]) );
  XNOR U13797 ( .A(a[1946]), .B(n11646), .Z(n11645) );
  IV U13798 ( .A(n11643), .Z(n11646) );
  XOR U13799 ( .A(n11647), .B(n11648), .Z(n11643) );
  ANDN U13800 ( .B(n11649), .A(n11650), .Z(n11647) );
  XNOR U13801 ( .A(b[1945]), .B(n11648), .Z(n11649) );
  XNOR U13802 ( .A(b[1945]), .B(n11650), .Z(c[1945]) );
  XNOR U13803 ( .A(a[1945]), .B(n11651), .Z(n11650) );
  IV U13804 ( .A(n11648), .Z(n11651) );
  XOR U13805 ( .A(n11652), .B(n11653), .Z(n11648) );
  ANDN U13806 ( .B(n11654), .A(n11655), .Z(n11652) );
  XNOR U13807 ( .A(b[1944]), .B(n11653), .Z(n11654) );
  XNOR U13808 ( .A(b[1944]), .B(n11655), .Z(c[1944]) );
  XNOR U13809 ( .A(a[1944]), .B(n11656), .Z(n11655) );
  IV U13810 ( .A(n11653), .Z(n11656) );
  XOR U13811 ( .A(n11657), .B(n11658), .Z(n11653) );
  ANDN U13812 ( .B(n11659), .A(n11660), .Z(n11657) );
  XNOR U13813 ( .A(b[1943]), .B(n11658), .Z(n11659) );
  XNOR U13814 ( .A(b[1943]), .B(n11660), .Z(c[1943]) );
  XNOR U13815 ( .A(a[1943]), .B(n11661), .Z(n11660) );
  IV U13816 ( .A(n11658), .Z(n11661) );
  XOR U13817 ( .A(n11662), .B(n11663), .Z(n11658) );
  ANDN U13818 ( .B(n11664), .A(n11665), .Z(n11662) );
  XNOR U13819 ( .A(b[1942]), .B(n11663), .Z(n11664) );
  XNOR U13820 ( .A(b[1942]), .B(n11665), .Z(c[1942]) );
  XNOR U13821 ( .A(a[1942]), .B(n11666), .Z(n11665) );
  IV U13822 ( .A(n11663), .Z(n11666) );
  XOR U13823 ( .A(n11667), .B(n11668), .Z(n11663) );
  ANDN U13824 ( .B(n11669), .A(n11670), .Z(n11667) );
  XNOR U13825 ( .A(b[1941]), .B(n11668), .Z(n11669) );
  XNOR U13826 ( .A(b[1941]), .B(n11670), .Z(c[1941]) );
  XNOR U13827 ( .A(a[1941]), .B(n11671), .Z(n11670) );
  IV U13828 ( .A(n11668), .Z(n11671) );
  XOR U13829 ( .A(n11672), .B(n11673), .Z(n11668) );
  ANDN U13830 ( .B(n11674), .A(n11675), .Z(n11672) );
  XNOR U13831 ( .A(b[1940]), .B(n11673), .Z(n11674) );
  XNOR U13832 ( .A(b[1940]), .B(n11675), .Z(c[1940]) );
  XNOR U13833 ( .A(a[1940]), .B(n11676), .Z(n11675) );
  IV U13834 ( .A(n11673), .Z(n11676) );
  XOR U13835 ( .A(n11677), .B(n11678), .Z(n11673) );
  ANDN U13836 ( .B(n11679), .A(n11680), .Z(n11677) );
  XNOR U13837 ( .A(b[1939]), .B(n11678), .Z(n11679) );
  XNOR U13838 ( .A(b[193]), .B(n11681), .Z(c[193]) );
  XNOR U13839 ( .A(b[1939]), .B(n11680), .Z(c[1939]) );
  XNOR U13840 ( .A(a[1939]), .B(n11682), .Z(n11680) );
  IV U13841 ( .A(n11678), .Z(n11682) );
  XOR U13842 ( .A(n11683), .B(n11684), .Z(n11678) );
  ANDN U13843 ( .B(n11685), .A(n11686), .Z(n11683) );
  XNOR U13844 ( .A(b[1938]), .B(n11684), .Z(n11685) );
  XNOR U13845 ( .A(b[1938]), .B(n11686), .Z(c[1938]) );
  XNOR U13846 ( .A(a[1938]), .B(n11687), .Z(n11686) );
  IV U13847 ( .A(n11684), .Z(n11687) );
  XOR U13848 ( .A(n11688), .B(n11689), .Z(n11684) );
  ANDN U13849 ( .B(n11690), .A(n11691), .Z(n11688) );
  XNOR U13850 ( .A(b[1937]), .B(n11689), .Z(n11690) );
  XNOR U13851 ( .A(b[1937]), .B(n11691), .Z(c[1937]) );
  XNOR U13852 ( .A(a[1937]), .B(n11692), .Z(n11691) );
  IV U13853 ( .A(n11689), .Z(n11692) );
  XOR U13854 ( .A(n11693), .B(n11694), .Z(n11689) );
  ANDN U13855 ( .B(n11695), .A(n11696), .Z(n11693) );
  XNOR U13856 ( .A(b[1936]), .B(n11694), .Z(n11695) );
  XNOR U13857 ( .A(b[1936]), .B(n11696), .Z(c[1936]) );
  XNOR U13858 ( .A(a[1936]), .B(n11697), .Z(n11696) );
  IV U13859 ( .A(n11694), .Z(n11697) );
  XOR U13860 ( .A(n11698), .B(n11699), .Z(n11694) );
  ANDN U13861 ( .B(n11700), .A(n11701), .Z(n11698) );
  XNOR U13862 ( .A(b[1935]), .B(n11699), .Z(n11700) );
  XNOR U13863 ( .A(b[1935]), .B(n11701), .Z(c[1935]) );
  XNOR U13864 ( .A(a[1935]), .B(n11702), .Z(n11701) );
  IV U13865 ( .A(n11699), .Z(n11702) );
  XOR U13866 ( .A(n11703), .B(n11704), .Z(n11699) );
  ANDN U13867 ( .B(n11705), .A(n11706), .Z(n11703) );
  XNOR U13868 ( .A(b[1934]), .B(n11704), .Z(n11705) );
  XNOR U13869 ( .A(b[1934]), .B(n11706), .Z(c[1934]) );
  XNOR U13870 ( .A(a[1934]), .B(n11707), .Z(n11706) );
  IV U13871 ( .A(n11704), .Z(n11707) );
  XOR U13872 ( .A(n11708), .B(n11709), .Z(n11704) );
  ANDN U13873 ( .B(n11710), .A(n11711), .Z(n11708) );
  XNOR U13874 ( .A(b[1933]), .B(n11709), .Z(n11710) );
  XNOR U13875 ( .A(b[1933]), .B(n11711), .Z(c[1933]) );
  XNOR U13876 ( .A(a[1933]), .B(n11712), .Z(n11711) );
  IV U13877 ( .A(n11709), .Z(n11712) );
  XOR U13878 ( .A(n11713), .B(n11714), .Z(n11709) );
  ANDN U13879 ( .B(n11715), .A(n11716), .Z(n11713) );
  XNOR U13880 ( .A(b[1932]), .B(n11714), .Z(n11715) );
  XNOR U13881 ( .A(b[1932]), .B(n11716), .Z(c[1932]) );
  XNOR U13882 ( .A(a[1932]), .B(n11717), .Z(n11716) );
  IV U13883 ( .A(n11714), .Z(n11717) );
  XOR U13884 ( .A(n11718), .B(n11719), .Z(n11714) );
  ANDN U13885 ( .B(n11720), .A(n11721), .Z(n11718) );
  XNOR U13886 ( .A(b[1931]), .B(n11719), .Z(n11720) );
  XNOR U13887 ( .A(b[1931]), .B(n11721), .Z(c[1931]) );
  XNOR U13888 ( .A(a[1931]), .B(n11722), .Z(n11721) );
  IV U13889 ( .A(n11719), .Z(n11722) );
  XOR U13890 ( .A(n11723), .B(n11724), .Z(n11719) );
  ANDN U13891 ( .B(n11725), .A(n11726), .Z(n11723) );
  XNOR U13892 ( .A(b[1930]), .B(n11724), .Z(n11725) );
  XNOR U13893 ( .A(b[1930]), .B(n11726), .Z(c[1930]) );
  XNOR U13894 ( .A(a[1930]), .B(n11727), .Z(n11726) );
  IV U13895 ( .A(n11724), .Z(n11727) );
  XOR U13896 ( .A(n11728), .B(n11729), .Z(n11724) );
  ANDN U13897 ( .B(n11730), .A(n11731), .Z(n11728) );
  XNOR U13898 ( .A(b[1929]), .B(n11729), .Z(n11730) );
  XNOR U13899 ( .A(b[192]), .B(n11732), .Z(c[192]) );
  XNOR U13900 ( .A(b[1929]), .B(n11731), .Z(c[1929]) );
  XNOR U13901 ( .A(a[1929]), .B(n11733), .Z(n11731) );
  IV U13902 ( .A(n11729), .Z(n11733) );
  XOR U13903 ( .A(n11734), .B(n11735), .Z(n11729) );
  ANDN U13904 ( .B(n11736), .A(n11737), .Z(n11734) );
  XNOR U13905 ( .A(b[1928]), .B(n11735), .Z(n11736) );
  XNOR U13906 ( .A(b[1928]), .B(n11737), .Z(c[1928]) );
  XNOR U13907 ( .A(a[1928]), .B(n11738), .Z(n11737) );
  IV U13908 ( .A(n11735), .Z(n11738) );
  XOR U13909 ( .A(n11739), .B(n11740), .Z(n11735) );
  ANDN U13910 ( .B(n11741), .A(n11742), .Z(n11739) );
  XNOR U13911 ( .A(b[1927]), .B(n11740), .Z(n11741) );
  XNOR U13912 ( .A(b[1927]), .B(n11742), .Z(c[1927]) );
  XNOR U13913 ( .A(a[1927]), .B(n11743), .Z(n11742) );
  IV U13914 ( .A(n11740), .Z(n11743) );
  XOR U13915 ( .A(n11744), .B(n11745), .Z(n11740) );
  ANDN U13916 ( .B(n11746), .A(n11747), .Z(n11744) );
  XNOR U13917 ( .A(b[1926]), .B(n11745), .Z(n11746) );
  XNOR U13918 ( .A(b[1926]), .B(n11747), .Z(c[1926]) );
  XNOR U13919 ( .A(a[1926]), .B(n11748), .Z(n11747) );
  IV U13920 ( .A(n11745), .Z(n11748) );
  XOR U13921 ( .A(n11749), .B(n11750), .Z(n11745) );
  ANDN U13922 ( .B(n11751), .A(n11752), .Z(n11749) );
  XNOR U13923 ( .A(b[1925]), .B(n11750), .Z(n11751) );
  XNOR U13924 ( .A(b[1925]), .B(n11752), .Z(c[1925]) );
  XNOR U13925 ( .A(a[1925]), .B(n11753), .Z(n11752) );
  IV U13926 ( .A(n11750), .Z(n11753) );
  XOR U13927 ( .A(n11754), .B(n11755), .Z(n11750) );
  ANDN U13928 ( .B(n11756), .A(n11757), .Z(n11754) );
  XNOR U13929 ( .A(b[1924]), .B(n11755), .Z(n11756) );
  XNOR U13930 ( .A(b[1924]), .B(n11757), .Z(c[1924]) );
  XNOR U13931 ( .A(a[1924]), .B(n11758), .Z(n11757) );
  IV U13932 ( .A(n11755), .Z(n11758) );
  XOR U13933 ( .A(n11759), .B(n11760), .Z(n11755) );
  ANDN U13934 ( .B(n11761), .A(n11762), .Z(n11759) );
  XNOR U13935 ( .A(b[1923]), .B(n11760), .Z(n11761) );
  XNOR U13936 ( .A(b[1923]), .B(n11762), .Z(c[1923]) );
  XNOR U13937 ( .A(a[1923]), .B(n11763), .Z(n11762) );
  IV U13938 ( .A(n11760), .Z(n11763) );
  XOR U13939 ( .A(n11764), .B(n11765), .Z(n11760) );
  ANDN U13940 ( .B(n11766), .A(n11767), .Z(n11764) );
  XNOR U13941 ( .A(b[1922]), .B(n11765), .Z(n11766) );
  XNOR U13942 ( .A(b[1922]), .B(n11767), .Z(c[1922]) );
  XNOR U13943 ( .A(a[1922]), .B(n11768), .Z(n11767) );
  IV U13944 ( .A(n11765), .Z(n11768) );
  XOR U13945 ( .A(n11769), .B(n11770), .Z(n11765) );
  ANDN U13946 ( .B(n11771), .A(n11772), .Z(n11769) );
  XNOR U13947 ( .A(b[1921]), .B(n11770), .Z(n11771) );
  XNOR U13948 ( .A(b[1921]), .B(n11772), .Z(c[1921]) );
  XNOR U13949 ( .A(a[1921]), .B(n11773), .Z(n11772) );
  IV U13950 ( .A(n11770), .Z(n11773) );
  XOR U13951 ( .A(n11774), .B(n11775), .Z(n11770) );
  ANDN U13952 ( .B(n11776), .A(n11777), .Z(n11774) );
  XNOR U13953 ( .A(b[1920]), .B(n11775), .Z(n11776) );
  XNOR U13954 ( .A(b[1920]), .B(n11777), .Z(c[1920]) );
  XNOR U13955 ( .A(a[1920]), .B(n11778), .Z(n11777) );
  IV U13956 ( .A(n11775), .Z(n11778) );
  XOR U13957 ( .A(n11779), .B(n11780), .Z(n11775) );
  ANDN U13958 ( .B(n11781), .A(n11782), .Z(n11779) );
  XNOR U13959 ( .A(b[1919]), .B(n11780), .Z(n11781) );
  XNOR U13960 ( .A(b[191]), .B(n11783), .Z(c[191]) );
  XNOR U13961 ( .A(b[1919]), .B(n11782), .Z(c[1919]) );
  XNOR U13962 ( .A(a[1919]), .B(n11784), .Z(n11782) );
  IV U13963 ( .A(n11780), .Z(n11784) );
  XOR U13964 ( .A(n11785), .B(n11786), .Z(n11780) );
  ANDN U13965 ( .B(n11787), .A(n11788), .Z(n11785) );
  XNOR U13966 ( .A(b[1918]), .B(n11786), .Z(n11787) );
  XNOR U13967 ( .A(b[1918]), .B(n11788), .Z(c[1918]) );
  XNOR U13968 ( .A(a[1918]), .B(n11789), .Z(n11788) );
  IV U13969 ( .A(n11786), .Z(n11789) );
  XOR U13970 ( .A(n11790), .B(n11791), .Z(n11786) );
  ANDN U13971 ( .B(n11792), .A(n11793), .Z(n11790) );
  XNOR U13972 ( .A(b[1917]), .B(n11791), .Z(n11792) );
  XNOR U13973 ( .A(b[1917]), .B(n11793), .Z(c[1917]) );
  XNOR U13974 ( .A(a[1917]), .B(n11794), .Z(n11793) );
  IV U13975 ( .A(n11791), .Z(n11794) );
  XOR U13976 ( .A(n11795), .B(n11796), .Z(n11791) );
  ANDN U13977 ( .B(n11797), .A(n11798), .Z(n11795) );
  XNOR U13978 ( .A(b[1916]), .B(n11796), .Z(n11797) );
  XNOR U13979 ( .A(b[1916]), .B(n11798), .Z(c[1916]) );
  XNOR U13980 ( .A(a[1916]), .B(n11799), .Z(n11798) );
  IV U13981 ( .A(n11796), .Z(n11799) );
  XOR U13982 ( .A(n11800), .B(n11801), .Z(n11796) );
  ANDN U13983 ( .B(n11802), .A(n11803), .Z(n11800) );
  XNOR U13984 ( .A(b[1915]), .B(n11801), .Z(n11802) );
  XNOR U13985 ( .A(b[1915]), .B(n11803), .Z(c[1915]) );
  XNOR U13986 ( .A(a[1915]), .B(n11804), .Z(n11803) );
  IV U13987 ( .A(n11801), .Z(n11804) );
  XOR U13988 ( .A(n11805), .B(n11806), .Z(n11801) );
  ANDN U13989 ( .B(n11807), .A(n11808), .Z(n11805) );
  XNOR U13990 ( .A(b[1914]), .B(n11806), .Z(n11807) );
  XNOR U13991 ( .A(b[1914]), .B(n11808), .Z(c[1914]) );
  XNOR U13992 ( .A(a[1914]), .B(n11809), .Z(n11808) );
  IV U13993 ( .A(n11806), .Z(n11809) );
  XOR U13994 ( .A(n11810), .B(n11811), .Z(n11806) );
  ANDN U13995 ( .B(n11812), .A(n11813), .Z(n11810) );
  XNOR U13996 ( .A(b[1913]), .B(n11811), .Z(n11812) );
  XNOR U13997 ( .A(b[1913]), .B(n11813), .Z(c[1913]) );
  XNOR U13998 ( .A(a[1913]), .B(n11814), .Z(n11813) );
  IV U13999 ( .A(n11811), .Z(n11814) );
  XOR U14000 ( .A(n11815), .B(n11816), .Z(n11811) );
  ANDN U14001 ( .B(n11817), .A(n11818), .Z(n11815) );
  XNOR U14002 ( .A(b[1912]), .B(n11816), .Z(n11817) );
  XNOR U14003 ( .A(b[1912]), .B(n11818), .Z(c[1912]) );
  XNOR U14004 ( .A(a[1912]), .B(n11819), .Z(n11818) );
  IV U14005 ( .A(n11816), .Z(n11819) );
  XOR U14006 ( .A(n11820), .B(n11821), .Z(n11816) );
  ANDN U14007 ( .B(n11822), .A(n11823), .Z(n11820) );
  XNOR U14008 ( .A(b[1911]), .B(n11821), .Z(n11822) );
  XNOR U14009 ( .A(b[1911]), .B(n11823), .Z(c[1911]) );
  XNOR U14010 ( .A(a[1911]), .B(n11824), .Z(n11823) );
  IV U14011 ( .A(n11821), .Z(n11824) );
  XOR U14012 ( .A(n11825), .B(n11826), .Z(n11821) );
  ANDN U14013 ( .B(n11827), .A(n11828), .Z(n11825) );
  XNOR U14014 ( .A(b[1910]), .B(n11826), .Z(n11827) );
  XNOR U14015 ( .A(b[1910]), .B(n11828), .Z(c[1910]) );
  XNOR U14016 ( .A(a[1910]), .B(n11829), .Z(n11828) );
  IV U14017 ( .A(n11826), .Z(n11829) );
  XOR U14018 ( .A(n11830), .B(n11831), .Z(n11826) );
  ANDN U14019 ( .B(n11832), .A(n11833), .Z(n11830) );
  XNOR U14020 ( .A(b[1909]), .B(n11831), .Z(n11832) );
  XNOR U14021 ( .A(b[190]), .B(n11834), .Z(c[190]) );
  XNOR U14022 ( .A(b[1909]), .B(n11833), .Z(c[1909]) );
  XNOR U14023 ( .A(a[1909]), .B(n11835), .Z(n11833) );
  IV U14024 ( .A(n11831), .Z(n11835) );
  XOR U14025 ( .A(n11836), .B(n11837), .Z(n11831) );
  ANDN U14026 ( .B(n11838), .A(n11839), .Z(n11836) );
  XNOR U14027 ( .A(b[1908]), .B(n11837), .Z(n11838) );
  XNOR U14028 ( .A(b[1908]), .B(n11839), .Z(c[1908]) );
  XNOR U14029 ( .A(a[1908]), .B(n11840), .Z(n11839) );
  IV U14030 ( .A(n11837), .Z(n11840) );
  XOR U14031 ( .A(n11841), .B(n11842), .Z(n11837) );
  ANDN U14032 ( .B(n11843), .A(n11844), .Z(n11841) );
  XNOR U14033 ( .A(b[1907]), .B(n11842), .Z(n11843) );
  XNOR U14034 ( .A(b[1907]), .B(n11844), .Z(c[1907]) );
  XNOR U14035 ( .A(a[1907]), .B(n11845), .Z(n11844) );
  IV U14036 ( .A(n11842), .Z(n11845) );
  XOR U14037 ( .A(n11846), .B(n11847), .Z(n11842) );
  ANDN U14038 ( .B(n11848), .A(n11849), .Z(n11846) );
  XNOR U14039 ( .A(b[1906]), .B(n11847), .Z(n11848) );
  XNOR U14040 ( .A(b[1906]), .B(n11849), .Z(c[1906]) );
  XNOR U14041 ( .A(a[1906]), .B(n11850), .Z(n11849) );
  IV U14042 ( .A(n11847), .Z(n11850) );
  XOR U14043 ( .A(n11851), .B(n11852), .Z(n11847) );
  ANDN U14044 ( .B(n11853), .A(n11854), .Z(n11851) );
  XNOR U14045 ( .A(b[1905]), .B(n11852), .Z(n11853) );
  XNOR U14046 ( .A(b[1905]), .B(n11854), .Z(c[1905]) );
  XNOR U14047 ( .A(a[1905]), .B(n11855), .Z(n11854) );
  IV U14048 ( .A(n11852), .Z(n11855) );
  XOR U14049 ( .A(n11856), .B(n11857), .Z(n11852) );
  ANDN U14050 ( .B(n11858), .A(n11859), .Z(n11856) );
  XNOR U14051 ( .A(b[1904]), .B(n11857), .Z(n11858) );
  XNOR U14052 ( .A(b[1904]), .B(n11859), .Z(c[1904]) );
  XNOR U14053 ( .A(a[1904]), .B(n11860), .Z(n11859) );
  IV U14054 ( .A(n11857), .Z(n11860) );
  XOR U14055 ( .A(n11861), .B(n11862), .Z(n11857) );
  ANDN U14056 ( .B(n11863), .A(n11864), .Z(n11861) );
  XNOR U14057 ( .A(b[1903]), .B(n11862), .Z(n11863) );
  XNOR U14058 ( .A(b[1903]), .B(n11864), .Z(c[1903]) );
  XNOR U14059 ( .A(a[1903]), .B(n11865), .Z(n11864) );
  IV U14060 ( .A(n11862), .Z(n11865) );
  XOR U14061 ( .A(n11866), .B(n11867), .Z(n11862) );
  ANDN U14062 ( .B(n11868), .A(n11869), .Z(n11866) );
  XNOR U14063 ( .A(b[1902]), .B(n11867), .Z(n11868) );
  XNOR U14064 ( .A(b[1902]), .B(n11869), .Z(c[1902]) );
  XNOR U14065 ( .A(a[1902]), .B(n11870), .Z(n11869) );
  IV U14066 ( .A(n11867), .Z(n11870) );
  XOR U14067 ( .A(n11871), .B(n11872), .Z(n11867) );
  ANDN U14068 ( .B(n11873), .A(n11874), .Z(n11871) );
  XNOR U14069 ( .A(b[1901]), .B(n11872), .Z(n11873) );
  XNOR U14070 ( .A(b[1901]), .B(n11874), .Z(c[1901]) );
  XNOR U14071 ( .A(a[1901]), .B(n11875), .Z(n11874) );
  IV U14072 ( .A(n11872), .Z(n11875) );
  XOR U14073 ( .A(n11876), .B(n11877), .Z(n11872) );
  ANDN U14074 ( .B(n11878), .A(n11879), .Z(n11876) );
  XNOR U14075 ( .A(b[1900]), .B(n11877), .Z(n11878) );
  XNOR U14076 ( .A(b[1900]), .B(n11879), .Z(c[1900]) );
  XNOR U14077 ( .A(a[1900]), .B(n11880), .Z(n11879) );
  IV U14078 ( .A(n11877), .Z(n11880) );
  XOR U14079 ( .A(n11881), .B(n11882), .Z(n11877) );
  ANDN U14080 ( .B(n11883), .A(n11884), .Z(n11881) );
  XNOR U14081 ( .A(b[1899]), .B(n11882), .Z(n11883) );
  XNOR U14082 ( .A(b[18]), .B(n11885), .Z(c[18]) );
  XNOR U14083 ( .A(b[189]), .B(n11886), .Z(c[189]) );
  XNOR U14084 ( .A(b[1899]), .B(n11884), .Z(c[1899]) );
  XNOR U14085 ( .A(a[1899]), .B(n11887), .Z(n11884) );
  IV U14086 ( .A(n11882), .Z(n11887) );
  XOR U14087 ( .A(n11888), .B(n11889), .Z(n11882) );
  ANDN U14088 ( .B(n11890), .A(n11891), .Z(n11888) );
  XNOR U14089 ( .A(b[1898]), .B(n11889), .Z(n11890) );
  XNOR U14090 ( .A(b[1898]), .B(n11891), .Z(c[1898]) );
  XNOR U14091 ( .A(a[1898]), .B(n11892), .Z(n11891) );
  IV U14092 ( .A(n11889), .Z(n11892) );
  XOR U14093 ( .A(n11893), .B(n11894), .Z(n11889) );
  ANDN U14094 ( .B(n11895), .A(n11896), .Z(n11893) );
  XNOR U14095 ( .A(b[1897]), .B(n11894), .Z(n11895) );
  XNOR U14096 ( .A(b[1897]), .B(n11896), .Z(c[1897]) );
  XNOR U14097 ( .A(a[1897]), .B(n11897), .Z(n11896) );
  IV U14098 ( .A(n11894), .Z(n11897) );
  XOR U14099 ( .A(n11898), .B(n11899), .Z(n11894) );
  ANDN U14100 ( .B(n11900), .A(n11901), .Z(n11898) );
  XNOR U14101 ( .A(b[1896]), .B(n11899), .Z(n11900) );
  XNOR U14102 ( .A(b[1896]), .B(n11901), .Z(c[1896]) );
  XNOR U14103 ( .A(a[1896]), .B(n11902), .Z(n11901) );
  IV U14104 ( .A(n11899), .Z(n11902) );
  XOR U14105 ( .A(n11903), .B(n11904), .Z(n11899) );
  ANDN U14106 ( .B(n11905), .A(n11906), .Z(n11903) );
  XNOR U14107 ( .A(b[1895]), .B(n11904), .Z(n11905) );
  XNOR U14108 ( .A(b[1895]), .B(n11906), .Z(c[1895]) );
  XNOR U14109 ( .A(a[1895]), .B(n11907), .Z(n11906) );
  IV U14110 ( .A(n11904), .Z(n11907) );
  XOR U14111 ( .A(n11908), .B(n11909), .Z(n11904) );
  ANDN U14112 ( .B(n11910), .A(n11911), .Z(n11908) );
  XNOR U14113 ( .A(b[1894]), .B(n11909), .Z(n11910) );
  XNOR U14114 ( .A(b[1894]), .B(n11911), .Z(c[1894]) );
  XNOR U14115 ( .A(a[1894]), .B(n11912), .Z(n11911) );
  IV U14116 ( .A(n11909), .Z(n11912) );
  XOR U14117 ( .A(n11913), .B(n11914), .Z(n11909) );
  ANDN U14118 ( .B(n11915), .A(n11916), .Z(n11913) );
  XNOR U14119 ( .A(b[1893]), .B(n11914), .Z(n11915) );
  XNOR U14120 ( .A(b[1893]), .B(n11916), .Z(c[1893]) );
  XNOR U14121 ( .A(a[1893]), .B(n11917), .Z(n11916) );
  IV U14122 ( .A(n11914), .Z(n11917) );
  XOR U14123 ( .A(n11918), .B(n11919), .Z(n11914) );
  ANDN U14124 ( .B(n11920), .A(n11921), .Z(n11918) );
  XNOR U14125 ( .A(b[1892]), .B(n11919), .Z(n11920) );
  XNOR U14126 ( .A(b[1892]), .B(n11921), .Z(c[1892]) );
  XNOR U14127 ( .A(a[1892]), .B(n11922), .Z(n11921) );
  IV U14128 ( .A(n11919), .Z(n11922) );
  XOR U14129 ( .A(n11923), .B(n11924), .Z(n11919) );
  ANDN U14130 ( .B(n11925), .A(n11926), .Z(n11923) );
  XNOR U14131 ( .A(b[1891]), .B(n11924), .Z(n11925) );
  XNOR U14132 ( .A(b[1891]), .B(n11926), .Z(c[1891]) );
  XNOR U14133 ( .A(a[1891]), .B(n11927), .Z(n11926) );
  IV U14134 ( .A(n11924), .Z(n11927) );
  XOR U14135 ( .A(n11928), .B(n11929), .Z(n11924) );
  ANDN U14136 ( .B(n11930), .A(n11931), .Z(n11928) );
  XNOR U14137 ( .A(b[1890]), .B(n11929), .Z(n11930) );
  XNOR U14138 ( .A(b[1890]), .B(n11931), .Z(c[1890]) );
  XNOR U14139 ( .A(a[1890]), .B(n11932), .Z(n11931) );
  IV U14140 ( .A(n11929), .Z(n11932) );
  XOR U14141 ( .A(n11933), .B(n11934), .Z(n11929) );
  ANDN U14142 ( .B(n11935), .A(n11936), .Z(n11933) );
  XNOR U14143 ( .A(b[1889]), .B(n11934), .Z(n11935) );
  XNOR U14144 ( .A(b[188]), .B(n11937), .Z(c[188]) );
  XNOR U14145 ( .A(b[1889]), .B(n11936), .Z(c[1889]) );
  XNOR U14146 ( .A(a[1889]), .B(n11938), .Z(n11936) );
  IV U14147 ( .A(n11934), .Z(n11938) );
  XOR U14148 ( .A(n11939), .B(n11940), .Z(n11934) );
  ANDN U14149 ( .B(n11941), .A(n11942), .Z(n11939) );
  XNOR U14150 ( .A(b[1888]), .B(n11940), .Z(n11941) );
  XNOR U14151 ( .A(b[1888]), .B(n11942), .Z(c[1888]) );
  XNOR U14152 ( .A(a[1888]), .B(n11943), .Z(n11942) );
  IV U14153 ( .A(n11940), .Z(n11943) );
  XOR U14154 ( .A(n11944), .B(n11945), .Z(n11940) );
  ANDN U14155 ( .B(n11946), .A(n11947), .Z(n11944) );
  XNOR U14156 ( .A(b[1887]), .B(n11945), .Z(n11946) );
  XNOR U14157 ( .A(b[1887]), .B(n11947), .Z(c[1887]) );
  XNOR U14158 ( .A(a[1887]), .B(n11948), .Z(n11947) );
  IV U14159 ( .A(n11945), .Z(n11948) );
  XOR U14160 ( .A(n11949), .B(n11950), .Z(n11945) );
  ANDN U14161 ( .B(n11951), .A(n11952), .Z(n11949) );
  XNOR U14162 ( .A(b[1886]), .B(n11950), .Z(n11951) );
  XNOR U14163 ( .A(b[1886]), .B(n11952), .Z(c[1886]) );
  XNOR U14164 ( .A(a[1886]), .B(n11953), .Z(n11952) );
  IV U14165 ( .A(n11950), .Z(n11953) );
  XOR U14166 ( .A(n11954), .B(n11955), .Z(n11950) );
  ANDN U14167 ( .B(n11956), .A(n11957), .Z(n11954) );
  XNOR U14168 ( .A(b[1885]), .B(n11955), .Z(n11956) );
  XNOR U14169 ( .A(b[1885]), .B(n11957), .Z(c[1885]) );
  XNOR U14170 ( .A(a[1885]), .B(n11958), .Z(n11957) );
  IV U14171 ( .A(n11955), .Z(n11958) );
  XOR U14172 ( .A(n11959), .B(n11960), .Z(n11955) );
  ANDN U14173 ( .B(n11961), .A(n11962), .Z(n11959) );
  XNOR U14174 ( .A(b[1884]), .B(n11960), .Z(n11961) );
  XNOR U14175 ( .A(b[1884]), .B(n11962), .Z(c[1884]) );
  XNOR U14176 ( .A(a[1884]), .B(n11963), .Z(n11962) );
  IV U14177 ( .A(n11960), .Z(n11963) );
  XOR U14178 ( .A(n11964), .B(n11965), .Z(n11960) );
  ANDN U14179 ( .B(n11966), .A(n11967), .Z(n11964) );
  XNOR U14180 ( .A(b[1883]), .B(n11965), .Z(n11966) );
  XNOR U14181 ( .A(b[1883]), .B(n11967), .Z(c[1883]) );
  XNOR U14182 ( .A(a[1883]), .B(n11968), .Z(n11967) );
  IV U14183 ( .A(n11965), .Z(n11968) );
  XOR U14184 ( .A(n11969), .B(n11970), .Z(n11965) );
  ANDN U14185 ( .B(n11971), .A(n11972), .Z(n11969) );
  XNOR U14186 ( .A(b[1882]), .B(n11970), .Z(n11971) );
  XNOR U14187 ( .A(b[1882]), .B(n11972), .Z(c[1882]) );
  XNOR U14188 ( .A(a[1882]), .B(n11973), .Z(n11972) );
  IV U14189 ( .A(n11970), .Z(n11973) );
  XOR U14190 ( .A(n11974), .B(n11975), .Z(n11970) );
  ANDN U14191 ( .B(n11976), .A(n11977), .Z(n11974) );
  XNOR U14192 ( .A(b[1881]), .B(n11975), .Z(n11976) );
  XNOR U14193 ( .A(b[1881]), .B(n11977), .Z(c[1881]) );
  XNOR U14194 ( .A(a[1881]), .B(n11978), .Z(n11977) );
  IV U14195 ( .A(n11975), .Z(n11978) );
  XOR U14196 ( .A(n11979), .B(n11980), .Z(n11975) );
  ANDN U14197 ( .B(n11981), .A(n11982), .Z(n11979) );
  XNOR U14198 ( .A(b[1880]), .B(n11980), .Z(n11981) );
  XNOR U14199 ( .A(b[1880]), .B(n11982), .Z(c[1880]) );
  XNOR U14200 ( .A(a[1880]), .B(n11983), .Z(n11982) );
  IV U14201 ( .A(n11980), .Z(n11983) );
  XOR U14202 ( .A(n11984), .B(n11985), .Z(n11980) );
  ANDN U14203 ( .B(n11986), .A(n11987), .Z(n11984) );
  XNOR U14204 ( .A(b[1879]), .B(n11985), .Z(n11986) );
  XNOR U14205 ( .A(b[187]), .B(n11988), .Z(c[187]) );
  XNOR U14206 ( .A(b[1879]), .B(n11987), .Z(c[1879]) );
  XNOR U14207 ( .A(a[1879]), .B(n11989), .Z(n11987) );
  IV U14208 ( .A(n11985), .Z(n11989) );
  XOR U14209 ( .A(n11990), .B(n11991), .Z(n11985) );
  ANDN U14210 ( .B(n11992), .A(n11993), .Z(n11990) );
  XNOR U14211 ( .A(b[1878]), .B(n11991), .Z(n11992) );
  XNOR U14212 ( .A(b[1878]), .B(n11993), .Z(c[1878]) );
  XNOR U14213 ( .A(a[1878]), .B(n11994), .Z(n11993) );
  IV U14214 ( .A(n11991), .Z(n11994) );
  XOR U14215 ( .A(n11995), .B(n11996), .Z(n11991) );
  ANDN U14216 ( .B(n11997), .A(n11998), .Z(n11995) );
  XNOR U14217 ( .A(b[1877]), .B(n11996), .Z(n11997) );
  XNOR U14218 ( .A(b[1877]), .B(n11998), .Z(c[1877]) );
  XNOR U14219 ( .A(a[1877]), .B(n11999), .Z(n11998) );
  IV U14220 ( .A(n11996), .Z(n11999) );
  XOR U14221 ( .A(n12000), .B(n12001), .Z(n11996) );
  ANDN U14222 ( .B(n12002), .A(n12003), .Z(n12000) );
  XNOR U14223 ( .A(b[1876]), .B(n12001), .Z(n12002) );
  XNOR U14224 ( .A(b[1876]), .B(n12003), .Z(c[1876]) );
  XNOR U14225 ( .A(a[1876]), .B(n12004), .Z(n12003) );
  IV U14226 ( .A(n12001), .Z(n12004) );
  XOR U14227 ( .A(n12005), .B(n12006), .Z(n12001) );
  ANDN U14228 ( .B(n12007), .A(n12008), .Z(n12005) );
  XNOR U14229 ( .A(b[1875]), .B(n12006), .Z(n12007) );
  XNOR U14230 ( .A(b[1875]), .B(n12008), .Z(c[1875]) );
  XNOR U14231 ( .A(a[1875]), .B(n12009), .Z(n12008) );
  IV U14232 ( .A(n12006), .Z(n12009) );
  XOR U14233 ( .A(n12010), .B(n12011), .Z(n12006) );
  ANDN U14234 ( .B(n12012), .A(n12013), .Z(n12010) );
  XNOR U14235 ( .A(b[1874]), .B(n12011), .Z(n12012) );
  XNOR U14236 ( .A(b[1874]), .B(n12013), .Z(c[1874]) );
  XNOR U14237 ( .A(a[1874]), .B(n12014), .Z(n12013) );
  IV U14238 ( .A(n12011), .Z(n12014) );
  XOR U14239 ( .A(n12015), .B(n12016), .Z(n12011) );
  ANDN U14240 ( .B(n12017), .A(n12018), .Z(n12015) );
  XNOR U14241 ( .A(b[1873]), .B(n12016), .Z(n12017) );
  XNOR U14242 ( .A(b[1873]), .B(n12018), .Z(c[1873]) );
  XNOR U14243 ( .A(a[1873]), .B(n12019), .Z(n12018) );
  IV U14244 ( .A(n12016), .Z(n12019) );
  XOR U14245 ( .A(n12020), .B(n12021), .Z(n12016) );
  ANDN U14246 ( .B(n12022), .A(n12023), .Z(n12020) );
  XNOR U14247 ( .A(b[1872]), .B(n12021), .Z(n12022) );
  XNOR U14248 ( .A(b[1872]), .B(n12023), .Z(c[1872]) );
  XNOR U14249 ( .A(a[1872]), .B(n12024), .Z(n12023) );
  IV U14250 ( .A(n12021), .Z(n12024) );
  XOR U14251 ( .A(n12025), .B(n12026), .Z(n12021) );
  ANDN U14252 ( .B(n12027), .A(n12028), .Z(n12025) );
  XNOR U14253 ( .A(b[1871]), .B(n12026), .Z(n12027) );
  XNOR U14254 ( .A(b[1871]), .B(n12028), .Z(c[1871]) );
  XNOR U14255 ( .A(a[1871]), .B(n12029), .Z(n12028) );
  IV U14256 ( .A(n12026), .Z(n12029) );
  XOR U14257 ( .A(n12030), .B(n12031), .Z(n12026) );
  ANDN U14258 ( .B(n12032), .A(n12033), .Z(n12030) );
  XNOR U14259 ( .A(b[1870]), .B(n12031), .Z(n12032) );
  XNOR U14260 ( .A(b[1870]), .B(n12033), .Z(c[1870]) );
  XNOR U14261 ( .A(a[1870]), .B(n12034), .Z(n12033) );
  IV U14262 ( .A(n12031), .Z(n12034) );
  XOR U14263 ( .A(n12035), .B(n12036), .Z(n12031) );
  ANDN U14264 ( .B(n12037), .A(n12038), .Z(n12035) );
  XNOR U14265 ( .A(b[1869]), .B(n12036), .Z(n12037) );
  XNOR U14266 ( .A(b[186]), .B(n12039), .Z(c[186]) );
  XNOR U14267 ( .A(b[1869]), .B(n12038), .Z(c[1869]) );
  XNOR U14268 ( .A(a[1869]), .B(n12040), .Z(n12038) );
  IV U14269 ( .A(n12036), .Z(n12040) );
  XOR U14270 ( .A(n12041), .B(n12042), .Z(n12036) );
  ANDN U14271 ( .B(n12043), .A(n12044), .Z(n12041) );
  XNOR U14272 ( .A(b[1868]), .B(n12042), .Z(n12043) );
  XNOR U14273 ( .A(b[1868]), .B(n12044), .Z(c[1868]) );
  XNOR U14274 ( .A(a[1868]), .B(n12045), .Z(n12044) );
  IV U14275 ( .A(n12042), .Z(n12045) );
  XOR U14276 ( .A(n12046), .B(n12047), .Z(n12042) );
  ANDN U14277 ( .B(n12048), .A(n12049), .Z(n12046) );
  XNOR U14278 ( .A(b[1867]), .B(n12047), .Z(n12048) );
  XNOR U14279 ( .A(b[1867]), .B(n12049), .Z(c[1867]) );
  XNOR U14280 ( .A(a[1867]), .B(n12050), .Z(n12049) );
  IV U14281 ( .A(n12047), .Z(n12050) );
  XOR U14282 ( .A(n12051), .B(n12052), .Z(n12047) );
  ANDN U14283 ( .B(n12053), .A(n12054), .Z(n12051) );
  XNOR U14284 ( .A(b[1866]), .B(n12052), .Z(n12053) );
  XNOR U14285 ( .A(b[1866]), .B(n12054), .Z(c[1866]) );
  XNOR U14286 ( .A(a[1866]), .B(n12055), .Z(n12054) );
  IV U14287 ( .A(n12052), .Z(n12055) );
  XOR U14288 ( .A(n12056), .B(n12057), .Z(n12052) );
  ANDN U14289 ( .B(n12058), .A(n12059), .Z(n12056) );
  XNOR U14290 ( .A(b[1865]), .B(n12057), .Z(n12058) );
  XNOR U14291 ( .A(b[1865]), .B(n12059), .Z(c[1865]) );
  XNOR U14292 ( .A(a[1865]), .B(n12060), .Z(n12059) );
  IV U14293 ( .A(n12057), .Z(n12060) );
  XOR U14294 ( .A(n12061), .B(n12062), .Z(n12057) );
  ANDN U14295 ( .B(n12063), .A(n12064), .Z(n12061) );
  XNOR U14296 ( .A(b[1864]), .B(n12062), .Z(n12063) );
  XNOR U14297 ( .A(b[1864]), .B(n12064), .Z(c[1864]) );
  XNOR U14298 ( .A(a[1864]), .B(n12065), .Z(n12064) );
  IV U14299 ( .A(n12062), .Z(n12065) );
  XOR U14300 ( .A(n12066), .B(n12067), .Z(n12062) );
  ANDN U14301 ( .B(n12068), .A(n12069), .Z(n12066) );
  XNOR U14302 ( .A(b[1863]), .B(n12067), .Z(n12068) );
  XNOR U14303 ( .A(b[1863]), .B(n12069), .Z(c[1863]) );
  XNOR U14304 ( .A(a[1863]), .B(n12070), .Z(n12069) );
  IV U14305 ( .A(n12067), .Z(n12070) );
  XOR U14306 ( .A(n12071), .B(n12072), .Z(n12067) );
  ANDN U14307 ( .B(n12073), .A(n12074), .Z(n12071) );
  XNOR U14308 ( .A(b[1862]), .B(n12072), .Z(n12073) );
  XNOR U14309 ( .A(b[1862]), .B(n12074), .Z(c[1862]) );
  XNOR U14310 ( .A(a[1862]), .B(n12075), .Z(n12074) );
  IV U14311 ( .A(n12072), .Z(n12075) );
  XOR U14312 ( .A(n12076), .B(n12077), .Z(n12072) );
  ANDN U14313 ( .B(n12078), .A(n12079), .Z(n12076) );
  XNOR U14314 ( .A(b[1861]), .B(n12077), .Z(n12078) );
  XNOR U14315 ( .A(b[1861]), .B(n12079), .Z(c[1861]) );
  XNOR U14316 ( .A(a[1861]), .B(n12080), .Z(n12079) );
  IV U14317 ( .A(n12077), .Z(n12080) );
  XOR U14318 ( .A(n12081), .B(n12082), .Z(n12077) );
  ANDN U14319 ( .B(n12083), .A(n12084), .Z(n12081) );
  XNOR U14320 ( .A(b[1860]), .B(n12082), .Z(n12083) );
  XNOR U14321 ( .A(b[1860]), .B(n12084), .Z(c[1860]) );
  XNOR U14322 ( .A(a[1860]), .B(n12085), .Z(n12084) );
  IV U14323 ( .A(n12082), .Z(n12085) );
  XOR U14324 ( .A(n12086), .B(n12087), .Z(n12082) );
  ANDN U14325 ( .B(n12088), .A(n12089), .Z(n12086) );
  XNOR U14326 ( .A(b[1859]), .B(n12087), .Z(n12088) );
  XNOR U14327 ( .A(b[185]), .B(n12090), .Z(c[185]) );
  XNOR U14328 ( .A(b[1859]), .B(n12089), .Z(c[1859]) );
  XNOR U14329 ( .A(a[1859]), .B(n12091), .Z(n12089) );
  IV U14330 ( .A(n12087), .Z(n12091) );
  XOR U14331 ( .A(n12092), .B(n12093), .Z(n12087) );
  ANDN U14332 ( .B(n12094), .A(n12095), .Z(n12092) );
  XNOR U14333 ( .A(b[1858]), .B(n12093), .Z(n12094) );
  XNOR U14334 ( .A(b[1858]), .B(n12095), .Z(c[1858]) );
  XNOR U14335 ( .A(a[1858]), .B(n12096), .Z(n12095) );
  IV U14336 ( .A(n12093), .Z(n12096) );
  XOR U14337 ( .A(n12097), .B(n12098), .Z(n12093) );
  ANDN U14338 ( .B(n12099), .A(n12100), .Z(n12097) );
  XNOR U14339 ( .A(b[1857]), .B(n12098), .Z(n12099) );
  XNOR U14340 ( .A(b[1857]), .B(n12100), .Z(c[1857]) );
  XNOR U14341 ( .A(a[1857]), .B(n12101), .Z(n12100) );
  IV U14342 ( .A(n12098), .Z(n12101) );
  XOR U14343 ( .A(n12102), .B(n12103), .Z(n12098) );
  ANDN U14344 ( .B(n12104), .A(n12105), .Z(n12102) );
  XNOR U14345 ( .A(b[1856]), .B(n12103), .Z(n12104) );
  XNOR U14346 ( .A(b[1856]), .B(n12105), .Z(c[1856]) );
  XNOR U14347 ( .A(a[1856]), .B(n12106), .Z(n12105) );
  IV U14348 ( .A(n12103), .Z(n12106) );
  XOR U14349 ( .A(n12107), .B(n12108), .Z(n12103) );
  ANDN U14350 ( .B(n12109), .A(n12110), .Z(n12107) );
  XNOR U14351 ( .A(b[1855]), .B(n12108), .Z(n12109) );
  XNOR U14352 ( .A(b[1855]), .B(n12110), .Z(c[1855]) );
  XNOR U14353 ( .A(a[1855]), .B(n12111), .Z(n12110) );
  IV U14354 ( .A(n12108), .Z(n12111) );
  XOR U14355 ( .A(n12112), .B(n12113), .Z(n12108) );
  ANDN U14356 ( .B(n12114), .A(n12115), .Z(n12112) );
  XNOR U14357 ( .A(b[1854]), .B(n12113), .Z(n12114) );
  XNOR U14358 ( .A(b[1854]), .B(n12115), .Z(c[1854]) );
  XNOR U14359 ( .A(a[1854]), .B(n12116), .Z(n12115) );
  IV U14360 ( .A(n12113), .Z(n12116) );
  XOR U14361 ( .A(n12117), .B(n12118), .Z(n12113) );
  ANDN U14362 ( .B(n12119), .A(n12120), .Z(n12117) );
  XNOR U14363 ( .A(b[1853]), .B(n12118), .Z(n12119) );
  XNOR U14364 ( .A(b[1853]), .B(n12120), .Z(c[1853]) );
  XNOR U14365 ( .A(a[1853]), .B(n12121), .Z(n12120) );
  IV U14366 ( .A(n12118), .Z(n12121) );
  XOR U14367 ( .A(n12122), .B(n12123), .Z(n12118) );
  ANDN U14368 ( .B(n12124), .A(n12125), .Z(n12122) );
  XNOR U14369 ( .A(b[1852]), .B(n12123), .Z(n12124) );
  XNOR U14370 ( .A(b[1852]), .B(n12125), .Z(c[1852]) );
  XNOR U14371 ( .A(a[1852]), .B(n12126), .Z(n12125) );
  IV U14372 ( .A(n12123), .Z(n12126) );
  XOR U14373 ( .A(n12127), .B(n12128), .Z(n12123) );
  ANDN U14374 ( .B(n12129), .A(n12130), .Z(n12127) );
  XNOR U14375 ( .A(b[1851]), .B(n12128), .Z(n12129) );
  XNOR U14376 ( .A(b[1851]), .B(n12130), .Z(c[1851]) );
  XNOR U14377 ( .A(a[1851]), .B(n12131), .Z(n12130) );
  IV U14378 ( .A(n12128), .Z(n12131) );
  XOR U14379 ( .A(n12132), .B(n12133), .Z(n12128) );
  ANDN U14380 ( .B(n12134), .A(n12135), .Z(n12132) );
  XNOR U14381 ( .A(b[1850]), .B(n12133), .Z(n12134) );
  XNOR U14382 ( .A(b[1850]), .B(n12135), .Z(c[1850]) );
  XNOR U14383 ( .A(a[1850]), .B(n12136), .Z(n12135) );
  IV U14384 ( .A(n12133), .Z(n12136) );
  XOR U14385 ( .A(n12137), .B(n12138), .Z(n12133) );
  ANDN U14386 ( .B(n12139), .A(n12140), .Z(n12137) );
  XNOR U14387 ( .A(b[1849]), .B(n12138), .Z(n12139) );
  XNOR U14388 ( .A(b[184]), .B(n12141), .Z(c[184]) );
  XNOR U14389 ( .A(b[1849]), .B(n12140), .Z(c[1849]) );
  XNOR U14390 ( .A(a[1849]), .B(n12142), .Z(n12140) );
  IV U14391 ( .A(n12138), .Z(n12142) );
  XOR U14392 ( .A(n12143), .B(n12144), .Z(n12138) );
  ANDN U14393 ( .B(n12145), .A(n12146), .Z(n12143) );
  XNOR U14394 ( .A(b[1848]), .B(n12144), .Z(n12145) );
  XNOR U14395 ( .A(b[1848]), .B(n12146), .Z(c[1848]) );
  XNOR U14396 ( .A(a[1848]), .B(n12147), .Z(n12146) );
  IV U14397 ( .A(n12144), .Z(n12147) );
  XOR U14398 ( .A(n12148), .B(n12149), .Z(n12144) );
  ANDN U14399 ( .B(n12150), .A(n12151), .Z(n12148) );
  XNOR U14400 ( .A(b[1847]), .B(n12149), .Z(n12150) );
  XNOR U14401 ( .A(b[1847]), .B(n12151), .Z(c[1847]) );
  XNOR U14402 ( .A(a[1847]), .B(n12152), .Z(n12151) );
  IV U14403 ( .A(n12149), .Z(n12152) );
  XOR U14404 ( .A(n12153), .B(n12154), .Z(n12149) );
  ANDN U14405 ( .B(n12155), .A(n12156), .Z(n12153) );
  XNOR U14406 ( .A(b[1846]), .B(n12154), .Z(n12155) );
  XNOR U14407 ( .A(b[1846]), .B(n12156), .Z(c[1846]) );
  XNOR U14408 ( .A(a[1846]), .B(n12157), .Z(n12156) );
  IV U14409 ( .A(n12154), .Z(n12157) );
  XOR U14410 ( .A(n12158), .B(n12159), .Z(n12154) );
  ANDN U14411 ( .B(n12160), .A(n12161), .Z(n12158) );
  XNOR U14412 ( .A(b[1845]), .B(n12159), .Z(n12160) );
  XNOR U14413 ( .A(b[1845]), .B(n12161), .Z(c[1845]) );
  XNOR U14414 ( .A(a[1845]), .B(n12162), .Z(n12161) );
  IV U14415 ( .A(n12159), .Z(n12162) );
  XOR U14416 ( .A(n12163), .B(n12164), .Z(n12159) );
  ANDN U14417 ( .B(n12165), .A(n12166), .Z(n12163) );
  XNOR U14418 ( .A(b[1844]), .B(n12164), .Z(n12165) );
  XNOR U14419 ( .A(b[1844]), .B(n12166), .Z(c[1844]) );
  XNOR U14420 ( .A(a[1844]), .B(n12167), .Z(n12166) );
  IV U14421 ( .A(n12164), .Z(n12167) );
  XOR U14422 ( .A(n12168), .B(n12169), .Z(n12164) );
  ANDN U14423 ( .B(n12170), .A(n12171), .Z(n12168) );
  XNOR U14424 ( .A(b[1843]), .B(n12169), .Z(n12170) );
  XNOR U14425 ( .A(b[1843]), .B(n12171), .Z(c[1843]) );
  XNOR U14426 ( .A(a[1843]), .B(n12172), .Z(n12171) );
  IV U14427 ( .A(n12169), .Z(n12172) );
  XOR U14428 ( .A(n12173), .B(n12174), .Z(n12169) );
  ANDN U14429 ( .B(n12175), .A(n12176), .Z(n12173) );
  XNOR U14430 ( .A(b[1842]), .B(n12174), .Z(n12175) );
  XNOR U14431 ( .A(b[1842]), .B(n12176), .Z(c[1842]) );
  XNOR U14432 ( .A(a[1842]), .B(n12177), .Z(n12176) );
  IV U14433 ( .A(n12174), .Z(n12177) );
  XOR U14434 ( .A(n12178), .B(n12179), .Z(n12174) );
  ANDN U14435 ( .B(n12180), .A(n12181), .Z(n12178) );
  XNOR U14436 ( .A(b[1841]), .B(n12179), .Z(n12180) );
  XNOR U14437 ( .A(b[1841]), .B(n12181), .Z(c[1841]) );
  XNOR U14438 ( .A(a[1841]), .B(n12182), .Z(n12181) );
  IV U14439 ( .A(n12179), .Z(n12182) );
  XOR U14440 ( .A(n12183), .B(n12184), .Z(n12179) );
  ANDN U14441 ( .B(n12185), .A(n12186), .Z(n12183) );
  XNOR U14442 ( .A(b[1840]), .B(n12184), .Z(n12185) );
  XNOR U14443 ( .A(b[1840]), .B(n12186), .Z(c[1840]) );
  XNOR U14444 ( .A(a[1840]), .B(n12187), .Z(n12186) );
  IV U14445 ( .A(n12184), .Z(n12187) );
  XOR U14446 ( .A(n12188), .B(n12189), .Z(n12184) );
  ANDN U14447 ( .B(n12190), .A(n12191), .Z(n12188) );
  XNOR U14448 ( .A(b[1839]), .B(n12189), .Z(n12190) );
  XNOR U14449 ( .A(b[183]), .B(n12192), .Z(c[183]) );
  XNOR U14450 ( .A(b[1839]), .B(n12191), .Z(c[1839]) );
  XNOR U14451 ( .A(a[1839]), .B(n12193), .Z(n12191) );
  IV U14452 ( .A(n12189), .Z(n12193) );
  XOR U14453 ( .A(n12194), .B(n12195), .Z(n12189) );
  ANDN U14454 ( .B(n12196), .A(n12197), .Z(n12194) );
  XNOR U14455 ( .A(b[1838]), .B(n12195), .Z(n12196) );
  XNOR U14456 ( .A(b[1838]), .B(n12197), .Z(c[1838]) );
  XNOR U14457 ( .A(a[1838]), .B(n12198), .Z(n12197) );
  IV U14458 ( .A(n12195), .Z(n12198) );
  XOR U14459 ( .A(n12199), .B(n12200), .Z(n12195) );
  ANDN U14460 ( .B(n12201), .A(n12202), .Z(n12199) );
  XNOR U14461 ( .A(b[1837]), .B(n12200), .Z(n12201) );
  XNOR U14462 ( .A(b[1837]), .B(n12202), .Z(c[1837]) );
  XNOR U14463 ( .A(a[1837]), .B(n12203), .Z(n12202) );
  IV U14464 ( .A(n12200), .Z(n12203) );
  XOR U14465 ( .A(n12204), .B(n12205), .Z(n12200) );
  ANDN U14466 ( .B(n12206), .A(n12207), .Z(n12204) );
  XNOR U14467 ( .A(b[1836]), .B(n12205), .Z(n12206) );
  XNOR U14468 ( .A(b[1836]), .B(n12207), .Z(c[1836]) );
  XNOR U14469 ( .A(a[1836]), .B(n12208), .Z(n12207) );
  IV U14470 ( .A(n12205), .Z(n12208) );
  XOR U14471 ( .A(n12209), .B(n12210), .Z(n12205) );
  ANDN U14472 ( .B(n12211), .A(n12212), .Z(n12209) );
  XNOR U14473 ( .A(b[1835]), .B(n12210), .Z(n12211) );
  XNOR U14474 ( .A(b[1835]), .B(n12212), .Z(c[1835]) );
  XNOR U14475 ( .A(a[1835]), .B(n12213), .Z(n12212) );
  IV U14476 ( .A(n12210), .Z(n12213) );
  XOR U14477 ( .A(n12214), .B(n12215), .Z(n12210) );
  ANDN U14478 ( .B(n12216), .A(n12217), .Z(n12214) );
  XNOR U14479 ( .A(b[1834]), .B(n12215), .Z(n12216) );
  XNOR U14480 ( .A(b[1834]), .B(n12217), .Z(c[1834]) );
  XNOR U14481 ( .A(a[1834]), .B(n12218), .Z(n12217) );
  IV U14482 ( .A(n12215), .Z(n12218) );
  XOR U14483 ( .A(n12219), .B(n12220), .Z(n12215) );
  ANDN U14484 ( .B(n12221), .A(n12222), .Z(n12219) );
  XNOR U14485 ( .A(b[1833]), .B(n12220), .Z(n12221) );
  XNOR U14486 ( .A(b[1833]), .B(n12222), .Z(c[1833]) );
  XNOR U14487 ( .A(a[1833]), .B(n12223), .Z(n12222) );
  IV U14488 ( .A(n12220), .Z(n12223) );
  XOR U14489 ( .A(n12224), .B(n12225), .Z(n12220) );
  ANDN U14490 ( .B(n12226), .A(n12227), .Z(n12224) );
  XNOR U14491 ( .A(b[1832]), .B(n12225), .Z(n12226) );
  XNOR U14492 ( .A(b[1832]), .B(n12227), .Z(c[1832]) );
  XNOR U14493 ( .A(a[1832]), .B(n12228), .Z(n12227) );
  IV U14494 ( .A(n12225), .Z(n12228) );
  XOR U14495 ( .A(n12229), .B(n12230), .Z(n12225) );
  ANDN U14496 ( .B(n12231), .A(n12232), .Z(n12229) );
  XNOR U14497 ( .A(b[1831]), .B(n12230), .Z(n12231) );
  XNOR U14498 ( .A(b[1831]), .B(n12232), .Z(c[1831]) );
  XNOR U14499 ( .A(a[1831]), .B(n12233), .Z(n12232) );
  IV U14500 ( .A(n12230), .Z(n12233) );
  XOR U14501 ( .A(n12234), .B(n12235), .Z(n12230) );
  ANDN U14502 ( .B(n12236), .A(n12237), .Z(n12234) );
  XNOR U14503 ( .A(b[1830]), .B(n12235), .Z(n12236) );
  XNOR U14504 ( .A(b[1830]), .B(n12237), .Z(c[1830]) );
  XNOR U14505 ( .A(a[1830]), .B(n12238), .Z(n12237) );
  IV U14506 ( .A(n12235), .Z(n12238) );
  XOR U14507 ( .A(n12239), .B(n12240), .Z(n12235) );
  ANDN U14508 ( .B(n12241), .A(n12242), .Z(n12239) );
  XNOR U14509 ( .A(b[1829]), .B(n12240), .Z(n12241) );
  XNOR U14510 ( .A(b[182]), .B(n12243), .Z(c[182]) );
  XNOR U14511 ( .A(b[1829]), .B(n12242), .Z(c[1829]) );
  XNOR U14512 ( .A(a[1829]), .B(n12244), .Z(n12242) );
  IV U14513 ( .A(n12240), .Z(n12244) );
  XOR U14514 ( .A(n12245), .B(n12246), .Z(n12240) );
  ANDN U14515 ( .B(n12247), .A(n12248), .Z(n12245) );
  XNOR U14516 ( .A(b[1828]), .B(n12246), .Z(n12247) );
  XNOR U14517 ( .A(b[1828]), .B(n12248), .Z(c[1828]) );
  XNOR U14518 ( .A(a[1828]), .B(n12249), .Z(n12248) );
  IV U14519 ( .A(n12246), .Z(n12249) );
  XOR U14520 ( .A(n12250), .B(n12251), .Z(n12246) );
  ANDN U14521 ( .B(n12252), .A(n12253), .Z(n12250) );
  XNOR U14522 ( .A(b[1827]), .B(n12251), .Z(n12252) );
  XNOR U14523 ( .A(b[1827]), .B(n12253), .Z(c[1827]) );
  XNOR U14524 ( .A(a[1827]), .B(n12254), .Z(n12253) );
  IV U14525 ( .A(n12251), .Z(n12254) );
  XOR U14526 ( .A(n12255), .B(n12256), .Z(n12251) );
  ANDN U14527 ( .B(n12257), .A(n12258), .Z(n12255) );
  XNOR U14528 ( .A(b[1826]), .B(n12256), .Z(n12257) );
  XNOR U14529 ( .A(b[1826]), .B(n12258), .Z(c[1826]) );
  XNOR U14530 ( .A(a[1826]), .B(n12259), .Z(n12258) );
  IV U14531 ( .A(n12256), .Z(n12259) );
  XOR U14532 ( .A(n12260), .B(n12261), .Z(n12256) );
  ANDN U14533 ( .B(n12262), .A(n12263), .Z(n12260) );
  XNOR U14534 ( .A(b[1825]), .B(n12261), .Z(n12262) );
  XNOR U14535 ( .A(b[1825]), .B(n12263), .Z(c[1825]) );
  XNOR U14536 ( .A(a[1825]), .B(n12264), .Z(n12263) );
  IV U14537 ( .A(n12261), .Z(n12264) );
  XOR U14538 ( .A(n12265), .B(n12266), .Z(n12261) );
  ANDN U14539 ( .B(n12267), .A(n12268), .Z(n12265) );
  XNOR U14540 ( .A(b[1824]), .B(n12266), .Z(n12267) );
  XNOR U14541 ( .A(b[1824]), .B(n12268), .Z(c[1824]) );
  XNOR U14542 ( .A(a[1824]), .B(n12269), .Z(n12268) );
  IV U14543 ( .A(n12266), .Z(n12269) );
  XOR U14544 ( .A(n12270), .B(n12271), .Z(n12266) );
  ANDN U14545 ( .B(n12272), .A(n12273), .Z(n12270) );
  XNOR U14546 ( .A(b[1823]), .B(n12271), .Z(n12272) );
  XNOR U14547 ( .A(b[1823]), .B(n12273), .Z(c[1823]) );
  XNOR U14548 ( .A(a[1823]), .B(n12274), .Z(n12273) );
  IV U14549 ( .A(n12271), .Z(n12274) );
  XOR U14550 ( .A(n12275), .B(n12276), .Z(n12271) );
  ANDN U14551 ( .B(n12277), .A(n12278), .Z(n12275) );
  XNOR U14552 ( .A(b[1822]), .B(n12276), .Z(n12277) );
  XNOR U14553 ( .A(b[1822]), .B(n12278), .Z(c[1822]) );
  XNOR U14554 ( .A(a[1822]), .B(n12279), .Z(n12278) );
  IV U14555 ( .A(n12276), .Z(n12279) );
  XOR U14556 ( .A(n12280), .B(n12281), .Z(n12276) );
  ANDN U14557 ( .B(n12282), .A(n12283), .Z(n12280) );
  XNOR U14558 ( .A(b[1821]), .B(n12281), .Z(n12282) );
  XNOR U14559 ( .A(b[1821]), .B(n12283), .Z(c[1821]) );
  XNOR U14560 ( .A(a[1821]), .B(n12284), .Z(n12283) );
  IV U14561 ( .A(n12281), .Z(n12284) );
  XOR U14562 ( .A(n12285), .B(n12286), .Z(n12281) );
  ANDN U14563 ( .B(n12287), .A(n12288), .Z(n12285) );
  XNOR U14564 ( .A(b[1820]), .B(n12286), .Z(n12287) );
  XNOR U14565 ( .A(b[1820]), .B(n12288), .Z(c[1820]) );
  XNOR U14566 ( .A(a[1820]), .B(n12289), .Z(n12288) );
  IV U14567 ( .A(n12286), .Z(n12289) );
  XOR U14568 ( .A(n12290), .B(n12291), .Z(n12286) );
  ANDN U14569 ( .B(n12292), .A(n12293), .Z(n12290) );
  XNOR U14570 ( .A(b[1819]), .B(n12291), .Z(n12292) );
  XNOR U14571 ( .A(b[181]), .B(n12294), .Z(c[181]) );
  XNOR U14572 ( .A(b[1819]), .B(n12293), .Z(c[1819]) );
  XNOR U14573 ( .A(a[1819]), .B(n12295), .Z(n12293) );
  IV U14574 ( .A(n12291), .Z(n12295) );
  XOR U14575 ( .A(n12296), .B(n12297), .Z(n12291) );
  ANDN U14576 ( .B(n12298), .A(n12299), .Z(n12296) );
  XNOR U14577 ( .A(b[1818]), .B(n12297), .Z(n12298) );
  XNOR U14578 ( .A(b[1818]), .B(n12299), .Z(c[1818]) );
  XNOR U14579 ( .A(a[1818]), .B(n12300), .Z(n12299) );
  IV U14580 ( .A(n12297), .Z(n12300) );
  XOR U14581 ( .A(n12301), .B(n12302), .Z(n12297) );
  ANDN U14582 ( .B(n12303), .A(n12304), .Z(n12301) );
  XNOR U14583 ( .A(b[1817]), .B(n12302), .Z(n12303) );
  XNOR U14584 ( .A(b[1817]), .B(n12304), .Z(c[1817]) );
  XNOR U14585 ( .A(a[1817]), .B(n12305), .Z(n12304) );
  IV U14586 ( .A(n12302), .Z(n12305) );
  XOR U14587 ( .A(n12306), .B(n12307), .Z(n12302) );
  ANDN U14588 ( .B(n12308), .A(n12309), .Z(n12306) );
  XNOR U14589 ( .A(b[1816]), .B(n12307), .Z(n12308) );
  XNOR U14590 ( .A(b[1816]), .B(n12309), .Z(c[1816]) );
  XNOR U14591 ( .A(a[1816]), .B(n12310), .Z(n12309) );
  IV U14592 ( .A(n12307), .Z(n12310) );
  XOR U14593 ( .A(n12311), .B(n12312), .Z(n12307) );
  ANDN U14594 ( .B(n12313), .A(n12314), .Z(n12311) );
  XNOR U14595 ( .A(b[1815]), .B(n12312), .Z(n12313) );
  XNOR U14596 ( .A(b[1815]), .B(n12314), .Z(c[1815]) );
  XNOR U14597 ( .A(a[1815]), .B(n12315), .Z(n12314) );
  IV U14598 ( .A(n12312), .Z(n12315) );
  XOR U14599 ( .A(n12316), .B(n12317), .Z(n12312) );
  ANDN U14600 ( .B(n12318), .A(n12319), .Z(n12316) );
  XNOR U14601 ( .A(b[1814]), .B(n12317), .Z(n12318) );
  XNOR U14602 ( .A(b[1814]), .B(n12319), .Z(c[1814]) );
  XNOR U14603 ( .A(a[1814]), .B(n12320), .Z(n12319) );
  IV U14604 ( .A(n12317), .Z(n12320) );
  XOR U14605 ( .A(n12321), .B(n12322), .Z(n12317) );
  ANDN U14606 ( .B(n12323), .A(n12324), .Z(n12321) );
  XNOR U14607 ( .A(b[1813]), .B(n12322), .Z(n12323) );
  XNOR U14608 ( .A(b[1813]), .B(n12324), .Z(c[1813]) );
  XNOR U14609 ( .A(a[1813]), .B(n12325), .Z(n12324) );
  IV U14610 ( .A(n12322), .Z(n12325) );
  XOR U14611 ( .A(n12326), .B(n12327), .Z(n12322) );
  ANDN U14612 ( .B(n12328), .A(n12329), .Z(n12326) );
  XNOR U14613 ( .A(b[1812]), .B(n12327), .Z(n12328) );
  XNOR U14614 ( .A(b[1812]), .B(n12329), .Z(c[1812]) );
  XNOR U14615 ( .A(a[1812]), .B(n12330), .Z(n12329) );
  IV U14616 ( .A(n12327), .Z(n12330) );
  XOR U14617 ( .A(n12331), .B(n12332), .Z(n12327) );
  ANDN U14618 ( .B(n12333), .A(n12334), .Z(n12331) );
  XNOR U14619 ( .A(b[1811]), .B(n12332), .Z(n12333) );
  XNOR U14620 ( .A(b[1811]), .B(n12334), .Z(c[1811]) );
  XNOR U14621 ( .A(a[1811]), .B(n12335), .Z(n12334) );
  IV U14622 ( .A(n12332), .Z(n12335) );
  XOR U14623 ( .A(n12336), .B(n12337), .Z(n12332) );
  ANDN U14624 ( .B(n12338), .A(n12339), .Z(n12336) );
  XNOR U14625 ( .A(b[1810]), .B(n12337), .Z(n12338) );
  XNOR U14626 ( .A(b[1810]), .B(n12339), .Z(c[1810]) );
  XNOR U14627 ( .A(a[1810]), .B(n12340), .Z(n12339) );
  IV U14628 ( .A(n12337), .Z(n12340) );
  XOR U14629 ( .A(n12341), .B(n12342), .Z(n12337) );
  ANDN U14630 ( .B(n12343), .A(n12344), .Z(n12341) );
  XNOR U14631 ( .A(b[1809]), .B(n12342), .Z(n12343) );
  XNOR U14632 ( .A(b[180]), .B(n12345), .Z(c[180]) );
  XNOR U14633 ( .A(b[1809]), .B(n12344), .Z(c[1809]) );
  XNOR U14634 ( .A(a[1809]), .B(n12346), .Z(n12344) );
  IV U14635 ( .A(n12342), .Z(n12346) );
  XOR U14636 ( .A(n12347), .B(n12348), .Z(n12342) );
  ANDN U14637 ( .B(n12349), .A(n12350), .Z(n12347) );
  XNOR U14638 ( .A(b[1808]), .B(n12348), .Z(n12349) );
  XNOR U14639 ( .A(b[1808]), .B(n12350), .Z(c[1808]) );
  XNOR U14640 ( .A(a[1808]), .B(n12351), .Z(n12350) );
  IV U14641 ( .A(n12348), .Z(n12351) );
  XOR U14642 ( .A(n12352), .B(n12353), .Z(n12348) );
  ANDN U14643 ( .B(n12354), .A(n12355), .Z(n12352) );
  XNOR U14644 ( .A(b[1807]), .B(n12353), .Z(n12354) );
  XNOR U14645 ( .A(b[1807]), .B(n12355), .Z(c[1807]) );
  XNOR U14646 ( .A(a[1807]), .B(n12356), .Z(n12355) );
  IV U14647 ( .A(n12353), .Z(n12356) );
  XOR U14648 ( .A(n12357), .B(n12358), .Z(n12353) );
  ANDN U14649 ( .B(n12359), .A(n12360), .Z(n12357) );
  XNOR U14650 ( .A(b[1806]), .B(n12358), .Z(n12359) );
  XNOR U14651 ( .A(b[1806]), .B(n12360), .Z(c[1806]) );
  XNOR U14652 ( .A(a[1806]), .B(n12361), .Z(n12360) );
  IV U14653 ( .A(n12358), .Z(n12361) );
  XOR U14654 ( .A(n12362), .B(n12363), .Z(n12358) );
  ANDN U14655 ( .B(n12364), .A(n12365), .Z(n12362) );
  XNOR U14656 ( .A(b[1805]), .B(n12363), .Z(n12364) );
  XNOR U14657 ( .A(b[1805]), .B(n12365), .Z(c[1805]) );
  XNOR U14658 ( .A(a[1805]), .B(n12366), .Z(n12365) );
  IV U14659 ( .A(n12363), .Z(n12366) );
  XOR U14660 ( .A(n12367), .B(n12368), .Z(n12363) );
  ANDN U14661 ( .B(n12369), .A(n12370), .Z(n12367) );
  XNOR U14662 ( .A(b[1804]), .B(n12368), .Z(n12369) );
  XNOR U14663 ( .A(b[1804]), .B(n12370), .Z(c[1804]) );
  XNOR U14664 ( .A(a[1804]), .B(n12371), .Z(n12370) );
  IV U14665 ( .A(n12368), .Z(n12371) );
  XOR U14666 ( .A(n12372), .B(n12373), .Z(n12368) );
  ANDN U14667 ( .B(n12374), .A(n12375), .Z(n12372) );
  XNOR U14668 ( .A(b[1803]), .B(n12373), .Z(n12374) );
  XNOR U14669 ( .A(b[1803]), .B(n12375), .Z(c[1803]) );
  XNOR U14670 ( .A(a[1803]), .B(n12376), .Z(n12375) );
  IV U14671 ( .A(n12373), .Z(n12376) );
  XOR U14672 ( .A(n12377), .B(n12378), .Z(n12373) );
  ANDN U14673 ( .B(n12379), .A(n12380), .Z(n12377) );
  XNOR U14674 ( .A(b[1802]), .B(n12378), .Z(n12379) );
  XNOR U14675 ( .A(b[1802]), .B(n12380), .Z(c[1802]) );
  XNOR U14676 ( .A(a[1802]), .B(n12381), .Z(n12380) );
  IV U14677 ( .A(n12378), .Z(n12381) );
  XOR U14678 ( .A(n12382), .B(n12383), .Z(n12378) );
  ANDN U14679 ( .B(n12384), .A(n12385), .Z(n12382) );
  XNOR U14680 ( .A(b[1801]), .B(n12383), .Z(n12384) );
  XNOR U14681 ( .A(b[1801]), .B(n12385), .Z(c[1801]) );
  XNOR U14682 ( .A(a[1801]), .B(n12386), .Z(n12385) );
  IV U14683 ( .A(n12383), .Z(n12386) );
  XOR U14684 ( .A(n12387), .B(n12388), .Z(n12383) );
  ANDN U14685 ( .B(n12389), .A(n12390), .Z(n12387) );
  XNOR U14686 ( .A(b[1800]), .B(n12388), .Z(n12389) );
  XNOR U14687 ( .A(b[1800]), .B(n12390), .Z(c[1800]) );
  XNOR U14688 ( .A(a[1800]), .B(n12391), .Z(n12390) );
  IV U14689 ( .A(n12388), .Z(n12391) );
  XOR U14690 ( .A(n12392), .B(n12393), .Z(n12388) );
  ANDN U14691 ( .B(n12394), .A(n12395), .Z(n12392) );
  XNOR U14692 ( .A(b[1799]), .B(n12393), .Z(n12394) );
  XNOR U14693 ( .A(b[17]), .B(n12396), .Z(c[17]) );
  XNOR U14694 ( .A(b[179]), .B(n12397), .Z(c[179]) );
  XNOR U14695 ( .A(b[1799]), .B(n12395), .Z(c[1799]) );
  XNOR U14696 ( .A(a[1799]), .B(n12398), .Z(n12395) );
  IV U14697 ( .A(n12393), .Z(n12398) );
  XOR U14698 ( .A(n12399), .B(n12400), .Z(n12393) );
  ANDN U14699 ( .B(n12401), .A(n12402), .Z(n12399) );
  XNOR U14700 ( .A(b[1798]), .B(n12400), .Z(n12401) );
  XNOR U14701 ( .A(b[1798]), .B(n12402), .Z(c[1798]) );
  XNOR U14702 ( .A(a[1798]), .B(n12403), .Z(n12402) );
  IV U14703 ( .A(n12400), .Z(n12403) );
  XOR U14704 ( .A(n12404), .B(n12405), .Z(n12400) );
  ANDN U14705 ( .B(n12406), .A(n12407), .Z(n12404) );
  XNOR U14706 ( .A(b[1797]), .B(n12405), .Z(n12406) );
  XNOR U14707 ( .A(b[1797]), .B(n12407), .Z(c[1797]) );
  XNOR U14708 ( .A(a[1797]), .B(n12408), .Z(n12407) );
  IV U14709 ( .A(n12405), .Z(n12408) );
  XOR U14710 ( .A(n12409), .B(n12410), .Z(n12405) );
  ANDN U14711 ( .B(n12411), .A(n12412), .Z(n12409) );
  XNOR U14712 ( .A(b[1796]), .B(n12410), .Z(n12411) );
  XNOR U14713 ( .A(b[1796]), .B(n12412), .Z(c[1796]) );
  XNOR U14714 ( .A(a[1796]), .B(n12413), .Z(n12412) );
  IV U14715 ( .A(n12410), .Z(n12413) );
  XOR U14716 ( .A(n12414), .B(n12415), .Z(n12410) );
  ANDN U14717 ( .B(n12416), .A(n12417), .Z(n12414) );
  XNOR U14718 ( .A(b[1795]), .B(n12415), .Z(n12416) );
  XNOR U14719 ( .A(b[1795]), .B(n12417), .Z(c[1795]) );
  XNOR U14720 ( .A(a[1795]), .B(n12418), .Z(n12417) );
  IV U14721 ( .A(n12415), .Z(n12418) );
  XOR U14722 ( .A(n12419), .B(n12420), .Z(n12415) );
  ANDN U14723 ( .B(n12421), .A(n12422), .Z(n12419) );
  XNOR U14724 ( .A(b[1794]), .B(n12420), .Z(n12421) );
  XNOR U14725 ( .A(b[1794]), .B(n12422), .Z(c[1794]) );
  XNOR U14726 ( .A(a[1794]), .B(n12423), .Z(n12422) );
  IV U14727 ( .A(n12420), .Z(n12423) );
  XOR U14728 ( .A(n12424), .B(n12425), .Z(n12420) );
  ANDN U14729 ( .B(n12426), .A(n12427), .Z(n12424) );
  XNOR U14730 ( .A(b[1793]), .B(n12425), .Z(n12426) );
  XNOR U14731 ( .A(b[1793]), .B(n12427), .Z(c[1793]) );
  XNOR U14732 ( .A(a[1793]), .B(n12428), .Z(n12427) );
  IV U14733 ( .A(n12425), .Z(n12428) );
  XOR U14734 ( .A(n12429), .B(n12430), .Z(n12425) );
  ANDN U14735 ( .B(n12431), .A(n12432), .Z(n12429) );
  XNOR U14736 ( .A(b[1792]), .B(n12430), .Z(n12431) );
  XNOR U14737 ( .A(b[1792]), .B(n12432), .Z(c[1792]) );
  XNOR U14738 ( .A(a[1792]), .B(n12433), .Z(n12432) );
  IV U14739 ( .A(n12430), .Z(n12433) );
  XOR U14740 ( .A(n12434), .B(n12435), .Z(n12430) );
  ANDN U14741 ( .B(n12436), .A(n12437), .Z(n12434) );
  XNOR U14742 ( .A(b[1791]), .B(n12435), .Z(n12436) );
  XNOR U14743 ( .A(b[1791]), .B(n12437), .Z(c[1791]) );
  XNOR U14744 ( .A(a[1791]), .B(n12438), .Z(n12437) );
  IV U14745 ( .A(n12435), .Z(n12438) );
  XOR U14746 ( .A(n12439), .B(n12440), .Z(n12435) );
  ANDN U14747 ( .B(n12441), .A(n12442), .Z(n12439) );
  XNOR U14748 ( .A(b[1790]), .B(n12440), .Z(n12441) );
  XNOR U14749 ( .A(b[1790]), .B(n12442), .Z(c[1790]) );
  XNOR U14750 ( .A(a[1790]), .B(n12443), .Z(n12442) );
  IV U14751 ( .A(n12440), .Z(n12443) );
  XOR U14752 ( .A(n12444), .B(n12445), .Z(n12440) );
  ANDN U14753 ( .B(n12446), .A(n12447), .Z(n12444) );
  XNOR U14754 ( .A(b[1789]), .B(n12445), .Z(n12446) );
  XNOR U14755 ( .A(b[178]), .B(n12448), .Z(c[178]) );
  XNOR U14756 ( .A(b[1789]), .B(n12447), .Z(c[1789]) );
  XNOR U14757 ( .A(a[1789]), .B(n12449), .Z(n12447) );
  IV U14758 ( .A(n12445), .Z(n12449) );
  XOR U14759 ( .A(n12450), .B(n12451), .Z(n12445) );
  ANDN U14760 ( .B(n12452), .A(n12453), .Z(n12450) );
  XNOR U14761 ( .A(b[1788]), .B(n12451), .Z(n12452) );
  XNOR U14762 ( .A(b[1788]), .B(n12453), .Z(c[1788]) );
  XNOR U14763 ( .A(a[1788]), .B(n12454), .Z(n12453) );
  IV U14764 ( .A(n12451), .Z(n12454) );
  XOR U14765 ( .A(n12455), .B(n12456), .Z(n12451) );
  ANDN U14766 ( .B(n12457), .A(n12458), .Z(n12455) );
  XNOR U14767 ( .A(b[1787]), .B(n12456), .Z(n12457) );
  XNOR U14768 ( .A(b[1787]), .B(n12458), .Z(c[1787]) );
  XNOR U14769 ( .A(a[1787]), .B(n12459), .Z(n12458) );
  IV U14770 ( .A(n12456), .Z(n12459) );
  XOR U14771 ( .A(n12460), .B(n12461), .Z(n12456) );
  ANDN U14772 ( .B(n12462), .A(n12463), .Z(n12460) );
  XNOR U14773 ( .A(b[1786]), .B(n12461), .Z(n12462) );
  XNOR U14774 ( .A(b[1786]), .B(n12463), .Z(c[1786]) );
  XNOR U14775 ( .A(a[1786]), .B(n12464), .Z(n12463) );
  IV U14776 ( .A(n12461), .Z(n12464) );
  XOR U14777 ( .A(n12465), .B(n12466), .Z(n12461) );
  ANDN U14778 ( .B(n12467), .A(n12468), .Z(n12465) );
  XNOR U14779 ( .A(b[1785]), .B(n12466), .Z(n12467) );
  XNOR U14780 ( .A(b[1785]), .B(n12468), .Z(c[1785]) );
  XNOR U14781 ( .A(a[1785]), .B(n12469), .Z(n12468) );
  IV U14782 ( .A(n12466), .Z(n12469) );
  XOR U14783 ( .A(n12470), .B(n12471), .Z(n12466) );
  ANDN U14784 ( .B(n12472), .A(n12473), .Z(n12470) );
  XNOR U14785 ( .A(b[1784]), .B(n12471), .Z(n12472) );
  XNOR U14786 ( .A(b[1784]), .B(n12473), .Z(c[1784]) );
  XNOR U14787 ( .A(a[1784]), .B(n12474), .Z(n12473) );
  IV U14788 ( .A(n12471), .Z(n12474) );
  XOR U14789 ( .A(n12475), .B(n12476), .Z(n12471) );
  ANDN U14790 ( .B(n12477), .A(n12478), .Z(n12475) );
  XNOR U14791 ( .A(b[1783]), .B(n12476), .Z(n12477) );
  XNOR U14792 ( .A(b[1783]), .B(n12478), .Z(c[1783]) );
  XNOR U14793 ( .A(a[1783]), .B(n12479), .Z(n12478) );
  IV U14794 ( .A(n12476), .Z(n12479) );
  XOR U14795 ( .A(n12480), .B(n12481), .Z(n12476) );
  ANDN U14796 ( .B(n12482), .A(n12483), .Z(n12480) );
  XNOR U14797 ( .A(b[1782]), .B(n12481), .Z(n12482) );
  XNOR U14798 ( .A(b[1782]), .B(n12483), .Z(c[1782]) );
  XNOR U14799 ( .A(a[1782]), .B(n12484), .Z(n12483) );
  IV U14800 ( .A(n12481), .Z(n12484) );
  XOR U14801 ( .A(n12485), .B(n12486), .Z(n12481) );
  ANDN U14802 ( .B(n12487), .A(n12488), .Z(n12485) );
  XNOR U14803 ( .A(b[1781]), .B(n12486), .Z(n12487) );
  XNOR U14804 ( .A(b[1781]), .B(n12488), .Z(c[1781]) );
  XNOR U14805 ( .A(a[1781]), .B(n12489), .Z(n12488) );
  IV U14806 ( .A(n12486), .Z(n12489) );
  XOR U14807 ( .A(n12490), .B(n12491), .Z(n12486) );
  ANDN U14808 ( .B(n12492), .A(n12493), .Z(n12490) );
  XNOR U14809 ( .A(b[1780]), .B(n12491), .Z(n12492) );
  XNOR U14810 ( .A(b[1780]), .B(n12493), .Z(c[1780]) );
  XNOR U14811 ( .A(a[1780]), .B(n12494), .Z(n12493) );
  IV U14812 ( .A(n12491), .Z(n12494) );
  XOR U14813 ( .A(n12495), .B(n12496), .Z(n12491) );
  ANDN U14814 ( .B(n12497), .A(n12498), .Z(n12495) );
  XNOR U14815 ( .A(b[1779]), .B(n12496), .Z(n12497) );
  XNOR U14816 ( .A(b[177]), .B(n12499), .Z(c[177]) );
  XNOR U14817 ( .A(b[1779]), .B(n12498), .Z(c[1779]) );
  XNOR U14818 ( .A(a[1779]), .B(n12500), .Z(n12498) );
  IV U14819 ( .A(n12496), .Z(n12500) );
  XOR U14820 ( .A(n12501), .B(n12502), .Z(n12496) );
  ANDN U14821 ( .B(n12503), .A(n12504), .Z(n12501) );
  XNOR U14822 ( .A(b[1778]), .B(n12502), .Z(n12503) );
  XNOR U14823 ( .A(b[1778]), .B(n12504), .Z(c[1778]) );
  XNOR U14824 ( .A(a[1778]), .B(n12505), .Z(n12504) );
  IV U14825 ( .A(n12502), .Z(n12505) );
  XOR U14826 ( .A(n12506), .B(n12507), .Z(n12502) );
  ANDN U14827 ( .B(n12508), .A(n12509), .Z(n12506) );
  XNOR U14828 ( .A(b[1777]), .B(n12507), .Z(n12508) );
  XNOR U14829 ( .A(b[1777]), .B(n12509), .Z(c[1777]) );
  XNOR U14830 ( .A(a[1777]), .B(n12510), .Z(n12509) );
  IV U14831 ( .A(n12507), .Z(n12510) );
  XOR U14832 ( .A(n12511), .B(n12512), .Z(n12507) );
  ANDN U14833 ( .B(n12513), .A(n12514), .Z(n12511) );
  XNOR U14834 ( .A(b[1776]), .B(n12512), .Z(n12513) );
  XNOR U14835 ( .A(b[1776]), .B(n12514), .Z(c[1776]) );
  XNOR U14836 ( .A(a[1776]), .B(n12515), .Z(n12514) );
  IV U14837 ( .A(n12512), .Z(n12515) );
  XOR U14838 ( .A(n12516), .B(n12517), .Z(n12512) );
  ANDN U14839 ( .B(n12518), .A(n12519), .Z(n12516) );
  XNOR U14840 ( .A(b[1775]), .B(n12517), .Z(n12518) );
  XNOR U14841 ( .A(b[1775]), .B(n12519), .Z(c[1775]) );
  XNOR U14842 ( .A(a[1775]), .B(n12520), .Z(n12519) );
  IV U14843 ( .A(n12517), .Z(n12520) );
  XOR U14844 ( .A(n12521), .B(n12522), .Z(n12517) );
  ANDN U14845 ( .B(n12523), .A(n12524), .Z(n12521) );
  XNOR U14846 ( .A(b[1774]), .B(n12522), .Z(n12523) );
  XNOR U14847 ( .A(b[1774]), .B(n12524), .Z(c[1774]) );
  XNOR U14848 ( .A(a[1774]), .B(n12525), .Z(n12524) );
  IV U14849 ( .A(n12522), .Z(n12525) );
  XOR U14850 ( .A(n12526), .B(n12527), .Z(n12522) );
  ANDN U14851 ( .B(n12528), .A(n12529), .Z(n12526) );
  XNOR U14852 ( .A(b[1773]), .B(n12527), .Z(n12528) );
  XNOR U14853 ( .A(b[1773]), .B(n12529), .Z(c[1773]) );
  XNOR U14854 ( .A(a[1773]), .B(n12530), .Z(n12529) );
  IV U14855 ( .A(n12527), .Z(n12530) );
  XOR U14856 ( .A(n12531), .B(n12532), .Z(n12527) );
  ANDN U14857 ( .B(n12533), .A(n12534), .Z(n12531) );
  XNOR U14858 ( .A(b[1772]), .B(n12532), .Z(n12533) );
  XNOR U14859 ( .A(b[1772]), .B(n12534), .Z(c[1772]) );
  XNOR U14860 ( .A(a[1772]), .B(n12535), .Z(n12534) );
  IV U14861 ( .A(n12532), .Z(n12535) );
  XOR U14862 ( .A(n12536), .B(n12537), .Z(n12532) );
  ANDN U14863 ( .B(n12538), .A(n12539), .Z(n12536) );
  XNOR U14864 ( .A(b[1771]), .B(n12537), .Z(n12538) );
  XNOR U14865 ( .A(b[1771]), .B(n12539), .Z(c[1771]) );
  XNOR U14866 ( .A(a[1771]), .B(n12540), .Z(n12539) );
  IV U14867 ( .A(n12537), .Z(n12540) );
  XOR U14868 ( .A(n12541), .B(n12542), .Z(n12537) );
  ANDN U14869 ( .B(n12543), .A(n12544), .Z(n12541) );
  XNOR U14870 ( .A(b[1770]), .B(n12542), .Z(n12543) );
  XNOR U14871 ( .A(b[1770]), .B(n12544), .Z(c[1770]) );
  XNOR U14872 ( .A(a[1770]), .B(n12545), .Z(n12544) );
  IV U14873 ( .A(n12542), .Z(n12545) );
  XOR U14874 ( .A(n12546), .B(n12547), .Z(n12542) );
  ANDN U14875 ( .B(n12548), .A(n12549), .Z(n12546) );
  XNOR U14876 ( .A(b[1769]), .B(n12547), .Z(n12548) );
  XNOR U14877 ( .A(b[176]), .B(n12550), .Z(c[176]) );
  XNOR U14878 ( .A(b[1769]), .B(n12549), .Z(c[1769]) );
  XNOR U14879 ( .A(a[1769]), .B(n12551), .Z(n12549) );
  IV U14880 ( .A(n12547), .Z(n12551) );
  XOR U14881 ( .A(n12552), .B(n12553), .Z(n12547) );
  ANDN U14882 ( .B(n12554), .A(n12555), .Z(n12552) );
  XNOR U14883 ( .A(b[1768]), .B(n12553), .Z(n12554) );
  XNOR U14884 ( .A(b[1768]), .B(n12555), .Z(c[1768]) );
  XNOR U14885 ( .A(a[1768]), .B(n12556), .Z(n12555) );
  IV U14886 ( .A(n12553), .Z(n12556) );
  XOR U14887 ( .A(n12557), .B(n12558), .Z(n12553) );
  ANDN U14888 ( .B(n12559), .A(n12560), .Z(n12557) );
  XNOR U14889 ( .A(b[1767]), .B(n12558), .Z(n12559) );
  XNOR U14890 ( .A(b[1767]), .B(n12560), .Z(c[1767]) );
  XNOR U14891 ( .A(a[1767]), .B(n12561), .Z(n12560) );
  IV U14892 ( .A(n12558), .Z(n12561) );
  XOR U14893 ( .A(n12562), .B(n12563), .Z(n12558) );
  ANDN U14894 ( .B(n12564), .A(n12565), .Z(n12562) );
  XNOR U14895 ( .A(b[1766]), .B(n12563), .Z(n12564) );
  XNOR U14896 ( .A(b[1766]), .B(n12565), .Z(c[1766]) );
  XNOR U14897 ( .A(a[1766]), .B(n12566), .Z(n12565) );
  IV U14898 ( .A(n12563), .Z(n12566) );
  XOR U14899 ( .A(n12567), .B(n12568), .Z(n12563) );
  ANDN U14900 ( .B(n12569), .A(n12570), .Z(n12567) );
  XNOR U14901 ( .A(b[1765]), .B(n12568), .Z(n12569) );
  XNOR U14902 ( .A(b[1765]), .B(n12570), .Z(c[1765]) );
  XNOR U14903 ( .A(a[1765]), .B(n12571), .Z(n12570) );
  IV U14904 ( .A(n12568), .Z(n12571) );
  XOR U14905 ( .A(n12572), .B(n12573), .Z(n12568) );
  ANDN U14906 ( .B(n12574), .A(n12575), .Z(n12572) );
  XNOR U14907 ( .A(b[1764]), .B(n12573), .Z(n12574) );
  XNOR U14908 ( .A(b[1764]), .B(n12575), .Z(c[1764]) );
  XNOR U14909 ( .A(a[1764]), .B(n12576), .Z(n12575) );
  IV U14910 ( .A(n12573), .Z(n12576) );
  XOR U14911 ( .A(n12577), .B(n12578), .Z(n12573) );
  ANDN U14912 ( .B(n12579), .A(n12580), .Z(n12577) );
  XNOR U14913 ( .A(b[1763]), .B(n12578), .Z(n12579) );
  XNOR U14914 ( .A(b[1763]), .B(n12580), .Z(c[1763]) );
  XNOR U14915 ( .A(a[1763]), .B(n12581), .Z(n12580) );
  IV U14916 ( .A(n12578), .Z(n12581) );
  XOR U14917 ( .A(n12582), .B(n12583), .Z(n12578) );
  ANDN U14918 ( .B(n12584), .A(n12585), .Z(n12582) );
  XNOR U14919 ( .A(b[1762]), .B(n12583), .Z(n12584) );
  XNOR U14920 ( .A(b[1762]), .B(n12585), .Z(c[1762]) );
  XNOR U14921 ( .A(a[1762]), .B(n12586), .Z(n12585) );
  IV U14922 ( .A(n12583), .Z(n12586) );
  XOR U14923 ( .A(n12587), .B(n12588), .Z(n12583) );
  ANDN U14924 ( .B(n12589), .A(n12590), .Z(n12587) );
  XNOR U14925 ( .A(b[1761]), .B(n12588), .Z(n12589) );
  XNOR U14926 ( .A(b[1761]), .B(n12590), .Z(c[1761]) );
  XNOR U14927 ( .A(a[1761]), .B(n12591), .Z(n12590) );
  IV U14928 ( .A(n12588), .Z(n12591) );
  XOR U14929 ( .A(n12592), .B(n12593), .Z(n12588) );
  ANDN U14930 ( .B(n12594), .A(n12595), .Z(n12592) );
  XNOR U14931 ( .A(b[1760]), .B(n12593), .Z(n12594) );
  XNOR U14932 ( .A(b[1760]), .B(n12595), .Z(c[1760]) );
  XNOR U14933 ( .A(a[1760]), .B(n12596), .Z(n12595) );
  IV U14934 ( .A(n12593), .Z(n12596) );
  XOR U14935 ( .A(n12597), .B(n12598), .Z(n12593) );
  ANDN U14936 ( .B(n12599), .A(n12600), .Z(n12597) );
  XNOR U14937 ( .A(b[1759]), .B(n12598), .Z(n12599) );
  XNOR U14938 ( .A(b[175]), .B(n12601), .Z(c[175]) );
  XNOR U14939 ( .A(b[1759]), .B(n12600), .Z(c[1759]) );
  XNOR U14940 ( .A(a[1759]), .B(n12602), .Z(n12600) );
  IV U14941 ( .A(n12598), .Z(n12602) );
  XOR U14942 ( .A(n12603), .B(n12604), .Z(n12598) );
  ANDN U14943 ( .B(n12605), .A(n12606), .Z(n12603) );
  XNOR U14944 ( .A(b[1758]), .B(n12604), .Z(n12605) );
  XNOR U14945 ( .A(b[1758]), .B(n12606), .Z(c[1758]) );
  XNOR U14946 ( .A(a[1758]), .B(n12607), .Z(n12606) );
  IV U14947 ( .A(n12604), .Z(n12607) );
  XOR U14948 ( .A(n12608), .B(n12609), .Z(n12604) );
  ANDN U14949 ( .B(n12610), .A(n12611), .Z(n12608) );
  XNOR U14950 ( .A(b[1757]), .B(n12609), .Z(n12610) );
  XNOR U14951 ( .A(b[1757]), .B(n12611), .Z(c[1757]) );
  XNOR U14952 ( .A(a[1757]), .B(n12612), .Z(n12611) );
  IV U14953 ( .A(n12609), .Z(n12612) );
  XOR U14954 ( .A(n12613), .B(n12614), .Z(n12609) );
  ANDN U14955 ( .B(n12615), .A(n12616), .Z(n12613) );
  XNOR U14956 ( .A(b[1756]), .B(n12614), .Z(n12615) );
  XNOR U14957 ( .A(b[1756]), .B(n12616), .Z(c[1756]) );
  XNOR U14958 ( .A(a[1756]), .B(n12617), .Z(n12616) );
  IV U14959 ( .A(n12614), .Z(n12617) );
  XOR U14960 ( .A(n12618), .B(n12619), .Z(n12614) );
  ANDN U14961 ( .B(n12620), .A(n12621), .Z(n12618) );
  XNOR U14962 ( .A(b[1755]), .B(n12619), .Z(n12620) );
  XNOR U14963 ( .A(b[1755]), .B(n12621), .Z(c[1755]) );
  XNOR U14964 ( .A(a[1755]), .B(n12622), .Z(n12621) );
  IV U14965 ( .A(n12619), .Z(n12622) );
  XOR U14966 ( .A(n12623), .B(n12624), .Z(n12619) );
  ANDN U14967 ( .B(n12625), .A(n12626), .Z(n12623) );
  XNOR U14968 ( .A(b[1754]), .B(n12624), .Z(n12625) );
  XNOR U14969 ( .A(b[1754]), .B(n12626), .Z(c[1754]) );
  XNOR U14970 ( .A(a[1754]), .B(n12627), .Z(n12626) );
  IV U14971 ( .A(n12624), .Z(n12627) );
  XOR U14972 ( .A(n12628), .B(n12629), .Z(n12624) );
  ANDN U14973 ( .B(n12630), .A(n12631), .Z(n12628) );
  XNOR U14974 ( .A(b[1753]), .B(n12629), .Z(n12630) );
  XNOR U14975 ( .A(b[1753]), .B(n12631), .Z(c[1753]) );
  XNOR U14976 ( .A(a[1753]), .B(n12632), .Z(n12631) );
  IV U14977 ( .A(n12629), .Z(n12632) );
  XOR U14978 ( .A(n12633), .B(n12634), .Z(n12629) );
  ANDN U14979 ( .B(n12635), .A(n12636), .Z(n12633) );
  XNOR U14980 ( .A(b[1752]), .B(n12634), .Z(n12635) );
  XNOR U14981 ( .A(b[1752]), .B(n12636), .Z(c[1752]) );
  XNOR U14982 ( .A(a[1752]), .B(n12637), .Z(n12636) );
  IV U14983 ( .A(n12634), .Z(n12637) );
  XOR U14984 ( .A(n12638), .B(n12639), .Z(n12634) );
  ANDN U14985 ( .B(n12640), .A(n12641), .Z(n12638) );
  XNOR U14986 ( .A(b[1751]), .B(n12639), .Z(n12640) );
  XNOR U14987 ( .A(b[1751]), .B(n12641), .Z(c[1751]) );
  XNOR U14988 ( .A(a[1751]), .B(n12642), .Z(n12641) );
  IV U14989 ( .A(n12639), .Z(n12642) );
  XOR U14990 ( .A(n12643), .B(n12644), .Z(n12639) );
  ANDN U14991 ( .B(n12645), .A(n12646), .Z(n12643) );
  XNOR U14992 ( .A(b[1750]), .B(n12644), .Z(n12645) );
  XNOR U14993 ( .A(b[1750]), .B(n12646), .Z(c[1750]) );
  XNOR U14994 ( .A(a[1750]), .B(n12647), .Z(n12646) );
  IV U14995 ( .A(n12644), .Z(n12647) );
  XOR U14996 ( .A(n12648), .B(n12649), .Z(n12644) );
  ANDN U14997 ( .B(n12650), .A(n12651), .Z(n12648) );
  XNOR U14998 ( .A(b[1749]), .B(n12649), .Z(n12650) );
  XNOR U14999 ( .A(b[174]), .B(n12652), .Z(c[174]) );
  XNOR U15000 ( .A(b[1749]), .B(n12651), .Z(c[1749]) );
  XNOR U15001 ( .A(a[1749]), .B(n12653), .Z(n12651) );
  IV U15002 ( .A(n12649), .Z(n12653) );
  XOR U15003 ( .A(n12654), .B(n12655), .Z(n12649) );
  ANDN U15004 ( .B(n12656), .A(n12657), .Z(n12654) );
  XNOR U15005 ( .A(b[1748]), .B(n12655), .Z(n12656) );
  XNOR U15006 ( .A(b[1748]), .B(n12657), .Z(c[1748]) );
  XNOR U15007 ( .A(a[1748]), .B(n12658), .Z(n12657) );
  IV U15008 ( .A(n12655), .Z(n12658) );
  XOR U15009 ( .A(n12659), .B(n12660), .Z(n12655) );
  ANDN U15010 ( .B(n12661), .A(n12662), .Z(n12659) );
  XNOR U15011 ( .A(b[1747]), .B(n12660), .Z(n12661) );
  XNOR U15012 ( .A(b[1747]), .B(n12662), .Z(c[1747]) );
  XNOR U15013 ( .A(a[1747]), .B(n12663), .Z(n12662) );
  IV U15014 ( .A(n12660), .Z(n12663) );
  XOR U15015 ( .A(n12664), .B(n12665), .Z(n12660) );
  ANDN U15016 ( .B(n12666), .A(n12667), .Z(n12664) );
  XNOR U15017 ( .A(b[1746]), .B(n12665), .Z(n12666) );
  XNOR U15018 ( .A(b[1746]), .B(n12667), .Z(c[1746]) );
  XNOR U15019 ( .A(a[1746]), .B(n12668), .Z(n12667) );
  IV U15020 ( .A(n12665), .Z(n12668) );
  XOR U15021 ( .A(n12669), .B(n12670), .Z(n12665) );
  ANDN U15022 ( .B(n12671), .A(n12672), .Z(n12669) );
  XNOR U15023 ( .A(b[1745]), .B(n12670), .Z(n12671) );
  XNOR U15024 ( .A(b[1745]), .B(n12672), .Z(c[1745]) );
  XNOR U15025 ( .A(a[1745]), .B(n12673), .Z(n12672) );
  IV U15026 ( .A(n12670), .Z(n12673) );
  XOR U15027 ( .A(n12674), .B(n12675), .Z(n12670) );
  ANDN U15028 ( .B(n12676), .A(n12677), .Z(n12674) );
  XNOR U15029 ( .A(b[1744]), .B(n12675), .Z(n12676) );
  XNOR U15030 ( .A(b[1744]), .B(n12677), .Z(c[1744]) );
  XNOR U15031 ( .A(a[1744]), .B(n12678), .Z(n12677) );
  IV U15032 ( .A(n12675), .Z(n12678) );
  XOR U15033 ( .A(n12679), .B(n12680), .Z(n12675) );
  ANDN U15034 ( .B(n12681), .A(n12682), .Z(n12679) );
  XNOR U15035 ( .A(b[1743]), .B(n12680), .Z(n12681) );
  XNOR U15036 ( .A(b[1743]), .B(n12682), .Z(c[1743]) );
  XNOR U15037 ( .A(a[1743]), .B(n12683), .Z(n12682) );
  IV U15038 ( .A(n12680), .Z(n12683) );
  XOR U15039 ( .A(n12684), .B(n12685), .Z(n12680) );
  ANDN U15040 ( .B(n12686), .A(n12687), .Z(n12684) );
  XNOR U15041 ( .A(b[1742]), .B(n12685), .Z(n12686) );
  XNOR U15042 ( .A(b[1742]), .B(n12687), .Z(c[1742]) );
  XNOR U15043 ( .A(a[1742]), .B(n12688), .Z(n12687) );
  IV U15044 ( .A(n12685), .Z(n12688) );
  XOR U15045 ( .A(n12689), .B(n12690), .Z(n12685) );
  ANDN U15046 ( .B(n12691), .A(n12692), .Z(n12689) );
  XNOR U15047 ( .A(b[1741]), .B(n12690), .Z(n12691) );
  XNOR U15048 ( .A(b[1741]), .B(n12692), .Z(c[1741]) );
  XNOR U15049 ( .A(a[1741]), .B(n12693), .Z(n12692) );
  IV U15050 ( .A(n12690), .Z(n12693) );
  XOR U15051 ( .A(n12694), .B(n12695), .Z(n12690) );
  ANDN U15052 ( .B(n12696), .A(n12697), .Z(n12694) );
  XNOR U15053 ( .A(b[1740]), .B(n12695), .Z(n12696) );
  XNOR U15054 ( .A(b[1740]), .B(n12697), .Z(c[1740]) );
  XNOR U15055 ( .A(a[1740]), .B(n12698), .Z(n12697) );
  IV U15056 ( .A(n12695), .Z(n12698) );
  XOR U15057 ( .A(n12699), .B(n12700), .Z(n12695) );
  ANDN U15058 ( .B(n12701), .A(n12702), .Z(n12699) );
  XNOR U15059 ( .A(b[1739]), .B(n12700), .Z(n12701) );
  XNOR U15060 ( .A(b[173]), .B(n12703), .Z(c[173]) );
  XNOR U15061 ( .A(b[1739]), .B(n12702), .Z(c[1739]) );
  XNOR U15062 ( .A(a[1739]), .B(n12704), .Z(n12702) );
  IV U15063 ( .A(n12700), .Z(n12704) );
  XOR U15064 ( .A(n12705), .B(n12706), .Z(n12700) );
  ANDN U15065 ( .B(n12707), .A(n12708), .Z(n12705) );
  XNOR U15066 ( .A(b[1738]), .B(n12706), .Z(n12707) );
  XNOR U15067 ( .A(b[1738]), .B(n12708), .Z(c[1738]) );
  XNOR U15068 ( .A(a[1738]), .B(n12709), .Z(n12708) );
  IV U15069 ( .A(n12706), .Z(n12709) );
  XOR U15070 ( .A(n12710), .B(n12711), .Z(n12706) );
  ANDN U15071 ( .B(n12712), .A(n12713), .Z(n12710) );
  XNOR U15072 ( .A(b[1737]), .B(n12711), .Z(n12712) );
  XNOR U15073 ( .A(b[1737]), .B(n12713), .Z(c[1737]) );
  XNOR U15074 ( .A(a[1737]), .B(n12714), .Z(n12713) );
  IV U15075 ( .A(n12711), .Z(n12714) );
  XOR U15076 ( .A(n12715), .B(n12716), .Z(n12711) );
  ANDN U15077 ( .B(n12717), .A(n12718), .Z(n12715) );
  XNOR U15078 ( .A(b[1736]), .B(n12716), .Z(n12717) );
  XNOR U15079 ( .A(b[1736]), .B(n12718), .Z(c[1736]) );
  XNOR U15080 ( .A(a[1736]), .B(n12719), .Z(n12718) );
  IV U15081 ( .A(n12716), .Z(n12719) );
  XOR U15082 ( .A(n12720), .B(n12721), .Z(n12716) );
  ANDN U15083 ( .B(n12722), .A(n12723), .Z(n12720) );
  XNOR U15084 ( .A(b[1735]), .B(n12721), .Z(n12722) );
  XNOR U15085 ( .A(b[1735]), .B(n12723), .Z(c[1735]) );
  XNOR U15086 ( .A(a[1735]), .B(n12724), .Z(n12723) );
  IV U15087 ( .A(n12721), .Z(n12724) );
  XOR U15088 ( .A(n12725), .B(n12726), .Z(n12721) );
  ANDN U15089 ( .B(n12727), .A(n12728), .Z(n12725) );
  XNOR U15090 ( .A(b[1734]), .B(n12726), .Z(n12727) );
  XNOR U15091 ( .A(b[1734]), .B(n12728), .Z(c[1734]) );
  XNOR U15092 ( .A(a[1734]), .B(n12729), .Z(n12728) );
  IV U15093 ( .A(n12726), .Z(n12729) );
  XOR U15094 ( .A(n12730), .B(n12731), .Z(n12726) );
  ANDN U15095 ( .B(n12732), .A(n12733), .Z(n12730) );
  XNOR U15096 ( .A(b[1733]), .B(n12731), .Z(n12732) );
  XNOR U15097 ( .A(b[1733]), .B(n12733), .Z(c[1733]) );
  XNOR U15098 ( .A(a[1733]), .B(n12734), .Z(n12733) );
  IV U15099 ( .A(n12731), .Z(n12734) );
  XOR U15100 ( .A(n12735), .B(n12736), .Z(n12731) );
  ANDN U15101 ( .B(n12737), .A(n12738), .Z(n12735) );
  XNOR U15102 ( .A(b[1732]), .B(n12736), .Z(n12737) );
  XNOR U15103 ( .A(b[1732]), .B(n12738), .Z(c[1732]) );
  XNOR U15104 ( .A(a[1732]), .B(n12739), .Z(n12738) );
  IV U15105 ( .A(n12736), .Z(n12739) );
  XOR U15106 ( .A(n12740), .B(n12741), .Z(n12736) );
  ANDN U15107 ( .B(n12742), .A(n12743), .Z(n12740) );
  XNOR U15108 ( .A(b[1731]), .B(n12741), .Z(n12742) );
  XNOR U15109 ( .A(b[1731]), .B(n12743), .Z(c[1731]) );
  XNOR U15110 ( .A(a[1731]), .B(n12744), .Z(n12743) );
  IV U15111 ( .A(n12741), .Z(n12744) );
  XOR U15112 ( .A(n12745), .B(n12746), .Z(n12741) );
  ANDN U15113 ( .B(n12747), .A(n12748), .Z(n12745) );
  XNOR U15114 ( .A(b[1730]), .B(n12746), .Z(n12747) );
  XNOR U15115 ( .A(b[1730]), .B(n12748), .Z(c[1730]) );
  XNOR U15116 ( .A(a[1730]), .B(n12749), .Z(n12748) );
  IV U15117 ( .A(n12746), .Z(n12749) );
  XOR U15118 ( .A(n12750), .B(n12751), .Z(n12746) );
  ANDN U15119 ( .B(n12752), .A(n12753), .Z(n12750) );
  XNOR U15120 ( .A(b[1729]), .B(n12751), .Z(n12752) );
  XNOR U15121 ( .A(b[172]), .B(n12754), .Z(c[172]) );
  XNOR U15122 ( .A(b[1729]), .B(n12753), .Z(c[1729]) );
  XNOR U15123 ( .A(a[1729]), .B(n12755), .Z(n12753) );
  IV U15124 ( .A(n12751), .Z(n12755) );
  XOR U15125 ( .A(n12756), .B(n12757), .Z(n12751) );
  ANDN U15126 ( .B(n12758), .A(n12759), .Z(n12756) );
  XNOR U15127 ( .A(b[1728]), .B(n12757), .Z(n12758) );
  XNOR U15128 ( .A(b[1728]), .B(n12759), .Z(c[1728]) );
  XNOR U15129 ( .A(a[1728]), .B(n12760), .Z(n12759) );
  IV U15130 ( .A(n12757), .Z(n12760) );
  XOR U15131 ( .A(n12761), .B(n12762), .Z(n12757) );
  ANDN U15132 ( .B(n12763), .A(n12764), .Z(n12761) );
  XNOR U15133 ( .A(b[1727]), .B(n12762), .Z(n12763) );
  XNOR U15134 ( .A(b[1727]), .B(n12764), .Z(c[1727]) );
  XNOR U15135 ( .A(a[1727]), .B(n12765), .Z(n12764) );
  IV U15136 ( .A(n12762), .Z(n12765) );
  XOR U15137 ( .A(n12766), .B(n12767), .Z(n12762) );
  ANDN U15138 ( .B(n12768), .A(n12769), .Z(n12766) );
  XNOR U15139 ( .A(b[1726]), .B(n12767), .Z(n12768) );
  XNOR U15140 ( .A(b[1726]), .B(n12769), .Z(c[1726]) );
  XNOR U15141 ( .A(a[1726]), .B(n12770), .Z(n12769) );
  IV U15142 ( .A(n12767), .Z(n12770) );
  XOR U15143 ( .A(n12771), .B(n12772), .Z(n12767) );
  ANDN U15144 ( .B(n12773), .A(n12774), .Z(n12771) );
  XNOR U15145 ( .A(b[1725]), .B(n12772), .Z(n12773) );
  XNOR U15146 ( .A(b[1725]), .B(n12774), .Z(c[1725]) );
  XNOR U15147 ( .A(a[1725]), .B(n12775), .Z(n12774) );
  IV U15148 ( .A(n12772), .Z(n12775) );
  XOR U15149 ( .A(n12776), .B(n12777), .Z(n12772) );
  ANDN U15150 ( .B(n12778), .A(n12779), .Z(n12776) );
  XNOR U15151 ( .A(b[1724]), .B(n12777), .Z(n12778) );
  XNOR U15152 ( .A(b[1724]), .B(n12779), .Z(c[1724]) );
  XNOR U15153 ( .A(a[1724]), .B(n12780), .Z(n12779) );
  IV U15154 ( .A(n12777), .Z(n12780) );
  XOR U15155 ( .A(n12781), .B(n12782), .Z(n12777) );
  ANDN U15156 ( .B(n12783), .A(n12784), .Z(n12781) );
  XNOR U15157 ( .A(b[1723]), .B(n12782), .Z(n12783) );
  XNOR U15158 ( .A(b[1723]), .B(n12784), .Z(c[1723]) );
  XNOR U15159 ( .A(a[1723]), .B(n12785), .Z(n12784) );
  IV U15160 ( .A(n12782), .Z(n12785) );
  XOR U15161 ( .A(n12786), .B(n12787), .Z(n12782) );
  ANDN U15162 ( .B(n12788), .A(n12789), .Z(n12786) );
  XNOR U15163 ( .A(b[1722]), .B(n12787), .Z(n12788) );
  XNOR U15164 ( .A(b[1722]), .B(n12789), .Z(c[1722]) );
  XNOR U15165 ( .A(a[1722]), .B(n12790), .Z(n12789) );
  IV U15166 ( .A(n12787), .Z(n12790) );
  XOR U15167 ( .A(n12791), .B(n12792), .Z(n12787) );
  ANDN U15168 ( .B(n12793), .A(n12794), .Z(n12791) );
  XNOR U15169 ( .A(b[1721]), .B(n12792), .Z(n12793) );
  XNOR U15170 ( .A(b[1721]), .B(n12794), .Z(c[1721]) );
  XNOR U15171 ( .A(a[1721]), .B(n12795), .Z(n12794) );
  IV U15172 ( .A(n12792), .Z(n12795) );
  XOR U15173 ( .A(n12796), .B(n12797), .Z(n12792) );
  ANDN U15174 ( .B(n12798), .A(n12799), .Z(n12796) );
  XNOR U15175 ( .A(b[1720]), .B(n12797), .Z(n12798) );
  XNOR U15176 ( .A(b[1720]), .B(n12799), .Z(c[1720]) );
  XNOR U15177 ( .A(a[1720]), .B(n12800), .Z(n12799) );
  IV U15178 ( .A(n12797), .Z(n12800) );
  XOR U15179 ( .A(n12801), .B(n12802), .Z(n12797) );
  ANDN U15180 ( .B(n12803), .A(n12804), .Z(n12801) );
  XNOR U15181 ( .A(b[1719]), .B(n12802), .Z(n12803) );
  XNOR U15182 ( .A(b[171]), .B(n12805), .Z(c[171]) );
  XNOR U15183 ( .A(b[1719]), .B(n12804), .Z(c[1719]) );
  XNOR U15184 ( .A(a[1719]), .B(n12806), .Z(n12804) );
  IV U15185 ( .A(n12802), .Z(n12806) );
  XOR U15186 ( .A(n12807), .B(n12808), .Z(n12802) );
  ANDN U15187 ( .B(n12809), .A(n12810), .Z(n12807) );
  XNOR U15188 ( .A(b[1718]), .B(n12808), .Z(n12809) );
  XNOR U15189 ( .A(b[1718]), .B(n12810), .Z(c[1718]) );
  XNOR U15190 ( .A(a[1718]), .B(n12811), .Z(n12810) );
  IV U15191 ( .A(n12808), .Z(n12811) );
  XOR U15192 ( .A(n12812), .B(n12813), .Z(n12808) );
  ANDN U15193 ( .B(n12814), .A(n12815), .Z(n12812) );
  XNOR U15194 ( .A(b[1717]), .B(n12813), .Z(n12814) );
  XNOR U15195 ( .A(b[1717]), .B(n12815), .Z(c[1717]) );
  XNOR U15196 ( .A(a[1717]), .B(n12816), .Z(n12815) );
  IV U15197 ( .A(n12813), .Z(n12816) );
  XOR U15198 ( .A(n12817), .B(n12818), .Z(n12813) );
  ANDN U15199 ( .B(n12819), .A(n12820), .Z(n12817) );
  XNOR U15200 ( .A(b[1716]), .B(n12818), .Z(n12819) );
  XNOR U15201 ( .A(b[1716]), .B(n12820), .Z(c[1716]) );
  XNOR U15202 ( .A(a[1716]), .B(n12821), .Z(n12820) );
  IV U15203 ( .A(n12818), .Z(n12821) );
  XOR U15204 ( .A(n12822), .B(n12823), .Z(n12818) );
  ANDN U15205 ( .B(n12824), .A(n12825), .Z(n12822) );
  XNOR U15206 ( .A(b[1715]), .B(n12823), .Z(n12824) );
  XNOR U15207 ( .A(b[1715]), .B(n12825), .Z(c[1715]) );
  XNOR U15208 ( .A(a[1715]), .B(n12826), .Z(n12825) );
  IV U15209 ( .A(n12823), .Z(n12826) );
  XOR U15210 ( .A(n12827), .B(n12828), .Z(n12823) );
  ANDN U15211 ( .B(n12829), .A(n12830), .Z(n12827) );
  XNOR U15212 ( .A(b[1714]), .B(n12828), .Z(n12829) );
  XNOR U15213 ( .A(b[1714]), .B(n12830), .Z(c[1714]) );
  XNOR U15214 ( .A(a[1714]), .B(n12831), .Z(n12830) );
  IV U15215 ( .A(n12828), .Z(n12831) );
  XOR U15216 ( .A(n12832), .B(n12833), .Z(n12828) );
  ANDN U15217 ( .B(n12834), .A(n12835), .Z(n12832) );
  XNOR U15218 ( .A(b[1713]), .B(n12833), .Z(n12834) );
  XNOR U15219 ( .A(b[1713]), .B(n12835), .Z(c[1713]) );
  XNOR U15220 ( .A(a[1713]), .B(n12836), .Z(n12835) );
  IV U15221 ( .A(n12833), .Z(n12836) );
  XOR U15222 ( .A(n12837), .B(n12838), .Z(n12833) );
  ANDN U15223 ( .B(n12839), .A(n12840), .Z(n12837) );
  XNOR U15224 ( .A(b[1712]), .B(n12838), .Z(n12839) );
  XNOR U15225 ( .A(b[1712]), .B(n12840), .Z(c[1712]) );
  XNOR U15226 ( .A(a[1712]), .B(n12841), .Z(n12840) );
  IV U15227 ( .A(n12838), .Z(n12841) );
  XOR U15228 ( .A(n12842), .B(n12843), .Z(n12838) );
  ANDN U15229 ( .B(n12844), .A(n12845), .Z(n12842) );
  XNOR U15230 ( .A(b[1711]), .B(n12843), .Z(n12844) );
  XNOR U15231 ( .A(b[1711]), .B(n12845), .Z(c[1711]) );
  XNOR U15232 ( .A(a[1711]), .B(n12846), .Z(n12845) );
  IV U15233 ( .A(n12843), .Z(n12846) );
  XOR U15234 ( .A(n12847), .B(n12848), .Z(n12843) );
  ANDN U15235 ( .B(n12849), .A(n12850), .Z(n12847) );
  XNOR U15236 ( .A(b[1710]), .B(n12848), .Z(n12849) );
  XNOR U15237 ( .A(b[1710]), .B(n12850), .Z(c[1710]) );
  XNOR U15238 ( .A(a[1710]), .B(n12851), .Z(n12850) );
  IV U15239 ( .A(n12848), .Z(n12851) );
  XOR U15240 ( .A(n12852), .B(n12853), .Z(n12848) );
  ANDN U15241 ( .B(n12854), .A(n12855), .Z(n12852) );
  XNOR U15242 ( .A(b[1709]), .B(n12853), .Z(n12854) );
  XNOR U15243 ( .A(b[170]), .B(n12856), .Z(c[170]) );
  XNOR U15244 ( .A(b[1709]), .B(n12855), .Z(c[1709]) );
  XNOR U15245 ( .A(a[1709]), .B(n12857), .Z(n12855) );
  IV U15246 ( .A(n12853), .Z(n12857) );
  XOR U15247 ( .A(n12858), .B(n12859), .Z(n12853) );
  ANDN U15248 ( .B(n12860), .A(n12861), .Z(n12858) );
  XNOR U15249 ( .A(b[1708]), .B(n12859), .Z(n12860) );
  XNOR U15250 ( .A(b[1708]), .B(n12861), .Z(c[1708]) );
  XNOR U15251 ( .A(a[1708]), .B(n12862), .Z(n12861) );
  IV U15252 ( .A(n12859), .Z(n12862) );
  XOR U15253 ( .A(n12863), .B(n12864), .Z(n12859) );
  ANDN U15254 ( .B(n12865), .A(n12866), .Z(n12863) );
  XNOR U15255 ( .A(b[1707]), .B(n12864), .Z(n12865) );
  XNOR U15256 ( .A(b[1707]), .B(n12866), .Z(c[1707]) );
  XNOR U15257 ( .A(a[1707]), .B(n12867), .Z(n12866) );
  IV U15258 ( .A(n12864), .Z(n12867) );
  XOR U15259 ( .A(n12868), .B(n12869), .Z(n12864) );
  ANDN U15260 ( .B(n12870), .A(n12871), .Z(n12868) );
  XNOR U15261 ( .A(b[1706]), .B(n12869), .Z(n12870) );
  XNOR U15262 ( .A(b[1706]), .B(n12871), .Z(c[1706]) );
  XNOR U15263 ( .A(a[1706]), .B(n12872), .Z(n12871) );
  IV U15264 ( .A(n12869), .Z(n12872) );
  XOR U15265 ( .A(n12873), .B(n12874), .Z(n12869) );
  ANDN U15266 ( .B(n12875), .A(n12876), .Z(n12873) );
  XNOR U15267 ( .A(b[1705]), .B(n12874), .Z(n12875) );
  XNOR U15268 ( .A(b[1705]), .B(n12876), .Z(c[1705]) );
  XNOR U15269 ( .A(a[1705]), .B(n12877), .Z(n12876) );
  IV U15270 ( .A(n12874), .Z(n12877) );
  XOR U15271 ( .A(n12878), .B(n12879), .Z(n12874) );
  ANDN U15272 ( .B(n12880), .A(n12881), .Z(n12878) );
  XNOR U15273 ( .A(b[1704]), .B(n12879), .Z(n12880) );
  XNOR U15274 ( .A(b[1704]), .B(n12881), .Z(c[1704]) );
  XNOR U15275 ( .A(a[1704]), .B(n12882), .Z(n12881) );
  IV U15276 ( .A(n12879), .Z(n12882) );
  XOR U15277 ( .A(n12883), .B(n12884), .Z(n12879) );
  ANDN U15278 ( .B(n12885), .A(n12886), .Z(n12883) );
  XNOR U15279 ( .A(b[1703]), .B(n12884), .Z(n12885) );
  XNOR U15280 ( .A(b[1703]), .B(n12886), .Z(c[1703]) );
  XNOR U15281 ( .A(a[1703]), .B(n12887), .Z(n12886) );
  IV U15282 ( .A(n12884), .Z(n12887) );
  XOR U15283 ( .A(n12888), .B(n12889), .Z(n12884) );
  ANDN U15284 ( .B(n12890), .A(n12891), .Z(n12888) );
  XNOR U15285 ( .A(b[1702]), .B(n12889), .Z(n12890) );
  XNOR U15286 ( .A(b[1702]), .B(n12891), .Z(c[1702]) );
  XNOR U15287 ( .A(a[1702]), .B(n12892), .Z(n12891) );
  IV U15288 ( .A(n12889), .Z(n12892) );
  XOR U15289 ( .A(n12893), .B(n12894), .Z(n12889) );
  ANDN U15290 ( .B(n12895), .A(n12896), .Z(n12893) );
  XNOR U15291 ( .A(b[1701]), .B(n12894), .Z(n12895) );
  XNOR U15292 ( .A(b[1701]), .B(n12896), .Z(c[1701]) );
  XNOR U15293 ( .A(a[1701]), .B(n12897), .Z(n12896) );
  IV U15294 ( .A(n12894), .Z(n12897) );
  XOR U15295 ( .A(n12898), .B(n12899), .Z(n12894) );
  ANDN U15296 ( .B(n12900), .A(n12901), .Z(n12898) );
  XNOR U15297 ( .A(b[1700]), .B(n12899), .Z(n12900) );
  XNOR U15298 ( .A(b[1700]), .B(n12901), .Z(c[1700]) );
  XNOR U15299 ( .A(a[1700]), .B(n12902), .Z(n12901) );
  IV U15300 ( .A(n12899), .Z(n12902) );
  XOR U15301 ( .A(n12903), .B(n12904), .Z(n12899) );
  ANDN U15302 ( .B(n12905), .A(n12906), .Z(n12903) );
  XNOR U15303 ( .A(b[1699]), .B(n12904), .Z(n12905) );
  XNOR U15304 ( .A(b[16]), .B(n12907), .Z(c[16]) );
  XNOR U15305 ( .A(b[169]), .B(n12908), .Z(c[169]) );
  XNOR U15306 ( .A(b[1699]), .B(n12906), .Z(c[1699]) );
  XNOR U15307 ( .A(a[1699]), .B(n12909), .Z(n12906) );
  IV U15308 ( .A(n12904), .Z(n12909) );
  XOR U15309 ( .A(n12910), .B(n12911), .Z(n12904) );
  ANDN U15310 ( .B(n12912), .A(n12913), .Z(n12910) );
  XNOR U15311 ( .A(b[1698]), .B(n12911), .Z(n12912) );
  XNOR U15312 ( .A(b[1698]), .B(n12913), .Z(c[1698]) );
  XNOR U15313 ( .A(a[1698]), .B(n12914), .Z(n12913) );
  IV U15314 ( .A(n12911), .Z(n12914) );
  XOR U15315 ( .A(n12915), .B(n12916), .Z(n12911) );
  ANDN U15316 ( .B(n12917), .A(n12918), .Z(n12915) );
  XNOR U15317 ( .A(b[1697]), .B(n12916), .Z(n12917) );
  XNOR U15318 ( .A(b[1697]), .B(n12918), .Z(c[1697]) );
  XNOR U15319 ( .A(a[1697]), .B(n12919), .Z(n12918) );
  IV U15320 ( .A(n12916), .Z(n12919) );
  XOR U15321 ( .A(n12920), .B(n12921), .Z(n12916) );
  ANDN U15322 ( .B(n12922), .A(n12923), .Z(n12920) );
  XNOR U15323 ( .A(b[1696]), .B(n12921), .Z(n12922) );
  XNOR U15324 ( .A(b[1696]), .B(n12923), .Z(c[1696]) );
  XNOR U15325 ( .A(a[1696]), .B(n12924), .Z(n12923) );
  IV U15326 ( .A(n12921), .Z(n12924) );
  XOR U15327 ( .A(n12925), .B(n12926), .Z(n12921) );
  ANDN U15328 ( .B(n12927), .A(n12928), .Z(n12925) );
  XNOR U15329 ( .A(b[1695]), .B(n12926), .Z(n12927) );
  XNOR U15330 ( .A(b[1695]), .B(n12928), .Z(c[1695]) );
  XNOR U15331 ( .A(a[1695]), .B(n12929), .Z(n12928) );
  IV U15332 ( .A(n12926), .Z(n12929) );
  XOR U15333 ( .A(n12930), .B(n12931), .Z(n12926) );
  ANDN U15334 ( .B(n12932), .A(n12933), .Z(n12930) );
  XNOR U15335 ( .A(b[1694]), .B(n12931), .Z(n12932) );
  XNOR U15336 ( .A(b[1694]), .B(n12933), .Z(c[1694]) );
  XNOR U15337 ( .A(a[1694]), .B(n12934), .Z(n12933) );
  IV U15338 ( .A(n12931), .Z(n12934) );
  XOR U15339 ( .A(n12935), .B(n12936), .Z(n12931) );
  ANDN U15340 ( .B(n12937), .A(n12938), .Z(n12935) );
  XNOR U15341 ( .A(b[1693]), .B(n12936), .Z(n12937) );
  XNOR U15342 ( .A(b[1693]), .B(n12938), .Z(c[1693]) );
  XNOR U15343 ( .A(a[1693]), .B(n12939), .Z(n12938) );
  IV U15344 ( .A(n12936), .Z(n12939) );
  XOR U15345 ( .A(n12940), .B(n12941), .Z(n12936) );
  ANDN U15346 ( .B(n12942), .A(n12943), .Z(n12940) );
  XNOR U15347 ( .A(b[1692]), .B(n12941), .Z(n12942) );
  XNOR U15348 ( .A(b[1692]), .B(n12943), .Z(c[1692]) );
  XNOR U15349 ( .A(a[1692]), .B(n12944), .Z(n12943) );
  IV U15350 ( .A(n12941), .Z(n12944) );
  XOR U15351 ( .A(n12945), .B(n12946), .Z(n12941) );
  ANDN U15352 ( .B(n12947), .A(n12948), .Z(n12945) );
  XNOR U15353 ( .A(b[1691]), .B(n12946), .Z(n12947) );
  XNOR U15354 ( .A(b[1691]), .B(n12948), .Z(c[1691]) );
  XNOR U15355 ( .A(a[1691]), .B(n12949), .Z(n12948) );
  IV U15356 ( .A(n12946), .Z(n12949) );
  XOR U15357 ( .A(n12950), .B(n12951), .Z(n12946) );
  ANDN U15358 ( .B(n12952), .A(n12953), .Z(n12950) );
  XNOR U15359 ( .A(b[1690]), .B(n12951), .Z(n12952) );
  XNOR U15360 ( .A(b[1690]), .B(n12953), .Z(c[1690]) );
  XNOR U15361 ( .A(a[1690]), .B(n12954), .Z(n12953) );
  IV U15362 ( .A(n12951), .Z(n12954) );
  XOR U15363 ( .A(n12955), .B(n12956), .Z(n12951) );
  ANDN U15364 ( .B(n12957), .A(n12958), .Z(n12955) );
  XNOR U15365 ( .A(b[1689]), .B(n12956), .Z(n12957) );
  XNOR U15366 ( .A(b[168]), .B(n12959), .Z(c[168]) );
  XNOR U15367 ( .A(b[1689]), .B(n12958), .Z(c[1689]) );
  XNOR U15368 ( .A(a[1689]), .B(n12960), .Z(n12958) );
  IV U15369 ( .A(n12956), .Z(n12960) );
  XOR U15370 ( .A(n12961), .B(n12962), .Z(n12956) );
  ANDN U15371 ( .B(n12963), .A(n12964), .Z(n12961) );
  XNOR U15372 ( .A(b[1688]), .B(n12962), .Z(n12963) );
  XNOR U15373 ( .A(b[1688]), .B(n12964), .Z(c[1688]) );
  XNOR U15374 ( .A(a[1688]), .B(n12965), .Z(n12964) );
  IV U15375 ( .A(n12962), .Z(n12965) );
  XOR U15376 ( .A(n12966), .B(n12967), .Z(n12962) );
  ANDN U15377 ( .B(n12968), .A(n12969), .Z(n12966) );
  XNOR U15378 ( .A(b[1687]), .B(n12967), .Z(n12968) );
  XNOR U15379 ( .A(b[1687]), .B(n12969), .Z(c[1687]) );
  XNOR U15380 ( .A(a[1687]), .B(n12970), .Z(n12969) );
  IV U15381 ( .A(n12967), .Z(n12970) );
  XOR U15382 ( .A(n12971), .B(n12972), .Z(n12967) );
  ANDN U15383 ( .B(n12973), .A(n12974), .Z(n12971) );
  XNOR U15384 ( .A(b[1686]), .B(n12972), .Z(n12973) );
  XNOR U15385 ( .A(b[1686]), .B(n12974), .Z(c[1686]) );
  XNOR U15386 ( .A(a[1686]), .B(n12975), .Z(n12974) );
  IV U15387 ( .A(n12972), .Z(n12975) );
  XOR U15388 ( .A(n12976), .B(n12977), .Z(n12972) );
  ANDN U15389 ( .B(n12978), .A(n12979), .Z(n12976) );
  XNOR U15390 ( .A(b[1685]), .B(n12977), .Z(n12978) );
  XNOR U15391 ( .A(b[1685]), .B(n12979), .Z(c[1685]) );
  XNOR U15392 ( .A(a[1685]), .B(n12980), .Z(n12979) );
  IV U15393 ( .A(n12977), .Z(n12980) );
  XOR U15394 ( .A(n12981), .B(n12982), .Z(n12977) );
  ANDN U15395 ( .B(n12983), .A(n12984), .Z(n12981) );
  XNOR U15396 ( .A(b[1684]), .B(n12982), .Z(n12983) );
  XNOR U15397 ( .A(b[1684]), .B(n12984), .Z(c[1684]) );
  XNOR U15398 ( .A(a[1684]), .B(n12985), .Z(n12984) );
  IV U15399 ( .A(n12982), .Z(n12985) );
  XOR U15400 ( .A(n12986), .B(n12987), .Z(n12982) );
  ANDN U15401 ( .B(n12988), .A(n12989), .Z(n12986) );
  XNOR U15402 ( .A(b[1683]), .B(n12987), .Z(n12988) );
  XNOR U15403 ( .A(b[1683]), .B(n12989), .Z(c[1683]) );
  XNOR U15404 ( .A(a[1683]), .B(n12990), .Z(n12989) );
  IV U15405 ( .A(n12987), .Z(n12990) );
  XOR U15406 ( .A(n12991), .B(n12992), .Z(n12987) );
  ANDN U15407 ( .B(n12993), .A(n12994), .Z(n12991) );
  XNOR U15408 ( .A(b[1682]), .B(n12992), .Z(n12993) );
  XNOR U15409 ( .A(b[1682]), .B(n12994), .Z(c[1682]) );
  XNOR U15410 ( .A(a[1682]), .B(n12995), .Z(n12994) );
  IV U15411 ( .A(n12992), .Z(n12995) );
  XOR U15412 ( .A(n12996), .B(n12997), .Z(n12992) );
  ANDN U15413 ( .B(n12998), .A(n12999), .Z(n12996) );
  XNOR U15414 ( .A(b[1681]), .B(n12997), .Z(n12998) );
  XNOR U15415 ( .A(b[1681]), .B(n12999), .Z(c[1681]) );
  XNOR U15416 ( .A(a[1681]), .B(n13000), .Z(n12999) );
  IV U15417 ( .A(n12997), .Z(n13000) );
  XOR U15418 ( .A(n13001), .B(n13002), .Z(n12997) );
  ANDN U15419 ( .B(n13003), .A(n13004), .Z(n13001) );
  XNOR U15420 ( .A(b[1680]), .B(n13002), .Z(n13003) );
  XNOR U15421 ( .A(b[1680]), .B(n13004), .Z(c[1680]) );
  XNOR U15422 ( .A(a[1680]), .B(n13005), .Z(n13004) );
  IV U15423 ( .A(n13002), .Z(n13005) );
  XOR U15424 ( .A(n13006), .B(n13007), .Z(n13002) );
  ANDN U15425 ( .B(n13008), .A(n13009), .Z(n13006) );
  XNOR U15426 ( .A(b[1679]), .B(n13007), .Z(n13008) );
  XNOR U15427 ( .A(b[167]), .B(n13010), .Z(c[167]) );
  XNOR U15428 ( .A(b[1679]), .B(n13009), .Z(c[1679]) );
  XNOR U15429 ( .A(a[1679]), .B(n13011), .Z(n13009) );
  IV U15430 ( .A(n13007), .Z(n13011) );
  XOR U15431 ( .A(n13012), .B(n13013), .Z(n13007) );
  ANDN U15432 ( .B(n13014), .A(n13015), .Z(n13012) );
  XNOR U15433 ( .A(b[1678]), .B(n13013), .Z(n13014) );
  XNOR U15434 ( .A(b[1678]), .B(n13015), .Z(c[1678]) );
  XNOR U15435 ( .A(a[1678]), .B(n13016), .Z(n13015) );
  IV U15436 ( .A(n13013), .Z(n13016) );
  XOR U15437 ( .A(n13017), .B(n13018), .Z(n13013) );
  ANDN U15438 ( .B(n13019), .A(n13020), .Z(n13017) );
  XNOR U15439 ( .A(b[1677]), .B(n13018), .Z(n13019) );
  XNOR U15440 ( .A(b[1677]), .B(n13020), .Z(c[1677]) );
  XNOR U15441 ( .A(a[1677]), .B(n13021), .Z(n13020) );
  IV U15442 ( .A(n13018), .Z(n13021) );
  XOR U15443 ( .A(n13022), .B(n13023), .Z(n13018) );
  ANDN U15444 ( .B(n13024), .A(n13025), .Z(n13022) );
  XNOR U15445 ( .A(b[1676]), .B(n13023), .Z(n13024) );
  XNOR U15446 ( .A(b[1676]), .B(n13025), .Z(c[1676]) );
  XNOR U15447 ( .A(a[1676]), .B(n13026), .Z(n13025) );
  IV U15448 ( .A(n13023), .Z(n13026) );
  XOR U15449 ( .A(n13027), .B(n13028), .Z(n13023) );
  ANDN U15450 ( .B(n13029), .A(n13030), .Z(n13027) );
  XNOR U15451 ( .A(b[1675]), .B(n13028), .Z(n13029) );
  XNOR U15452 ( .A(b[1675]), .B(n13030), .Z(c[1675]) );
  XNOR U15453 ( .A(a[1675]), .B(n13031), .Z(n13030) );
  IV U15454 ( .A(n13028), .Z(n13031) );
  XOR U15455 ( .A(n13032), .B(n13033), .Z(n13028) );
  ANDN U15456 ( .B(n13034), .A(n13035), .Z(n13032) );
  XNOR U15457 ( .A(b[1674]), .B(n13033), .Z(n13034) );
  XNOR U15458 ( .A(b[1674]), .B(n13035), .Z(c[1674]) );
  XNOR U15459 ( .A(a[1674]), .B(n13036), .Z(n13035) );
  IV U15460 ( .A(n13033), .Z(n13036) );
  XOR U15461 ( .A(n13037), .B(n13038), .Z(n13033) );
  ANDN U15462 ( .B(n13039), .A(n13040), .Z(n13037) );
  XNOR U15463 ( .A(b[1673]), .B(n13038), .Z(n13039) );
  XNOR U15464 ( .A(b[1673]), .B(n13040), .Z(c[1673]) );
  XNOR U15465 ( .A(a[1673]), .B(n13041), .Z(n13040) );
  IV U15466 ( .A(n13038), .Z(n13041) );
  XOR U15467 ( .A(n13042), .B(n13043), .Z(n13038) );
  ANDN U15468 ( .B(n13044), .A(n13045), .Z(n13042) );
  XNOR U15469 ( .A(b[1672]), .B(n13043), .Z(n13044) );
  XNOR U15470 ( .A(b[1672]), .B(n13045), .Z(c[1672]) );
  XNOR U15471 ( .A(a[1672]), .B(n13046), .Z(n13045) );
  IV U15472 ( .A(n13043), .Z(n13046) );
  XOR U15473 ( .A(n13047), .B(n13048), .Z(n13043) );
  ANDN U15474 ( .B(n13049), .A(n13050), .Z(n13047) );
  XNOR U15475 ( .A(b[1671]), .B(n13048), .Z(n13049) );
  XNOR U15476 ( .A(b[1671]), .B(n13050), .Z(c[1671]) );
  XNOR U15477 ( .A(a[1671]), .B(n13051), .Z(n13050) );
  IV U15478 ( .A(n13048), .Z(n13051) );
  XOR U15479 ( .A(n13052), .B(n13053), .Z(n13048) );
  ANDN U15480 ( .B(n13054), .A(n13055), .Z(n13052) );
  XNOR U15481 ( .A(b[1670]), .B(n13053), .Z(n13054) );
  XNOR U15482 ( .A(b[1670]), .B(n13055), .Z(c[1670]) );
  XNOR U15483 ( .A(a[1670]), .B(n13056), .Z(n13055) );
  IV U15484 ( .A(n13053), .Z(n13056) );
  XOR U15485 ( .A(n13057), .B(n13058), .Z(n13053) );
  ANDN U15486 ( .B(n13059), .A(n13060), .Z(n13057) );
  XNOR U15487 ( .A(b[1669]), .B(n13058), .Z(n13059) );
  XNOR U15488 ( .A(b[166]), .B(n13061), .Z(c[166]) );
  XNOR U15489 ( .A(b[1669]), .B(n13060), .Z(c[1669]) );
  XNOR U15490 ( .A(a[1669]), .B(n13062), .Z(n13060) );
  IV U15491 ( .A(n13058), .Z(n13062) );
  XOR U15492 ( .A(n13063), .B(n13064), .Z(n13058) );
  ANDN U15493 ( .B(n13065), .A(n13066), .Z(n13063) );
  XNOR U15494 ( .A(b[1668]), .B(n13064), .Z(n13065) );
  XNOR U15495 ( .A(b[1668]), .B(n13066), .Z(c[1668]) );
  XNOR U15496 ( .A(a[1668]), .B(n13067), .Z(n13066) );
  IV U15497 ( .A(n13064), .Z(n13067) );
  XOR U15498 ( .A(n13068), .B(n13069), .Z(n13064) );
  ANDN U15499 ( .B(n13070), .A(n13071), .Z(n13068) );
  XNOR U15500 ( .A(b[1667]), .B(n13069), .Z(n13070) );
  XNOR U15501 ( .A(b[1667]), .B(n13071), .Z(c[1667]) );
  XNOR U15502 ( .A(a[1667]), .B(n13072), .Z(n13071) );
  IV U15503 ( .A(n13069), .Z(n13072) );
  XOR U15504 ( .A(n13073), .B(n13074), .Z(n13069) );
  ANDN U15505 ( .B(n13075), .A(n13076), .Z(n13073) );
  XNOR U15506 ( .A(b[1666]), .B(n13074), .Z(n13075) );
  XNOR U15507 ( .A(b[1666]), .B(n13076), .Z(c[1666]) );
  XNOR U15508 ( .A(a[1666]), .B(n13077), .Z(n13076) );
  IV U15509 ( .A(n13074), .Z(n13077) );
  XOR U15510 ( .A(n13078), .B(n13079), .Z(n13074) );
  ANDN U15511 ( .B(n13080), .A(n13081), .Z(n13078) );
  XNOR U15512 ( .A(b[1665]), .B(n13079), .Z(n13080) );
  XNOR U15513 ( .A(b[1665]), .B(n13081), .Z(c[1665]) );
  XNOR U15514 ( .A(a[1665]), .B(n13082), .Z(n13081) );
  IV U15515 ( .A(n13079), .Z(n13082) );
  XOR U15516 ( .A(n13083), .B(n13084), .Z(n13079) );
  ANDN U15517 ( .B(n13085), .A(n13086), .Z(n13083) );
  XNOR U15518 ( .A(b[1664]), .B(n13084), .Z(n13085) );
  XNOR U15519 ( .A(b[1664]), .B(n13086), .Z(c[1664]) );
  XNOR U15520 ( .A(a[1664]), .B(n13087), .Z(n13086) );
  IV U15521 ( .A(n13084), .Z(n13087) );
  XOR U15522 ( .A(n13088), .B(n13089), .Z(n13084) );
  ANDN U15523 ( .B(n13090), .A(n13091), .Z(n13088) );
  XNOR U15524 ( .A(b[1663]), .B(n13089), .Z(n13090) );
  XNOR U15525 ( .A(b[1663]), .B(n13091), .Z(c[1663]) );
  XNOR U15526 ( .A(a[1663]), .B(n13092), .Z(n13091) );
  IV U15527 ( .A(n13089), .Z(n13092) );
  XOR U15528 ( .A(n13093), .B(n13094), .Z(n13089) );
  ANDN U15529 ( .B(n13095), .A(n13096), .Z(n13093) );
  XNOR U15530 ( .A(b[1662]), .B(n13094), .Z(n13095) );
  XNOR U15531 ( .A(b[1662]), .B(n13096), .Z(c[1662]) );
  XNOR U15532 ( .A(a[1662]), .B(n13097), .Z(n13096) );
  IV U15533 ( .A(n13094), .Z(n13097) );
  XOR U15534 ( .A(n13098), .B(n13099), .Z(n13094) );
  ANDN U15535 ( .B(n13100), .A(n13101), .Z(n13098) );
  XNOR U15536 ( .A(b[1661]), .B(n13099), .Z(n13100) );
  XNOR U15537 ( .A(b[1661]), .B(n13101), .Z(c[1661]) );
  XNOR U15538 ( .A(a[1661]), .B(n13102), .Z(n13101) );
  IV U15539 ( .A(n13099), .Z(n13102) );
  XOR U15540 ( .A(n13103), .B(n13104), .Z(n13099) );
  ANDN U15541 ( .B(n13105), .A(n13106), .Z(n13103) );
  XNOR U15542 ( .A(b[1660]), .B(n13104), .Z(n13105) );
  XNOR U15543 ( .A(b[1660]), .B(n13106), .Z(c[1660]) );
  XNOR U15544 ( .A(a[1660]), .B(n13107), .Z(n13106) );
  IV U15545 ( .A(n13104), .Z(n13107) );
  XOR U15546 ( .A(n13108), .B(n13109), .Z(n13104) );
  ANDN U15547 ( .B(n13110), .A(n13111), .Z(n13108) );
  XNOR U15548 ( .A(b[1659]), .B(n13109), .Z(n13110) );
  XNOR U15549 ( .A(b[165]), .B(n13112), .Z(c[165]) );
  XNOR U15550 ( .A(b[1659]), .B(n13111), .Z(c[1659]) );
  XNOR U15551 ( .A(a[1659]), .B(n13113), .Z(n13111) );
  IV U15552 ( .A(n13109), .Z(n13113) );
  XOR U15553 ( .A(n13114), .B(n13115), .Z(n13109) );
  ANDN U15554 ( .B(n13116), .A(n13117), .Z(n13114) );
  XNOR U15555 ( .A(b[1658]), .B(n13115), .Z(n13116) );
  XNOR U15556 ( .A(b[1658]), .B(n13117), .Z(c[1658]) );
  XNOR U15557 ( .A(a[1658]), .B(n13118), .Z(n13117) );
  IV U15558 ( .A(n13115), .Z(n13118) );
  XOR U15559 ( .A(n13119), .B(n13120), .Z(n13115) );
  ANDN U15560 ( .B(n13121), .A(n13122), .Z(n13119) );
  XNOR U15561 ( .A(b[1657]), .B(n13120), .Z(n13121) );
  XNOR U15562 ( .A(b[1657]), .B(n13122), .Z(c[1657]) );
  XNOR U15563 ( .A(a[1657]), .B(n13123), .Z(n13122) );
  IV U15564 ( .A(n13120), .Z(n13123) );
  XOR U15565 ( .A(n13124), .B(n13125), .Z(n13120) );
  ANDN U15566 ( .B(n13126), .A(n13127), .Z(n13124) );
  XNOR U15567 ( .A(b[1656]), .B(n13125), .Z(n13126) );
  XNOR U15568 ( .A(b[1656]), .B(n13127), .Z(c[1656]) );
  XNOR U15569 ( .A(a[1656]), .B(n13128), .Z(n13127) );
  IV U15570 ( .A(n13125), .Z(n13128) );
  XOR U15571 ( .A(n13129), .B(n13130), .Z(n13125) );
  ANDN U15572 ( .B(n13131), .A(n13132), .Z(n13129) );
  XNOR U15573 ( .A(b[1655]), .B(n13130), .Z(n13131) );
  XNOR U15574 ( .A(b[1655]), .B(n13132), .Z(c[1655]) );
  XNOR U15575 ( .A(a[1655]), .B(n13133), .Z(n13132) );
  IV U15576 ( .A(n13130), .Z(n13133) );
  XOR U15577 ( .A(n13134), .B(n13135), .Z(n13130) );
  ANDN U15578 ( .B(n13136), .A(n13137), .Z(n13134) );
  XNOR U15579 ( .A(b[1654]), .B(n13135), .Z(n13136) );
  XNOR U15580 ( .A(b[1654]), .B(n13137), .Z(c[1654]) );
  XNOR U15581 ( .A(a[1654]), .B(n13138), .Z(n13137) );
  IV U15582 ( .A(n13135), .Z(n13138) );
  XOR U15583 ( .A(n13139), .B(n13140), .Z(n13135) );
  ANDN U15584 ( .B(n13141), .A(n13142), .Z(n13139) );
  XNOR U15585 ( .A(b[1653]), .B(n13140), .Z(n13141) );
  XNOR U15586 ( .A(b[1653]), .B(n13142), .Z(c[1653]) );
  XNOR U15587 ( .A(a[1653]), .B(n13143), .Z(n13142) );
  IV U15588 ( .A(n13140), .Z(n13143) );
  XOR U15589 ( .A(n13144), .B(n13145), .Z(n13140) );
  ANDN U15590 ( .B(n13146), .A(n13147), .Z(n13144) );
  XNOR U15591 ( .A(b[1652]), .B(n13145), .Z(n13146) );
  XNOR U15592 ( .A(b[1652]), .B(n13147), .Z(c[1652]) );
  XNOR U15593 ( .A(a[1652]), .B(n13148), .Z(n13147) );
  IV U15594 ( .A(n13145), .Z(n13148) );
  XOR U15595 ( .A(n13149), .B(n13150), .Z(n13145) );
  ANDN U15596 ( .B(n13151), .A(n13152), .Z(n13149) );
  XNOR U15597 ( .A(b[1651]), .B(n13150), .Z(n13151) );
  XNOR U15598 ( .A(b[1651]), .B(n13152), .Z(c[1651]) );
  XNOR U15599 ( .A(a[1651]), .B(n13153), .Z(n13152) );
  IV U15600 ( .A(n13150), .Z(n13153) );
  XOR U15601 ( .A(n13154), .B(n13155), .Z(n13150) );
  ANDN U15602 ( .B(n13156), .A(n13157), .Z(n13154) );
  XNOR U15603 ( .A(b[1650]), .B(n13155), .Z(n13156) );
  XNOR U15604 ( .A(b[1650]), .B(n13157), .Z(c[1650]) );
  XNOR U15605 ( .A(a[1650]), .B(n13158), .Z(n13157) );
  IV U15606 ( .A(n13155), .Z(n13158) );
  XOR U15607 ( .A(n13159), .B(n13160), .Z(n13155) );
  ANDN U15608 ( .B(n13161), .A(n13162), .Z(n13159) );
  XNOR U15609 ( .A(b[1649]), .B(n13160), .Z(n13161) );
  XNOR U15610 ( .A(b[164]), .B(n13163), .Z(c[164]) );
  XNOR U15611 ( .A(b[1649]), .B(n13162), .Z(c[1649]) );
  XNOR U15612 ( .A(a[1649]), .B(n13164), .Z(n13162) );
  IV U15613 ( .A(n13160), .Z(n13164) );
  XOR U15614 ( .A(n13165), .B(n13166), .Z(n13160) );
  ANDN U15615 ( .B(n13167), .A(n13168), .Z(n13165) );
  XNOR U15616 ( .A(b[1648]), .B(n13166), .Z(n13167) );
  XNOR U15617 ( .A(b[1648]), .B(n13168), .Z(c[1648]) );
  XNOR U15618 ( .A(a[1648]), .B(n13169), .Z(n13168) );
  IV U15619 ( .A(n13166), .Z(n13169) );
  XOR U15620 ( .A(n13170), .B(n13171), .Z(n13166) );
  ANDN U15621 ( .B(n13172), .A(n13173), .Z(n13170) );
  XNOR U15622 ( .A(b[1647]), .B(n13171), .Z(n13172) );
  XNOR U15623 ( .A(b[1647]), .B(n13173), .Z(c[1647]) );
  XNOR U15624 ( .A(a[1647]), .B(n13174), .Z(n13173) );
  IV U15625 ( .A(n13171), .Z(n13174) );
  XOR U15626 ( .A(n13175), .B(n13176), .Z(n13171) );
  ANDN U15627 ( .B(n13177), .A(n13178), .Z(n13175) );
  XNOR U15628 ( .A(b[1646]), .B(n13176), .Z(n13177) );
  XNOR U15629 ( .A(b[1646]), .B(n13178), .Z(c[1646]) );
  XNOR U15630 ( .A(a[1646]), .B(n13179), .Z(n13178) );
  IV U15631 ( .A(n13176), .Z(n13179) );
  XOR U15632 ( .A(n13180), .B(n13181), .Z(n13176) );
  ANDN U15633 ( .B(n13182), .A(n13183), .Z(n13180) );
  XNOR U15634 ( .A(b[1645]), .B(n13181), .Z(n13182) );
  XNOR U15635 ( .A(b[1645]), .B(n13183), .Z(c[1645]) );
  XNOR U15636 ( .A(a[1645]), .B(n13184), .Z(n13183) );
  IV U15637 ( .A(n13181), .Z(n13184) );
  XOR U15638 ( .A(n13185), .B(n13186), .Z(n13181) );
  ANDN U15639 ( .B(n13187), .A(n13188), .Z(n13185) );
  XNOR U15640 ( .A(b[1644]), .B(n13186), .Z(n13187) );
  XNOR U15641 ( .A(b[1644]), .B(n13188), .Z(c[1644]) );
  XNOR U15642 ( .A(a[1644]), .B(n13189), .Z(n13188) );
  IV U15643 ( .A(n13186), .Z(n13189) );
  XOR U15644 ( .A(n13190), .B(n13191), .Z(n13186) );
  ANDN U15645 ( .B(n13192), .A(n13193), .Z(n13190) );
  XNOR U15646 ( .A(b[1643]), .B(n13191), .Z(n13192) );
  XNOR U15647 ( .A(b[1643]), .B(n13193), .Z(c[1643]) );
  XNOR U15648 ( .A(a[1643]), .B(n13194), .Z(n13193) );
  IV U15649 ( .A(n13191), .Z(n13194) );
  XOR U15650 ( .A(n13195), .B(n13196), .Z(n13191) );
  ANDN U15651 ( .B(n13197), .A(n13198), .Z(n13195) );
  XNOR U15652 ( .A(b[1642]), .B(n13196), .Z(n13197) );
  XNOR U15653 ( .A(b[1642]), .B(n13198), .Z(c[1642]) );
  XNOR U15654 ( .A(a[1642]), .B(n13199), .Z(n13198) );
  IV U15655 ( .A(n13196), .Z(n13199) );
  XOR U15656 ( .A(n13200), .B(n13201), .Z(n13196) );
  ANDN U15657 ( .B(n13202), .A(n13203), .Z(n13200) );
  XNOR U15658 ( .A(b[1641]), .B(n13201), .Z(n13202) );
  XNOR U15659 ( .A(b[1641]), .B(n13203), .Z(c[1641]) );
  XNOR U15660 ( .A(a[1641]), .B(n13204), .Z(n13203) );
  IV U15661 ( .A(n13201), .Z(n13204) );
  XOR U15662 ( .A(n13205), .B(n13206), .Z(n13201) );
  ANDN U15663 ( .B(n13207), .A(n13208), .Z(n13205) );
  XNOR U15664 ( .A(b[1640]), .B(n13206), .Z(n13207) );
  XNOR U15665 ( .A(b[1640]), .B(n13208), .Z(c[1640]) );
  XNOR U15666 ( .A(a[1640]), .B(n13209), .Z(n13208) );
  IV U15667 ( .A(n13206), .Z(n13209) );
  XOR U15668 ( .A(n13210), .B(n13211), .Z(n13206) );
  ANDN U15669 ( .B(n13212), .A(n13213), .Z(n13210) );
  XNOR U15670 ( .A(b[1639]), .B(n13211), .Z(n13212) );
  XNOR U15671 ( .A(b[163]), .B(n13214), .Z(c[163]) );
  XNOR U15672 ( .A(b[1639]), .B(n13213), .Z(c[1639]) );
  XNOR U15673 ( .A(a[1639]), .B(n13215), .Z(n13213) );
  IV U15674 ( .A(n13211), .Z(n13215) );
  XOR U15675 ( .A(n13216), .B(n13217), .Z(n13211) );
  ANDN U15676 ( .B(n13218), .A(n13219), .Z(n13216) );
  XNOR U15677 ( .A(b[1638]), .B(n13217), .Z(n13218) );
  XNOR U15678 ( .A(b[1638]), .B(n13219), .Z(c[1638]) );
  XNOR U15679 ( .A(a[1638]), .B(n13220), .Z(n13219) );
  IV U15680 ( .A(n13217), .Z(n13220) );
  XOR U15681 ( .A(n13221), .B(n13222), .Z(n13217) );
  ANDN U15682 ( .B(n13223), .A(n13224), .Z(n13221) );
  XNOR U15683 ( .A(b[1637]), .B(n13222), .Z(n13223) );
  XNOR U15684 ( .A(b[1637]), .B(n13224), .Z(c[1637]) );
  XNOR U15685 ( .A(a[1637]), .B(n13225), .Z(n13224) );
  IV U15686 ( .A(n13222), .Z(n13225) );
  XOR U15687 ( .A(n13226), .B(n13227), .Z(n13222) );
  ANDN U15688 ( .B(n13228), .A(n13229), .Z(n13226) );
  XNOR U15689 ( .A(b[1636]), .B(n13227), .Z(n13228) );
  XNOR U15690 ( .A(b[1636]), .B(n13229), .Z(c[1636]) );
  XNOR U15691 ( .A(a[1636]), .B(n13230), .Z(n13229) );
  IV U15692 ( .A(n13227), .Z(n13230) );
  XOR U15693 ( .A(n13231), .B(n13232), .Z(n13227) );
  ANDN U15694 ( .B(n13233), .A(n13234), .Z(n13231) );
  XNOR U15695 ( .A(b[1635]), .B(n13232), .Z(n13233) );
  XNOR U15696 ( .A(b[1635]), .B(n13234), .Z(c[1635]) );
  XNOR U15697 ( .A(a[1635]), .B(n13235), .Z(n13234) );
  IV U15698 ( .A(n13232), .Z(n13235) );
  XOR U15699 ( .A(n13236), .B(n13237), .Z(n13232) );
  ANDN U15700 ( .B(n13238), .A(n13239), .Z(n13236) );
  XNOR U15701 ( .A(b[1634]), .B(n13237), .Z(n13238) );
  XNOR U15702 ( .A(b[1634]), .B(n13239), .Z(c[1634]) );
  XNOR U15703 ( .A(a[1634]), .B(n13240), .Z(n13239) );
  IV U15704 ( .A(n13237), .Z(n13240) );
  XOR U15705 ( .A(n13241), .B(n13242), .Z(n13237) );
  ANDN U15706 ( .B(n13243), .A(n13244), .Z(n13241) );
  XNOR U15707 ( .A(b[1633]), .B(n13242), .Z(n13243) );
  XNOR U15708 ( .A(b[1633]), .B(n13244), .Z(c[1633]) );
  XNOR U15709 ( .A(a[1633]), .B(n13245), .Z(n13244) );
  IV U15710 ( .A(n13242), .Z(n13245) );
  XOR U15711 ( .A(n13246), .B(n13247), .Z(n13242) );
  ANDN U15712 ( .B(n13248), .A(n13249), .Z(n13246) );
  XNOR U15713 ( .A(b[1632]), .B(n13247), .Z(n13248) );
  XNOR U15714 ( .A(b[1632]), .B(n13249), .Z(c[1632]) );
  XNOR U15715 ( .A(a[1632]), .B(n13250), .Z(n13249) );
  IV U15716 ( .A(n13247), .Z(n13250) );
  XOR U15717 ( .A(n13251), .B(n13252), .Z(n13247) );
  ANDN U15718 ( .B(n13253), .A(n13254), .Z(n13251) );
  XNOR U15719 ( .A(b[1631]), .B(n13252), .Z(n13253) );
  XNOR U15720 ( .A(b[1631]), .B(n13254), .Z(c[1631]) );
  XNOR U15721 ( .A(a[1631]), .B(n13255), .Z(n13254) );
  IV U15722 ( .A(n13252), .Z(n13255) );
  XOR U15723 ( .A(n13256), .B(n13257), .Z(n13252) );
  ANDN U15724 ( .B(n13258), .A(n13259), .Z(n13256) );
  XNOR U15725 ( .A(b[1630]), .B(n13257), .Z(n13258) );
  XNOR U15726 ( .A(b[1630]), .B(n13259), .Z(c[1630]) );
  XNOR U15727 ( .A(a[1630]), .B(n13260), .Z(n13259) );
  IV U15728 ( .A(n13257), .Z(n13260) );
  XOR U15729 ( .A(n13261), .B(n13262), .Z(n13257) );
  ANDN U15730 ( .B(n13263), .A(n13264), .Z(n13261) );
  XNOR U15731 ( .A(b[1629]), .B(n13262), .Z(n13263) );
  XNOR U15732 ( .A(b[162]), .B(n13265), .Z(c[162]) );
  XNOR U15733 ( .A(b[1629]), .B(n13264), .Z(c[1629]) );
  XNOR U15734 ( .A(a[1629]), .B(n13266), .Z(n13264) );
  IV U15735 ( .A(n13262), .Z(n13266) );
  XOR U15736 ( .A(n13267), .B(n13268), .Z(n13262) );
  ANDN U15737 ( .B(n13269), .A(n13270), .Z(n13267) );
  XNOR U15738 ( .A(b[1628]), .B(n13268), .Z(n13269) );
  XNOR U15739 ( .A(b[1628]), .B(n13270), .Z(c[1628]) );
  XNOR U15740 ( .A(a[1628]), .B(n13271), .Z(n13270) );
  IV U15741 ( .A(n13268), .Z(n13271) );
  XOR U15742 ( .A(n13272), .B(n13273), .Z(n13268) );
  ANDN U15743 ( .B(n13274), .A(n13275), .Z(n13272) );
  XNOR U15744 ( .A(b[1627]), .B(n13273), .Z(n13274) );
  XNOR U15745 ( .A(b[1627]), .B(n13275), .Z(c[1627]) );
  XNOR U15746 ( .A(a[1627]), .B(n13276), .Z(n13275) );
  IV U15747 ( .A(n13273), .Z(n13276) );
  XOR U15748 ( .A(n13277), .B(n13278), .Z(n13273) );
  ANDN U15749 ( .B(n13279), .A(n13280), .Z(n13277) );
  XNOR U15750 ( .A(b[1626]), .B(n13278), .Z(n13279) );
  XNOR U15751 ( .A(b[1626]), .B(n13280), .Z(c[1626]) );
  XNOR U15752 ( .A(a[1626]), .B(n13281), .Z(n13280) );
  IV U15753 ( .A(n13278), .Z(n13281) );
  XOR U15754 ( .A(n13282), .B(n13283), .Z(n13278) );
  ANDN U15755 ( .B(n13284), .A(n13285), .Z(n13282) );
  XNOR U15756 ( .A(b[1625]), .B(n13283), .Z(n13284) );
  XNOR U15757 ( .A(b[1625]), .B(n13285), .Z(c[1625]) );
  XNOR U15758 ( .A(a[1625]), .B(n13286), .Z(n13285) );
  IV U15759 ( .A(n13283), .Z(n13286) );
  XOR U15760 ( .A(n13287), .B(n13288), .Z(n13283) );
  ANDN U15761 ( .B(n13289), .A(n13290), .Z(n13287) );
  XNOR U15762 ( .A(b[1624]), .B(n13288), .Z(n13289) );
  XNOR U15763 ( .A(b[1624]), .B(n13290), .Z(c[1624]) );
  XNOR U15764 ( .A(a[1624]), .B(n13291), .Z(n13290) );
  IV U15765 ( .A(n13288), .Z(n13291) );
  XOR U15766 ( .A(n13292), .B(n13293), .Z(n13288) );
  ANDN U15767 ( .B(n13294), .A(n13295), .Z(n13292) );
  XNOR U15768 ( .A(b[1623]), .B(n13293), .Z(n13294) );
  XNOR U15769 ( .A(b[1623]), .B(n13295), .Z(c[1623]) );
  XNOR U15770 ( .A(a[1623]), .B(n13296), .Z(n13295) );
  IV U15771 ( .A(n13293), .Z(n13296) );
  XOR U15772 ( .A(n13297), .B(n13298), .Z(n13293) );
  ANDN U15773 ( .B(n13299), .A(n13300), .Z(n13297) );
  XNOR U15774 ( .A(b[1622]), .B(n13298), .Z(n13299) );
  XNOR U15775 ( .A(b[1622]), .B(n13300), .Z(c[1622]) );
  XNOR U15776 ( .A(a[1622]), .B(n13301), .Z(n13300) );
  IV U15777 ( .A(n13298), .Z(n13301) );
  XOR U15778 ( .A(n13302), .B(n13303), .Z(n13298) );
  ANDN U15779 ( .B(n13304), .A(n13305), .Z(n13302) );
  XNOR U15780 ( .A(b[1621]), .B(n13303), .Z(n13304) );
  XNOR U15781 ( .A(b[1621]), .B(n13305), .Z(c[1621]) );
  XNOR U15782 ( .A(a[1621]), .B(n13306), .Z(n13305) );
  IV U15783 ( .A(n13303), .Z(n13306) );
  XOR U15784 ( .A(n13307), .B(n13308), .Z(n13303) );
  ANDN U15785 ( .B(n13309), .A(n13310), .Z(n13307) );
  XNOR U15786 ( .A(b[1620]), .B(n13308), .Z(n13309) );
  XNOR U15787 ( .A(b[1620]), .B(n13310), .Z(c[1620]) );
  XNOR U15788 ( .A(a[1620]), .B(n13311), .Z(n13310) );
  IV U15789 ( .A(n13308), .Z(n13311) );
  XOR U15790 ( .A(n13312), .B(n13313), .Z(n13308) );
  ANDN U15791 ( .B(n13314), .A(n13315), .Z(n13312) );
  XNOR U15792 ( .A(b[1619]), .B(n13313), .Z(n13314) );
  XNOR U15793 ( .A(b[161]), .B(n13316), .Z(c[161]) );
  XNOR U15794 ( .A(b[1619]), .B(n13315), .Z(c[1619]) );
  XNOR U15795 ( .A(a[1619]), .B(n13317), .Z(n13315) );
  IV U15796 ( .A(n13313), .Z(n13317) );
  XOR U15797 ( .A(n13318), .B(n13319), .Z(n13313) );
  ANDN U15798 ( .B(n13320), .A(n13321), .Z(n13318) );
  XNOR U15799 ( .A(b[1618]), .B(n13319), .Z(n13320) );
  XNOR U15800 ( .A(b[1618]), .B(n13321), .Z(c[1618]) );
  XNOR U15801 ( .A(a[1618]), .B(n13322), .Z(n13321) );
  IV U15802 ( .A(n13319), .Z(n13322) );
  XOR U15803 ( .A(n13323), .B(n13324), .Z(n13319) );
  ANDN U15804 ( .B(n13325), .A(n13326), .Z(n13323) );
  XNOR U15805 ( .A(b[1617]), .B(n13324), .Z(n13325) );
  XNOR U15806 ( .A(b[1617]), .B(n13326), .Z(c[1617]) );
  XNOR U15807 ( .A(a[1617]), .B(n13327), .Z(n13326) );
  IV U15808 ( .A(n13324), .Z(n13327) );
  XOR U15809 ( .A(n13328), .B(n13329), .Z(n13324) );
  ANDN U15810 ( .B(n13330), .A(n13331), .Z(n13328) );
  XNOR U15811 ( .A(b[1616]), .B(n13329), .Z(n13330) );
  XNOR U15812 ( .A(b[1616]), .B(n13331), .Z(c[1616]) );
  XNOR U15813 ( .A(a[1616]), .B(n13332), .Z(n13331) );
  IV U15814 ( .A(n13329), .Z(n13332) );
  XOR U15815 ( .A(n13333), .B(n13334), .Z(n13329) );
  ANDN U15816 ( .B(n13335), .A(n13336), .Z(n13333) );
  XNOR U15817 ( .A(b[1615]), .B(n13334), .Z(n13335) );
  XNOR U15818 ( .A(b[1615]), .B(n13336), .Z(c[1615]) );
  XNOR U15819 ( .A(a[1615]), .B(n13337), .Z(n13336) );
  IV U15820 ( .A(n13334), .Z(n13337) );
  XOR U15821 ( .A(n13338), .B(n13339), .Z(n13334) );
  ANDN U15822 ( .B(n13340), .A(n13341), .Z(n13338) );
  XNOR U15823 ( .A(b[1614]), .B(n13339), .Z(n13340) );
  XNOR U15824 ( .A(b[1614]), .B(n13341), .Z(c[1614]) );
  XNOR U15825 ( .A(a[1614]), .B(n13342), .Z(n13341) );
  IV U15826 ( .A(n13339), .Z(n13342) );
  XOR U15827 ( .A(n13343), .B(n13344), .Z(n13339) );
  ANDN U15828 ( .B(n13345), .A(n13346), .Z(n13343) );
  XNOR U15829 ( .A(b[1613]), .B(n13344), .Z(n13345) );
  XNOR U15830 ( .A(b[1613]), .B(n13346), .Z(c[1613]) );
  XNOR U15831 ( .A(a[1613]), .B(n13347), .Z(n13346) );
  IV U15832 ( .A(n13344), .Z(n13347) );
  XOR U15833 ( .A(n13348), .B(n13349), .Z(n13344) );
  ANDN U15834 ( .B(n13350), .A(n13351), .Z(n13348) );
  XNOR U15835 ( .A(b[1612]), .B(n13349), .Z(n13350) );
  XNOR U15836 ( .A(b[1612]), .B(n13351), .Z(c[1612]) );
  XNOR U15837 ( .A(a[1612]), .B(n13352), .Z(n13351) );
  IV U15838 ( .A(n13349), .Z(n13352) );
  XOR U15839 ( .A(n13353), .B(n13354), .Z(n13349) );
  ANDN U15840 ( .B(n13355), .A(n13356), .Z(n13353) );
  XNOR U15841 ( .A(b[1611]), .B(n13354), .Z(n13355) );
  XNOR U15842 ( .A(b[1611]), .B(n13356), .Z(c[1611]) );
  XNOR U15843 ( .A(a[1611]), .B(n13357), .Z(n13356) );
  IV U15844 ( .A(n13354), .Z(n13357) );
  XOR U15845 ( .A(n13358), .B(n13359), .Z(n13354) );
  ANDN U15846 ( .B(n13360), .A(n13361), .Z(n13358) );
  XNOR U15847 ( .A(b[1610]), .B(n13359), .Z(n13360) );
  XNOR U15848 ( .A(b[1610]), .B(n13361), .Z(c[1610]) );
  XNOR U15849 ( .A(a[1610]), .B(n13362), .Z(n13361) );
  IV U15850 ( .A(n13359), .Z(n13362) );
  XOR U15851 ( .A(n13363), .B(n13364), .Z(n13359) );
  ANDN U15852 ( .B(n13365), .A(n13366), .Z(n13363) );
  XNOR U15853 ( .A(b[1609]), .B(n13364), .Z(n13365) );
  XNOR U15854 ( .A(b[160]), .B(n13367), .Z(c[160]) );
  XNOR U15855 ( .A(b[1609]), .B(n13366), .Z(c[1609]) );
  XNOR U15856 ( .A(a[1609]), .B(n13368), .Z(n13366) );
  IV U15857 ( .A(n13364), .Z(n13368) );
  XOR U15858 ( .A(n13369), .B(n13370), .Z(n13364) );
  ANDN U15859 ( .B(n13371), .A(n13372), .Z(n13369) );
  XNOR U15860 ( .A(b[1608]), .B(n13370), .Z(n13371) );
  XNOR U15861 ( .A(b[1608]), .B(n13372), .Z(c[1608]) );
  XNOR U15862 ( .A(a[1608]), .B(n13373), .Z(n13372) );
  IV U15863 ( .A(n13370), .Z(n13373) );
  XOR U15864 ( .A(n13374), .B(n13375), .Z(n13370) );
  ANDN U15865 ( .B(n13376), .A(n13377), .Z(n13374) );
  XNOR U15866 ( .A(b[1607]), .B(n13375), .Z(n13376) );
  XNOR U15867 ( .A(b[1607]), .B(n13377), .Z(c[1607]) );
  XNOR U15868 ( .A(a[1607]), .B(n13378), .Z(n13377) );
  IV U15869 ( .A(n13375), .Z(n13378) );
  XOR U15870 ( .A(n13379), .B(n13380), .Z(n13375) );
  ANDN U15871 ( .B(n13381), .A(n13382), .Z(n13379) );
  XNOR U15872 ( .A(b[1606]), .B(n13380), .Z(n13381) );
  XNOR U15873 ( .A(b[1606]), .B(n13382), .Z(c[1606]) );
  XNOR U15874 ( .A(a[1606]), .B(n13383), .Z(n13382) );
  IV U15875 ( .A(n13380), .Z(n13383) );
  XOR U15876 ( .A(n13384), .B(n13385), .Z(n13380) );
  ANDN U15877 ( .B(n13386), .A(n13387), .Z(n13384) );
  XNOR U15878 ( .A(b[1605]), .B(n13385), .Z(n13386) );
  XNOR U15879 ( .A(b[1605]), .B(n13387), .Z(c[1605]) );
  XNOR U15880 ( .A(a[1605]), .B(n13388), .Z(n13387) );
  IV U15881 ( .A(n13385), .Z(n13388) );
  XOR U15882 ( .A(n13389), .B(n13390), .Z(n13385) );
  ANDN U15883 ( .B(n13391), .A(n13392), .Z(n13389) );
  XNOR U15884 ( .A(b[1604]), .B(n13390), .Z(n13391) );
  XNOR U15885 ( .A(b[1604]), .B(n13392), .Z(c[1604]) );
  XNOR U15886 ( .A(a[1604]), .B(n13393), .Z(n13392) );
  IV U15887 ( .A(n13390), .Z(n13393) );
  XOR U15888 ( .A(n13394), .B(n13395), .Z(n13390) );
  ANDN U15889 ( .B(n13396), .A(n13397), .Z(n13394) );
  XNOR U15890 ( .A(b[1603]), .B(n13395), .Z(n13396) );
  XNOR U15891 ( .A(b[1603]), .B(n13397), .Z(c[1603]) );
  XNOR U15892 ( .A(a[1603]), .B(n13398), .Z(n13397) );
  IV U15893 ( .A(n13395), .Z(n13398) );
  XOR U15894 ( .A(n13399), .B(n13400), .Z(n13395) );
  ANDN U15895 ( .B(n13401), .A(n13402), .Z(n13399) );
  XNOR U15896 ( .A(b[1602]), .B(n13400), .Z(n13401) );
  XNOR U15897 ( .A(b[1602]), .B(n13402), .Z(c[1602]) );
  XNOR U15898 ( .A(a[1602]), .B(n13403), .Z(n13402) );
  IV U15899 ( .A(n13400), .Z(n13403) );
  XOR U15900 ( .A(n13404), .B(n13405), .Z(n13400) );
  ANDN U15901 ( .B(n13406), .A(n13407), .Z(n13404) );
  XNOR U15902 ( .A(b[1601]), .B(n13405), .Z(n13406) );
  XNOR U15903 ( .A(b[1601]), .B(n13407), .Z(c[1601]) );
  XNOR U15904 ( .A(a[1601]), .B(n13408), .Z(n13407) );
  IV U15905 ( .A(n13405), .Z(n13408) );
  XOR U15906 ( .A(n13409), .B(n13410), .Z(n13405) );
  ANDN U15907 ( .B(n13411), .A(n13412), .Z(n13409) );
  XNOR U15908 ( .A(b[1600]), .B(n13410), .Z(n13411) );
  XNOR U15909 ( .A(b[1600]), .B(n13412), .Z(c[1600]) );
  XNOR U15910 ( .A(a[1600]), .B(n13413), .Z(n13412) );
  IV U15911 ( .A(n13410), .Z(n13413) );
  XOR U15912 ( .A(n13414), .B(n13415), .Z(n13410) );
  ANDN U15913 ( .B(n13416), .A(n13417), .Z(n13414) );
  XNOR U15914 ( .A(b[1599]), .B(n13415), .Z(n13416) );
  XNOR U15915 ( .A(b[15]), .B(n13418), .Z(c[15]) );
  XNOR U15916 ( .A(b[159]), .B(n13419), .Z(c[159]) );
  XNOR U15917 ( .A(b[1599]), .B(n13417), .Z(c[1599]) );
  XNOR U15918 ( .A(a[1599]), .B(n13420), .Z(n13417) );
  IV U15919 ( .A(n13415), .Z(n13420) );
  XOR U15920 ( .A(n13421), .B(n13422), .Z(n13415) );
  ANDN U15921 ( .B(n13423), .A(n13424), .Z(n13421) );
  XNOR U15922 ( .A(b[1598]), .B(n13422), .Z(n13423) );
  XNOR U15923 ( .A(b[1598]), .B(n13424), .Z(c[1598]) );
  XNOR U15924 ( .A(a[1598]), .B(n13425), .Z(n13424) );
  IV U15925 ( .A(n13422), .Z(n13425) );
  XOR U15926 ( .A(n13426), .B(n13427), .Z(n13422) );
  ANDN U15927 ( .B(n13428), .A(n13429), .Z(n13426) );
  XNOR U15928 ( .A(b[1597]), .B(n13427), .Z(n13428) );
  XNOR U15929 ( .A(b[1597]), .B(n13429), .Z(c[1597]) );
  XNOR U15930 ( .A(a[1597]), .B(n13430), .Z(n13429) );
  IV U15931 ( .A(n13427), .Z(n13430) );
  XOR U15932 ( .A(n13431), .B(n13432), .Z(n13427) );
  ANDN U15933 ( .B(n13433), .A(n13434), .Z(n13431) );
  XNOR U15934 ( .A(b[1596]), .B(n13432), .Z(n13433) );
  XNOR U15935 ( .A(b[1596]), .B(n13434), .Z(c[1596]) );
  XNOR U15936 ( .A(a[1596]), .B(n13435), .Z(n13434) );
  IV U15937 ( .A(n13432), .Z(n13435) );
  XOR U15938 ( .A(n13436), .B(n13437), .Z(n13432) );
  ANDN U15939 ( .B(n13438), .A(n13439), .Z(n13436) );
  XNOR U15940 ( .A(b[1595]), .B(n13437), .Z(n13438) );
  XNOR U15941 ( .A(b[1595]), .B(n13439), .Z(c[1595]) );
  XNOR U15942 ( .A(a[1595]), .B(n13440), .Z(n13439) );
  IV U15943 ( .A(n13437), .Z(n13440) );
  XOR U15944 ( .A(n13441), .B(n13442), .Z(n13437) );
  ANDN U15945 ( .B(n13443), .A(n13444), .Z(n13441) );
  XNOR U15946 ( .A(b[1594]), .B(n13442), .Z(n13443) );
  XNOR U15947 ( .A(b[1594]), .B(n13444), .Z(c[1594]) );
  XNOR U15948 ( .A(a[1594]), .B(n13445), .Z(n13444) );
  IV U15949 ( .A(n13442), .Z(n13445) );
  XOR U15950 ( .A(n13446), .B(n13447), .Z(n13442) );
  ANDN U15951 ( .B(n13448), .A(n13449), .Z(n13446) );
  XNOR U15952 ( .A(b[1593]), .B(n13447), .Z(n13448) );
  XNOR U15953 ( .A(b[1593]), .B(n13449), .Z(c[1593]) );
  XNOR U15954 ( .A(a[1593]), .B(n13450), .Z(n13449) );
  IV U15955 ( .A(n13447), .Z(n13450) );
  XOR U15956 ( .A(n13451), .B(n13452), .Z(n13447) );
  ANDN U15957 ( .B(n13453), .A(n13454), .Z(n13451) );
  XNOR U15958 ( .A(b[1592]), .B(n13452), .Z(n13453) );
  XNOR U15959 ( .A(b[1592]), .B(n13454), .Z(c[1592]) );
  XNOR U15960 ( .A(a[1592]), .B(n13455), .Z(n13454) );
  IV U15961 ( .A(n13452), .Z(n13455) );
  XOR U15962 ( .A(n13456), .B(n13457), .Z(n13452) );
  ANDN U15963 ( .B(n13458), .A(n13459), .Z(n13456) );
  XNOR U15964 ( .A(b[1591]), .B(n13457), .Z(n13458) );
  XNOR U15965 ( .A(b[1591]), .B(n13459), .Z(c[1591]) );
  XNOR U15966 ( .A(a[1591]), .B(n13460), .Z(n13459) );
  IV U15967 ( .A(n13457), .Z(n13460) );
  XOR U15968 ( .A(n13461), .B(n13462), .Z(n13457) );
  ANDN U15969 ( .B(n13463), .A(n13464), .Z(n13461) );
  XNOR U15970 ( .A(b[1590]), .B(n13462), .Z(n13463) );
  XNOR U15971 ( .A(b[1590]), .B(n13464), .Z(c[1590]) );
  XNOR U15972 ( .A(a[1590]), .B(n13465), .Z(n13464) );
  IV U15973 ( .A(n13462), .Z(n13465) );
  XOR U15974 ( .A(n13466), .B(n13467), .Z(n13462) );
  ANDN U15975 ( .B(n13468), .A(n13469), .Z(n13466) );
  XNOR U15976 ( .A(b[1589]), .B(n13467), .Z(n13468) );
  XNOR U15977 ( .A(b[158]), .B(n13470), .Z(c[158]) );
  XNOR U15978 ( .A(b[1589]), .B(n13469), .Z(c[1589]) );
  XNOR U15979 ( .A(a[1589]), .B(n13471), .Z(n13469) );
  IV U15980 ( .A(n13467), .Z(n13471) );
  XOR U15981 ( .A(n13472), .B(n13473), .Z(n13467) );
  ANDN U15982 ( .B(n13474), .A(n13475), .Z(n13472) );
  XNOR U15983 ( .A(b[1588]), .B(n13473), .Z(n13474) );
  XNOR U15984 ( .A(b[1588]), .B(n13475), .Z(c[1588]) );
  XNOR U15985 ( .A(a[1588]), .B(n13476), .Z(n13475) );
  IV U15986 ( .A(n13473), .Z(n13476) );
  XOR U15987 ( .A(n13477), .B(n13478), .Z(n13473) );
  ANDN U15988 ( .B(n13479), .A(n13480), .Z(n13477) );
  XNOR U15989 ( .A(b[1587]), .B(n13478), .Z(n13479) );
  XNOR U15990 ( .A(b[1587]), .B(n13480), .Z(c[1587]) );
  XNOR U15991 ( .A(a[1587]), .B(n13481), .Z(n13480) );
  IV U15992 ( .A(n13478), .Z(n13481) );
  XOR U15993 ( .A(n13482), .B(n13483), .Z(n13478) );
  ANDN U15994 ( .B(n13484), .A(n13485), .Z(n13482) );
  XNOR U15995 ( .A(b[1586]), .B(n13483), .Z(n13484) );
  XNOR U15996 ( .A(b[1586]), .B(n13485), .Z(c[1586]) );
  XNOR U15997 ( .A(a[1586]), .B(n13486), .Z(n13485) );
  IV U15998 ( .A(n13483), .Z(n13486) );
  XOR U15999 ( .A(n13487), .B(n13488), .Z(n13483) );
  ANDN U16000 ( .B(n13489), .A(n13490), .Z(n13487) );
  XNOR U16001 ( .A(b[1585]), .B(n13488), .Z(n13489) );
  XNOR U16002 ( .A(b[1585]), .B(n13490), .Z(c[1585]) );
  XNOR U16003 ( .A(a[1585]), .B(n13491), .Z(n13490) );
  IV U16004 ( .A(n13488), .Z(n13491) );
  XOR U16005 ( .A(n13492), .B(n13493), .Z(n13488) );
  ANDN U16006 ( .B(n13494), .A(n13495), .Z(n13492) );
  XNOR U16007 ( .A(b[1584]), .B(n13493), .Z(n13494) );
  XNOR U16008 ( .A(b[1584]), .B(n13495), .Z(c[1584]) );
  XNOR U16009 ( .A(a[1584]), .B(n13496), .Z(n13495) );
  IV U16010 ( .A(n13493), .Z(n13496) );
  XOR U16011 ( .A(n13497), .B(n13498), .Z(n13493) );
  ANDN U16012 ( .B(n13499), .A(n13500), .Z(n13497) );
  XNOR U16013 ( .A(b[1583]), .B(n13498), .Z(n13499) );
  XNOR U16014 ( .A(b[1583]), .B(n13500), .Z(c[1583]) );
  XNOR U16015 ( .A(a[1583]), .B(n13501), .Z(n13500) );
  IV U16016 ( .A(n13498), .Z(n13501) );
  XOR U16017 ( .A(n13502), .B(n13503), .Z(n13498) );
  ANDN U16018 ( .B(n13504), .A(n13505), .Z(n13502) );
  XNOR U16019 ( .A(b[1582]), .B(n13503), .Z(n13504) );
  XNOR U16020 ( .A(b[1582]), .B(n13505), .Z(c[1582]) );
  XNOR U16021 ( .A(a[1582]), .B(n13506), .Z(n13505) );
  IV U16022 ( .A(n13503), .Z(n13506) );
  XOR U16023 ( .A(n13507), .B(n13508), .Z(n13503) );
  ANDN U16024 ( .B(n13509), .A(n13510), .Z(n13507) );
  XNOR U16025 ( .A(b[1581]), .B(n13508), .Z(n13509) );
  XNOR U16026 ( .A(b[1581]), .B(n13510), .Z(c[1581]) );
  XNOR U16027 ( .A(a[1581]), .B(n13511), .Z(n13510) );
  IV U16028 ( .A(n13508), .Z(n13511) );
  XOR U16029 ( .A(n13512), .B(n13513), .Z(n13508) );
  ANDN U16030 ( .B(n13514), .A(n13515), .Z(n13512) );
  XNOR U16031 ( .A(b[1580]), .B(n13513), .Z(n13514) );
  XNOR U16032 ( .A(b[1580]), .B(n13515), .Z(c[1580]) );
  XNOR U16033 ( .A(a[1580]), .B(n13516), .Z(n13515) );
  IV U16034 ( .A(n13513), .Z(n13516) );
  XOR U16035 ( .A(n13517), .B(n13518), .Z(n13513) );
  ANDN U16036 ( .B(n13519), .A(n13520), .Z(n13517) );
  XNOR U16037 ( .A(b[1579]), .B(n13518), .Z(n13519) );
  XNOR U16038 ( .A(b[157]), .B(n13521), .Z(c[157]) );
  XNOR U16039 ( .A(b[1579]), .B(n13520), .Z(c[1579]) );
  XNOR U16040 ( .A(a[1579]), .B(n13522), .Z(n13520) );
  IV U16041 ( .A(n13518), .Z(n13522) );
  XOR U16042 ( .A(n13523), .B(n13524), .Z(n13518) );
  ANDN U16043 ( .B(n13525), .A(n13526), .Z(n13523) );
  XNOR U16044 ( .A(b[1578]), .B(n13524), .Z(n13525) );
  XNOR U16045 ( .A(b[1578]), .B(n13526), .Z(c[1578]) );
  XNOR U16046 ( .A(a[1578]), .B(n13527), .Z(n13526) );
  IV U16047 ( .A(n13524), .Z(n13527) );
  XOR U16048 ( .A(n13528), .B(n13529), .Z(n13524) );
  ANDN U16049 ( .B(n13530), .A(n13531), .Z(n13528) );
  XNOR U16050 ( .A(b[1577]), .B(n13529), .Z(n13530) );
  XNOR U16051 ( .A(b[1577]), .B(n13531), .Z(c[1577]) );
  XNOR U16052 ( .A(a[1577]), .B(n13532), .Z(n13531) );
  IV U16053 ( .A(n13529), .Z(n13532) );
  XOR U16054 ( .A(n13533), .B(n13534), .Z(n13529) );
  ANDN U16055 ( .B(n13535), .A(n13536), .Z(n13533) );
  XNOR U16056 ( .A(b[1576]), .B(n13534), .Z(n13535) );
  XNOR U16057 ( .A(b[1576]), .B(n13536), .Z(c[1576]) );
  XNOR U16058 ( .A(a[1576]), .B(n13537), .Z(n13536) );
  IV U16059 ( .A(n13534), .Z(n13537) );
  XOR U16060 ( .A(n13538), .B(n13539), .Z(n13534) );
  ANDN U16061 ( .B(n13540), .A(n13541), .Z(n13538) );
  XNOR U16062 ( .A(b[1575]), .B(n13539), .Z(n13540) );
  XNOR U16063 ( .A(b[1575]), .B(n13541), .Z(c[1575]) );
  XNOR U16064 ( .A(a[1575]), .B(n13542), .Z(n13541) );
  IV U16065 ( .A(n13539), .Z(n13542) );
  XOR U16066 ( .A(n13543), .B(n13544), .Z(n13539) );
  ANDN U16067 ( .B(n13545), .A(n13546), .Z(n13543) );
  XNOR U16068 ( .A(b[1574]), .B(n13544), .Z(n13545) );
  XNOR U16069 ( .A(b[1574]), .B(n13546), .Z(c[1574]) );
  XNOR U16070 ( .A(a[1574]), .B(n13547), .Z(n13546) );
  IV U16071 ( .A(n13544), .Z(n13547) );
  XOR U16072 ( .A(n13548), .B(n13549), .Z(n13544) );
  ANDN U16073 ( .B(n13550), .A(n13551), .Z(n13548) );
  XNOR U16074 ( .A(b[1573]), .B(n13549), .Z(n13550) );
  XNOR U16075 ( .A(b[1573]), .B(n13551), .Z(c[1573]) );
  XNOR U16076 ( .A(a[1573]), .B(n13552), .Z(n13551) );
  IV U16077 ( .A(n13549), .Z(n13552) );
  XOR U16078 ( .A(n13553), .B(n13554), .Z(n13549) );
  ANDN U16079 ( .B(n13555), .A(n13556), .Z(n13553) );
  XNOR U16080 ( .A(b[1572]), .B(n13554), .Z(n13555) );
  XNOR U16081 ( .A(b[1572]), .B(n13556), .Z(c[1572]) );
  XNOR U16082 ( .A(a[1572]), .B(n13557), .Z(n13556) );
  IV U16083 ( .A(n13554), .Z(n13557) );
  XOR U16084 ( .A(n13558), .B(n13559), .Z(n13554) );
  ANDN U16085 ( .B(n13560), .A(n13561), .Z(n13558) );
  XNOR U16086 ( .A(b[1571]), .B(n13559), .Z(n13560) );
  XNOR U16087 ( .A(b[1571]), .B(n13561), .Z(c[1571]) );
  XNOR U16088 ( .A(a[1571]), .B(n13562), .Z(n13561) );
  IV U16089 ( .A(n13559), .Z(n13562) );
  XOR U16090 ( .A(n13563), .B(n13564), .Z(n13559) );
  ANDN U16091 ( .B(n13565), .A(n13566), .Z(n13563) );
  XNOR U16092 ( .A(b[1570]), .B(n13564), .Z(n13565) );
  XNOR U16093 ( .A(b[1570]), .B(n13566), .Z(c[1570]) );
  XNOR U16094 ( .A(a[1570]), .B(n13567), .Z(n13566) );
  IV U16095 ( .A(n13564), .Z(n13567) );
  XOR U16096 ( .A(n13568), .B(n13569), .Z(n13564) );
  ANDN U16097 ( .B(n13570), .A(n13571), .Z(n13568) );
  XNOR U16098 ( .A(b[1569]), .B(n13569), .Z(n13570) );
  XNOR U16099 ( .A(b[156]), .B(n13572), .Z(c[156]) );
  XNOR U16100 ( .A(b[1569]), .B(n13571), .Z(c[1569]) );
  XNOR U16101 ( .A(a[1569]), .B(n13573), .Z(n13571) );
  IV U16102 ( .A(n13569), .Z(n13573) );
  XOR U16103 ( .A(n13574), .B(n13575), .Z(n13569) );
  ANDN U16104 ( .B(n13576), .A(n13577), .Z(n13574) );
  XNOR U16105 ( .A(b[1568]), .B(n13575), .Z(n13576) );
  XNOR U16106 ( .A(b[1568]), .B(n13577), .Z(c[1568]) );
  XNOR U16107 ( .A(a[1568]), .B(n13578), .Z(n13577) );
  IV U16108 ( .A(n13575), .Z(n13578) );
  XOR U16109 ( .A(n13579), .B(n13580), .Z(n13575) );
  ANDN U16110 ( .B(n13581), .A(n13582), .Z(n13579) );
  XNOR U16111 ( .A(b[1567]), .B(n13580), .Z(n13581) );
  XNOR U16112 ( .A(b[1567]), .B(n13582), .Z(c[1567]) );
  XNOR U16113 ( .A(a[1567]), .B(n13583), .Z(n13582) );
  IV U16114 ( .A(n13580), .Z(n13583) );
  XOR U16115 ( .A(n13584), .B(n13585), .Z(n13580) );
  ANDN U16116 ( .B(n13586), .A(n13587), .Z(n13584) );
  XNOR U16117 ( .A(b[1566]), .B(n13585), .Z(n13586) );
  XNOR U16118 ( .A(b[1566]), .B(n13587), .Z(c[1566]) );
  XNOR U16119 ( .A(a[1566]), .B(n13588), .Z(n13587) );
  IV U16120 ( .A(n13585), .Z(n13588) );
  XOR U16121 ( .A(n13589), .B(n13590), .Z(n13585) );
  ANDN U16122 ( .B(n13591), .A(n13592), .Z(n13589) );
  XNOR U16123 ( .A(b[1565]), .B(n13590), .Z(n13591) );
  XNOR U16124 ( .A(b[1565]), .B(n13592), .Z(c[1565]) );
  XNOR U16125 ( .A(a[1565]), .B(n13593), .Z(n13592) );
  IV U16126 ( .A(n13590), .Z(n13593) );
  XOR U16127 ( .A(n13594), .B(n13595), .Z(n13590) );
  ANDN U16128 ( .B(n13596), .A(n13597), .Z(n13594) );
  XNOR U16129 ( .A(b[1564]), .B(n13595), .Z(n13596) );
  XNOR U16130 ( .A(b[1564]), .B(n13597), .Z(c[1564]) );
  XNOR U16131 ( .A(a[1564]), .B(n13598), .Z(n13597) );
  IV U16132 ( .A(n13595), .Z(n13598) );
  XOR U16133 ( .A(n13599), .B(n13600), .Z(n13595) );
  ANDN U16134 ( .B(n13601), .A(n13602), .Z(n13599) );
  XNOR U16135 ( .A(b[1563]), .B(n13600), .Z(n13601) );
  XNOR U16136 ( .A(b[1563]), .B(n13602), .Z(c[1563]) );
  XNOR U16137 ( .A(a[1563]), .B(n13603), .Z(n13602) );
  IV U16138 ( .A(n13600), .Z(n13603) );
  XOR U16139 ( .A(n13604), .B(n13605), .Z(n13600) );
  ANDN U16140 ( .B(n13606), .A(n13607), .Z(n13604) );
  XNOR U16141 ( .A(b[1562]), .B(n13605), .Z(n13606) );
  XNOR U16142 ( .A(b[1562]), .B(n13607), .Z(c[1562]) );
  XNOR U16143 ( .A(a[1562]), .B(n13608), .Z(n13607) );
  IV U16144 ( .A(n13605), .Z(n13608) );
  XOR U16145 ( .A(n13609), .B(n13610), .Z(n13605) );
  ANDN U16146 ( .B(n13611), .A(n13612), .Z(n13609) );
  XNOR U16147 ( .A(b[1561]), .B(n13610), .Z(n13611) );
  XNOR U16148 ( .A(b[1561]), .B(n13612), .Z(c[1561]) );
  XNOR U16149 ( .A(a[1561]), .B(n13613), .Z(n13612) );
  IV U16150 ( .A(n13610), .Z(n13613) );
  XOR U16151 ( .A(n13614), .B(n13615), .Z(n13610) );
  ANDN U16152 ( .B(n13616), .A(n13617), .Z(n13614) );
  XNOR U16153 ( .A(b[1560]), .B(n13615), .Z(n13616) );
  XNOR U16154 ( .A(b[1560]), .B(n13617), .Z(c[1560]) );
  XNOR U16155 ( .A(a[1560]), .B(n13618), .Z(n13617) );
  IV U16156 ( .A(n13615), .Z(n13618) );
  XOR U16157 ( .A(n13619), .B(n13620), .Z(n13615) );
  ANDN U16158 ( .B(n13621), .A(n13622), .Z(n13619) );
  XNOR U16159 ( .A(b[1559]), .B(n13620), .Z(n13621) );
  XNOR U16160 ( .A(b[155]), .B(n13623), .Z(c[155]) );
  XNOR U16161 ( .A(b[1559]), .B(n13622), .Z(c[1559]) );
  XNOR U16162 ( .A(a[1559]), .B(n13624), .Z(n13622) );
  IV U16163 ( .A(n13620), .Z(n13624) );
  XOR U16164 ( .A(n13625), .B(n13626), .Z(n13620) );
  ANDN U16165 ( .B(n13627), .A(n13628), .Z(n13625) );
  XNOR U16166 ( .A(b[1558]), .B(n13626), .Z(n13627) );
  XNOR U16167 ( .A(b[1558]), .B(n13628), .Z(c[1558]) );
  XNOR U16168 ( .A(a[1558]), .B(n13629), .Z(n13628) );
  IV U16169 ( .A(n13626), .Z(n13629) );
  XOR U16170 ( .A(n13630), .B(n13631), .Z(n13626) );
  ANDN U16171 ( .B(n13632), .A(n13633), .Z(n13630) );
  XNOR U16172 ( .A(b[1557]), .B(n13631), .Z(n13632) );
  XNOR U16173 ( .A(b[1557]), .B(n13633), .Z(c[1557]) );
  XNOR U16174 ( .A(a[1557]), .B(n13634), .Z(n13633) );
  IV U16175 ( .A(n13631), .Z(n13634) );
  XOR U16176 ( .A(n13635), .B(n13636), .Z(n13631) );
  ANDN U16177 ( .B(n13637), .A(n13638), .Z(n13635) );
  XNOR U16178 ( .A(b[1556]), .B(n13636), .Z(n13637) );
  XNOR U16179 ( .A(b[1556]), .B(n13638), .Z(c[1556]) );
  XNOR U16180 ( .A(a[1556]), .B(n13639), .Z(n13638) );
  IV U16181 ( .A(n13636), .Z(n13639) );
  XOR U16182 ( .A(n13640), .B(n13641), .Z(n13636) );
  ANDN U16183 ( .B(n13642), .A(n13643), .Z(n13640) );
  XNOR U16184 ( .A(b[1555]), .B(n13641), .Z(n13642) );
  XNOR U16185 ( .A(b[1555]), .B(n13643), .Z(c[1555]) );
  XNOR U16186 ( .A(a[1555]), .B(n13644), .Z(n13643) );
  IV U16187 ( .A(n13641), .Z(n13644) );
  XOR U16188 ( .A(n13645), .B(n13646), .Z(n13641) );
  ANDN U16189 ( .B(n13647), .A(n13648), .Z(n13645) );
  XNOR U16190 ( .A(b[1554]), .B(n13646), .Z(n13647) );
  XNOR U16191 ( .A(b[1554]), .B(n13648), .Z(c[1554]) );
  XNOR U16192 ( .A(a[1554]), .B(n13649), .Z(n13648) );
  IV U16193 ( .A(n13646), .Z(n13649) );
  XOR U16194 ( .A(n13650), .B(n13651), .Z(n13646) );
  ANDN U16195 ( .B(n13652), .A(n13653), .Z(n13650) );
  XNOR U16196 ( .A(b[1553]), .B(n13651), .Z(n13652) );
  XNOR U16197 ( .A(b[1553]), .B(n13653), .Z(c[1553]) );
  XNOR U16198 ( .A(a[1553]), .B(n13654), .Z(n13653) );
  IV U16199 ( .A(n13651), .Z(n13654) );
  XOR U16200 ( .A(n13655), .B(n13656), .Z(n13651) );
  ANDN U16201 ( .B(n13657), .A(n13658), .Z(n13655) );
  XNOR U16202 ( .A(b[1552]), .B(n13656), .Z(n13657) );
  XNOR U16203 ( .A(b[1552]), .B(n13658), .Z(c[1552]) );
  XNOR U16204 ( .A(a[1552]), .B(n13659), .Z(n13658) );
  IV U16205 ( .A(n13656), .Z(n13659) );
  XOR U16206 ( .A(n13660), .B(n13661), .Z(n13656) );
  ANDN U16207 ( .B(n13662), .A(n13663), .Z(n13660) );
  XNOR U16208 ( .A(b[1551]), .B(n13661), .Z(n13662) );
  XNOR U16209 ( .A(b[1551]), .B(n13663), .Z(c[1551]) );
  XNOR U16210 ( .A(a[1551]), .B(n13664), .Z(n13663) );
  IV U16211 ( .A(n13661), .Z(n13664) );
  XOR U16212 ( .A(n13665), .B(n13666), .Z(n13661) );
  ANDN U16213 ( .B(n13667), .A(n13668), .Z(n13665) );
  XNOR U16214 ( .A(b[1550]), .B(n13666), .Z(n13667) );
  XNOR U16215 ( .A(b[1550]), .B(n13668), .Z(c[1550]) );
  XNOR U16216 ( .A(a[1550]), .B(n13669), .Z(n13668) );
  IV U16217 ( .A(n13666), .Z(n13669) );
  XOR U16218 ( .A(n13670), .B(n13671), .Z(n13666) );
  ANDN U16219 ( .B(n13672), .A(n13673), .Z(n13670) );
  XNOR U16220 ( .A(b[1549]), .B(n13671), .Z(n13672) );
  XNOR U16221 ( .A(b[154]), .B(n13674), .Z(c[154]) );
  XNOR U16222 ( .A(b[1549]), .B(n13673), .Z(c[1549]) );
  XNOR U16223 ( .A(a[1549]), .B(n13675), .Z(n13673) );
  IV U16224 ( .A(n13671), .Z(n13675) );
  XOR U16225 ( .A(n13676), .B(n13677), .Z(n13671) );
  ANDN U16226 ( .B(n13678), .A(n13679), .Z(n13676) );
  XNOR U16227 ( .A(b[1548]), .B(n13677), .Z(n13678) );
  XNOR U16228 ( .A(b[1548]), .B(n13679), .Z(c[1548]) );
  XNOR U16229 ( .A(a[1548]), .B(n13680), .Z(n13679) );
  IV U16230 ( .A(n13677), .Z(n13680) );
  XOR U16231 ( .A(n13681), .B(n13682), .Z(n13677) );
  ANDN U16232 ( .B(n13683), .A(n13684), .Z(n13681) );
  XNOR U16233 ( .A(b[1547]), .B(n13682), .Z(n13683) );
  XNOR U16234 ( .A(b[1547]), .B(n13684), .Z(c[1547]) );
  XNOR U16235 ( .A(a[1547]), .B(n13685), .Z(n13684) );
  IV U16236 ( .A(n13682), .Z(n13685) );
  XOR U16237 ( .A(n13686), .B(n13687), .Z(n13682) );
  ANDN U16238 ( .B(n13688), .A(n13689), .Z(n13686) );
  XNOR U16239 ( .A(b[1546]), .B(n13687), .Z(n13688) );
  XNOR U16240 ( .A(b[1546]), .B(n13689), .Z(c[1546]) );
  XNOR U16241 ( .A(a[1546]), .B(n13690), .Z(n13689) );
  IV U16242 ( .A(n13687), .Z(n13690) );
  XOR U16243 ( .A(n13691), .B(n13692), .Z(n13687) );
  ANDN U16244 ( .B(n13693), .A(n13694), .Z(n13691) );
  XNOR U16245 ( .A(b[1545]), .B(n13692), .Z(n13693) );
  XNOR U16246 ( .A(b[1545]), .B(n13694), .Z(c[1545]) );
  XNOR U16247 ( .A(a[1545]), .B(n13695), .Z(n13694) );
  IV U16248 ( .A(n13692), .Z(n13695) );
  XOR U16249 ( .A(n13696), .B(n13697), .Z(n13692) );
  ANDN U16250 ( .B(n13698), .A(n13699), .Z(n13696) );
  XNOR U16251 ( .A(b[1544]), .B(n13697), .Z(n13698) );
  XNOR U16252 ( .A(b[1544]), .B(n13699), .Z(c[1544]) );
  XNOR U16253 ( .A(a[1544]), .B(n13700), .Z(n13699) );
  IV U16254 ( .A(n13697), .Z(n13700) );
  XOR U16255 ( .A(n13701), .B(n13702), .Z(n13697) );
  ANDN U16256 ( .B(n13703), .A(n13704), .Z(n13701) );
  XNOR U16257 ( .A(b[1543]), .B(n13702), .Z(n13703) );
  XNOR U16258 ( .A(b[1543]), .B(n13704), .Z(c[1543]) );
  XNOR U16259 ( .A(a[1543]), .B(n13705), .Z(n13704) );
  IV U16260 ( .A(n13702), .Z(n13705) );
  XOR U16261 ( .A(n13706), .B(n13707), .Z(n13702) );
  ANDN U16262 ( .B(n13708), .A(n13709), .Z(n13706) );
  XNOR U16263 ( .A(b[1542]), .B(n13707), .Z(n13708) );
  XNOR U16264 ( .A(b[1542]), .B(n13709), .Z(c[1542]) );
  XNOR U16265 ( .A(a[1542]), .B(n13710), .Z(n13709) );
  IV U16266 ( .A(n13707), .Z(n13710) );
  XOR U16267 ( .A(n13711), .B(n13712), .Z(n13707) );
  ANDN U16268 ( .B(n13713), .A(n13714), .Z(n13711) );
  XNOR U16269 ( .A(b[1541]), .B(n13712), .Z(n13713) );
  XNOR U16270 ( .A(b[1541]), .B(n13714), .Z(c[1541]) );
  XNOR U16271 ( .A(a[1541]), .B(n13715), .Z(n13714) );
  IV U16272 ( .A(n13712), .Z(n13715) );
  XOR U16273 ( .A(n13716), .B(n13717), .Z(n13712) );
  ANDN U16274 ( .B(n13718), .A(n13719), .Z(n13716) );
  XNOR U16275 ( .A(b[1540]), .B(n13717), .Z(n13718) );
  XNOR U16276 ( .A(b[1540]), .B(n13719), .Z(c[1540]) );
  XNOR U16277 ( .A(a[1540]), .B(n13720), .Z(n13719) );
  IV U16278 ( .A(n13717), .Z(n13720) );
  XOR U16279 ( .A(n13721), .B(n13722), .Z(n13717) );
  ANDN U16280 ( .B(n13723), .A(n13724), .Z(n13721) );
  XNOR U16281 ( .A(b[1539]), .B(n13722), .Z(n13723) );
  XNOR U16282 ( .A(b[153]), .B(n13725), .Z(c[153]) );
  XNOR U16283 ( .A(b[1539]), .B(n13724), .Z(c[1539]) );
  XNOR U16284 ( .A(a[1539]), .B(n13726), .Z(n13724) );
  IV U16285 ( .A(n13722), .Z(n13726) );
  XOR U16286 ( .A(n13727), .B(n13728), .Z(n13722) );
  ANDN U16287 ( .B(n13729), .A(n13730), .Z(n13727) );
  XNOR U16288 ( .A(b[1538]), .B(n13728), .Z(n13729) );
  XNOR U16289 ( .A(b[1538]), .B(n13730), .Z(c[1538]) );
  XNOR U16290 ( .A(a[1538]), .B(n13731), .Z(n13730) );
  IV U16291 ( .A(n13728), .Z(n13731) );
  XOR U16292 ( .A(n13732), .B(n13733), .Z(n13728) );
  ANDN U16293 ( .B(n13734), .A(n13735), .Z(n13732) );
  XNOR U16294 ( .A(b[1537]), .B(n13733), .Z(n13734) );
  XNOR U16295 ( .A(b[1537]), .B(n13735), .Z(c[1537]) );
  XNOR U16296 ( .A(a[1537]), .B(n13736), .Z(n13735) );
  IV U16297 ( .A(n13733), .Z(n13736) );
  XOR U16298 ( .A(n13737), .B(n13738), .Z(n13733) );
  ANDN U16299 ( .B(n13739), .A(n13740), .Z(n13737) );
  XNOR U16300 ( .A(b[1536]), .B(n13738), .Z(n13739) );
  XNOR U16301 ( .A(b[1536]), .B(n13740), .Z(c[1536]) );
  XNOR U16302 ( .A(a[1536]), .B(n13741), .Z(n13740) );
  IV U16303 ( .A(n13738), .Z(n13741) );
  XOR U16304 ( .A(n13742), .B(n13743), .Z(n13738) );
  ANDN U16305 ( .B(n13744), .A(n13745), .Z(n13742) );
  XNOR U16306 ( .A(b[1535]), .B(n13743), .Z(n13744) );
  XNOR U16307 ( .A(b[1535]), .B(n13745), .Z(c[1535]) );
  XNOR U16308 ( .A(a[1535]), .B(n13746), .Z(n13745) );
  IV U16309 ( .A(n13743), .Z(n13746) );
  XOR U16310 ( .A(n13747), .B(n13748), .Z(n13743) );
  ANDN U16311 ( .B(n13749), .A(n13750), .Z(n13747) );
  XNOR U16312 ( .A(b[1534]), .B(n13748), .Z(n13749) );
  XNOR U16313 ( .A(b[1534]), .B(n13750), .Z(c[1534]) );
  XNOR U16314 ( .A(a[1534]), .B(n13751), .Z(n13750) );
  IV U16315 ( .A(n13748), .Z(n13751) );
  XOR U16316 ( .A(n13752), .B(n13753), .Z(n13748) );
  ANDN U16317 ( .B(n13754), .A(n13755), .Z(n13752) );
  XNOR U16318 ( .A(b[1533]), .B(n13753), .Z(n13754) );
  XNOR U16319 ( .A(b[1533]), .B(n13755), .Z(c[1533]) );
  XNOR U16320 ( .A(a[1533]), .B(n13756), .Z(n13755) );
  IV U16321 ( .A(n13753), .Z(n13756) );
  XOR U16322 ( .A(n13757), .B(n13758), .Z(n13753) );
  ANDN U16323 ( .B(n13759), .A(n13760), .Z(n13757) );
  XNOR U16324 ( .A(b[1532]), .B(n13758), .Z(n13759) );
  XNOR U16325 ( .A(b[1532]), .B(n13760), .Z(c[1532]) );
  XNOR U16326 ( .A(a[1532]), .B(n13761), .Z(n13760) );
  IV U16327 ( .A(n13758), .Z(n13761) );
  XOR U16328 ( .A(n13762), .B(n13763), .Z(n13758) );
  ANDN U16329 ( .B(n13764), .A(n13765), .Z(n13762) );
  XNOR U16330 ( .A(b[1531]), .B(n13763), .Z(n13764) );
  XNOR U16331 ( .A(b[1531]), .B(n13765), .Z(c[1531]) );
  XNOR U16332 ( .A(a[1531]), .B(n13766), .Z(n13765) );
  IV U16333 ( .A(n13763), .Z(n13766) );
  XOR U16334 ( .A(n13767), .B(n13768), .Z(n13763) );
  ANDN U16335 ( .B(n13769), .A(n13770), .Z(n13767) );
  XNOR U16336 ( .A(b[1530]), .B(n13768), .Z(n13769) );
  XNOR U16337 ( .A(b[1530]), .B(n13770), .Z(c[1530]) );
  XNOR U16338 ( .A(a[1530]), .B(n13771), .Z(n13770) );
  IV U16339 ( .A(n13768), .Z(n13771) );
  XOR U16340 ( .A(n13772), .B(n13773), .Z(n13768) );
  ANDN U16341 ( .B(n13774), .A(n13775), .Z(n13772) );
  XNOR U16342 ( .A(b[1529]), .B(n13773), .Z(n13774) );
  XNOR U16343 ( .A(b[152]), .B(n13776), .Z(c[152]) );
  XNOR U16344 ( .A(b[1529]), .B(n13775), .Z(c[1529]) );
  XNOR U16345 ( .A(a[1529]), .B(n13777), .Z(n13775) );
  IV U16346 ( .A(n13773), .Z(n13777) );
  XOR U16347 ( .A(n13778), .B(n13779), .Z(n13773) );
  ANDN U16348 ( .B(n13780), .A(n13781), .Z(n13778) );
  XNOR U16349 ( .A(b[1528]), .B(n13779), .Z(n13780) );
  XNOR U16350 ( .A(b[1528]), .B(n13781), .Z(c[1528]) );
  XNOR U16351 ( .A(a[1528]), .B(n13782), .Z(n13781) );
  IV U16352 ( .A(n13779), .Z(n13782) );
  XOR U16353 ( .A(n13783), .B(n13784), .Z(n13779) );
  ANDN U16354 ( .B(n13785), .A(n13786), .Z(n13783) );
  XNOR U16355 ( .A(b[1527]), .B(n13784), .Z(n13785) );
  XNOR U16356 ( .A(b[1527]), .B(n13786), .Z(c[1527]) );
  XNOR U16357 ( .A(a[1527]), .B(n13787), .Z(n13786) );
  IV U16358 ( .A(n13784), .Z(n13787) );
  XOR U16359 ( .A(n13788), .B(n13789), .Z(n13784) );
  ANDN U16360 ( .B(n13790), .A(n13791), .Z(n13788) );
  XNOR U16361 ( .A(b[1526]), .B(n13789), .Z(n13790) );
  XNOR U16362 ( .A(b[1526]), .B(n13791), .Z(c[1526]) );
  XNOR U16363 ( .A(a[1526]), .B(n13792), .Z(n13791) );
  IV U16364 ( .A(n13789), .Z(n13792) );
  XOR U16365 ( .A(n13793), .B(n13794), .Z(n13789) );
  ANDN U16366 ( .B(n13795), .A(n13796), .Z(n13793) );
  XNOR U16367 ( .A(b[1525]), .B(n13794), .Z(n13795) );
  XNOR U16368 ( .A(b[1525]), .B(n13796), .Z(c[1525]) );
  XNOR U16369 ( .A(a[1525]), .B(n13797), .Z(n13796) );
  IV U16370 ( .A(n13794), .Z(n13797) );
  XOR U16371 ( .A(n13798), .B(n13799), .Z(n13794) );
  ANDN U16372 ( .B(n13800), .A(n13801), .Z(n13798) );
  XNOR U16373 ( .A(b[1524]), .B(n13799), .Z(n13800) );
  XNOR U16374 ( .A(b[1524]), .B(n13801), .Z(c[1524]) );
  XNOR U16375 ( .A(a[1524]), .B(n13802), .Z(n13801) );
  IV U16376 ( .A(n13799), .Z(n13802) );
  XOR U16377 ( .A(n13803), .B(n13804), .Z(n13799) );
  ANDN U16378 ( .B(n13805), .A(n13806), .Z(n13803) );
  XNOR U16379 ( .A(b[1523]), .B(n13804), .Z(n13805) );
  XNOR U16380 ( .A(b[1523]), .B(n13806), .Z(c[1523]) );
  XNOR U16381 ( .A(a[1523]), .B(n13807), .Z(n13806) );
  IV U16382 ( .A(n13804), .Z(n13807) );
  XOR U16383 ( .A(n13808), .B(n13809), .Z(n13804) );
  ANDN U16384 ( .B(n13810), .A(n13811), .Z(n13808) );
  XNOR U16385 ( .A(b[1522]), .B(n13809), .Z(n13810) );
  XNOR U16386 ( .A(b[1522]), .B(n13811), .Z(c[1522]) );
  XNOR U16387 ( .A(a[1522]), .B(n13812), .Z(n13811) );
  IV U16388 ( .A(n13809), .Z(n13812) );
  XOR U16389 ( .A(n13813), .B(n13814), .Z(n13809) );
  ANDN U16390 ( .B(n13815), .A(n13816), .Z(n13813) );
  XNOR U16391 ( .A(b[1521]), .B(n13814), .Z(n13815) );
  XNOR U16392 ( .A(b[1521]), .B(n13816), .Z(c[1521]) );
  XNOR U16393 ( .A(a[1521]), .B(n13817), .Z(n13816) );
  IV U16394 ( .A(n13814), .Z(n13817) );
  XOR U16395 ( .A(n13818), .B(n13819), .Z(n13814) );
  ANDN U16396 ( .B(n13820), .A(n13821), .Z(n13818) );
  XNOR U16397 ( .A(b[1520]), .B(n13819), .Z(n13820) );
  XNOR U16398 ( .A(b[1520]), .B(n13821), .Z(c[1520]) );
  XNOR U16399 ( .A(a[1520]), .B(n13822), .Z(n13821) );
  IV U16400 ( .A(n13819), .Z(n13822) );
  XOR U16401 ( .A(n13823), .B(n13824), .Z(n13819) );
  ANDN U16402 ( .B(n13825), .A(n13826), .Z(n13823) );
  XNOR U16403 ( .A(b[1519]), .B(n13824), .Z(n13825) );
  XNOR U16404 ( .A(b[151]), .B(n13827), .Z(c[151]) );
  XNOR U16405 ( .A(b[1519]), .B(n13826), .Z(c[1519]) );
  XNOR U16406 ( .A(a[1519]), .B(n13828), .Z(n13826) );
  IV U16407 ( .A(n13824), .Z(n13828) );
  XOR U16408 ( .A(n13829), .B(n13830), .Z(n13824) );
  ANDN U16409 ( .B(n13831), .A(n13832), .Z(n13829) );
  XNOR U16410 ( .A(b[1518]), .B(n13830), .Z(n13831) );
  XNOR U16411 ( .A(b[1518]), .B(n13832), .Z(c[1518]) );
  XNOR U16412 ( .A(a[1518]), .B(n13833), .Z(n13832) );
  IV U16413 ( .A(n13830), .Z(n13833) );
  XOR U16414 ( .A(n13834), .B(n13835), .Z(n13830) );
  ANDN U16415 ( .B(n13836), .A(n13837), .Z(n13834) );
  XNOR U16416 ( .A(b[1517]), .B(n13835), .Z(n13836) );
  XNOR U16417 ( .A(b[1517]), .B(n13837), .Z(c[1517]) );
  XNOR U16418 ( .A(a[1517]), .B(n13838), .Z(n13837) );
  IV U16419 ( .A(n13835), .Z(n13838) );
  XOR U16420 ( .A(n13839), .B(n13840), .Z(n13835) );
  ANDN U16421 ( .B(n13841), .A(n13842), .Z(n13839) );
  XNOR U16422 ( .A(b[1516]), .B(n13840), .Z(n13841) );
  XNOR U16423 ( .A(b[1516]), .B(n13842), .Z(c[1516]) );
  XNOR U16424 ( .A(a[1516]), .B(n13843), .Z(n13842) );
  IV U16425 ( .A(n13840), .Z(n13843) );
  XOR U16426 ( .A(n13844), .B(n13845), .Z(n13840) );
  ANDN U16427 ( .B(n13846), .A(n13847), .Z(n13844) );
  XNOR U16428 ( .A(b[1515]), .B(n13845), .Z(n13846) );
  XNOR U16429 ( .A(b[1515]), .B(n13847), .Z(c[1515]) );
  XNOR U16430 ( .A(a[1515]), .B(n13848), .Z(n13847) );
  IV U16431 ( .A(n13845), .Z(n13848) );
  XOR U16432 ( .A(n13849), .B(n13850), .Z(n13845) );
  ANDN U16433 ( .B(n13851), .A(n13852), .Z(n13849) );
  XNOR U16434 ( .A(b[1514]), .B(n13850), .Z(n13851) );
  XNOR U16435 ( .A(b[1514]), .B(n13852), .Z(c[1514]) );
  XNOR U16436 ( .A(a[1514]), .B(n13853), .Z(n13852) );
  IV U16437 ( .A(n13850), .Z(n13853) );
  XOR U16438 ( .A(n13854), .B(n13855), .Z(n13850) );
  ANDN U16439 ( .B(n13856), .A(n13857), .Z(n13854) );
  XNOR U16440 ( .A(b[1513]), .B(n13855), .Z(n13856) );
  XNOR U16441 ( .A(b[1513]), .B(n13857), .Z(c[1513]) );
  XNOR U16442 ( .A(a[1513]), .B(n13858), .Z(n13857) );
  IV U16443 ( .A(n13855), .Z(n13858) );
  XOR U16444 ( .A(n13859), .B(n13860), .Z(n13855) );
  ANDN U16445 ( .B(n13861), .A(n13862), .Z(n13859) );
  XNOR U16446 ( .A(b[1512]), .B(n13860), .Z(n13861) );
  XNOR U16447 ( .A(b[1512]), .B(n13862), .Z(c[1512]) );
  XNOR U16448 ( .A(a[1512]), .B(n13863), .Z(n13862) );
  IV U16449 ( .A(n13860), .Z(n13863) );
  XOR U16450 ( .A(n13864), .B(n13865), .Z(n13860) );
  ANDN U16451 ( .B(n13866), .A(n13867), .Z(n13864) );
  XNOR U16452 ( .A(b[1511]), .B(n13865), .Z(n13866) );
  XNOR U16453 ( .A(b[1511]), .B(n13867), .Z(c[1511]) );
  XNOR U16454 ( .A(a[1511]), .B(n13868), .Z(n13867) );
  IV U16455 ( .A(n13865), .Z(n13868) );
  XOR U16456 ( .A(n13869), .B(n13870), .Z(n13865) );
  ANDN U16457 ( .B(n13871), .A(n13872), .Z(n13869) );
  XNOR U16458 ( .A(b[1510]), .B(n13870), .Z(n13871) );
  XNOR U16459 ( .A(b[1510]), .B(n13872), .Z(c[1510]) );
  XNOR U16460 ( .A(a[1510]), .B(n13873), .Z(n13872) );
  IV U16461 ( .A(n13870), .Z(n13873) );
  XOR U16462 ( .A(n13874), .B(n13875), .Z(n13870) );
  ANDN U16463 ( .B(n13876), .A(n13877), .Z(n13874) );
  XNOR U16464 ( .A(b[1509]), .B(n13875), .Z(n13876) );
  XNOR U16465 ( .A(b[150]), .B(n13878), .Z(c[150]) );
  XNOR U16466 ( .A(b[1509]), .B(n13877), .Z(c[1509]) );
  XNOR U16467 ( .A(a[1509]), .B(n13879), .Z(n13877) );
  IV U16468 ( .A(n13875), .Z(n13879) );
  XOR U16469 ( .A(n13880), .B(n13881), .Z(n13875) );
  ANDN U16470 ( .B(n13882), .A(n13883), .Z(n13880) );
  XNOR U16471 ( .A(b[1508]), .B(n13881), .Z(n13882) );
  XNOR U16472 ( .A(b[1508]), .B(n13883), .Z(c[1508]) );
  XNOR U16473 ( .A(a[1508]), .B(n13884), .Z(n13883) );
  IV U16474 ( .A(n13881), .Z(n13884) );
  XOR U16475 ( .A(n13885), .B(n13886), .Z(n13881) );
  ANDN U16476 ( .B(n13887), .A(n13888), .Z(n13885) );
  XNOR U16477 ( .A(b[1507]), .B(n13886), .Z(n13887) );
  XNOR U16478 ( .A(b[1507]), .B(n13888), .Z(c[1507]) );
  XNOR U16479 ( .A(a[1507]), .B(n13889), .Z(n13888) );
  IV U16480 ( .A(n13886), .Z(n13889) );
  XOR U16481 ( .A(n13890), .B(n13891), .Z(n13886) );
  ANDN U16482 ( .B(n13892), .A(n13893), .Z(n13890) );
  XNOR U16483 ( .A(b[1506]), .B(n13891), .Z(n13892) );
  XNOR U16484 ( .A(b[1506]), .B(n13893), .Z(c[1506]) );
  XNOR U16485 ( .A(a[1506]), .B(n13894), .Z(n13893) );
  IV U16486 ( .A(n13891), .Z(n13894) );
  XOR U16487 ( .A(n13895), .B(n13896), .Z(n13891) );
  ANDN U16488 ( .B(n13897), .A(n13898), .Z(n13895) );
  XNOR U16489 ( .A(b[1505]), .B(n13896), .Z(n13897) );
  XNOR U16490 ( .A(b[1505]), .B(n13898), .Z(c[1505]) );
  XNOR U16491 ( .A(a[1505]), .B(n13899), .Z(n13898) );
  IV U16492 ( .A(n13896), .Z(n13899) );
  XOR U16493 ( .A(n13900), .B(n13901), .Z(n13896) );
  ANDN U16494 ( .B(n13902), .A(n13903), .Z(n13900) );
  XNOR U16495 ( .A(b[1504]), .B(n13901), .Z(n13902) );
  XNOR U16496 ( .A(b[1504]), .B(n13903), .Z(c[1504]) );
  XNOR U16497 ( .A(a[1504]), .B(n13904), .Z(n13903) );
  IV U16498 ( .A(n13901), .Z(n13904) );
  XOR U16499 ( .A(n13905), .B(n13906), .Z(n13901) );
  ANDN U16500 ( .B(n13907), .A(n13908), .Z(n13905) );
  XNOR U16501 ( .A(b[1503]), .B(n13906), .Z(n13907) );
  XNOR U16502 ( .A(b[1503]), .B(n13908), .Z(c[1503]) );
  XNOR U16503 ( .A(a[1503]), .B(n13909), .Z(n13908) );
  IV U16504 ( .A(n13906), .Z(n13909) );
  XOR U16505 ( .A(n13910), .B(n13911), .Z(n13906) );
  ANDN U16506 ( .B(n13912), .A(n13913), .Z(n13910) );
  XNOR U16507 ( .A(b[1502]), .B(n13911), .Z(n13912) );
  XNOR U16508 ( .A(b[1502]), .B(n13913), .Z(c[1502]) );
  XNOR U16509 ( .A(a[1502]), .B(n13914), .Z(n13913) );
  IV U16510 ( .A(n13911), .Z(n13914) );
  XOR U16511 ( .A(n13915), .B(n13916), .Z(n13911) );
  ANDN U16512 ( .B(n13917), .A(n13918), .Z(n13915) );
  XNOR U16513 ( .A(b[1501]), .B(n13916), .Z(n13917) );
  XNOR U16514 ( .A(b[1501]), .B(n13918), .Z(c[1501]) );
  XNOR U16515 ( .A(a[1501]), .B(n13919), .Z(n13918) );
  IV U16516 ( .A(n13916), .Z(n13919) );
  XOR U16517 ( .A(n13920), .B(n13921), .Z(n13916) );
  ANDN U16518 ( .B(n13922), .A(n13923), .Z(n13920) );
  XNOR U16519 ( .A(b[1500]), .B(n13921), .Z(n13922) );
  XNOR U16520 ( .A(b[1500]), .B(n13923), .Z(c[1500]) );
  XNOR U16521 ( .A(a[1500]), .B(n13924), .Z(n13923) );
  IV U16522 ( .A(n13921), .Z(n13924) );
  XOR U16523 ( .A(n13925), .B(n13926), .Z(n13921) );
  ANDN U16524 ( .B(n13927), .A(n13928), .Z(n13925) );
  XNOR U16525 ( .A(b[1499]), .B(n13926), .Z(n13927) );
  XNOR U16526 ( .A(b[14]), .B(n13929), .Z(c[14]) );
  XNOR U16527 ( .A(b[149]), .B(n13930), .Z(c[149]) );
  XNOR U16528 ( .A(b[1499]), .B(n13928), .Z(c[1499]) );
  XNOR U16529 ( .A(a[1499]), .B(n13931), .Z(n13928) );
  IV U16530 ( .A(n13926), .Z(n13931) );
  XOR U16531 ( .A(n13932), .B(n13933), .Z(n13926) );
  ANDN U16532 ( .B(n13934), .A(n13935), .Z(n13932) );
  XNOR U16533 ( .A(b[1498]), .B(n13933), .Z(n13934) );
  XNOR U16534 ( .A(b[1498]), .B(n13935), .Z(c[1498]) );
  XNOR U16535 ( .A(a[1498]), .B(n13936), .Z(n13935) );
  IV U16536 ( .A(n13933), .Z(n13936) );
  XOR U16537 ( .A(n13937), .B(n13938), .Z(n13933) );
  ANDN U16538 ( .B(n13939), .A(n13940), .Z(n13937) );
  XNOR U16539 ( .A(b[1497]), .B(n13938), .Z(n13939) );
  XNOR U16540 ( .A(b[1497]), .B(n13940), .Z(c[1497]) );
  XNOR U16541 ( .A(a[1497]), .B(n13941), .Z(n13940) );
  IV U16542 ( .A(n13938), .Z(n13941) );
  XOR U16543 ( .A(n13942), .B(n13943), .Z(n13938) );
  ANDN U16544 ( .B(n13944), .A(n13945), .Z(n13942) );
  XNOR U16545 ( .A(b[1496]), .B(n13943), .Z(n13944) );
  XNOR U16546 ( .A(b[1496]), .B(n13945), .Z(c[1496]) );
  XNOR U16547 ( .A(a[1496]), .B(n13946), .Z(n13945) );
  IV U16548 ( .A(n13943), .Z(n13946) );
  XOR U16549 ( .A(n13947), .B(n13948), .Z(n13943) );
  ANDN U16550 ( .B(n13949), .A(n13950), .Z(n13947) );
  XNOR U16551 ( .A(b[1495]), .B(n13948), .Z(n13949) );
  XNOR U16552 ( .A(b[1495]), .B(n13950), .Z(c[1495]) );
  XNOR U16553 ( .A(a[1495]), .B(n13951), .Z(n13950) );
  IV U16554 ( .A(n13948), .Z(n13951) );
  XOR U16555 ( .A(n13952), .B(n13953), .Z(n13948) );
  ANDN U16556 ( .B(n13954), .A(n13955), .Z(n13952) );
  XNOR U16557 ( .A(b[1494]), .B(n13953), .Z(n13954) );
  XNOR U16558 ( .A(b[1494]), .B(n13955), .Z(c[1494]) );
  XNOR U16559 ( .A(a[1494]), .B(n13956), .Z(n13955) );
  IV U16560 ( .A(n13953), .Z(n13956) );
  XOR U16561 ( .A(n13957), .B(n13958), .Z(n13953) );
  ANDN U16562 ( .B(n13959), .A(n13960), .Z(n13957) );
  XNOR U16563 ( .A(b[1493]), .B(n13958), .Z(n13959) );
  XNOR U16564 ( .A(b[1493]), .B(n13960), .Z(c[1493]) );
  XNOR U16565 ( .A(a[1493]), .B(n13961), .Z(n13960) );
  IV U16566 ( .A(n13958), .Z(n13961) );
  XOR U16567 ( .A(n13962), .B(n13963), .Z(n13958) );
  ANDN U16568 ( .B(n13964), .A(n13965), .Z(n13962) );
  XNOR U16569 ( .A(b[1492]), .B(n13963), .Z(n13964) );
  XNOR U16570 ( .A(b[1492]), .B(n13965), .Z(c[1492]) );
  XNOR U16571 ( .A(a[1492]), .B(n13966), .Z(n13965) );
  IV U16572 ( .A(n13963), .Z(n13966) );
  XOR U16573 ( .A(n13967), .B(n13968), .Z(n13963) );
  ANDN U16574 ( .B(n13969), .A(n13970), .Z(n13967) );
  XNOR U16575 ( .A(b[1491]), .B(n13968), .Z(n13969) );
  XNOR U16576 ( .A(b[1491]), .B(n13970), .Z(c[1491]) );
  XNOR U16577 ( .A(a[1491]), .B(n13971), .Z(n13970) );
  IV U16578 ( .A(n13968), .Z(n13971) );
  XOR U16579 ( .A(n13972), .B(n13973), .Z(n13968) );
  ANDN U16580 ( .B(n13974), .A(n13975), .Z(n13972) );
  XNOR U16581 ( .A(b[1490]), .B(n13973), .Z(n13974) );
  XNOR U16582 ( .A(b[1490]), .B(n13975), .Z(c[1490]) );
  XNOR U16583 ( .A(a[1490]), .B(n13976), .Z(n13975) );
  IV U16584 ( .A(n13973), .Z(n13976) );
  XOR U16585 ( .A(n13977), .B(n13978), .Z(n13973) );
  ANDN U16586 ( .B(n13979), .A(n13980), .Z(n13977) );
  XNOR U16587 ( .A(b[1489]), .B(n13978), .Z(n13979) );
  XNOR U16588 ( .A(b[148]), .B(n13981), .Z(c[148]) );
  XNOR U16589 ( .A(b[1489]), .B(n13980), .Z(c[1489]) );
  XNOR U16590 ( .A(a[1489]), .B(n13982), .Z(n13980) );
  IV U16591 ( .A(n13978), .Z(n13982) );
  XOR U16592 ( .A(n13983), .B(n13984), .Z(n13978) );
  ANDN U16593 ( .B(n13985), .A(n13986), .Z(n13983) );
  XNOR U16594 ( .A(b[1488]), .B(n13984), .Z(n13985) );
  XNOR U16595 ( .A(b[1488]), .B(n13986), .Z(c[1488]) );
  XNOR U16596 ( .A(a[1488]), .B(n13987), .Z(n13986) );
  IV U16597 ( .A(n13984), .Z(n13987) );
  XOR U16598 ( .A(n13988), .B(n13989), .Z(n13984) );
  ANDN U16599 ( .B(n13990), .A(n13991), .Z(n13988) );
  XNOR U16600 ( .A(b[1487]), .B(n13989), .Z(n13990) );
  XNOR U16601 ( .A(b[1487]), .B(n13991), .Z(c[1487]) );
  XNOR U16602 ( .A(a[1487]), .B(n13992), .Z(n13991) );
  IV U16603 ( .A(n13989), .Z(n13992) );
  XOR U16604 ( .A(n13993), .B(n13994), .Z(n13989) );
  ANDN U16605 ( .B(n13995), .A(n13996), .Z(n13993) );
  XNOR U16606 ( .A(b[1486]), .B(n13994), .Z(n13995) );
  XNOR U16607 ( .A(b[1486]), .B(n13996), .Z(c[1486]) );
  XNOR U16608 ( .A(a[1486]), .B(n13997), .Z(n13996) );
  IV U16609 ( .A(n13994), .Z(n13997) );
  XOR U16610 ( .A(n13998), .B(n13999), .Z(n13994) );
  ANDN U16611 ( .B(n14000), .A(n14001), .Z(n13998) );
  XNOR U16612 ( .A(b[1485]), .B(n13999), .Z(n14000) );
  XNOR U16613 ( .A(b[1485]), .B(n14001), .Z(c[1485]) );
  XNOR U16614 ( .A(a[1485]), .B(n14002), .Z(n14001) );
  IV U16615 ( .A(n13999), .Z(n14002) );
  XOR U16616 ( .A(n14003), .B(n14004), .Z(n13999) );
  ANDN U16617 ( .B(n14005), .A(n14006), .Z(n14003) );
  XNOR U16618 ( .A(b[1484]), .B(n14004), .Z(n14005) );
  XNOR U16619 ( .A(b[1484]), .B(n14006), .Z(c[1484]) );
  XNOR U16620 ( .A(a[1484]), .B(n14007), .Z(n14006) );
  IV U16621 ( .A(n14004), .Z(n14007) );
  XOR U16622 ( .A(n14008), .B(n14009), .Z(n14004) );
  ANDN U16623 ( .B(n14010), .A(n14011), .Z(n14008) );
  XNOR U16624 ( .A(b[1483]), .B(n14009), .Z(n14010) );
  XNOR U16625 ( .A(b[1483]), .B(n14011), .Z(c[1483]) );
  XNOR U16626 ( .A(a[1483]), .B(n14012), .Z(n14011) );
  IV U16627 ( .A(n14009), .Z(n14012) );
  XOR U16628 ( .A(n14013), .B(n14014), .Z(n14009) );
  ANDN U16629 ( .B(n14015), .A(n14016), .Z(n14013) );
  XNOR U16630 ( .A(b[1482]), .B(n14014), .Z(n14015) );
  XNOR U16631 ( .A(b[1482]), .B(n14016), .Z(c[1482]) );
  XNOR U16632 ( .A(a[1482]), .B(n14017), .Z(n14016) );
  IV U16633 ( .A(n14014), .Z(n14017) );
  XOR U16634 ( .A(n14018), .B(n14019), .Z(n14014) );
  ANDN U16635 ( .B(n14020), .A(n14021), .Z(n14018) );
  XNOR U16636 ( .A(b[1481]), .B(n14019), .Z(n14020) );
  XNOR U16637 ( .A(b[1481]), .B(n14021), .Z(c[1481]) );
  XNOR U16638 ( .A(a[1481]), .B(n14022), .Z(n14021) );
  IV U16639 ( .A(n14019), .Z(n14022) );
  XOR U16640 ( .A(n14023), .B(n14024), .Z(n14019) );
  ANDN U16641 ( .B(n14025), .A(n14026), .Z(n14023) );
  XNOR U16642 ( .A(b[1480]), .B(n14024), .Z(n14025) );
  XNOR U16643 ( .A(b[1480]), .B(n14026), .Z(c[1480]) );
  XNOR U16644 ( .A(a[1480]), .B(n14027), .Z(n14026) );
  IV U16645 ( .A(n14024), .Z(n14027) );
  XOR U16646 ( .A(n14028), .B(n14029), .Z(n14024) );
  ANDN U16647 ( .B(n14030), .A(n14031), .Z(n14028) );
  XNOR U16648 ( .A(b[1479]), .B(n14029), .Z(n14030) );
  XNOR U16649 ( .A(b[147]), .B(n14032), .Z(c[147]) );
  XNOR U16650 ( .A(b[1479]), .B(n14031), .Z(c[1479]) );
  XNOR U16651 ( .A(a[1479]), .B(n14033), .Z(n14031) );
  IV U16652 ( .A(n14029), .Z(n14033) );
  XOR U16653 ( .A(n14034), .B(n14035), .Z(n14029) );
  ANDN U16654 ( .B(n14036), .A(n14037), .Z(n14034) );
  XNOR U16655 ( .A(b[1478]), .B(n14035), .Z(n14036) );
  XNOR U16656 ( .A(b[1478]), .B(n14037), .Z(c[1478]) );
  XNOR U16657 ( .A(a[1478]), .B(n14038), .Z(n14037) );
  IV U16658 ( .A(n14035), .Z(n14038) );
  XOR U16659 ( .A(n14039), .B(n14040), .Z(n14035) );
  ANDN U16660 ( .B(n14041), .A(n14042), .Z(n14039) );
  XNOR U16661 ( .A(b[1477]), .B(n14040), .Z(n14041) );
  XNOR U16662 ( .A(b[1477]), .B(n14042), .Z(c[1477]) );
  XNOR U16663 ( .A(a[1477]), .B(n14043), .Z(n14042) );
  IV U16664 ( .A(n14040), .Z(n14043) );
  XOR U16665 ( .A(n14044), .B(n14045), .Z(n14040) );
  ANDN U16666 ( .B(n14046), .A(n14047), .Z(n14044) );
  XNOR U16667 ( .A(b[1476]), .B(n14045), .Z(n14046) );
  XNOR U16668 ( .A(b[1476]), .B(n14047), .Z(c[1476]) );
  XNOR U16669 ( .A(a[1476]), .B(n14048), .Z(n14047) );
  IV U16670 ( .A(n14045), .Z(n14048) );
  XOR U16671 ( .A(n14049), .B(n14050), .Z(n14045) );
  ANDN U16672 ( .B(n14051), .A(n14052), .Z(n14049) );
  XNOR U16673 ( .A(b[1475]), .B(n14050), .Z(n14051) );
  XNOR U16674 ( .A(b[1475]), .B(n14052), .Z(c[1475]) );
  XNOR U16675 ( .A(a[1475]), .B(n14053), .Z(n14052) );
  IV U16676 ( .A(n14050), .Z(n14053) );
  XOR U16677 ( .A(n14054), .B(n14055), .Z(n14050) );
  ANDN U16678 ( .B(n14056), .A(n14057), .Z(n14054) );
  XNOR U16679 ( .A(b[1474]), .B(n14055), .Z(n14056) );
  XNOR U16680 ( .A(b[1474]), .B(n14057), .Z(c[1474]) );
  XNOR U16681 ( .A(a[1474]), .B(n14058), .Z(n14057) );
  IV U16682 ( .A(n14055), .Z(n14058) );
  XOR U16683 ( .A(n14059), .B(n14060), .Z(n14055) );
  ANDN U16684 ( .B(n14061), .A(n14062), .Z(n14059) );
  XNOR U16685 ( .A(b[1473]), .B(n14060), .Z(n14061) );
  XNOR U16686 ( .A(b[1473]), .B(n14062), .Z(c[1473]) );
  XNOR U16687 ( .A(a[1473]), .B(n14063), .Z(n14062) );
  IV U16688 ( .A(n14060), .Z(n14063) );
  XOR U16689 ( .A(n14064), .B(n14065), .Z(n14060) );
  ANDN U16690 ( .B(n14066), .A(n14067), .Z(n14064) );
  XNOR U16691 ( .A(b[1472]), .B(n14065), .Z(n14066) );
  XNOR U16692 ( .A(b[1472]), .B(n14067), .Z(c[1472]) );
  XNOR U16693 ( .A(a[1472]), .B(n14068), .Z(n14067) );
  IV U16694 ( .A(n14065), .Z(n14068) );
  XOR U16695 ( .A(n14069), .B(n14070), .Z(n14065) );
  ANDN U16696 ( .B(n14071), .A(n14072), .Z(n14069) );
  XNOR U16697 ( .A(b[1471]), .B(n14070), .Z(n14071) );
  XNOR U16698 ( .A(b[1471]), .B(n14072), .Z(c[1471]) );
  XNOR U16699 ( .A(a[1471]), .B(n14073), .Z(n14072) );
  IV U16700 ( .A(n14070), .Z(n14073) );
  XOR U16701 ( .A(n14074), .B(n14075), .Z(n14070) );
  ANDN U16702 ( .B(n14076), .A(n14077), .Z(n14074) );
  XNOR U16703 ( .A(b[1470]), .B(n14075), .Z(n14076) );
  XNOR U16704 ( .A(b[1470]), .B(n14077), .Z(c[1470]) );
  XNOR U16705 ( .A(a[1470]), .B(n14078), .Z(n14077) );
  IV U16706 ( .A(n14075), .Z(n14078) );
  XOR U16707 ( .A(n14079), .B(n14080), .Z(n14075) );
  ANDN U16708 ( .B(n14081), .A(n14082), .Z(n14079) );
  XNOR U16709 ( .A(b[1469]), .B(n14080), .Z(n14081) );
  XNOR U16710 ( .A(b[146]), .B(n14083), .Z(c[146]) );
  XNOR U16711 ( .A(b[1469]), .B(n14082), .Z(c[1469]) );
  XNOR U16712 ( .A(a[1469]), .B(n14084), .Z(n14082) );
  IV U16713 ( .A(n14080), .Z(n14084) );
  XOR U16714 ( .A(n14085), .B(n14086), .Z(n14080) );
  ANDN U16715 ( .B(n14087), .A(n14088), .Z(n14085) );
  XNOR U16716 ( .A(b[1468]), .B(n14086), .Z(n14087) );
  XNOR U16717 ( .A(b[1468]), .B(n14088), .Z(c[1468]) );
  XNOR U16718 ( .A(a[1468]), .B(n14089), .Z(n14088) );
  IV U16719 ( .A(n14086), .Z(n14089) );
  XOR U16720 ( .A(n14090), .B(n14091), .Z(n14086) );
  ANDN U16721 ( .B(n14092), .A(n14093), .Z(n14090) );
  XNOR U16722 ( .A(b[1467]), .B(n14091), .Z(n14092) );
  XNOR U16723 ( .A(b[1467]), .B(n14093), .Z(c[1467]) );
  XNOR U16724 ( .A(a[1467]), .B(n14094), .Z(n14093) );
  IV U16725 ( .A(n14091), .Z(n14094) );
  XOR U16726 ( .A(n14095), .B(n14096), .Z(n14091) );
  ANDN U16727 ( .B(n14097), .A(n14098), .Z(n14095) );
  XNOR U16728 ( .A(b[1466]), .B(n14096), .Z(n14097) );
  XNOR U16729 ( .A(b[1466]), .B(n14098), .Z(c[1466]) );
  XNOR U16730 ( .A(a[1466]), .B(n14099), .Z(n14098) );
  IV U16731 ( .A(n14096), .Z(n14099) );
  XOR U16732 ( .A(n14100), .B(n14101), .Z(n14096) );
  ANDN U16733 ( .B(n14102), .A(n14103), .Z(n14100) );
  XNOR U16734 ( .A(b[1465]), .B(n14101), .Z(n14102) );
  XNOR U16735 ( .A(b[1465]), .B(n14103), .Z(c[1465]) );
  XNOR U16736 ( .A(a[1465]), .B(n14104), .Z(n14103) );
  IV U16737 ( .A(n14101), .Z(n14104) );
  XOR U16738 ( .A(n14105), .B(n14106), .Z(n14101) );
  ANDN U16739 ( .B(n14107), .A(n14108), .Z(n14105) );
  XNOR U16740 ( .A(b[1464]), .B(n14106), .Z(n14107) );
  XNOR U16741 ( .A(b[1464]), .B(n14108), .Z(c[1464]) );
  XNOR U16742 ( .A(a[1464]), .B(n14109), .Z(n14108) );
  IV U16743 ( .A(n14106), .Z(n14109) );
  XOR U16744 ( .A(n14110), .B(n14111), .Z(n14106) );
  ANDN U16745 ( .B(n14112), .A(n14113), .Z(n14110) );
  XNOR U16746 ( .A(b[1463]), .B(n14111), .Z(n14112) );
  XNOR U16747 ( .A(b[1463]), .B(n14113), .Z(c[1463]) );
  XNOR U16748 ( .A(a[1463]), .B(n14114), .Z(n14113) );
  IV U16749 ( .A(n14111), .Z(n14114) );
  XOR U16750 ( .A(n14115), .B(n14116), .Z(n14111) );
  ANDN U16751 ( .B(n14117), .A(n14118), .Z(n14115) );
  XNOR U16752 ( .A(b[1462]), .B(n14116), .Z(n14117) );
  XNOR U16753 ( .A(b[1462]), .B(n14118), .Z(c[1462]) );
  XNOR U16754 ( .A(a[1462]), .B(n14119), .Z(n14118) );
  IV U16755 ( .A(n14116), .Z(n14119) );
  XOR U16756 ( .A(n14120), .B(n14121), .Z(n14116) );
  ANDN U16757 ( .B(n14122), .A(n14123), .Z(n14120) );
  XNOR U16758 ( .A(b[1461]), .B(n14121), .Z(n14122) );
  XNOR U16759 ( .A(b[1461]), .B(n14123), .Z(c[1461]) );
  XNOR U16760 ( .A(a[1461]), .B(n14124), .Z(n14123) );
  IV U16761 ( .A(n14121), .Z(n14124) );
  XOR U16762 ( .A(n14125), .B(n14126), .Z(n14121) );
  ANDN U16763 ( .B(n14127), .A(n14128), .Z(n14125) );
  XNOR U16764 ( .A(b[1460]), .B(n14126), .Z(n14127) );
  XNOR U16765 ( .A(b[1460]), .B(n14128), .Z(c[1460]) );
  XNOR U16766 ( .A(a[1460]), .B(n14129), .Z(n14128) );
  IV U16767 ( .A(n14126), .Z(n14129) );
  XOR U16768 ( .A(n14130), .B(n14131), .Z(n14126) );
  ANDN U16769 ( .B(n14132), .A(n14133), .Z(n14130) );
  XNOR U16770 ( .A(b[1459]), .B(n14131), .Z(n14132) );
  XNOR U16771 ( .A(b[145]), .B(n14134), .Z(c[145]) );
  XNOR U16772 ( .A(b[1459]), .B(n14133), .Z(c[1459]) );
  XNOR U16773 ( .A(a[1459]), .B(n14135), .Z(n14133) );
  IV U16774 ( .A(n14131), .Z(n14135) );
  XOR U16775 ( .A(n14136), .B(n14137), .Z(n14131) );
  ANDN U16776 ( .B(n14138), .A(n14139), .Z(n14136) );
  XNOR U16777 ( .A(b[1458]), .B(n14137), .Z(n14138) );
  XNOR U16778 ( .A(b[1458]), .B(n14139), .Z(c[1458]) );
  XNOR U16779 ( .A(a[1458]), .B(n14140), .Z(n14139) );
  IV U16780 ( .A(n14137), .Z(n14140) );
  XOR U16781 ( .A(n14141), .B(n14142), .Z(n14137) );
  ANDN U16782 ( .B(n14143), .A(n14144), .Z(n14141) );
  XNOR U16783 ( .A(b[1457]), .B(n14142), .Z(n14143) );
  XNOR U16784 ( .A(b[1457]), .B(n14144), .Z(c[1457]) );
  XNOR U16785 ( .A(a[1457]), .B(n14145), .Z(n14144) );
  IV U16786 ( .A(n14142), .Z(n14145) );
  XOR U16787 ( .A(n14146), .B(n14147), .Z(n14142) );
  ANDN U16788 ( .B(n14148), .A(n14149), .Z(n14146) );
  XNOR U16789 ( .A(b[1456]), .B(n14147), .Z(n14148) );
  XNOR U16790 ( .A(b[1456]), .B(n14149), .Z(c[1456]) );
  XNOR U16791 ( .A(a[1456]), .B(n14150), .Z(n14149) );
  IV U16792 ( .A(n14147), .Z(n14150) );
  XOR U16793 ( .A(n14151), .B(n14152), .Z(n14147) );
  ANDN U16794 ( .B(n14153), .A(n14154), .Z(n14151) );
  XNOR U16795 ( .A(b[1455]), .B(n14152), .Z(n14153) );
  XNOR U16796 ( .A(b[1455]), .B(n14154), .Z(c[1455]) );
  XNOR U16797 ( .A(a[1455]), .B(n14155), .Z(n14154) );
  IV U16798 ( .A(n14152), .Z(n14155) );
  XOR U16799 ( .A(n14156), .B(n14157), .Z(n14152) );
  ANDN U16800 ( .B(n14158), .A(n14159), .Z(n14156) );
  XNOR U16801 ( .A(b[1454]), .B(n14157), .Z(n14158) );
  XNOR U16802 ( .A(b[1454]), .B(n14159), .Z(c[1454]) );
  XNOR U16803 ( .A(a[1454]), .B(n14160), .Z(n14159) );
  IV U16804 ( .A(n14157), .Z(n14160) );
  XOR U16805 ( .A(n14161), .B(n14162), .Z(n14157) );
  ANDN U16806 ( .B(n14163), .A(n14164), .Z(n14161) );
  XNOR U16807 ( .A(b[1453]), .B(n14162), .Z(n14163) );
  XNOR U16808 ( .A(b[1453]), .B(n14164), .Z(c[1453]) );
  XNOR U16809 ( .A(a[1453]), .B(n14165), .Z(n14164) );
  IV U16810 ( .A(n14162), .Z(n14165) );
  XOR U16811 ( .A(n14166), .B(n14167), .Z(n14162) );
  ANDN U16812 ( .B(n14168), .A(n14169), .Z(n14166) );
  XNOR U16813 ( .A(b[1452]), .B(n14167), .Z(n14168) );
  XNOR U16814 ( .A(b[1452]), .B(n14169), .Z(c[1452]) );
  XNOR U16815 ( .A(a[1452]), .B(n14170), .Z(n14169) );
  IV U16816 ( .A(n14167), .Z(n14170) );
  XOR U16817 ( .A(n14171), .B(n14172), .Z(n14167) );
  ANDN U16818 ( .B(n14173), .A(n14174), .Z(n14171) );
  XNOR U16819 ( .A(b[1451]), .B(n14172), .Z(n14173) );
  XNOR U16820 ( .A(b[1451]), .B(n14174), .Z(c[1451]) );
  XNOR U16821 ( .A(a[1451]), .B(n14175), .Z(n14174) );
  IV U16822 ( .A(n14172), .Z(n14175) );
  XOR U16823 ( .A(n14176), .B(n14177), .Z(n14172) );
  ANDN U16824 ( .B(n14178), .A(n14179), .Z(n14176) );
  XNOR U16825 ( .A(b[1450]), .B(n14177), .Z(n14178) );
  XNOR U16826 ( .A(b[1450]), .B(n14179), .Z(c[1450]) );
  XNOR U16827 ( .A(a[1450]), .B(n14180), .Z(n14179) );
  IV U16828 ( .A(n14177), .Z(n14180) );
  XOR U16829 ( .A(n14181), .B(n14182), .Z(n14177) );
  ANDN U16830 ( .B(n14183), .A(n14184), .Z(n14181) );
  XNOR U16831 ( .A(b[1449]), .B(n14182), .Z(n14183) );
  XNOR U16832 ( .A(b[144]), .B(n14185), .Z(c[144]) );
  XNOR U16833 ( .A(b[1449]), .B(n14184), .Z(c[1449]) );
  XNOR U16834 ( .A(a[1449]), .B(n14186), .Z(n14184) );
  IV U16835 ( .A(n14182), .Z(n14186) );
  XOR U16836 ( .A(n14187), .B(n14188), .Z(n14182) );
  ANDN U16837 ( .B(n14189), .A(n14190), .Z(n14187) );
  XNOR U16838 ( .A(b[1448]), .B(n14188), .Z(n14189) );
  XNOR U16839 ( .A(b[1448]), .B(n14190), .Z(c[1448]) );
  XNOR U16840 ( .A(a[1448]), .B(n14191), .Z(n14190) );
  IV U16841 ( .A(n14188), .Z(n14191) );
  XOR U16842 ( .A(n14192), .B(n14193), .Z(n14188) );
  ANDN U16843 ( .B(n14194), .A(n14195), .Z(n14192) );
  XNOR U16844 ( .A(b[1447]), .B(n14193), .Z(n14194) );
  XNOR U16845 ( .A(b[1447]), .B(n14195), .Z(c[1447]) );
  XNOR U16846 ( .A(a[1447]), .B(n14196), .Z(n14195) );
  IV U16847 ( .A(n14193), .Z(n14196) );
  XOR U16848 ( .A(n14197), .B(n14198), .Z(n14193) );
  ANDN U16849 ( .B(n14199), .A(n14200), .Z(n14197) );
  XNOR U16850 ( .A(b[1446]), .B(n14198), .Z(n14199) );
  XNOR U16851 ( .A(b[1446]), .B(n14200), .Z(c[1446]) );
  XNOR U16852 ( .A(a[1446]), .B(n14201), .Z(n14200) );
  IV U16853 ( .A(n14198), .Z(n14201) );
  XOR U16854 ( .A(n14202), .B(n14203), .Z(n14198) );
  ANDN U16855 ( .B(n14204), .A(n14205), .Z(n14202) );
  XNOR U16856 ( .A(b[1445]), .B(n14203), .Z(n14204) );
  XNOR U16857 ( .A(b[1445]), .B(n14205), .Z(c[1445]) );
  XNOR U16858 ( .A(a[1445]), .B(n14206), .Z(n14205) );
  IV U16859 ( .A(n14203), .Z(n14206) );
  XOR U16860 ( .A(n14207), .B(n14208), .Z(n14203) );
  ANDN U16861 ( .B(n14209), .A(n14210), .Z(n14207) );
  XNOR U16862 ( .A(b[1444]), .B(n14208), .Z(n14209) );
  XNOR U16863 ( .A(b[1444]), .B(n14210), .Z(c[1444]) );
  XNOR U16864 ( .A(a[1444]), .B(n14211), .Z(n14210) );
  IV U16865 ( .A(n14208), .Z(n14211) );
  XOR U16866 ( .A(n14212), .B(n14213), .Z(n14208) );
  ANDN U16867 ( .B(n14214), .A(n14215), .Z(n14212) );
  XNOR U16868 ( .A(b[1443]), .B(n14213), .Z(n14214) );
  XNOR U16869 ( .A(b[1443]), .B(n14215), .Z(c[1443]) );
  XNOR U16870 ( .A(a[1443]), .B(n14216), .Z(n14215) );
  IV U16871 ( .A(n14213), .Z(n14216) );
  XOR U16872 ( .A(n14217), .B(n14218), .Z(n14213) );
  ANDN U16873 ( .B(n14219), .A(n14220), .Z(n14217) );
  XNOR U16874 ( .A(b[1442]), .B(n14218), .Z(n14219) );
  XNOR U16875 ( .A(b[1442]), .B(n14220), .Z(c[1442]) );
  XNOR U16876 ( .A(a[1442]), .B(n14221), .Z(n14220) );
  IV U16877 ( .A(n14218), .Z(n14221) );
  XOR U16878 ( .A(n14222), .B(n14223), .Z(n14218) );
  ANDN U16879 ( .B(n14224), .A(n14225), .Z(n14222) );
  XNOR U16880 ( .A(b[1441]), .B(n14223), .Z(n14224) );
  XNOR U16881 ( .A(b[1441]), .B(n14225), .Z(c[1441]) );
  XNOR U16882 ( .A(a[1441]), .B(n14226), .Z(n14225) );
  IV U16883 ( .A(n14223), .Z(n14226) );
  XOR U16884 ( .A(n14227), .B(n14228), .Z(n14223) );
  ANDN U16885 ( .B(n14229), .A(n14230), .Z(n14227) );
  XNOR U16886 ( .A(b[1440]), .B(n14228), .Z(n14229) );
  XNOR U16887 ( .A(b[1440]), .B(n14230), .Z(c[1440]) );
  XNOR U16888 ( .A(a[1440]), .B(n14231), .Z(n14230) );
  IV U16889 ( .A(n14228), .Z(n14231) );
  XOR U16890 ( .A(n14232), .B(n14233), .Z(n14228) );
  ANDN U16891 ( .B(n14234), .A(n14235), .Z(n14232) );
  XNOR U16892 ( .A(b[1439]), .B(n14233), .Z(n14234) );
  XNOR U16893 ( .A(b[143]), .B(n14236), .Z(c[143]) );
  XNOR U16894 ( .A(b[1439]), .B(n14235), .Z(c[1439]) );
  XNOR U16895 ( .A(a[1439]), .B(n14237), .Z(n14235) );
  IV U16896 ( .A(n14233), .Z(n14237) );
  XOR U16897 ( .A(n14238), .B(n14239), .Z(n14233) );
  ANDN U16898 ( .B(n14240), .A(n14241), .Z(n14238) );
  XNOR U16899 ( .A(b[1438]), .B(n14239), .Z(n14240) );
  XNOR U16900 ( .A(b[1438]), .B(n14241), .Z(c[1438]) );
  XNOR U16901 ( .A(a[1438]), .B(n14242), .Z(n14241) );
  IV U16902 ( .A(n14239), .Z(n14242) );
  XOR U16903 ( .A(n14243), .B(n14244), .Z(n14239) );
  ANDN U16904 ( .B(n14245), .A(n14246), .Z(n14243) );
  XNOR U16905 ( .A(b[1437]), .B(n14244), .Z(n14245) );
  XNOR U16906 ( .A(b[1437]), .B(n14246), .Z(c[1437]) );
  XNOR U16907 ( .A(a[1437]), .B(n14247), .Z(n14246) );
  IV U16908 ( .A(n14244), .Z(n14247) );
  XOR U16909 ( .A(n14248), .B(n14249), .Z(n14244) );
  ANDN U16910 ( .B(n14250), .A(n14251), .Z(n14248) );
  XNOR U16911 ( .A(b[1436]), .B(n14249), .Z(n14250) );
  XNOR U16912 ( .A(b[1436]), .B(n14251), .Z(c[1436]) );
  XNOR U16913 ( .A(a[1436]), .B(n14252), .Z(n14251) );
  IV U16914 ( .A(n14249), .Z(n14252) );
  XOR U16915 ( .A(n14253), .B(n14254), .Z(n14249) );
  ANDN U16916 ( .B(n14255), .A(n14256), .Z(n14253) );
  XNOR U16917 ( .A(b[1435]), .B(n14254), .Z(n14255) );
  XNOR U16918 ( .A(b[1435]), .B(n14256), .Z(c[1435]) );
  XNOR U16919 ( .A(a[1435]), .B(n14257), .Z(n14256) );
  IV U16920 ( .A(n14254), .Z(n14257) );
  XOR U16921 ( .A(n14258), .B(n14259), .Z(n14254) );
  ANDN U16922 ( .B(n14260), .A(n14261), .Z(n14258) );
  XNOR U16923 ( .A(b[1434]), .B(n14259), .Z(n14260) );
  XNOR U16924 ( .A(b[1434]), .B(n14261), .Z(c[1434]) );
  XNOR U16925 ( .A(a[1434]), .B(n14262), .Z(n14261) );
  IV U16926 ( .A(n14259), .Z(n14262) );
  XOR U16927 ( .A(n14263), .B(n14264), .Z(n14259) );
  ANDN U16928 ( .B(n14265), .A(n14266), .Z(n14263) );
  XNOR U16929 ( .A(b[1433]), .B(n14264), .Z(n14265) );
  XNOR U16930 ( .A(b[1433]), .B(n14266), .Z(c[1433]) );
  XNOR U16931 ( .A(a[1433]), .B(n14267), .Z(n14266) );
  IV U16932 ( .A(n14264), .Z(n14267) );
  XOR U16933 ( .A(n14268), .B(n14269), .Z(n14264) );
  ANDN U16934 ( .B(n14270), .A(n14271), .Z(n14268) );
  XNOR U16935 ( .A(b[1432]), .B(n14269), .Z(n14270) );
  XNOR U16936 ( .A(b[1432]), .B(n14271), .Z(c[1432]) );
  XNOR U16937 ( .A(a[1432]), .B(n14272), .Z(n14271) );
  IV U16938 ( .A(n14269), .Z(n14272) );
  XOR U16939 ( .A(n14273), .B(n14274), .Z(n14269) );
  ANDN U16940 ( .B(n14275), .A(n14276), .Z(n14273) );
  XNOR U16941 ( .A(b[1431]), .B(n14274), .Z(n14275) );
  XNOR U16942 ( .A(b[1431]), .B(n14276), .Z(c[1431]) );
  XNOR U16943 ( .A(a[1431]), .B(n14277), .Z(n14276) );
  IV U16944 ( .A(n14274), .Z(n14277) );
  XOR U16945 ( .A(n14278), .B(n14279), .Z(n14274) );
  ANDN U16946 ( .B(n14280), .A(n14281), .Z(n14278) );
  XNOR U16947 ( .A(b[1430]), .B(n14279), .Z(n14280) );
  XNOR U16948 ( .A(b[1430]), .B(n14281), .Z(c[1430]) );
  XNOR U16949 ( .A(a[1430]), .B(n14282), .Z(n14281) );
  IV U16950 ( .A(n14279), .Z(n14282) );
  XOR U16951 ( .A(n14283), .B(n14284), .Z(n14279) );
  ANDN U16952 ( .B(n14285), .A(n14286), .Z(n14283) );
  XNOR U16953 ( .A(b[1429]), .B(n14284), .Z(n14285) );
  XNOR U16954 ( .A(b[142]), .B(n14287), .Z(c[142]) );
  XNOR U16955 ( .A(b[1429]), .B(n14286), .Z(c[1429]) );
  XNOR U16956 ( .A(a[1429]), .B(n14288), .Z(n14286) );
  IV U16957 ( .A(n14284), .Z(n14288) );
  XOR U16958 ( .A(n14289), .B(n14290), .Z(n14284) );
  ANDN U16959 ( .B(n14291), .A(n14292), .Z(n14289) );
  XNOR U16960 ( .A(b[1428]), .B(n14290), .Z(n14291) );
  XNOR U16961 ( .A(b[1428]), .B(n14292), .Z(c[1428]) );
  XNOR U16962 ( .A(a[1428]), .B(n14293), .Z(n14292) );
  IV U16963 ( .A(n14290), .Z(n14293) );
  XOR U16964 ( .A(n14294), .B(n14295), .Z(n14290) );
  ANDN U16965 ( .B(n14296), .A(n14297), .Z(n14294) );
  XNOR U16966 ( .A(b[1427]), .B(n14295), .Z(n14296) );
  XNOR U16967 ( .A(b[1427]), .B(n14297), .Z(c[1427]) );
  XNOR U16968 ( .A(a[1427]), .B(n14298), .Z(n14297) );
  IV U16969 ( .A(n14295), .Z(n14298) );
  XOR U16970 ( .A(n14299), .B(n14300), .Z(n14295) );
  ANDN U16971 ( .B(n14301), .A(n14302), .Z(n14299) );
  XNOR U16972 ( .A(b[1426]), .B(n14300), .Z(n14301) );
  XNOR U16973 ( .A(b[1426]), .B(n14302), .Z(c[1426]) );
  XNOR U16974 ( .A(a[1426]), .B(n14303), .Z(n14302) );
  IV U16975 ( .A(n14300), .Z(n14303) );
  XOR U16976 ( .A(n14304), .B(n14305), .Z(n14300) );
  ANDN U16977 ( .B(n14306), .A(n14307), .Z(n14304) );
  XNOR U16978 ( .A(b[1425]), .B(n14305), .Z(n14306) );
  XNOR U16979 ( .A(b[1425]), .B(n14307), .Z(c[1425]) );
  XNOR U16980 ( .A(a[1425]), .B(n14308), .Z(n14307) );
  IV U16981 ( .A(n14305), .Z(n14308) );
  XOR U16982 ( .A(n14309), .B(n14310), .Z(n14305) );
  ANDN U16983 ( .B(n14311), .A(n14312), .Z(n14309) );
  XNOR U16984 ( .A(b[1424]), .B(n14310), .Z(n14311) );
  XNOR U16985 ( .A(b[1424]), .B(n14312), .Z(c[1424]) );
  XNOR U16986 ( .A(a[1424]), .B(n14313), .Z(n14312) );
  IV U16987 ( .A(n14310), .Z(n14313) );
  XOR U16988 ( .A(n14314), .B(n14315), .Z(n14310) );
  ANDN U16989 ( .B(n14316), .A(n14317), .Z(n14314) );
  XNOR U16990 ( .A(b[1423]), .B(n14315), .Z(n14316) );
  XNOR U16991 ( .A(b[1423]), .B(n14317), .Z(c[1423]) );
  XNOR U16992 ( .A(a[1423]), .B(n14318), .Z(n14317) );
  IV U16993 ( .A(n14315), .Z(n14318) );
  XOR U16994 ( .A(n14319), .B(n14320), .Z(n14315) );
  ANDN U16995 ( .B(n14321), .A(n14322), .Z(n14319) );
  XNOR U16996 ( .A(b[1422]), .B(n14320), .Z(n14321) );
  XNOR U16997 ( .A(b[1422]), .B(n14322), .Z(c[1422]) );
  XNOR U16998 ( .A(a[1422]), .B(n14323), .Z(n14322) );
  IV U16999 ( .A(n14320), .Z(n14323) );
  XOR U17000 ( .A(n14324), .B(n14325), .Z(n14320) );
  ANDN U17001 ( .B(n14326), .A(n14327), .Z(n14324) );
  XNOR U17002 ( .A(b[1421]), .B(n14325), .Z(n14326) );
  XNOR U17003 ( .A(b[1421]), .B(n14327), .Z(c[1421]) );
  XNOR U17004 ( .A(a[1421]), .B(n14328), .Z(n14327) );
  IV U17005 ( .A(n14325), .Z(n14328) );
  XOR U17006 ( .A(n14329), .B(n14330), .Z(n14325) );
  ANDN U17007 ( .B(n14331), .A(n14332), .Z(n14329) );
  XNOR U17008 ( .A(b[1420]), .B(n14330), .Z(n14331) );
  XNOR U17009 ( .A(b[1420]), .B(n14332), .Z(c[1420]) );
  XNOR U17010 ( .A(a[1420]), .B(n14333), .Z(n14332) );
  IV U17011 ( .A(n14330), .Z(n14333) );
  XOR U17012 ( .A(n14334), .B(n14335), .Z(n14330) );
  ANDN U17013 ( .B(n14336), .A(n14337), .Z(n14334) );
  XNOR U17014 ( .A(b[1419]), .B(n14335), .Z(n14336) );
  XNOR U17015 ( .A(b[141]), .B(n14338), .Z(c[141]) );
  XNOR U17016 ( .A(b[1419]), .B(n14337), .Z(c[1419]) );
  XNOR U17017 ( .A(a[1419]), .B(n14339), .Z(n14337) );
  IV U17018 ( .A(n14335), .Z(n14339) );
  XOR U17019 ( .A(n14340), .B(n14341), .Z(n14335) );
  ANDN U17020 ( .B(n14342), .A(n14343), .Z(n14340) );
  XNOR U17021 ( .A(b[1418]), .B(n14341), .Z(n14342) );
  XNOR U17022 ( .A(b[1418]), .B(n14343), .Z(c[1418]) );
  XNOR U17023 ( .A(a[1418]), .B(n14344), .Z(n14343) );
  IV U17024 ( .A(n14341), .Z(n14344) );
  XOR U17025 ( .A(n14345), .B(n14346), .Z(n14341) );
  ANDN U17026 ( .B(n14347), .A(n14348), .Z(n14345) );
  XNOR U17027 ( .A(b[1417]), .B(n14346), .Z(n14347) );
  XNOR U17028 ( .A(b[1417]), .B(n14348), .Z(c[1417]) );
  XNOR U17029 ( .A(a[1417]), .B(n14349), .Z(n14348) );
  IV U17030 ( .A(n14346), .Z(n14349) );
  XOR U17031 ( .A(n14350), .B(n14351), .Z(n14346) );
  ANDN U17032 ( .B(n14352), .A(n14353), .Z(n14350) );
  XNOR U17033 ( .A(b[1416]), .B(n14351), .Z(n14352) );
  XNOR U17034 ( .A(b[1416]), .B(n14353), .Z(c[1416]) );
  XNOR U17035 ( .A(a[1416]), .B(n14354), .Z(n14353) );
  IV U17036 ( .A(n14351), .Z(n14354) );
  XOR U17037 ( .A(n14355), .B(n14356), .Z(n14351) );
  ANDN U17038 ( .B(n14357), .A(n14358), .Z(n14355) );
  XNOR U17039 ( .A(b[1415]), .B(n14356), .Z(n14357) );
  XNOR U17040 ( .A(b[1415]), .B(n14358), .Z(c[1415]) );
  XNOR U17041 ( .A(a[1415]), .B(n14359), .Z(n14358) );
  IV U17042 ( .A(n14356), .Z(n14359) );
  XOR U17043 ( .A(n14360), .B(n14361), .Z(n14356) );
  ANDN U17044 ( .B(n14362), .A(n14363), .Z(n14360) );
  XNOR U17045 ( .A(b[1414]), .B(n14361), .Z(n14362) );
  XNOR U17046 ( .A(b[1414]), .B(n14363), .Z(c[1414]) );
  XNOR U17047 ( .A(a[1414]), .B(n14364), .Z(n14363) );
  IV U17048 ( .A(n14361), .Z(n14364) );
  XOR U17049 ( .A(n14365), .B(n14366), .Z(n14361) );
  ANDN U17050 ( .B(n14367), .A(n14368), .Z(n14365) );
  XNOR U17051 ( .A(b[1413]), .B(n14366), .Z(n14367) );
  XNOR U17052 ( .A(b[1413]), .B(n14368), .Z(c[1413]) );
  XNOR U17053 ( .A(a[1413]), .B(n14369), .Z(n14368) );
  IV U17054 ( .A(n14366), .Z(n14369) );
  XOR U17055 ( .A(n14370), .B(n14371), .Z(n14366) );
  ANDN U17056 ( .B(n14372), .A(n14373), .Z(n14370) );
  XNOR U17057 ( .A(b[1412]), .B(n14371), .Z(n14372) );
  XNOR U17058 ( .A(b[1412]), .B(n14373), .Z(c[1412]) );
  XNOR U17059 ( .A(a[1412]), .B(n14374), .Z(n14373) );
  IV U17060 ( .A(n14371), .Z(n14374) );
  XOR U17061 ( .A(n14375), .B(n14376), .Z(n14371) );
  ANDN U17062 ( .B(n14377), .A(n14378), .Z(n14375) );
  XNOR U17063 ( .A(b[1411]), .B(n14376), .Z(n14377) );
  XNOR U17064 ( .A(b[1411]), .B(n14378), .Z(c[1411]) );
  XNOR U17065 ( .A(a[1411]), .B(n14379), .Z(n14378) );
  IV U17066 ( .A(n14376), .Z(n14379) );
  XOR U17067 ( .A(n14380), .B(n14381), .Z(n14376) );
  ANDN U17068 ( .B(n14382), .A(n14383), .Z(n14380) );
  XNOR U17069 ( .A(b[1410]), .B(n14381), .Z(n14382) );
  XNOR U17070 ( .A(b[1410]), .B(n14383), .Z(c[1410]) );
  XNOR U17071 ( .A(a[1410]), .B(n14384), .Z(n14383) );
  IV U17072 ( .A(n14381), .Z(n14384) );
  XOR U17073 ( .A(n14385), .B(n14386), .Z(n14381) );
  ANDN U17074 ( .B(n14387), .A(n14388), .Z(n14385) );
  XNOR U17075 ( .A(b[1409]), .B(n14386), .Z(n14387) );
  XNOR U17076 ( .A(b[140]), .B(n14389), .Z(c[140]) );
  XNOR U17077 ( .A(b[1409]), .B(n14388), .Z(c[1409]) );
  XNOR U17078 ( .A(a[1409]), .B(n14390), .Z(n14388) );
  IV U17079 ( .A(n14386), .Z(n14390) );
  XOR U17080 ( .A(n14391), .B(n14392), .Z(n14386) );
  ANDN U17081 ( .B(n14393), .A(n14394), .Z(n14391) );
  XNOR U17082 ( .A(b[1408]), .B(n14392), .Z(n14393) );
  XNOR U17083 ( .A(b[1408]), .B(n14394), .Z(c[1408]) );
  XNOR U17084 ( .A(a[1408]), .B(n14395), .Z(n14394) );
  IV U17085 ( .A(n14392), .Z(n14395) );
  XOR U17086 ( .A(n14396), .B(n14397), .Z(n14392) );
  ANDN U17087 ( .B(n14398), .A(n14399), .Z(n14396) );
  XNOR U17088 ( .A(b[1407]), .B(n14397), .Z(n14398) );
  XNOR U17089 ( .A(b[1407]), .B(n14399), .Z(c[1407]) );
  XNOR U17090 ( .A(a[1407]), .B(n14400), .Z(n14399) );
  IV U17091 ( .A(n14397), .Z(n14400) );
  XOR U17092 ( .A(n14401), .B(n14402), .Z(n14397) );
  ANDN U17093 ( .B(n14403), .A(n14404), .Z(n14401) );
  XNOR U17094 ( .A(b[1406]), .B(n14402), .Z(n14403) );
  XNOR U17095 ( .A(b[1406]), .B(n14404), .Z(c[1406]) );
  XNOR U17096 ( .A(a[1406]), .B(n14405), .Z(n14404) );
  IV U17097 ( .A(n14402), .Z(n14405) );
  XOR U17098 ( .A(n14406), .B(n14407), .Z(n14402) );
  ANDN U17099 ( .B(n14408), .A(n14409), .Z(n14406) );
  XNOR U17100 ( .A(b[1405]), .B(n14407), .Z(n14408) );
  XNOR U17101 ( .A(b[1405]), .B(n14409), .Z(c[1405]) );
  XNOR U17102 ( .A(a[1405]), .B(n14410), .Z(n14409) );
  IV U17103 ( .A(n14407), .Z(n14410) );
  XOR U17104 ( .A(n14411), .B(n14412), .Z(n14407) );
  ANDN U17105 ( .B(n14413), .A(n14414), .Z(n14411) );
  XNOR U17106 ( .A(b[1404]), .B(n14412), .Z(n14413) );
  XNOR U17107 ( .A(b[1404]), .B(n14414), .Z(c[1404]) );
  XNOR U17108 ( .A(a[1404]), .B(n14415), .Z(n14414) );
  IV U17109 ( .A(n14412), .Z(n14415) );
  XOR U17110 ( .A(n14416), .B(n14417), .Z(n14412) );
  ANDN U17111 ( .B(n14418), .A(n14419), .Z(n14416) );
  XNOR U17112 ( .A(b[1403]), .B(n14417), .Z(n14418) );
  XNOR U17113 ( .A(b[1403]), .B(n14419), .Z(c[1403]) );
  XNOR U17114 ( .A(a[1403]), .B(n14420), .Z(n14419) );
  IV U17115 ( .A(n14417), .Z(n14420) );
  XOR U17116 ( .A(n14421), .B(n14422), .Z(n14417) );
  ANDN U17117 ( .B(n14423), .A(n14424), .Z(n14421) );
  XNOR U17118 ( .A(b[1402]), .B(n14422), .Z(n14423) );
  XNOR U17119 ( .A(b[1402]), .B(n14424), .Z(c[1402]) );
  XNOR U17120 ( .A(a[1402]), .B(n14425), .Z(n14424) );
  IV U17121 ( .A(n14422), .Z(n14425) );
  XOR U17122 ( .A(n14426), .B(n14427), .Z(n14422) );
  ANDN U17123 ( .B(n14428), .A(n14429), .Z(n14426) );
  XNOR U17124 ( .A(b[1401]), .B(n14427), .Z(n14428) );
  XNOR U17125 ( .A(b[1401]), .B(n14429), .Z(c[1401]) );
  XNOR U17126 ( .A(a[1401]), .B(n14430), .Z(n14429) );
  IV U17127 ( .A(n14427), .Z(n14430) );
  XOR U17128 ( .A(n14431), .B(n14432), .Z(n14427) );
  ANDN U17129 ( .B(n14433), .A(n14434), .Z(n14431) );
  XNOR U17130 ( .A(b[1400]), .B(n14432), .Z(n14433) );
  XNOR U17131 ( .A(b[1400]), .B(n14434), .Z(c[1400]) );
  XNOR U17132 ( .A(a[1400]), .B(n14435), .Z(n14434) );
  IV U17133 ( .A(n14432), .Z(n14435) );
  XOR U17134 ( .A(n14436), .B(n14437), .Z(n14432) );
  ANDN U17135 ( .B(n14438), .A(n14439), .Z(n14436) );
  XNOR U17136 ( .A(b[1399]), .B(n14437), .Z(n14438) );
  XNOR U17137 ( .A(b[13]), .B(n14440), .Z(c[13]) );
  XNOR U17138 ( .A(b[139]), .B(n14441), .Z(c[139]) );
  XNOR U17139 ( .A(b[1399]), .B(n14439), .Z(c[1399]) );
  XNOR U17140 ( .A(a[1399]), .B(n14442), .Z(n14439) );
  IV U17141 ( .A(n14437), .Z(n14442) );
  XOR U17142 ( .A(n14443), .B(n14444), .Z(n14437) );
  ANDN U17143 ( .B(n14445), .A(n14446), .Z(n14443) );
  XNOR U17144 ( .A(b[1398]), .B(n14444), .Z(n14445) );
  XNOR U17145 ( .A(b[1398]), .B(n14446), .Z(c[1398]) );
  XNOR U17146 ( .A(a[1398]), .B(n14447), .Z(n14446) );
  IV U17147 ( .A(n14444), .Z(n14447) );
  XOR U17148 ( .A(n14448), .B(n14449), .Z(n14444) );
  ANDN U17149 ( .B(n14450), .A(n14451), .Z(n14448) );
  XNOR U17150 ( .A(b[1397]), .B(n14449), .Z(n14450) );
  XNOR U17151 ( .A(b[1397]), .B(n14451), .Z(c[1397]) );
  XNOR U17152 ( .A(a[1397]), .B(n14452), .Z(n14451) );
  IV U17153 ( .A(n14449), .Z(n14452) );
  XOR U17154 ( .A(n14453), .B(n14454), .Z(n14449) );
  ANDN U17155 ( .B(n14455), .A(n14456), .Z(n14453) );
  XNOR U17156 ( .A(b[1396]), .B(n14454), .Z(n14455) );
  XNOR U17157 ( .A(b[1396]), .B(n14456), .Z(c[1396]) );
  XNOR U17158 ( .A(a[1396]), .B(n14457), .Z(n14456) );
  IV U17159 ( .A(n14454), .Z(n14457) );
  XOR U17160 ( .A(n14458), .B(n14459), .Z(n14454) );
  ANDN U17161 ( .B(n14460), .A(n14461), .Z(n14458) );
  XNOR U17162 ( .A(b[1395]), .B(n14459), .Z(n14460) );
  XNOR U17163 ( .A(b[1395]), .B(n14461), .Z(c[1395]) );
  XNOR U17164 ( .A(a[1395]), .B(n14462), .Z(n14461) );
  IV U17165 ( .A(n14459), .Z(n14462) );
  XOR U17166 ( .A(n14463), .B(n14464), .Z(n14459) );
  ANDN U17167 ( .B(n14465), .A(n14466), .Z(n14463) );
  XNOR U17168 ( .A(b[1394]), .B(n14464), .Z(n14465) );
  XNOR U17169 ( .A(b[1394]), .B(n14466), .Z(c[1394]) );
  XNOR U17170 ( .A(a[1394]), .B(n14467), .Z(n14466) );
  IV U17171 ( .A(n14464), .Z(n14467) );
  XOR U17172 ( .A(n14468), .B(n14469), .Z(n14464) );
  ANDN U17173 ( .B(n14470), .A(n14471), .Z(n14468) );
  XNOR U17174 ( .A(b[1393]), .B(n14469), .Z(n14470) );
  XNOR U17175 ( .A(b[1393]), .B(n14471), .Z(c[1393]) );
  XNOR U17176 ( .A(a[1393]), .B(n14472), .Z(n14471) );
  IV U17177 ( .A(n14469), .Z(n14472) );
  XOR U17178 ( .A(n14473), .B(n14474), .Z(n14469) );
  ANDN U17179 ( .B(n14475), .A(n14476), .Z(n14473) );
  XNOR U17180 ( .A(b[1392]), .B(n14474), .Z(n14475) );
  XNOR U17181 ( .A(b[1392]), .B(n14476), .Z(c[1392]) );
  XNOR U17182 ( .A(a[1392]), .B(n14477), .Z(n14476) );
  IV U17183 ( .A(n14474), .Z(n14477) );
  XOR U17184 ( .A(n14478), .B(n14479), .Z(n14474) );
  ANDN U17185 ( .B(n14480), .A(n14481), .Z(n14478) );
  XNOR U17186 ( .A(b[1391]), .B(n14479), .Z(n14480) );
  XNOR U17187 ( .A(b[1391]), .B(n14481), .Z(c[1391]) );
  XNOR U17188 ( .A(a[1391]), .B(n14482), .Z(n14481) );
  IV U17189 ( .A(n14479), .Z(n14482) );
  XOR U17190 ( .A(n14483), .B(n14484), .Z(n14479) );
  ANDN U17191 ( .B(n14485), .A(n14486), .Z(n14483) );
  XNOR U17192 ( .A(b[1390]), .B(n14484), .Z(n14485) );
  XNOR U17193 ( .A(b[1390]), .B(n14486), .Z(c[1390]) );
  XNOR U17194 ( .A(a[1390]), .B(n14487), .Z(n14486) );
  IV U17195 ( .A(n14484), .Z(n14487) );
  XOR U17196 ( .A(n14488), .B(n14489), .Z(n14484) );
  ANDN U17197 ( .B(n14490), .A(n14491), .Z(n14488) );
  XNOR U17198 ( .A(b[1389]), .B(n14489), .Z(n14490) );
  XNOR U17199 ( .A(b[138]), .B(n14492), .Z(c[138]) );
  XNOR U17200 ( .A(b[1389]), .B(n14491), .Z(c[1389]) );
  XNOR U17201 ( .A(a[1389]), .B(n14493), .Z(n14491) );
  IV U17202 ( .A(n14489), .Z(n14493) );
  XOR U17203 ( .A(n14494), .B(n14495), .Z(n14489) );
  ANDN U17204 ( .B(n14496), .A(n14497), .Z(n14494) );
  XNOR U17205 ( .A(b[1388]), .B(n14495), .Z(n14496) );
  XNOR U17206 ( .A(b[1388]), .B(n14497), .Z(c[1388]) );
  XNOR U17207 ( .A(a[1388]), .B(n14498), .Z(n14497) );
  IV U17208 ( .A(n14495), .Z(n14498) );
  XOR U17209 ( .A(n14499), .B(n14500), .Z(n14495) );
  ANDN U17210 ( .B(n14501), .A(n14502), .Z(n14499) );
  XNOR U17211 ( .A(b[1387]), .B(n14500), .Z(n14501) );
  XNOR U17212 ( .A(b[1387]), .B(n14502), .Z(c[1387]) );
  XNOR U17213 ( .A(a[1387]), .B(n14503), .Z(n14502) );
  IV U17214 ( .A(n14500), .Z(n14503) );
  XOR U17215 ( .A(n14504), .B(n14505), .Z(n14500) );
  ANDN U17216 ( .B(n14506), .A(n14507), .Z(n14504) );
  XNOR U17217 ( .A(b[1386]), .B(n14505), .Z(n14506) );
  XNOR U17218 ( .A(b[1386]), .B(n14507), .Z(c[1386]) );
  XNOR U17219 ( .A(a[1386]), .B(n14508), .Z(n14507) );
  IV U17220 ( .A(n14505), .Z(n14508) );
  XOR U17221 ( .A(n14509), .B(n14510), .Z(n14505) );
  ANDN U17222 ( .B(n14511), .A(n14512), .Z(n14509) );
  XNOR U17223 ( .A(b[1385]), .B(n14510), .Z(n14511) );
  XNOR U17224 ( .A(b[1385]), .B(n14512), .Z(c[1385]) );
  XNOR U17225 ( .A(a[1385]), .B(n14513), .Z(n14512) );
  IV U17226 ( .A(n14510), .Z(n14513) );
  XOR U17227 ( .A(n14514), .B(n14515), .Z(n14510) );
  ANDN U17228 ( .B(n14516), .A(n14517), .Z(n14514) );
  XNOR U17229 ( .A(b[1384]), .B(n14515), .Z(n14516) );
  XNOR U17230 ( .A(b[1384]), .B(n14517), .Z(c[1384]) );
  XNOR U17231 ( .A(a[1384]), .B(n14518), .Z(n14517) );
  IV U17232 ( .A(n14515), .Z(n14518) );
  XOR U17233 ( .A(n14519), .B(n14520), .Z(n14515) );
  ANDN U17234 ( .B(n14521), .A(n14522), .Z(n14519) );
  XNOR U17235 ( .A(b[1383]), .B(n14520), .Z(n14521) );
  XNOR U17236 ( .A(b[1383]), .B(n14522), .Z(c[1383]) );
  XNOR U17237 ( .A(a[1383]), .B(n14523), .Z(n14522) );
  IV U17238 ( .A(n14520), .Z(n14523) );
  XOR U17239 ( .A(n14524), .B(n14525), .Z(n14520) );
  ANDN U17240 ( .B(n14526), .A(n14527), .Z(n14524) );
  XNOR U17241 ( .A(b[1382]), .B(n14525), .Z(n14526) );
  XNOR U17242 ( .A(b[1382]), .B(n14527), .Z(c[1382]) );
  XNOR U17243 ( .A(a[1382]), .B(n14528), .Z(n14527) );
  IV U17244 ( .A(n14525), .Z(n14528) );
  XOR U17245 ( .A(n14529), .B(n14530), .Z(n14525) );
  ANDN U17246 ( .B(n14531), .A(n14532), .Z(n14529) );
  XNOR U17247 ( .A(b[1381]), .B(n14530), .Z(n14531) );
  XNOR U17248 ( .A(b[1381]), .B(n14532), .Z(c[1381]) );
  XNOR U17249 ( .A(a[1381]), .B(n14533), .Z(n14532) );
  IV U17250 ( .A(n14530), .Z(n14533) );
  XOR U17251 ( .A(n14534), .B(n14535), .Z(n14530) );
  ANDN U17252 ( .B(n14536), .A(n14537), .Z(n14534) );
  XNOR U17253 ( .A(b[1380]), .B(n14535), .Z(n14536) );
  XNOR U17254 ( .A(b[1380]), .B(n14537), .Z(c[1380]) );
  XNOR U17255 ( .A(a[1380]), .B(n14538), .Z(n14537) );
  IV U17256 ( .A(n14535), .Z(n14538) );
  XOR U17257 ( .A(n14539), .B(n14540), .Z(n14535) );
  ANDN U17258 ( .B(n14541), .A(n14542), .Z(n14539) );
  XNOR U17259 ( .A(b[1379]), .B(n14540), .Z(n14541) );
  XNOR U17260 ( .A(b[137]), .B(n14543), .Z(c[137]) );
  XNOR U17261 ( .A(b[1379]), .B(n14542), .Z(c[1379]) );
  XNOR U17262 ( .A(a[1379]), .B(n14544), .Z(n14542) );
  IV U17263 ( .A(n14540), .Z(n14544) );
  XOR U17264 ( .A(n14545), .B(n14546), .Z(n14540) );
  ANDN U17265 ( .B(n14547), .A(n14548), .Z(n14545) );
  XNOR U17266 ( .A(b[1378]), .B(n14546), .Z(n14547) );
  XNOR U17267 ( .A(b[1378]), .B(n14548), .Z(c[1378]) );
  XNOR U17268 ( .A(a[1378]), .B(n14549), .Z(n14548) );
  IV U17269 ( .A(n14546), .Z(n14549) );
  XOR U17270 ( .A(n14550), .B(n14551), .Z(n14546) );
  ANDN U17271 ( .B(n14552), .A(n14553), .Z(n14550) );
  XNOR U17272 ( .A(b[1377]), .B(n14551), .Z(n14552) );
  XNOR U17273 ( .A(b[1377]), .B(n14553), .Z(c[1377]) );
  XNOR U17274 ( .A(a[1377]), .B(n14554), .Z(n14553) );
  IV U17275 ( .A(n14551), .Z(n14554) );
  XOR U17276 ( .A(n14555), .B(n14556), .Z(n14551) );
  ANDN U17277 ( .B(n14557), .A(n14558), .Z(n14555) );
  XNOR U17278 ( .A(b[1376]), .B(n14556), .Z(n14557) );
  XNOR U17279 ( .A(b[1376]), .B(n14558), .Z(c[1376]) );
  XNOR U17280 ( .A(a[1376]), .B(n14559), .Z(n14558) );
  IV U17281 ( .A(n14556), .Z(n14559) );
  XOR U17282 ( .A(n14560), .B(n14561), .Z(n14556) );
  ANDN U17283 ( .B(n14562), .A(n14563), .Z(n14560) );
  XNOR U17284 ( .A(b[1375]), .B(n14561), .Z(n14562) );
  XNOR U17285 ( .A(b[1375]), .B(n14563), .Z(c[1375]) );
  XNOR U17286 ( .A(a[1375]), .B(n14564), .Z(n14563) );
  IV U17287 ( .A(n14561), .Z(n14564) );
  XOR U17288 ( .A(n14565), .B(n14566), .Z(n14561) );
  ANDN U17289 ( .B(n14567), .A(n14568), .Z(n14565) );
  XNOR U17290 ( .A(b[1374]), .B(n14566), .Z(n14567) );
  XNOR U17291 ( .A(b[1374]), .B(n14568), .Z(c[1374]) );
  XNOR U17292 ( .A(a[1374]), .B(n14569), .Z(n14568) );
  IV U17293 ( .A(n14566), .Z(n14569) );
  XOR U17294 ( .A(n14570), .B(n14571), .Z(n14566) );
  ANDN U17295 ( .B(n14572), .A(n14573), .Z(n14570) );
  XNOR U17296 ( .A(b[1373]), .B(n14571), .Z(n14572) );
  XNOR U17297 ( .A(b[1373]), .B(n14573), .Z(c[1373]) );
  XNOR U17298 ( .A(a[1373]), .B(n14574), .Z(n14573) );
  IV U17299 ( .A(n14571), .Z(n14574) );
  XOR U17300 ( .A(n14575), .B(n14576), .Z(n14571) );
  ANDN U17301 ( .B(n14577), .A(n14578), .Z(n14575) );
  XNOR U17302 ( .A(b[1372]), .B(n14576), .Z(n14577) );
  XNOR U17303 ( .A(b[1372]), .B(n14578), .Z(c[1372]) );
  XNOR U17304 ( .A(a[1372]), .B(n14579), .Z(n14578) );
  IV U17305 ( .A(n14576), .Z(n14579) );
  XOR U17306 ( .A(n14580), .B(n14581), .Z(n14576) );
  ANDN U17307 ( .B(n14582), .A(n14583), .Z(n14580) );
  XNOR U17308 ( .A(b[1371]), .B(n14581), .Z(n14582) );
  XNOR U17309 ( .A(b[1371]), .B(n14583), .Z(c[1371]) );
  XNOR U17310 ( .A(a[1371]), .B(n14584), .Z(n14583) );
  IV U17311 ( .A(n14581), .Z(n14584) );
  XOR U17312 ( .A(n14585), .B(n14586), .Z(n14581) );
  ANDN U17313 ( .B(n14587), .A(n14588), .Z(n14585) );
  XNOR U17314 ( .A(b[1370]), .B(n14586), .Z(n14587) );
  XNOR U17315 ( .A(b[1370]), .B(n14588), .Z(c[1370]) );
  XNOR U17316 ( .A(a[1370]), .B(n14589), .Z(n14588) );
  IV U17317 ( .A(n14586), .Z(n14589) );
  XOR U17318 ( .A(n14590), .B(n14591), .Z(n14586) );
  ANDN U17319 ( .B(n14592), .A(n14593), .Z(n14590) );
  XNOR U17320 ( .A(b[1369]), .B(n14591), .Z(n14592) );
  XNOR U17321 ( .A(b[136]), .B(n14594), .Z(c[136]) );
  XNOR U17322 ( .A(b[1369]), .B(n14593), .Z(c[1369]) );
  XNOR U17323 ( .A(a[1369]), .B(n14595), .Z(n14593) );
  IV U17324 ( .A(n14591), .Z(n14595) );
  XOR U17325 ( .A(n14596), .B(n14597), .Z(n14591) );
  ANDN U17326 ( .B(n14598), .A(n14599), .Z(n14596) );
  XNOR U17327 ( .A(b[1368]), .B(n14597), .Z(n14598) );
  XNOR U17328 ( .A(b[1368]), .B(n14599), .Z(c[1368]) );
  XNOR U17329 ( .A(a[1368]), .B(n14600), .Z(n14599) );
  IV U17330 ( .A(n14597), .Z(n14600) );
  XOR U17331 ( .A(n14601), .B(n14602), .Z(n14597) );
  ANDN U17332 ( .B(n14603), .A(n14604), .Z(n14601) );
  XNOR U17333 ( .A(b[1367]), .B(n14602), .Z(n14603) );
  XNOR U17334 ( .A(b[1367]), .B(n14604), .Z(c[1367]) );
  XNOR U17335 ( .A(a[1367]), .B(n14605), .Z(n14604) );
  IV U17336 ( .A(n14602), .Z(n14605) );
  XOR U17337 ( .A(n14606), .B(n14607), .Z(n14602) );
  ANDN U17338 ( .B(n14608), .A(n14609), .Z(n14606) );
  XNOR U17339 ( .A(b[1366]), .B(n14607), .Z(n14608) );
  XNOR U17340 ( .A(b[1366]), .B(n14609), .Z(c[1366]) );
  XNOR U17341 ( .A(a[1366]), .B(n14610), .Z(n14609) );
  IV U17342 ( .A(n14607), .Z(n14610) );
  XOR U17343 ( .A(n14611), .B(n14612), .Z(n14607) );
  ANDN U17344 ( .B(n14613), .A(n14614), .Z(n14611) );
  XNOR U17345 ( .A(b[1365]), .B(n14612), .Z(n14613) );
  XNOR U17346 ( .A(b[1365]), .B(n14614), .Z(c[1365]) );
  XNOR U17347 ( .A(a[1365]), .B(n14615), .Z(n14614) );
  IV U17348 ( .A(n14612), .Z(n14615) );
  XOR U17349 ( .A(n14616), .B(n14617), .Z(n14612) );
  ANDN U17350 ( .B(n14618), .A(n14619), .Z(n14616) );
  XNOR U17351 ( .A(b[1364]), .B(n14617), .Z(n14618) );
  XNOR U17352 ( .A(b[1364]), .B(n14619), .Z(c[1364]) );
  XNOR U17353 ( .A(a[1364]), .B(n14620), .Z(n14619) );
  IV U17354 ( .A(n14617), .Z(n14620) );
  XOR U17355 ( .A(n14621), .B(n14622), .Z(n14617) );
  ANDN U17356 ( .B(n14623), .A(n14624), .Z(n14621) );
  XNOR U17357 ( .A(b[1363]), .B(n14622), .Z(n14623) );
  XNOR U17358 ( .A(b[1363]), .B(n14624), .Z(c[1363]) );
  XNOR U17359 ( .A(a[1363]), .B(n14625), .Z(n14624) );
  IV U17360 ( .A(n14622), .Z(n14625) );
  XOR U17361 ( .A(n14626), .B(n14627), .Z(n14622) );
  ANDN U17362 ( .B(n14628), .A(n14629), .Z(n14626) );
  XNOR U17363 ( .A(b[1362]), .B(n14627), .Z(n14628) );
  XNOR U17364 ( .A(b[1362]), .B(n14629), .Z(c[1362]) );
  XNOR U17365 ( .A(a[1362]), .B(n14630), .Z(n14629) );
  IV U17366 ( .A(n14627), .Z(n14630) );
  XOR U17367 ( .A(n14631), .B(n14632), .Z(n14627) );
  ANDN U17368 ( .B(n14633), .A(n14634), .Z(n14631) );
  XNOR U17369 ( .A(b[1361]), .B(n14632), .Z(n14633) );
  XNOR U17370 ( .A(b[1361]), .B(n14634), .Z(c[1361]) );
  XNOR U17371 ( .A(a[1361]), .B(n14635), .Z(n14634) );
  IV U17372 ( .A(n14632), .Z(n14635) );
  XOR U17373 ( .A(n14636), .B(n14637), .Z(n14632) );
  ANDN U17374 ( .B(n14638), .A(n14639), .Z(n14636) );
  XNOR U17375 ( .A(b[1360]), .B(n14637), .Z(n14638) );
  XNOR U17376 ( .A(b[1360]), .B(n14639), .Z(c[1360]) );
  XNOR U17377 ( .A(a[1360]), .B(n14640), .Z(n14639) );
  IV U17378 ( .A(n14637), .Z(n14640) );
  XOR U17379 ( .A(n14641), .B(n14642), .Z(n14637) );
  ANDN U17380 ( .B(n14643), .A(n14644), .Z(n14641) );
  XNOR U17381 ( .A(b[1359]), .B(n14642), .Z(n14643) );
  XNOR U17382 ( .A(b[135]), .B(n14645), .Z(c[135]) );
  XNOR U17383 ( .A(b[1359]), .B(n14644), .Z(c[1359]) );
  XNOR U17384 ( .A(a[1359]), .B(n14646), .Z(n14644) );
  IV U17385 ( .A(n14642), .Z(n14646) );
  XOR U17386 ( .A(n14647), .B(n14648), .Z(n14642) );
  ANDN U17387 ( .B(n14649), .A(n14650), .Z(n14647) );
  XNOR U17388 ( .A(b[1358]), .B(n14648), .Z(n14649) );
  XNOR U17389 ( .A(b[1358]), .B(n14650), .Z(c[1358]) );
  XNOR U17390 ( .A(a[1358]), .B(n14651), .Z(n14650) );
  IV U17391 ( .A(n14648), .Z(n14651) );
  XOR U17392 ( .A(n14652), .B(n14653), .Z(n14648) );
  ANDN U17393 ( .B(n14654), .A(n14655), .Z(n14652) );
  XNOR U17394 ( .A(b[1357]), .B(n14653), .Z(n14654) );
  XNOR U17395 ( .A(b[1357]), .B(n14655), .Z(c[1357]) );
  XNOR U17396 ( .A(a[1357]), .B(n14656), .Z(n14655) );
  IV U17397 ( .A(n14653), .Z(n14656) );
  XOR U17398 ( .A(n14657), .B(n14658), .Z(n14653) );
  ANDN U17399 ( .B(n14659), .A(n14660), .Z(n14657) );
  XNOR U17400 ( .A(b[1356]), .B(n14658), .Z(n14659) );
  XNOR U17401 ( .A(b[1356]), .B(n14660), .Z(c[1356]) );
  XNOR U17402 ( .A(a[1356]), .B(n14661), .Z(n14660) );
  IV U17403 ( .A(n14658), .Z(n14661) );
  XOR U17404 ( .A(n14662), .B(n14663), .Z(n14658) );
  ANDN U17405 ( .B(n14664), .A(n14665), .Z(n14662) );
  XNOR U17406 ( .A(b[1355]), .B(n14663), .Z(n14664) );
  XNOR U17407 ( .A(b[1355]), .B(n14665), .Z(c[1355]) );
  XNOR U17408 ( .A(a[1355]), .B(n14666), .Z(n14665) );
  IV U17409 ( .A(n14663), .Z(n14666) );
  XOR U17410 ( .A(n14667), .B(n14668), .Z(n14663) );
  ANDN U17411 ( .B(n14669), .A(n14670), .Z(n14667) );
  XNOR U17412 ( .A(b[1354]), .B(n14668), .Z(n14669) );
  XNOR U17413 ( .A(b[1354]), .B(n14670), .Z(c[1354]) );
  XNOR U17414 ( .A(a[1354]), .B(n14671), .Z(n14670) );
  IV U17415 ( .A(n14668), .Z(n14671) );
  XOR U17416 ( .A(n14672), .B(n14673), .Z(n14668) );
  ANDN U17417 ( .B(n14674), .A(n14675), .Z(n14672) );
  XNOR U17418 ( .A(b[1353]), .B(n14673), .Z(n14674) );
  XNOR U17419 ( .A(b[1353]), .B(n14675), .Z(c[1353]) );
  XNOR U17420 ( .A(a[1353]), .B(n14676), .Z(n14675) );
  IV U17421 ( .A(n14673), .Z(n14676) );
  XOR U17422 ( .A(n14677), .B(n14678), .Z(n14673) );
  ANDN U17423 ( .B(n14679), .A(n14680), .Z(n14677) );
  XNOR U17424 ( .A(b[1352]), .B(n14678), .Z(n14679) );
  XNOR U17425 ( .A(b[1352]), .B(n14680), .Z(c[1352]) );
  XNOR U17426 ( .A(a[1352]), .B(n14681), .Z(n14680) );
  IV U17427 ( .A(n14678), .Z(n14681) );
  XOR U17428 ( .A(n14682), .B(n14683), .Z(n14678) );
  ANDN U17429 ( .B(n14684), .A(n14685), .Z(n14682) );
  XNOR U17430 ( .A(b[1351]), .B(n14683), .Z(n14684) );
  XNOR U17431 ( .A(b[1351]), .B(n14685), .Z(c[1351]) );
  XNOR U17432 ( .A(a[1351]), .B(n14686), .Z(n14685) );
  IV U17433 ( .A(n14683), .Z(n14686) );
  XOR U17434 ( .A(n14687), .B(n14688), .Z(n14683) );
  ANDN U17435 ( .B(n14689), .A(n14690), .Z(n14687) );
  XNOR U17436 ( .A(b[1350]), .B(n14688), .Z(n14689) );
  XNOR U17437 ( .A(b[1350]), .B(n14690), .Z(c[1350]) );
  XNOR U17438 ( .A(a[1350]), .B(n14691), .Z(n14690) );
  IV U17439 ( .A(n14688), .Z(n14691) );
  XOR U17440 ( .A(n14692), .B(n14693), .Z(n14688) );
  ANDN U17441 ( .B(n14694), .A(n14695), .Z(n14692) );
  XNOR U17442 ( .A(b[1349]), .B(n14693), .Z(n14694) );
  XNOR U17443 ( .A(b[134]), .B(n14696), .Z(c[134]) );
  XNOR U17444 ( .A(b[1349]), .B(n14695), .Z(c[1349]) );
  XNOR U17445 ( .A(a[1349]), .B(n14697), .Z(n14695) );
  IV U17446 ( .A(n14693), .Z(n14697) );
  XOR U17447 ( .A(n14698), .B(n14699), .Z(n14693) );
  ANDN U17448 ( .B(n14700), .A(n14701), .Z(n14698) );
  XNOR U17449 ( .A(b[1348]), .B(n14699), .Z(n14700) );
  XNOR U17450 ( .A(b[1348]), .B(n14701), .Z(c[1348]) );
  XNOR U17451 ( .A(a[1348]), .B(n14702), .Z(n14701) );
  IV U17452 ( .A(n14699), .Z(n14702) );
  XOR U17453 ( .A(n14703), .B(n14704), .Z(n14699) );
  ANDN U17454 ( .B(n14705), .A(n14706), .Z(n14703) );
  XNOR U17455 ( .A(b[1347]), .B(n14704), .Z(n14705) );
  XNOR U17456 ( .A(b[1347]), .B(n14706), .Z(c[1347]) );
  XNOR U17457 ( .A(a[1347]), .B(n14707), .Z(n14706) );
  IV U17458 ( .A(n14704), .Z(n14707) );
  XOR U17459 ( .A(n14708), .B(n14709), .Z(n14704) );
  ANDN U17460 ( .B(n14710), .A(n14711), .Z(n14708) );
  XNOR U17461 ( .A(b[1346]), .B(n14709), .Z(n14710) );
  XNOR U17462 ( .A(b[1346]), .B(n14711), .Z(c[1346]) );
  XNOR U17463 ( .A(a[1346]), .B(n14712), .Z(n14711) );
  IV U17464 ( .A(n14709), .Z(n14712) );
  XOR U17465 ( .A(n14713), .B(n14714), .Z(n14709) );
  ANDN U17466 ( .B(n14715), .A(n14716), .Z(n14713) );
  XNOR U17467 ( .A(b[1345]), .B(n14714), .Z(n14715) );
  XNOR U17468 ( .A(b[1345]), .B(n14716), .Z(c[1345]) );
  XNOR U17469 ( .A(a[1345]), .B(n14717), .Z(n14716) );
  IV U17470 ( .A(n14714), .Z(n14717) );
  XOR U17471 ( .A(n14718), .B(n14719), .Z(n14714) );
  ANDN U17472 ( .B(n14720), .A(n14721), .Z(n14718) );
  XNOR U17473 ( .A(b[1344]), .B(n14719), .Z(n14720) );
  XNOR U17474 ( .A(b[1344]), .B(n14721), .Z(c[1344]) );
  XNOR U17475 ( .A(a[1344]), .B(n14722), .Z(n14721) );
  IV U17476 ( .A(n14719), .Z(n14722) );
  XOR U17477 ( .A(n14723), .B(n14724), .Z(n14719) );
  ANDN U17478 ( .B(n14725), .A(n14726), .Z(n14723) );
  XNOR U17479 ( .A(b[1343]), .B(n14724), .Z(n14725) );
  XNOR U17480 ( .A(b[1343]), .B(n14726), .Z(c[1343]) );
  XNOR U17481 ( .A(a[1343]), .B(n14727), .Z(n14726) );
  IV U17482 ( .A(n14724), .Z(n14727) );
  XOR U17483 ( .A(n14728), .B(n14729), .Z(n14724) );
  ANDN U17484 ( .B(n14730), .A(n14731), .Z(n14728) );
  XNOR U17485 ( .A(b[1342]), .B(n14729), .Z(n14730) );
  XNOR U17486 ( .A(b[1342]), .B(n14731), .Z(c[1342]) );
  XNOR U17487 ( .A(a[1342]), .B(n14732), .Z(n14731) );
  IV U17488 ( .A(n14729), .Z(n14732) );
  XOR U17489 ( .A(n14733), .B(n14734), .Z(n14729) );
  ANDN U17490 ( .B(n14735), .A(n14736), .Z(n14733) );
  XNOR U17491 ( .A(b[1341]), .B(n14734), .Z(n14735) );
  XNOR U17492 ( .A(b[1341]), .B(n14736), .Z(c[1341]) );
  XNOR U17493 ( .A(a[1341]), .B(n14737), .Z(n14736) );
  IV U17494 ( .A(n14734), .Z(n14737) );
  XOR U17495 ( .A(n14738), .B(n14739), .Z(n14734) );
  ANDN U17496 ( .B(n14740), .A(n14741), .Z(n14738) );
  XNOR U17497 ( .A(b[1340]), .B(n14739), .Z(n14740) );
  XNOR U17498 ( .A(b[1340]), .B(n14741), .Z(c[1340]) );
  XNOR U17499 ( .A(a[1340]), .B(n14742), .Z(n14741) );
  IV U17500 ( .A(n14739), .Z(n14742) );
  XOR U17501 ( .A(n14743), .B(n14744), .Z(n14739) );
  ANDN U17502 ( .B(n14745), .A(n14746), .Z(n14743) );
  XNOR U17503 ( .A(b[1339]), .B(n14744), .Z(n14745) );
  XNOR U17504 ( .A(b[133]), .B(n14747), .Z(c[133]) );
  XNOR U17505 ( .A(b[1339]), .B(n14746), .Z(c[1339]) );
  XNOR U17506 ( .A(a[1339]), .B(n14748), .Z(n14746) );
  IV U17507 ( .A(n14744), .Z(n14748) );
  XOR U17508 ( .A(n14749), .B(n14750), .Z(n14744) );
  ANDN U17509 ( .B(n14751), .A(n14752), .Z(n14749) );
  XNOR U17510 ( .A(b[1338]), .B(n14750), .Z(n14751) );
  XNOR U17511 ( .A(b[1338]), .B(n14752), .Z(c[1338]) );
  XNOR U17512 ( .A(a[1338]), .B(n14753), .Z(n14752) );
  IV U17513 ( .A(n14750), .Z(n14753) );
  XOR U17514 ( .A(n14754), .B(n14755), .Z(n14750) );
  ANDN U17515 ( .B(n14756), .A(n14757), .Z(n14754) );
  XNOR U17516 ( .A(b[1337]), .B(n14755), .Z(n14756) );
  XNOR U17517 ( .A(b[1337]), .B(n14757), .Z(c[1337]) );
  XNOR U17518 ( .A(a[1337]), .B(n14758), .Z(n14757) );
  IV U17519 ( .A(n14755), .Z(n14758) );
  XOR U17520 ( .A(n14759), .B(n14760), .Z(n14755) );
  ANDN U17521 ( .B(n14761), .A(n14762), .Z(n14759) );
  XNOR U17522 ( .A(b[1336]), .B(n14760), .Z(n14761) );
  XNOR U17523 ( .A(b[1336]), .B(n14762), .Z(c[1336]) );
  XNOR U17524 ( .A(a[1336]), .B(n14763), .Z(n14762) );
  IV U17525 ( .A(n14760), .Z(n14763) );
  XOR U17526 ( .A(n14764), .B(n14765), .Z(n14760) );
  ANDN U17527 ( .B(n14766), .A(n14767), .Z(n14764) );
  XNOR U17528 ( .A(b[1335]), .B(n14765), .Z(n14766) );
  XNOR U17529 ( .A(b[1335]), .B(n14767), .Z(c[1335]) );
  XNOR U17530 ( .A(a[1335]), .B(n14768), .Z(n14767) );
  IV U17531 ( .A(n14765), .Z(n14768) );
  XOR U17532 ( .A(n14769), .B(n14770), .Z(n14765) );
  ANDN U17533 ( .B(n14771), .A(n14772), .Z(n14769) );
  XNOR U17534 ( .A(b[1334]), .B(n14770), .Z(n14771) );
  XNOR U17535 ( .A(b[1334]), .B(n14772), .Z(c[1334]) );
  XNOR U17536 ( .A(a[1334]), .B(n14773), .Z(n14772) );
  IV U17537 ( .A(n14770), .Z(n14773) );
  XOR U17538 ( .A(n14774), .B(n14775), .Z(n14770) );
  ANDN U17539 ( .B(n14776), .A(n14777), .Z(n14774) );
  XNOR U17540 ( .A(b[1333]), .B(n14775), .Z(n14776) );
  XNOR U17541 ( .A(b[1333]), .B(n14777), .Z(c[1333]) );
  XNOR U17542 ( .A(a[1333]), .B(n14778), .Z(n14777) );
  IV U17543 ( .A(n14775), .Z(n14778) );
  XOR U17544 ( .A(n14779), .B(n14780), .Z(n14775) );
  ANDN U17545 ( .B(n14781), .A(n14782), .Z(n14779) );
  XNOR U17546 ( .A(b[1332]), .B(n14780), .Z(n14781) );
  XNOR U17547 ( .A(b[1332]), .B(n14782), .Z(c[1332]) );
  XNOR U17548 ( .A(a[1332]), .B(n14783), .Z(n14782) );
  IV U17549 ( .A(n14780), .Z(n14783) );
  XOR U17550 ( .A(n14784), .B(n14785), .Z(n14780) );
  ANDN U17551 ( .B(n14786), .A(n14787), .Z(n14784) );
  XNOR U17552 ( .A(b[1331]), .B(n14785), .Z(n14786) );
  XNOR U17553 ( .A(b[1331]), .B(n14787), .Z(c[1331]) );
  XNOR U17554 ( .A(a[1331]), .B(n14788), .Z(n14787) );
  IV U17555 ( .A(n14785), .Z(n14788) );
  XOR U17556 ( .A(n14789), .B(n14790), .Z(n14785) );
  ANDN U17557 ( .B(n14791), .A(n14792), .Z(n14789) );
  XNOR U17558 ( .A(b[1330]), .B(n14790), .Z(n14791) );
  XNOR U17559 ( .A(b[1330]), .B(n14792), .Z(c[1330]) );
  XNOR U17560 ( .A(a[1330]), .B(n14793), .Z(n14792) );
  IV U17561 ( .A(n14790), .Z(n14793) );
  XOR U17562 ( .A(n14794), .B(n14795), .Z(n14790) );
  ANDN U17563 ( .B(n14796), .A(n14797), .Z(n14794) );
  XNOR U17564 ( .A(b[1329]), .B(n14795), .Z(n14796) );
  XNOR U17565 ( .A(b[132]), .B(n14798), .Z(c[132]) );
  XNOR U17566 ( .A(b[1329]), .B(n14797), .Z(c[1329]) );
  XNOR U17567 ( .A(a[1329]), .B(n14799), .Z(n14797) );
  IV U17568 ( .A(n14795), .Z(n14799) );
  XOR U17569 ( .A(n14800), .B(n14801), .Z(n14795) );
  ANDN U17570 ( .B(n14802), .A(n14803), .Z(n14800) );
  XNOR U17571 ( .A(b[1328]), .B(n14801), .Z(n14802) );
  XNOR U17572 ( .A(b[1328]), .B(n14803), .Z(c[1328]) );
  XNOR U17573 ( .A(a[1328]), .B(n14804), .Z(n14803) );
  IV U17574 ( .A(n14801), .Z(n14804) );
  XOR U17575 ( .A(n14805), .B(n14806), .Z(n14801) );
  ANDN U17576 ( .B(n14807), .A(n14808), .Z(n14805) );
  XNOR U17577 ( .A(b[1327]), .B(n14806), .Z(n14807) );
  XNOR U17578 ( .A(b[1327]), .B(n14808), .Z(c[1327]) );
  XNOR U17579 ( .A(a[1327]), .B(n14809), .Z(n14808) );
  IV U17580 ( .A(n14806), .Z(n14809) );
  XOR U17581 ( .A(n14810), .B(n14811), .Z(n14806) );
  ANDN U17582 ( .B(n14812), .A(n14813), .Z(n14810) );
  XNOR U17583 ( .A(b[1326]), .B(n14811), .Z(n14812) );
  XNOR U17584 ( .A(b[1326]), .B(n14813), .Z(c[1326]) );
  XNOR U17585 ( .A(a[1326]), .B(n14814), .Z(n14813) );
  IV U17586 ( .A(n14811), .Z(n14814) );
  XOR U17587 ( .A(n14815), .B(n14816), .Z(n14811) );
  ANDN U17588 ( .B(n14817), .A(n14818), .Z(n14815) );
  XNOR U17589 ( .A(b[1325]), .B(n14816), .Z(n14817) );
  XNOR U17590 ( .A(b[1325]), .B(n14818), .Z(c[1325]) );
  XNOR U17591 ( .A(a[1325]), .B(n14819), .Z(n14818) );
  IV U17592 ( .A(n14816), .Z(n14819) );
  XOR U17593 ( .A(n14820), .B(n14821), .Z(n14816) );
  ANDN U17594 ( .B(n14822), .A(n14823), .Z(n14820) );
  XNOR U17595 ( .A(b[1324]), .B(n14821), .Z(n14822) );
  XNOR U17596 ( .A(b[1324]), .B(n14823), .Z(c[1324]) );
  XNOR U17597 ( .A(a[1324]), .B(n14824), .Z(n14823) );
  IV U17598 ( .A(n14821), .Z(n14824) );
  XOR U17599 ( .A(n14825), .B(n14826), .Z(n14821) );
  ANDN U17600 ( .B(n14827), .A(n14828), .Z(n14825) );
  XNOR U17601 ( .A(b[1323]), .B(n14826), .Z(n14827) );
  XNOR U17602 ( .A(b[1323]), .B(n14828), .Z(c[1323]) );
  XNOR U17603 ( .A(a[1323]), .B(n14829), .Z(n14828) );
  IV U17604 ( .A(n14826), .Z(n14829) );
  XOR U17605 ( .A(n14830), .B(n14831), .Z(n14826) );
  ANDN U17606 ( .B(n14832), .A(n14833), .Z(n14830) );
  XNOR U17607 ( .A(b[1322]), .B(n14831), .Z(n14832) );
  XNOR U17608 ( .A(b[1322]), .B(n14833), .Z(c[1322]) );
  XNOR U17609 ( .A(a[1322]), .B(n14834), .Z(n14833) );
  IV U17610 ( .A(n14831), .Z(n14834) );
  XOR U17611 ( .A(n14835), .B(n14836), .Z(n14831) );
  ANDN U17612 ( .B(n14837), .A(n14838), .Z(n14835) );
  XNOR U17613 ( .A(b[1321]), .B(n14836), .Z(n14837) );
  XNOR U17614 ( .A(b[1321]), .B(n14838), .Z(c[1321]) );
  XNOR U17615 ( .A(a[1321]), .B(n14839), .Z(n14838) );
  IV U17616 ( .A(n14836), .Z(n14839) );
  XOR U17617 ( .A(n14840), .B(n14841), .Z(n14836) );
  ANDN U17618 ( .B(n14842), .A(n14843), .Z(n14840) );
  XNOR U17619 ( .A(b[1320]), .B(n14841), .Z(n14842) );
  XNOR U17620 ( .A(b[1320]), .B(n14843), .Z(c[1320]) );
  XNOR U17621 ( .A(a[1320]), .B(n14844), .Z(n14843) );
  IV U17622 ( .A(n14841), .Z(n14844) );
  XOR U17623 ( .A(n14845), .B(n14846), .Z(n14841) );
  ANDN U17624 ( .B(n14847), .A(n14848), .Z(n14845) );
  XNOR U17625 ( .A(b[1319]), .B(n14846), .Z(n14847) );
  XNOR U17626 ( .A(b[131]), .B(n14849), .Z(c[131]) );
  XNOR U17627 ( .A(b[1319]), .B(n14848), .Z(c[1319]) );
  XNOR U17628 ( .A(a[1319]), .B(n14850), .Z(n14848) );
  IV U17629 ( .A(n14846), .Z(n14850) );
  XOR U17630 ( .A(n14851), .B(n14852), .Z(n14846) );
  ANDN U17631 ( .B(n14853), .A(n14854), .Z(n14851) );
  XNOR U17632 ( .A(b[1318]), .B(n14852), .Z(n14853) );
  XNOR U17633 ( .A(b[1318]), .B(n14854), .Z(c[1318]) );
  XNOR U17634 ( .A(a[1318]), .B(n14855), .Z(n14854) );
  IV U17635 ( .A(n14852), .Z(n14855) );
  XOR U17636 ( .A(n14856), .B(n14857), .Z(n14852) );
  ANDN U17637 ( .B(n14858), .A(n14859), .Z(n14856) );
  XNOR U17638 ( .A(b[1317]), .B(n14857), .Z(n14858) );
  XNOR U17639 ( .A(b[1317]), .B(n14859), .Z(c[1317]) );
  XNOR U17640 ( .A(a[1317]), .B(n14860), .Z(n14859) );
  IV U17641 ( .A(n14857), .Z(n14860) );
  XOR U17642 ( .A(n14861), .B(n14862), .Z(n14857) );
  ANDN U17643 ( .B(n14863), .A(n14864), .Z(n14861) );
  XNOR U17644 ( .A(b[1316]), .B(n14862), .Z(n14863) );
  XNOR U17645 ( .A(b[1316]), .B(n14864), .Z(c[1316]) );
  XNOR U17646 ( .A(a[1316]), .B(n14865), .Z(n14864) );
  IV U17647 ( .A(n14862), .Z(n14865) );
  XOR U17648 ( .A(n14866), .B(n14867), .Z(n14862) );
  ANDN U17649 ( .B(n14868), .A(n14869), .Z(n14866) );
  XNOR U17650 ( .A(b[1315]), .B(n14867), .Z(n14868) );
  XNOR U17651 ( .A(b[1315]), .B(n14869), .Z(c[1315]) );
  XNOR U17652 ( .A(a[1315]), .B(n14870), .Z(n14869) );
  IV U17653 ( .A(n14867), .Z(n14870) );
  XOR U17654 ( .A(n14871), .B(n14872), .Z(n14867) );
  ANDN U17655 ( .B(n14873), .A(n14874), .Z(n14871) );
  XNOR U17656 ( .A(b[1314]), .B(n14872), .Z(n14873) );
  XNOR U17657 ( .A(b[1314]), .B(n14874), .Z(c[1314]) );
  XNOR U17658 ( .A(a[1314]), .B(n14875), .Z(n14874) );
  IV U17659 ( .A(n14872), .Z(n14875) );
  XOR U17660 ( .A(n14876), .B(n14877), .Z(n14872) );
  ANDN U17661 ( .B(n14878), .A(n14879), .Z(n14876) );
  XNOR U17662 ( .A(b[1313]), .B(n14877), .Z(n14878) );
  XNOR U17663 ( .A(b[1313]), .B(n14879), .Z(c[1313]) );
  XNOR U17664 ( .A(a[1313]), .B(n14880), .Z(n14879) );
  IV U17665 ( .A(n14877), .Z(n14880) );
  XOR U17666 ( .A(n14881), .B(n14882), .Z(n14877) );
  ANDN U17667 ( .B(n14883), .A(n14884), .Z(n14881) );
  XNOR U17668 ( .A(b[1312]), .B(n14882), .Z(n14883) );
  XNOR U17669 ( .A(b[1312]), .B(n14884), .Z(c[1312]) );
  XNOR U17670 ( .A(a[1312]), .B(n14885), .Z(n14884) );
  IV U17671 ( .A(n14882), .Z(n14885) );
  XOR U17672 ( .A(n14886), .B(n14887), .Z(n14882) );
  ANDN U17673 ( .B(n14888), .A(n14889), .Z(n14886) );
  XNOR U17674 ( .A(b[1311]), .B(n14887), .Z(n14888) );
  XNOR U17675 ( .A(b[1311]), .B(n14889), .Z(c[1311]) );
  XNOR U17676 ( .A(a[1311]), .B(n14890), .Z(n14889) );
  IV U17677 ( .A(n14887), .Z(n14890) );
  XOR U17678 ( .A(n14891), .B(n14892), .Z(n14887) );
  ANDN U17679 ( .B(n14893), .A(n14894), .Z(n14891) );
  XNOR U17680 ( .A(b[1310]), .B(n14892), .Z(n14893) );
  XNOR U17681 ( .A(b[1310]), .B(n14894), .Z(c[1310]) );
  XNOR U17682 ( .A(a[1310]), .B(n14895), .Z(n14894) );
  IV U17683 ( .A(n14892), .Z(n14895) );
  XOR U17684 ( .A(n14896), .B(n14897), .Z(n14892) );
  ANDN U17685 ( .B(n14898), .A(n14899), .Z(n14896) );
  XNOR U17686 ( .A(b[1309]), .B(n14897), .Z(n14898) );
  XNOR U17687 ( .A(b[130]), .B(n14900), .Z(c[130]) );
  XNOR U17688 ( .A(b[1309]), .B(n14899), .Z(c[1309]) );
  XNOR U17689 ( .A(a[1309]), .B(n14901), .Z(n14899) );
  IV U17690 ( .A(n14897), .Z(n14901) );
  XOR U17691 ( .A(n14902), .B(n14903), .Z(n14897) );
  ANDN U17692 ( .B(n14904), .A(n14905), .Z(n14902) );
  XNOR U17693 ( .A(b[1308]), .B(n14903), .Z(n14904) );
  XNOR U17694 ( .A(b[1308]), .B(n14905), .Z(c[1308]) );
  XNOR U17695 ( .A(a[1308]), .B(n14906), .Z(n14905) );
  IV U17696 ( .A(n14903), .Z(n14906) );
  XOR U17697 ( .A(n14907), .B(n14908), .Z(n14903) );
  ANDN U17698 ( .B(n14909), .A(n14910), .Z(n14907) );
  XNOR U17699 ( .A(b[1307]), .B(n14908), .Z(n14909) );
  XNOR U17700 ( .A(b[1307]), .B(n14910), .Z(c[1307]) );
  XNOR U17701 ( .A(a[1307]), .B(n14911), .Z(n14910) );
  IV U17702 ( .A(n14908), .Z(n14911) );
  XOR U17703 ( .A(n14912), .B(n14913), .Z(n14908) );
  ANDN U17704 ( .B(n14914), .A(n14915), .Z(n14912) );
  XNOR U17705 ( .A(b[1306]), .B(n14913), .Z(n14914) );
  XNOR U17706 ( .A(b[1306]), .B(n14915), .Z(c[1306]) );
  XNOR U17707 ( .A(a[1306]), .B(n14916), .Z(n14915) );
  IV U17708 ( .A(n14913), .Z(n14916) );
  XOR U17709 ( .A(n14917), .B(n14918), .Z(n14913) );
  ANDN U17710 ( .B(n14919), .A(n14920), .Z(n14917) );
  XNOR U17711 ( .A(b[1305]), .B(n14918), .Z(n14919) );
  XNOR U17712 ( .A(b[1305]), .B(n14920), .Z(c[1305]) );
  XNOR U17713 ( .A(a[1305]), .B(n14921), .Z(n14920) );
  IV U17714 ( .A(n14918), .Z(n14921) );
  XOR U17715 ( .A(n14922), .B(n14923), .Z(n14918) );
  ANDN U17716 ( .B(n14924), .A(n14925), .Z(n14922) );
  XNOR U17717 ( .A(b[1304]), .B(n14923), .Z(n14924) );
  XNOR U17718 ( .A(b[1304]), .B(n14925), .Z(c[1304]) );
  XNOR U17719 ( .A(a[1304]), .B(n14926), .Z(n14925) );
  IV U17720 ( .A(n14923), .Z(n14926) );
  XOR U17721 ( .A(n14927), .B(n14928), .Z(n14923) );
  ANDN U17722 ( .B(n14929), .A(n14930), .Z(n14927) );
  XNOR U17723 ( .A(b[1303]), .B(n14928), .Z(n14929) );
  XNOR U17724 ( .A(b[1303]), .B(n14930), .Z(c[1303]) );
  XNOR U17725 ( .A(a[1303]), .B(n14931), .Z(n14930) );
  IV U17726 ( .A(n14928), .Z(n14931) );
  XOR U17727 ( .A(n14932), .B(n14933), .Z(n14928) );
  ANDN U17728 ( .B(n14934), .A(n14935), .Z(n14932) );
  XNOR U17729 ( .A(b[1302]), .B(n14933), .Z(n14934) );
  XNOR U17730 ( .A(b[1302]), .B(n14935), .Z(c[1302]) );
  XNOR U17731 ( .A(a[1302]), .B(n14936), .Z(n14935) );
  IV U17732 ( .A(n14933), .Z(n14936) );
  XOR U17733 ( .A(n14937), .B(n14938), .Z(n14933) );
  ANDN U17734 ( .B(n14939), .A(n14940), .Z(n14937) );
  XNOR U17735 ( .A(b[1301]), .B(n14938), .Z(n14939) );
  XNOR U17736 ( .A(b[1301]), .B(n14940), .Z(c[1301]) );
  XNOR U17737 ( .A(a[1301]), .B(n14941), .Z(n14940) );
  IV U17738 ( .A(n14938), .Z(n14941) );
  XOR U17739 ( .A(n14942), .B(n14943), .Z(n14938) );
  ANDN U17740 ( .B(n14944), .A(n14945), .Z(n14942) );
  XNOR U17741 ( .A(b[1300]), .B(n14943), .Z(n14944) );
  XNOR U17742 ( .A(b[1300]), .B(n14945), .Z(c[1300]) );
  XNOR U17743 ( .A(a[1300]), .B(n14946), .Z(n14945) );
  IV U17744 ( .A(n14943), .Z(n14946) );
  XOR U17745 ( .A(n14947), .B(n14948), .Z(n14943) );
  ANDN U17746 ( .B(n14949), .A(n14950), .Z(n14947) );
  XNOR U17747 ( .A(b[1299]), .B(n14948), .Z(n14949) );
  XNOR U17748 ( .A(b[12]), .B(n14951), .Z(c[12]) );
  XNOR U17749 ( .A(b[129]), .B(n14952), .Z(c[129]) );
  XNOR U17750 ( .A(b[1299]), .B(n14950), .Z(c[1299]) );
  XNOR U17751 ( .A(a[1299]), .B(n14953), .Z(n14950) );
  IV U17752 ( .A(n14948), .Z(n14953) );
  XOR U17753 ( .A(n14954), .B(n14955), .Z(n14948) );
  ANDN U17754 ( .B(n14956), .A(n14957), .Z(n14954) );
  XNOR U17755 ( .A(b[1298]), .B(n14955), .Z(n14956) );
  XNOR U17756 ( .A(b[1298]), .B(n14957), .Z(c[1298]) );
  XNOR U17757 ( .A(a[1298]), .B(n14958), .Z(n14957) );
  IV U17758 ( .A(n14955), .Z(n14958) );
  XOR U17759 ( .A(n14959), .B(n14960), .Z(n14955) );
  ANDN U17760 ( .B(n14961), .A(n14962), .Z(n14959) );
  XNOR U17761 ( .A(b[1297]), .B(n14960), .Z(n14961) );
  XNOR U17762 ( .A(b[1297]), .B(n14962), .Z(c[1297]) );
  XNOR U17763 ( .A(a[1297]), .B(n14963), .Z(n14962) );
  IV U17764 ( .A(n14960), .Z(n14963) );
  XOR U17765 ( .A(n14964), .B(n14965), .Z(n14960) );
  ANDN U17766 ( .B(n14966), .A(n14967), .Z(n14964) );
  XNOR U17767 ( .A(b[1296]), .B(n14965), .Z(n14966) );
  XNOR U17768 ( .A(b[1296]), .B(n14967), .Z(c[1296]) );
  XNOR U17769 ( .A(a[1296]), .B(n14968), .Z(n14967) );
  IV U17770 ( .A(n14965), .Z(n14968) );
  XOR U17771 ( .A(n14969), .B(n14970), .Z(n14965) );
  ANDN U17772 ( .B(n14971), .A(n14972), .Z(n14969) );
  XNOR U17773 ( .A(b[1295]), .B(n14970), .Z(n14971) );
  XNOR U17774 ( .A(b[1295]), .B(n14972), .Z(c[1295]) );
  XNOR U17775 ( .A(a[1295]), .B(n14973), .Z(n14972) );
  IV U17776 ( .A(n14970), .Z(n14973) );
  XOR U17777 ( .A(n14974), .B(n14975), .Z(n14970) );
  ANDN U17778 ( .B(n14976), .A(n14977), .Z(n14974) );
  XNOR U17779 ( .A(b[1294]), .B(n14975), .Z(n14976) );
  XNOR U17780 ( .A(b[1294]), .B(n14977), .Z(c[1294]) );
  XNOR U17781 ( .A(a[1294]), .B(n14978), .Z(n14977) );
  IV U17782 ( .A(n14975), .Z(n14978) );
  XOR U17783 ( .A(n14979), .B(n14980), .Z(n14975) );
  ANDN U17784 ( .B(n14981), .A(n14982), .Z(n14979) );
  XNOR U17785 ( .A(b[1293]), .B(n14980), .Z(n14981) );
  XNOR U17786 ( .A(b[1293]), .B(n14982), .Z(c[1293]) );
  XNOR U17787 ( .A(a[1293]), .B(n14983), .Z(n14982) );
  IV U17788 ( .A(n14980), .Z(n14983) );
  XOR U17789 ( .A(n14984), .B(n14985), .Z(n14980) );
  ANDN U17790 ( .B(n14986), .A(n14987), .Z(n14984) );
  XNOR U17791 ( .A(b[1292]), .B(n14985), .Z(n14986) );
  XNOR U17792 ( .A(b[1292]), .B(n14987), .Z(c[1292]) );
  XNOR U17793 ( .A(a[1292]), .B(n14988), .Z(n14987) );
  IV U17794 ( .A(n14985), .Z(n14988) );
  XOR U17795 ( .A(n14989), .B(n14990), .Z(n14985) );
  ANDN U17796 ( .B(n14991), .A(n14992), .Z(n14989) );
  XNOR U17797 ( .A(b[1291]), .B(n14990), .Z(n14991) );
  XNOR U17798 ( .A(b[1291]), .B(n14992), .Z(c[1291]) );
  XNOR U17799 ( .A(a[1291]), .B(n14993), .Z(n14992) );
  IV U17800 ( .A(n14990), .Z(n14993) );
  XOR U17801 ( .A(n14994), .B(n14995), .Z(n14990) );
  ANDN U17802 ( .B(n14996), .A(n14997), .Z(n14994) );
  XNOR U17803 ( .A(b[1290]), .B(n14995), .Z(n14996) );
  XNOR U17804 ( .A(b[1290]), .B(n14997), .Z(c[1290]) );
  XNOR U17805 ( .A(a[1290]), .B(n14998), .Z(n14997) );
  IV U17806 ( .A(n14995), .Z(n14998) );
  XOR U17807 ( .A(n14999), .B(n15000), .Z(n14995) );
  ANDN U17808 ( .B(n15001), .A(n15002), .Z(n14999) );
  XNOR U17809 ( .A(b[1289]), .B(n15000), .Z(n15001) );
  XNOR U17810 ( .A(b[128]), .B(n15003), .Z(c[128]) );
  XNOR U17811 ( .A(b[1289]), .B(n15002), .Z(c[1289]) );
  XNOR U17812 ( .A(a[1289]), .B(n15004), .Z(n15002) );
  IV U17813 ( .A(n15000), .Z(n15004) );
  XOR U17814 ( .A(n15005), .B(n15006), .Z(n15000) );
  ANDN U17815 ( .B(n15007), .A(n15008), .Z(n15005) );
  XNOR U17816 ( .A(b[1288]), .B(n15006), .Z(n15007) );
  XNOR U17817 ( .A(b[1288]), .B(n15008), .Z(c[1288]) );
  XNOR U17818 ( .A(a[1288]), .B(n15009), .Z(n15008) );
  IV U17819 ( .A(n15006), .Z(n15009) );
  XOR U17820 ( .A(n15010), .B(n15011), .Z(n15006) );
  ANDN U17821 ( .B(n15012), .A(n15013), .Z(n15010) );
  XNOR U17822 ( .A(b[1287]), .B(n15011), .Z(n15012) );
  XNOR U17823 ( .A(b[1287]), .B(n15013), .Z(c[1287]) );
  XNOR U17824 ( .A(a[1287]), .B(n15014), .Z(n15013) );
  IV U17825 ( .A(n15011), .Z(n15014) );
  XOR U17826 ( .A(n15015), .B(n15016), .Z(n15011) );
  ANDN U17827 ( .B(n15017), .A(n15018), .Z(n15015) );
  XNOR U17828 ( .A(b[1286]), .B(n15016), .Z(n15017) );
  XNOR U17829 ( .A(b[1286]), .B(n15018), .Z(c[1286]) );
  XNOR U17830 ( .A(a[1286]), .B(n15019), .Z(n15018) );
  IV U17831 ( .A(n15016), .Z(n15019) );
  XOR U17832 ( .A(n15020), .B(n15021), .Z(n15016) );
  ANDN U17833 ( .B(n15022), .A(n15023), .Z(n15020) );
  XNOR U17834 ( .A(b[1285]), .B(n15021), .Z(n15022) );
  XNOR U17835 ( .A(b[1285]), .B(n15023), .Z(c[1285]) );
  XNOR U17836 ( .A(a[1285]), .B(n15024), .Z(n15023) );
  IV U17837 ( .A(n15021), .Z(n15024) );
  XOR U17838 ( .A(n15025), .B(n15026), .Z(n15021) );
  ANDN U17839 ( .B(n15027), .A(n15028), .Z(n15025) );
  XNOR U17840 ( .A(b[1284]), .B(n15026), .Z(n15027) );
  XNOR U17841 ( .A(b[1284]), .B(n15028), .Z(c[1284]) );
  XNOR U17842 ( .A(a[1284]), .B(n15029), .Z(n15028) );
  IV U17843 ( .A(n15026), .Z(n15029) );
  XOR U17844 ( .A(n15030), .B(n15031), .Z(n15026) );
  ANDN U17845 ( .B(n15032), .A(n15033), .Z(n15030) );
  XNOR U17846 ( .A(b[1283]), .B(n15031), .Z(n15032) );
  XNOR U17847 ( .A(b[1283]), .B(n15033), .Z(c[1283]) );
  XNOR U17848 ( .A(a[1283]), .B(n15034), .Z(n15033) );
  IV U17849 ( .A(n15031), .Z(n15034) );
  XOR U17850 ( .A(n15035), .B(n15036), .Z(n15031) );
  ANDN U17851 ( .B(n15037), .A(n15038), .Z(n15035) );
  XNOR U17852 ( .A(b[1282]), .B(n15036), .Z(n15037) );
  XNOR U17853 ( .A(b[1282]), .B(n15038), .Z(c[1282]) );
  XNOR U17854 ( .A(a[1282]), .B(n15039), .Z(n15038) );
  IV U17855 ( .A(n15036), .Z(n15039) );
  XOR U17856 ( .A(n15040), .B(n15041), .Z(n15036) );
  ANDN U17857 ( .B(n15042), .A(n15043), .Z(n15040) );
  XNOR U17858 ( .A(b[1281]), .B(n15041), .Z(n15042) );
  XNOR U17859 ( .A(b[1281]), .B(n15043), .Z(c[1281]) );
  XNOR U17860 ( .A(a[1281]), .B(n15044), .Z(n15043) );
  IV U17861 ( .A(n15041), .Z(n15044) );
  XOR U17862 ( .A(n15045), .B(n15046), .Z(n15041) );
  ANDN U17863 ( .B(n15047), .A(n15048), .Z(n15045) );
  XNOR U17864 ( .A(b[1280]), .B(n15046), .Z(n15047) );
  XNOR U17865 ( .A(b[1280]), .B(n15048), .Z(c[1280]) );
  XNOR U17866 ( .A(a[1280]), .B(n15049), .Z(n15048) );
  IV U17867 ( .A(n15046), .Z(n15049) );
  XOR U17868 ( .A(n15050), .B(n15051), .Z(n15046) );
  ANDN U17869 ( .B(n15052), .A(n15053), .Z(n15050) );
  XNOR U17870 ( .A(b[1279]), .B(n15051), .Z(n15052) );
  XNOR U17871 ( .A(b[127]), .B(n15054), .Z(c[127]) );
  XNOR U17872 ( .A(b[1279]), .B(n15053), .Z(c[1279]) );
  XNOR U17873 ( .A(a[1279]), .B(n15055), .Z(n15053) );
  IV U17874 ( .A(n15051), .Z(n15055) );
  XOR U17875 ( .A(n15056), .B(n15057), .Z(n15051) );
  ANDN U17876 ( .B(n15058), .A(n15059), .Z(n15056) );
  XNOR U17877 ( .A(b[1278]), .B(n15057), .Z(n15058) );
  XNOR U17878 ( .A(b[1278]), .B(n15059), .Z(c[1278]) );
  XNOR U17879 ( .A(a[1278]), .B(n15060), .Z(n15059) );
  IV U17880 ( .A(n15057), .Z(n15060) );
  XOR U17881 ( .A(n15061), .B(n15062), .Z(n15057) );
  ANDN U17882 ( .B(n15063), .A(n15064), .Z(n15061) );
  XNOR U17883 ( .A(b[1277]), .B(n15062), .Z(n15063) );
  XNOR U17884 ( .A(b[1277]), .B(n15064), .Z(c[1277]) );
  XNOR U17885 ( .A(a[1277]), .B(n15065), .Z(n15064) );
  IV U17886 ( .A(n15062), .Z(n15065) );
  XOR U17887 ( .A(n15066), .B(n15067), .Z(n15062) );
  ANDN U17888 ( .B(n15068), .A(n15069), .Z(n15066) );
  XNOR U17889 ( .A(b[1276]), .B(n15067), .Z(n15068) );
  XNOR U17890 ( .A(b[1276]), .B(n15069), .Z(c[1276]) );
  XNOR U17891 ( .A(a[1276]), .B(n15070), .Z(n15069) );
  IV U17892 ( .A(n15067), .Z(n15070) );
  XOR U17893 ( .A(n15071), .B(n15072), .Z(n15067) );
  ANDN U17894 ( .B(n15073), .A(n15074), .Z(n15071) );
  XNOR U17895 ( .A(b[1275]), .B(n15072), .Z(n15073) );
  XNOR U17896 ( .A(b[1275]), .B(n15074), .Z(c[1275]) );
  XNOR U17897 ( .A(a[1275]), .B(n15075), .Z(n15074) );
  IV U17898 ( .A(n15072), .Z(n15075) );
  XOR U17899 ( .A(n15076), .B(n15077), .Z(n15072) );
  ANDN U17900 ( .B(n15078), .A(n15079), .Z(n15076) );
  XNOR U17901 ( .A(b[1274]), .B(n15077), .Z(n15078) );
  XNOR U17902 ( .A(b[1274]), .B(n15079), .Z(c[1274]) );
  XNOR U17903 ( .A(a[1274]), .B(n15080), .Z(n15079) );
  IV U17904 ( .A(n15077), .Z(n15080) );
  XOR U17905 ( .A(n15081), .B(n15082), .Z(n15077) );
  ANDN U17906 ( .B(n15083), .A(n15084), .Z(n15081) );
  XNOR U17907 ( .A(b[1273]), .B(n15082), .Z(n15083) );
  XNOR U17908 ( .A(b[1273]), .B(n15084), .Z(c[1273]) );
  XNOR U17909 ( .A(a[1273]), .B(n15085), .Z(n15084) );
  IV U17910 ( .A(n15082), .Z(n15085) );
  XOR U17911 ( .A(n15086), .B(n15087), .Z(n15082) );
  ANDN U17912 ( .B(n15088), .A(n15089), .Z(n15086) );
  XNOR U17913 ( .A(b[1272]), .B(n15087), .Z(n15088) );
  XNOR U17914 ( .A(b[1272]), .B(n15089), .Z(c[1272]) );
  XNOR U17915 ( .A(a[1272]), .B(n15090), .Z(n15089) );
  IV U17916 ( .A(n15087), .Z(n15090) );
  XOR U17917 ( .A(n15091), .B(n15092), .Z(n15087) );
  ANDN U17918 ( .B(n15093), .A(n15094), .Z(n15091) );
  XNOR U17919 ( .A(b[1271]), .B(n15092), .Z(n15093) );
  XNOR U17920 ( .A(b[1271]), .B(n15094), .Z(c[1271]) );
  XNOR U17921 ( .A(a[1271]), .B(n15095), .Z(n15094) );
  IV U17922 ( .A(n15092), .Z(n15095) );
  XOR U17923 ( .A(n15096), .B(n15097), .Z(n15092) );
  ANDN U17924 ( .B(n15098), .A(n15099), .Z(n15096) );
  XNOR U17925 ( .A(b[1270]), .B(n15097), .Z(n15098) );
  XNOR U17926 ( .A(b[1270]), .B(n15099), .Z(c[1270]) );
  XNOR U17927 ( .A(a[1270]), .B(n15100), .Z(n15099) );
  IV U17928 ( .A(n15097), .Z(n15100) );
  XOR U17929 ( .A(n15101), .B(n15102), .Z(n15097) );
  ANDN U17930 ( .B(n15103), .A(n15104), .Z(n15101) );
  XNOR U17931 ( .A(b[1269]), .B(n15102), .Z(n15103) );
  XNOR U17932 ( .A(b[126]), .B(n15105), .Z(c[126]) );
  XNOR U17933 ( .A(b[1269]), .B(n15104), .Z(c[1269]) );
  XNOR U17934 ( .A(a[1269]), .B(n15106), .Z(n15104) );
  IV U17935 ( .A(n15102), .Z(n15106) );
  XOR U17936 ( .A(n15107), .B(n15108), .Z(n15102) );
  ANDN U17937 ( .B(n15109), .A(n15110), .Z(n15107) );
  XNOR U17938 ( .A(b[1268]), .B(n15108), .Z(n15109) );
  XNOR U17939 ( .A(b[1268]), .B(n15110), .Z(c[1268]) );
  XNOR U17940 ( .A(a[1268]), .B(n15111), .Z(n15110) );
  IV U17941 ( .A(n15108), .Z(n15111) );
  XOR U17942 ( .A(n15112), .B(n15113), .Z(n15108) );
  ANDN U17943 ( .B(n15114), .A(n15115), .Z(n15112) );
  XNOR U17944 ( .A(b[1267]), .B(n15113), .Z(n15114) );
  XNOR U17945 ( .A(b[1267]), .B(n15115), .Z(c[1267]) );
  XNOR U17946 ( .A(a[1267]), .B(n15116), .Z(n15115) );
  IV U17947 ( .A(n15113), .Z(n15116) );
  XOR U17948 ( .A(n15117), .B(n15118), .Z(n15113) );
  ANDN U17949 ( .B(n15119), .A(n15120), .Z(n15117) );
  XNOR U17950 ( .A(b[1266]), .B(n15118), .Z(n15119) );
  XNOR U17951 ( .A(b[1266]), .B(n15120), .Z(c[1266]) );
  XNOR U17952 ( .A(a[1266]), .B(n15121), .Z(n15120) );
  IV U17953 ( .A(n15118), .Z(n15121) );
  XOR U17954 ( .A(n15122), .B(n15123), .Z(n15118) );
  ANDN U17955 ( .B(n15124), .A(n15125), .Z(n15122) );
  XNOR U17956 ( .A(b[1265]), .B(n15123), .Z(n15124) );
  XNOR U17957 ( .A(b[1265]), .B(n15125), .Z(c[1265]) );
  XNOR U17958 ( .A(a[1265]), .B(n15126), .Z(n15125) );
  IV U17959 ( .A(n15123), .Z(n15126) );
  XOR U17960 ( .A(n15127), .B(n15128), .Z(n15123) );
  ANDN U17961 ( .B(n15129), .A(n15130), .Z(n15127) );
  XNOR U17962 ( .A(b[1264]), .B(n15128), .Z(n15129) );
  XNOR U17963 ( .A(b[1264]), .B(n15130), .Z(c[1264]) );
  XNOR U17964 ( .A(a[1264]), .B(n15131), .Z(n15130) );
  IV U17965 ( .A(n15128), .Z(n15131) );
  XOR U17966 ( .A(n15132), .B(n15133), .Z(n15128) );
  ANDN U17967 ( .B(n15134), .A(n15135), .Z(n15132) );
  XNOR U17968 ( .A(b[1263]), .B(n15133), .Z(n15134) );
  XNOR U17969 ( .A(b[1263]), .B(n15135), .Z(c[1263]) );
  XNOR U17970 ( .A(a[1263]), .B(n15136), .Z(n15135) );
  IV U17971 ( .A(n15133), .Z(n15136) );
  XOR U17972 ( .A(n15137), .B(n15138), .Z(n15133) );
  ANDN U17973 ( .B(n15139), .A(n15140), .Z(n15137) );
  XNOR U17974 ( .A(b[1262]), .B(n15138), .Z(n15139) );
  XNOR U17975 ( .A(b[1262]), .B(n15140), .Z(c[1262]) );
  XNOR U17976 ( .A(a[1262]), .B(n15141), .Z(n15140) );
  IV U17977 ( .A(n15138), .Z(n15141) );
  XOR U17978 ( .A(n15142), .B(n15143), .Z(n15138) );
  ANDN U17979 ( .B(n15144), .A(n15145), .Z(n15142) );
  XNOR U17980 ( .A(b[1261]), .B(n15143), .Z(n15144) );
  XNOR U17981 ( .A(b[1261]), .B(n15145), .Z(c[1261]) );
  XNOR U17982 ( .A(a[1261]), .B(n15146), .Z(n15145) );
  IV U17983 ( .A(n15143), .Z(n15146) );
  XOR U17984 ( .A(n15147), .B(n15148), .Z(n15143) );
  ANDN U17985 ( .B(n15149), .A(n15150), .Z(n15147) );
  XNOR U17986 ( .A(b[1260]), .B(n15148), .Z(n15149) );
  XNOR U17987 ( .A(b[1260]), .B(n15150), .Z(c[1260]) );
  XNOR U17988 ( .A(a[1260]), .B(n15151), .Z(n15150) );
  IV U17989 ( .A(n15148), .Z(n15151) );
  XOR U17990 ( .A(n15152), .B(n15153), .Z(n15148) );
  ANDN U17991 ( .B(n15154), .A(n15155), .Z(n15152) );
  XNOR U17992 ( .A(b[1259]), .B(n15153), .Z(n15154) );
  XNOR U17993 ( .A(b[125]), .B(n15156), .Z(c[125]) );
  XNOR U17994 ( .A(b[1259]), .B(n15155), .Z(c[1259]) );
  XNOR U17995 ( .A(a[1259]), .B(n15157), .Z(n15155) );
  IV U17996 ( .A(n15153), .Z(n15157) );
  XOR U17997 ( .A(n15158), .B(n15159), .Z(n15153) );
  ANDN U17998 ( .B(n15160), .A(n15161), .Z(n15158) );
  XNOR U17999 ( .A(b[1258]), .B(n15159), .Z(n15160) );
  XNOR U18000 ( .A(b[1258]), .B(n15161), .Z(c[1258]) );
  XNOR U18001 ( .A(a[1258]), .B(n15162), .Z(n15161) );
  IV U18002 ( .A(n15159), .Z(n15162) );
  XOR U18003 ( .A(n15163), .B(n15164), .Z(n15159) );
  ANDN U18004 ( .B(n15165), .A(n15166), .Z(n15163) );
  XNOR U18005 ( .A(b[1257]), .B(n15164), .Z(n15165) );
  XNOR U18006 ( .A(b[1257]), .B(n15166), .Z(c[1257]) );
  XNOR U18007 ( .A(a[1257]), .B(n15167), .Z(n15166) );
  IV U18008 ( .A(n15164), .Z(n15167) );
  XOR U18009 ( .A(n15168), .B(n15169), .Z(n15164) );
  ANDN U18010 ( .B(n15170), .A(n15171), .Z(n15168) );
  XNOR U18011 ( .A(b[1256]), .B(n15169), .Z(n15170) );
  XNOR U18012 ( .A(b[1256]), .B(n15171), .Z(c[1256]) );
  XNOR U18013 ( .A(a[1256]), .B(n15172), .Z(n15171) );
  IV U18014 ( .A(n15169), .Z(n15172) );
  XOR U18015 ( .A(n15173), .B(n15174), .Z(n15169) );
  ANDN U18016 ( .B(n15175), .A(n15176), .Z(n15173) );
  XNOR U18017 ( .A(b[1255]), .B(n15174), .Z(n15175) );
  XNOR U18018 ( .A(b[1255]), .B(n15176), .Z(c[1255]) );
  XNOR U18019 ( .A(a[1255]), .B(n15177), .Z(n15176) );
  IV U18020 ( .A(n15174), .Z(n15177) );
  XOR U18021 ( .A(n15178), .B(n15179), .Z(n15174) );
  ANDN U18022 ( .B(n15180), .A(n15181), .Z(n15178) );
  XNOR U18023 ( .A(b[1254]), .B(n15179), .Z(n15180) );
  XNOR U18024 ( .A(b[1254]), .B(n15181), .Z(c[1254]) );
  XNOR U18025 ( .A(a[1254]), .B(n15182), .Z(n15181) );
  IV U18026 ( .A(n15179), .Z(n15182) );
  XOR U18027 ( .A(n15183), .B(n15184), .Z(n15179) );
  ANDN U18028 ( .B(n15185), .A(n15186), .Z(n15183) );
  XNOR U18029 ( .A(b[1253]), .B(n15184), .Z(n15185) );
  XNOR U18030 ( .A(b[1253]), .B(n15186), .Z(c[1253]) );
  XNOR U18031 ( .A(a[1253]), .B(n15187), .Z(n15186) );
  IV U18032 ( .A(n15184), .Z(n15187) );
  XOR U18033 ( .A(n15188), .B(n15189), .Z(n15184) );
  ANDN U18034 ( .B(n15190), .A(n15191), .Z(n15188) );
  XNOR U18035 ( .A(b[1252]), .B(n15189), .Z(n15190) );
  XNOR U18036 ( .A(b[1252]), .B(n15191), .Z(c[1252]) );
  XNOR U18037 ( .A(a[1252]), .B(n15192), .Z(n15191) );
  IV U18038 ( .A(n15189), .Z(n15192) );
  XOR U18039 ( .A(n15193), .B(n15194), .Z(n15189) );
  ANDN U18040 ( .B(n15195), .A(n15196), .Z(n15193) );
  XNOR U18041 ( .A(b[1251]), .B(n15194), .Z(n15195) );
  XNOR U18042 ( .A(b[1251]), .B(n15196), .Z(c[1251]) );
  XNOR U18043 ( .A(a[1251]), .B(n15197), .Z(n15196) );
  IV U18044 ( .A(n15194), .Z(n15197) );
  XOR U18045 ( .A(n15198), .B(n15199), .Z(n15194) );
  ANDN U18046 ( .B(n15200), .A(n15201), .Z(n15198) );
  XNOR U18047 ( .A(b[1250]), .B(n15199), .Z(n15200) );
  XNOR U18048 ( .A(b[1250]), .B(n15201), .Z(c[1250]) );
  XNOR U18049 ( .A(a[1250]), .B(n15202), .Z(n15201) );
  IV U18050 ( .A(n15199), .Z(n15202) );
  XOR U18051 ( .A(n15203), .B(n15204), .Z(n15199) );
  ANDN U18052 ( .B(n15205), .A(n15206), .Z(n15203) );
  XNOR U18053 ( .A(b[1249]), .B(n15204), .Z(n15205) );
  XNOR U18054 ( .A(b[124]), .B(n15207), .Z(c[124]) );
  XNOR U18055 ( .A(b[1249]), .B(n15206), .Z(c[1249]) );
  XNOR U18056 ( .A(a[1249]), .B(n15208), .Z(n15206) );
  IV U18057 ( .A(n15204), .Z(n15208) );
  XOR U18058 ( .A(n15209), .B(n15210), .Z(n15204) );
  ANDN U18059 ( .B(n15211), .A(n15212), .Z(n15209) );
  XNOR U18060 ( .A(b[1248]), .B(n15210), .Z(n15211) );
  XNOR U18061 ( .A(b[1248]), .B(n15212), .Z(c[1248]) );
  XNOR U18062 ( .A(a[1248]), .B(n15213), .Z(n15212) );
  IV U18063 ( .A(n15210), .Z(n15213) );
  XOR U18064 ( .A(n15214), .B(n15215), .Z(n15210) );
  ANDN U18065 ( .B(n15216), .A(n15217), .Z(n15214) );
  XNOR U18066 ( .A(b[1247]), .B(n15215), .Z(n15216) );
  XNOR U18067 ( .A(b[1247]), .B(n15217), .Z(c[1247]) );
  XNOR U18068 ( .A(a[1247]), .B(n15218), .Z(n15217) );
  IV U18069 ( .A(n15215), .Z(n15218) );
  XOR U18070 ( .A(n15219), .B(n15220), .Z(n15215) );
  ANDN U18071 ( .B(n15221), .A(n15222), .Z(n15219) );
  XNOR U18072 ( .A(b[1246]), .B(n15220), .Z(n15221) );
  XNOR U18073 ( .A(b[1246]), .B(n15222), .Z(c[1246]) );
  XNOR U18074 ( .A(a[1246]), .B(n15223), .Z(n15222) );
  IV U18075 ( .A(n15220), .Z(n15223) );
  XOR U18076 ( .A(n15224), .B(n15225), .Z(n15220) );
  ANDN U18077 ( .B(n15226), .A(n15227), .Z(n15224) );
  XNOR U18078 ( .A(b[1245]), .B(n15225), .Z(n15226) );
  XNOR U18079 ( .A(b[1245]), .B(n15227), .Z(c[1245]) );
  XNOR U18080 ( .A(a[1245]), .B(n15228), .Z(n15227) );
  IV U18081 ( .A(n15225), .Z(n15228) );
  XOR U18082 ( .A(n15229), .B(n15230), .Z(n15225) );
  ANDN U18083 ( .B(n15231), .A(n15232), .Z(n15229) );
  XNOR U18084 ( .A(b[1244]), .B(n15230), .Z(n15231) );
  XNOR U18085 ( .A(b[1244]), .B(n15232), .Z(c[1244]) );
  XNOR U18086 ( .A(a[1244]), .B(n15233), .Z(n15232) );
  IV U18087 ( .A(n15230), .Z(n15233) );
  XOR U18088 ( .A(n15234), .B(n15235), .Z(n15230) );
  ANDN U18089 ( .B(n15236), .A(n15237), .Z(n15234) );
  XNOR U18090 ( .A(b[1243]), .B(n15235), .Z(n15236) );
  XNOR U18091 ( .A(b[1243]), .B(n15237), .Z(c[1243]) );
  XNOR U18092 ( .A(a[1243]), .B(n15238), .Z(n15237) );
  IV U18093 ( .A(n15235), .Z(n15238) );
  XOR U18094 ( .A(n15239), .B(n15240), .Z(n15235) );
  ANDN U18095 ( .B(n15241), .A(n15242), .Z(n15239) );
  XNOR U18096 ( .A(b[1242]), .B(n15240), .Z(n15241) );
  XNOR U18097 ( .A(b[1242]), .B(n15242), .Z(c[1242]) );
  XNOR U18098 ( .A(a[1242]), .B(n15243), .Z(n15242) );
  IV U18099 ( .A(n15240), .Z(n15243) );
  XOR U18100 ( .A(n15244), .B(n15245), .Z(n15240) );
  ANDN U18101 ( .B(n15246), .A(n15247), .Z(n15244) );
  XNOR U18102 ( .A(b[1241]), .B(n15245), .Z(n15246) );
  XNOR U18103 ( .A(b[1241]), .B(n15247), .Z(c[1241]) );
  XNOR U18104 ( .A(a[1241]), .B(n15248), .Z(n15247) );
  IV U18105 ( .A(n15245), .Z(n15248) );
  XOR U18106 ( .A(n15249), .B(n15250), .Z(n15245) );
  ANDN U18107 ( .B(n15251), .A(n15252), .Z(n15249) );
  XNOR U18108 ( .A(b[1240]), .B(n15250), .Z(n15251) );
  XNOR U18109 ( .A(b[1240]), .B(n15252), .Z(c[1240]) );
  XNOR U18110 ( .A(a[1240]), .B(n15253), .Z(n15252) );
  IV U18111 ( .A(n15250), .Z(n15253) );
  XOR U18112 ( .A(n15254), .B(n15255), .Z(n15250) );
  ANDN U18113 ( .B(n15256), .A(n15257), .Z(n15254) );
  XNOR U18114 ( .A(b[1239]), .B(n15255), .Z(n15256) );
  XNOR U18115 ( .A(b[123]), .B(n15258), .Z(c[123]) );
  XNOR U18116 ( .A(b[1239]), .B(n15257), .Z(c[1239]) );
  XNOR U18117 ( .A(a[1239]), .B(n15259), .Z(n15257) );
  IV U18118 ( .A(n15255), .Z(n15259) );
  XOR U18119 ( .A(n15260), .B(n15261), .Z(n15255) );
  ANDN U18120 ( .B(n15262), .A(n15263), .Z(n15260) );
  XNOR U18121 ( .A(b[1238]), .B(n15261), .Z(n15262) );
  XNOR U18122 ( .A(b[1238]), .B(n15263), .Z(c[1238]) );
  XNOR U18123 ( .A(a[1238]), .B(n15264), .Z(n15263) );
  IV U18124 ( .A(n15261), .Z(n15264) );
  XOR U18125 ( .A(n15265), .B(n15266), .Z(n15261) );
  ANDN U18126 ( .B(n15267), .A(n15268), .Z(n15265) );
  XNOR U18127 ( .A(b[1237]), .B(n15266), .Z(n15267) );
  XNOR U18128 ( .A(b[1237]), .B(n15268), .Z(c[1237]) );
  XNOR U18129 ( .A(a[1237]), .B(n15269), .Z(n15268) );
  IV U18130 ( .A(n15266), .Z(n15269) );
  XOR U18131 ( .A(n15270), .B(n15271), .Z(n15266) );
  ANDN U18132 ( .B(n15272), .A(n15273), .Z(n15270) );
  XNOR U18133 ( .A(b[1236]), .B(n15271), .Z(n15272) );
  XNOR U18134 ( .A(b[1236]), .B(n15273), .Z(c[1236]) );
  XNOR U18135 ( .A(a[1236]), .B(n15274), .Z(n15273) );
  IV U18136 ( .A(n15271), .Z(n15274) );
  XOR U18137 ( .A(n15275), .B(n15276), .Z(n15271) );
  ANDN U18138 ( .B(n15277), .A(n15278), .Z(n15275) );
  XNOR U18139 ( .A(b[1235]), .B(n15276), .Z(n15277) );
  XNOR U18140 ( .A(b[1235]), .B(n15278), .Z(c[1235]) );
  XNOR U18141 ( .A(a[1235]), .B(n15279), .Z(n15278) );
  IV U18142 ( .A(n15276), .Z(n15279) );
  XOR U18143 ( .A(n15280), .B(n15281), .Z(n15276) );
  ANDN U18144 ( .B(n15282), .A(n15283), .Z(n15280) );
  XNOR U18145 ( .A(b[1234]), .B(n15281), .Z(n15282) );
  XNOR U18146 ( .A(b[1234]), .B(n15283), .Z(c[1234]) );
  XNOR U18147 ( .A(a[1234]), .B(n15284), .Z(n15283) );
  IV U18148 ( .A(n15281), .Z(n15284) );
  XOR U18149 ( .A(n15285), .B(n15286), .Z(n15281) );
  ANDN U18150 ( .B(n15287), .A(n15288), .Z(n15285) );
  XNOR U18151 ( .A(b[1233]), .B(n15286), .Z(n15287) );
  XNOR U18152 ( .A(b[1233]), .B(n15288), .Z(c[1233]) );
  XNOR U18153 ( .A(a[1233]), .B(n15289), .Z(n15288) );
  IV U18154 ( .A(n15286), .Z(n15289) );
  XOR U18155 ( .A(n15290), .B(n15291), .Z(n15286) );
  ANDN U18156 ( .B(n15292), .A(n15293), .Z(n15290) );
  XNOR U18157 ( .A(b[1232]), .B(n15291), .Z(n15292) );
  XNOR U18158 ( .A(b[1232]), .B(n15293), .Z(c[1232]) );
  XNOR U18159 ( .A(a[1232]), .B(n15294), .Z(n15293) );
  IV U18160 ( .A(n15291), .Z(n15294) );
  XOR U18161 ( .A(n15295), .B(n15296), .Z(n15291) );
  ANDN U18162 ( .B(n15297), .A(n15298), .Z(n15295) );
  XNOR U18163 ( .A(b[1231]), .B(n15296), .Z(n15297) );
  XNOR U18164 ( .A(b[1231]), .B(n15298), .Z(c[1231]) );
  XNOR U18165 ( .A(a[1231]), .B(n15299), .Z(n15298) );
  IV U18166 ( .A(n15296), .Z(n15299) );
  XOR U18167 ( .A(n15300), .B(n15301), .Z(n15296) );
  ANDN U18168 ( .B(n15302), .A(n15303), .Z(n15300) );
  XNOR U18169 ( .A(b[1230]), .B(n15301), .Z(n15302) );
  XNOR U18170 ( .A(b[1230]), .B(n15303), .Z(c[1230]) );
  XNOR U18171 ( .A(a[1230]), .B(n15304), .Z(n15303) );
  IV U18172 ( .A(n15301), .Z(n15304) );
  XOR U18173 ( .A(n15305), .B(n15306), .Z(n15301) );
  ANDN U18174 ( .B(n15307), .A(n15308), .Z(n15305) );
  XNOR U18175 ( .A(b[1229]), .B(n15306), .Z(n15307) );
  XNOR U18176 ( .A(b[122]), .B(n15309), .Z(c[122]) );
  XNOR U18177 ( .A(b[1229]), .B(n15308), .Z(c[1229]) );
  XNOR U18178 ( .A(a[1229]), .B(n15310), .Z(n15308) );
  IV U18179 ( .A(n15306), .Z(n15310) );
  XOR U18180 ( .A(n15311), .B(n15312), .Z(n15306) );
  ANDN U18181 ( .B(n15313), .A(n15314), .Z(n15311) );
  XNOR U18182 ( .A(b[1228]), .B(n15312), .Z(n15313) );
  XNOR U18183 ( .A(b[1228]), .B(n15314), .Z(c[1228]) );
  XNOR U18184 ( .A(a[1228]), .B(n15315), .Z(n15314) );
  IV U18185 ( .A(n15312), .Z(n15315) );
  XOR U18186 ( .A(n15316), .B(n15317), .Z(n15312) );
  ANDN U18187 ( .B(n15318), .A(n15319), .Z(n15316) );
  XNOR U18188 ( .A(b[1227]), .B(n15317), .Z(n15318) );
  XNOR U18189 ( .A(b[1227]), .B(n15319), .Z(c[1227]) );
  XNOR U18190 ( .A(a[1227]), .B(n15320), .Z(n15319) );
  IV U18191 ( .A(n15317), .Z(n15320) );
  XOR U18192 ( .A(n15321), .B(n15322), .Z(n15317) );
  ANDN U18193 ( .B(n15323), .A(n15324), .Z(n15321) );
  XNOR U18194 ( .A(b[1226]), .B(n15322), .Z(n15323) );
  XNOR U18195 ( .A(b[1226]), .B(n15324), .Z(c[1226]) );
  XNOR U18196 ( .A(a[1226]), .B(n15325), .Z(n15324) );
  IV U18197 ( .A(n15322), .Z(n15325) );
  XOR U18198 ( .A(n15326), .B(n15327), .Z(n15322) );
  ANDN U18199 ( .B(n15328), .A(n15329), .Z(n15326) );
  XNOR U18200 ( .A(b[1225]), .B(n15327), .Z(n15328) );
  XNOR U18201 ( .A(b[1225]), .B(n15329), .Z(c[1225]) );
  XNOR U18202 ( .A(a[1225]), .B(n15330), .Z(n15329) );
  IV U18203 ( .A(n15327), .Z(n15330) );
  XOR U18204 ( .A(n15331), .B(n15332), .Z(n15327) );
  ANDN U18205 ( .B(n15333), .A(n15334), .Z(n15331) );
  XNOR U18206 ( .A(b[1224]), .B(n15332), .Z(n15333) );
  XNOR U18207 ( .A(b[1224]), .B(n15334), .Z(c[1224]) );
  XNOR U18208 ( .A(a[1224]), .B(n15335), .Z(n15334) );
  IV U18209 ( .A(n15332), .Z(n15335) );
  XOR U18210 ( .A(n15336), .B(n15337), .Z(n15332) );
  ANDN U18211 ( .B(n15338), .A(n15339), .Z(n15336) );
  XNOR U18212 ( .A(b[1223]), .B(n15337), .Z(n15338) );
  XNOR U18213 ( .A(b[1223]), .B(n15339), .Z(c[1223]) );
  XNOR U18214 ( .A(a[1223]), .B(n15340), .Z(n15339) );
  IV U18215 ( .A(n15337), .Z(n15340) );
  XOR U18216 ( .A(n15341), .B(n15342), .Z(n15337) );
  ANDN U18217 ( .B(n15343), .A(n15344), .Z(n15341) );
  XNOR U18218 ( .A(b[1222]), .B(n15342), .Z(n15343) );
  XNOR U18219 ( .A(b[1222]), .B(n15344), .Z(c[1222]) );
  XNOR U18220 ( .A(a[1222]), .B(n15345), .Z(n15344) );
  IV U18221 ( .A(n15342), .Z(n15345) );
  XOR U18222 ( .A(n15346), .B(n15347), .Z(n15342) );
  ANDN U18223 ( .B(n15348), .A(n15349), .Z(n15346) );
  XNOR U18224 ( .A(b[1221]), .B(n15347), .Z(n15348) );
  XNOR U18225 ( .A(b[1221]), .B(n15349), .Z(c[1221]) );
  XNOR U18226 ( .A(a[1221]), .B(n15350), .Z(n15349) );
  IV U18227 ( .A(n15347), .Z(n15350) );
  XOR U18228 ( .A(n15351), .B(n15352), .Z(n15347) );
  ANDN U18229 ( .B(n15353), .A(n15354), .Z(n15351) );
  XNOR U18230 ( .A(b[1220]), .B(n15352), .Z(n15353) );
  XNOR U18231 ( .A(b[1220]), .B(n15354), .Z(c[1220]) );
  XNOR U18232 ( .A(a[1220]), .B(n15355), .Z(n15354) );
  IV U18233 ( .A(n15352), .Z(n15355) );
  XOR U18234 ( .A(n15356), .B(n15357), .Z(n15352) );
  ANDN U18235 ( .B(n15358), .A(n15359), .Z(n15356) );
  XNOR U18236 ( .A(b[1219]), .B(n15357), .Z(n15358) );
  XNOR U18237 ( .A(b[121]), .B(n15360), .Z(c[121]) );
  XNOR U18238 ( .A(b[1219]), .B(n15359), .Z(c[1219]) );
  XNOR U18239 ( .A(a[1219]), .B(n15361), .Z(n15359) );
  IV U18240 ( .A(n15357), .Z(n15361) );
  XOR U18241 ( .A(n15362), .B(n15363), .Z(n15357) );
  ANDN U18242 ( .B(n15364), .A(n15365), .Z(n15362) );
  XNOR U18243 ( .A(b[1218]), .B(n15363), .Z(n15364) );
  XNOR U18244 ( .A(b[1218]), .B(n15365), .Z(c[1218]) );
  XNOR U18245 ( .A(a[1218]), .B(n15366), .Z(n15365) );
  IV U18246 ( .A(n15363), .Z(n15366) );
  XOR U18247 ( .A(n15367), .B(n15368), .Z(n15363) );
  ANDN U18248 ( .B(n15369), .A(n15370), .Z(n15367) );
  XNOR U18249 ( .A(b[1217]), .B(n15368), .Z(n15369) );
  XNOR U18250 ( .A(b[1217]), .B(n15370), .Z(c[1217]) );
  XNOR U18251 ( .A(a[1217]), .B(n15371), .Z(n15370) );
  IV U18252 ( .A(n15368), .Z(n15371) );
  XOR U18253 ( .A(n15372), .B(n15373), .Z(n15368) );
  ANDN U18254 ( .B(n15374), .A(n15375), .Z(n15372) );
  XNOR U18255 ( .A(b[1216]), .B(n15373), .Z(n15374) );
  XNOR U18256 ( .A(b[1216]), .B(n15375), .Z(c[1216]) );
  XNOR U18257 ( .A(a[1216]), .B(n15376), .Z(n15375) );
  IV U18258 ( .A(n15373), .Z(n15376) );
  XOR U18259 ( .A(n15377), .B(n15378), .Z(n15373) );
  ANDN U18260 ( .B(n15379), .A(n15380), .Z(n15377) );
  XNOR U18261 ( .A(b[1215]), .B(n15378), .Z(n15379) );
  XNOR U18262 ( .A(b[1215]), .B(n15380), .Z(c[1215]) );
  XNOR U18263 ( .A(a[1215]), .B(n15381), .Z(n15380) );
  IV U18264 ( .A(n15378), .Z(n15381) );
  XOR U18265 ( .A(n15382), .B(n15383), .Z(n15378) );
  ANDN U18266 ( .B(n15384), .A(n15385), .Z(n15382) );
  XNOR U18267 ( .A(b[1214]), .B(n15383), .Z(n15384) );
  XNOR U18268 ( .A(b[1214]), .B(n15385), .Z(c[1214]) );
  XNOR U18269 ( .A(a[1214]), .B(n15386), .Z(n15385) );
  IV U18270 ( .A(n15383), .Z(n15386) );
  XOR U18271 ( .A(n15387), .B(n15388), .Z(n15383) );
  ANDN U18272 ( .B(n15389), .A(n15390), .Z(n15387) );
  XNOR U18273 ( .A(b[1213]), .B(n15388), .Z(n15389) );
  XNOR U18274 ( .A(b[1213]), .B(n15390), .Z(c[1213]) );
  XNOR U18275 ( .A(a[1213]), .B(n15391), .Z(n15390) );
  IV U18276 ( .A(n15388), .Z(n15391) );
  XOR U18277 ( .A(n15392), .B(n15393), .Z(n15388) );
  ANDN U18278 ( .B(n15394), .A(n15395), .Z(n15392) );
  XNOR U18279 ( .A(b[1212]), .B(n15393), .Z(n15394) );
  XNOR U18280 ( .A(b[1212]), .B(n15395), .Z(c[1212]) );
  XNOR U18281 ( .A(a[1212]), .B(n15396), .Z(n15395) );
  IV U18282 ( .A(n15393), .Z(n15396) );
  XOR U18283 ( .A(n15397), .B(n15398), .Z(n15393) );
  ANDN U18284 ( .B(n15399), .A(n15400), .Z(n15397) );
  XNOR U18285 ( .A(b[1211]), .B(n15398), .Z(n15399) );
  XNOR U18286 ( .A(b[1211]), .B(n15400), .Z(c[1211]) );
  XNOR U18287 ( .A(a[1211]), .B(n15401), .Z(n15400) );
  IV U18288 ( .A(n15398), .Z(n15401) );
  XOR U18289 ( .A(n15402), .B(n15403), .Z(n15398) );
  ANDN U18290 ( .B(n15404), .A(n15405), .Z(n15402) );
  XNOR U18291 ( .A(b[1210]), .B(n15403), .Z(n15404) );
  XNOR U18292 ( .A(b[1210]), .B(n15405), .Z(c[1210]) );
  XNOR U18293 ( .A(a[1210]), .B(n15406), .Z(n15405) );
  IV U18294 ( .A(n15403), .Z(n15406) );
  XOR U18295 ( .A(n15407), .B(n15408), .Z(n15403) );
  ANDN U18296 ( .B(n15409), .A(n15410), .Z(n15407) );
  XNOR U18297 ( .A(b[1209]), .B(n15408), .Z(n15409) );
  XNOR U18298 ( .A(b[120]), .B(n15411), .Z(c[120]) );
  XNOR U18299 ( .A(b[1209]), .B(n15410), .Z(c[1209]) );
  XNOR U18300 ( .A(a[1209]), .B(n15412), .Z(n15410) );
  IV U18301 ( .A(n15408), .Z(n15412) );
  XOR U18302 ( .A(n15413), .B(n15414), .Z(n15408) );
  ANDN U18303 ( .B(n15415), .A(n15416), .Z(n15413) );
  XNOR U18304 ( .A(b[1208]), .B(n15414), .Z(n15415) );
  XNOR U18305 ( .A(b[1208]), .B(n15416), .Z(c[1208]) );
  XNOR U18306 ( .A(a[1208]), .B(n15417), .Z(n15416) );
  IV U18307 ( .A(n15414), .Z(n15417) );
  XOR U18308 ( .A(n15418), .B(n15419), .Z(n15414) );
  ANDN U18309 ( .B(n15420), .A(n15421), .Z(n15418) );
  XNOR U18310 ( .A(b[1207]), .B(n15419), .Z(n15420) );
  XNOR U18311 ( .A(b[1207]), .B(n15421), .Z(c[1207]) );
  XNOR U18312 ( .A(a[1207]), .B(n15422), .Z(n15421) );
  IV U18313 ( .A(n15419), .Z(n15422) );
  XOR U18314 ( .A(n15423), .B(n15424), .Z(n15419) );
  ANDN U18315 ( .B(n15425), .A(n15426), .Z(n15423) );
  XNOR U18316 ( .A(b[1206]), .B(n15424), .Z(n15425) );
  XNOR U18317 ( .A(b[1206]), .B(n15426), .Z(c[1206]) );
  XNOR U18318 ( .A(a[1206]), .B(n15427), .Z(n15426) );
  IV U18319 ( .A(n15424), .Z(n15427) );
  XOR U18320 ( .A(n15428), .B(n15429), .Z(n15424) );
  ANDN U18321 ( .B(n15430), .A(n15431), .Z(n15428) );
  XNOR U18322 ( .A(b[1205]), .B(n15429), .Z(n15430) );
  XNOR U18323 ( .A(b[1205]), .B(n15431), .Z(c[1205]) );
  XNOR U18324 ( .A(a[1205]), .B(n15432), .Z(n15431) );
  IV U18325 ( .A(n15429), .Z(n15432) );
  XOR U18326 ( .A(n15433), .B(n15434), .Z(n15429) );
  ANDN U18327 ( .B(n15435), .A(n15436), .Z(n15433) );
  XNOR U18328 ( .A(b[1204]), .B(n15434), .Z(n15435) );
  XNOR U18329 ( .A(b[1204]), .B(n15436), .Z(c[1204]) );
  XNOR U18330 ( .A(a[1204]), .B(n15437), .Z(n15436) );
  IV U18331 ( .A(n15434), .Z(n15437) );
  XOR U18332 ( .A(n15438), .B(n15439), .Z(n15434) );
  ANDN U18333 ( .B(n15440), .A(n15441), .Z(n15438) );
  XNOR U18334 ( .A(b[1203]), .B(n15439), .Z(n15440) );
  XNOR U18335 ( .A(b[1203]), .B(n15441), .Z(c[1203]) );
  XNOR U18336 ( .A(a[1203]), .B(n15442), .Z(n15441) );
  IV U18337 ( .A(n15439), .Z(n15442) );
  XOR U18338 ( .A(n15443), .B(n15444), .Z(n15439) );
  ANDN U18339 ( .B(n15445), .A(n15446), .Z(n15443) );
  XNOR U18340 ( .A(b[1202]), .B(n15444), .Z(n15445) );
  XNOR U18341 ( .A(b[1202]), .B(n15446), .Z(c[1202]) );
  XNOR U18342 ( .A(a[1202]), .B(n15447), .Z(n15446) );
  IV U18343 ( .A(n15444), .Z(n15447) );
  XOR U18344 ( .A(n15448), .B(n15449), .Z(n15444) );
  ANDN U18345 ( .B(n15450), .A(n15451), .Z(n15448) );
  XNOR U18346 ( .A(b[1201]), .B(n15449), .Z(n15450) );
  XNOR U18347 ( .A(b[1201]), .B(n15451), .Z(c[1201]) );
  XNOR U18348 ( .A(a[1201]), .B(n15452), .Z(n15451) );
  IV U18349 ( .A(n15449), .Z(n15452) );
  XOR U18350 ( .A(n15453), .B(n15454), .Z(n15449) );
  ANDN U18351 ( .B(n15455), .A(n15456), .Z(n15453) );
  XNOR U18352 ( .A(b[1200]), .B(n15454), .Z(n15455) );
  XNOR U18353 ( .A(b[1200]), .B(n15456), .Z(c[1200]) );
  XNOR U18354 ( .A(a[1200]), .B(n15457), .Z(n15456) );
  IV U18355 ( .A(n15454), .Z(n15457) );
  XOR U18356 ( .A(n15458), .B(n15459), .Z(n15454) );
  ANDN U18357 ( .B(n15460), .A(n15461), .Z(n15458) );
  XNOR U18358 ( .A(b[1199]), .B(n15459), .Z(n15460) );
  XNOR U18359 ( .A(b[11]), .B(n15462), .Z(c[11]) );
  XNOR U18360 ( .A(b[119]), .B(n15463), .Z(c[119]) );
  XNOR U18361 ( .A(b[1199]), .B(n15461), .Z(c[1199]) );
  XNOR U18362 ( .A(a[1199]), .B(n15464), .Z(n15461) );
  IV U18363 ( .A(n15459), .Z(n15464) );
  XOR U18364 ( .A(n15465), .B(n15466), .Z(n15459) );
  ANDN U18365 ( .B(n15467), .A(n15468), .Z(n15465) );
  XNOR U18366 ( .A(b[1198]), .B(n15466), .Z(n15467) );
  XNOR U18367 ( .A(b[1198]), .B(n15468), .Z(c[1198]) );
  XNOR U18368 ( .A(a[1198]), .B(n15469), .Z(n15468) );
  IV U18369 ( .A(n15466), .Z(n15469) );
  XOR U18370 ( .A(n15470), .B(n15471), .Z(n15466) );
  ANDN U18371 ( .B(n15472), .A(n15473), .Z(n15470) );
  XNOR U18372 ( .A(b[1197]), .B(n15471), .Z(n15472) );
  XNOR U18373 ( .A(b[1197]), .B(n15473), .Z(c[1197]) );
  XNOR U18374 ( .A(a[1197]), .B(n15474), .Z(n15473) );
  IV U18375 ( .A(n15471), .Z(n15474) );
  XOR U18376 ( .A(n15475), .B(n15476), .Z(n15471) );
  ANDN U18377 ( .B(n15477), .A(n15478), .Z(n15475) );
  XNOR U18378 ( .A(b[1196]), .B(n15476), .Z(n15477) );
  XNOR U18379 ( .A(b[1196]), .B(n15478), .Z(c[1196]) );
  XNOR U18380 ( .A(a[1196]), .B(n15479), .Z(n15478) );
  IV U18381 ( .A(n15476), .Z(n15479) );
  XOR U18382 ( .A(n15480), .B(n15481), .Z(n15476) );
  ANDN U18383 ( .B(n15482), .A(n15483), .Z(n15480) );
  XNOR U18384 ( .A(b[1195]), .B(n15481), .Z(n15482) );
  XNOR U18385 ( .A(b[1195]), .B(n15483), .Z(c[1195]) );
  XNOR U18386 ( .A(a[1195]), .B(n15484), .Z(n15483) );
  IV U18387 ( .A(n15481), .Z(n15484) );
  XOR U18388 ( .A(n15485), .B(n15486), .Z(n15481) );
  ANDN U18389 ( .B(n15487), .A(n15488), .Z(n15485) );
  XNOR U18390 ( .A(b[1194]), .B(n15486), .Z(n15487) );
  XNOR U18391 ( .A(b[1194]), .B(n15488), .Z(c[1194]) );
  XNOR U18392 ( .A(a[1194]), .B(n15489), .Z(n15488) );
  IV U18393 ( .A(n15486), .Z(n15489) );
  XOR U18394 ( .A(n15490), .B(n15491), .Z(n15486) );
  ANDN U18395 ( .B(n15492), .A(n15493), .Z(n15490) );
  XNOR U18396 ( .A(b[1193]), .B(n15491), .Z(n15492) );
  XNOR U18397 ( .A(b[1193]), .B(n15493), .Z(c[1193]) );
  XNOR U18398 ( .A(a[1193]), .B(n15494), .Z(n15493) );
  IV U18399 ( .A(n15491), .Z(n15494) );
  XOR U18400 ( .A(n15495), .B(n15496), .Z(n15491) );
  ANDN U18401 ( .B(n15497), .A(n15498), .Z(n15495) );
  XNOR U18402 ( .A(b[1192]), .B(n15496), .Z(n15497) );
  XNOR U18403 ( .A(b[1192]), .B(n15498), .Z(c[1192]) );
  XNOR U18404 ( .A(a[1192]), .B(n15499), .Z(n15498) );
  IV U18405 ( .A(n15496), .Z(n15499) );
  XOR U18406 ( .A(n15500), .B(n15501), .Z(n15496) );
  ANDN U18407 ( .B(n15502), .A(n15503), .Z(n15500) );
  XNOR U18408 ( .A(b[1191]), .B(n15501), .Z(n15502) );
  XNOR U18409 ( .A(b[1191]), .B(n15503), .Z(c[1191]) );
  XNOR U18410 ( .A(a[1191]), .B(n15504), .Z(n15503) );
  IV U18411 ( .A(n15501), .Z(n15504) );
  XOR U18412 ( .A(n15505), .B(n15506), .Z(n15501) );
  ANDN U18413 ( .B(n15507), .A(n15508), .Z(n15505) );
  XNOR U18414 ( .A(b[1190]), .B(n15506), .Z(n15507) );
  XNOR U18415 ( .A(b[1190]), .B(n15508), .Z(c[1190]) );
  XNOR U18416 ( .A(a[1190]), .B(n15509), .Z(n15508) );
  IV U18417 ( .A(n15506), .Z(n15509) );
  XOR U18418 ( .A(n15510), .B(n15511), .Z(n15506) );
  ANDN U18419 ( .B(n15512), .A(n15513), .Z(n15510) );
  XNOR U18420 ( .A(b[1189]), .B(n15511), .Z(n15512) );
  XNOR U18421 ( .A(b[118]), .B(n15514), .Z(c[118]) );
  XNOR U18422 ( .A(b[1189]), .B(n15513), .Z(c[1189]) );
  XNOR U18423 ( .A(a[1189]), .B(n15515), .Z(n15513) );
  IV U18424 ( .A(n15511), .Z(n15515) );
  XOR U18425 ( .A(n15516), .B(n15517), .Z(n15511) );
  ANDN U18426 ( .B(n15518), .A(n15519), .Z(n15516) );
  XNOR U18427 ( .A(b[1188]), .B(n15517), .Z(n15518) );
  XNOR U18428 ( .A(b[1188]), .B(n15519), .Z(c[1188]) );
  XNOR U18429 ( .A(a[1188]), .B(n15520), .Z(n15519) );
  IV U18430 ( .A(n15517), .Z(n15520) );
  XOR U18431 ( .A(n15521), .B(n15522), .Z(n15517) );
  ANDN U18432 ( .B(n15523), .A(n15524), .Z(n15521) );
  XNOR U18433 ( .A(b[1187]), .B(n15522), .Z(n15523) );
  XNOR U18434 ( .A(b[1187]), .B(n15524), .Z(c[1187]) );
  XNOR U18435 ( .A(a[1187]), .B(n15525), .Z(n15524) );
  IV U18436 ( .A(n15522), .Z(n15525) );
  XOR U18437 ( .A(n15526), .B(n15527), .Z(n15522) );
  ANDN U18438 ( .B(n15528), .A(n15529), .Z(n15526) );
  XNOR U18439 ( .A(b[1186]), .B(n15527), .Z(n15528) );
  XNOR U18440 ( .A(b[1186]), .B(n15529), .Z(c[1186]) );
  XNOR U18441 ( .A(a[1186]), .B(n15530), .Z(n15529) );
  IV U18442 ( .A(n15527), .Z(n15530) );
  XOR U18443 ( .A(n15531), .B(n15532), .Z(n15527) );
  ANDN U18444 ( .B(n15533), .A(n15534), .Z(n15531) );
  XNOR U18445 ( .A(b[1185]), .B(n15532), .Z(n15533) );
  XNOR U18446 ( .A(b[1185]), .B(n15534), .Z(c[1185]) );
  XNOR U18447 ( .A(a[1185]), .B(n15535), .Z(n15534) );
  IV U18448 ( .A(n15532), .Z(n15535) );
  XOR U18449 ( .A(n15536), .B(n15537), .Z(n15532) );
  ANDN U18450 ( .B(n15538), .A(n15539), .Z(n15536) );
  XNOR U18451 ( .A(b[1184]), .B(n15537), .Z(n15538) );
  XNOR U18452 ( .A(b[1184]), .B(n15539), .Z(c[1184]) );
  XNOR U18453 ( .A(a[1184]), .B(n15540), .Z(n15539) );
  IV U18454 ( .A(n15537), .Z(n15540) );
  XOR U18455 ( .A(n15541), .B(n15542), .Z(n15537) );
  ANDN U18456 ( .B(n15543), .A(n15544), .Z(n15541) );
  XNOR U18457 ( .A(b[1183]), .B(n15542), .Z(n15543) );
  XNOR U18458 ( .A(b[1183]), .B(n15544), .Z(c[1183]) );
  XNOR U18459 ( .A(a[1183]), .B(n15545), .Z(n15544) );
  IV U18460 ( .A(n15542), .Z(n15545) );
  XOR U18461 ( .A(n15546), .B(n15547), .Z(n15542) );
  ANDN U18462 ( .B(n15548), .A(n15549), .Z(n15546) );
  XNOR U18463 ( .A(b[1182]), .B(n15547), .Z(n15548) );
  XNOR U18464 ( .A(b[1182]), .B(n15549), .Z(c[1182]) );
  XNOR U18465 ( .A(a[1182]), .B(n15550), .Z(n15549) );
  IV U18466 ( .A(n15547), .Z(n15550) );
  XOR U18467 ( .A(n15551), .B(n15552), .Z(n15547) );
  ANDN U18468 ( .B(n15553), .A(n15554), .Z(n15551) );
  XNOR U18469 ( .A(b[1181]), .B(n15552), .Z(n15553) );
  XNOR U18470 ( .A(b[1181]), .B(n15554), .Z(c[1181]) );
  XNOR U18471 ( .A(a[1181]), .B(n15555), .Z(n15554) );
  IV U18472 ( .A(n15552), .Z(n15555) );
  XOR U18473 ( .A(n15556), .B(n15557), .Z(n15552) );
  ANDN U18474 ( .B(n15558), .A(n15559), .Z(n15556) );
  XNOR U18475 ( .A(b[1180]), .B(n15557), .Z(n15558) );
  XNOR U18476 ( .A(b[1180]), .B(n15559), .Z(c[1180]) );
  XNOR U18477 ( .A(a[1180]), .B(n15560), .Z(n15559) );
  IV U18478 ( .A(n15557), .Z(n15560) );
  XOR U18479 ( .A(n15561), .B(n15562), .Z(n15557) );
  ANDN U18480 ( .B(n15563), .A(n15564), .Z(n15561) );
  XNOR U18481 ( .A(b[1179]), .B(n15562), .Z(n15563) );
  XNOR U18482 ( .A(b[117]), .B(n15565), .Z(c[117]) );
  XNOR U18483 ( .A(b[1179]), .B(n15564), .Z(c[1179]) );
  XNOR U18484 ( .A(a[1179]), .B(n15566), .Z(n15564) );
  IV U18485 ( .A(n15562), .Z(n15566) );
  XOR U18486 ( .A(n15567), .B(n15568), .Z(n15562) );
  ANDN U18487 ( .B(n15569), .A(n15570), .Z(n15567) );
  XNOR U18488 ( .A(b[1178]), .B(n15568), .Z(n15569) );
  XNOR U18489 ( .A(b[1178]), .B(n15570), .Z(c[1178]) );
  XNOR U18490 ( .A(a[1178]), .B(n15571), .Z(n15570) );
  IV U18491 ( .A(n15568), .Z(n15571) );
  XOR U18492 ( .A(n15572), .B(n15573), .Z(n15568) );
  ANDN U18493 ( .B(n15574), .A(n15575), .Z(n15572) );
  XNOR U18494 ( .A(b[1177]), .B(n15573), .Z(n15574) );
  XNOR U18495 ( .A(b[1177]), .B(n15575), .Z(c[1177]) );
  XNOR U18496 ( .A(a[1177]), .B(n15576), .Z(n15575) );
  IV U18497 ( .A(n15573), .Z(n15576) );
  XOR U18498 ( .A(n15577), .B(n15578), .Z(n15573) );
  ANDN U18499 ( .B(n15579), .A(n15580), .Z(n15577) );
  XNOR U18500 ( .A(b[1176]), .B(n15578), .Z(n15579) );
  XNOR U18501 ( .A(b[1176]), .B(n15580), .Z(c[1176]) );
  XNOR U18502 ( .A(a[1176]), .B(n15581), .Z(n15580) );
  IV U18503 ( .A(n15578), .Z(n15581) );
  XOR U18504 ( .A(n15582), .B(n15583), .Z(n15578) );
  ANDN U18505 ( .B(n15584), .A(n15585), .Z(n15582) );
  XNOR U18506 ( .A(b[1175]), .B(n15583), .Z(n15584) );
  XNOR U18507 ( .A(b[1175]), .B(n15585), .Z(c[1175]) );
  XNOR U18508 ( .A(a[1175]), .B(n15586), .Z(n15585) );
  IV U18509 ( .A(n15583), .Z(n15586) );
  XOR U18510 ( .A(n15587), .B(n15588), .Z(n15583) );
  ANDN U18511 ( .B(n15589), .A(n15590), .Z(n15587) );
  XNOR U18512 ( .A(b[1174]), .B(n15588), .Z(n15589) );
  XNOR U18513 ( .A(b[1174]), .B(n15590), .Z(c[1174]) );
  XNOR U18514 ( .A(a[1174]), .B(n15591), .Z(n15590) );
  IV U18515 ( .A(n15588), .Z(n15591) );
  XOR U18516 ( .A(n15592), .B(n15593), .Z(n15588) );
  ANDN U18517 ( .B(n15594), .A(n15595), .Z(n15592) );
  XNOR U18518 ( .A(b[1173]), .B(n15593), .Z(n15594) );
  XNOR U18519 ( .A(b[1173]), .B(n15595), .Z(c[1173]) );
  XNOR U18520 ( .A(a[1173]), .B(n15596), .Z(n15595) );
  IV U18521 ( .A(n15593), .Z(n15596) );
  XOR U18522 ( .A(n15597), .B(n15598), .Z(n15593) );
  ANDN U18523 ( .B(n15599), .A(n15600), .Z(n15597) );
  XNOR U18524 ( .A(b[1172]), .B(n15598), .Z(n15599) );
  XNOR U18525 ( .A(b[1172]), .B(n15600), .Z(c[1172]) );
  XNOR U18526 ( .A(a[1172]), .B(n15601), .Z(n15600) );
  IV U18527 ( .A(n15598), .Z(n15601) );
  XOR U18528 ( .A(n15602), .B(n15603), .Z(n15598) );
  ANDN U18529 ( .B(n15604), .A(n15605), .Z(n15602) );
  XNOR U18530 ( .A(b[1171]), .B(n15603), .Z(n15604) );
  XNOR U18531 ( .A(b[1171]), .B(n15605), .Z(c[1171]) );
  XNOR U18532 ( .A(a[1171]), .B(n15606), .Z(n15605) );
  IV U18533 ( .A(n15603), .Z(n15606) );
  XOR U18534 ( .A(n15607), .B(n15608), .Z(n15603) );
  ANDN U18535 ( .B(n15609), .A(n15610), .Z(n15607) );
  XNOR U18536 ( .A(b[1170]), .B(n15608), .Z(n15609) );
  XNOR U18537 ( .A(b[1170]), .B(n15610), .Z(c[1170]) );
  XNOR U18538 ( .A(a[1170]), .B(n15611), .Z(n15610) );
  IV U18539 ( .A(n15608), .Z(n15611) );
  XOR U18540 ( .A(n15612), .B(n15613), .Z(n15608) );
  ANDN U18541 ( .B(n15614), .A(n15615), .Z(n15612) );
  XNOR U18542 ( .A(b[1169]), .B(n15613), .Z(n15614) );
  XNOR U18543 ( .A(b[116]), .B(n15616), .Z(c[116]) );
  XNOR U18544 ( .A(b[1169]), .B(n15615), .Z(c[1169]) );
  XNOR U18545 ( .A(a[1169]), .B(n15617), .Z(n15615) );
  IV U18546 ( .A(n15613), .Z(n15617) );
  XOR U18547 ( .A(n15618), .B(n15619), .Z(n15613) );
  ANDN U18548 ( .B(n15620), .A(n15621), .Z(n15618) );
  XNOR U18549 ( .A(b[1168]), .B(n15619), .Z(n15620) );
  XNOR U18550 ( .A(b[1168]), .B(n15621), .Z(c[1168]) );
  XNOR U18551 ( .A(a[1168]), .B(n15622), .Z(n15621) );
  IV U18552 ( .A(n15619), .Z(n15622) );
  XOR U18553 ( .A(n15623), .B(n15624), .Z(n15619) );
  ANDN U18554 ( .B(n15625), .A(n15626), .Z(n15623) );
  XNOR U18555 ( .A(b[1167]), .B(n15624), .Z(n15625) );
  XNOR U18556 ( .A(b[1167]), .B(n15626), .Z(c[1167]) );
  XNOR U18557 ( .A(a[1167]), .B(n15627), .Z(n15626) );
  IV U18558 ( .A(n15624), .Z(n15627) );
  XOR U18559 ( .A(n15628), .B(n15629), .Z(n15624) );
  ANDN U18560 ( .B(n15630), .A(n15631), .Z(n15628) );
  XNOR U18561 ( .A(b[1166]), .B(n15629), .Z(n15630) );
  XNOR U18562 ( .A(b[1166]), .B(n15631), .Z(c[1166]) );
  XNOR U18563 ( .A(a[1166]), .B(n15632), .Z(n15631) );
  IV U18564 ( .A(n15629), .Z(n15632) );
  XOR U18565 ( .A(n15633), .B(n15634), .Z(n15629) );
  ANDN U18566 ( .B(n15635), .A(n15636), .Z(n15633) );
  XNOR U18567 ( .A(b[1165]), .B(n15634), .Z(n15635) );
  XNOR U18568 ( .A(b[1165]), .B(n15636), .Z(c[1165]) );
  XNOR U18569 ( .A(a[1165]), .B(n15637), .Z(n15636) );
  IV U18570 ( .A(n15634), .Z(n15637) );
  XOR U18571 ( .A(n15638), .B(n15639), .Z(n15634) );
  ANDN U18572 ( .B(n15640), .A(n15641), .Z(n15638) );
  XNOR U18573 ( .A(b[1164]), .B(n15639), .Z(n15640) );
  XNOR U18574 ( .A(b[1164]), .B(n15641), .Z(c[1164]) );
  XNOR U18575 ( .A(a[1164]), .B(n15642), .Z(n15641) );
  IV U18576 ( .A(n15639), .Z(n15642) );
  XOR U18577 ( .A(n15643), .B(n15644), .Z(n15639) );
  ANDN U18578 ( .B(n15645), .A(n15646), .Z(n15643) );
  XNOR U18579 ( .A(b[1163]), .B(n15644), .Z(n15645) );
  XNOR U18580 ( .A(b[1163]), .B(n15646), .Z(c[1163]) );
  XNOR U18581 ( .A(a[1163]), .B(n15647), .Z(n15646) );
  IV U18582 ( .A(n15644), .Z(n15647) );
  XOR U18583 ( .A(n15648), .B(n15649), .Z(n15644) );
  ANDN U18584 ( .B(n15650), .A(n15651), .Z(n15648) );
  XNOR U18585 ( .A(b[1162]), .B(n15649), .Z(n15650) );
  XNOR U18586 ( .A(b[1162]), .B(n15651), .Z(c[1162]) );
  XNOR U18587 ( .A(a[1162]), .B(n15652), .Z(n15651) );
  IV U18588 ( .A(n15649), .Z(n15652) );
  XOR U18589 ( .A(n15653), .B(n15654), .Z(n15649) );
  ANDN U18590 ( .B(n15655), .A(n15656), .Z(n15653) );
  XNOR U18591 ( .A(b[1161]), .B(n15654), .Z(n15655) );
  XNOR U18592 ( .A(b[1161]), .B(n15656), .Z(c[1161]) );
  XNOR U18593 ( .A(a[1161]), .B(n15657), .Z(n15656) );
  IV U18594 ( .A(n15654), .Z(n15657) );
  XOR U18595 ( .A(n15658), .B(n15659), .Z(n15654) );
  ANDN U18596 ( .B(n15660), .A(n15661), .Z(n15658) );
  XNOR U18597 ( .A(b[1160]), .B(n15659), .Z(n15660) );
  XNOR U18598 ( .A(b[1160]), .B(n15661), .Z(c[1160]) );
  XNOR U18599 ( .A(a[1160]), .B(n15662), .Z(n15661) );
  IV U18600 ( .A(n15659), .Z(n15662) );
  XOR U18601 ( .A(n15663), .B(n15664), .Z(n15659) );
  ANDN U18602 ( .B(n15665), .A(n15666), .Z(n15663) );
  XNOR U18603 ( .A(b[1159]), .B(n15664), .Z(n15665) );
  XNOR U18604 ( .A(b[115]), .B(n15667), .Z(c[115]) );
  XNOR U18605 ( .A(b[1159]), .B(n15666), .Z(c[1159]) );
  XNOR U18606 ( .A(a[1159]), .B(n15668), .Z(n15666) );
  IV U18607 ( .A(n15664), .Z(n15668) );
  XOR U18608 ( .A(n15669), .B(n15670), .Z(n15664) );
  ANDN U18609 ( .B(n15671), .A(n15672), .Z(n15669) );
  XNOR U18610 ( .A(b[1158]), .B(n15670), .Z(n15671) );
  XNOR U18611 ( .A(b[1158]), .B(n15672), .Z(c[1158]) );
  XNOR U18612 ( .A(a[1158]), .B(n15673), .Z(n15672) );
  IV U18613 ( .A(n15670), .Z(n15673) );
  XOR U18614 ( .A(n15674), .B(n15675), .Z(n15670) );
  ANDN U18615 ( .B(n15676), .A(n15677), .Z(n15674) );
  XNOR U18616 ( .A(b[1157]), .B(n15675), .Z(n15676) );
  XNOR U18617 ( .A(b[1157]), .B(n15677), .Z(c[1157]) );
  XNOR U18618 ( .A(a[1157]), .B(n15678), .Z(n15677) );
  IV U18619 ( .A(n15675), .Z(n15678) );
  XOR U18620 ( .A(n15679), .B(n15680), .Z(n15675) );
  ANDN U18621 ( .B(n15681), .A(n15682), .Z(n15679) );
  XNOR U18622 ( .A(b[1156]), .B(n15680), .Z(n15681) );
  XNOR U18623 ( .A(b[1156]), .B(n15682), .Z(c[1156]) );
  XNOR U18624 ( .A(a[1156]), .B(n15683), .Z(n15682) );
  IV U18625 ( .A(n15680), .Z(n15683) );
  XOR U18626 ( .A(n15684), .B(n15685), .Z(n15680) );
  ANDN U18627 ( .B(n15686), .A(n15687), .Z(n15684) );
  XNOR U18628 ( .A(b[1155]), .B(n15685), .Z(n15686) );
  XNOR U18629 ( .A(b[1155]), .B(n15687), .Z(c[1155]) );
  XNOR U18630 ( .A(a[1155]), .B(n15688), .Z(n15687) );
  IV U18631 ( .A(n15685), .Z(n15688) );
  XOR U18632 ( .A(n15689), .B(n15690), .Z(n15685) );
  ANDN U18633 ( .B(n15691), .A(n15692), .Z(n15689) );
  XNOR U18634 ( .A(b[1154]), .B(n15690), .Z(n15691) );
  XNOR U18635 ( .A(b[1154]), .B(n15692), .Z(c[1154]) );
  XNOR U18636 ( .A(a[1154]), .B(n15693), .Z(n15692) );
  IV U18637 ( .A(n15690), .Z(n15693) );
  XOR U18638 ( .A(n15694), .B(n15695), .Z(n15690) );
  ANDN U18639 ( .B(n15696), .A(n15697), .Z(n15694) );
  XNOR U18640 ( .A(b[1153]), .B(n15695), .Z(n15696) );
  XNOR U18641 ( .A(b[1153]), .B(n15697), .Z(c[1153]) );
  XNOR U18642 ( .A(a[1153]), .B(n15698), .Z(n15697) );
  IV U18643 ( .A(n15695), .Z(n15698) );
  XOR U18644 ( .A(n15699), .B(n15700), .Z(n15695) );
  ANDN U18645 ( .B(n15701), .A(n15702), .Z(n15699) );
  XNOR U18646 ( .A(b[1152]), .B(n15700), .Z(n15701) );
  XNOR U18647 ( .A(b[1152]), .B(n15702), .Z(c[1152]) );
  XNOR U18648 ( .A(a[1152]), .B(n15703), .Z(n15702) );
  IV U18649 ( .A(n15700), .Z(n15703) );
  XOR U18650 ( .A(n15704), .B(n15705), .Z(n15700) );
  ANDN U18651 ( .B(n15706), .A(n15707), .Z(n15704) );
  XNOR U18652 ( .A(b[1151]), .B(n15705), .Z(n15706) );
  XNOR U18653 ( .A(b[1151]), .B(n15707), .Z(c[1151]) );
  XNOR U18654 ( .A(a[1151]), .B(n15708), .Z(n15707) );
  IV U18655 ( .A(n15705), .Z(n15708) );
  XOR U18656 ( .A(n15709), .B(n15710), .Z(n15705) );
  ANDN U18657 ( .B(n15711), .A(n15712), .Z(n15709) );
  XNOR U18658 ( .A(b[1150]), .B(n15710), .Z(n15711) );
  XNOR U18659 ( .A(b[1150]), .B(n15712), .Z(c[1150]) );
  XNOR U18660 ( .A(a[1150]), .B(n15713), .Z(n15712) );
  IV U18661 ( .A(n15710), .Z(n15713) );
  XOR U18662 ( .A(n15714), .B(n15715), .Z(n15710) );
  ANDN U18663 ( .B(n15716), .A(n15717), .Z(n15714) );
  XNOR U18664 ( .A(b[1149]), .B(n15715), .Z(n15716) );
  XNOR U18665 ( .A(b[114]), .B(n15718), .Z(c[114]) );
  XNOR U18666 ( .A(b[1149]), .B(n15717), .Z(c[1149]) );
  XNOR U18667 ( .A(a[1149]), .B(n15719), .Z(n15717) );
  IV U18668 ( .A(n15715), .Z(n15719) );
  XOR U18669 ( .A(n15720), .B(n15721), .Z(n15715) );
  ANDN U18670 ( .B(n15722), .A(n15723), .Z(n15720) );
  XNOR U18671 ( .A(b[1148]), .B(n15721), .Z(n15722) );
  XNOR U18672 ( .A(b[1148]), .B(n15723), .Z(c[1148]) );
  XNOR U18673 ( .A(a[1148]), .B(n15724), .Z(n15723) );
  IV U18674 ( .A(n15721), .Z(n15724) );
  XOR U18675 ( .A(n15725), .B(n15726), .Z(n15721) );
  ANDN U18676 ( .B(n15727), .A(n15728), .Z(n15725) );
  XNOR U18677 ( .A(b[1147]), .B(n15726), .Z(n15727) );
  XNOR U18678 ( .A(b[1147]), .B(n15728), .Z(c[1147]) );
  XNOR U18679 ( .A(a[1147]), .B(n15729), .Z(n15728) );
  IV U18680 ( .A(n15726), .Z(n15729) );
  XOR U18681 ( .A(n15730), .B(n15731), .Z(n15726) );
  ANDN U18682 ( .B(n15732), .A(n15733), .Z(n15730) );
  XNOR U18683 ( .A(b[1146]), .B(n15731), .Z(n15732) );
  XNOR U18684 ( .A(b[1146]), .B(n15733), .Z(c[1146]) );
  XNOR U18685 ( .A(a[1146]), .B(n15734), .Z(n15733) );
  IV U18686 ( .A(n15731), .Z(n15734) );
  XOR U18687 ( .A(n15735), .B(n15736), .Z(n15731) );
  ANDN U18688 ( .B(n15737), .A(n15738), .Z(n15735) );
  XNOR U18689 ( .A(b[1145]), .B(n15736), .Z(n15737) );
  XNOR U18690 ( .A(b[1145]), .B(n15738), .Z(c[1145]) );
  XNOR U18691 ( .A(a[1145]), .B(n15739), .Z(n15738) );
  IV U18692 ( .A(n15736), .Z(n15739) );
  XOR U18693 ( .A(n15740), .B(n15741), .Z(n15736) );
  ANDN U18694 ( .B(n15742), .A(n15743), .Z(n15740) );
  XNOR U18695 ( .A(b[1144]), .B(n15741), .Z(n15742) );
  XNOR U18696 ( .A(b[1144]), .B(n15743), .Z(c[1144]) );
  XNOR U18697 ( .A(a[1144]), .B(n15744), .Z(n15743) );
  IV U18698 ( .A(n15741), .Z(n15744) );
  XOR U18699 ( .A(n15745), .B(n15746), .Z(n15741) );
  ANDN U18700 ( .B(n15747), .A(n15748), .Z(n15745) );
  XNOR U18701 ( .A(b[1143]), .B(n15746), .Z(n15747) );
  XNOR U18702 ( .A(b[1143]), .B(n15748), .Z(c[1143]) );
  XNOR U18703 ( .A(a[1143]), .B(n15749), .Z(n15748) );
  IV U18704 ( .A(n15746), .Z(n15749) );
  XOR U18705 ( .A(n15750), .B(n15751), .Z(n15746) );
  ANDN U18706 ( .B(n15752), .A(n15753), .Z(n15750) );
  XNOR U18707 ( .A(b[1142]), .B(n15751), .Z(n15752) );
  XNOR U18708 ( .A(b[1142]), .B(n15753), .Z(c[1142]) );
  XNOR U18709 ( .A(a[1142]), .B(n15754), .Z(n15753) );
  IV U18710 ( .A(n15751), .Z(n15754) );
  XOR U18711 ( .A(n15755), .B(n15756), .Z(n15751) );
  ANDN U18712 ( .B(n15757), .A(n15758), .Z(n15755) );
  XNOR U18713 ( .A(b[1141]), .B(n15756), .Z(n15757) );
  XNOR U18714 ( .A(b[1141]), .B(n15758), .Z(c[1141]) );
  XNOR U18715 ( .A(a[1141]), .B(n15759), .Z(n15758) );
  IV U18716 ( .A(n15756), .Z(n15759) );
  XOR U18717 ( .A(n15760), .B(n15761), .Z(n15756) );
  ANDN U18718 ( .B(n15762), .A(n15763), .Z(n15760) );
  XNOR U18719 ( .A(b[1140]), .B(n15761), .Z(n15762) );
  XNOR U18720 ( .A(b[1140]), .B(n15763), .Z(c[1140]) );
  XNOR U18721 ( .A(a[1140]), .B(n15764), .Z(n15763) );
  IV U18722 ( .A(n15761), .Z(n15764) );
  XOR U18723 ( .A(n15765), .B(n15766), .Z(n15761) );
  ANDN U18724 ( .B(n15767), .A(n15768), .Z(n15765) );
  XNOR U18725 ( .A(b[1139]), .B(n15766), .Z(n15767) );
  XNOR U18726 ( .A(b[113]), .B(n15769), .Z(c[113]) );
  XNOR U18727 ( .A(b[1139]), .B(n15768), .Z(c[1139]) );
  XNOR U18728 ( .A(a[1139]), .B(n15770), .Z(n15768) );
  IV U18729 ( .A(n15766), .Z(n15770) );
  XOR U18730 ( .A(n15771), .B(n15772), .Z(n15766) );
  ANDN U18731 ( .B(n15773), .A(n15774), .Z(n15771) );
  XNOR U18732 ( .A(b[1138]), .B(n15772), .Z(n15773) );
  XNOR U18733 ( .A(b[1138]), .B(n15774), .Z(c[1138]) );
  XNOR U18734 ( .A(a[1138]), .B(n15775), .Z(n15774) );
  IV U18735 ( .A(n15772), .Z(n15775) );
  XOR U18736 ( .A(n15776), .B(n15777), .Z(n15772) );
  ANDN U18737 ( .B(n15778), .A(n15779), .Z(n15776) );
  XNOR U18738 ( .A(b[1137]), .B(n15777), .Z(n15778) );
  XNOR U18739 ( .A(b[1137]), .B(n15779), .Z(c[1137]) );
  XNOR U18740 ( .A(a[1137]), .B(n15780), .Z(n15779) );
  IV U18741 ( .A(n15777), .Z(n15780) );
  XOR U18742 ( .A(n15781), .B(n15782), .Z(n15777) );
  ANDN U18743 ( .B(n15783), .A(n15784), .Z(n15781) );
  XNOR U18744 ( .A(b[1136]), .B(n15782), .Z(n15783) );
  XNOR U18745 ( .A(b[1136]), .B(n15784), .Z(c[1136]) );
  XNOR U18746 ( .A(a[1136]), .B(n15785), .Z(n15784) );
  IV U18747 ( .A(n15782), .Z(n15785) );
  XOR U18748 ( .A(n15786), .B(n15787), .Z(n15782) );
  ANDN U18749 ( .B(n15788), .A(n15789), .Z(n15786) );
  XNOR U18750 ( .A(b[1135]), .B(n15787), .Z(n15788) );
  XNOR U18751 ( .A(b[1135]), .B(n15789), .Z(c[1135]) );
  XNOR U18752 ( .A(a[1135]), .B(n15790), .Z(n15789) );
  IV U18753 ( .A(n15787), .Z(n15790) );
  XOR U18754 ( .A(n15791), .B(n15792), .Z(n15787) );
  ANDN U18755 ( .B(n15793), .A(n15794), .Z(n15791) );
  XNOR U18756 ( .A(b[1134]), .B(n15792), .Z(n15793) );
  XNOR U18757 ( .A(b[1134]), .B(n15794), .Z(c[1134]) );
  XNOR U18758 ( .A(a[1134]), .B(n15795), .Z(n15794) );
  IV U18759 ( .A(n15792), .Z(n15795) );
  XOR U18760 ( .A(n15796), .B(n15797), .Z(n15792) );
  ANDN U18761 ( .B(n15798), .A(n15799), .Z(n15796) );
  XNOR U18762 ( .A(b[1133]), .B(n15797), .Z(n15798) );
  XNOR U18763 ( .A(b[1133]), .B(n15799), .Z(c[1133]) );
  XNOR U18764 ( .A(a[1133]), .B(n15800), .Z(n15799) );
  IV U18765 ( .A(n15797), .Z(n15800) );
  XOR U18766 ( .A(n15801), .B(n15802), .Z(n15797) );
  ANDN U18767 ( .B(n15803), .A(n15804), .Z(n15801) );
  XNOR U18768 ( .A(b[1132]), .B(n15802), .Z(n15803) );
  XNOR U18769 ( .A(b[1132]), .B(n15804), .Z(c[1132]) );
  XNOR U18770 ( .A(a[1132]), .B(n15805), .Z(n15804) );
  IV U18771 ( .A(n15802), .Z(n15805) );
  XOR U18772 ( .A(n15806), .B(n15807), .Z(n15802) );
  ANDN U18773 ( .B(n15808), .A(n15809), .Z(n15806) );
  XNOR U18774 ( .A(b[1131]), .B(n15807), .Z(n15808) );
  XNOR U18775 ( .A(b[1131]), .B(n15809), .Z(c[1131]) );
  XNOR U18776 ( .A(a[1131]), .B(n15810), .Z(n15809) );
  IV U18777 ( .A(n15807), .Z(n15810) );
  XOR U18778 ( .A(n15811), .B(n15812), .Z(n15807) );
  ANDN U18779 ( .B(n15813), .A(n15814), .Z(n15811) );
  XNOR U18780 ( .A(b[1130]), .B(n15812), .Z(n15813) );
  XNOR U18781 ( .A(b[1130]), .B(n15814), .Z(c[1130]) );
  XNOR U18782 ( .A(a[1130]), .B(n15815), .Z(n15814) );
  IV U18783 ( .A(n15812), .Z(n15815) );
  XOR U18784 ( .A(n15816), .B(n15817), .Z(n15812) );
  ANDN U18785 ( .B(n15818), .A(n15819), .Z(n15816) );
  XNOR U18786 ( .A(b[1129]), .B(n15817), .Z(n15818) );
  XNOR U18787 ( .A(b[112]), .B(n15820), .Z(c[112]) );
  XNOR U18788 ( .A(b[1129]), .B(n15819), .Z(c[1129]) );
  XNOR U18789 ( .A(a[1129]), .B(n15821), .Z(n15819) );
  IV U18790 ( .A(n15817), .Z(n15821) );
  XOR U18791 ( .A(n15822), .B(n15823), .Z(n15817) );
  ANDN U18792 ( .B(n15824), .A(n15825), .Z(n15822) );
  XNOR U18793 ( .A(b[1128]), .B(n15823), .Z(n15824) );
  XNOR U18794 ( .A(b[1128]), .B(n15825), .Z(c[1128]) );
  XNOR U18795 ( .A(a[1128]), .B(n15826), .Z(n15825) );
  IV U18796 ( .A(n15823), .Z(n15826) );
  XOR U18797 ( .A(n15827), .B(n15828), .Z(n15823) );
  ANDN U18798 ( .B(n15829), .A(n15830), .Z(n15827) );
  XNOR U18799 ( .A(b[1127]), .B(n15828), .Z(n15829) );
  XNOR U18800 ( .A(b[1127]), .B(n15830), .Z(c[1127]) );
  XNOR U18801 ( .A(a[1127]), .B(n15831), .Z(n15830) );
  IV U18802 ( .A(n15828), .Z(n15831) );
  XOR U18803 ( .A(n15832), .B(n15833), .Z(n15828) );
  ANDN U18804 ( .B(n15834), .A(n15835), .Z(n15832) );
  XNOR U18805 ( .A(b[1126]), .B(n15833), .Z(n15834) );
  XNOR U18806 ( .A(b[1126]), .B(n15835), .Z(c[1126]) );
  XNOR U18807 ( .A(a[1126]), .B(n15836), .Z(n15835) );
  IV U18808 ( .A(n15833), .Z(n15836) );
  XOR U18809 ( .A(n15837), .B(n15838), .Z(n15833) );
  ANDN U18810 ( .B(n15839), .A(n15840), .Z(n15837) );
  XNOR U18811 ( .A(b[1125]), .B(n15838), .Z(n15839) );
  XNOR U18812 ( .A(b[1125]), .B(n15840), .Z(c[1125]) );
  XNOR U18813 ( .A(a[1125]), .B(n15841), .Z(n15840) );
  IV U18814 ( .A(n15838), .Z(n15841) );
  XOR U18815 ( .A(n15842), .B(n15843), .Z(n15838) );
  ANDN U18816 ( .B(n15844), .A(n15845), .Z(n15842) );
  XNOR U18817 ( .A(b[1124]), .B(n15843), .Z(n15844) );
  XNOR U18818 ( .A(b[1124]), .B(n15845), .Z(c[1124]) );
  XNOR U18819 ( .A(a[1124]), .B(n15846), .Z(n15845) );
  IV U18820 ( .A(n15843), .Z(n15846) );
  XOR U18821 ( .A(n15847), .B(n15848), .Z(n15843) );
  ANDN U18822 ( .B(n15849), .A(n15850), .Z(n15847) );
  XNOR U18823 ( .A(b[1123]), .B(n15848), .Z(n15849) );
  XNOR U18824 ( .A(b[1123]), .B(n15850), .Z(c[1123]) );
  XNOR U18825 ( .A(a[1123]), .B(n15851), .Z(n15850) );
  IV U18826 ( .A(n15848), .Z(n15851) );
  XOR U18827 ( .A(n15852), .B(n15853), .Z(n15848) );
  ANDN U18828 ( .B(n15854), .A(n15855), .Z(n15852) );
  XNOR U18829 ( .A(b[1122]), .B(n15853), .Z(n15854) );
  XNOR U18830 ( .A(b[1122]), .B(n15855), .Z(c[1122]) );
  XNOR U18831 ( .A(a[1122]), .B(n15856), .Z(n15855) );
  IV U18832 ( .A(n15853), .Z(n15856) );
  XOR U18833 ( .A(n15857), .B(n15858), .Z(n15853) );
  ANDN U18834 ( .B(n15859), .A(n15860), .Z(n15857) );
  XNOR U18835 ( .A(b[1121]), .B(n15858), .Z(n15859) );
  XNOR U18836 ( .A(b[1121]), .B(n15860), .Z(c[1121]) );
  XNOR U18837 ( .A(a[1121]), .B(n15861), .Z(n15860) );
  IV U18838 ( .A(n15858), .Z(n15861) );
  XOR U18839 ( .A(n15862), .B(n15863), .Z(n15858) );
  ANDN U18840 ( .B(n15864), .A(n15865), .Z(n15862) );
  XNOR U18841 ( .A(b[1120]), .B(n15863), .Z(n15864) );
  XNOR U18842 ( .A(b[1120]), .B(n15865), .Z(c[1120]) );
  XNOR U18843 ( .A(a[1120]), .B(n15866), .Z(n15865) );
  IV U18844 ( .A(n15863), .Z(n15866) );
  XOR U18845 ( .A(n15867), .B(n15868), .Z(n15863) );
  ANDN U18846 ( .B(n15869), .A(n15870), .Z(n15867) );
  XNOR U18847 ( .A(b[1119]), .B(n15868), .Z(n15869) );
  XNOR U18848 ( .A(b[111]), .B(n15871), .Z(c[111]) );
  XNOR U18849 ( .A(b[1119]), .B(n15870), .Z(c[1119]) );
  XNOR U18850 ( .A(a[1119]), .B(n15872), .Z(n15870) );
  IV U18851 ( .A(n15868), .Z(n15872) );
  XOR U18852 ( .A(n15873), .B(n15874), .Z(n15868) );
  ANDN U18853 ( .B(n15875), .A(n15876), .Z(n15873) );
  XNOR U18854 ( .A(b[1118]), .B(n15874), .Z(n15875) );
  XNOR U18855 ( .A(b[1118]), .B(n15876), .Z(c[1118]) );
  XNOR U18856 ( .A(a[1118]), .B(n15877), .Z(n15876) );
  IV U18857 ( .A(n15874), .Z(n15877) );
  XOR U18858 ( .A(n15878), .B(n15879), .Z(n15874) );
  ANDN U18859 ( .B(n15880), .A(n15881), .Z(n15878) );
  XNOR U18860 ( .A(b[1117]), .B(n15879), .Z(n15880) );
  XNOR U18861 ( .A(b[1117]), .B(n15881), .Z(c[1117]) );
  XNOR U18862 ( .A(a[1117]), .B(n15882), .Z(n15881) );
  IV U18863 ( .A(n15879), .Z(n15882) );
  XOR U18864 ( .A(n15883), .B(n15884), .Z(n15879) );
  ANDN U18865 ( .B(n15885), .A(n15886), .Z(n15883) );
  XNOR U18866 ( .A(b[1116]), .B(n15884), .Z(n15885) );
  XNOR U18867 ( .A(b[1116]), .B(n15886), .Z(c[1116]) );
  XNOR U18868 ( .A(a[1116]), .B(n15887), .Z(n15886) );
  IV U18869 ( .A(n15884), .Z(n15887) );
  XOR U18870 ( .A(n15888), .B(n15889), .Z(n15884) );
  ANDN U18871 ( .B(n15890), .A(n15891), .Z(n15888) );
  XNOR U18872 ( .A(b[1115]), .B(n15889), .Z(n15890) );
  XNOR U18873 ( .A(b[1115]), .B(n15891), .Z(c[1115]) );
  XNOR U18874 ( .A(a[1115]), .B(n15892), .Z(n15891) );
  IV U18875 ( .A(n15889), .Z(n15892) );
  XOR U18876 ( .A(n15893), .B(n15894), .Z(n15889) );
  ANDN U18877 ( .B(n15895), .A(n15896), .Z(n15893) );
  XNOR U18878 ( .A(b[1114]), .B(n15894), .Z(n15895) );
  XNOR U18879 ( .A(b[1114]), .B(n15896), .Z(c[1114]) );
  XNOR U18880 ( .A(a[1114]), .B(n15897), .Z(n15896) );
  IV U18881 ( .A(n15894), .Z(n15897) );
  XOR U18882 ( .A(n15898), .B(n15899), .Z(n15894) );
  ANDN U18883 ( .B(n15900), .A(n15901), .Z(n15898) );
  XNOR U18884 ( .A(b[1113]), .B(n15899), .Z(n15900) );
  XNOR U18885 ( .A(b[1113]), .B(n15901), .Z(c[1113]) );
  XNOR U18886 ( .A(a[1113]), .B(n15902), .Z(n15901) );
  IV U18887 ( .A(n15899), .Z(n15902) );
  XOR U18888 ( .A(n15903), .B(n15904), .Z(n15899) );
  ANDN U18889 ( .B(n15905), .A(n15906), .Z(n15903) );
  XNOR U18890 ( .A(b[1112]), .B(n15904), .Z(n15905) );
  XNOR U18891 ( .A(b[1112]), .B(n15906), .Z(c[1112]) );
  XNOR U18892 ( .A(a[1112]), .B(n15907), .Z(n15906) );
  IV U18893 ( .A(n15904), .Z(n15907) );
  XOR U18894 ( .A(n15908), .B(n15909), .Z(n15904) );
  ANDN U18895 ( .B(n15910), .A(n15911), .Z(n15908) );
  XNOR U18896 ( .A(b[1111]), .B(n15909), .Z(n15910) );
  XNOR U18897 ( .A(b[1111]), .B(n15911), .Z(c[1111]) );
  XNOR U18898 ( .A(a[1111]), .B(n15912), .Z(n15911) );
  IV U18899 ( .A(n15909), .Z(n15912) );
  XOR U18900 ( .A(n15913), .B(n15914), .Z(n15909) );
  ANDN U18901 ( .B(n15915), .A(n15916), .Z(n15913) );
  XNOR U18902 ( .A(b[1110]), .B(n15914), .Z(n15915) );
  XNOR U18903 ( .A(b[1110]), .B(n15916), .Z(c[1110]) );
  XNOR U18904 ( .A(a[1110]), .B(n15917), .Z(n15916) );
  IV U18905 ( .A(n15914), .Z(n15917) );
  XOR U18906 ( .A(n15918), .B(n15919), .Z(n15914) );
  ANDN U18907 ( .B(n15920), .A(n15921), .Z(n15918) );
  XNOR U18908 ( .A(b[1109]), .B(n15919), .Z(n15920) );
  XNOR U18909 ( .A(b[110]), .B(n15922), .Z(c[110]) );
  XNOR U18910 ( .A(b[1109]), .B(n15921), .Z(c[1109]) );
  XNOR U18911 ( .A(a[1109]), .B(n15923), .Z(n15921) );
  IV U18912 ( .A(n15919), .Z(n15923) );
  XOR U18913 ( .A(n15924), .B(n15925), .Z(n15919) );
  ANDN U18914 ( .B(n15926), .A(n15927), .Z(n15924) );
  XNOR U18915 ( .A(b[1108]), .B(n15925), .Z(n15926) );
  XNOR U18916 ( .A(b[1108]), .B(n15927), .Z(c[1108]) );
  XNOR U18917 ( .A(a[1108]), .B(n15928), .Z(n15927) );
  IV U18918 ( .A(n15925), .Z(n15928) );
  XOR U18919 ( .A(n15929), .B(n15930), .Z(n15925) );
  ANDN U18920 ( .B(n15931), .A(n15932), .Z(n15929) );
  XNOR U18921 ( .A(b[1107]), .B(n15930), .Z(n15931) );
  XNOR U18922 ( .A(b[1107]), .B(n15932), .Z(c[1107]) );
  XNOR U18923 ( .A(a[1107]), .B(n15933), .Z(n15932) );
  IV U18924 ( .A(n15930), .Z(n15933) );
  XOR U18925 ( .A(n15934), .B(n15935), .Z(n15930) );
  ANDN U18926 ( .B(n15936), .A(n15937), .Z(n15934) );
  XNOR U18927 ( .A(b[1106]), .B(n15935), .Z(n15936) );
  XNOR U18928 ( .A(b[1106]), .B(n15937), .Z(c[1106]) );
  XNOR U18929 ( .A(a[1106]), .B(n15938), .Z(n15937) );
  IV U18930 ( .A(n15935), .Z(n15938) );
  XOR U18931 ( .A(n15939), .B(n15940), .Z(n15935) );
  ANDN U18932 ( .B(n15941), .A(n15942), .Z(n15939) );
  XNOR U18933 ( .A(b[1105]), .B(n15940), .Z(n15941) );
  XNOR U18934 ( .A(b[1105]), .B(n15942), .Z(c[1105]) );
  XNOR U18935 ( .A(a[1105]), .B(n15943), .Z(n15942) );
  IV U18936 ( .A(n15940), .Z(n15943) );
  XOR U18937 ( .A(n15944), .B(n15945), .Z(n15940) );
  ANDN U18938 ( .B(n15946), .A(n15947), .Z(n15944) );
  XNOR U18939 ( .A(b[1104]), .B(n15945), .Z(n15946) );
  XNOR U18940 ( .A(b[1104]), .B(n15947), .Z(c[1104]) );
  XNOR U18941 ( .A(a[1104]), .B(n15948), .Z(n15947) );
  IV U18942 ( .A(n15945), .Z(n15948) );
  XOR U18943 ( .A(n15949), .B(n15950), .Z(n15945) );
  ANDN U18944 ( .B(n15951), .A(n15952), .Z(n15949) );
  XNOR U18945 ( .A(b[1103]), .B(n15950), .Z(n15951) );
  XNOR U18946 ( .A(b[1103]), .B(n15952), .Z(c[1103]) );
  XNOR U18947 ( .A(a[1103]), .B(n15953), .Z(n15952) );
  IV U18948 ( .A(n15950), .Z(n15953) );
  XOR U18949 ( .A(n15954), .B(n15955), .Z(n15950) );
  ANDN U18950 ( .B(n15956), .A(n15957), .Z(n15954) );
  XNOR U18951 ( .A(b[1102]), .B(n15955), .Z(n15956) );
  XNOR U18952 ( .A(b[1102]), .B(n15957), .Z(c[1102]) );
  XNOR U18953 ( .A(a[1102]), .B(n15958), .Z(n15957) );
  IV U18954 ( .A(n15955), .Z(n15958) );
  XOR U18955 ( .A(n15959), .B(n15960), .Z(n15955) );
  ANDN U18956 ( .B(n15961), .A(n15962), .Z(n15959) );
  XNOR U18957 ( .A(b[1101]), .B(n15960), .Z(n15961) );
  XNOR U18958 ( .A(b[1101]), .B(n15962), .Z(c[1101]) );
  XNOR U18959 ( .A(a[1101]), .B(n15963), .Z(n15962) );
  IV U18960 ( .A(n15960), .Z(n15963) );
  XOR U18961 ( .A(n15964), .B(n15965), .Z(n15960) );
  ANDN U18962 ( .B(n15966), .A(n15967), .Z(n15964) );
  XNOR U18963 ( .A(b[1100]), .B(n15965), .Z(n15966) );
  XNOR U18964 ( .A(b[1100]), .B(n15967), .Z(c[1100]) );
  XNOR U18965 ( .A(a[1100]), .B(n15968), .Z(n15967) );
  IV U18966 ( .A(n15965), .Z(n15968) );
  XOR U18967 ( .A(n15969), .B(n15970), .Z(n15965) );
  ANDN U18968 ( .B(n15971), .A(n15972), .Z(n15969) );
  XNOR U18969 ( .A(b[1099]), .B(n15970), .Z(n15971) );
  XNOR U18970 ( .A(b[10]), .B(n15973), .Z(c[10]) );
  XNOR U18971 ( .A(b[109]), .B(n15974), .Z(c[109]) );
  XNOR U18972 ( .A(b[1099]), .B(n15972), .Z(c[1099]) );
  XNOR U18973 ( .A(a[1099]), .B(n15975), .Z(n15972) );
  IV U18974 ( .A(n15970), .Z(n15975) );
  XOR U18975 ( .A(n15976), .B(n15977), .Z(n15970) );
  ANDN U18976 ( .B(n15978), .A(n15979), .Z(n15976) );
  XNOR U18977 ( .A(b[1098]), .B(n15977), .Z(n15978) );
  XNOR U18978 ( .A(b[1098]), .B(n15979), .Z(c[1098]) );
  XNOR U18979 ( .A(a[1098]), .B(n15980), .Z(n15979) );
  IV U18980 ( .A(n15977), .Z(n15980) );
  XOR U18981 ( .A(n15981), .B(n15982), .Z(n15977) );
  ANDN U18982 ( .B(n15983), .A(n15984), .Z(n15981) );
  XNOR U18983 ( .A(b[1097]), .B(n15982), .Z(n15983) );
  XNOR U18984 ( .A(b[1097]), .B(n15984), .Z(c[1097]) );
  XNOR U18985 ( .A(a[1097]), .B(n15985), .Z(n15984) );
  IV U18986 ( .A(n15982), .Z(n15985) );
  XOR U18987 ( .A(n15986), .B(n15987), .Z(n15982) );
  ANDN U18988 ( .B(n15988), .A(n15989), .Z(n15986) );
  XNOR U18989 ( .A(b[1096]), .B(n15987), .Z(n15988) );
  XNOR U18990 ( .A(b[1096]), .B(n15989), .Z(c[1096]) );
  XNOR U18991 ( .A(a[1096]), .B(n15990), .Z(n15989) );
  IV U18992 ( .A(n15987), .Z(n15990) );
  XOR U18993 ( .A(n15991), .B(n15992), .Z(n15987) );
  ANDN U18994 ( .B(n15993), .A(n15994), .Z(n15991) );
  XNOR U18995 ( .A(b[1095]), .B(n15992), .Z(n15993) );
  XNOR U18996 ( .A(b[1095]), .B(n15994), .Z(c[1095]) );
  XNOR U18997 ( .A(a[1095]), .B(n15995), .Z(n15994) );
  IV U18998 ( .A(n15992), .Z(n15995) );
  XOR U18999 ( .A(n15996), .B(n15997), .Z(n15992) );
  ANDN U19000 ( .B(n15998), .A(n15999), .Z(n15996) );
  XNOR U19001 ( .A(b[1094]), .B(n15997), .Z(n15998) );
  XNOR U19002 ( .A(b[1094]), .B(n15999), .Z(c[1094]) );
  XNOR U19003 ( .A(a[1094]), .B(n16000), .Z(n15999) );
  IV U19004 ( .A(n15997), .Z(n16000) );
  XOR U19005 ( .A(n16001), .B(n16002), .Z(n15997) );
  ANDN U19006 ( .B(n16003), .A(n16004), .Z(n16001) );
  XNOR U19007 ( .A(b[1093]), .B(n16002), .Z(n16003) );
  XNOR U19008 ( .A(b[1093]), .B(n16004), .Z(c[1093]) );
  XNOR U19009 ( .A(a[1093]), .B(n16005), .Z(n16004) );
  IV U19010 ( .A(n16002), .Z(n16005) );
  XOR U19011 ( .A(n16006), .B(n16007), .Z(n16002) );
  ANDN U19012 ( .B(n16008), .A(n16009), .Z(n16006) );
  XNOR U19013 ( .A(b[1092]), .B(n16007), .Z(n16008) );
  XNOR U19014 ( .A(b[1092]), .B(n16009), .Z(c[1092]) );
  XNOR U19015 ( .A(a[1092]), .B(n16010), .Z(n16009) );
  IV U19016 ( .A(n16007), .Z(n16010) );
  XOR U19017 ( .A(n16011), .B(n16012), .Z(n16007) );
  ANDN U19018 ( .B(n16013), .A(n16014), .Z(n16011) );
  XNOR U19019 ( .A(b[1091]), .B(n16012), .Z(n16013) );
  XNOR U19020 ( .A(b[1091]), .B(n16014), .Z(c[1091]) );
  XNOR U19021 ( .A(a[1091]), .B(n16015), .Z(n16014) );
  IV U19022 ( .A(n16012), .Z(n16015) );
  XOR U19023 ( .A(n16016), .B(n16017), .Z(n16012) );
  ANDN U19024 ( .B(n16018), .A(n16019), .Z(n16016) );
  XNOR U19025 ( .A(b[1090]), .B(n16017), .Z(n16018) );
  XNOR U19026 ( .A(b[1090]), .B(n16019), .Z(c[1090]) );
  XNOR U19027 ( .A(a[1090]), .B(n16020), .Z(n16019) );
  IV U19028 ( .A(n16017), .Z(n16020) );
  XOR U19029 ( .A(n16021), .B(n16022), .Z(n16017) );
  ANDN U19030 ( .B(n16023), .A(n16024), .Z(n16021) );
  XNOR U19031 ( .A(b[1089]), .B(n16022), .Z(n16023) );
  XNOR U19032 ( .A(b[108]), .B(n16025), .Z(c[108]) );
  XNOR U19033 ( .A(b[1089]), .B(n16024), .Z(c[1089]) );
  XNOR U19034 ( .A(a[1089]), .B(n16026), .Z(n16024) );
  IV U19035 ( .A(n16022), .Z(n16026) );
  XOR U19036 ( .A(n16027), .B(n16028), .Z(n16022) );
  ANDN U19037 ( .B(n16029), .A(n16030), .Z(n16027) );
  XNOR U19038 ( .A(b[1088]), .B(n16028), .Z(n16029) );
  XNOR U19039 ( .A(b[1088]), .B(n16030), .Z(c[1088]) );
  XNOR U19040 ( .A(a[1088]), .B(n16031), .Z(n16030) );
  IV U19041 ( .A(n16028), .Z(n16031) );
  XOR U19042 ( .A(n16032), .B(n16033), .Z(n16028) );
  ANDN U19043 ( .B(n16034), .A(n16035), .Z(n16032) );
  XNOR U19044 ( .A(b[1087]), .B(n16033), .Z(n16034) );
  XNOR U19045 ( .A(b[1087]), .B(n16035), .Z(c[1087]) );
  XNOR U19046 ( .A(a[1087]), .B(n16036), .Z(n16035) );
  IV U19047 ( .A(n16033), .Z(n16036) );
  XOR U19048 ( .A(n16037), .B(n16038), .Z(n16033) );
  ANDN U19049 ( .B(n16039), .A(n16040), .Z(n16037) );
  XNOR U19050 ( .A(b[1086]), .B(n16038), .Z(n16039) );
  XNOR U19051 ( .A(b[1086]), .B(n16040), .Z(c[1086]) );
  XNOR U19052 ( .A(a[1086]), .B(n16041), .Z(n16040) );
  IV U19053 ( .A(n16038), .Z(n16041) );
  XOR U19054 ( .A(n16042), .B(n16043), .Z(n16038) );
  ANDN U19055 ( .B(n16044), .A(n16045), .Z(n16042) );
  XNOR U19056 ( .A(b[1085]), .B(n16043), .Z(n16044) );
  XNOR U19057 ( .A(b[1085]), .B(n16045), .Z(c[1085]) );
  XNOR U19058 ( .A(a[1085]), .B(n16046), .Z(n16045) );
  IV U19059 ( .A(n16043), .Z(n16046) );
  XOR U19060 ( .A(n16047), .B(n16048), .Z(n16043) );
  ANDN U19061 ( .B(n16049), .A(n16050), .Z(n16047) );
  XNOR U19062 ( .A(b[1084]), .B(n16048), .Z(n16049) );
  XNOR U19063 ( .A(b[1084]), .B(n16050), .Z(c[1084]) );
  XNOR U19064 ( .A(a[1084]), .B(n16051), .Z(n16050) );
  IV U19065 ( .A(n16048), .Z(n16051) );
  XOR U19066 ( .A(n16052), .B(n16053), .Z(n16048) );
  ANDN U19067 ( .B(n16054), .A(n16055), .Z(n16052) );
  XNOR U19068 ( .A(b[1083]), .B(n16053), .Z(n16054) );
  XNOR U19069 ( .A(b[1083]), .B(n16055), .Z(c[1083]) );
  XNOR U19070 ( .A(a[1083]), .B(n16056), .Z(n16055) );
  IV U19071 ( .A(n16053), .Z(n16056) );
  XOR U19072 ( .A(n16057), .B(n16058), .Z(n16053) );
  ANDN U19073 ( .B(n16059), .A(n16060), .Z(n16057) );
  XNOR U19074 ( .A(b[1082]), .B(n16058), .Z(n16059) );
  XNOR U19075 ( .A(b[1082]), .B(n16060), .Z(c[1082]) );
  XNOR U19076 ( .A(a[1082]), .B(n16061), .Z(n16060) );
  IV U19077 ( .A(n16058), .Z(n16061) );
  XOR U19078 ( .A(n16062), .B(n16063), .Z(n16058) );
  ANDN U19079 ( .B(n16064), .A(n16065), .Z(n16062) );
  XNOR U19080 ( .A(b[1081]), .B(n16063), .Z(n16064) );
  XNOR U19081 ( .A(b[1081]), .B(n16065), .Z(c[1081]) );
  XNOR U19082 ( .A(a[1081]), .B(n16066), .Z(n16065) );
  IV U19083 ( .A(n16063), .Z(n16066) );
  XOR U19084 ( .A(n16067), .B(n16068), .Z(n16063) );
  ANDN U19085 ( .B(n16069), .A(n16070), .Z(n16067) );
  XNOR U19086 ( .A(b[1080]), .B(n16068), .Z(n16069) );
  XNOR U19087 ( .A(b[1080]), .B(n16070), .Z(c[1080]) );
  XNOR U19088 ( .A(a[1080]), .B(n16071), .Z(n16070) );
  IV U19089 ( .A(n16068), .Z(n16071) );
  XOR U19090 ( .A(n16072), .B(n16073), .Z(n16068) );
  ANDN U19091 ( .B(n16074), .A(n16075), .Z(n16072) );
  XNOR U19092 ( .A(b[1079]), .B(n16073), .Z(n16074) );
  XNOR U19093 ( .A(b[107]), .B(n16076), .Z(c[107]) );
  XNOR U19094 ( .A(b[1079]), .B(n16075), .Z(c[1079]) );
  XNOR U19095 ( .A(a[1079]), .B(n16077), .Z(n16075) );
  IV U19096 ( .A(n16073), .Z(n16077) );
  XOR U19097 ( .A(n16078), .B(n16079), .Z(n16073) );
  ANDN U19098 ( .B(n16080), .A(n16081), .Z(n16078) );
  XNOR U19099 ( .A(b[1078]), .B(n16079), .Z(n16080) );
  XNOR U19100 ( .A(b[1078]), .B(n16081), .Z(c[1078]) );
  XNOR U19101 ( .A(a[1078]), .B(n16082), .Z(n16081) );
  IV U19102 ( .A(n16079), .Z(n16082) );
  XOR U19103 ( .A(n16083), .B(n16084), .Z(n16079) );
  ANDN U19104 ( .B(n16085), .A(n16086), .Z(n16083) );
  XNOR U19105 ( .A(b[1077]), .B(n16084), .Z(n16085) );
  XNOR U19106 ( .A(b[1077]), .B(n16086), .Z(c[1077]) );
  XNOR U19107 ( .A(a[1077]), .B(n16087), .Z(n16086) );
  IV U19108 ( .A(n16084), .Z(n16087) );
  XOR U19109 ( .A(n16088), .B(n16089), .Z(n16084) );
  ANDN U19110 ( .B(n16090), .A(n16091), .Z(n16088) );
  XNOR U19111 ( .A(b[1076]), .B(n16089), .Z(n16090) );
  XNOR U19112 ( .A(b[1076]), .B(n16091), .Z(c[1076]) );
  XNOR U19113 ( .A(a[1076]), .B(n16092), .Z(n16091) );
  IV U19114 ( .A(n16089), .Z(n16092) );
  XOR U19115 ( .A(n16093), .B(n16094), .Z(n16089) );
  ANDN U19116 ( .B(n16095), .A(n16096), .Z(n16093) );
  XNOR U19117 ( .A(b[1075]), .B(n16094), .Z(n16095) );
  XNOR U19118 ( .A(b[1075]), .B(n16096), .Z(c[1075]) );
  XNOR U19119 ( .A(a[1075]), .B(n16097), .Z(n16096) );
  IV U19120 ( .A(n16094), .Z(n16097) );
  XOR U19121 ( .A(n16098), .B(n16099), .Z(n16094) );
  ANDN U19122 ( .B(n16100), .A(n16101), .Z(n16098) );
  XNOR U19123 ( .A(b[1074]), .B(n16099), .Z(n16100) );
  XNOR U19124 ( .A(b[1074]), .B(n16101), .Z(c[1074]) );
  XNOR U19125 ( .A(a[1074]), .B(n16102), .Z(n16101) );
  IV U19126 ( .A(n16099), .Z(n16102) );
  XOR U19127 ( .A(n16103), .B(n16104), .Z(n16099) );
  ANDN U19128 ( .B(n16105), .A(n16106), .Z(n16103) );
  XNOR U19129 ( .A(b[1073]), .B(n16104), .Z(n16105) );
  XNOR U19130 ( .A(b[1073]), .B(n16106), .Z(c[1073]) );
  XNOR U19131 ( .A(a[1073]), .B(n16107), .Z(n16106) );
  IV U19132 ( .A(n16104), .Z(n16107) );
  XOR U19133 ( .A(n16108), .B(n16109), .Z(n16104) );
  ANDN U19134 ( .B(n16110), .A(n16111), .Z(n16108) );
  XNOR U19135 ( .A(b[1072]), .B(n16109), .Z(n16110) );
  XNOR U19136 ( .A(b[1072]), .B(n16111), .Z(c[1072]) );
  XNOR U19137 ( .A(a[1072]), .B(n16112), .Z(n16111) );
  IV U19138 ( .A(n16109), .Z(n16112) );
  XOR U19139 ( .A(n16113), .B(n16114), .Z(n16109) );
  ANDN U19140 ( .B(n16115), .A(n16116), .Z(n16113) );
  XNOR U19141 ( .A(b[1071]), .B(n16114), .Z(n16115) );
  XNOR U19142 ( .A(b[1071]), .B(n16116), .Z(c[1071]) );
  XNOR U19143 ( .A(a[1071]), .B(n16117), .Z(n16116) );
  IV U19144 ( .A(n16114), .Z(n16117) );
  XOR U19145 ( .A(n16118), .B(n16119), .Z(n16114) );
  ANDN U19146 ( .B(n16120), .A(n16121), .Z(n16118) );
  XNOR U19147 ( .A(b[1070]), .B(n16119), .Z(n16120) );
  XNOR U19148 ( .A(b[1070]), .B(n16121), .Z(c[1070]) );
  XNOR U19149 ( .A(a[1070]), .B(n16122), .Z(n16121) );
  IV U19150 ( .A(n16119), .Z(n16122) );
  XOR U19151 ( .A(n16123), .B(n16124), .Z(n16119) );
  ANDN U19152 ( .B(n16125), .A(n16126), .Z(n16123) );
  XNOR U19153 ( .A(b[1069]), .B(n16124), .Z(n16125) );
  XNOR U19154 ( .A(b[106]), .B(n16127), .Z(c[106]) );
  XNOR U19155 ( .A(b[1069]), .B(n16126), .Z(c[1069]) );
  XNOR U19156 ( .A(a[1069]), .B(n16128), .Z(n16126) );
  IV U19157 ( .A(n16124), .Z(n16128) );
  XOR U19158 ( .A(n16129), .B(n16130), .Z(n16124) );
  ANDN U19159 ( .B(n16131), .A(n16132), .Z(n16129) );
  XNOR U19160 ( .A(b[1068]), .B(n16130), .Z(n16131) );
  XNOR U19161 ( .A(b[1068]), .B(n16132), .Z(c[1068]) );
  XNOR U19162 ( .A(a[1068]), .B(n16133), .Z(n16132) );
  IV U19163 ( .A(n16130), .Z(n16133) );
  XOR U19164 ( .A(n16134), .B(n16135), .Z(n16130) );
  ANDN U19165 ( .B(n16136), .A(n16137), .Z(n16134) );
  XNOR U19166 ( .A(b[1067]), .B(n16135), .Z(n16136) );
  XNOR U19167 ( .A(b[1067]), .B(n16137), .Z(c[1067]) );
  XNOR U19168 ( .A(a[1067]), .B(n16138), .Z(n16137) );
  IV U19169 ( .A(n16135), .Z(n16138) );
  XOR U19170 ( .A(n16139), .B(n16140), .Z(n16135) );
  ANDN U19171 ( .B(n16141), .A(n16142), .Z(n16139) );
  XNOR U19172 ( .A(b[1066]), .B(n16140), .Z(n16141) );
  XNOR U19173 ( .A(b[1066]), .B(n16142), .Z(c[1066]) );
  XNOR U19174 ( .A(a[1066]), .B(n16143), .Z(n16142) );
  IV U19175 ( .A(n16140), .Z(n16143) );
  XOR U19176 ( .A(n16144), .B(n16145), .Z(n16140) );
  ANDN U19177 ( .B(n16146), .A(n16147), .Z(n16144) );
  XNOR U19178 ( .A(b[1065]), .B(n16145), .Z(n16146) );
  XNOR U19179 ( .A(b[1065]), .B(n16147), .Z(c[1065]) );
  XNOR U19180 ( .A(a[1065]), .B(n16148), .Z(n16147) );
  IV U19181 ( .A(n16145), .Z(n16148) );
  XOR U19182 ( .A(n16149), .B(n16150), .Z(n16145) );
  ANDN U19183 ( .B(n16151), .A(n16152), .Z(n16149) );
  XNOR U19184 ( .A(b[1064]), .B(n16150), .Z(n16151) );
  XNOR U19185 ( .A(b[1064]), .B(n16152), .Z(c[1064]) );
  XNOR U19186 ( .A(a[1064]), .B(n16153), .Z(n16152) );
  IV U19187 ( .A(n16150), .Z(n16153) );
  XOR U19188 ( .A(n16154), .B(n16155), .Z(n16150) );
  ANDN U19189 ( .B(n16156), .A(n16157), .Z(n16154) );
  XNOR U19190 ( .A(b[1063]), .B(n16155), .Z(n16156) );
  XNOR U19191 ( .A(b[1063]), .B(n16157), .Z(c[1063]) );
  XNOR U19192 ( .A(a[1063]), .B(n16158), .Z(n16157) );
  IV U19193 ( .A(n16155), .Z(n16158) );
  XOR U19194 ( .A(n16159), .B(n16160), .Z(n16155) );
  ANDN U19195 ( .B(n16161), .A(n16162), .Z(n16159) );
  XNOR U19196 ( .A(b[1062]), .B(n16160), .Z(n16161) );
  XNOR U19197 ( .A(b[1062]), .B(n16162), .Z(c[1062]) );
  XNOR U19198 ( .A(a[1062]), .B(n16163), .Z(n16162) );
  IV U19199 ( .A(n16160), .Z(n16163) );
  XOR U19200 ( .A(n16164), .B(n16165), .Z(n16160) );
  ANDN U19201 ( .B(n16166), .A(n16167), .Z(n16164) );
  XNOR U19202 ( .A(b[1061]), .B(n16165), .Z(n16166) );
  XNOR U19203 ( .A(b[1061]), .B(n16167), .Z(c[1061]) );
  XNOR U19204 ( .A(a[1061]), .B(n16168), .Z(n16167) );
  IV U19205 ( .A(n16165), .Z(n16168) );
  XOR U19206 ( .A(n16169), .B(n16170), .Z(n16165) );
  ANDN U19207 ( .B(n16171), .A(n16172), .Z(n16169) );
  XNOR U19208 ( .A(b[1060]), .B(n16170), .Z(n16171) );
  XNOR U19209 ( .A(b[1060]), .B(n16172), .Z(c[1060]) );
  XNOR U19210 ( .A(a[1060]), .B(n16173), .Z(n16172) );
  IV U19211 ( .A(n16170), .Z(n16173) );
  XOR U19212 ( .A(n16174), .B(n16175), .Z(n16170) );
  ANDN U19213 ( .B(n16176), .A(n16177), .Z(n16174) );
  XNOR U19214 ( .A(b[1059]), .B(n16175), .Z(n16176) );
  XNOR U19215 ( .A(b[105]), .B(n16178), .Z(c[105]) );
  XNOR U19216 ( .A(b[1059]), .B(n16177), .Z(c[1059]) );
  XNOR U19217 ( .A(a[1059]), .B(n16179), .Z(n16177) );
  IV U19218 ( .A(n16175), .Z(n16179) );
  XOR U19219 ( .A(n16180), .B(n16181), .Z(n16175) );
  ANDN U19220 ( .B(n16182), .A(n16183), .Z(n16180) );
  XNOR U19221 ( .A(b[1058]), .B(n16181), .Z(n16182) );
  XNOR U19222 ( .A(b[1058]), .B(n16183), .Z(c[1058]) );
  XNOR U19223 ( .A(a[1058]), .B(n16184), .Z(n16183) );
  IV U19224 ( .A(n16181), .Z(n16184) );
  XOR U19225 ( .A(n16185), .B(n16186), .Z(n16181) );
  ANDN U19226 ( .B(n16187), .A(n16188), .Z(n16185) );
  XNOR U19227 ( .A(b[1057]), .B(n16186), .Z(n16187) );
  XNOR U19228 ( .A(b[1057]), .B(n16188), .Z(c[1057]) );
  XNOR U19229 ( .A(a[1057]), .B(n16189), .Z(n16188) );
  IV U19230 ( .A(n16186), .Z(n16189) );
  XOR U19231 ( .A(n16190), .B(n16191), .Z(n16186) );
  ANDN U19232 ( .B(n16192), .A(n16193), .Z(n16190) );
  XNOR U19233 ( .A(b[1056]), .B(n16191), .Z(n16192) );
  XNOR U19234 ( .A(b[1056]), .B(n16193), .Z(c[1056]) );
  XNOR U19235 ( .A(a[1056]), .B(n16194), .Z(n16193) );
  IV U19236 ( .A(n16191), .Z(n16194) );
  XOR U19237 ( .A(n16195), .B(n16196), .Z(n16191) );
  ANDN U19238 ( .B(n16197), .A(n16198), .Z(n16195) );
  XNOR U19239 ( .A(b[1055]), .B(n16196), .Z(n16197) );
  XNOR U19240 ( .A(b[1055]), .B(n16198), .Z(c[1055]) );
  XNOR U19241 ( .A(a[1055]), .B(n16199), .Z(n16198) );
  IV U19242 ( .A(n16196), .Z(n16199) );
  XOR U19243 ( .A(n16200), .B(n16201), .Z(n16196) );
  ANDN U19244 ( .B(n16202), .A(n16203), .Z(n16200) );
  XNOR U19245 ( .A(b[1054]), .B(n16201), .Z(n16202) );
  XNOR U19246 ( .A(b[1054]), .B(n16203), .Z(c[1054]) );
  XNOR U19247 ( .A(a[1054]), .B(n16204), .Z(n16203) );
  IV U19248 ( .A(n16201), .Z(n16204) );
  XOR U19249 ( .A(n16205), .B(n16206), .Z(n16201) );
  ANDN U19250 ( .B(n16207), .A(n16208), .Z(n16205) );
  XNOR U19251 ( .A(b[1053]), .B(n16206), .Z(n16207) );
  XNOR U19252 ( .A(b[1053]), .B(n16208), .Z(c[1053]) );
  XNOR U19253 ( .A(a[1053]), .B(n16209), .Z(n16208) );
  IV U19254 ( .A(n16206), .Z(n16209) );
  XOR U19255 ( .A(n16210), .B(n16211), .Z(n16206) );
  ANDN U19256 ( .B(n16212), .A(n16213), .Z(n16210) );
  XNOR U19257 ( .A(b[1052]), .B(n16211), .Z(n16212) );
  XNOR U19258 ( .A(b[1052]), .B(n16213), .Z(c[1052]) );
  XNOR U19259 ( .A(a[1052]), .B(n16214), .Z(n16213) );
  IV U19260 ( .A(n16211), .Z(n16214) );
  XOR U19261 ( .A(n16215), .B(n16216), .Z(n16211) );
  ANDN U19262 ( .B(n16217), .A(n16218), .Z(n16215) );
  XNOR U19263 ( .A(b[1051]), .B(n16216), .Z(n16217) );
  XNOR U19264 ( .A(b[1051]), .B(n16218), .Z(c[1051]) );
  XNOR U19265 ( .A(a[1051]), .B(n16219), .Z(n16218) );
  IV U19266 ( .A(n16216), .Z(n16219) );
  XOR U19267 ( .A(n16220), .B(n16221), .Z(n16216) );
  ANDN U19268 ( .B(n16222), .A(n16223), .Z(n16220) );
  XNOR U19269 ( .A(b[1050]), .B(n16221), .Z(n16222) );
  XNOR U19270 ( .A(b[1050]), .B(n16223), .Z(c[1050]) );
  XNOR U19271 ( .A(a[1050]), .B(n16224), .Z(n16223) );
  IV U19272 ( .A(n16221), .Z(n16224) );
  XOR U19273 ( .A(n16225), .B(n16226), .Z(n16221) );
  ANDN U19274 ( .B(n16227), .A(n16228), .Z(n16225) );
  XNOR U19275 ( .A(b[1049]), .B(n16226), .Z(n16227) );
  XNOR U19276 ( .A(b[104]), .B(n16229), .Z(c[104]) );
  XNOR U19277 ( .A(b[1049]), .B(n16228), .Z(c[1049]) );
  XNOR U19278 ( .A(a[1049]), .B(n16230), .Z(n16228) );
  IV U19279 ( .A(n16226), .Z(n16230) );
  XOR U19280 ( .A(n16231), .B(n16232), .Z(n16226) );
  ANDN U19281 ( .B(n16233), .A(n16234), .Z(n16231) );
  XNOR U19282 ( .A(b[1048]), .B(n16232), .Z(n16233) );
  XNOR U19283 ( .A(b[1048]), .B(n16234), .Z(c[1048]) );
  XNOR U19284 ( .A(a[1048]), .B(n16235), .Z(n16234) );
  IV U19285 ( .A(n16232), .Z(n16235) );
  XOR U19286 ( .A(n16236), .B(n16237), .Z(n16232) );
  ANDN U19287 ( .B(n16238), .A(n16239), .Z(n16236) );
  XNOR U19288 ( .A(b[1047]), .B(n16237), .Z(n16238) );
  XNOR U19289 ( .A(b[1047]), .B(n16239), .Z(c[1047]) );
  XNOR U19290 ( .A(a[1047]), .B(n16240), .Z(n16239) );
  IV U19291 ( .A(n16237), .Z(n16240) );
  XOR U19292 ( .A(n16241), .B(n16242), .Z(n16237) );
  ANDN U19293 ( .B(n16243), .A(n16244), .Z(n16241) );
  XNOR U19294 ( .A(b[1046]), .B(n16242), .Z(n16243) );
  XNOR U19295 ( .A(b[1046]), .B(n16244), .Z(c[1046]) );
  XNOR U19296 ( .A(a[1046]), .B(n16245), .Z(n16244) );
  IV U19297 ( .A(n16242), .Z(n16245) );
  XOR U19298 ( .A(n16246), .B(n16247), .Z(n16242) );
  ANDN U19299 ( .B(n16248), .A(n16249), .Z(n16246) );
  XNOR U19300 ( .A(b[1045]), .B(n16247), .Z(n16248) );
  XNOR U19301 ( .A(b[1045]), .B(n16249), .Z(c[1045]) );
  XNOR U19302 ( .A(a[1045]), .B(n16250), .Z(n16249) );
  IV U19303 ( .A(n16247), .Z(n16250) );
  XOR U19304 ( .A(n16251), .B(n16252), .Z(n16247) );
  ANDN U19305 ( .B(n16253), .A(n16254), .Z(n16251) );
  XNOR U19306 ( .A(b[1044]), .B(n16252), .Z(n16253) );
  XNOR U19307 ( .A(b[1044]), .B(n16254), .Z(c[1044]) );
  XNOR U19308 ( .A(a[1044]), .B(n16255), .Z(n16254) );
  IV U19309 ( .A(n16252), .Z(n16255) );
  XOR U19310 ( .A(n16256), .B(n16257), .Z(n16252) );
  ANDN U19311 ( .B(n16258), .A(n16259), .Z(n16256) );
  XNOR U19312 ( .A(b[1043]), .B(n16257), .Z(n16258) );
  XNOR U19313 ( .A(b[1043]), .B(n16259), .Z(c[1043]) );
  XNOR U19314 ( .A(a[1043]), .B(n16260), .Z(n16259) );
  IV U19315 ( .A(n16257), .Z(n16260) );
  XOR U19316 ( .A(n16261), .B(n16262), .Z(n16257) );
  ANDN U19317 ( .B(n16263), .A(n16264), .Z(n16261) );
  XNOR U19318 ( .A(b[1042]), .B(n16262), .Z(n16263) );
  XNOR U19319 ( .A(b[1042]), .B(n16264), .Z(c[1042]) );
  XNOR U19320 ( .A(a[1042]), .B(n16265), .Z(n16264) );
  IV U19321 ( .A(n16262), .Z(n16265) );
  XOR U19322 ( .A(n16266), .B(n16267), .Z(n16262) );
  ANDN U19323 ( .B(n16268), .A(n16269), .Z(n16266) );
  XNOR U19324 ( .A(b[1041]), .B(n16267), .Z(n16268) );
  XNOR U19325 ( .A(b[1041]), .B(n16269), .Z(c[1041]) );
  XNOR U19326 ( .A(a[1041]), .B(n16270), .Z(n16269) );
  IV U19327 ( .A(n16267), .Z(n16270) );
  XOR U19328 ( .A(n16271), .B(n16272), .Z(n16267) );
  ANDN U19329 ( .B(n16273), .A(n16274), .Z(n16271) );
  XNOR U19330 ( .A(b[1040]), .B(n16272), .Z(n16273) );
  XNOR U19331 ( .A(b[1040]), .B(n16274), .Z(c[1040]) );
  XNOR U19332 ( .A(a[1040]), .B(n16275), .Z(n16274) );
  IV U19333 ( .A(n16272), .Z(n16275) );
  XOR U19334 ( .A(n16276), .B(n16277), .Z(n16272) );
  ANDN U19335 ( .B(n16278), .A(n16279), .Z(n16276) );
  XNOR U19336 ( .A(b[1039]), .B(n16277), .Z(n16278) );
  XNOR U19337 ( .A(b[103]), .B(n16280), .Z(c[103]) );
  XNOR U19338 ( .A(b[1039]), .B(n16279), .Z(c[1039]) );
  XNOR U19339 ( .A(a[1039]), .B(n16281), .Z(n16279) );
  IV U19340 ( .A(n16277), .Z(n16281) );
  XOR U19341 ( .A(n16282), .B(n16283), .Z(n16277) );
  ANDN U19342 ( .B(n16284), .A(n16285), .Z(n16282) );
  XNOR U19343 ( .A(b[1038]), .B(n16283), .Z(n16284) );
  XNOR U19344 ( .A(b[1038]), .B(n16285), .Z(c[1038]) );
  XNOR U19345 ( .A(a[1038]), .B(n16286), .Z(n16285) );
  IV U19346 ( .A(n16283), .Z(n16286) );
  XOR U19347 ( .A(n16287), .B(n16288), .Z(n16283) );
  ANDN U19348 ( .B(n16289), .A(n16290), .Z(n16287) );
  XNOR U19349 ( .A(b[1037]), .B(n16288), .Z(n16289) );
  XNOR U19350 ( .A(b[1037]), .B(n16290), .Z(c[1037]) );
  XNOR U19351 ( .A(a[1037]), .B(n16291), .Z(n16290) );
  IV U19352 ( .A(n16288), .Z(n16291) );
  XOR U19353 ( .A(n16292), .B(n16293), .Z(n16288) );
  ANDN U19354 ( .B(n16294), .A(n16295), .Z(n16292) );
  XNOR U19355 ( .A(b[1036]), .B(n16293), .Z(n16294) );
  XNOR U19356 ( .A(b[1036]), .B(n16295), .Z(c[1036]) );
  XNOR U19357 ( .A(a[1036]), .B(n16296), .Z(n16295) );
  IV U19358 ( .A(n16293), .Z(n16296) );
  XOR U19359 ( .A(n16297), .B(n16298), .Z(n16293) );
  ANDN U19360 ( .B(n16299), .A(n16300), .Z(n16297) );
  XNOR U19361 ( .A(b[1035]), .B(n16298), .Z(n16299) );
  XNOR U19362 ( .A(b[1035]), .B(n16300), .Z(c[1035]) );
  XNOR U19363 ( .A(a[1035]), .B(n16301), .Z(n16300) );
  IV U19364 ( .A(n16298), .Z(n16301) );
  XOR U19365 ( .A(n16302), .B(n16303), .Z(n16298) );
  ANDN U19366 ( .B(n16304), .A(n16305), .Z(n16302) );
  XNOR U19367 ( .A(b[1034]), .B(n16303), .Z(n16304) );
  XNOR U19368 ( .A(b[1034]), .B(n16305), .Z(c[1034]) );
  XNOR U19369 ( .A(a[1034]), .B(n16306), .Z(n16305) );
  IV U19370 ( .A(n16303), .Z(n16306) );
  XOR U19371 ( .A(n16307), .B(n16308), .Z(n16303) );
  ANDN U19372 ( .B(n16309), .A(n16310), .Z(n16307) );
  XNOR U19373 ( .A(b[1033]), .B(n16308), .Z(n16309) );
  XNOR U19374 ( .A(b[1033]), .B(n16310), .Z(c[1033]) );
  XNOR U19375 ( .A(a[1033]), .B(n16311), .Z(n16310) );
  IV U19376 ( .A(n16308), .Z(n16311) );
  XOR U19377 ( .A(n16312), .B(n16313), .Z(n16308) );
  ANDN U19378 ( .B(n16314), .A(n16315), .Z(n16312) );
  XNOR U19379 ( .A(b[1032]), .B(n16313), .Z(n16314) );
  XNOR U19380 ( .A(b[1032]), .B(n16315), .Z(c[1032]) );
  XNOR U19381 ( .A(a[1032]), .B(n16316), .Z(n16315) );
  IV U19382 ( .A(n16313), .Z(n16316) );
  XOR U19383 ( .A(n16317), .B(n16318), .Z(n16313) );
  ANDN U19384 ( .B(n16319), .A(n16320), .Z(n16317) );
  XNOR U19385 ( .A(b[1031]), .B(n16318), .Z(n16319) );
  XNOR U19386 ( .A(b[1031]), .B(n16320), .Z(c[1031]) );
  XNOR U19387 ( .A(a[1031]), .B(n16321), .Z(n16320) );
  IV U19388 ( .A(n16318), .Z(n16321) );
  XOR U19389 ( .A(n16322), .B(n16323), .Z(n16318) );
  ANDN U19390 ( .B(n16324), .A(n16325), .Z(n16322) );
  XNOR U19391 ( .A(b[1030]), .B(n16323), .Z(n16324) );
  XNOR U19392 ( .A(b[1030]), .B(n16325), .Z(c[1030]) );
  XNOR U19393 ( .A(a[1030]), .B(n16326), .Z(n16325) );
  IV U19394 ( .A(n16323), .Z(n16326) );
  XOR U19395 ( .A(n16327), .B(n16328), .Z(n16323) );
  ANDN U19396 ( .B(n16329), .A(n16330), .Z(n16327) );
  XNOR U19397 ( .A(b[1029]), .B(n16328), .Z(n16329) );
  XNOR U19398 ( .A(b[102]), .B(n16331), .Z(c[102]) );
  XNOR U19399 ( .A(b[1029]), .B(n16330), .Z(c[1029]) );
  XNOR U19400 ( .A(a[1029]), .B(n16332), .Z(n16330) );
  IV U19401 ( .A(n16328), .Z(n16332) );
  XOR U19402 ( .A(n16333), .B(n16334), .Z(n16328) );
  ANDN U19403 ( .B(n16335), .A(n16336), .Z(n16333) );
  XNOR U19404 ( .A(b[1028]), .B(n16334), .Z(n16335) );
  XNOR U19405 ( .A(b[1028]), .B(n16336), .Z(c[1028]) );
  XNOR U19406 ( .A(a[1028]), .B(n16337), .Z(n16336) );
  IV U19407 ( .A(n16334), .Z(n16337) );
  XOR U19408 ( .A(n16338), .B(n16339), .Z(n16334) );
  ANDN U19409 ( .B(n16340), .A(n16341), .Z(n16338) );
  XNOR U19410 ( .A(b[1027]), .B(n16339), .Z(n16340) );
  XNOR U19411 ( .A(b[1027]), .B(n16341), .Z(c[1027]) );
  XNOR U19412 ( .A(a[1027]), .B(n16342), .Z(n16341) );
  IV U19413 ( .A(n16339), .Z(n16342) );
  XOR U19414 ( .A(n16343), .B(n16344), .Z(n16339) );
  ANDN U19415 ( .B(n16345), .A(n16346), .Z(n16343) );
  XNOR U19416 ( .A(b[1026]), .B(n16344), .Z(n16345) );
  XNOR U19417 ( .A(b[1026]), .B(n16346), .Z(c[1026]) );
  XNOR U19418 ( .A(a[1026]), .B(n16347), .Z(n16346) );
  IV U19419 ( .A(n16344), .Z(n16347) );
  XOR U19420 ( .A(n16348), .B(n16349), .Z(n16344) );
  ANDN U19421 ( .B(n16350), .A(n16351), .Z(n16348) );
  XNOR U19422 ( .A(b[1025]), .B(n16349), .Z(n16350) );
  XNOR U19423 ( .A(b[1025]), .B(n16351), .Z(c[1025]) );
  XNOR U19424 ( .A(a[1025]), .B(n16352), .Z(n16351) );
  IV U19425 ( .A(n16349), .Z(n16352) );
  XOR U19426 ( .A(n16353), .B(n16354), .Z(n16349) );
  ANDN U19427 ( .B(n16355), .A(n16356), .Z(n16353) );
  XNOR U19428 ( .A(b[1024]), .B(n16354), .Z(n16355) );
  XNOR U19429 ( .A(b[1024]), .B(n16356), .Z(c[1024]) );
  XNOR U19430 ( .A(a[1024]), .B(n16357), .Z(n16356) );
  IV U19431 ( .A(n16354), .Z(n16357) );
  XOR U19432 ( .A(n16358), .B(n16359), .Z(n16354) );
  ANDN U19433 ( .B(n16360), .A(n16361), .Z(n16358) );
  XNOR U19434 ( .A(b[1023]), .B(n16359), .Z(n16360) );
  XNOR U19435 ( .A(b[1023]), .B(n16361), .Z(c[1023]) );
  XNOR U19436 ( .A(a[1023]), .B(n16362), .Z(n16361) );
  IV U19437 ( .A(n16359), .Z(n16362) );
  XOR U19438 ( .A(n16363), .B(n16364), .Z(n16359) );
  ANDN U19439 ( .B(n16365), .A(n16366), .Z(n16363) );
  XNOR U19440 ( .A(b[1022]), .B(n16364), .Z(n16365) );
  XNOR U19441 ( .A(b[1022]), .B(n16366), .Z(c[1022]) );
  XNOR U19442 ( .A(a[1022]), .B(n16367), .Z(n16366) );
  IV U19443 ( .A(n16364), .Z(n16367) );
  XOR U19444 ( .A(n16368), .B(n16369), .Z(n16364) );
  ANDN U19445 ( .B(n16370), .A(n16371), .Z(n16368) );
  XNOR U19446 ( .A(b[1021]), .B(n16369), .Z(n16370) );
  XNOR U19447 ( .A(b[1021]), .B(n16371), .Z(c[1021]) );
  XNOR U19448 ( .A(a[1021]), .B(n16372), .Z(n16371) );
  IV U19449 ( .A(n16369), .Z(n16372) );
  XOR U19450 ( .A(n16373), .B(n16374), .Z(n16369) );
  ANDN U19451 ( .B(n16375), .A(n16376), .Z(n16373) );
  XNOR U19452 ( .A(b[1020]), .B(n16374), .Z(n16375) );
  XNOR U19453 ( .A(b[1020]), .B(n16376), .Z(c[1020]) );
  XNOR U19454 ( .A(a[1020]), .B(n16377), .Z(n16376) );
  IV U19455 ( .A(n16374), .Z(n16377) );
  XOR U19456 ( .A(n16378), .B(n16379), .Z(n16374) );
  ANDN U19457 ( .B(n16380), .A(n16381), .Z(n16378) );
  XNOR U19458 ( .A(b[1019]), .B(n16379), .Z(n16380) );
  XNOR U19459 ( .A(b[101]), .B(n16382), .Z(c[101]) );
  XNOR U19460 ( .A(b[1019]), .B(n16381), .Z(c[1019]) );
  XNOR U19461 ( .A(a[1019]), .B(n16383), .Z(n16381) );
  IV U19462 ( .A(n16379), .Z(n16383) );
  XOR U19463 ( .A(n16384), .B(n16385), .Z(n16379) );
  ANDN U19464 ( .B(n16386), .A(n16387), .Z(n16384) );
  XNOR U19465 ( .A(b[1018]), .B(n16385), .Z(n16386) );
  XNOR U19466 ( .A(b[1018]), .B(n16387), .Z(c[1018]) );
  XNOR U19467 ( .A(a[1018]), .B(n16388), .Z(n16387) );
  IV U19468 ( .A(n16385), .Z(n16388) );
  XOR U19469 ( .A(n16389), .B(n16390), .Z(n16385) );
  ANDN U19470 ( .B(n16391), .A(n16392), .Z(n16389) );
  XNOR U19471 ( .A(b[1017]), .B(n16390), .Z(n16391) );
  XNOR U19472 ( .A(b[1017]), .B(n16392), .Z(c[1017]) );
  XNOR U19473 ( .A(a[1017]), .B(n16393), .Z(n16392) );
  IV U19474 ( .A(n16390), .Z(n16393) );
  XOR U19475 ( .A(n16394), .B(n16395), .Z(n16390) );
  ANDN U19476 ( .B(n16396), .A(n16397), .Z(n16394) );
  XNOR U19477 ( .A(b[1016]), .B(n16395), .Z(n16396) );
  XNOR U19478 ( .A(b[1016]), .B(n16397), .Z(c[1016]) );
  XNOR U19479 ( .A(a[1016]), .B(n16398), .Z(n16397) );
  IV U19480 ( .A(n16395), .Z(n16398) );
  XOR U19481 ( .A(n16399), .B(n16400), .Z(n16395) );
  ANDN U19482 ( .B(n16401), .A(n16402), .Z(n16399) );
  XNOR U19483 ( .A(b[1015]), .B(n16400), .Z(n16401) );
  XNOR U19484 ( .A(b[1015]), .B(n16402), .Z(c[1015]) );
  XNOR U19485 ( .A(a[1015]), .B(n16403), .Z(n16402) );
  IV U19486 ( .A(n16400), .Z(n16403) );
  XOR U19487 ( .A(n16404), .B(n16405), .Z(n16400) );
  ANDN U19488 ( .B(n16406), .A(n16407), .Z(n16404) );
  XNOR U19489 ( .A(b[1014]), .B(n16405), .Z(n16406) );
  XNOR U19490 ( .A(b[1014]), .B(n16407), .Z(c[1014]) );
  XNOR U19491 ( .A(a[1014]), .B(n16408), .Z(n16407) );
  IV U19492 ( .A(n16405), .Z(n16408) );
  XOR U19493 ( .A(n16409), .B(n16410), .Z(n16405) );
  ANDN U19494 ( .B(n16411), .A(n16412), .Z(n16409) );
  XNOR U19495 ( .A(b[1013]), .B(n16410), .Z(n16411) );
  XNOR U19496 ( .A(b[1013]), .B(n16412), .Z(c[1013]) );
  XNOR U19497 ( .A(a[1013]), .B(n16413), .Z(n16412) );
  IV U19498 ( .A(n16410), .Z(n16413) );
  XOR U19499 ( .A(n16414), .B(n16415), .Z(n16410) );
  ANDN U19500 ( .B(n16416), .A(n16417), .Z(n16414) );
  XNOR U19501 ( .A(b[1012]), .B(n16415), .Z(n16416) );
  XNOR U19502 ( .A(b[1012]), .B(n16417), .Z(c[1012]) );
  XNOR U19503 ( .A(a[1012]), .B(n16418), .Z(n16417) );
  IV U19504 ( .A(n16415), .Z(n16418) );
  XOR U19505 ( .A(n16419), .B(n16420), .Z(n16415) );
  ANDN U19506 ( .B(n16421), .A(n16422), .Z(n16419) );
  XNOR U19507 ( .A(b[1011]), .B(n16420), .Z(n16421) );
  XNOR U19508 ( .A(b[1011]), .B(n16422), .Z(c[1011]) );
  XNOR U19509 ( .A(a[1011]), .B(n16423), .Z(n16422) );
  IV U19510 ( .A(n16420), .Z(n16423) );
  XOR U19511 ( .A(n16424), .B(n16425), .Z(n16420) );
  ANDN U19512 ( .B(n16426), .A(n16427), .Z(n16424) );
  XNOR U19513 ( .A(b[1010]), .B(n16425), .Z(n16426) );
  XNOR U19514 ( .A(b[1010]), .B(n16427), .Z(c[1010]) );
  XNOR U19515 ( .A(a[1010]), .B(n16428), .Z(n16427) );
  IV U19516 ( .A(n16425), .Z(n16428) );
  XOR U19517 ( .A(n16429), .B(n16430), .Z(n16425) );
  ANDN U19518 ( .B(n16431), .A(n16432), .Z(n16429) );
  XNOR U19519 ( .A(b[1009]), .B(n16430), .Z(n16431) );
  XNOR U19520 ( .A(b[100]), .B(n16433), .Z(c[100]) );
  XNOR U19521 ( .A(b[1009]), .B(n16432), .Z(c[1009]) );
  XNOR U19522 ( .A(a[1009]), .B(n16434), .Z(n16432) );
  IV U19523 ( .A(n16430), .Z(n16434) );
  XOR U19524 ( .A(n16435), .B(n16436), .Z(n16430) );
  ANDN U19525 ( .B(n16437), .A(n16438), .Z(n16435) );
  XNOR U19526 ( .A(b[1008]), .B(n16436), .Z(n16437) );
  XNOR U19527 ( .A(b[1008]), .B(n16438), .Z(c[1008]) );
  XNOR U19528 ( .A(a[1008]), .B(n16439), .Z(n16438) );
  IV U19529 ( .A(n16436), .Z(n16439) );
  XOR U19530 ( .A(n16440), .B(n16441), .Z(n16436) );
  ANDN U19531 ( .B(n16442), .A(n16443), .Z(n16440) );
  XNOR U19532 ( .A(b[1007]), .B(n16441), .Z(n16442) );
  XNOR U19533 ( .A(b[1007]), .B(n16443), .Z(c[1007]) );
  XNOR U19534 ( .A(a[1007]), .B(n16444), .Z(n16443) );
  IV U19535 ( .A(n16441), .Z(n16444) );
  XOR U19536 ( .A(n16445), .B(n16446), .Z(n16441) );
  ANDN U19537 ( .B(n16447), .A(n16448), .Z(n16445) );
  XNOR U19538 ( .A(b[1006]), .B(n16446), .Z(n16447) );
  XNOR U19539 ( .A(b[1006]), .B(n16448), .Z(c[1006]) );
  XNOR U19540 ( .A(a[1006]), .B(n16449), .Z(n16448) );
  IV U19541 ( .A(n16446), .Z(n16449) );
  XOR U19542 ( .A(n16450), .B(n16451), .Z(n16446) );
  ANDN U19543 ( .B(n16452), .A(n16453), .Z(n16450) );
  XNOR U19544 ( .A(b[1005]), .B(n16451), .Z(n16452) );
  XNOR U19545 ( .A(b[1005]), .B(n16453), .Z(c[1005]) );
  XNOR U19546 ( .A(a[1005]), .B(n16454), .Z(n16453) );
  IV U19547 ( .A(n16451), .Z(n16454) );
  XOR U19548 ( .A(n16455), .B(n16456), .Z(n16451) );
  ANDN U19549 ( .B(n16457), .A(n16458), .Z(n16455) );
  XNOR U19550 ( .A(b[1004]), .B(n16456), .Z(n16457) );
  XNOR U19551 ( .A(b[1004]), .B(n16458), .Z(c[1004]) );
  XNOR U19552 ( .A(a[1004]), .B(n16459), .Z(n16458) );
  IV U19553 ( .A(n16456), .Z(n16459) );
  XOR U19554 ( .A(n16460), .B(n16461), .Z(n16456) );
  ANDN U19555 ( .B(n16462), .A(n16463), .Z(n16460) );
  XNOR U19556 ( .A(b[1003]), .B(n16461), .Z(n16462) );
  XNOR U19557 ( .A(b[1003]), .B(n16463), .Z(c[1003]) );
  XNOR U19558 ( .A(a[1003]), .B(n16464), .Z(n16463) );
  IV U19559 ( .A(n16461), .Z(n16464) );
  XOR U19560 ( .A(n16465), .B(n16466), .Z(n16461) );
  ANDN U19561 ( .B(n16467), .A(n16468), .Z(n16465) );
  XNOR U19562 ( .A(b[1002]), .B(n16466), .Z(n16467) );
  XNOR U19563 ( .A(b[1002]), .B(n16468), .Z(c[1002]) );
  XNOR U19564 ( .A(a[1002]), .B(n16469), .Z(n16468) );
  IV U19565 ( .A(n16466), .Z(n16469) );
  XOR U19566 ( .A(n16470), .B(n16471), .Z(n16466) );
  ANDN U19567 ( .B(n16472), .A(n16473), .Z(n16470) );
  XNOR U19568 ( .A(b[1001]), .B(n16471), .Z(n16472) );
  XNOR U19569 ( .A(b[1001]), .B(n16473), .Z(c[1001]) );
  XNOR U19570 ( .A(a[1001]), .B(n16474), .Z(n16473) );
  IV U19571 ( .A(n16471), .Z(n16474) );
  XOR U19572 ( .A(n16475), .B(n16476), .Z(n16471) );
  ANDN U19573 ( .B(n16477), .A(n16478), .Z(n16475) );
  XNOR U19574 ( .A(b[1000]), .B(n16476), .Z(n16477) );
  XNOR U19575 ( .A(b[1000]), .B(n16478), .Z(c[1000]) );
  XNOR U19576 ( .A(a[1000]), .B(n16479), .Z(n16478) );
  IV U19577 ( .A(n16476), .Z(n16479) );
  XOR U19578 ( .A(n16480), .B(n16481), .Z(n16476) );
  ANDN U19579 ( .B(n16482), .A(n8), .Z(n16480) );
  XNOR U19580 ( .A(a[999]), .B(n16483), .Z(n8) );
  IV U19581 ( .A(n16481), .Z(n16483) );
  XNOR U19582 ( .A(b[999]), .B(n16481), .Z(n16482) );
  XOR U19583 ( .A(n16484), .B(n16485), .Z(n16481) );
  ANDN U19584 ( .B(n16486), .A(n9), .Z(n16484) );
  XNOR U19585 ( .A(a[998]), .B(n16487), .Z(n9) );
  IV U19586 ( .A(n16485), .Z(n16487) );
  XNOR U19587 ( .A(b[998]), .B(n16485), .Z(n16486) );
  XOR U19588 ( .A(n16488), .B(n16489), .Z(n16485) );
  ANDN U19589 ( .B(n16490), .A(n10), .Z(n16488) );
  XNOR U19590 ( .A(a[997]), .B(n16491), .Z(n10) );
  IV U19591 ( .A(n16489), .Z(n16491) );
  XNOR U19592 ( .A(b[997]), .B(n16489), .Z(n16490) );
  XOR U19593 ( .A(n16492), .B(n16493), .Z(n16489) );
  ANDN U19594 ( .B(n16494), .A(n11), .Z(n16492) );
  XNOR U19595 ( .A(a[996]), .B(n16495), .Z(n11) );
  IV U19596 ( .A(n16493), .Z(n16495) );
  XNOR U19597 ( .A(b[996]), .B(n16493), .Z(n16494) );
  XOR U19598 ( .A(n16496), .B(n16497), .Z(n16493) );
  ANDN U19599 ( .B(n16498), .A(n12), .Z(n16496) );
  XNOR U19600 ( .A(a[995]), .B(n16499), .Z(n12) );
  IV U19601 ( .A(n16497), .Z(n16499) );
  XNOR U19602 ( .A(b[995]), .B(n16497), .Z(n16498) );
  XOR U19603 ( .A(n16500), .B(n16501), .Z(n16497) );
  ANDN U19604 ( .B(n16502), .A(n13), .Z(n16500) );
  XNOR U19605 ( .A(a[994]), .B(n16503), .Z(n13) );
  IV U19606 ( .A(n16501), .Z(n16503) );
  XNOR U19607 ( .A(b[994]), .B(n16501), .Z(n16502) );
  XOR U19608 ( .A(n16504), .B(n16505), .Z(n16501) );
  ANDN U19609 ( .B(n16506), .A(n14), .Z(n16504) );
  XNOR U19610 ( .A(a[993]), .B(n16507), .Z(n14) );
  IV U19611 ( .A(n16505), .Z(n16507) );
  XNOR U19612 ( .A(b[993]), .B(n16505), .Z(n16506) );
  XOR U19613 ( .A(n16508), .B(n16509), .Z(n16505) );
  ANDN U19614 ( .B(n16510), .A(n15), .Z(n16508) );
  XNOR U19615 ( .A(a[992]), .B(n16511), .Z(n15) );
  IV U19616 ( .A(n16509), .Z(n16511) );
  XNOR U19617 ( .A(b[992]), .B(n16509), .Z(n16510) );
  XOR U19618 ( .A(n16512), .B(n16513), .Z(n16509) );
  ANDN U19619 ( .B(n16514), .A(n16), .Z(n16512) );
  XNOR U19620 ( .A(a[991]), .B(n16515), .Z(n16) );
  IV U19621 ( .A(n16513), .Z(n16515) );
  XNOR U19622 ( .A(b[991]), .B(n16513), .Z(n16514) );
  XOR U19623 ( .A(n16516), .B(n16517), .Z(n16513) );
  ANDN U19624 ( .B(n16518), .A(n17), .Z(n16516) );
  XNOR U19625 ( .A(a[990]), .B(n16519), .Z(n17) );
  IV U19626 ( .A(n16517), .Z(n16519) );
  XNOR U19627 ( .A(b[990]), .B(n16517), .Z(n16518) );
  XOR U19628 ( .A(n16520), .B(n16521), .Z(n16517) );
  ANDN U19629 ( .B(n16522), .A(n19), .Z(n16520) );
  XNOR U19630 ( .A(a[989]), .B(n16523), .Z(n19) );
  IV U19631 ( .A(n16521), .Z(n16523) );
  XNOR U19632 ( .A(b[989]), .B(n16521), .Z(n16522) );
  XOR U19633 ( .A(n16524), .B(n16525), .Z(n16521) );
  ANDN U19634 ( .B(n16526), .A(n20), .Z(n16524) );
  XNOR U19635 ( .A(a[988]), .B(n16527), .Z(n20) );
  IV U19636 ( .A(n16525), .Z(n16527) );
  XNOR U19637 ( .A(b[988]), .B(n16525), .Z(n16526) );
  XOR U19638 ( .A(n16528), .B(n16529), .Z(n16525) );
  ANDN U19639 ( .B(n16530), .A(n21), .Z(n16528) );
  XNOR U19640 ( .A(a[987]), .B(n16531), .Z(n21) );
  IV U19641 ( .A(n16529), .Z(n16531) );
  XNOR U19642 ( .A(b[987]), .B(n16529), .Z(n16530) );
  XOR U19643 ( .A(n16532), .B(n16533), .Z(n16529) );
  ANDN U19644 ( .B(n16534), .A(n22), .Z(n16532) );
  XNOR U19645 ( .A(a[986]), .B(n16535), .Z(n22) );
  IV U19646 ( .A(n16533), .Z(n16535) );
  XNOR U19647 ( .A(b[986]), .B(n16533), .Z(n16534) );
  XOR U19648 ( .A(n16536), .B(n16537), .Z(n16533) );
  ANDN U19649 ( .B(n16538), .A(n23), .Z(n16536) );
  XNOR U19650 ( .A(a[985]), .B(n16539), .Z(n23) );
  IV U19651 ( .A(n16537), .Z(n16539) );
  XNOR U19652 ( .A(b[985]), .B(n16537), .Z(n16538) );
  XOR U19653 ( .A(n16540), .B(n16541), .Z(n16537) );
  ANDN U19654 ( .B(n16542), .A(n24), .Z(n16540) );
  XNOR U19655 ( .A(a[984]), .B(n16543), .Z(n24) );
  IV U19656 ( .A(n16541), .Z(n16543) );
  XNOR U19657 ( .A(b[984]), .B(n16541), .Z(n16542) );
  XOR U19658 ( .A(n16544), .B(n16545), .Z(n16541) );
  ANDN U19659 ( .B(n16546), .A(n25), .Z(n16544) );
  XNOR U19660 ( .A(a[983]), .B(n16547), .Z(n25) );
  IV U19661 ( .A(n16545), .Z(n16547) );
  XNOR U19662 ( .A(b[983]), .B(n16545), .Z(n16546) );
  XOR U19663 ( .A(n16548), .B(n16549), .Z(n16545) );
  ANDN U19664 ( .B(n16550), .A(n26), .Z(n16548) );
  XNOR U19665 ( .A(a[982]), .B(n16551), .Z(n26) );
  IV U19666 ( .A(n16549), .Z(n16551) );
  XNOR U19667 ( .A(b[982]), .B(n16549), .Z(n16550) );
  XOR U19668 ( .A(n16552), .B(n16553), .Z(n16549) );
  ANDN U19669 ( .B(n16554), .A(n27), .Z(n16552) );
  XNOR U19670 ( .A(a[981]), .B(n16555), .Z(n27) );
  IV U19671 ( .A(n16553), .Z(n16555) );
  XNOR U19672 ( .A(b[981]), .B(n16553), .Z(n16554) );
  XOR U19673 ( .A(n16556), .B(n16557), .Z(n16553) );
  ANDN U19674 ( .B(n16558), .A(n28), .Z(n16556) );
  XNOR U19675 ( .A(a[980]), .B(n16559), .Z(n28) );
  IV U19676 ( .A(n16557), .Z(n16559) );
  XNOR U19677 ( .A(b[980]), .B(n16557), .Z(n16558) );
  XOR U19678 ( .A(n16560), .B(n16561), .Z(n16557) );
  ANDN U19679 ( .B(n16562), .A(n30), .Z(n16560) );
  XNOR U19680 ( .A(a[979]), .B(n16563), .Z(n30) );
  IV U19681 ( .A(n16561), .Z(n16563) );
  XNOR U19682 ( .A(b[979]), .B(n16561), .Z(n16562) );
  XOR U19683 ( .A(n16564), .B(n16565), .Z(n16561) );
  ANDN U19684 ( .B(n16566), .A(n31), .Z(n16564) );
  XNOR U19685 ( .A(a[978]), .B(n16567), .Z(n31) );
  IV U19686 ( .A(n16565), .Z(n16567) );
  XNOR U19687 ( .A(b[978]), .B(n16565), .Z(n16566) );
  XOR U19688 ( .A(n16568), .B(n16569), .Z(n16565) );
  ANDN U19689 ( .B(n16570), .A(n32), .Z(n16568) );
  XNOR U19690 ( .A(a[977]), .B(n16571), .Z(n32) );
  IV U19691 ( .A(n16569), .Z(n16571) );
  XNOR U19692 ( .A(b[977]), .B(n16569), .Z(n16570) );
  XOR U19693 ( .A(n16572), .B(n16573), .Z(n16569) );
  ANDN U19694 ( .B(n16574), .A(n33), .Z(n16572) );
  XNOR U19695 ( .A(a[976]), .B(n16575), .Z(n33) );
  IV U19696 ( .A(n16573), .Z(n16575) );
  XNOR U19697 ( .A(b[976]), .B(n16573), .Z(n16574) );
  XOR U19698 ( .A(n16576), .B(n16577), .Z(n16573) );
  ANDN U19699 ( .B(n16578), .A(n34), .Z(n16576) );
  XNOR U19700 ( .A(a[975]), .B(n16579), .Z(n34) );
  IV U19701 ( .A(n16577), .Z(n16579) );
  XNOR U19702 ( .A(b[975]), .B(n16577), .Z(n16578) );
  XOR U19703 ( .A(n16580), .B(n16581), .Z(n16577) );
  ANDN U19704 ( .B(n16582), .A(n35), .Z(n16580) );
  XNOR U19705 ( .A(a[974]), .B(n16583), .Z(n35) );
  IV U19706 ( .A(n16581), .Z(n16583) );
  XNOR U19707 ( .A(b[974]), .B(n16581), .Z(n16582) );
  XOR U19708 ( .A(n16584), .B(n16585), .Z(n16581) );
  ANDN U19709 ( .B(n16586), .A(n36), .Z(n16584) );
  XNOR U19710 ( .A(a[973]), .B(n16587), .Z(n36) );
  IV U19711 ( .A(n16585), .Z(n16587) );
  XNOR U19712 ( .A(b[973]), .B(n16585), .Z(n16586) );
  XOR U19713 ( .A(n16588), .B(n16589), .Z(n16585) );
  ANDN U19714 ( .B(n16590), .A(n37), .Z(n16588) );
  XNOR U19715 ( .A(a[972]), .B(n16591), .Z(n37) );
  IV U19716 ( .A(n16589), .Z(n16591) );
  XNOR U19717 ( .A(b[972]), .B(n16589), .Z(n16590) );
  XOR U19718 ( .A(n16592), .B(n16593), .Z(n16589) );
  ANDN U19719 ( .B(n16594), .A(n38), .Z(n16592) );
  XNOR U19720 ( .A(a[971]), .B(n16595), .Z(n38) );
  IV U19721 ( .A(n16593), .Z(n16595) );
  XNOR U19722 ( .A(b[971]), .B(n16593), .Z(n16594) );
  XOR U19723 ( .A(n16596), .B(n16597), .Z(n16593) );
  ANDN U19724 ( .B(n16598), .A(n39), .Z(n16596) );
  XNOR U19725 ( .A(a[970]), .B(n16599), .Z(n39) );
  IV U19726 ( .A(n16597), .Z(n16599) );
  XNOR U19727 ( .A(b[970]), .B(n16597), .Z(n16598) );
  XOR U19728 ( .A(n16600), .B(n16601), .Z(n16597) );
  ANDN U19729 ( .B(n16602), .A(n41), .Z(n16600) );
  XNOR U19730 ( .A(a[969]), .B(n16603), .Z(n41) );
  IV U19731 ( .A(n16601), .Z(n16603) );
  XNOR U19732 ( .A(b[969]), .B(n16601), .Z(n16602) );
  XOR U19733 ( .A(n16604), .B(n16605), .Z(n16601) );
  ANDN U19734 ( .B(n16606), .A(n42), .Z(n16604) );
  XNOR U19735 ( .A(a[968]), .B(n16607), .Z(n42) );
  IV U19736 ( .A(n16605), .Z(n16607) );
  XNOR U19737 ( .A(b[968]), .B(n16605), .Z(n16606) );
  XOR U19738 ( .A(n16608), .B(n16609), .Z(n16605) );
  ANDN U19739 ( .B(n16610), .A(n43), .Z(n16608) );
  XNOR U19740 ( .A(a[967]), .B(n16611), .Z(n43) );
  IV U19741 ( .A(n16609), .Z(n16611) );
  XNOR U19742 ( .A(b[967]), .B(n16609), .Z(n16610) );
  XOR U19743 ( .A(n16612), .B(n16613), .Z(n16609) );
  ANDN U19744 ( .B(n16614), .A(n44), .Z(n16612) );
  XNOR U19745 ( .A(a[966]), .B(n16615), .Z(n44) );
  IV U19746 ( .A(n16613), .Z(n16615) );
  XNOR U19747 ( .A(b[966]), .B(n16613), .Z(n16614) );
  XOR U19748 ( .A(n16616), .B(n16617), .Z(n16613) );
  ANDN U19749 ( .B(n16618), .A(n45), .Z(n16616) );
  XNOR U19750 ( .A(a[965]), .B(n16619), .Z(n45) );
  IV U19751 ( .A(n16617), .Z(n16619) );
  XNOR U19752 ( .A(b[965]), .B(n16617), .Z(n16618) );
  XOR U19753 ( .A(n16620), .B(n16621), .Z(n16617) );
  ANDN U19754 ( .B(n16622), .A(n46), .Z(n16620) );
  XNOR U19755 ( .A(a[964]), .B(n16623), .Z(n46) );
  IV U19756 ( .A(n16621), .Z(n16623) );
  XNOR U19757 ( .A(b[964]), .B(n16621), .Z(n16622) );
  XOR U19758 ( .A(n16624), .B(n16625), .Z(n16621) );
  ANDN U19759 ( .B(n16626), .A(n47), .Z(n16624) );
  XNOR U19760 ( .A(a[963]), .B(n16627), .Z(n47) );
  IV U19761 ( .A(n16625), .Z(n16627) );
  XNOR U19762 ( .A(b[963]), .B(n16625), .Z(n16626) );
  XOR U19763 ( .A(n16628), .B(n16629), .Z(n16625) );
  ANDN U19764 ( .B(n16630), .A(n48), .Z(n16628) );
  XNOR U19765 ( .A(a[962]), .B(n16631), .Z(n48) );
  IV U19766 ( .A(n16629), .Z(n16631) );
  XNOR U19767 ( .A(b[962]), .B(n16629), .Z(n16630) );
  XOR U19768 ( .A(n16632), .B(n16633), .Z(n16629) );
  ANDN U19769 ( .B(n16634), .A(n49), .Z(n16632) );
  XNOR U19770 ( .A(a[961]), .B(n16635), .Z(n49) );
  IV U19771 ( .A(n16633), .Z(n16635) );
  XNOR U19772 ( .A(b[961]), .B(n16633), .Z(n16634) );
  XOR U19773 ( .A(n16636), .B(n16637), .Z(n16633) );
  ANDN U19774 ( .B(n16638), .A(n50), .Z(n16636) );
  XNOR U19775 ( .A(a[960]), .B(n16639), .Z(n50) );
  IV U19776 ( .A(n16637), .Z(n16639) );
  XNOR U19777 ( .A(b[960]), .B(n16637), .Z(n16638) );
  XOR U19778 ( .A(n16640), .B(n16641), .Z(n16637) );
  ANDN U19779 ( .B(n16642), .A(n52), .Z(n16640) );
  XNOR U19780 ( .A(a[959]), .B(n16643), .Z(n52) );
  IV U19781 ( .A(n16641), .Z(n16643) );
  XNOR U19782 ( .A(b[959]), .B(n16641), .Z(n16642) );
  XOR U19783 ( .A(n16644), .B(n16645), .Z(n16641) );
  ANDN U19784 ( .B(n16646), .A(n53), .Z(n16644) );
  XNOR U19785 ( .A(a[958]), .B(n16647), .Z(n53) );
  IV U19786 ( .A(n16645), .Z(n16647) );
  XNOR U19787 ( .A(b[958]), .B(n16645), .Z(n16646) );
  XOR U19788 ( .A(n16648), .B(n16649), .Z(n16645) );
  ANDN U19789 ( .B(n16650), .A(n54), .Z(n16648) );
  XNOR U19790 ( .A(a[957]), .B(n16651), .Z(n54) );
  IV U19791 ( .A(n16649), .Z(n16651) );
  XNOR U19792 ( .A(b[957]), .B(n16649), .Z(n16650) );
  XOR U19793 ( .A(n16652), .B(n16653), .Z(n16649) );
  ANDN U19794 ( .B(n16654), .A(n55), .Z(n16652) );
  XNOR U19795 ( .A(a[956]), .B(n16655), .Z(n55) );
  IV U19796 ( .A(n16653), .Z(n16655) );
  XNOR U19797 ( .A(b[956]), .B(n16653), .Z(n16654) );
  XOR U19798 ( .A(n16656), .B(n16657), .Z(n16653) );
  ANDN U19799 ( .B(n16658), .A(n56), .Z(n16656) );
  XNOR U19800 ( .A(a[955]), .B(n16659), .Z(n56) );
  IV U19801 ( .A(n16657), .Z(n16659) );
  XNOR U19802 ( .A(b[955]), .B(n16657), .Z(n16658) );
  XOR U19803 ( .A(n16660), .B(n16661), .Z(n16657) );
  ANDN U19804 ( .B(n16662), .A(n57), .Z(n16660) );
  XNOR U19805 ( .A(a[954]), .B(n16663), .Z(n57) );
  IV U19806 ( .A(n16661), .Z(n16663) );
  XNOR U19807 ( .A(b[954]), .B(n16661), .Z(n16662) );
  XOR U19808 ( .A(n16664), .B(n16665), .Z(n16661) );
  ANDN U19809 ( .B(n16666), .A(n58), .Z(n16664) );
  XNOR U19810 ( .A(a[953]), .B(n16667), .Z(n58) );
  IV U19811 ( .A(n16665), .Z(n16667) );
  XNOR U19812 ( .A(b[953]), .B(n16665), .Z(n16666) );
  XOR U19813 ( .A(n16668), .B(n16669), .Z(n16665) );
  ANDN U19814 ( .B(n16670), .A(n59), .Z(n16668) );
  XNOR U19815 ( .A(a[952]), .B(n16671), .Z(n59) );
  IV U19816 ( .A(n16669), .Z(n16671) );
  XNOR U19817 ( .A(b[952]), .B(n16669), .Z(n16670) );
  XOR U19818 ( .A(n16672), .B(n16673), .Z(n16669) );
  ANDN U19819 ( .B(n16674), .A(n60), .Z(n16672) );
  XNOR U19820 ( .A(a[951]), .B(n16675), .Z(n60) );
  IV U19821 ( .A(n16673), .Z(n16675) );
  XNOR U19822 ( .A(b[951]), .B(n16673), .Z(n16674) );
  XOR U19823 ( .A(n16676), .B(n16677), .Z(n16673) );
  ANDN U19824 ( .B(n16678), .A(n61), .Z(n16676) );
  XNOR U19825 ( .A(a[950]), .B(n16679), .Z(n61) );
  IV U19826 ( .A(n16677), .Z(n16679) );
  XNOR U19827 ( .A(b[950]), .B(n16677), .Z(n16678) );
  XOR U19828 ( .A(n16680), .B(n16681), .Z(n16677) );
  ANDN U19829 ( .B(n16682), .A(n63), .Z(n16680) );
  XNOR U19830 ( .A(a[949]), .B(n16683), .Z(n63) );
  IV U19831 ( .A(n16681), .Z(n16683) );
  XNOR U19832 ( .A(b[949]), .B(n16681), .Z(n16682) );
  XOR U19833 ( .A(n16684), .B(n16685), .Z(n16681) );
  ANDN U19834 ( .B(n16686), .A(n64), .Z(n16684) );
  XNOR U19835 ( .A(a[948]), .B(n16687), .Z(n64) );
  IV U19836 ( .A(n16685), .Z(n16687) );
  XNOR U19837 ( .A(b[948]), .B(n16685), .Z(n16686) );
  XOR U19838 ( .A(n16688), .B(n16689), .Z(n16685) );
  ANDN U19839 ( .B(n16690), .A(n65), .Z(n16688) );
  XNOR U19840 ( .A(a[947]), .B(n16691), .Z(n65) );
  IV U19841 ( .A(n16689), .Z(n16691) );
  XNOR U19842 ( .A(b[947]), .B(n16689), .Z(n16690) );
  XOR U19843 ( .A(n16692), .B(n16693), .Z(n16689) );
  ANDN U19844 ( .B(n16694), .A(n66), .Z(n16692) );
  XNOR U19845 ( .A(a[946]), .B(n16695), .Z(n66) );
  IV U19846 ( .A(n16693), .Z(n16695) );
  XNOR U19847 ( .A(b[946]), .B(n16693), .Z(n16694) );
  XOR U19848 ( .A(n16696), .B(n16697), .Z(n16693) );
  ANDN U19849 ( .B(n16698), .A(n67), .Z(n16696) );
  XNOR U19850 ( .A(a[945]), .B(n16699), .Z(n67) );
  IV U19851 ( .A(n16697), .Z(n16699) );
  XNOR U19852 ( .A(b[945]), .B(n16697), .Z(n16698) );
  XOR U19853 ( .A(n16700), .B(n16701), .Z(n16697) );
  ANDN U19854 ( .B(n16702), .A(n68), .Z(n16700) );
  XNOR U19855 ( .A(a[944]), .B(n16703), .Z(n68) );
  IV U19856 ( .A(n16701), .Z(n16703) );
  XNOR U19857 ( .A(b[944]), .B(n16701), .Z(n16702) );
  XOR U19858 ( .A(n16704), .B(n16705), .Z(n16701) );
  ANDN U19859 ( .B(n16706), .A(n69), .Z(n16704) );
  XNOR U19860 ( .A(a[943]), .B(n16707), .Z(n69) );
  IV U19861 ( .A(n16705), .Z(n16707) );
  XNOR U19862 ( .A(b[943]), .B(n16705), .Z(n16706) );
  XOR U19863 ( .A(n16708), .B(n16709), .Z(n16705) );
  ANDN U19864 ( .B(n16710), .A(n70), .Z(n16708) );
  XNOR U19865 ( .A(a[942]), .B(n16711), .Z(n70) );
  IV U19866 ( .A(n16709), .Z(n16711) );
  XNOR U19867 ( .A(b[942]), .B(n16709), .Z(n16710) );
  XOR U19868 ( .A(n16712), .B(n16713), .Z(n16709) );
  ANDN U19869 ( .B(n16714), .A(n71), .Z(n16712) );
  XNOR U19870 ( .A(a[941]), .B(n16715), .Z(n71) );
  IV U19871 ( .A(n16713), .Z(n16715) );
  XNOR U19872 ( .A(b[941]), .B(n16713), .Z(n16714) );
  XOR U19873 ( .A(n16716), .B(n16717), .Z(n16713) );
  ANDN U19874 ( .B(n16718), .A(n72), .Z(n16716) );
  XNOR U19875 ( .A(a[940]), .B(n16719), .Z(n72) );
  IV U19876 ( .A(n16717), .Z(n16719) );
  XNOR U19877 ( .A(b[940]), .B(n16717), .Z(n16718) );
  XOR U19878 ( .A(n16720), .B(n16721), .Z(n16717) );
  ANDN U19879 ( .B(n16722), .A(n74), .Z(n16720) );
  XNOR U19880 ( .A(a[939]), .B(n16723), .Z(n74) );
  IV U19881 ( .A(n16721), .Z(n16723) );
  XNOR U19882 ( .A(b[939]), .B(n16721), .Z(n16722) );
  XOR U19883 ( .A(n16724), .B(n16725), .Z(n16721) );
  ANDN U19884 ( .B(n16726), .A(n75), .Z(n16724) );
  XNOR U19885 ( .A(a[938]), .B(n16727), .Z(n75) );
  IV U19886 ( .A(n16725), .Z(n16727) );
  XNOR U19887 ( .A(b[938]), .B(n16725), .Z(n16726) );
  XOR U19888 ( .A(n16728), .B(n16729), .Z(n16725) );
  ANDN U19889 ( .B(n16730), .A(n76), .Z(n16728) );
  XNOR U19890 ( .A(a[937]), .B(n16731), .Z(n76) );
  IV U19891 ( .A(n16729), .Z(n16731) );
  XNOR U19892 ( .A(b[937]), .B(n16729), .Z(n16730) );
  XOR U19893 ( .A(n16732), .B(n16733), .Z(n16729) );
  ANDN U19894 ( .B(n16734), .A(n77), .Z(n16732) );
  XNOR U19895 ( .A(a[936]), .B(n16735), .Z(n77) );
  IV U19896 ( .A(n16733), .Z(n16735) );
  XNOR U19897 ( .A(b[936]), .B(n16733), .Z(n16734) );
  XOR U19898 ( .A(n16736), .B(n16737), .Z(n16733) );
  ANDN U19899 ( .B(n16738), .A(n78), .Z(n16736) );
  XNOR U19900 ( .A(a[935]), .B(n16739), .Z(n78) );
  IV U19901 ( .A(n16737), .Z(n16739) );
  XNOR U19902 ( .A(b[935]), .B(n16737), .Z(n16738) );
  XOR U19903 ( .A(n16740), .B(n16741), .Z(n16737) );
  ANDN U19904 ( .B(n16742), .A(n79), .Z(n16740) );
  XNOR U19905 ( .A(a[934]), .B(n16743), .Z(n79) );
  IV U19906 ( .A(n16741), .Z(n16743) );
  XNOR U19907 ( .A(b[934]), .B(n16741), .Z(n16742) );
  XOR U19908 ( .A(n16744), .B(n16745), .Z(n16741) );
  ANDN U19909 ( .B(n16746), .A(n80), .Z(n16744) );
  XNOR U19910 ( .A(a[933]), .B(n16747), .Z(n80) );
  IV U19911 ( .A(n16745), .Z(n16747) );
  XNOR U19912 ( .A(b[933]), .B(n16745), .Z(n16746) );
  XOR U19913 ( .A(n16748), .B(n16749), .Z(n16745) );
  ANDN U19914 ( .B(n16750), .A(n81), .Z(n16748) );
  XNOR U19915 ( .A(a[932]), .B(n16751), .Z(n81) );
  IV U19916 ( .A(n16749), .Z(n16751) );
  XNOR U19917 ( .A(b[932]), .B(n16749), .Z(n16750) );
  XOR U19918 ( .A(n16752), .B(n16753), .Z(n16749) );
  ANDN U19919 ( .B(n16754), .A(n82), .Z(n16752) );
  XNOR U19920 ( .A(a[931]), .B(n16755), .Z(n82) );
  IV U19921 ( .A(n16753), .Z(n16755) );
  XNOR U19922 ( .A(b[931]), .B(n16753), .Z(n16754) );
  XOR U19923 ( .A(n16756), .B(n16757), .Z(n16753) );
  ANDN U19924 ( .B(n16758), .A(n83), .Z(n16756) );
  XNOR U19925 ( .A(a[930]), .B(n16759), .Z(n83) );
  IV U19926 ( .A(n16757), .Z(n16759) );
  XNOR U19927 ( .A(b[930]), .B(n16757), .Z(n16758) );
  XOR U19928 ( .A(n16760), .B(n16761), .Z(n16757) );
  ANDN U19929 ( .B(n16762), .A(n85), .Z(n16760) );
  XNOR U19930 ( .A(a[929]), .B(n16763), .Z(n85) );
  IV U19931 ( .A(n16761), .Z(n16763) );
  XNOR U19932 ( .A(b[929]), .B(n16761), .Z(n16762) );
  XOR U19933 ( .A(n16764), .B(n16765), .Z(n16761) );
  ANDN U19934 ( .B(n16766), .A(n86), .Z(n16764) );
  XNOR U19935 ( .A(a[928]), .B(n16767), .Z(n86) );
  IV U19936 ( .A(n16765), .Z(n16767) );
  XNOR U19937 ( .A(b[928]), .B(n16765), .Z(n16766) );
  XOR U19938 ( .A(n16768), .B(n16769), .Z(n16765) );
  ANDN U19939 ( .B(n16770), .A(n87), .Z(n16768) );
  XNOR U19940 ( .A(a[927]), .B(n16771), .Z(n87) );
  IV U19941 ( .A(n16769), .Z(n16771) );
  XNOR U19942 ( .A(b[927]), .B(n16769), .Z(n16770) );
  XOR U19943 ( .A(n16772), .B(n16773), .Z(n16769) );
  ANDN U19944 ( .B(n16774), .A(n88), .Z(n16772) );
  XNOR U19945 ( .A(a[926]), .B(n16775), .Z(n88) );
  IV U19946 ( .A(n16773), .Z(n16775) );
  XNOR U19947 ( .A(b[926]), .B(n16773), .Z(n16774) );
  XOR U19948 ( .A(n16776), .B(n16777), .Z(n16773) );
  ANDN U19949 ( .B(n16778), .A(n89), .Z(n16776) );
  XNOR U19950 ( .A(a[925]), .B(n16779), .Z(n89) );
  IV U19951 ( .A(n16777), .Z(n16779) );
  XNOR U19952 ( .A(b[925]), .B(n16777), .Z(n16778) );
  XOR U19953 ( .A(n16780), .B(n16781), .Z(n16777) );
  ANDN U19954 ( .B(n16782), .A(n90), .Z(n16780) );
  XNOR U19955 ( .A(a[924]), .B(n16783), .Z(n90) );
  IV U19956 ( .A(n16781), .Z(n16783) );
  XNOR U19957 ( .A(b[924]), .B(n16781), .Z(n16782) );
  XOR U19958 ( .A(n16784), .B(n16785), .Z(n16781) );
  ANDN U19959 ( .B(n16786), .A(n91), .Z(n16784) );
  XNOR U19960 ( .A(a[923]), .B(n16787), .Z(n91) );
  IV U19961 ( .A(n16785), .Z(n16787) );
  XNOR U19962 ( .A(b[923]), .B(n16785), .Z(n16786) );
  XOR U19963 ( .A(n16788), .B(n16789), .Z(n16785) );
  ANDN U19964 ( .B(n16790), .A(n92), .Z(n16788) );
  XNOR U19965 ( .A(a[922]), .B(n16791), .Z(n92) );
  IV U19966 ( .A(n16789), .Z(n16791) );
  XNOR U19967 ( .A(b[922]), .B(n16789), .Z(n16790) );
  XOR U19968 ( .A(n16792), .B(n16793), .Z(n16789) );
  ANDN U19969 ( .B(n16794), .A(n93), .Z(n16792) );
  XNOR U19970 ( .A(a[921]), .B(n16795), .Z(n93) );
  IV U19971 ( .A(n16793), .Z(n16795) );
  XNOR U19972 ( .A(b[921]), .B(n16793), .Z(n16794) );
  XOR U19973 ( .A(n16796), .B(n16797), .Z(n16793) );
  ANDN U19974 ( .B(n16798), .A(n94), .Z(n16796) );
  XNOR U19975 ( .A(a[920]), .B(n16799), .Z(n94) );
  IV U19976 ( .A(n16797), .Z(n16799) );
  XNOR U19977 ( .A(b[920]), .B(n16797), .Z(n16798) );
  XOR U19978 ( .A(n16800), .B(n16801), .Z(n16797) );
  ANDN U19979 ( .B(n16802), .A(n96), .Z(n16800) );
  XNOR U19980 ( .A(a[919]), .B(n16803), .Z(n96) );
  IV U19981 ( .A(n16801), .Z(n16803) );
  XNOR U19982 ( .A(b[919]), .B(n16801), .Z(n16802) );
  XOR U19983 ( .A(n16804), .B(n16805), .Z(n16801) );
  ANDN U19984 ( .B(n16806), .A(n97), .Z(n16804) );
  XNOR U19985 ( .A(a[918]), .B(n16807), .Z(n97) );
  IV U19986 ( .A(n16805), .Z(n16807) );
  XNOR U19987 ( .A(b[918]), .B(n16805), .Z(n16806) );
  XOR U19988 ( .A(n16808), .B(n16809), .Z(n16805) );
  ANDN U19989 ( .B(n16810), .A(n98), .Z(n16808) );
  XNOR U19990 ( .A(a[917]), .B(n16811), .Z(n98) );
  IV U19991 ( .A(n16809), .Z(n16811) );
  XNOR U19992 ( .A(b[917]), .B(n16809), .Z(n16810) );
  XOR U19993 ( .A(n16812), .B(n16813), .Z(n16809) );
  ANDN U19994 ( .B(n16814), .A(n99), .Z(n16812) );
  XNOR U19995 ( .A(a[916]), .B(n16815), .Z(n99) );
  IV U19996 ( .A(n16813), .Z(n16815) );
  XNOR U19997 ( .A(b[916]), .B(n16813), .Z(n16814) );
  XOR U19998 ( .A(n16816), .B(n16817), .Z(n16813) );
  ANDN U19999 ( .B(n16818), .A(n100), .Z(n16816) );
  XNOR U20000 ( .A(a[915]), .B(n16819), .Z(n100) );
  IV U20001 ( .A(n16817), .Z(n16819) );
  XNOR U20002 ( .A(b[915]), .B(n16817), .Z(n16818) );
  XOR U20003 ( .A(n16820), .B(n16821), .Z(n16817) );
  ANDN U20004 ( .B(n16822), .A(n101), .Z(n16820) );
  XNOR U20005 ( .A(a[914]), .B(n16823), .Z(n101) );
  IV U20006 ( .A(n16821), .Z(n16823) );
  XNOR U20007 ( .A(b[914]), .B(n16821), .Z(n16822) );
  XOR U20008 ( .A(n16824), .B(n16825), .Z(n16821) );
  ANDN U20009 ( .B(n16826), .A(n102), .Z(n16824) );
  XNOR U20010 ( .A(a[913]), .B(n16827), .Z(n102) );
  IV U20011 ( .A(n16825), .Z(n16827) );
  XNOR U20012 ( .A(b[913]), .B(n16825), .Z(n16826) );
  XOR U20013 ( .A(n16828), .B(n16829), .Z(n16825) );
  ANDN U20014 ( .B(n16830), .A(n103), .Z(n16828) );
  XNOR U20015 ( .A(a[912]), .B(n16831), .Z(n103) );
  IV U20016 ( .A(n16829), .Z(n16831) );
  XNOR U20017 ( .A(b[912]), .B(n16829), .Z(n16830) );
  XOR U20018 ( .A(n16832), .B(n16833), .Z(n16829) );
  ANDN U20019 ( .B(n16834), .A(n104), .Z(n16832) );
  XNOR U20020 ( .A(a[911]), .B(n16835), .Z(n104) );
  IV U20021 ( .A(n16833), .Z(n16835) );
  XNOR U20022 ( .A(b[911]), .B(n16833), .Z(n16834) );
  XOR U20023 ( .A(n16836), .B(n16837), .Z(n16833) );
  ANDN U20024 ( .B(n16838), .A(n105), .Z(n16836) );
  XNOR U20025 ( .A(a[910]), .B(n16839), .Z(n105) );
  IV U20026 ( .A(n16837), .Z(n16839) );
  XNOR U20027 ( .A(b[910]), .B(n16837), .Z(n16838) );
  XOR U20028 ( .A(n16840), .B(n16841), .Z(n16837) );
  ANDN U20029 ( .B(n16842), .A(n107), .Z(n16840) );
  XNOR U20030 ( .A(a[909]), .B(n16843), .Z(n107) );
  IV U20031 ( .A(n16841), .Z(n16843) );
  XNOR U20032 ( .A(b[909]), .B(n16841), .Z(n16842) );
  XOR U20033 ( .A(n16844), .B(n16845), .Z(n16841) );
  ANDN U20034 ( .B(n16846), .A(n108), .Z(n16844) );
  XNOR U20035 ( .A(a[908]), .B(n16847), .Z(n108) );
  IV U20036 ( .A(n16845), .Z(n16847) );
  XNOR U20037 ( .A(b[908]), .B(n16845), .Z(n16846) );
  XOR U20038 ( .A(n16848), .B(n16849), .Z(n16845) );
  ANDN U20039 ( .B(n16850), .A(n109), .Z(n16848) );
  XNOR U20040 ( .A(a[907]), .B(n16851), .Z(n109) );
  IV U20041 ( .A(n16849), .Z(n16851) );
  XNOR U20042 ( .A(b[907]), .B(n16849), .Z(n16850) );
  XOR U20043 ( .A(n16852), .B(n16853), .Z(n16849) );
  ANDN U20044 ( .B(n16854), .A(n110), .Z(n16852) );
  XNOR U20045 ( .A(a[906]), .B(n16855), .Z(n110) );
  IV U20046 ( .A(n16853), .Z(n16855) );
  XNOR U20047 ( .A(b[906]), .B(n16853), .Z(n16854) );
  XOR U20048 ( .A(n16856), .B(n16857), .Z(n16853) );
  ANDN U20049 ( .B(n16858), .A(n111), .Z(n16856) );
  XNOR U20050 ( .A(a[905]), .B(n16859), .Z(n111) );
  IV U20051 ( .A(n16857), .Z(n16859) );
  XNOR U20052 ( .A(b[905]), .B(n16857), .Z(n16858) );
  XOR U20053 ( .A(n16860), .B(n16861), .Z(n16857) );
  ANDN U20054 ( .B(n16862), .A(n112), .Z(n16860) );
  XNOR U20055 ( .A(a[904]), .B(n16863), .Z(n112) );
  IV U20056 ( .A(n16861), .Z(n16863) );
  XNOR U20057 ( .A(b[904]), .B(n16861), .Z(n16862) );
  XOR U20058 ( .A(n16864), .B(n16865), .Z(n16861) );
  ANDN U20059 ( .B(n16866), .A(n113), .Z(n16864) );
  XNOR U20060 ( .A(a[903]), .B(n16867), .Z(n113) );
  IV U20061 ( .A(n16865), .Z(n16867) );
  XNOR U20062 ( .A(b[903]), .B(n16865), .Z(n16866) );
  XOR U20063 ( .A(n16868), .B(n16869), .Z(n16865) );
  ANDN U20064 ( .B(n16870), .A(n114), .Z(n16868) );
  XNOR U20065 ( .A(a[902]), .B(n16871), .Z(n114) );
  IV U20066 ( .A(n16869), .Z(n16871) );
  XNOR U20067 ( .A(b[902]), .B(n16869), .Z(n16870) );
  XOR U20068 ( .A(n16872), .B(n16873), .Z(n16869) );
  ANDN U20069 ( .B(n16874), .A(n115), .Z(n16872) );
  XNOR U20070 ( .A(a[901]), .B(n16875), .Z(n115) );
  IV U20071 ( .A(n16873), .Z(n16875) );
  XNOR U20072 ( .A(b[901]), .B(n16873), .Z(n16874) );
  XOR U20073 ( .A(n16876), .B(n16877), .Z(n16873) );
  ANDN U20074 ( .B(n16878), .A(n116), .Z(n16876) );
  XNOR U20075 ( .A(a[900]), .B(n16879), .Z(n116) );
  IV U20076 ( .A(n16877), .Z(n16879) );
  XNOR U20077 ( .A(b[900]), .B(n16877), .Z(n16878) );
  XOR U20078 ( .A(n16880), .B(n16881), .Z(n16877) );
  ANDN U20079 ( .B(n16882), .A(n119), .Z(n16880) );
  XNOR U20080 ( .A(a[899]), .B(n16883), .Z(n119) );
  IV U20081 ( .A(n16881), .Z(n16883) );
  XNOR U20082 ( .A(b[899]), .B(n16881), .Z(n16882) );
  XOR U20083 ( .A(n16884), .B(n16885), .Z(n16881) );
  ANDN U20084 ( .B(n16886), .A(n120), .Z(n16884) );
  XNOR U20085 ( .A(a[898]), .B(n16887), .Z(n120) );
  IV U20086 ( .A(n16885), .Z(n16887) );
  XNOR U20087 ( .A(b[898]), .B(n16885), .Z(n16886) );
  XOR U20088 ( .A(n16888), .B(n16889), .Z(n16885) );
  ANDN U20089 ( .B(n16890), .A(n121), .Z(n16888) );
  XNOR U20090 ( .A(a[897]), .B(n16891), .Z(n121) );
  IV U20091 ( .A(n16889), .Z(n16891) );
  XNOR U20092 ( .A(b[897]), .B(n16889), .Z(n16890) );
  XOR U20093 ( .A(n16892), .B(n16893), .Z(n16889) );
  ANDN U20094 ( .B(n16894), .A(n122), .Z(n16892) );
  XNOR U20095 ( .A(a[896]), .B(n16895), .Z(n122) );
  IV U20096 ( .A(n16893), .Z(n16895) );
  XNOR U20097 ( .A(b[896]), .B(n16893), .Z(n16894) );
  XOR U20098 ( .A(n16896), .B(n16897), .Z(n16893) );
  ANDN U20099 ( .B(n16898), .A(n123), .Z(n16896) );
  XNOR U20100 ( .A(a[895]), .B(n16899), .Z(n123) );
  IV U20101 ( .A(n16897), .Z(n16899) );
  XNOR U20102 ( .A(b[895]), .B(n16897), .Z(n16898) );
  XOR U20103 ( .A(n16900), .B(n16901), .Z(n16897) );
  ANDN U20104 ( .B(n16902), .A(n124), .Z(n16900) );
  XNOR U20105 ( .A(a[894]), .B(n16903), .Z(n124) );
  IV U20106 ( .A(n16901), .Z(n16903) );
  XNOR U20107 ( .A(b[894]), .B(n16901), .Z(n16902) );
  XOR U20108 ( .A(n16904), .B(n16905), .Z(n16901) );
  ANDN U20109 ( .B(n16906), .A(n125), .Z(n16904) );
  XNOR U20110 ( .A(a[893]), .B(n16907), .Z(n125) );
  IV U20111 ( .A(n16905), .Z(n16907) );
  XNOR U20112 ( .A(b[893]), .B(n16905), .Z(n16906) );
  XOR U20113 ( .A(n16908), .B(n16909), .Z(n16905) );
  ANDN U20114 ( .B(n16910), .A(n126), .Z(n16908) );
  XNOR U20115 ( .A(a[892]), .B(n16911), .Z(n126) );
  IV U20116 ( .A(n16909), .Z(n16911) );
  XNOR U20117 ( .A(b[892]), .B(n16909), .Z(n16910) );
  XOR U20118 ( .A(n16912), .B(n16913), .Z(n16909) );
  ANDN U20119 ( .B(n16914), .A(n127), .Z(n16912) );
  XNOR U20120 ( .A(a[891]), .B(n16915), .Z(n127) );
  IV U20121 ( .A(n16913), .Z(n16915) );
  XNOR U20122 ( .A(b[891]), .B(n16913), .Z(n16914) );
  XOR U20123 ( .A(n16916), .B(n16917), .Z(n16913) );
  ANDN U20124 ( .B(n16918), .A(n128), .Z(n16916) );
  XNOR U20125 ( .A(a[890]), .B(n16919), .Z(n128) );
  IV U20126 ( .A(n16917), .Z(n16919) );
  XNOR U20127 ( .A(b[890]), .B(n16917), .Z(n16918) );
  XOR U20128 ( .A(n16920), .B(n16921), .Z(n16917) );
  ANDN U20129 ( .B(n16922), .A(n130), .Z(n16920) );
  XNOR U20130 ( .A(a[889]), .B(n16923), .Z(n130) );
  IV U20131 ( .A(n16921), .Z(n16923) );
  XNOR U20132 ( .A(b[889]), .B(n16921), .Z(n16922) );
  XOR U20133 ( .A(n16924), .B(n16925), .Z(n16921) );
  ANDN U20134 ( .B(n16926), .A(n131), .Z(n16924) );
  XNOR U20135 ( .A(a[888]), .B(n16927), .Z(n131) );
  IV U20136 ( .A(n16925), .Z(n16927) );
  XNOR U20137 ( .A(b[888]), .B(n16925), .Z(n16926) );
  XOR U20138 ( .A(n16928), .B(n16929), .Z(n16925) );
  ANDN U20139 ( .B(n16930), .A(n132), .Z(n16928) );
  XNOR U20140 ( .A(a[887]), .B(n16931), .Z(n132) );
  IV U20141 ( .A(n16929), .Z(n16931) );
  XNOR U20142 ( .A(b[887]), .B(n16929), .Z(n16930) );
  XOR U20143 ( .A(n16932), .B(n16933), .Z(n16929) );
  ANDN U20144 ( .B(n16934), .A(n133), .Z(n16932) );
  XNOR U20145 ( .A(a[886]), .B(n16935), .Z(n133) );
  IV U20146 ( .A(n16933), .Z(n16935) );
  XNOR U20147 ( .A(b[886]), .B(n16933), .Z(n16934) );
  XOR U20148 ( .A(n16936), .B(n16937), .Z(n16933) );
  ANDN U20149 ( .B(n16938), .A(n134), .Z(n16936) );
  XNOR U20150 ( .A(a[885]), .B(n16939), .Z(n134) );
  IV U20151 ( .A(n16937), .Z(n16939) );
  XNOR U20152 ( .A(b[885]), .B(n16937), .Z(n16938) );
  XOR U20153 ( .A(n16940), .B(n16941), .Z(n16937) );
  ANDN U20154 ( .B(n16942), .A(n135), .Z(n16940) );
  XNOR U20155 ( .A(a[884]), .B(n16943), .Z(n135) );
  IV U20156 ( .A(n16941), .Z(n16943) );
  XNOR U20157 ( .A(b[884]), .B(n16941), .Z(n16942) );
  XOR U20158 ( .A(n16944), .B(n16945), .Z(n16941) );
  ANDN U20159 ( .B(n16946), .A(n136), .Z(n16944) );
  XNOR U20160 ( .A(a[883]), .B(n16947), .Z(n136) );
  IV U20161 ( .A(n16945), .Z(n16947) );
  XNOR U20162 ( .A(b[883]), .B(n16945), .Z(n16946) );
  XOR U20163 ( .A(n16948), .B(n16949), .Z(n16945) );
  ANDN U20164 ( .B(n16950), .A(n137), .Z(n16948) );
  XNOR U20165 ( .A(a[882]), .B(n16951), .Z(n137) );
  IV U20166 ( .A(n16949), .Z(n16951) );
  XNOR U20167 ( .A(b[882]), .B(n16949), .Z(n16950) );
  XOR U20168 ( .A(n16952), .B(n16953), .Z(n16949) );
  ANDN U20169 ( .B(n16954), .A(n138), .Z(n16952) );
  XNOR U20170 ( .A(a[881]), .B(n16955), .Z(n138) );
  IV U20171 ( .A(n16953), .Z(n16955) );
  XNOR U20172 ( .A(b[881]), .B(n16953), .Z(n16954) );
  XOR U20173 ( .A(n16956), .B(n16957), .Z(n16953) );
  ANDN U20174 ( .B(n16958), .A(n139), .Z(n16956) );
  XNOR U20175 ( .A(a[880]), .B(n16959), .Z(n139) );
  IV U20176 ( .A(n16957), .Z(n16959) );
  XNOR U20177 ( .A(b[880]), .B(n16957), .Z(n16958) );
  XOR U20178 ( .A(n16960), .B(n16961), .Z(n16957) );
  ANDN U20179 ( .B(n16962), .A(n141), .Z(n16960) );
  XNOR U20180 ( .A(a[879]), .B(n16963), .Z(n141) );
  IV U20181 ( .A(n16961), .Z(n16963) );
  XNOR U20182 ( .A(b[879]), .B(n16961), .Z(n16962) );
  XOR U20183 ( .A(n16964), .B(n16965), .Z(n16961) );
  ANDN U20184 ( .B(n16966), .A(n142), .Z(n16964) );
  XNOR U20185 ( .A(a[878]), .B(n16967), .Z(n142) );
  IV U20186 ( .A(n16965), .Z(n16967) );
  XNOR U20187 ( .A(b[878]), .B(n16965), .Z(n16966) );
  XOR U20188 ( .A(n16968), .B(n16969), .Z(n16965) );
  ANDN U20189 ( .B(n16970), .A(n143), .Z(n16968) );
  XNOR U20190 ( .A(a[877]), .B(n16971), .Z(n143) );
  IV U20191 ( .A(n16969), .Z(n16971) );
  XNOR U20192 ( .A(b[877]), .B(n16969), .Z(n16970) );
  XOR U20193 ( .A(n16972), .B(n16973), .Z(n16969) );
  ANDN U20194 ( .B(n16974), .A(n144), .Z(n16972) );
  XNOR U20195 ( .A(a[876]), .B(n16975), .Z(n144) );
  IV U20196 ( .A(n16973), .Z(n16975) );
  XNOR U20197 ( .A(b[876]), .B(n16973), .Z(n16974) );
  XOR U20198 ( .A(n16976), .B(n16977), .Z(n16973) );
  ANDN U20199 ( .B(n16978), .A(n145), .Z(n16976) );
  XNOR U20200 ( .A(a[875]), .B(n16979), .Z(n145) );
  IV U20201 ( .A(n16977), .Z(n16979) );
  XNOR U20202 ( .A(b[875]), .B(n16977), .Z(n16978) );
  XOR U20203 ( .A(n16980), .B(n16981), .Z(n16977) );
  ANDN U20204 ( .B(n16982), .A(n146), .Z(n16980) );
  XNOR U20205 ( .A(a[874]), .B(n16983), .Z(n146) );
  IV U20206 ( .A(n16981), .Z(n16983) );
  XNOR U20207 ( .A(b[874]), .B(n16981), .Z(n16982) );
  XOR U20208 ( .A(n16984), .B(n16985), .Z(n16981) );
  ANDN U20209 ( .B(n16986), .A(n147), .Z(n16984) );
  XNOR U20210 ( .A(a[873]), .B(n16987), .Z(n147) );
  IV U20211 ( .A(n16985), .Z(n16987) );
  XNOR U20212 ( .A(b[873]), .B(n16985), .Z(n16986) );
  XOR U20213 ( .A(n16988), .B(n16989), .Z(n16985) );
  ANDN U20214 ( .B(n16990), .A(n148), .Z(n16988) );
  XNOR U20215 ( .A(a[872]), .B(n16991), .Z(n148) );
  IV U20216 ( .A(n16989), .Z(n16991) );
  XNOR U20217 ( .A(b[872]), .B(n16989), .Z(n16990) );
  XOR U20218 ( .A(n16992), .B(n16993), .Z(n16989) );
  ANDN U20219 ( .B(n16994), .A(n149), .Z(n16992) );
  XNOR U20220 ( .A(a[871]), .B(n16995), .Z(n149) );
  IV U20221 ( .A(n16993), .Z(n16995) );
  XNOR U20222 ( .A(b[871]), .B(n16993), .Z(n16994) );
  XOR U20223 ( .A(n16996), .B(n16997), .Z(n16993) );
  ANDN U20224 ( .B(n16998), .A(n150), .Z(n16996) );
  XNOR U20225 ( .A(a[870]), .B(n16999), .Z(n150) );
  IV U20226 ( .A(n16997), .Z(n16999) );
  XNOR U20227 ( .A(b[870]), .B(n16997), .Z(n16998) );
  XOR U20228 ( .A(n17000), .B(n17001), .Z(n16997) );
  ANDN U20229 ( .B(n17002), .A(n152), .Z(n17000) );
  XNOR U20230 ( .A(a[869]), .B(n17003), .Z(n152) );
  IV U20231 ( .A(n17001), .Z(n17003) );
  XNOR U20232 ( .A(b[869]), .B(n17001), .Z(n17002) );
  XOR U20233 ( .A(n17004), .B(n17005), .Z(n17001) );
  ANDN U20234 ( .B(n17006), .A(n153), .Z(n17004) );
  XNOR U20235 ( .A(a[868]), .B(n17007), .Z(n153) );
  IV U20236 ( .A(n17005), .Z(n17007) );
  XNOR U20237 ( .A(b[868]), .B(n17005), .Z(n17006) );
  XOR U20238 ( .A(n17008), .B(n17009), .Z(n17005) );
  ANDN U20239 ( .B(n17010), .A(n154), .Z(n17008) );
  XNOR U20240 ( .A(a[867]), .B(n17011), .Z(n154) );
  IV U20241 ( .A(n17009), .Z(n17011) );
  XNOR U20242 ( .A(b[867]), .B(n17009), .Z(n17010) );
  XOR U20243 ( .A(n17012), .B(n17013), .Z(n17009) );
  ANDN U20244 ( .B(n17014), .A(n155), .Z(n17012) );
  XNOR U20245 ( .A(a[866]), .B(n17015), .Z(n155) );
  IV U20246 ( .A(n17013), .Z(n17015) );
  XNOR U20247 ( .A(b[866]), .B(n17013), .Z(n17014) );
  XOR U20248 ( .A(n17016), .B(n17017), .Z(n17013) );
  ANDN U20249 ( .B(n17018), .A(n156), .Z(n17016) );
  XNOR U20250 ( .A(a[865]), .B(n17019), .Z(n156) );
  IV U20251 ( .A(n17017), .Z(n17019) );
  XNOR U20252 ( .A(b[865]), .B(n17017), .Z(n17018) );
  XOR U20253 ( .A(n17020), .B(n17021), .Z(n17017) );
  ANDN U20254 ( .B(n17022), .A(n157), .Z(n17020) );
  XNOR U20255 ( .A(a[864]), .B(n17023), .Z(n157) );
  IV U20256 ( .A(n17021), .Z(n17023) );
  XNOR U20257 ( .A(b[864]), .B(n17021), .Z(n17022) );
  XOR U20258 ( .A(n17024), .B(n17025), .Z(n17021) );
  ANDN U20259 ( .B(n17026), .A(n158), .Z(n17024) );
  XNOR U20260 ( .A(a[863]), .B(n17027), .Z(n158) );
  IV U20261 ( .A(n17025), .Z(n17027) );
  XNOR U20262 ( .A(b[863]), .B(n17025), .Z(n17026) );
  XOR U20263 ( .A(n17028), .B(n17029), .Z(n17025) );
  ANDN U20264 ( .B(n17030), .A(n159), .Z(n17028) );
  XNOR U20265 ( .A(a[862]), .B(n17031), .Z(n159) );
  IV U20266 ( .A(n17029), .Z(n17031) );
  XNOR U20267 ( .A(b[862]), .B(n17029), .Z(n17030) );
  XOR U20268 ( .A(n17032), .B(n17033), .Z(n17029) );
  ANDN U20269 ( .B(n17034), .A(n160), .Z(n17032) );
  XNOR U20270 ( .A(a[861]), .B(n17035), .Z(n160) );
  IV U20271 ( .A(n17033), .Z(n17035) );
  XNOR U20272 ( .A(b[861]), .B(n17033), .Z(n17034) );
  XOR U20273 ( .A(n17036), .B(n17037), .Z(n17033) );
  ANDN U20274 ( .B(n17038), .A(n161), .Z(n17036) );
  XNOR U20275 ( .A(a[860]), .B(n17039), .Z(n161) );
  IV U20276 ( .A(n17037), .Z(n17039) );
  XNOR U20277 ( .A(b[860]), .B(n17037), .Z(n17038) );
  XOR U20278 ( .A(n17040), .B(n17041), .Z(n17037) );
  ANDN U20279 ( .B(n17042), .A(n163), .Z(n17040) );
  XNOR U20280 ( .A(a[859]), .B(n17043), .Z(n163) );
  IV U20281 ( .A(n17041), .Z(n17043) );
  XNOR U20282 ( .A(b[859]), .B(n17041), .Z(n17042) );
  XOR U20283 ( .A(n17044), .B(n17045), .Z(n17041) );
  ANDN U20284 ( .B(n17046), .A(n164), .Z(n17044) );
  XNOR U20285 ( .A(a[858]), .B(n17047), .Z(n164) );
  IV U20286 ( .A(n17045), .Z(n17047) );
  XNOR U20287 ( .A(b[858]), .B(n17045), .Z(n17046) );
  XOR U20288 ( .A(n17048), .B(n17049), .Z(n17045) );
  ANDN U20289 ( .B(n17050), .A(n165), .Z(n17048) );
  XNOR U20290 ( .A(a[857]), .B(n17051), .Z(n165) );
  IV U20291 ( .A(n17049), .Z(n17051) );
  XNOR U20292 ( .A(b[857]), .B(n17049), .Z(n17050) );
  XOR U20293 ( .A(n17052), .B(n17053), .Z(n17049) );
  ANDN U20294 ( .B(n17054), .A(n166), .Z(n17052) );
  XNOR U20295 ( .A(a[856]), .B(n17055), .Z(n166) );
  IV U20296 ( .A(n17053), .Z(n17055) );
  XNOR U20297 ( .A(b[856]), .B(n17053), .Z(n17054) );
  XOR U20298 ( .A(n17056), .B(n17057), .Z(n17053) );
  ANDN U20299 ( .B(n17058), .A(n167), .Z(n17056) );
  XNOR U20300 ( .A(a[855]), .B(n17059), .Z(n167) );
  IV U20301 ( .A(n17057), .Z(n17059) );
  XNOR U20302 ( .A(b[855]), .B(n17057), .Z(n17058) );
  XOR U20303 ( .A(n17060), .B(n17061), .Z(n17057) );
  ANDN U20304 ( .B(n17062), .A(n168), .Z(n17060) );
  XNOR U20305 ( .A(a[854]), .B(n17063), .Z(n168) );
  IV U20306 ( .A(n17061), .Z(n17063) );
  XNOR U20307 ( .A(b[854]), .B(n17061), .Z(n17062) );
  XOR U20308 ( .A(n17064), .B(n17065), .Z(n17061) );
  ANDN U20309 ( .B(n17066), .A(n169), .Z(n17064) );
  XNOR U20310 ( .A(a[853]), .B(n17067), .Z(n169) );
  IV U20311 ( .A(n17065), .Z(n17067) );
  XNOR U20312 ( .A(b[853]), .B(n17065), .Z(n17066) );
  XOR U20313 ( .A(n17068), .B(n17069), .Z(n17065) );
  ANDN U20314 ( .B(n17070), .A(n170), .Z(n17068) );
  XNOR U20315 ( .A(a[852]), .B(n17071), .Z(n170) );
  IV U20316 ( .A(n17069), .Z(n17071) );
  XNOR U20317 ( .A(b[852]), .B(n17069), .Z(n17070) );
  XOR U20318 ( .A(n17072), .B(n17073), .Z(n17069) );
  ANDN U20319 ( .B(n17074), .A(n171), .Z(n17072) );
  XNOR U20320 ( .A(a[851]), .B(n17075), .Z(n171) );
  IV U20321 ( .A(n17073), .Z(n17075) );
  XNOR U20322 ( .A(b[851]), .B(n17073), .Z(n17074) );
  XOR U20323 ( .A(n17076), .B(n17077), .Z(n17073) );
  ANDN U20324 ( .B(n17078), .A(n172), .Z(n17076) );
  XNOR U20325 ( .A(a[850]), .B(n17079), .Z(n172) );
  IV U20326 ( .A(n17077), .Z(n17079) );
  XNOR U20327 ( .A(b[850]), .B(n17077), .Z(n17078) );
  XOR U20328 ( .A(n17080), .B(n17081), .Z(n17077) );
  ANDN U20329 ( .B(n17082), .A(n174), .Z(n17080) );
  XNOR U20330 ( .A(a[849]), .B(n17083), .Z(n174) );
  IV U20331 ( .A(n17081), .Z(n17083) );
  XNOR U20332 ( .A(b[849]), .B(n17081), .Z(n17082) );
  XOR U20333 ( .A(n17084), .B(n17085), .Z(n17081) );
  ANDN U20334 ( .B(n17086), .A(n175), .Z(n17084) );
  XNOR U20335 ( .A(a[848]), .B(n17087), .Z(n175) );
  IV U20336 ( .A(n17085), .Z(n17087) );
  XNOR U20337 ( .A(b[848]), .B(n17085), .Z(n17086) );
  XOR U20338 ( .A(n17088), .B(n17089), .Z(n17085) );
  ANDN U20339 ( .B(n17090), .A(n176), .Z(n17088) );
  XNOR U20340 ( .A(a[847]), .B(n17091), .Z(n176) );
  IV U20341 ( .A(n17089), .Z(n17091) );
  XNOR U20342 ( .A(b[847]), .B(n17089), .Z(n17090) );
  XOR U20343 ( .A(n17092), .B(n17093), .Z(n17089) );
  ANDN U20344 ( .B(n17094), .A(n177), .Z(n17092) );
  XNOR U20345 ( .A(a[846]), .B(n17095), .Z(n177) );
  IV U20346 ( .A(n17093), .Z(n17095) );
  XNOR U20347 ( .A(b[846]), .B(n17093), .Z(n17094) );
  XOR U20348 ( .A(n17096), .B(n17097), .Z(n17093) );
  ANDN U20349 ( .B(n17098), .A(n178), .Z(n17096) );
  XNOR U20350 ( .A(a[845]), .B(n17099), .Z(n178) );
  IV U20351 ( .A(n17097), .Z(n17099) );
  XNOR U20352 ( .A(b[845]), .B(n17097), .Z(n17098) );
  XOR U20353 ( .A(n17100), .B(n17101), .Z(n17097) );
  ANDN U20354 ( .B(n17102), .A(n179), .Z(n17100) );
  XNOR U20355 ( .A(a[844]), .B(n17103), .Z(n179) );
  IV U20356 ( .A(n17101), .Z(n17103) );
  XNOR U20357 ( .A(b[844]), .B(n17101), .Z(n17102) );
  XOR U20358 ( .A(n17104), .B(n17105), .Z(n17101) );
  ANDN U20359 ( .B(n17106), .A(n180), .Z(n17104) );
  XNOR U20360 ( .A(a[843]), .B(n17107), .Z(n180) );
  IV U20361 ( .A(n17105), .Z(n17107) );
  XNOR U20362 ( .A(b[843]), .B(n17105), .Z(n17106) );
  XOR U20363 ( .A(n17108), .B(n17109), .Z(n17105) );
  ANDN U20364 ( .B(n17110), .A(n181), .Z(n17108) );
  XNOR U20365 ( .A(a[842]), .B(n17111), .Z(n181) );
  IV U20366 ( .A(n17109), .Z(n17111) );
  XNOR U20367 ( .A(b[842]), .B(n17109), .Z(n17110) );
  XOR U20368 ( .A(n17112), .B(n17113), .Z(n17109) );
  ANDN U20369 ( .B(n17114), .A(n182), .Z(n17112) );
  XNOR U20370 ( .A(a[841]), .B(n17115), .Z(n182) );
  IV U20371 ( .A(n17113), .Z(n17115) );
  XNOR U20372 ( .A(b[841]), .B(n17113), .Z(n17114) );
  XOR U20373 ( .A(n17116), .B(n17117), .Z(n17113) );
  ANDN U20374 ( .B(n17118), .A(n183), .Z(n17116) );
  XNOR U20375 ( .A(a[840]), .B(n17119), .Z(n183) );
  IV U20376 ( .A(n17117), .Z(n17119) );
  XNOR U20377 ( .A(b[840]), .B(n17117), .Z(n17118) );
  XOR U20378 ( .A(n17120), .B(n17121), .Z(n17117) );
  ANDN U20379 ( .B(n17122), .A(n185), .Z(n17120) );
  XNOR U20380 ( .A(a[839]), .B(n17123), .Z(n185) );
  IV U20381 ( .A(n17121), .Z(n17123) );
  XNOR U20382 ( .A(b[839]), .B(n17121), .Z(n17122) );
  XOR U20383 ( .A(n17124), .B(n17125), .Z(n17121) );
  ANDN U20384 ( .B(n17126), .A(n186), .Z(n17124) );
  XNOR U20385 ( .A(a[838]), .B(n17127), .Z(n186) );
  IV U20386 ( .A(n17125), .Z(n17127) );
  XNOR U20387 ( .A(b[838]), .B(n17125), .Z(n17126) );
  XOR U20388 ( .A(n17128), .B(n17129), .Z(n17125) );
  ANDN U20389 ( .B(n17130), .A(n187), .Z(n17128) );
  XNOR U20390 ( .A(a[837]), .B(n17131), .Z(n187) );
  IV U20391 ( .A(n17129), .Z(n17131) );
  XNOR U20392 ( .A(b[837]), .B(n17129), .Z(n17130) );
  XOR U20393 ( .A(n17132), .B(n17133), .Z(n17129) );
  ANDN U20394 ( .B(n17134), .A(n188), .Z(n17132) );
  XNOR U20395 ( .A(a[836]), .B(n17135), .Z(n188) );
  IV U20396 ( .A(n17133), .Z(n17135) );
  XNOR U20397 ( .A(b[836]), .B(n17133), .Z(n17134) );
  XOR U20398 ( .A(n17136), .B(n17137), .Z(n17133) );
  ANDN U20399 ( .B(n17138), .A(n189), .Z(n17136) );
  XNOR U20400 ( .A(a[835]), .B(n17139), .Z(n189) );
  IV U20401 ( .A(n17137), .Z(n17139) );
  XNOR U20402 ( .A(b[835]), .B(n17137), .Z(n17138) );
  XOR U20403 ( .A(n17140), .B(n17141), .Z(n17137) );
  ANDN U20404 ( .B(n17142), .A(n190), .Z(n17140) );
  XNOR U20405 ( .A(a[834]), .B(n17143), .Z(n190) );
  IV U20406 ( .A(n17141), .Z(n17143) );
  XNOR U20407 ( .A(b[834]), .B(n17141), .Z(n17142) );
  XOR U20408 ( .A(n17144), .B(n17145), .Z(n17141) );
  ANDN U20409 ( .B(n17146), .A(n191), .Z(n17144) );
  XNOR U20410 ( .A(a[833]), .B(n17147), .Z(n191) );
  IV U20411 ( .A(n17145), .Z(n17147) );
  XNOR U20412 ( .A(b[833]), .B(n17145), .Z(n17146) );
  XOR U20413 ( .A(n17148), .B(n17149), .Z(n17145) );
  ANDN U20414 ( .B(n17150), .A(n192), .Z(n17148) );
  XNOR U20415 ( .A(a[832]), .B(n17151), .Z(n192) );
  IV U20416 ( .A(n17149), .Z(n17151) );
  XNOR U20417 ( .A(b[832]), .B(n17149), .Z(n17150) );
  XOR U20418 ( .A(n17152), .B(n17153), .Z(n17149) );
  ANDN U20419 ( .B(n17154), .A(n193), .Z(n17152) );
  XNOR U20420 ( .A(a[831]), .B(n17155), .Z(n193) );
  IV U20421 ( .A(n17153), .Z(n17155) );
  XNOR U20422 ( .A(b[831]), .B(n17153), .Z(n17154) );
  XOR U20423 ( .A(n17156), .B(n17157), .Z(n17153) );
  ANDN U20424 ( .B(n17158), .A(n194), .Z(n17156) );
  XNOR U20425 ( .A(a[830]), .B(n17159), .Z(n194) );
  IV U20426 ( .A(n17157), .Z(n17159) );
  XNOR U20427 ( .A(b[830]), .B(n17157), .Z(n17158) );
  XOR U20428 ( .A(n17160), .B(n17161), .Z(n17157) );
  ANDN U20429 ( .B(n17162), .A(n196), .Z(n17160) );
  XNOR U20430 ( .A(a[829]), .B(n17163), .Z(n196) );
  IV U20431 ( .A(n17161), .Z(n17163) );
  XNOR U20432 ( .A(b[829]), .B(n17161), .Z(n17162) );
  XOR U20433 ( .A(n17164), .B(n17165), .Z(n17161) );
  ANDN U20434 ( .B(n17166), .A(n197), .Z(n17164) );
  XNOR U20435 ( .A(a[828]), .B(n17167), .Z(n197) );
  IV U20436 ( .A(n17165), .Z(n17167) );
  XNOR U20437 ( .A(b[828]), .B(n17165), .Z(n17166) );
  XOR U20438 ( .A(n17168), .B(n17169), .Z(n17165) );
  ANDN U20439 ( .B(n17170), .A(n198), .Z(n17168) );
  XNOR U20440 ( .A(a[827]), .B(n17171), .Z(n198) );
  IV U20441 ( .A(n17169), .Z(n17171) );
  XNOR U20442 ( .A(b[827]), .B(n17169), .Z(n17170) );
  XOR U20443 ( .A(n17172), .B(n17173), .Z(n17169) );
  ANDN U20444 ( .B(n17174), .A(n199), .Z(n17172) );
  XNOR U20445 ( .A(a[826]), .B(n17175), .Z(n199) );
  IV U20446 ( .A(n17173), .Z(n17175) );
  XNOR U20447 ( .A(b[826]), .B(n17173), .Z(n17174) );
  XOR U20448 ( .A(n17176), .B(n17177), .Z(n17173) );
  ANDN U20449 ( .B(n17178), .A(n200), .Z(n17176) );
  XNOR U20450 ( .A(a[825]), .B(n17179), .Z(n200) );
  IV U20451 ( .A(n17177), .Z(n17179) );
  XNOR U20452 ( .A(b[825]), .B(n17177), .Z(n17178) );
  XOR U20453 ( .A(n17180), .B(n17181), .Z(n17177) );
  ANDN U20454 ( .B(n17182), .A(n201), .Z(n17180) );
  XNOR U20455 ( .A(a[824]), .B(n17183), .Z(n201) );
  IV U20456 ( .A(n17181), .Z(n17183) );
  XNOR U20457 ( .A(b[824]), .B(n17181), .Z(n17182) );
  XOR U20458 ( .A(n17184), .B(n17185), .Z(n17181) );
  ANDN U20459 ( .B(n17186), .A(n202), .Z(n17184) );
  XNOR U20460 ( .A(a[823]), .B(n17187), .Z(n202) );
  IV U20461 ( .A(n17185), .Z(n17187) );
  XNOR U20462 ( .A(b[823]), .B(n17185), .Z(n17186) );
  XOR U20463 ( .A(n17188), .B(n17189), .Z(n17185) );
  ANDN U20464 ( .B(n17190), .A(n203), .Z(n17188) );
  XNOR U20465 ( .A(a[822]), .B(n17191), .Z(n203) );
  IV U20466 ( .A(n17189), .Z(n17191) );
  XNOR U20467 ( .A(b[822]), .B(n17189), .Z(n17190) );
  XOR U20468 ( .A(n17192), .B(n17193), .Z(n17189) );
  ANDN U20469 ( .B(n17194), .A(n204), .Z(n17192) );
  XNOR U20470 ( .A(a[821]), .B(n17195), .Z(n204) );
  IV U20471 ( .A(n17193), .Z(n17195) );
  XNOR U20472 ( .A(b[821]), .B(n17193), .Z(n17194) );
  XOR U20473 ( .A(n17196), .B(n17197), .Z(n17193) );
  ANDN U20474 ( .B(n17198), .A(n205), .Z(n17196) );
  XNOR U20475 ( .A(a[820]), .B(n17199), .Z(n205) );
  IV U20476 ( .A(n17197), .Z(n17199) );
  XNOR U20477 ( .A(b[820]), .B(n17197), .Z(n17198) );
  XOR U20478 ( .A(n17200), .B(n17201), .Z(n17197) );
  ANDN U20479 ( .B(n17202), .A(n207), .Z(n17200) );
  XNOR U20480 ( .A(a[819]), .B(n17203), .Z(n207) );
  IV U20481 ( .A(n17201), .Z(n17203) );
  XNOR U20482 ( .A(b[819]), .B(n17201), .Z(n17202) );
  XOR U20483 ( .A(n17204), .B(n17205), .Z(n17201) );
  ANDN U20484 ( .B(n17206), .A(n208), .Z(n17204) );
  XNOR U20485 ( .A(a[818]), .B(n17207), .Z(n208) );
  IV U20486 ( .A(n17205), .Z(n17207) );
  XNOR U20487 ( .A(b[818]), .B(n17205), .Z(n17206) );
  XOR U20488 ( .A(n17208), .B(n17209), .Z(n17205) );
  ANDN U20489 ( .B(n17210), .A(n209), .Z(n17208) );
  XNOR U20490 ( .A(a[817]), .B(n17211), .Z(n209) );
  IV U20491 ( .A(n17209), .Z(n17211) );
  XNOR U20492 ( .A(b[817]), .B(n17209), .Z(n17210) );
  XOR U20493 ( .A(n17212), .B(n17213), .Z(n17209) );
  ANDN U20494 ( .B(n17214), .A(n210), .Z(n17212) );
  XNOR U20495 ( .A(a[816]), .B(n17215), .Z(n210) );
  IV U20496 ( .A(n17213), .Z(n17215) );
  XNOR U20497 ( .A(b[816]), .B(n17213), .Z(n17214) );
  XOR U20498 ( .A(n17216), .B(n17217), .Z(n17213) );
  ANDN U20499 ( .B(n17218), .A(n211), .Z(n17216) );
  XNOR U20500 ( .A(a[815]), .B(n17219), .Z(n211) );
  IV U20501 ( .A(n17217), .Z(n17219) );
  XNOR U20502 ( .A(b[815]), .B(n17217), .Z(n17218) );
  XOR U20503 ( .A(n17220), .B(n17221), .Z(n17217) );
  ANDN U20504 ( .B(n17222), .A(n212), .Z(n17220) );
  XNOR U20505 ( .A(a[814]), .B(n17223), .Z(n212) );
  IV U20506 ( .A(n17221), .Z(n17223) );
  XNOR U20507 ( .A(b[814]), .B(n17221), .Z(n17222) );
  XOR U20508 ( .A(n17224), .B(n17225), .Z(n17221) );
  ANDN U20509 ( .B(n17226), .A(n213), .Z(n17224) );
  XNOR U20510 ( .A(a[813]), .B(n17227), .Z(n213) );
  IV U20511 ( .A(n17225), .Z(n17227) );
  XNOR U20512 ( .A(b[813]), .B(n17225), .Z(n17226) );
  XOR U20513 ( .A(n17228), .B(n17229), .Z(n17225) );
  ANDN U20514 ( .B(n17230), .A(n214), .Z(n17228) );
  XNOR U20515 ( .A(a[812]), .B(n17231), .Z(n214) );
  IV U20516 ( .A(n17229), .Z(n17231) );
  XNOR U20517 ( .A(b[812]), .B(n17229), .Z(n17230) );
  XOR U20518 ( .A(n17232), .B(n17233), .Z(n17229) );
  ANDN U20519 ( .B(n17234), .A(n215), .Z(n17232) );
  XNOR U20520 ( .A(a[811]), .B(n17235), .Z(n215) );
  IV U20521 ( .A(n17233), .Z(n17235) );
  XNOR U20522 ( .A(b[811]), .B(n17233), .Z(n17234) );
  XOR U20523 ( .A(n17236), .B(n17237), .Z(n17233) );
  ANDN U20524 ( .B(n17238), .A(n216), .Z(n17236) );
  XNOR U20525 ( .A(a[810]), .B(n17239), .Z(n216) );
  IV U20526 ( .A(n17237), .Z(n17239) );
  XNOR U20527 ( .A(b[810]), .B(n17237), .Z(n17238) );
  XOR U20528 ( .A(n17240), .B(n17241), .Z(n17237) );
  ANDN U20529 ( .B(n17242), .A(n218), .Z(n17240) );
  XNOR U20530 ( .A(a[809]), .B(n17243), .Z(n218) );
  IV U20531 ( .A(n17241), .Z(n17243) );
  XNOR U20532 ( .A(b[809]), .B(n17241), .Z(n17242) );
  XOR U20533 ( .A(n17244), .B(n17245), .Z(n17241) );
  ANDN U20534 ( .B(n17246), .A(n219), .Z(n17244) );
  XNOR U20535 ( .A(a[808]), .B(n17247), .Z(n219) );
  IV U20536 ( .A(n17245), .Z(n17247) );
  XNOR U20537 ( .A(b[808]), .B(n17245), .Z(n17246) );
  XOR U20538 ( .A(n17248), .B(n17249), .Z(n17245) );
  ANDN U20539 ( .B(n17250), .A(n220), .Z(n17248) );
  XNOR U20540 ( .A(a[807]), .B(n17251), .Z(n220) );
  IV U20541 ( .A(n17249), .Z(n17251) );
  XNOR U20542 ( .A(b[807]), .B(n17249), .Z(n17250) );
  XOR U20543 ( .A(n17252), .B(n17253), .Z(n17249) );
  ANDN U20544 ( .B(n17254), .A(n221), .Z(n17252) );
  XNOR U20545 ( .A(a[806]), .B(n17255), .Z(n221) );
  IV U20546 ( .A(n17253), .Z(n17255) );
  XNOR U20547 ( .A(b[806]), .B(n17253), .Z(n17254) );
  XOR U20548 ( .A(n17256), .B(n17257), .Z(n17253) );
  ANDN U20549 ( .B(n17258), .A(n222), .Z(n17256) );
  XNOR U20550 ( .A(a[805]), .B(n17259), .Z(n222) );
  IV U20551 ( .A(n17257), .Z(n17259) );
  XNOR U20552 ( .A(b[805]), .B(n17257), .Z(n17258) );
  XOR U20553 ( .A(n17260), .B(n17261), .Z(n17257) );
  ANDN U20554 ( .B(n17262), .A(n223), .Z(n17260) );
  XNOR U20555 ( .A(a[804]), .B(n17263), .Z(n223) );
  IV U20556 ( .A(n17261), .Z(n17263) );
  XNOR U20557 ( .A(b[804]), .B(n17261), .Z(n17262) );
  XOR U20558 ( .A(n17264), .B(n17265), .Z(n17261) );
  ANDN U20559 ( .B(n17266), .A(n224), .Z(n17264) );
  XNOR U20560 ( .A(a[803]), .B(n17267), .Z(n224) );
  IV U20561 ( .A(n17265), .Z(n17267) );
  XNOR U20562 ( .A(b[803]), .B(n17265), .Z(n17266) );
  XOR U20563 ( .A(n17268), .B(n17269), .Z(n17265) );
  ANDN U20564 ( .B(n17270), .A(n225), .Z(n17268) );
  XNOR U20565 ( .A(a[802]), .B(n17271), .Z(n225) );
  IV U20566 ( .A(n17269), .Z(n17271) );
  XNOR U20567 ( .A(b[802]), .B(n17269), .Z(n17270) );
  XOR U20568 ( .A(n17272), .B(n17273), .Z(n17269) );
  ANDN U20569 ( .B(n17274), .A(n226), .Z(n17272) );
  XNOR U20570 ( .A(a[801]), .B(n17275), .Z(n226) );
  IV U20571 ( .A(n17273), .Z(n17275) );
  XNOR U20572 ( .A(b[801]), .B(n17273), .Z(n17274) );
  XOR U20573 ( .A(n17276), .B(n17277), .Z(n17273) );
  ANDN U20574 ( .B(n17278), .A(n227), .Z(n17276) );
  XNOR U20575 ( .A(a[800]), .B(n17279), .Z(n227) );
  IV U20576 ( .A(n17277), .Z(n17279) );
  XNOR U20577 ( .A(b[800]), .B(n17277), .Z(n17278) );
  XOR U20578 ( .A(n17280), .B(n17281), .Z(n17277) );
  ANDN U20579 ( .B(n17282), .A(n230), .Z(n17280) );
  XNOR U20580 ( .A(a[799]), .B(n17283), .Z(n230) );
  IV U20581 ( .A(n17281), .Z(n17283) );
  XNOR U20582 ( .A(b[799]), .B(n17281), .Z(n17282) );
  XOR U20583 ( .A(n17284), .B(n17285), .Z(n17281) );
  ANDN U20584 ( .B(n17286), .A(n231), .Z(n17284) );
  XNOR U20585 ( .A(a[798]), .B(n17287), .Z(n231) );
  IV U20586 ( .A(n17285), .Z(n17287) );
  XNOR U20587 ( .A(b[798]), .B(n17285), .Z(n17286) );
  XOR U20588 ( .A(n17288), .B(n17289), .Z(n17285) );
  ANDN U20589 ( .B(n17290), .A(n232), .Z(n17288) );
  XNOR U20590 ( .A(a[797]), .B(n17291), .Z(n232) );
  IV U20591 ( .A(n17289), .Z(n17291) );
  XNOR U20592 ( .A(b[797]), .B(n17289), .Z(n17290) );
  XOR U20593 ( .A(n17292), .B(n17293), .Z(n17289) );
  ANDN U20594 ( .B(n17294), .A(n233), .Z(n17292) );
  XNOR U20595 ( .A(a[796]), .B(n17295), .Z(n233) );
  IV U20596 ( .A(n17293), .Z(n17295) );
  XNOR U20597 ( .A(b[796]), .B(n17293), .Z(n17294) );
  XOR U20598 ( .A(n17296), .B(n17297), .Z(n17293) );
  ANDN U20599 ( .B(n17298), .A(n234), .Z(n17296) );
  XNOR U20600 ( .A(a[795]), .B(n17299), .Z(n234) );
  IV U20601 ( .A(n17297), .Z(n17299) );
  XNOR U20602 ( .A(b[795]), .B(n17297), .Z(n17298) );
  XOR U20603 ( .A(n17300), .B(n17301), .Z(n17297) );
  ANDN U20604 ( .B(n17302), .A(n235), .Z(n17300) );
  XNOR U20605 ( .A(a[794]), .B(n17303), .Z(n235) );
  IV U20606 ( .A(n17301), .Z(n17303) );
  XNOR U20607 ( .A(b[794]), .B(n17301), .Z(n17302) );
  XOR U20608 ( .A(n17304), .B(n17305), .Z(n17301) );
  ANDN U20609 ( .B(n17306), .A(n236), .Z(n17304) );
  XNOR U20610 ( .A(a[793]), .B(n17307), .Z(n236) );
  IV U20611 ( .A(n17305), .Z(n17307) );
  XNOR U20612 ( .A(b[793]), .B(n17305), .Z(n17306) );
  XOR U20613 ( .A(n17308), .B(n17309), .Z(n17305) );
  ANDN U20614 ( .B(n17310), .A(n237), .Z(n17308) );
  XNOR U20615 ( .A(a[792]), .B(n17311), .Z(n237) );
  IV U20616 ( .A(n17309), .Z(n17311) );
  XNOR U20617 ( .A(b[792]), .B(n17309), .Z(n17310) );
  XOR U20618 ( .A(n17312), .B(n17313), .Z(n17309) );
  ANDN U20619 ( .B(n17314), .A(n238), .Z(n17312) );
  XNOR U20620 ( .A(a[791]), .B(n17315), .Z(n238) );
  IV U20621 ( .A(n17313), .Z(n17315) );
  XNOR U20622 ( .A(b[791]), .B(n17313), .Z(n17314) );
  XOR U20623 ( .A(n17316), .B(n17317), .Z(n17313) );
  ANDN U20624 ( .B(n17318), .A(n239), .Z(n17316) );
  XNOR U20625 ( .A(a[790]), .B(n17319), .Z(n239) );
  IV U20626 ( .A(n17317), .Z(n17319) );
  XNOR U20627 ( .A(b[790]), .B(n17317), .Z(n17318) );
  XOR U20628 ( .A(n17320), .B(n17321), .Z(n17317) );
  ANDN U20629 ( .B(n17322), .A(n241), .Z(n17320) );
  XNOR U20630 ( .A(a[789]), .B(n17323), .Z(n241) );
  IV U20631 ( .A(n17321), .Z(n17323) );
  XNOR U20632 ( .A(b[789]), .B(n17321), .Z(n17322) );
  XOR U20633 ( .A(n17324), .B(n17325), .Z(n17321) );
  ANDN U20634 ( .B(n17326), .A(n242), .Z(n17324) );
  XNOR U20635 ( .A(a[788]), .B(n17327), .Z(n242) );
  IV U20636 ( .A(n17325), .Z(n17327) );
  XNOR U20637 ( .A(b[788]), .B(n17325), .Z(n17326) );
  XOR U20638 ( .A(n17328), .B(n17329), .Z(n17325) );
  ANDN U20639 ( .B(n17330), .A(n243), .Z(n17328) );
  XNOR U20640 ( .A(a[787]), .B(n17331), .Z(n243) );
  IV U20641 ( .A(n17329), .Z(n17331) );
  XNOR U20642 ( .A(b[787]), .B(n17329), .Z(n17330) );
  XOR U20643 ( .A(n17332), .B(n17333), .Z(n17329) );
  ANDN U20644 ( .B(n17334), .A(n244), .Z(n17332) );
  XNOR U20645 ( .A(a[786]), .B(n17335), .Z(n244) );
  IV U20646 ( .A(n17333), .Z(n17335) );
  XNOR U20647 ( .A(b[786]), .B(n17333), .Z(n17334) );
  XOR U20648 ( .A(n17336), .B(n17337), .Z(n17333) );
  ANDN U20649 ( .B(n17338), .A(n245), .Z(n17336) );
  XNOR U20650 ( .A(a[785]), .B(n17339), .Z(n245) );
  IV U20651 ( .A(n17337), .Z(n17339) );
  XNOR U20652 ( .A(b[785]), .B(n17337), .Z(n17338) );
  XOR U20653 ( .A(n17340), .B(n17341), .Z(n17337) );
  ANDN U20654 ( .B(n17342), .A(n246), .Z(n17340) );
  XNOR U20655 ( .A(a[784]), .B(n17343), .Z(n246) );
  IV U20656 ( .A(n17341), .Z(n17343) );
  XNOR U20657 ( .A(b[784]), .B(n17341), .Z(n17342) );
  XOR U20658 ( .A(n17344), .B(n17345), .Z(n17341) );
  ANDN U20659 ( .B(n17346), .A(n247), .Z(n17344) );
  XNOR U20660 ( .A(a[783]), .B(n17347), .Z(n247) );
  IV U20661 ( .A(n17345), .Z(n17347) );
  XNOR U20662 ( .A(b[783]), .B(n17345), .Z(n17346) );
  XOR U20663 ( .A(n17348), .B(n17349), .Z(n17345) );
  ANDN U20664 ( .B(n17350), .A(n248), .Z(n17348) );
  XNOR U20665 ( .A(a[782]), .B(n17351), .Z(n248) );
  IV U20666 ( .A(n17349), .Z(n17351) );
  XNOR U20667 ( .A(b[782]), .B(n17349), .Z(n17350) );
  XOR U20668 ( .A(n17352), .B(n17353), .Z(n17349) );
  ANDN U20669 ( .B(n17354), .A(n249), .Z(n17352) );
  XNOR U20670 ( .A(a[781]), .B(n17355), .Z(n249) );
  IV U20671 ( .A(n17353), .Z(n17355) );
  XNOR U20672 ( .A(b[781]), .B(n17353), .Z(n17354) );
  XOR U20673 ( .A(n17356), .B(n17357), .Z(n17353) );
  ANDN U20674 ( .B(n17358), .A(n250), .Z(n17356) );
  XNOR U20675 ( .A(a[780]), .B(n17359), .Z(n250) );
  IV U20676 ( .A(n17357), .Z(n17359) );
  XNOR U20677 ( .A(b[780]), .B(n17357), .Z(n17358) );
  XOR U20678 ( .A(n17360), .B(n17361), .Z(n17357) );
  ANDN U20679 ( .B(n17362), .A(n252), .Z(n17360) );
  XNOR U20680 ( .A(a[779]), .B(n17363), .Z(n252) );
  IV U20681 ( .A(n17361), .Z(n17363) );
  XNOR U20682 ( .A(b[779]), .B(n17361), .Z(n17362) );
  XOR U20683 ( .A(n17364), .B(n17365), .Z(n17361) );
  ANDN U20684 ( .B(n17366), .A(n253), .Z(n17364) );
  XNOR U20685 ( .A(a[778]), .B(n17367), .Z(n253) );
  IV U20686 ( .A(n17365), .Z(n17367) );
  XNOR U20687 ( .A(b[778]), .B(n17365), .Z(n17366) );
  XOR U20688 ( .A(n17368), .B(n17369), .Z(n17365) );
  ANDN U20689 ( .B(n17370), .A(n254), .Z(n17368) );
  XNOR U20690 ( .A(a[777]), .B(n17371), .Z(n254) );
  IV U20691 ( .A(n17369), .Z(n17371) );
  XNOR U20692 ( .A(b[777]), .B(n17369), .Z(n17370) );
  XOR U20693 ( .A(n17372), .B(n17373), .Z(n17369) );
  ANDN U20694 ( .B(n17374), .A(n255), .Z(n17372) );
  XNOR U20695 ( .A(a[776]), .B(n17375), .Z(n255) );
  IV U20696 ( .A(n17373), .Z(n17375) );
  XNOR U20697 ( .A(b[776]), .B(n17373), .Z(n17374) );
  XOR U20698 ( .A(n17376), .B(n17377), .Z(n17373) );
  ANDN U20699 ( .B(n17378), .A(n256), .Z(n17376) );
  XNOR U20700 ( .A(a[775]), .B(n17379), .Z(n256) );
  IV U20701 ( .A(n17377), .Z(n17379) );
  XNOR U20702 ( .A(b[775]), .B(n17377), .Z(n17378) );
  XOR U20703 ( .A(n17380), .B(n17381), .Z(n17377) );
  ANDN U20704 ( .B(n17382), .A(n257), .Z(n17380) );
  XNOR U20705 ( .A(a[774]), .B(n17383), .Z(n257) );
  IV U20706 ( .A(n17381), .Z(n17383) );
  XNOR U20707 ( .A(b[774]), .B(n17381), .Z(n17382) );
  XOR U20708 ( .A(n17384), .B(n17385), .Z(n17381) );
  ANDN U20709 ( .B(n17386), .A(n258), .Z(n17384) );
  XNOR U20710 ( .A(a[773]), .B(n17387), .Z(n258) );
  IV U20711 ( .A(n17385), .Z(n17387) );
  XNOR U20712 ( .A(b[773]), .B(n17385), .Z(n17386) );
  XOR U20713 ( .A(n17388), .B(n17389), .Z(n17385) );
  ANDN U20714 ( .B(n17390), .A(n259), .Z(n17388) );
  XNOR U20715 ( .A(a[772]), .B(n17391), .Z(n259) );
  IV U20716 ( .A(n17389), .Z(n17391) );
  XNOR U20717 ( .A(b[772]), .B(n17389), .Z(n17390) );
  XOR U20718 ( .A(n17392), .B(n17393), .Z(n17389) );
  ANDN U20719 ( .B(n17394), .A(n260), .Z(n17392) );
  XNOR U20720 ( .A(a[771]), .B(n17395), .Z(n260) );
  IV U20721 ( .A(n17393), .Z(n17395) );
  XNOR U20722 ( .A(b[771]), .B(n17393), .Z(n17394) );
  XOR U20723 ( .A(n17396), .B(n17397), .Z(n17393) );
  ANDN U20724 ( .B(n17398), .A(n261), .Z(n17396) );
  XNOR U20725 ( .A(a[770]), .B(n17399), .Z(n261) );
  IV U20726 ( .A(n17397), .Z(n17399) );
  XNOR U20727 ( .A(b[770]), .B(n17397), .Z(n17398) );
  XOR U20728 ( .A(n17400), .B(n17401), .Z(n17397) );
  ANDN U20729 ( .B(n17402), .A(n263), .Z(n17400) );
  XNOR U20730 ( .A(a[769]), .B(n17403), .Z(n263) );
  IV U20731 ( .A(n17401), .Z(n17403) );
  XNOR U20732 ( .A(b[769]), .B(n17401), .Z(n17402) );
  XOR U20733 ( .A(n17404), .B(n17405), .Z(n17401) );
  ANDN U20734 ( .B(n17406), .A(n264), .Z(n17404) );
  XNOR U20735 ( .A(a[768]), .B(n17407), .Z(n264) );
  IV U20736 ( .A(n17405), .Z(n17407) );
  XNOR U20737 ( .A(b[768]), .B(n17405), .Z(n17406) );
  XOR U20738 ( .A(n17408), .B(n17409), .Z(n17405) );
  ANDN U20739 ( .B(n17410), .A(n265), .Z(n17408) );
  XNOR U20740 ( .A(a[767]), .B(n17411), .Z(n265) );
  IV U20741 ( .A(n17409), .Z(n17411) );
  XNOR U20742 ( .A(b[767]), .B(n17409), .Z(n17410) );
  XOR U20743 ( .A(n17412), .B(n17413), .Z(n17409) );
  ANDN U20744 ( .B(n17414), .A(n266), .Z(n17412) );
  XNOR U20745 ( .A(a[766]), .B(n17415), .Z(n266) );
  IV U20746 ( .A(n17413), .Z(n17415) );
  XNOR U20747 ( .A(b[766]), .B(n17413), .Z(n17414) );
  XOR U20748 ( .A(n17416), .B(n17417), .Z(n17413) );
  ANDN U20749 ( .B(n17418), .A(n267), .Z(n17416) );
  XNOR U20750 ( .A(a[765]), .B(n17419), .Z(n267) );
  IV U20751 ( .A(n17417), .Z(n17419) );
  XNOR U20752 ( .A(b[765]), .B(n17417), .Z(n17418) );
  XOR U20753 ( .A(n17420), .B(n17421), .Z(n17417) );
  ANDN U20754 ( .B(n17422), .A(n268), .Z(n17420) );
  XNOR U20755 ( .A(a[764]), .B(n17423), .Z(n268) );
  IV U20756 ( .A(n17421), .Z(n17423) );
  XNOR U20757 ( .A(b[764]), .B(n17421), .Z(n17422) );
  XOR U20758 ( .A(n17424), .B(n17425), .Z(n17421) );
  ANDN U20759 ( .B(n17426), .A(n269), .Z(n17424) );
  XNOR U20760 ( .A(a[763]), .B(n17427), .Z(n269) );
  IV U20761 ( .A(n17425), .Z(n17427) );
  XNOR U20762 ( .A(b[763]), .B(n17425), .Z(n17426) );
  XOR U20763 ( .A(n17428), .B(n17429), .Z(n17425) );
  ANDN U20764 ( .B(n17430), .A(n270), .Z(n17428) );
  XNOR U20765 ( .A(a[762]), .B(n17431), .Z(n270) );
  IV U20766 ( .A(n17429), .Z(n17431) );
  XNOR U20767 ( .A(b[762]), .B(n17429), .Z(n17430) );
  XOR U20768 ( .A(n17432), .B(n17433), .Z(n17429) );
  ANDN U20769 ( .B(n17434), .A(n271), .Z(n17432) );
  XNOR U20770 ( .A(a[761]), .B(n17435), .Z(n271) );
  IV U20771 ( .A(n17433), .Z(n17435) );
  XNOR U20772 ( .A(b[761]), .B(n17433), .Z(n17434) );
  XOR U20773 ( .A(n17436), .B(n17437), .Z(n17433) );
  ANDN U20774 ( .B(n17438), .A(n272), .Z(n17436) );
  XNOR U20775 ( .A(a[760]), .B(n17439), .Z(n272) );
  IV U20776 ( .A(n17437), .Z(n17439) );
  XNOR U20777 ( .A(b[760]), .B(n17437), .Z(n17438) );
  XOR U20778 ( .A(n17440), .B(n17441), .Z(n17437) );
  ANDN U20779 ( .B(n17442), .A(n274), .Z(n17440) );
  XNOR U20780 ( .A(a[759]), .B(n17443), .Z(n274) );
  IV U20781 ( .A(n17441), .Z(n17443) );
  XNOR U20782 ( .A(b[759]), .B(n17441), .Z(n17442) );
  XOR U20783 ( .A(n17444), .B(n17445), .Z(n17441) );
  ANDN U20784 ( .B(n17446), .A(n275), .Z(n17444) );
  XNOR U20785 ( .A(a[758]), .B(n17447), .Z(n275) );
  IV U20786 ( .A(n17445), .Z(n17447) );
  XNOR U20787 ( .A(b[758]), .B(n17445), .Z(n17446) );
  XOR U20788 ( .A(n17448), .B(n17449), .Z(n17445) );
  ANDN U20789 ( .B(n17450), .A(n276), .Z(n17448) );
  XNOR U20790 ( .A(a[757]), .B(n17451), .Z(n276) );
  IV U20791 ( .A(n17449), .Z(n17451) );
  XNOR U20792 ( .A(b[757]), .B(n17449), .Z(n17450) );
  XOR U20793 ( .A(n17452), .B(n17453), .Z(n17449) );
  ANDN U20794 ( .B(n17454), .A(n277), .Z(n17452) );
  XNOR U20795 ( .A(a[756]), .B(n17455), .Z(n277) );
  IV U20796 ( .A(n17453), .Z(n17455) );
  XNOR U20797 ( .A(b[756]), .B(n17453), .Z(n17454) );
  XOR U20798 ( .A(n17456), .B(n17457), .Z(n17453) );
  ANDN U20799 ( .B(n17458), .A(n278), .Z(n17456) );
  XNOR U20800 ( .A(a[755]), .B(n17459), .Z(n278) );
  IV U20801 ( .A(n17457), .Z(n17459) );
  XNOR U20802 ( .A(b[755]), .B(n17457), .Z(n17458) );
  XOR U20803 ( .A(n17460), .B(n17461), .Z(n17457) );
  ANDN U20804 ( .B(n17462), .A(n279), .Z(n17460) );
  XNOR U20805 ( .A(a[754]), .B(n17463), .Z(n279) );
  IV U20806 ( .A(n17461), .Z(n17463) );
  XNOR U20807 ( .A(b[754]), .B(n17461), .Z(n17462) );
  XOR U20808 ( .A(n17464), .B(n17465), .Z(n17461) );
  ANDN U20809 ( .B(n17466), .A(n280), .Z(n17464) );
  XNOR U20810 ( .A(a[753]), .B(n17467), .Z(n280) );
  IV U20811 ( .A(n17465), .Z(n17467) );
  XNOR U20812 ( .A(b[753]), .B(n17465), .Z(n17466) );
  XOR U20813 ( .A(n17468), .B(n17469), .Z(n17465) );
  ANDN U20814 ( .B(n17470), .A(n281), .Z(n17468) );
  XNOR U20815 ( .A(a[752]), .B(n17471), .Z(n281) );
  IV U20816 ( .A(n17469), .Z(n17471) );
  XNOR U20817 ( .A(b[752]), .B(n17469), .Z(n17470) );
  XOR U20818 ( .A(n17472), .B(n17473), .Z(n17469) );
  ANDN U20819 ( .B(n17474), .A(n282), .Z(n17472) );
  XNOR U20820 ( .A(a[751]), .B(n17475), .Z(n282) );
  IV U20821 ( .A(n17473), .Z(n17475) );
  XNOR U20822 ( .A(b[751]), .B(n17473), .Z(n17474) );
  XOR U20823 ( .A(n17476), .B(n17477), .Z(n17473) );
  ANDN U20824 ( .B(n17478), .A(n283), .Z(n17476) );
  XNOR U20825 ( .A(a[750]), .B(n17479), .Z(n283) );
  IV U20826 ( .A(n17477), .Z(n17479) );
  XNOR U20827 ( .A(b[750]), .B(n17477), .Z(n17478) );
  XOR U20828 ( .A(n17480), .B(n17481), .Z(n17477) );
  ANDN U20829 ( .B(n17482), .A(n285), .Z(n17480) );
  XNOR U20830 ( .A(a[749]), .B(n17483), .Z(n285) );
  IV U20831 ( .A(n17481), .Z(n17483) );
  XNOR U20832 ( .A(b[749]), .B(n17481), .Z(n17482) );
  XOR U20833 ( .A(n17484), .B(n17485), .Z(n17481) );
  ANDN U20834 ( .B(n17486), .A(n286), .Z(n17484) );
  XNOR U20835 ( .A(a[748]), .B(n17487), .Z(n286) );
  IV U20836 ( .A(n17485), .Z(n17487) );
  XNOR U20837 ( .A(b[748]), .B(n17485), .Z(n17486) );
  XOR U20838 ( .A(n17488), .B(n17489), .Z(n17485) );
  ANDN U20839 ( .B(n17490), .A(n287), .Z(n17488) );
  XNOR U20840 ( .A(a[747]), .B(n17491), .Z(n287) );
  IV U20841 ( .A(n17489), .Z(n17491) );
  XNOR U20842 ( .A(b[747]), .B(n17489), .Z(n17490) );
  XOR U20843 ( .A(n17492), .B(n17493), .Z(n17489) );
  ANDN U20844 ( .B(n17494), .A(n288), .Z(n17492) );
  XNOR U20845 ( .A(a[746]), .B(n17495), .Z(n288) );
  IV U20846 ( .A(n17493), .Z(n17495) );
  XNOR U20847 ( .A(b[746]), .B(n17493), .Z(n17494) );
  XOR U20848 ( .A(n17496), .B(n17497), .Z(n17493) );
  ANDN U20849 ( .B(n17498), .A(n289), .Z(n17496) );
  XNOR U20850 ( .A(a[745]), .B(n17499), .Z(n289) );
  IV U20851 ( .A(n17497), .Z(n17499) );
  XNOR U20852 ( .A(b[745]), .B(n17497), .Z(n17498) );
  XOR U20853 ( .A(n17500), .B(n17501), .Z(n17497) );
  ANDN U20854 ( .B(n17502), .A(n290), .Z(n17500) );
  XNOR U20855 ( .A(a[744]), .B(n17503), .Z(n290) );
  IV U20856 ( .A(n17501), .Z(n17503) );
  XNOR U20857 ( .A(b[744]), .B(n17501), .Z(n17502) );
  XOR U20858 ( .A(n17504), .B(n17505), .Z(n17501) );
  ANDN U20859 ( .B(n17506), .A(n291), .Z(n17504) );
  XNOR U20860 ( .A(a[743]), .B(n17507), .Z(n291) );
  IV U20861 ( .A(n17505), .Z(n17507) );
  XNOR U20862 ( .A(b[743]), .B(n17505), .Z(n17506) );
  XOR U20863 ( .A(n17508), .B(n17509), .Z(n17505) );
  ANDN U20864 ( .B(n17510), .A(n292), .Z(n17508) );
  XNOR U20865 ( .A(a[742]), .B(n17511), .Z(n292) );
  IV U20866 ( .A(n17509), .Z(n17511) );
  XNOR U20867 ( .A(b[742]), .B(n17509), .Z(n17510) );
  XOR U20868 ( .A(n17512), .B(n17513), .Z(n17509) );
  ANDN U20869 ( .B(n17514), .A(n293), .Z(n17512) );
  XNOR U20870 ( .A(a[741]), .B(n17515), .Z(n293) );
  IV U20871 ( .A(n17513), .Z(n17515) );
  XNOR U20872 ( .A(b[741]), .B(n17513), .Z(n17514) );
  XOR U20873 ( .A(n17516), .B(n17517), .Z(n17513) );
  ANDN U20874 ( .B(n17518), .A(n294), .Z(n17516) );
  XNOR U20875 ( .A(a[740]), .B(n17519), .Z(n294) );
  IV U20876 ( .A(n17517), .Z(n17519) );
  XNOR U20877 ( .A(b[740]), .B(n17517), .Z(n17518) );
  XOR U20878 ( .A(n17520), .B(n17521), .Z(n17517) );
  ANDN U20879 ( .B(n17522), .A(n296), .Z(n17520) );
  XNOR U20880 ( .A(a[739]), .B(n17523), .Z(n296) );
  IV U20881 ( .A(n17521), .Z(n17523) );
  XNOR U20882 ( .A(b[739]), .B(n17521), .Z(n17522) );
  XOR U20883 ( .A(n17524), .B(n17525), .Z(n17521) );
  ANDN U20884 ( .B(n17526), .A(n297), .Z(n17524) );
  XNOR U20885 ( .A(a[738]), .B(n17527), .Z(n297) );
  IV U20886 ( .A(n17525), .Z(n17527) );
  XNOR U20887 ( .A(b[738]), .B(n17525), .Z(n17526) );
  XOR U20888 ( .A(n17528), .B(n17529), .Z(n17525) );
  ANDN U20889 ( .B(n17530), .A(n298), .Z(n17528) );
  XNOR U20890 ( .A(a[737]), .B(n17531), .Z(n298) );
  IV U20891 ( .A(n17529), .Z(n17531) );
  XNOR U20892 ( .A(b[737]), .B(n17529), .Z(n17530) );
  XOR U20893 ( .A(n17532), .B(n17533), .Z(n17529) );
  ANDN U20894 ( .B(n17534), .A(n299), .Z(n17532) );
  XNOR U20895 ( .A(a[736]), .B(n17535), .Z(n299) );
  IV U20896 ( .A(n17533), .Z(n17535) );
  XNOR U20897 ( .A(b[736]), .B(n17533), .Z(n17534) );
  XOR U20898 ( .A(n17536), .B(n17537), .Z(n17533) );
  ANDN U20899 ( .B(n17538), .A(n300), .Z(n17536) );
  XNOR U20900 ( .A(a[735]), .B(n17539), .Z(n300) );
  IV U20901 ( .A(n17537), .Z(n17539) );
  XNOR U20902 ( .A(b[735]), .B(n17537), .Z(n17538) );
  XOR U20903 ( .A(n17540), .B(n17541), .Z(n17537) );
  ANDN U20904 ( .B(n17542), .A(n301), .Z(n17540) );
  XNOR U20905 ( .A(a[734]), .B(n17543), .Z(n301) );
  IV U20906 ( .A(n17541), .Z(n17543) );
  XNOR U20907 ( .A(b[734]), .B(n17541), .Z(n17542) );
  XOR U20908 ( .A(n17544), .B(n17545), .Z(n17541) );
  ANDN U20909 ( .B(n17546), .A(n302), .Z(n17544) );
  XNOR U20910 ( .A(a[733]), .B(n17547), .Z(n302) );
  IV U20911 ( .A(n17545), .Z(n17547) );
  XNOR U20912 ( .A(b[733]), .B(n17545), .Z(n17546) );
  XOR U20913 ( .A(n17548), .B(n17549), .Z(n17545) );
  ANDN U20914 ( .B(n17550), .A(n303), .Z(n17548) );
  XNOR U20915 ( .A(a[732]), .B(n17551), .Z(n303) );
  IV U20916 ( .A(n17549), .Z(n17551) );
  XNOR U20917 ( .A(b[732]), .B(n17549), .Z(n17550) );
  XOR U20918 ( .A(n17552), .B(n17553), .Z(n17549) );
  ANDN U20919 ( .B(n17554), .A(n304), .Z(n17552) );
  XNOR U20920 ( .A(a[731]), .B(n17555), .Z(n304) );
  IV U20921 ( .A(n17553), .Z(n17555) );
  XNOR U20922 ( .A(b[731]), .B(n17553), .Z(n17554) );
  XOR U20923 ( .A(n17556), .B(n17557), .Z(n17553) );
  ANDN U20924 ( .B(n17558), .A(n305), .Z(n17556) );
  XNOR U20925 ( .A(a[730]), .B(n17559), .Z(n305) );
  IV U20926 ( .A(n17557), .Z(n17559) );
  XNOR U20927 ( .A(b[730]), .B(n17557), .Z(n17558) );
  XOR U20928 ( .A(n17560), .B(n17561), .Z(n17557) );
  ANDN U20929 ( .B(n17562), .A(n307), .Z(n17560) );
  XNOR U20930 ( .A(a[729]), .B(n17563), .Z(n307) );
  IV U20931 ( .A(n17561), .Z(n17563) );
  XNOR U20932 ( .A(b[729]), .B(n17561), .Z(n17562) );
  XOR U20933 ( .A(n17564), .B(n17565), .Z(n17561) );
  ANDN U20934 ( .B(n17566), .A(n308), .Z(n17564) );
  XNOR U20935 ( .A(a[728]), .B(n17567), .Z(n308) );
  IV U20936 ( .A(n17565), .Z(n17567) );
  XNOR U20937 ( .A(b[728]), .B(n17565), .Z(n17566) );
  XOR U20938 ( .A(n17568), .B(n17569), .Z(n17565) );
  ANDN U20939 ( .B(n17570), .A(n309), .Z(n17568) );
  XNOR U20940 ( .A(a[727]), .B(n17571), .Z(n309) );
  IV U20941 ( .A(n17569), .Z(n17571) );
  XNOR U20942 ( .A(b[727]), .B(n17569), .Z(n17570) );
  XOR U20943 ( .A(n17572), .B(n17573), .Z(n17569) );
  ANDN U20944 ( .B(n17574), .A(n310), .Z(n17572) );
  XNOR U20945 ( .A(a[726]), .B(n17575), .Z(n310) );
  IV U20946 ( .A(n17573), .Z(n17575) );
  XNOR U20947 ( .A(b[726]), .B(n17573), .Z(n17574) );
  XOR U20948 ( .A(n17576), .B(n17577), .Z(n17573) );
  ANDN U20949 ( .B(n17578), .A(n311), .Z(n17576) );
  XNOR U20950 ( .A(a[725]), .B(n17579), .Z(n311) );
  IV U20951 ( .A(n17577), .Z(n17579) );
  XNOR U20952 ( .A(b[725]), .B(n17577), .Z(n17578) );
  XOR U20953 ( .A(n17580), .B(n17581), .Z(n17577) );
  ANDN U20954 ( .B(n17582), .A(n312), .Z(n17580) );
  XNOR U20955 ( .A(a[724]), .B(n17583), .Z(n312) );
  IV U20956 ( .A(n17581), .Z(n17583) );
  XNOR U20957 ( .A(b[724]), .B(n17581), .Z(n17582) );
  XOR U20958 ( .A(n17584), .B(n17585), .Z(n17581) );
  ANDN U20959 ( .B(n17586), .A(n313), .Z(n17584) );
  XNOR U20960 ( .A(a[723]), .B(n17587), .Z(n313) );
  IV U20961 ( .A(n17585), .Z(n17587) );
  XNOR U20962 ( .A(b[723]), .B(n17585), .Z(n17586) );
  XOR U20963 ( .A(n17588), .B(n17589), .Z(n17585) );
  ANDN U20964 ( .B(n17590), .A(n314), .Z(n17588) );
  XNOR U20965 ( .A(a[722]), .B(n17591), .Z(n314) );
  IV U20966 ( .A(n17589), .Z(n17591) );
  XNOR U20967 ( .A(b[722]), .B(n17589), .Z(n17590) );
  XOR U20968 ( .A(n17592), .B(n17593), .Z(n17589) );
  ANDN U20969 ( .B(n17594), .A(n315), .Z(n17592) );
  XNOR U20970 ( .A(a[721]), .B(n17595), .Z(n315) );
  IV U20971 ( .A(n17593), .Z(n17595) );
  XNOR U20972 ( .A(b[721]), .B(n17593), .Z(n17594) );
  XOR U20973 ( .A(n17596), .B(n17597), .Z(n17593) );
  ANDN U20974 ( .B(n17598), .A(n316), .Z(n17596) );
  XNOR U20975 ( .A(a[720]), .B(n17599), .Z(n316) );
  IV U20976 ( .A(n17597), .Z(n17599) );
  XNOR U20977 ( .A(b[720]), .B(n17597), .Z(n17598) );
  XOR U20978 ( .A(n17600), .B(n17601), .Z(n17597) );
  ANDN U20979 ( .B(n17602), .A(n318), .Z(n17600) );
  XNOR U20980 ( .A(a[719]), .B(n17603), .Z(n318) );
  IV U20981 ( .A(n17601), .Z(n17603) );
  XNOR U20982 ( .A(b[719]), .B(n17601), .Z(n17602) );
  XOR U20983 ( .A(n17604), .B(n17605), .Z(n17601) );
  ANDN U20984 ( .B(n17606), .A(n319), .Z(n17604) );
  XNOR U20985 ( .A(a[718]), .B(n17607), .Z(n319) );
  IV U20986 ( .A(n17605), .Z(n17607) );
  XNOR U20987 ( .A(b[718]), .B(n17605), .Z(n17606) );
  XOR U20988 ( .A(n17608), .B(n17609), .Z(n17605) );
  ANDN U20989 ( .B(n17610), .A(n320), .Z(n17608) );
  XNOR U20990 ( .A(a[717]), .B(n17611), .Z(n320) );
  IV U20991 ( .A(n17609), .Z(n17611) );
  XNOR U20992 ( .A(b[717]), .B(n17609), .Z(n17610) );
  XOR U20993 ( .A(n17612), .B(n17613), .Z(n17609) );
  ANDN U20994 ( .B(n17614), .A(n321), .Z(n17612) );
  XNOR U20995 ( .A(a[716]), .B(n17615), .Z(n321) );
  IV U20996 ( .A(n17613), .Z(n17615) );
  XNOR U20997 ( .A(b[716]), .B(n17613), .Z(n17614) );
  XOR U20998 ( .A(n17616), .B(n17617), .Z(n17613) );
  ANDN U20999 ( .B(n17618), .A(n322), .Z(n17616) );
  XNOR U21000 ( .A(a[715]), .B(n17619), .Z(n322) );
  IV U21001 ( .A(n17617), .Z(n17619) );
  XNOR U21002 ( .A(b[715]), .B(n17617), .Z(n17618) );
  XOR U21003 ( .A(n17620), .B(n17621), .Z(n17617) );
  ANDN U21004 ( .B(n17622), .A(n323), .Z(n17620) );
  XNOR U21005 ( .A(a[714]), .B(n17623), .Z(n323) );
  IV U21006 ( .A(n17621), .Z(n17623) );
  XNOR U21007 ( .A(b[714]), .B(n17621), .Z(n17622) );
  XOR U21008 ( .A(n17624), .B(n17625), .Z(n17621) );
  ANDN U21009 ( .B(n17626), .A(n324), .Z(n17624) );
  XNOR U21010 ( .A(a[713]), .B(n17627), .Z(n324) );
  IV U21011 ( .A(n17625), .Z(n17627) );
  XNOR U21012 ( .A(b[713]), .B(n17625), .Z(n17626) );
  XOR U21013 ( .A(n17628), .B(n17629), .Z(n17625) );
  ANDN U21014 ( .B(n17630), .A(n325), .Z(n17628) );
  XNOR U21015 ( .A(a[712]), .B(n17631), .Z(n325) );
  IV U21016 ( .A(n17629), .Z(n17631) );
  XNOR U21017 ( .A(b[712]), .B(n17629), .Z(n17630) );
  XOR U21018 ( .A(n17632), .B(n17633), .Z(n17629) );
  ANDN U21019 ( .B(n17634), .A(n326), .Z(n17632) );
  XNOR U21020 ( .A(a[711]), .B(n17635), .Z(n326) );
  IV U21021 ( .A(n17633), .Z(n17635) );
  XNOR U21022 ( .A(b[711]), .B(n17633), .Z(n17634) );
  XOR U21023 ( .A(n17636), .B(n17637), .Z(n17633) );
  ANDN U21024 ( .B(n17638), .A(n327), .Z(n17636) );
  XNOR U21025 ( .A(a[710]), .B(n17639), .Z(n327) );
  IV U21026 ( .A(n17637), .Z(n17639) );
  XNOR U21027 ( .A(b[710]), .B(n17637), .Z(n17638) );
  XOR U21028 ( .A(n17640), .B(n17641), .Z(n17637) );
  ANDN U21029 ( .B(n17642), .A(n329), .Z(n17640) );
  XNOR U21030 ( .A(a[709]), .B(n17643), .Z(n329) );
  IV U21031 ( .A(n17641), .Z(n17643) );
  XNOR U21032 ( .A(b[709]), .B(n17641), .Z(n17642) );
  XOR U21033 ( .A(n17644), .B(n17645), .Z(n17641) );
  ANDN U21034 ( .B(n17646), .A(n330), .Z(n17644) );
  XNOR U21035 ( .A(a[708]), .B(n17647), .Z(n330) );
  IV U21036 ( .A(n17645), .Z(n17647) );
  XNOR U21037 ( .A(b[708]), .B(n17645), .Z(n17646) );
  XOR U21038 ( .A(n17648), .B(n17649), .Z(n17645) );
  ANDN U21039 ( .B(n17650), .A(n331), .Z(n17648) );
  XNOR U21040 ( .A(a[707]), .B(n17651), .Z(n331) );
  IV U21041 ( .A(n17649), .Z(n17651) );
  XNOR U21042 ( .A(b[707]), .B(n17649), .Z(n17650) );
  XOR U21043 ( .A(n17652), .B(n17653), .Z(n17649) );
  ANDN U21044 ( .B(n17654), .A(n332), .Z(n17652) );
  XNOR U21045 ( .A(a[706]), .B(n17655), .Z(n332) );
  IV U21046 ( .A(n17653), .Z(n17655) );
  XNOR U21047 ( .A(b[706]), .B(n17653), .Z(n17654) );
  XOR U21048 ( .A(n17656), .B(n17657), .Z(n17653) );
  ANDN U21049 ( .B(n17658), .A(n333), .Z(n17656) );
  XNOR U21050 ( .A(a[705]), .B(n17659), .Z(n333) );
  IV U21051 ( .A(n17657), .Z(n17659) );
  XNOR U21052 ( .A(b[705]), .B(n17657), .Z(n17658) );
  XOR U21053 ( .A(n17660), .B(n17661), .Z(n17657) );
  ANDN U21054 ( .B(n17662), .A(n334), .Z(n17660) );
  XNOR U21055 ( .A(a[704]), .B(n17663), .Z(n334) );
  IV U21056 ( .A(n17661), .Z(n17663) );
  XNOR U21057 ( .A(b[704]), .B(n17661), .Z(n17662) );
  XOR U21058 ( .A(n17664), .B(n17665), .Z(n17661) );
  ANDN U21059 ( .B(n17666), .A(n335), .Z(n17664) );
  XNOR U21060 ( .A(a[703]), .B(n17667), .Z(n335) );
  IV U21061 ( .A(n17665), .Z(n17667) );
  XNOR U21062 ( .A(b[703]), .B(n17665), .Z(n17666) );
  XOR U21063 ( .A(n17668), .B(n17669), .Z(n17665) );
  ANDN U21064 ( .B(n17670), .A(n336), .Z(n17668) );
  XNOR U21065 ( .A(a[702]), .B(n17671), .Z(n336) );
  IV U21066 ( .A(n17669), .Z(n17671) );
  XNOR U21067 ( .A(b[702]), .B(n17669), .Z(n17670) );
  XOR U21068 ( .A(n17672), .B(n17673), .Z(n17669) );
  ANDN U21069 ( .B(n17674), .A(n337), .Z(n17672) );
  XNOR U21070 ( .A(a[701]), .B(n17675), .Z(n337) );
  IV U21071 ( .A(n17673), .Z(n17675) );
  XNOR U21072 ( .A(b[701]), .B(n17673), .Z(n17674) );
  XOR U21073 ( .A(n17676), .B(n17677), .Z(n17673) );
  ANDN U21074 ( .B(n17678), .A(n338), .Z(n17676) );
  XNOR U21075 ( .A(a[700]), .B(n17679), .Z(n338) );
  IV U21076 ( .A(n17677), .Z(n17679) );
  XNOR U21077 ( .A(b[700]), .B(n17677), .Z(n17678) );
  XOR U21078 ( .A(n17680), .B(n17681), .Z(n17677) );
  ANDN U21079 ( .B(n17682), .A(n341), .Z(n17680) );
  XNOR U21080 ( .A(a[699]), .B(n17683), .Z(n341) );
  IV U21081 ( .A(n17681), .Z(n17683) );
  XNOR U21082 ( .A(b[699]), .B(n17681), .Z(n17682) );
  XOR U21083 ( .A(n17684), .B(n17685), .Z(n17681) );
  ANDN U21084 ( .B(n17686), .A(n342), .Z(n17684) );
  XNOR U21085 ( .A(a[698]), .B(n17687), .Z(n342) );
  IV U21086 ( .A(n17685), .Z(n17687) );
  XNOR U21087 ( .A(b[698]), .B(n17685), .Z(n17686) );
  XOR U21088 ( .A(n17688), .B(n17689), .Z(n17685) );
  ANDN U21089 ( .B(n17690), .A(n343), .Z(n17688) );
  XNOR U21090 ( .A(a[697]), .B(n17691), .Z(n343) );
  IV U21091 ( .A(n17689), .Z(n17691) );
  XNOR U21092 ( .A(b[697]), .B(n17689), .Z(n17690) );
  XOR U21093 ( .A(n17692), .B(n17693), .Z(n17689) );
  ANDN U21094 ( .B(n17694), .A(n344), .Z(n17692) );
  XNOR U21095 ( .A(a[696]), .B(n17695), .Z(n344) );
  IV U21096 ( .A(n17693), .Z(n17695) );
  XNOR U21097 ( .A(b[696]), .B(n17693), .Z(n17694) );
  XOR U21098 ( .A(n17696), .B(n17697), .Z(n17693) );
  ANDN U21099 ( .B(n17698), .A(n345), .Z(n17696) );
  XNOR U21100 ( .A(a[695]), .B(n17699), .Z(n345) );
  IV U21101 ( .A(n17697), .Z(n17699) );
  XNOR U21102 ( .A(b[695]), .B(n17697), .Z(n17698) );
  XOR U21103 ( .A(n17700), .B(n17701), .Z(n17697) );
  ANDN U21104 ( .B(n17702), .A(n346), .Z(n17700) );
  XNOR U21105 ( .A(a[694]), .B(n17703), .Z(n346) );
  IV U21106 ( .A(n17701), .Z(n17703) );
  XNOR U21107 ( .A(b[694]), .B(n17701), .Z(n17702) );
  XOR U21108 ( .A(n17704), .B(n17705), .Z(n17701) );
  ANDN U21109 ( .B(n17706), .A(n347), .Z(n17704) );
  XNOR U21110 ( .A(a[693]), .B(n17707), .Z(n347) );
  IV U21111 ( .A(n17705), .Z(n17707) );
  XNOR U21112 ( .A(b[693]), .B(n17705), .Z(n17706) );
  XOR U21113 ( .A(n17708), .B(n17709), .Z(n17705) );
  ANDN U21114 ( .B(n17710), .A(n348), .Z(n17708) );
  XNOR U21115 ( .A(a[692]), .B(n17711), .Z(n348) );
  IV U21116 ( .A(n17709), .Z(n17711) );
  XNOR U21117 ( .A(b[692]), .B(n17709), .Z(n17710) );
  XOR U21118 ( .A(n17712), .B(n17713), .Z(n17709) );
  ANDN U21119 ( .B(n17714), .A(n349), .Z(n17712) );
  XNOR U21120 ( .A(a[691]), .B(n17715), .Z(n349) );
  IV U21121 ( .A(n17713), .Z(n17715) );
  XNOR U21122 ( .A(b[691]), .B(n17713), .Z(n17714) );
  XOR U21123 ( .A(n17716), .B(n17717), .Z(n17713) );
  ANDN U21124 ( .B(n17718), .A(n350), .Z(n17716) );
  XNOR U21125 ( .A(a[690]), .B(n17719), .Z(n350) );
  IV U21126 ( .A(n17717), .Z(n17719) );
  XNOR U21127 ( .A(b[690]), .B(n17717), .Z(n17718) );
  XOR U21128 ( .A(n17720), .B(n17721), .Z(n17717) );
  ANDN U21129 ( .B(n17722), .A(n352), .Z(n17720) );
  XNOR U21130 ( .A(a[689]), .B(n17723), .Z(n352) );
  IV U21131 ( .A(n17721), .Z(n17723) );
  XNOR U21132 ( .A(b[689]), .B(n17721), .Z(n17722) );
  XOR U21133 ( .A(n17724), .B(n17725), .Z(n17721) );
  ANDN U21134 ( .B(n17726), .A(n353), .Z(n17724) );
  XNOR U21135 ( .A(a[688]), .B(n17727), .Z(n353) );
  IV U21136 ( .A(n17725), .Z(n17727) );
  XNOR U21137 ( .A(b[688]), .B(n17725), .Z(n17726) );
  XOR U21138 ( .A(n17728), .B(n17729), .Z(n17725) );
  ANDN U21139 ( .B(n17730), .A(n354), .Z(n17728) );
  XNOR U21140 ( .A(a[687]), .B(n17731), .Z(n354) );
  IV U21141 ( .A(n17729), .Z(n17731) );
  XNOR U21142 ( .A(b[687]), .B(n17729), .Z(n17730) );
  XOR U21143 ( .A(n17732), .B(n17733), .Z(n17729) );
  ANDN U21144 ( .B(n17734), .A(n355), .Z(n17732) );
  XNOR U21145 ( .A(a[686]), .B(n17735), .Z(n355) );
  IV U21146 ( .A(n17733), .Z(n17735) );
  XNOR U21147 ( .A(b[686]), .B(n17733), .Z(n17734) );
  XOR U21148 ( .A(n17736), .B(n17737), .Z(n17733) );
  ANDN U21149 ( .B(n17738), .A(n356), .Z(n17736) );
  XNOR U21150 ( .A(a[685]), .B(n17739), .Z(n356) );
  IV U21151 ( .A(n17737), .Z(n17739) );
  XNOR U21152 ( .A(b[685]), .B(n17737), .Z(n17738) );
  XOR U21153 ( .A(n17740), .B(n17741), .Z(n17737) );
  ANDN U21154 ( .B(n17742), .A(n357), .Z(n17740) );
  XNOR U21155 ( .A(a[684]), .B(n17743), .Z(n357) );
  IV U21156 ( .A(n17741), .Z(n17743) );
  XNOR U21157 ( .A(b[684]), .B(n17741), .Z(n17742) );
  XOR U21158 ( .A(n17744), .B(n17745), .Z(n17741) );
  ANDN U21159 ( .B(n17746), .A(n358), .Z(n17744) );
  XNOR U21160 ( .A(a[683]), .B(n17747), .Z(n358) );
  IV U21161 ( .A(n17745), .Z(n17747) );
  XNOR U21162 ( .A(b[683]), .B(n17745), .Z(n17746) );
  XOR U21163 ( .A(n17748), .B(n17749), .Z(n17745) );
  ANDN U21164 ( .B(n17750), .A(n359), .Z(n17748) );
  XNOR U21165 ( .A(a[682]), .B(n17751), .Z(n359) );
  IV U21166 ( .A(n17749), .Z(n17751) );
  XNOR U21167 ( .A(b[682]), .B(n17749), .Z(n17750) );
  XOR U21168 ( .A(n17752), .B(n17753), .Z(n17749) );
  ANDN U21169 ( .B(n17754), .A(n360), .Z(n17752) );
  XNOR U21170 ( .A(a[681]), .B(n17755), .Z(n360) );
  IV U21171 ( .A(n17753), .Z(n17755) );
  XNOR U21172 ( .A(b[681]), .B(n17753), .Z(n17754) );
  XOR U21173 ( .A(n17756), .B(n17757), .Z(n17753) );
  ANDN U21174 ( .B(n17758), .A(n361), .Z(n17756) );
  XNOR U21175 ( .A(a[680]), .B(n17759), .Z(n361) );
  IV U21176 ( .A(n17757), .Z(n17759) );
  XNOR U21177 ( .A(b[680]), .B(n17757), .Z(n17758) );
  XOR U21178 ( .A(n17760), .B(n17761), .Z(n17757) );
  ANDN U21179 ( .B(n17762), .A(n363), .Z(n17760) );
  XNOR U21180 ( .A(a[679]), .B(n17763), .Z(n363) );
  IV U21181 ( .A(n17761), .Z(n17763) );
  XNOR U21182 ( .A(b[679]), .B(n17761), .Z(n17762) );
  XOR U21183 ( .A(n17764), .B(n17765), .Z(n17761) );
  ANDN U21184 ( .B(n17766), .A(n364), .Z(n17764) );
  XNOR U21185 ( .A(a[678]), .B(n17767), .Z(n364) );
  IV U21186 ( .A(n17765), .Z(n17767) );
  XNOR U21187 ( .A(b[678]), .B(n17765), .Z(n17766) );
  XOR U21188 ( .A(n17768), .B(n17769), .Z(n17765) );
  ANDN U21189 ( .B(n17770), .A(n365), .Z(n17768) );
  XNOR U21190 ( .A(a[677]), .B(n17771), .Z(n365) );
  IV U21191 ( .A(n17769), .Z(n17771) );
  XNOR U21192 ( .A(b[677]), .B(n17769), .Z(n17770) );
  XOR U21193 ( .A(n17772), .B(n17773), .Z(n17769) );
  ANDN U21194 ( .B(n17774), .A(n366), .Z(n17772) );
  XNOR U21195 ( .A(a[676]), .B(n17775), .Z(n366) );
  IV U21196 ( .A(n17773), .Z(n17775) );
  XNOR U21197 ( .A(b[676]), .B(n17773), .Z(n17774) );
  XOR U21198 ( .A(n17776), .B(n17777), .Z(n17773) );
  ANDN U21199 ( .B(n17778), .A(n367), .Z(n17776) );
  XNOR U21200 ( .A(a[675]), .B(n17779), .Z(n367) );
  IV U21201 ( .A(n17777), .Z(n17779) );
  XNOR U21202 ( .A(b[675]), .B(n17777), .Z(n17778) );
  XOR U21203 ( .A(n17780), .B(n17781), .Z(n17777) );
  ANDN U21204 ( .B(n17782), .A(n368), .Z(n17780) );
  XNOR U21205 ( .A(a[674]), .B(n17783), .Z(n368) );
  IV U21206 ( .A(n17781), .Z(n17783) );
  XNOR U21207 ( .A(b[674]), .B(n17781), .Z(n17782) );
  XOR U21208 ( .A(n17784), .B(n17785), .Z(n17781) );
  ANDN U21209 ( .B(n17786), .A(n369), .Z(n17784) );
  XNOR U21210 ( .A(a[673]), .B(n17787), .Z(n369) );
  IV U21211 ( .A(n17785), .Z(n17787) );
  XNOR U21212 ( .A(b[673]), .B(n17785), .Z(n17786) );
  XOR U21213 ( .A(n17788), .B(n17789), .Z(n17785) );
  ANDN U21214 ( .B(n17790), .A(n370), .Z(n17788) );
  XNOR U21215 ( .A(a[672]), .B(n17791), .Z(n370) );
  IV U21216 ( .A(n17789), .Z(n17791) );
  XNOR U21217 ( .A(b[672]), .B(n17789), .Z(n17790) );
  XOR U21218 ( .A(n17792), .B(n17793), .Z(n17789) );
  ANDN U21219 ( .B(n17794), .A(n371), .Z(n17792) );
  XNOR U21220 ( .A(a[671]), .B(n17795), .Z(n371) );
  IV U21221 ( .A(n17793), .Z(n17795) );
  XNOR U21222 ( .A(b[671]), .B(n17793), .Z(n17794) );
  XOR U21223 ( .A(n17796), .B(n17797), .Z(n17793) );
  ANDN U21224 ( .B(n17798), .A(n372), .Z(n17796) );
  XNOR U21225 ( .A(a[670]), .B(n17799), .Z(n372) );
  IV U21226 ( .A(n17797), .Z(n17799) );
  XNOR U21227 ( .A(b[670]), .B(n17797), .Z(n17798) );
  XOR U21228 ( .A(n17800), .B(n17801), .Z(n17797) );
  ANDN U21229 ( .B(n17802), .A(n374), .Z(n17800) );
  XNOR U21230 ( .A(a[669]), .B(n17803), .Z(n374) );
  IV U21231 ( .A(n17801), .Z(n17803) );
  XNOR U21232 ( .A(b[669]), .B(n17801), .Z(n17802) );
  XOR U21233 ( .A(n17804), .B(n17805), .Z(n17801) );
  ANDN U21234 ( .B(n17806), .A(n375), .Z(n17804) );
  XNOR U21235 ( .A(a[668]), .B(n17807), .Z(n375) );
  IV U21236 ( .A(n17805), .Z(n17807) );
  XNOR U21237 ( .A(b[668]), .B(n17805), .Z(n17806) );
  XOR U21238 ( .A(n17808), .B(n17809), .Z(n17805) );
  ANDN U21239 ( .B(n17810), .A(n376), .Z(n17808) );
  XNOR U21240 ( .A(a[667]), .B(n17811), .Z(n376) );
  IV U21241 ( .A(n17809), .Z(n17811) );
  XNOR U21242 ( .A(b[667]), .B(n17809), .Z(n17810) );
  XOR U21243 ( .A(n17812), .B(n17813), .Z(n17809) );
  ANDN U21244 ( .B(n17814), .A(n377), .Z(n17812) );
  XNOR U21245 ( .A(a[666]), .B(n17815), .Z(n377) );
  IV U21246 ( .A(n17813), .Z(n17815) );
  XNOR U21247 ( .A(b[666]), .B(n17813), .Z(n17814) );
  XOR U21248 ( .A(n17816), .B(n17817), .Z(n17813) );
  ANDN U21249 ( .B(n17818), .A(n378), .Z(n17816) );
  XNOR U21250 ( .A(a[665]), .B(n17819), .Z(n378) );
  IV U21251 ( .A(n17817), .Z(n17819) );
  XNOR U21252 ( .A(b[665]), .B(n17817), .Z(n17818) );
  XOR U21253 ( .A(n17820), .B(n17821), .Z(n17817) );
  ANDN U21254 ( .B(n17822), .A(n379), .Z(n17820) );
  XNOR U21255 ( .A(a[664]), .B(n17823), .Z(n379) );
  IV U21256 ( .A(n17821), .Z(n17823) );
  XNOR U21257 ( .A(b[664]), .B(n17821), .Z(n17822) );
  XOR U21258 ( .A(n17824), .B(n17825), .Z(n17821) );
  ANDN U21259 ( .B(n17826), .A(n380), .Z(n17824) );
  XNOR U21260 ( .A(a[663]), .B(n17827), .Z(n380) );
  IV U21261 ( .A(n17825), .Z(n17827) );
  XNOR U21262 ( .A(b[663]), .B(n17825), .Z(n17826) );
  XOR U21263 ( .A(n17828), .B(n17829), .Z(n17825) );
  ANDN U21264 ( .B(n17830), .A(n381), .Z(n17828) );
  XNOR U21265 ( .A(a[662]), .B(n17831), .Z(n381) );
  IV U21266 ( .A(n17829), .Z(n17831) );
  XNOR U21267 ( .A(b[662]), .B(n17829), .Z(n17830) );
  XOR U21268 ( .A(n17832), .B(n17833), .Z(n17829) );
  ANDN U21269 ( .B(n17834), .A(n382), .Z(n17832) );
  XNOR U21270 ( .A(a[661]), .B(n17835), .Z(n382) );
  IV U21271 ( .A(n17833), .Z(n17835) );
  XNOR U21272 ( .A(b[661]), .B(n17833), .Z(n17834) );
  XOR U21273 ( .A(n17836), .B(n17837), .Z(n17833) );
  ANDN U21274 ( .B(n17838), .A(n383), .Z(n17836) );
  XNOR U21275 ( .A(a[660]), .B(n17839), .Z(n383) );
  IV U21276 ( .A(n17837), .Z(n17839) );
  XNOR U21277 ( .A(b[660]), .B(n17837), .Z(n17838) );
  XOR U21278 ( .A(n17840), .B(n17841), .Z(n17837) );
  ANDN U21279 ( .B(n17842), .A(n385), .Z(n17840) );
  XNOR U21280 ( .A(a[659]), .B(n17843), .Z(n385) );
  IV U21281 ( .A(n17841), .Z(n17843) );
  XNOR U21282 ( .A(b[659]), .B(n17841), .Z(n17842) );
  XOR U21283 ( .A(n17844), .B(n17845), .Z(n17841) );
  ANDN U21284 ( .B(n17846), .A(n386), .Z(n17844) );
  XNOR U21285 ( .A(a[658]), .B(n17847), .Z(n386) );
  IV U21286 ( .A(n17845), .Z(n17847) );
  XNOR U21287 ( .A(b[658]), .B(n17845), .Z(n17846) );
  XOR U21288 ( .A(n17848), .B(n17849), .Z(n17845) );
  ANDN U21289 ( .B(n17850), .A(n387), .Z(n17848) );
  XNOR U21290 ( .A(a[657]), .B(n17851), .Z(n387) );
  IV U21291 ( .A(n17849), .Z(n17851) );
  XNOR U21292 ( .A(b[657]), .B(n17849), .Z(n17850) );
  XOR U21293 ( .A(n17852), .B(n17853), .Z(n17849) );
  ANDN U21294 ( .B(n17854), .A(n388), .Z(n17852) );
  XNOR U21295 ( .A(a[656]), .B(n17855), .Z(n388) );
  IV U21296 ( .A(n17853), .Z(n17855) );
  XNOR U21297 ( .A(b[656]), .B(n17853), .Z(n17854) );
  XOR U21298 ( .A(n17856), .B(n17857), .Z(n17853) );
  ANDN U21299 ( .B(n17858), .A(n389), .Z(n17856) );
  XNOR U21300 ( .A(a[655]), .B(n17859), .Z(n389) );
  IV U21301 ( .A(n17857), .Z(n17859) );
  XNOR U21302 ( .A(b[655]), .B(n17857), .Z(n17858) );
  XOR U21303 ( .A(n17860), .B(n17861), .Z(n17857) );
  ANDN U21304 ( .B(n17862), .A(n390), .Z(n17860) );
  XNOR U21305 ( .A(a[654]), .B(n17863), .Z(n390) );
  IV U21306 ( .A(n17861), .Z(n17863) );
  XNOR U21307 ( .A(b[654]), .B(n17861), .Z(n17862) );
  XOR U21308 ( .A(n17864), .B(n17865), .Z(n17861) );
  ANDN U21309 ( .B(n17866), .A(n391), .Z(n17864) );
  XNOR U21310 ( .A(a[653]), .B(n17867), .Z(n391) );
  IV U21311 ( .A(n17865), .Z(n17867) );
  XNOR U21312 ( .A(b[653]), .B(n17865), .Z(n17866) );
  XOR U21313 ( .A(n17868), .B(n17869), .Z(n17865) );
  ANDN U21314 ( .B(n17870), .A(n392), .Z(n17868) );
  XNOR U21315 ( .A(a[652]), .B(n17871), .Z(n392) );
  IV U21316 ( .A(n17869), .Z(n17871) );
  XNOR U21317 ( .A(b[652]), .B(n17869), .Z(n17870) );
  XOR U21318 ( .A(n17872), .B(n17873), .Z(n17869) );
  ANDN U21319 ( .B(n17874), .A(n393), .Z(n17872) );
  XNOR U21320 ( .A(a[651]), .B(n17875), .Z(n393) );
  IV U21321 ( .A(n17873), .Z(n17875) );
  XNOR U21322 ( .A(b[651]), .B(n17873), .Z(n17874) );
  XOR U21323 ( .A(n17876), .B(n17877), .Z(n17873) );
  ANDN U21324 ( .B(n17878), .A(n394), .Z(n17876) );
  XNOR U21325 ( .A(a[650]), .B(n17879), .Z(n394) );
  IV U21326 ( .A(n17877), .Z(n17879) );
  XNOR U21327 ( .A(b[650]), .B(n17877), .Z(n17878) );
  XOR U21328 ( .A(n17880), .B(n17881), .Z(n17877) );
  ANDN U21329 ( .B(n17882), .A(n396), .Z(n17880) );
  XNOR U21330 ( .A(a[649]), .B(n17883), .Z(n396) );
  IV U21331 ( .A(n17881), .Z(n17883) );
  XNOR U21332 ( .A(b[649]), .B(n17881), .Z(n17882) );
  XOR U21333 ( .A(n17884), .B(n17885), .Z(n17881) );
  ANDN U21334 ( .B(n17886), .A(n397), .Z(n17884) );
  XNOR U21335 ( .A(a[648]), .B(n17887), .Z(n397) );
  IV U21336 ( .A(n17885), .Z(n17887) );
  XNOR U21337 ( .A(b[648]), .B(n17885), .Z(n17886) );
  XOR U21338 ( .A(n17888), .B(n17889), .Z(n17885) );
  ANDN U21339 ( .B(n17890), .A(n398), .Z(n17888) );
  XNOR U21340 ( .A(a[647]), .B(n17891), .Z(n398) );
  IV U21341 ( .A(n17889), .Z(n17891) );
  XNOR U21342 ( .A(b[647]), .B(n17889), .Z(n17890) );
  XOR U21343 ( .A(n17892), .B(n17893), .Z(n17889) );
  ANDN U21344 ( .B(n17894), .A(n399), .Z(n17892) );
  XNOR U21345 ( .A(a[646]), .B(n17895), .Z(n399) );
  IV U21346 ( .A(n17893), .Z(n17895) );
  XNOR U21347 ( .A(b[646]), .B(n17893), .Z(n17894) );
  XOR U21348 ( .A(n17896), .B(n17897), .Z(n17893) );
  ANDN U21349 ( .B(n17898), .A(n400), .Z(n17896) );
  XNOR U21350 ( .A(a[645]), .B(n17899), .Z(n400) );
  IV U21351 ( .A(n17897), .Z(n17899) );
  XNOR U21352 ( .A(b[645]), .B(n17897), .Z(n17898) );
  XOR U21353 ( .A(n17900), .B(n17901), .Z(n17897) );
  ANDN U21354 ( .B(n17902), .A(n401), .Z(n17900) );
  XNOR U21355 ( .A(a[644]), .B(n17903), .Z(n401) );
  IV U21356 ( .A(n17901), .Z(n17903) );
  XNOR U21357 ( .A(b[644]), .B(n17901), .Z(n17902) );
  XOR U21358 ( .A(n17904), .B(n17905), .Z(n17901) );
  ANDN U21359 ( .B(n17906), .A(n402), .Z(n17904) );
  XNOR U21360 ( .A(a[643]), .B(n17907), .Z(n402) );
  IV U21361 ( .A(n17905), .Z(n17907) );
  XNOR U21362 ( .A(b[643]), .B(n17905), .Z(n17906) );
  XOR U21363 ( .A(n17908), .B(n17909), .Z(n17905) );
  ANDN U21364 ( .B(n17910), .A(n403), .Z(n17908) );
  XNOR U21365 ( .A(a[642]), .B(n17911), .Z(n403) );
  IV U21366 ( .A(n17909), .Z(n17911) );
  XNOR U21367 ( .A(b[642]), .B(n17909), .Z(n17910) );
  XOR U21368 ( .A(n17912), .B(n17913), .Z(n17909) );
  ANDN U21369 ( .B(n17914), .A(n404), .Z(n17912) );
  XNOR U21370 ( .A(a[641]), .B(n17915), .Z(n404) );
  IV U21371 ( .A(n17913), .Z(n17915) );
  XNOR U21372 ( .A(b[641]), .B(n17913), .Z(n17914) );
  XOR U21373 ( .A(n17916), .B(n17917), .Z(n17913) );
  ANDN U21374 ( .B(n17918), .A(n405), .Z(n17916) );
  XNOR U21375 ( .A(a[640]), .B(n17919), .Z(n405) );
  IV U21376 ( .A(n17917), .Z(n17919) );
  XNOR U21377 ( .A(b[640]), .B(n17917), .Z(n17918) );
  XOR U21378 ( .A(n17920), .B(n17921), .Z(n17917) );
  ANDN U21379 ( .B(n17922), .A(n407), .Z(n17920) );
  XNOR U21380 ( .A(a[639]), .B(n17923), .Z(n407) );
  IV U21381 ( .A(n17921), .Z(n17923) );
  XNOR U21382 ( .A(b[639]), .B(n17921), .Z(n17922) );
  XOR U21383 ( .A(n17924), .B(n17925), .Z(n17921) );
  ANDN U21384 ( .B(n17926), .A(n408), .Z(n17924) );
  XNOR U21385 ( .A(a[638]), .B(n17927), .Z(n408) );
  IV U21386 ( .A(n17925), .Z(n17927) );
  XNOR U21387 ( .A(b[638]), .B(n17925), .Z(n17926) );
  XOR U21388 ( .A(n17928), .B(n17929), .Z(n17925) );
  ANDN U21389 ( .B(n17930), .A(n409), .Z(n17928) );
  XNOR U21390 ( .A(a[637]), .B(n17931), .Z(n409) );
  IV U21391 ( .A(n17929), .Z(n17931) );
  XNOR U21392 ( .A(b[637]), .B(n17929), .Z(n17930) );
  XOR U21393 ( .A(n17932), .B(n17933), .Z(n17929) );
  ANDN U21394 ( .B(n17934), .A(n410), .Z(n17932) );
  XNOR U21395 ( .A(a[636]), .B(n17935), .Z(n410) );
  IV U21396 ( .A(n17933), .Z(n17935) );
  XNOR U21397 ( .A(b[636]), .B(n17933), .Z(n17934) );
  XOR U21398 ( .A(n17936), .B(n17937), .Z(n17933) );
  ANDN U21399 ( .B(n17938), .A(n411), .Z(n17936) );
  XNOR U21400 ( .A(a[635]), .B(n17939), .Z(n411) );
  IV U21401 ( .A(n17937), .Z(n17939) );
  XNOR U21402 ( .A(b[635]), .B(n17937), .Z(n17938) );
  XOR U21403 ( .A(n17940), .B(n17941), .Z(n17937) );
  ANDN U21404 ( .B(n17942), .A(n412), .Z(n17940) );
  XNOR U21405 ( .A(a[634]), .B(n17943), .Z(n412) );
  IV U21406 ( .A(n17941), .Z(n17943) );
  XNOR U21407 ( .A(b[634]), .B(n17941), .Z(n17942) );
  XOR U21408 ( .A(n17944), .B(n17945), .Z(n17941) );
  ANDN U21409 ( .B(n17946), .A(n413), .Z(n17944) );
  XNOR U21410 ( .A(a[633]), .B(n17947), .Z(n413) );
  IV U21411 ( .A(n17945), .Z(n17947) );
  XNOR U21412 ( .A(b[633]), .B(n17945), .Z(n17946) );
  XOR U21413 ( .A(n17948), .B(n17949), .Z(n17945) );
  ANDN U21414 ( .B(n17950), .A(n414), .Z(n17948) );
  XNOR U21415 ( .A(a[632]), .B(n17951), .Z(n414) );
  IV U21416 ( .A(n17949), .Z(n17951) );
  XNOR U21417 ( .A(b[632]), .B(n17949), .Z(n17950) );
  XOR U21418 ( .A(n17952), .B(n17953), .Z(n17949) );
  ANDN U21419 ( .B(n17954), .A(n415), .Z(n17952) );
  XNOR U21420 ( .A(a[631]), .B(n17955), .Z(n415) );
  IV U21421 ( .A(n17953), .Z(n17955) );
  XNOR U21422 ( .A(b[631]), .B(n17953), .Z(n17954) );
  XOR U21423 ( .A(n17956), .B(n17957), .Z(n17953) );
  ANDN U21424 ( .B(n17958), .A(n416), .Z(n17956) );
  XNOR U21425 ( .A(a[630]), .B(n17959), .Z(n416) );
  IV U21426 ( .A(n17957), .Z(n17959) );
  XNOR U21427 ( .A(b[630]), .B(n17957), .Z(n17958) );
  XOR U21428 ( .A(n17960), .B(n17961), .Z(n17957) );
  ANDN U21429 ( .B(n17962), .A(n418), .Z(n17960) );
  XNOR U21430 ( .A(a[629]), .B(n17963), .Z(n418) );
  IV U21431 ( .A(n17961), .Z(n17963) );
  XNOR U21432 ( .A(b[629]), .B(n17961), .Z(n17962) );
  XOR U21433 ( .A(n17964), .B(n17965), .Z(n17961) );
  ANDN U21434 ( .B(n17966), .A(n419), .Z(n17964) );
  XNOR U21435 ( .A(a[628]), .B(n17967), .Z(n419) );
  IV U21436 ( .A(n17965), .Z(n17967) );
  XNOR U21437 ( .A(b[628]), .B(n17965), .Z(n17966) );
  XOR U21438 ( .A(n17968), .B(n17969), .Z(n17965) );
  ANDN U21439 ( .B(n17970), .A(n420), .Z(n17968) );
  XNOR U21440 ( .A(a[627]), .B(n17971), .Z(n420) );
  IV U21441 ( .A(n17969), .Z(n17971) );
  XNOR U21442 ( .A(b[627]), .B(n17969), .Z(n17970) );
  XOR U21443 ( .A(n17972), .B(n17973), .Z(n17969) );
  ANDN U21444 ( .B(n17974), .A(n421), .Z(n17972) );
  XNOR U21445 ( .A(a[626]), .B(n17975), .Z(n421) );
  IV U21446 ( .A(n17973), .Z(n17975) );
  XNOR U21447 ( .A(b[626]), .B(n17973), .Z(n17974) );
  XOR U21448 ( .A(n17976), .B(n17977), .Z(n17973) );
  ANDN U21449 ( .B(n17978), .A(n422), .Z(n17976) );
  XNOR U21450 ( .A(a[625]), .B(n17979), .Z(n422) );
  IV U21451 ( .A(n17977), .Z(n17979) );
  XNOR U21452 ( .A(b[625]), .B(n17977), .Z(n17978) );
  XOR U21453 ( .A(n17980), .B(n17981), .Z(n17977) );
  ANDN U21454 ( .B(n17982), .A(n423), .Z(n17980) );
  XNOR U21455 ( .A(a[624]), .B(n17983), .Z(n423) );
  IV U21456 ( .A(n17981), .Z(n17983) );
  XNOR U21457 ( .A(b[624]), .B(n17981), .Z(n17982) );
  XOR U21458 ( .A(n17984), .B(n17985), .Z(n17981) );
  ANDN U21459 ( .B(n17986), .A(n424), .Z(n17984) );
  XNOR U21460 ( .A(a[623]), .B(n17987), .Z(n424) );
  IV U21461 ( .A(n17985), .Z(n17987) );
  XNOR U21462 ( .A(b[623]), .B(n17985), .Z(n17986) );
  XOR U21463 ( .A(n17988), .B(n17989), .Z(n17985) );
  ANDN U21464 ( .B(n17990), .A(n425), .Z(n17988) );
  XNOR U21465 ( .A(a[622]), .B(n17991), .Z(n425) );
  IV U21466 ( .A(n17989), .Z(n17991) );
  XNOR U21467 ( .A(b[622]), .B(n17989), .Z(n17990) );
  XOR U21468 ( .A(n17992), .B(n17993), .Z(n17989) );
  ANDN U21469 ( .B(n17994), .A(n426), .Z(n17992) );
  XNOR U21470 ( .A(a[621]), .B(n17995), .Z(n426) );
  IV U21471 ( .A(n17993), .Z(n17995) );
  XNOR U21472 ( .A(b[621]), .B(n17993), .Z(n17994) );
  XOR U21473 ( .A(n17996), .B(n17997), .Z(n17993) );
  ANDN U21474 ( .B(n17998), .A(n427), .Z(n17996) );
  XNOR U21475 ( .A(a[620]), .B(n17999), .Z(n427) );
  IV U21476 ( .A(n17997), .Z(n17999) );
  XNOR U21477 ( .A(b[620]), .B(n17997), .Z(n17998) );
  XOR U21478 ( .A(n18000), .B(n18001), .Z(n17997) );
  ANDN U21479 ( .B(n18002), .A(n429), .Z(n18000) );
  XNOR U21480 ( .A(a[619]), .B(n18003), .Z(n429) );
  IV U21481 ( .A(n18001), .Z(n18003) );
  XNOR U21482 ( .A(b[619]), .B(n18001), .Z(n18002) );
  XOR U21483 ( .A(n18004), .B(n18005), .Z(n18001) );
  ANDN U21484 ( .B(n18006), .A(n430), .Z(n18004) );
  XNOR U21485 ( .A(a[618]), .B(n18007), .Z(n430) );
  IV U21486 ( .A(n18005), .Z(n18007) );
  XNOR U21487 ( .A(b[618]), .B(n18005), .Z(n18006) );
  XOR U21488 ( .A(n18008), .B(n18009), .Z(n18005) );
  ANDN U21489 ( .B(n18010), .A(n431), .Z(n18008) );
  XNOR U21490 ( .A(a[617]), .B(n18011), .Z(n431) );
  IV U21491 ( .A(n18009), .Z(n18011) );
  XNOR U21492 ( .A(b[617]), .B(n18009), .Z(n18010) );
  XOR U21493 ( .A(n18012), .B(n18013), .Z(n18009) );
  ANDN U21494 ( .B(n18014), .A(n432), .Z(n18012) );
  XNOR U21495 ( .A(a[616]), .B(n18015), .Z(n432) );
  IV U21496 ( .A(n18013), .Z(n18015) );
  XNOR U21497 ( .A(b[616]), .B(n18013), .Z(n18014) );
  XOR U21498 ( .A(n18016), .B(n18017), .Z(n18013) );
  ANDN U21499 ( .B(n18018), .A(n433), .Z(n18016) );
  XNOR U21500 ( .A(a[615]), .B(n18019), .Z(n433) );
  IV U21501 ( .A(n18017), .Z(n18019) );
  XNOR U21502 ( .A(b[615]), .B(n18017), .Z(n18018) );
  XOR U21503 ( .A(n18020), .B(n18021), .Z(n18017) );
  ANDN U21504 ( .B(n18022), .A(n434), .Z(n18020) );
  XNOR U21505 ( .A(a[614]), .B(n18023), .Z(n434) );
  IV U21506 ( .A(n18021), .Z(n18023) );
  XNOR U21507 ( .A(b[614]), .B(n18021), .Z(n18022) );
  XOR U21508 ( .A(n18024), .B(n18025), .Z(n18021) );
  ANDN U21509 ( .B(n18026), .A(n435), .Z(n18024) );
  XNOR U21510 ( .A(a[613]), .B(n18027), .Z(n435) );
  IV U21511 ( .A(n18025), .Z(n18027) );
  XNOR U21512 ( .A(b[613]), .B(n18025), .Z(n18026) );
  XOR U21513 ( .A(n18028), .B(n18029), .Z(n18025) );
  ANDN U21514 ( .B(n18030), .A(n436), .Z(n18028) );
  XNOR U21515 ( .A(a[612]), .B(n18031), .Z(n436) );
  IV U21516 ( .A(n18029), .Z(n18031) );
  XNOR U21517 ( .A(b[612]), .B(n18029), .Z(n18030) );
  XOR U21518 ( .A(n18032), .B(n18033), .Z(n18029) );
  ANDN U21519 ( .B(n18034), .A(n437), .Z(n18032) );
  XNOR U21520 ( .A(a[611]), .B(n18035), .Z(n437) );
  IV U21521 ( .A(n18033), .Z(n18035) );
  XNOR U21522 ( .A(b[611]), .B(n18033), .Z(n18034) );
  XOR U21523 ( .A(n18036), .B(n18037), .Z(n18033) );
  ANDN U21524 ( .B(n18038), .A(n438), .Z(n18036) );
  XNOR U21525 ( .A(a[610]), .B(n18039), .Z(n438) );
  IV U21526 ( .A(n18037), .Z(n18039) );
  XNOR U21527 ( .A(b[610]), .B(n18037), .Z(n18038) );
  XOR U21528 ( .A(n18040), .B(n18041), .Z(n18037) );
  ANDN U21529 ( .B(n18042), .A(n440), .Z(n18040) );
  XNOR U21530 ( .A(a[609]), .B(n18043), .Z(n440) );
  IV U21531 ( .A(n18041), .Z(n18043) );
  XNOR U21532 ( .A(b[609]), .B(n18041), .Z(n18042) );
  XOR U21533 ( .A(n18044), .B(n18045), .Z(n18041) );
  ANDN U21534 ( .B(n18046), .A(n441), .Z(n18044) );
  XNOR U21535 ( .A(a[608]), .B(n18047), .Z(n441) );
  IV U21536 ( .A(n18045), .Z(n18047) );
  XNOR U21537 ( .A(b[608]), .B(n18045), .Z(n18046) );
  XOR U21538 ( .A(n18048), .B(n18049), .Z(n18045) );
  ANDN U21539 ( .B(n18050), .A(n442), .Z(n18048) );
  XNOR U21540 ( .A(a[607]), .B(n18051), .Z(n442) );
  IV U21541 ( .A(n18049), .Z(n18051) );
  XNOR U21542 ( .A(b[607]), .B(n18049), .Z(n18050) );
  XOR U21543 ( .A(n18052), .B(n18053), .Z(n18049) );
  ANDN U21544 ( .B(n18054), .A(n443), .Z(n18052) );
  XNOR U21545 ( .A(a[606]), .B(n18055), .Z(n443) );
  IV U21546 ( .A(n18053), .Z(n18055) );
  XNOR U21547 ( .A(b[606]), .B(n18053), .Z(n18054) );
  XOR U21548 ( .A(n18056), .B(n18057), .Z(n18053) );
  ANDN U21549 ( .B(n18058), .A(n444), .Z(n18056) );
  XNOR U21550 ( .A(a[605]), .B(n18059), .Z(n444) );
  IV U21551 ( .A(n18057), .Z(n18059) );
  XNOR U21552 ( .A(b[605]), .B(n18057), .Z(n18058) );
  XOR U21553 ( .A(n18060), .B(n18061), .Z(n18057) );
  ANDN U21554 ( .B(n18062), .A(n445), .Z(n18060) );
  XNOR U21555 ( .A(a[604]), .B(n18063), .Z(n445) );
  IV U21556 ( .A(n18061), .Z(n18063) );
  XNOR U21557 ( .A(b[604]), .B(n18061), .Z(n18062) );
  XOR U21558 ( .A(n18064), .B(n18065), .Z(n18061) );
  ANDN U21559 ( .B(n18066), .A(n446), .Z(n18064) );
  XNOR U21560 ( .A(a[603]), .B(n18067), .Z(n446) );
  IV U21561 ( .A(n18065), .Z(n18067) );
  XNOR U21562 ( .A(b[603]), .B(n18065), .Z(n18066) );
  XOR U21563 ( .A(n18068), .B(n18069), .Z(n18065) );
  ANDN U21564 ( .B(n18070), .A(n447), .Z(n18068) );
  XNOR U21565 ( .A(a[602]), .B(n18071), .Z(n447) );
  IV U21566 ( .A(n18069), .Z(n18071) );
  XNOR U21567 ( .A(b[602]), .B(n18069), .Z(n18070) );
  XOR U21568 ( .A(n18072), .B(n18073), .Z(n18069) );
  ANDN U21569 ( .B(n18074), .A(n448), .Z(n18072) );
  XNOR U21570 ( .A(a[601]), .B(n18075), .Z(n448) );
  IV U21571 ( .A(n18073), .Z(n18075) );
  XNOR U21572 ( .A(b[601]), .B(n18073), .Z(n18074) );
  XOR U21573 ( .A(n18076), .B(n18077), .Z(n18073) );
  ANDN U21574 ( .B(n18078), .A(n449), .Z(n18076) );
  XNOR U21575 ( .A(a[600]), .B(n18079), .Z(n449) );
  IV U21576 ( .A(n18077), .Z(n18079) );
  XNOR U21577 ( .A(b[600]), .B(n18077), .Z(n18078) );
  XOR U21578 ( .A(n18080), .B(n18081), .Z(n18077) );
  ANDN U21579 ( .B(n18082), .A(n452), .Z(n18080) );
  XNOR U21580 ( .A(a[599]), .B(n18083), .Z(n452) );
  IV U21581 ( .A(n18081), .Z(n18083) );
  XNOR U21582 ( .A(b[599]), .B(n18081), .Z(n18082) );
  XOR U21583 ( .A(n18084), .B(n18085), .Z(n18081) );
  ANDN U21584 ( .B(n18086), .A(n453), .Z(n18084) );
  XNOR U21585 ( .A(a[598]), .B(n18087), .Z(n453) );
  IV U21586 ( .A(n18085), .Z(n18087) );
  XNOR U21587 ( .A(b[598]), .B(n18085), .Z(n18086) );
  XOR U21588 ( .A(n18088), .B(n18089), .Z(n18085) );
  ANDN U21589 ( .B(n18090), .A(n454), .Z(n18088) );
  XNOR U21590 ( .A(a[597]), .B(n18091), .Z(n454) );
  IV U21591 ( .A(n18089), .Z(n18091) );
  XNOR U21592 ( .A(b[597]), .B(n18089), .Z(n18090) );
  XOR U21593 ( .A(n18092), .B(n18093), .Z(n18089) );
  ANDN U21594 ( .B(n18094), .A(n455), .Z(n18092) );
  XNOR U21595 ( .A(a[596]), .B(n18095), .Z(n455) );
  IV U21596 ( .A(n18093), .Z(n18095) );
  XNOR U21597 ( .A(b[596]), .B(n18093), .Z(n18094) );
  XOR U21598 ( .A(n18096), .B(n18097), .Z(n18093) );
  ANDN U21599 ( .B(n18098), .A(n456), .Z(n18096) );
  XNOR U21600 ( .A(a[595]), .B(n18099), .Z(n456) );
  IV U21601 ( .A(n18097), .Z(n18099) );
  XNOR U21602 ( .A(b[595]), .B(n18097), .Z(n18098) );
  XOR U21603 ( .A(n18100), .B(n18101), .Z(n18097) );
  ANDN U21604 ( .B(n18102), .A(n457), .Z(n18100) );
  XNOR U21605 ( .A(a[594]), .B(n18103), .Z(n457) );
  IV U21606 ( .A(n18101), .Z(n18103) );
  XNOR U21607 ( .A(b[594]), .B(n18101), .Z(n18102) );
  XOR U21608 ( .A(n18104), .B(n18105), .Z(n18101) );
  ANDN U21609 ( .B(n18106), .A(n458), .Z(n18104) );
  XNOR U21610 ( .A(a[593]), .B(n18107), .Z(n458) );
  IV U21611 ( .A(n18105), .Z(n18107) );
  XNOR U21612 ( .A(b[593]), .B(n18105), .Z(n18106) );
  XOR U21613 ( .A(n18108), .B(n18109), .Z(n18105) );
  ANDN U21614 ( .B(n18110), .A(n459), .Z(n18108) );
  XNOR U21615 ( .A(a[592]), .B(n18111), .Z(n459) );
  IV U21616 ( .A(n18109), .Z(n18111) );
  XNOR U21617 ( .A(b[592]), .B(n18109), .Z(n18110) );
  XOR U21618 ( .A(n18112), .B(n18113), .Z(n18109) );
  ANDN U21619 ( .B(n18114), .A(n460), .Z(n18112) );
  XNOR U21620 ( .A(a[591]), .B(n18115), .Z(n460) );
  IV U21621 ( .A(n18113), .Z(n18115) );
  XNOR U21622 ( .A(b[591]), .B(n18113), .Z(n18114) );
  XOR U21623 ( .A(n18116), .B(n18117), .Z(n18113) );
  ANDN U21624 ( .B(n18118), .A(n461), .Z(n18116) );
  XNOR U21625 ( .A(a[590]), .B(n18119), .Z(n461) );
  IV U21626 ( .A(n18117), .Z(n18119) );
  XNOR U21627 ( .A(b[590]), .B(n18117), .Z(n18118) );
  XOR U21628 ( .A(n18120), .B(n18121), .Z(n18117) );
  ANDN U21629 ( .B(n18122), .A(n463), .Z(n18120) );
  XNOR U21630 ( .A(a[589]), .B(n18123), .Z(n463) );
  IV U21631 ( .A(n18121), .Z(n18123) );
  XNOR U21632 ( .A(b[589]), .B(n18121), .Z(n18122) );
  XOR U21633 ( .A(n18124), .B(n18125), .Z(n18121) );
  ANDN U21634 ( .B(n18126), .A(n464), .Z(n18124) );
  XNOR U21635 ( .A(a[588]), .B(n18127), .Z(n464) );
  IV U21636 ( .A(n18125), .Z(n18127) );
  XNOR U21637 ( .A(b[588]), .B(n18125), .Z(n18126) );
  XOR U21638 ( .A(n18128), .B(n18129), .Z(n18125) );
  ANDN U21639 ( .B(n18130), .A(n465), .Z(n18128) );
  XNOR U21640 ( .A(a[587]), .B(n18131), .Z(n465) );
  IV U21641 ( .A(n18129), .Z(n18131) );
  XNOR U21642 ( .A(b[587]), .B(n18129), .Z(n18130) );
  XOR U21643 ( .A(n18132), .B(n18133), .Z(n18129) );
  ANDN U21644 ( .B(n18134), .A(n466), .Z(n18132) );
  XNOR U21645 ( .A(a[586]), .B(n18135), .Z(n466) );
  IV U21646 ( .A(n18133), .Z(n18135) );
  XNOR U21647 ( .A(b[586]), .B(n18133), .Z(n18134) );
  XOR U21648 ( .A(n18136), .B(n18137), .Z(n18133) );
  ANDN U21649 ( .B(n18138), .A(n467), .Z(n18136) );
  XNOR U21650 ( .A(a[585]), .B(n18139), .Z(n467) );
  IV U21651 ( .A(n18137), .Z(n18139) );
  XNOR U21652 ( .A(b[585]), .B(n18137), .Z(n18138) );
  XOR U21653 ( .A(n18140), .B(n18141), .Z(n18137) );
  ANDN U21654 ( .B(n18142), .A(n468), .Z(n18140) );
  XNOR U21655 ( .A(a[584]), .B(n18143), .Z(n468) );
  IV U21656 ( .A(n18141), .Z(n18143) );
  XNOR U21657 ( .A(b[584]), .B(n18141), .Z(n18142) );
  XOR U21658 ( .A(n18144), .B(n18145), .Z(n18141) );
  ANDN U21659 ( .B(n18146), .A(n469), .Z(n18144) );
  XNOR U21660 ( .A(a[583]), .B(n18147), .Z(n469) );
  IV U21661 ( .A(n18145), .Z(n18147) );
  XNOR U21662 ( .A(b[583]), .B(n18145), .Z(n18146) );
  XOR U21663 ( .A(n18148), .B(n18149), .Z(n18145) );
  ANDN U21664 ( .B(n18150), .A(n470), .Z(n18148) );
  XNOR U21665 ( .A(a[582]), .B(n18151), .Z(n470) );
  IV U21666 ( .A(n18149), .Z(n18151) );
  XNOR U21667 ( .A(b[582]), .B(n18149), .Z(n18150) );
  XOR U21668 ( .A(n18152), .B(n18153), .Z(n18149) );
  ANDN U21669 ( .B(n18154), .A(n471), .Z(n18152) );
  XNOR U21670 ( .A(a[581]), .B(n18155), .Z(n471) );
  IV U21671 ( .A(n18153), .Z(n18155) );
  XNOR U21672 ( .A(b[581]), .B(n18153), .Z(n18154) );
  XOR U21673 ( .A(n18156), .B(n18157), .Z(n18153) );
  ANDN U21674 ( .B(n18158), .A(n472), .Z(n18156) );
  XNOR U21675 ( .A(a[580]), .B(n18159), .Z(n472) );
  IV U21676 ( .A(n18157), .Z(n18159) );
  XNOR U21677 ( .A(b[580]), .B(n18157), .Z(n18158) );
  XOR U21678 ( .A(n18160), .B(n18161), .Z(n18157) );
  ANDN U21679 ( .B(n18162), .A(n474), .Z(n18160) );
  XNOR U21680 ( .A(a[579]), .B(n18163), .Z(n474) );
  IV U21681 ( .A(n18161), .Z(n18163) );
  XNOR U21682 ( .A(b[579]), .B(n18161), .Z(n18162) );
  XOR U21683 ( .A(n18164), .B(n18165), .Z(n18161) );
  ANDN U21684 ( .B(n18166), .A(n475), .Z(n18164) );
  XNOR U21685 ( .A(a[578]), .B(n18167), .Z(n475) );
  IV U21686 ( .A(n18165), .Z(n18167) );
  XNOR U21687 ( .A(b[578]), .B(n18165), .Z(n18166) );
  XOR U21688 ( .A(n18168), .B(n18169), .Z(n18165) );
  ANDN U21689 ( .B(n18170), .A(n476), .Z(n18168) );
  XNOR U21690 ( .A(a[577]), .B(n18171), .Z(n476) );
  IV U21691 ( .A(n18169), .Z(n18171) );
  XNOR U21692 ( .A(b[577]), .B(n18169), .Z(n18170) );
  XOR U21693 ( .A(n18172), .B(n18173), .Z(n18169) );
  ANDN U21694 ( .B(n18174), .A(n477), .Z(n18172) );
  XNOR U21695 ( .A(a[576]), .B(n18175), .Z(n477) );
  IV U21696 ( .A(n18173), .Z(n18175) );
  XNOR U21697 ( .A(b[576]), .B(n18173), .Z(n18174) );
  XOR U21698 ( .A(n18176), .B(n18177), .Z(n18173) );
  ANDN U21699 ( .B(n18178), .A(n478), .Z(n18176) );
  XNOR U21700 ( .A(a[575]), .B(n18179), .Z(n478) );
  IV U21701 ( .A(n18177), .Z(n18179) );
  XNOR U21702 ( .A(b[575]), .B(n18177), .Z(n18178) );
  XOR U21703 ( .A(n18180), .B(n18181), .Z(n18177) );
  ANDN U21704 ( .B(n18182), .A(n479), .Z(n18180) );
  XNOR U21705 ( .A(a[574]), .B(n18183), .Z(n479) );
  IV U21706 ( .A(n18181), .Z(n18183) );
  XNOR U21707 ( .A(b[574]), .B(n18181), .Z(n18182) );
  XOR U21708 ( .A(n18184), .B(n18185), .Z(n18181) );
  ANDN U21709 ( .B(n18186), .A(n480), .Z(n18184) );
  XNOR U21710 ( .A(a[573]), .B(n18187), .Z(n480) );
  IV U21711 ( .A(n18185), .Z(n18187) );
  XNOR U21712 ( .A(b[573]), .B(n18185), .Z(n18186) );
  XOR U21713 ( .A(n18188), .B(n18189), .Z(n18185) );
  ANDN U21714 ( .B(n18190), .A(n481), .Z(n18188) );
  XNOR U21715 ( .A(a[572]), .B(n18191), .Z(n481) );
  IV U21716 ( .A(n18189), .Z(n18191) );
  XNOR U21717 ( .A(b[572]), .B(n18189), .Z(n18190) );
  XOR U21718 ( .A(n18192), .B(n18193), .Z(n18189) );
  ANDN U21719 ( .B(n18194), .A(n482), .Z(n18192) );
  XNOR U21720 ( .A(a[571]), .B(n18195), .Z(n482) );
  IV U21721 ( .A(n18193), .Z(n18195) );
  XNOR U21722 ( .A(b[571]), .B(n18193), .Z(n18194) );
  XOR U21723 ( .A(n18196), .B(n18197), .Z(n18193) );
  ANDN U21724 ( .B(n18198), .A(n483), .Z(n18196) );
  XNOR U21725 ( .A(a[570]), .B(n18199), .Z(n483) );
  IV U21726 ( .A(n18197), .Z(n18199) );
  XNOR U21727 ( .A(b[570]), .B(n18197), .Z(n18198) );
  XOR U21728 ( .A(n18200), .B(n18201), .Z(n18197) );
  ANDN U21729 ( .B(n18202), .A(n485), .Z(n18200) );
  XNOR U21730 ( .A(a[569]), .B(n18203), .Z(n485) );
  IV U21731 ( .A(n18201), .Z(n18203) );
  XNOR U21732 ( .A(b[569]), .B(n18201), .Z(n18202) );
  XOR U21733 ( .A(n18204), .B(n18205), .Z(n18201) );
  ANDN U21734 ( .B(n18206), .A(n486), .Z(n18204) );
  XNOR U21735 ( .A(a[568]), .B(n18207), .Z(n486) );
  IV U21736 ( .A(n18205), .Z(n18207) );
  XNOR U21737 ( .A(b[568]), .B(n18205), .Z(n18206) );
  XOR U21738 ( .A(n18208), .B(n18209), .Z(n18205) );
  ANDN U21739 ( .B(n18210), .A(n487), .Z(n18208) );
  XNOR U21740 ( .A(a[567]), .B(n18211), .Z(n487) );
  IV U21741 ( .A(n18209), .Z(n18211) );
  XNOR U21742 ( .A(b[567]), .B(n18209), .Z(n18210) );
  XOR U21743 ( .A(n18212), .B(n18213), .Z(n18209) );
  ANDN U21744 ( .B(n18214), .A(n488), .Z(n18212) );
  XNOR U21745 ( .A(a[566]), .B(n18215), .Z(n488) );
  IV U21746 ( .A(n18213), .Z(n18215) );
  XNOR U21747 ( .A(b[566]), .B(n18213), .Z(n18214) );
  XOR U21748 ( .A(n18216), .B(n18217), .Z(n18213) );
  ANDN U21749 ( .B(n18218), .A(n489), .Z(n18216) );
  XNOR U21750 ( .A(a[565]), .B(n18219), .Z(n489) );
  IV U21751 ( .A(n18217), .Z(n18219) );
  XNOR U21752 ( .A(b[565]), .B(n18217), .Z(n18218) );
  XOR U21753 ( .A(n18220), .B(n18221), .Z(n18217) );
  ANDN U21754 ( .B(n18222), .A(n490), .Z(n18220) );
  XNOR U21755 ( .A(a[564]), .B(n18223), .Z(n490) );
  IV U21756 ( .A(n18221), .Z(n18223) );
  XNOR U21757 ( .A(b[564]), .B(n18221), .Z(n18222) );
  XOR U21758 ( .A(n18224), .B(n18225), .Z(n18221) );
  ANDN U21759 ( .B(n18226), .A(n491), .Z(n18224) );
  XNOR U21760 ( .A(a[563]), .B(n18227), .Z(n491) );
  IV U21761 ( .A(n18225), .Z(n18227) );
  XNOR U21762 ( .A(b[563]), .B(n18225), .Z(n18226) );
  XOR U21763 ( .A(n18228), .B(n18229), .Z(n18225) );
  ANDN U21764 ( .B(n18230), .A(n492), .Z(n18228) );
  XNOR U21765 ( .A(a[562]), .B(n18231), .Z(n492) );
  IV U21766 ( .A(n18229), .Z(n18231) );
  XNOR U21767 ( .A(b[562]), .B(n18229), .Z(n18230) );
  XOR U21768 ( .A(n18232), .B(n18233), .Z(n18229) );
  ANDN U21769 ( .B(n18234), .A(n493), .Z(n18232) );
  XNOR U21770 ( .A(a[561]), .B(n18235), .Z(n493) );
  IV U21771 ( .A(n18233), .Z(n18235) );
  XNOR U21772 ( .A(b[561]), .B(n18233), .Z(n18234) );
  XOR U21773 ( .A(n18236), .B(n18237), .Z(n18233) );
  ANDN U21774 ( .B(n18238), .A(n494), .Z(n18236) );
  XNOR U21775 ( .A(a[560]), .B(n18239), .Z(n494) );
  IV U21776 ( .A(n18237), .Z(n18239) );
  XNOR U21777 ( .A(b[560]), .B(n18237), .Z(n18238) );
  XOR U21778 ( .A(n18240), .B(n18241), .Z(n18237) );
  ANDN U21779 ( .B(n18242), .A(n496), .Z(n18240) );
  XNOR U21780 ( .A(a[559]), .B(n18243), .Z(n496) );
  IV U21781 ( .A(n18241), .Z(n18243) );
  XNOR U21782 ( .A(b[559]), .B(n18241), .Z(n18242) );
  XOR U21783 ( .A(n18244), .B(n18245), .Z(n18241) );
  ANDN U21784 ( .B(n18246), .A(n497), .Z(n18244) );
  XNOR U21785 ( .A(a[558]), .B(n18247), .Z(n497) );
  IV U21786 ( .A(n18245), .Z(n18247) );
  XNOR U21787 ( .A(b[558]), .B(n18245), .Z(n18246) );
  XOR U21788 ( .A(n18248), .B(n18249), .Z(n18245) );
  ANDN U21789 ( .B(n18250), .A(n498), .Z(n18248) );
  XNOR U21790 ( .A(a[557]), .B(n18251), .Z(n498) );
  IV U21791 ( .A(n18249), .Z(n18251) );
  XNOR U21792 ( .A(b[557]), .B(n18249), .Z(n18250) );
  XOR U21793 ( .A(n18252), .B(n18253), .Z(n18249) );
  ANDN U21794 ( .B(n18254), .A(n499), .Z(n18252) );
  XNOR U21795 ( .A(a[556]), .B(n18255), .Z(n499) );
  IV U21796 ( .A(n18253), .Z(n18255) );
  XNOR U21797 ( .A(b[556]), .B(n18253), .Z(n18254) );
  XOR U21798 ( .A(n18256), .B(n18257), .Z(n18253) );
  ANDN U21799 ( .B(n18258), .A(n500), .Z(n18256) );
  XNOR U21800 ( .A(a[555]), .B(n18259), .Z(n500) );
  IV U21801 ( .A(n18257), .Z(n18259) );
  XNOR U21802 ( .A(b[555]), .B(n18257), .Z(n18258) );
  XOR U21803 ( .A(n18260), .B(n18261), .Z(n18257) );
  ANDN U21804 ( .B(n18262), .A(n501), .Z(n18260) );
  XNOR U21805 ( .A(a[554]), .B(n18263), .Z(n501) );
  IV U21806 ( .A(n18261), .Z(n18263) );
  XNOR U21807 ( .A(b[554]), .B(n18261), .Z(n18262) );
  XOR U21808 ( .A(n18264), .B(n18265), .Z(n18261) );
  ANDN U21809 ( .B(n18266), .A(n502), .Z(n18264) );
  XNOR U21810 ( .A(a[553]), .B(n18267), .Z(n502) );
  IV U21811 ( .A(n18265), .Z(n18267) );
  XNOR U21812 ( .A(b[553]), .B(n18265), .Z(n18266) );
  XOR U21813 ( .A(n18268), .B(n18269), .Z(n18265) );
  ANDN U21814 ( .B(n18270), .A(n503), .Z(n18268) );
  XNOR U21815 ( .A(a[552]), .B(n18271), .Z(n503) );
  IV U21816 ( .A(n18269), .Z(n18271) );
  XNOR U21817 ( .A(b[552]), .B(n18269), .Z(n18270) );
  XOR U21818 ( .A(n18272), .B(n18273), .Z(n18269) );
  ANDN U21819 ( .B(n18274), .A(n504), .Z(n18272) );
  XNOR U21820 ( .A(a[551]), .B(n18275), .Z(n504) );
  IV U21821 ( .A(n18273), .Z(n18275) );
  XNOR U21822 ( .A(b[551]), .B(n18273), .Z(n18274) );
  XOR U21823 ( .A(n18276), .B(n18277), .Z(n18273) );
  ANDN U21824 ( .B(n18278), .A(n505), .Z(n18276) );
  XNOR U21825 ( .A(a[550]), .B(n18279), .Z(n505) );
  IV U21826 ( .A(n18277), .Z(n18279) );
  XNOR U21827 ( .A(b[550]), .B(n18277), .Z(n18278) );
  XOR U21828 ( .A(n18280), .B(n18281), .Z(n18277) );
  ANDN U21829 ( .B(n18282), .A(n507), .Z(n18280) );
  XNOR U21830 ( .A(a[549]), .B(n18283), .Z(n507) );
  IV U21831 ( .A(n18281), .Z(n18283) );
  XNOR U21832 ( .A(b[549]), .B(n18281), .Z(n18282) );
  XOR U21833 ( .A(n18284), .B(n18285), .Z(n18281) );
  ANDN U21834 ( .B(n18286), .A(n508), .Z(n18284) );
  XNOR U21835 ( .A(a[548]), .B(n18287), .Z(n508) );
  IV U21836 ( .A(n18285), .Z(n18287) );
  XNOR U21837 ( .A(b[548]), .B(n18285), .Z(n18286) );
  XOR U21838 ( .A(n18288), .B(n18289), .Z(n18285) );
  ANDN U21839 ( .B(n18290), .A(n509), .Z(n18288) );
  XNOR U21840 ( .A(a[547]), .B(n18291), .Z(n509) );
  IV U21841 ( .A(n18289), .Z(n18291) );
  XNOR U21842 ( .A(b[547]), .B(n18289), .Z(n18290) );
  XOR U21843 ( .A(n18292), .B(n18293), .Z(n18289) );
  ANDN U21844 ( .B(n18294), .A(n510), .Z(n18292) );
  XNOR U21845 ( .A(a[546]), .B(n18295), .Z(n510) );
  IV U21846 ( .A(n18293), .Z(n18295) );
  XNOR U21847 ( .A(b[546]), .B(n18293), .Z(n18294) );
  XOR U21848 ( .A(n18296), .B(n18297), .Z(n18293) );
  ANDN U21849 ( .B(n18298), .A(n511), .Z(n18296) );
  XNOR U21850 ( .A(a[545]), .B(n18299), .Z(n511) );
  IV U21851 ( .A(n18297), .Z(n18299) );
  XNOR U21852 ( .A(b[545]), .B(n18297), .Z(n18298) );
  XOR U21853 ( .A(n18300), .B(n18301), .Z(n18297) );
  ANDN U21854 ( .B(n18302), .A(n512), .Z(n18300) );
  XNOR U21855 ( .A(a[544]), .B(n18303), .Z(n512) );
  IV U21856 ( .A(n18301), .Z(n18303) );
  XNOR U21857 ( .A(b[544]), .B(n18301), .Z(n18302) );
  XOR U21858 ( .A(n18304), .B(n18305), .Z(n18301) );
  ANDN U21859 ( .B(n18306), .A(n513), .Z(n18304) );
  XNOR U21860 ( .A(a[543]), .B(n18307), .Z(n513) );
  IV U21861 ( .A(n18305), .Z(n18307) );
  XNOR U21862 ( .A(b[543]), .B(n18305), .Z(n18306) );
  XOR U21863 ( .A(n18308), .B(n18309), .Z(n18305) );
  ANDN U21864 ( .B(n18310), .A(n514), .Z(n18308) );
  XNOR U21865 ( .A(a[542]), .B(n18311), .Z(n514) );
  IV U21866 ( .A(n18309), .Z(n18311) );
  XNOR U21867 ( .A(b[542]), .B(n18309), .Z(n18310) );
  XOR U21868 ( .A(n18312), .B(n18313), .Z(n18309) );
  ANDN U21869 ( .B(n18314), .A(n515), .Z(n18312) );
  XNOR U21870 ( .A(a[541]), .B(n18315), .Z(n515) );
  IV U21871 ( .A(n18313), .Z(n18315) );
  XNOR U21872 ( .A(b[541]), .B(n18313), .Z(n18314) );
  XOR U21873 ( .A(n18316), .B(n18317), .Z(n18313) );
  ANDN U21874 ( .B(n18318), .A(n516), .Z(n18316) );
  XNOR U21875 ( .A(a[540]), .B(n18319), .Z(n516) );
  IV U21876 ( .A(n18317), .Z(n18319) );
  XNOR U21877 ( .A(b[540]), .B(n18317), .Z(n18318) );
  XOR U21878 ( .A(n18320), .B(n18321), .Z(n18317) );
  ANDN U21879 ( .B(n18322), .A(n518), .Z(n18320) );
  XNOR U21880 ( .A(a[539]), .B(n18323), .Z(n518) );
  IV U21881 ( .A(n18321), .Z(n18323) );
  XNOR U21882 ( .A(b[539]), .B(n18321), .Z(n18322) );
  XOR U21883 ( .A(n18324), .B(n18325), .Z(n18321) );
  ANDN U21884 ( .B(n18326), .A(n519), .Z(n18324) );
  XNOR U21885 ( .A(a[538]), .B(n18327), .Z(n519) );
  IV U21886 ( .A(n18325), .Z(n18327) );
  XNOR U21887 ( .A(b[538]), .B(n18325), .Z(n18326) );
  XOR U21888 ( .A(n18328), .B(n18329), .Z(n18325) );
  ANDN U21889 ( .B(n18330), .A(n520), .Z(n18328) );
  XNOR U21890 ( .A(a[537]), .B(n18331), .Z(n520) );
  IV U21891 ( .A(n18329), .Z(n18331) );
  XNOR U21892 ( .A(b[537]), .B(n18329), .Z(n18330) );
  XOR U21893 ( .A(n18332), .B(n18333), .Z(n18329) );
  ANDN U21894 ( .B(n18334), .A(n521), .Z(n18332) );
  XNOR U21895 ( .A(a[536]), .B(n18335), .Z(n521) );
  IV U21896 ( .A(n18333), .Z(n18335) );
  XNOR U21897 ( .A(b[536]), .B(n18333), .Z(n18334) );
  XOR U21898 ( .A(n18336), .B(n18337), .Z(n18333) );
  ANDN U21899 ( .B(n18338), .A(n522), .Z(n18336) );
  XNOR U21900 ( .A(a[535]), .B(n18339), .Z(n522) );
  IV U21901 ( .A(n18337), .Z(n18339) );
  XNOR U21902 ( .A(b[535]), .B(n18337), .Z(n18338) );
  XOR U21903 ( .A(n18340), .B(n18341), .Z(n18337) );
  ANDN U21904 ( .B(n18342), .A(n523), .Z(n18340) );
  XNOR U21905 ( .A(a[534]), .B(n18343), .Z(n523) );
  IV U21906 ( .A(n18341), .Z(n18343) );
  XNOR U21907 ( .A(b[534]), .B(n18341), .Z(n18342) );
  XOR U21908 ( .A(n18344), .B(n18345), .Z(n18341) );
  ANDN U21909 ( .B(n18346), .A(n524), .Z(n18344) );
  XNOR U21910 ( .A(a[533]), .B(n18347), .Z(n524) );
  IV U21911 ( .A(n18345), .Z(n18347) );
  XNOR U21912 ( .A(b[533]), .B(n18345), .Z(n18346) );
  XOR U21913 ( .A(n18348), .B(n18349), .Z(n18345) );
  ANDN U21914 ( .B(n18350), .A(n525), .Z(n18348) );
  XNOR U21915 ( .A(a[532]), .B(n18351), .Z(n525) );
  IV U21916 ( .A(n18349), .Z(n18351) );
  XNOR U21917 ( .A(b[532]), .B(n18349), .Z(n18350) );
  XOR U21918 ( .A(n18352), .B(n18353), .Z(n18349) );
  ANDN U21919 ( .B(n18354), .A(n526), .Z(n18352) );
  XNOR U21920 ( .A(a[531]), .B(n18355), .Z(n526) );
  IV U21921 ( .A(n18353), .Z(n18355) );
  XNOR U21922 ( .A(b[531]), .B(n18353), .Z(n18354) );
  XOR U21923 ( .A(n18356), .B(n18357), .Z(n18353) );
  ANDN U21924 ( .B(n18358), .A(n527), .Z(n18356) );
  XNOR U21925 ( .A(a[530]), .B(n18359), .Z(n527) );
  IV U21926 ( .A(n18357), .Z(n18359) );
  XNOR U21927 ( .A(b[530]), .B(n18357), .Z(n18358) );
  XOR U21928 ( .A(n18360), .B(n18361), .Z(n18357) );
  ANDN U21929 ( .B(n18362), .A(n529), .Z(n18360) );
  XNOR U21930 ( .A(a[529]), .B(n18363), .Z(n529) );
  IV U21931 ( .A(n18361), .Z(n18363) );
  XNOR U21932 ( .A(b[529]), .B(n18361), .Z(n18362) );
  XOR U21933 ( .A(n18364), .B(n18365), .Z(n18361) );
  ANDN U21934 ( .B(n18366), .A(n530), .Z(n18364) );
  XNOR U21935 ( .A(a[528]), .B(n18367), .Z(n530) );
  IV U21936 ( .A(n18365), .Z(n18367) );
  XNOR U21937 ( .A(b[528]), .B(n18365), .Z(n18366) );
  XOR U21938 ( .A(n18368), .B(n18369), .Z(n18365) );
  ANDN U21939 ( .B(n18370), .A(n531), .Z(n18368) );
  XNOR U21940 ( .A(a[527]), .B(n18371), .Z(n531) );
  IV U21941 ( .A(n18369), .Z(n18371) );
  XNOR U21942 ( .A(b[527]), .B(n18369), .Z(n18370) );
  XOR U21943 ( .A(n18372), .B(n18373), .Z(n18369) );
  ANDN U21944 ( .B(n18374), .A(n532), .Z(n18372) );
  XNOR U21945 ( .A(a[526]), .B(n18375), .Z(n532) );
  IV U21946 ( .A(n18373), .Z(n18375) );
  XNOR U21947 ( .A(b[526]), .B(n18373), .Z(n18374) );
  XOR U21948 ( .A(n18376), .B(n18377), .Z(n18373) );
  ANDN U21949 ( .B(n18378), .A(n533), .Z(n18376) );
  XNOR U21950 ( .A(a[525]), .B(n18379), .Z(n533) );
  IV U21951 ( .A(n18377), .Z(n18379) );
  XNOR U21952 ( .A(b[525]), .B(n18377), .Z(n18378) );
  XOR U21953 ( .A(n18380), .B(n18381), .Z(n18377) );
  ANDN U21954 ( .B(n18382), .A(n534), .Z(n18380) );
  XNOR U21955 ( .A(a[524]), .B(n18383), .Z(n534) );
  IV U21956 ( .A(n18381), .Z(n18383) );
  XNOR U21957 ( .A(b[524]), .B(n18381), .Z(n18382) );
  XOR U21958 ( .A(n18384), .B(n18385), .Z(n18381) );
  ANDN U21959 ( .B(n18386), .A(n535), .Z(n18384) );
  XNOR U21960 ( .A(a[523]), .B(n18387), .Z(n535) );
  IV U21961 ( .A(n18385), .Z(n18387) );
  XNOR U21962 ( .A(b[523]), .B(n18385), .Z(n18386) );
  XOR U21963 ( .A(n18388), .B(n18389), .Z(n18385) );
  ANDN U21964 ( .B(n18390), .A(n536), .Z(n18388) );
  XNOR U21965 ( .A(a[522]), .B(n18391), .Z(n536) );
  IV U21966 ( .A(n18389), .Z(n18391) );
  XNOR U21967 ( .A(b[522]), .B(n18389), .Z(n18390) );
  XOR U21968 ( .A(n18392), .B(n18393), .Z(n18389) );
  ANDN U21969 ( .B(n18394), .A(n537), .Z(n18392) );
  XNOR U21970 ( .A(a[521]), .B(n18395), .Z(n537) );
  IV U21971 ( .A(n18393), .Z(n18395) );
  XNOR U21972 ( .A(b[521]), .B(n18393), .Z(n18394) );
  XOR U21973 ( .A(n18396), .B(n18397), .Z(n18393) );
  ANDN U21974 ( .B(n18398), .A(n538), .Z(n18396) );
  XNOR U21975 ( .A(a[520]), .B(n18399), .Z(n538) );
  IV U21976 ( .A(n18397), .Z(n18399) );
  XNOR U21977 ( .A(b[520]), .B(n18397), .Z(n18398) );
  XOR U21978 ( .A(n18400), .B(n18401), .Z(n18397) );
  ANDN U21979 ( .B(n18402), .A(n540), .Z(n18400) );
  XNOR U21980 ( .A(a[519]), .B(n18403), .Z(n540) );
  IV U21981 ( .A(n18401), .Z(n18403) );
  XNOR U21982 ( .A(b[519]), .B(n18401), .Z(n18402) );
  XOR U21983 ( .A(n18404), .B(n18405), .Z(n18401) );
  ANDN U21984 ( .B(n18406), .A(n541), .Z(n18404) );
  XNOR U21985 ( .A(a[518]), .B(n18407), .Z(n541) );
  IV U21986 ( .A(n18405), .Z(n18407) );
  XNOR U21987 ( .A(b[518]), .B(n18405), .Z(n18406) );
  XOR U21988 ( .A(n18408), .B(n18409), .Z(n18405) );
  ANDN U21989 ( .B(n18410), .A(n542), .Z(n18408) );
  XNOR U21990 ( .A(a[517]), .B(n18411), .Z(n542) );
  IV U21991 ( .A(n18409), .Z(n18411) );
  XNOR U21992 ( .A(b[517]), .B(n18409), .Z(n18410) );
  XOR U21993 ( .A(n18412), .B(n18413), .Z(n18409) );
  ANDN U21994 ( .B(n18414), .A(n543), .Z(n18412) );
  XNOR U21995 ( .A(a[516]), .B(n18415), .Z(n543) );
  IV U21996 ( .A(n18413), .Z(n18415) );
  XNOR U21997 ( .A(b[516]), .B(n18413), .Z(n18414) );
  XOR U21998 ( .A(n18416), .B(n18417), .Z(n18413) );
  ANDN U21999 ( .B(n18418), .A(n544), .Z(n18416) );
  XNOR U22000 ( .A(a[515]), .B(n18419), .Z(n544) );
  IV U22001 ( .A(n18417), .Z(n18419) );
  XNOR U22002 ( .A(b[515]), .B(n18417), .Z(n18418) );
  XOR U22003 ( .A(n18420), .B(n18421), .Z(n18417) );
  ANDN U22004 ( .B(n18422), .A(n545), .Z(n18420) );
  XNOR U22005 ( .A(a[514]), .B(n18423), .Z(n545) );
  IV U22006 ( .A(n18421), .Z(n18423) );
  XNOR U22007 ( .A(b[514]), .B(n18421), .Z(n18422) );
  XOR U22008 ( .A(n18424), .B(n18425), .Z(n18421) );
  ANDN U22009 ( .B(n18426), .A(n546), .Z(n18424) );
  XNOR U22010 ( .A(a[513]), .B(n18427), .Z(n546) );
  IV U22011 ( .A(n18425), .Z(n18427) );
  XNOR U22012 ( .A(b[513]), .B(n18425), .Z(n18426) );
  XOR U22013 ( .A(n18428), .B(n18429), .Z(n18425) );
  ANDN U22014 ( .B(n18430), .A(n547), .Z(n18428) );
  XNOR U22015 ( .A(a[512]), .B(n18431), .Z(n547) );
  IV U22016 ( .A(n18429), .Z(n18431) );
  XNOR U22017 ( .A(b[512]), .B(n18429), .Z(n18430) );
  XOR U22018 ( .A(n18432), .B(n18433), .Z(n18429) );
  ANDN U22019 ( .B(n18434), .A(n548), .Z(n18432) );
  XNOR U22020 ( .A(a[511]), .B(n18435), .Z(n548) );
  IV U22021 ( .A(n18433), .Z(n18435) );
  XNOR U22022 ( .A(b[511]), .B(n18433), .Z(n18434) );
  XOR U22023 ( .A(n18436), .B(n18437), .Z(n18433) );
  ANDN U22024 ( .B(n18438), .A(n549), .Z(n18436) );
  XNOR U22025 ( .A(a[510]), .B(n18439), .Z(n549) );
  IV U22026 ( .A(n18437), .Z(n18439) );
  XNOR U22027 ( .A(b[510]), .B(n18437), .Z(n18438) );
  XOR U22028 ( .A(n18440), .B(n18441), .Z(n18437) );
  ANDN U22029 ( .B(n18442), .A(n551), .Z(n18440) );
  XNOR U22030 ( .A(a[509]), .B(n18443), .Z(n551) );
  IV U22031 ( .A(n18441), .Z(n18443) );
  XNOR U22032 ( .A(b[509]), .B(n18441), .Z(n18442) );
  XOR U22033 ( .A(n18444), .B(n18445), .Z(n18441) );
  ANDN U22034 ( .B(n18446), .A(n552), .Z(n18444) );
  XNOR U22035 ( .A(a[508]), .B(n18447), .Z(n552) );
  IV U22036 ( .A(n18445), .Z(n18447) );
  XNOR U22037 ( .A(b[508]), .B(n18445), .Z(n18446) );
  XOR U22038 ( .A(n18448), .B(n18449), .Z(n18445) );
  ANDN U22039 ( .B(n18450), .A(n553), .Z(n18448) );
  XNOR U22040 ( .A(a[507]), .B(n18451), .Z(n553) );
  IV U22041 ( .A(n18449), .Z(n18451) );
  XNOR U22042 ( .A(b[507]), .B(n18449), .Z(n18450) );
  XOR U22043 ( .A(n18452), .B(n18453), .Z(n18449) );
  ANDN U22044 ( .B(n18454), .A(n554), .Z(n18452) );
  XNOR U22045 ( .A(a[506]), .B(n18455), .Z(n554) );
  IV U22046 ( .A(n18453), .Z(n18455) );
  XNOR U22047 ( .A(b[506]), .B(n18453), .Z(n18454) );
  XOR U22048 ( .A(n18456), .B(n18457), .Z(n18453) );
  ANDN U22049 ( .B(n18458), .A(n555), .Z(n18456) );
  XNOR U22050 ( .A(a[505]), .B(n18459), .Z(n555) );
  IV U22051 ( .A(n18457), .Z(n18459) );
  XNOR U22052 ( .A(b[505]), .B(n18457), .Z(n18458) );
  XOR U22053 ( .A(n18460), .B(n18461), .Z(n18457) );
  ANDN U22054 ( .B(n18462), .A(n556), .Z(n18460) );
  XNOR U22055 ( .A(a[504]), .B(n18463), .Z(n556) );
  IV U22056 ( .A(n18461), .Z(n18463) );
  XNOR U22057 ( .A(b[504]), .B(n18461), .Z(n18462) );
  XOR U22058 ( .A(n18464), .B(n18465), .Z(n18461) );
  ANDN U22059 ( .B(n18466), .A(n557), .Z(n18464) );
  XNOR U22060 ( .A(a[503]), .B(n18467), .Z(n557) );
  IV U22061 ( .A(n18465), .Z(n18467) );
  XNOR U22062 ( .A(b[503]), .B(n18465), .Z(n18466) );
  XOR U22063 ( .A(n18468), .B(n18469), .Z(n18465) );
  ANDN U22064 ( .B(n18470), .A(n558), .Z(n18468) );
  XNOR U22065 ( .A(a[502]), .B(n18471), .Z(n558) );
  IV U22066 ( .A(n18469), .Z(n18471) );
  XNOR U22067 ( .A(b[502]), .B(n18469), .Z(n18470) );
  XOR U22068 ( .A(n18472), .B(n18473), .Z(n18469) );
  ANDN U22069 ( .B(n18474), .A(n559), .Z(n18472) );
  XNOR U22070 ( .A(a[501]), .B(n18475), .Z(n559) );
  IV U22071 ( .A(n18473), .Z(n18475) );
  XNOR U22072 ( .A(b[501]), .B(n18473), .Z(n18474) );
  XOR U22073 ( .A(n18476), .B(n18477), .Z(n18473) );
  ANDN U22074 ( .B(n18478), .A(n560), .Z(n18476) );
  XNOR U22075 ( .A(a[500]), .B(n18479), .Z(n560) );
  IV U22076 ( .A(n18477), .Z(n18479) );
  XNOR U22077 ( .A(b[500]), .B(n18477), .Z(n18478) );
  XOR U22078 ( .A(n18480), .B(n18481), .Z(n18477) );
  ANDN U22079 ( .B(n18482), .A(n563), .Z(n18480) );
  XNOR U22080 ( .A(a[499]), .B(n18483), .Z(n563) );
  IV U22081 ( .A(n18481), .Z(n18483) );
  XNOR U22082 ( .A(b[499]), .B(n18481), .Z(n18482) );
  XOR U22083 ( .A(n18484), .B(n18485), .Z(n18481) );
  ANDN U22084 ( .B(n18486), .A(n564), .Z(n18484) );
  XNOR U22085 ( .A(a[498]), .B(n18487), .Z(n564) );
  IV U22086 ( .A(n18485), .Z(n18487) );
  XNOR U22087 ( .A(b[498]), .B(n18485), .Z(n18486) );
  XOR U22088 ( .A(n18488), .B(n18489), .Z(n18485) );
  ANDN U22089 ( .B(n18490), .A(n565), .Z(n18488) );
  XNOR U22090 ( .A(a[497]), .B(n18491), .Z(n565) );
  IV U22091 ( .A(n18489), .Z(n18491) );
  XNOR U22092 ( .A(b[497]), .B(n18489), .Z(n18490) );
  XOR U22093 ( .A(n18492), .B(n18493), .Z(n18489) );
  ANDN U22094 ( .B(n18494), .A(n566), .Z(n18492) );
  XNOR U22095 ( .A(a[496]), .B(n18495), .Z(n566) );
  IV U22096 ( .A(n18493), .Z(n18495) );
  XNOR U22097 ( .A(b[496]), .B(n18493), .Z(n18494) );
  XOR U22098 ( .A(n18496), .B(n18497), .Z(n18493) );
  ANDN U22099 ( .B(n18498), .A(n567), .Z(n18496) );
  XNOR U22100 ( .A(a[495]), .B(n18499), .Z(n567) );
  IV U22101 ( .A(n18497), .Z(n18499) );
  XNOR U22102 ( .A(b[495]), .B(n18497), .Z(n18498) );
  XOR U22103 ( .A(n18500), .B(n18501), .Z(n18497) );
  ANDN U22104 ( .B(n18502), .A(n568), .Z(n18500) );
  XNOR U22105 ( .A(a[494]), .B(n18503), .Z(n568) );
  IV U22106 ( .A(n18501), .Z(n18503) );
  XNOR U22107 ( .A(b[494]), .B(n18501), .Z(n18502) );
  XOR U22108 ( .A(n18504), .B(n18505), .Z(n18501) );
  ANDN U22109 ( .B(n18506), .A(n569), .Z(n18504) );
  XNOR U22110 ( .A(a[493]), .B(n18507), .Z(n569) );
  IV U22111 ( .A(n18505), .Z(n18507) );
  XNOR U22112 ( .A(b[493]), .B(n18505), .Z(n18506) );
  XOR U22113 ( .A(n18508), .B(n18509), .Z(n18505) );
  ANDN U22114 ( .B(n18510), .A(n570), .Z(n18508) );
  XNOR U22115 ( .A(a[492]), .B(n18511), .Z(n570) );
  IV U22116 ( .A(n18509), .Z(n18511) );
  XNOR U22117 ( .A(b[492]), .B(n18509), .Z(n18510) );
  XOR U22118 ( .A(n18512), .B(n18513), .Z(n18509) );
  ANDN U22119 ( .B(n18514), .A(n571), .Z(n18512) );
  XNOR U22120 ( .A(a[491]), .B(n18515), .Z(n571) );
  IV U22121 ( .A(n18513), .Z(n18515) );
  XNOR U22122 ( .A(b[491]), .B(n18513), .Z(n18514) );
  XOR U22123 ( .A(n18516), .B(n18517), .Z(n18513) );
  ANDN U22124 ( .B(n18518), .A(n572), .Z(n18516) );
  XNOR U22125 ( .A(a[490]), .B(n18519), .Z(n572) );
  IV U22126 ( .A(n18517), .Z(n18519) );
  XNOR U22127 ( .A(b[490]), .B(n18517), .Z(n18518) );
  XOR U22128 ( .A(n18520), .B(n18521), .Z(n18517) );
  ANDN U22129 ( .B(n18522), .A(n574), .Z(n18520) );
  XNOR U22130 ( .A(a[489]), .B(n18523), .Z(n574) );
  IV U22131 ( .A(n18521), .Z(n18523) );
  XNOR U22132 ( .A(b[489]), .B(n18521), .Z(n18522) );
  XOR U22133 ( .A(n18524), .B(n18525), .Z(n18521) );
  ANDN U22134 ( .B(n18526), .A(n575), .Z(n18524) );
  XNOR U22135 ( .A(a[488]), .B(n18527), .Z(n575) );
  IV U22136 ( .A(n18525), .Z(n18527) );
  XNOR U22137 ( .A(b[488]), .B(n18525), .Z(n18526) );
  XOR U22138 ( .A(n18528), .B(n18529), .Z(n18525) );
  ANDN U22139 ( .B(n18530), .A(n576), .Z(n18528) );
  XNOR U22140 ( .A(a[487]), .B(n18531), .Z(n576) );
  IV U22141 ( .A(n18529), .Z(n18531) );
  XNOR U22142 ( .A(b[487]), .B(n18529), .Z(n18530) );
  XOR U22143 ( .A(n18532), .B(n18533), .Z(n18529) );
  ANDN U22144 ( .B(n18534), .A(n577), .Z(n18532) );
  XNOR U22145 ( .A(a[486]), .B(n18535), .Z(n577) );
  IV U22146 ( .A(n18533), .Z(n18535) );
  XNOR U22147 ( .A(b[486]), .B(n18533), .Z(n18534) );
  XOR U22148 ( .A(n18536), .B(n18537), .Z(n18533) );
  ANDN U22149 ( .B(n18538), .A(n578), .Z(n18536) );
  XNOR U22150 ( .A(a[485]), .B(n18539), .Z(n578) );
  IV U22151 ( .A(n18537), .Z(n18539) );
  XNOR U22152 ( .A(b[485]), .B(n18537), .Z(n18538) );
  XOR U22153 ( .A(n18540), .B(n18541), .Z(n18537) );
  ANDN U22154 ( .B(n18542), .A(n579), .Z(n18540) );
  XNOR U22155 ( .A(a[484]), .B(n18543), .Z(n579) );
  IV U22156 ( .A(n18541), .Z(n18543) );
  XNOR U22157 ( .A(b[484]), .B(n18541), .Z(n18542) );
  XOR U22158 ( .A(n18544), .B(n18545), .Z(n18541) );
  ANDN U22159 ( .B(n18546), .A(n580), .Z(n18544) );
  XNOR U22160 ( .A(a[483]), .B(n18547), .Z(n580) );
  IV U22161 ( .A(n18545), .Z(n18547) );
  XNOR U22162 ( .A(b[483]), .B(n18545), .Z(n18546) );
  XOR U22163 ( .A(n18548), .B(n18549), .Z(n18545) );
  ANDN U22164 ( .B(n18550), .A(n581), .Z(n18548) );
  XNOR U22165 ( .A(a[482]), .B(n18551), .Z(n581) );
  IV U22166 ( .A(n18549), .Z(n18551) );
  XNOR U22167 ( .A(b[482]), .B(n18549), .Z(n18550) );
  XOR U22168 ( .A(n18552), .B(n18553), .Z(n18549) );
  ANDN U22169 ( .B(n18554), .A(n582), .Z(n18552) );
  XNOR U22170 ( .A(a[481]), .B(n18555), .Z(n582) );
  IV U22171 ( .A(n18553), .Z(n18555) );
  XNOR U22172 ( .A(b[481]), .B(n18553), .Z(n18554) );
  XOR U22173 ( .A(n18556), .B(n18557), .Z(n18553) );
  ANDN U22174 ( .B(n18558), .A(n583), .Z(n18556) );
  XNOR U22175 ( .A(a[480]), .B(n18559), .Z(n583) );
  IV U22176 ( .A(n18557), .Z(n18559) );
  XNOR U22177 ( .A(b[480]), .B(n18557), .Z(n18558) );
  XOR U22178 ( .A(n18560), .B(n18561), .Z(n18557) );
  ANDN U22179 ( .B(n18562), .A(n585), .Z(n18560) );
  XNOR U22180 ( .A(a[479]), .B(n18563), .Z(n585) );
  IV U22181 ( .A(n18561), .Z(n18563) );
  XNOR U22182 ( .A(b[479]), .B(n18561), .Z(n18562) );
  XOR U22183 ( .A(n18564), .B(n18565), .Z(n18561) );
  ANDN U22184 ( .B(n18566), .A(n586), .Z(n18564) );
  XNOR U22185 ( .A(a[478]), .B(n18567), .Z(n586) );
  IV U22186 ( .A(n18565), .Z(n18567) );
  XNOR U22187 ( .A(b[478]), .B(n18565), .Z(n18566) );
  XOR U22188 ( .A(n18568), .B(n18569), .Z(n18565) );
  ANDN U22189 ( .B(n18570), .A(n587), .Z(n18568) );
  XNOR U22190 ( .A(a[477]), .B(n18571), .Z(n587) );
  IV U22191 ( .A(n18569), .Z(n18571) );
  XNOR U22192 ( .A(b[477]), .B(n18569), .Z(n18570) );
  XOR U22193 ( .A(n18572), .B(n18573), .Z(n18569) );
  ANDN U22194 ( .B(n18574), .A(n588), .Z(n18572) );
  XNOR U22195 ( .A(a[476]), .B(n18575), .Z(n588) );
  IV U22196 ( .A(n18573), .Z(n18575) );
  XNOR U22197 ( .A(b[476]), .B(n18573), .Z(n18574) );
  XOR U22198 ( .A(n18576), .B(n18577), .Z(n18573) );
  ANDN U22199 ( .B(n18578), .A(n589), .Z(n18576) );
  XNOR U22200 ( .A(a[475]), .B(n18579), .Z(n589) );
  IV U22201 ( .A(n18577), .Z(n18579) );
  XNOR U22202 ( .A(b[475]), .B(n18577), .Z(n18578) );
  XOR U22203 ( .A(n18580), .B(n18581), .Z(n18577) );
  ANDN U22204 ( .B(n18582), .A(n590), .Z(n18580) );
  XNOR U22205 ( .A(a[474]), .B(n18583), .Z(n590) );
  IV U22206 ( .A(n18581), .Z(n18583) );
  XNOR U22207 ( .A(b[474]), .B(n18581), .Z(n18582) );
  XOR U22208 ( .A(n18584), .B(n18585), .Z(n18581) );
  ANDN U22209 ( .B(n18586), .A(n591), .Z(n18584) );
  XNOR U22210 ( .A(a[473]), .B(n18587), .Z(n591) );
  IV U22211 ( .A(n18585), .Z(n18587) );
  XNOR U22212 ( .A(b[473]), .B(n18585), .Z(n18586) );
  XOR U22213 ( .A(n18588), .B(n18589), .Z(n18585) );
  ANDN U22214 ( .B(n18590), .A(n592), .Z(n18588) );
  XNOR U22215 ( .A(a[472]), .B(n18591), .Z(n592) );
  IV U22216 ( .A(n18589), .Z(n18591) );
  XNOR U22217 ( .A(b[472]), .B(n18589), .Z(n18590) );
  XOR U22218 ( .A(n18592), .B(n18593), .Z(n18589) );
  ANDN U22219 ( .B(n18594), .A(n593), .Z(n18592) );
  XNOR U22220 ( .A(a[471]), .B(n18595), .Z(n593) );
  IV U22221 ( .A(n18593), .Z(n18595) );
  XNOR U22222 ( .A(b[471]), .B(n18593), .Z(n18594) );
  XOR U22223 ( .A(n18596), .B(n18597), .Z(n18593) );
  ANDN U22224 ( .B(n18598), .A(n594), .Z(n18596) );
  XNOR U22225 ( .A(a[470]), .B(n18599), .Z(n594) );
  IV U22226 ( .A(n18597), .Z(n18599) );
  XNOR U22227 ( .A(b[470]), .B(n18597), .Z(n18598) );
  XOR U22228 ( .A(n18600), .B(n18601), .Z(n18597) );
  ANDN U22229 ( .B(n18602), .A(n596), .Z(n18600) );
  XNOR U22230 ( .A(a[469]), .B(n18603), .Z(n596) );
  IV U22231 ( .A(n18601), .Z(n18603) );
  XNOR U22232 ( .A(b[469]), .B(n18601), .Z(n18602) );
  XOR U22233 ( .A(n18604), .B(n18605), .Z(n18601) );
  ANDN U22234 ( .B(n18606), .A(n597), .Z(n18604) );
  XNOR U22235 ( .A(a[468]), .B(n18607), .Z(n597) );
  IV U22236 ( .A(n18605), .Z(n18607) );
  XNOR U22237 ( .A(b[468]), .B(n18605), .Z(n18606) );
  XOR U22238 ( .A(n18608), .B(n18609), .Z(n18605) );
  ANDN U22239 ( .B(n18610), .A(n598), .Z(n18608) );
  XNOR U22240 ( .A(a[467]), .B(n18611), .Z(n598) );
  IV U22241 ( .A(n18609), .Z(n18611) );
  XNOR U22242 ( .A(b[467]), .B(n18609), .Z(n18610) );
  XOR U22243 ( .A(n18612), .B(n18613), .Z(n18609) );
  ANDN U22244 ( .B(n18614), .A(n599), .Z(n18612) );
  XNOR U22245 ( .A(a[466]), .B(n18615), .Z(n599) );
  IV U22246 ( .A(n18613), .Z(n18615) );
  XNOR U22247 ( .A(b[466]), .B(n18613), .Z(n18614) );
  XOR U22248 ( .A(n18616), .B(n18617), .Z(n18613) );
  ANDN U22249 ( .B(n18618), .A(n600), .Z(n18616) );
  XNOR U22250 ( .A(a[465]), .B(n18619), .Z(n600) );
  IV U22251 ( .A(n18617), .Z(n18619) );
  XNOR U22252 ( .A(b[465]), .B(n18617), .Z(n18618) );
  XOR U22253 ( .A(n18620), .B(n18621), .Z(n18617) );
  ANDN U22254 ( .B(n18622), .A(n601), .Z(n18620) );
  XNOR U22255 ( .A(a[464]), .B(n18623), .Z(n601) );
  IV U22256 ( .A(n18621), .Z(n18623) );
  XNOR U22257 ( .A(b[464]), .B(n18621), .Z(n18622) );
  XOR U22258 ( .A(n18624), .B(n18625), .Z(n18621) );
  ANDN U22259 ( .B(n18626), .A(n602), .Z(n18624) );
  XNOR U22260 ( .A(a[463]), .B(n18627), .Z(n602) );
  IV U22261 ( .A(n18625), .Z(n18627) );
  XNOR U22262 ( .A(b[463]), .B(n18625), .Z(n18626) );
  XOR U22263 ( .A(n18628), .B(n18629), .Z(n18625) );
  ANDN U22264 ( .B(n18630), .A(n603), .Z(n18628) );
  XNOR U22265 ( .A(a[462]), .B(n18631), .Z(n603) );
  IV U22266 ( .A(n18629), .Z(n18631) );
  XNOR U22267 ( .A(b[462]), .B(n18629), .Z(n18630) );
  XOR U22268 ( .A(n18632), .B(n18633), .Z(n18629) );
  ANDN U22269 ( .B(n18634), .A(n604), .Z(n18632) );
  XNOR U22270 ( .A(a[461]), .B(n18635), .Z(n604) );
  IV U22271 ( .A(n18633), .Z(n18635) );
  XNOR U22272 ( .A(b[461]), .B(n18633), .Z(n18634) );
  XOR U22273 ( .A(n18636), .B(n18637), .Z(n18633) );
  ANDN U22274 ( .B(n18638), .A(n605), .Z(n18636) );
  XNOR U22275 ( .A(a[460]), .B(n18639), .Z(n605) );
  IV U22276 ( .A(n18637), .Z(n18639) );
  XNOR U22277 ( .A(b[460]), .B(n18637), .Z(n18638) );
  XOR U22278 ( .A(n18640), .B(n18641), .Z(n18637) );
  ANDN U22279 ( .B(n18642), .A(n607), .Z(n18640) );
  XNOR U22280 ( .A(a[459]), .B(n18643), .Z(n607) );
  IV U22281 ( .A(n18641), .Z(n18643) );
  XNOR U22282 ( .A(b[459]), .B(n18641), .Z(n18642) );
  XOR U22283 ( .A(n18644), .B(n18645), .Z(n18641) );
  ANDN U22284 ( .B(n18646), .A(n608), .Z(n18644) );
  XNOR U22285 ( .A(a[458]), .B(n18647), .Z(n608) );
  IV U22286 ( .A(n18645), .Z(n18647) );
  XNOR U22287 ( .A(b[458]), .B(n18645), .Z(n18646) );
  XOR U22288 ( .A(n18648), .B(n18649), .Z(n18645) );
  ANDN U22289 ( .B(n18650), .A(n609), .Z(n18648) );
  XNOR U22290 ( .A(a[457]), .B(n18651), .Z(n609) );
  IV U22291 ( .A(n18649), .Z(n18651) );
  XNOR U22292 ( .A(b[457]), .B(n18649), .Z(n18650) );
  XOR U22293 ( .A(n18652), .B(n18653), .Z(n18649) );
  ANDN U22294 ( .B(n18654), .A(n610), .Z(n18652) );
  XNOR U22295 ( .A(a[456]), .B(n18655), .Z(n610) );
  IV U22296 ( .A(n18653), .Z(n18655) );
  XNOR U22297 ( .A(b[456]), .B(n18653), .Z(n18654) );
  XOR U22298 ( .A(n18656), .B(n18657), .Z(n18653) );
  ANDN U22299 ( .B(n18658), .A(n611), .Z(n18656) );
  XNOR U22300 ( .A(a[455]), .B(n18659), .Z(n611) );
  IV U22301 ( .A(n18657), .Z(n18659) );
  XNOR U22302 ( .A(b[455]), .B(n18657), .Z(n18658) );
  XOR U22303 ( .A(n18660), .B(n18661), .Z(n18657) );
  ANDN U22304 ( .B(n18662), .A(n612), .Z(n18660) );
  XNOR U22305 ( .A(a[454]), .B(n18663), .Z(n612) );
  IV U22306 ( .A(n18661), .Z(n18663) );
  XNOR U22307 ( .A(b[454]), .B(n18661), .Z(n18662) );
  XOR U22308 ( .A(n18664), .B(n18665), .Z(n18661) );
  ANDN U22309 ( .B(n18666), .A(n613), .Z(n18664) );
  XNOR U22310 ( .A(a[453]), .B(n18667), .Z(n613) );
  IV U22311 ( .A(n18665), .Z(n18667) );
  XNOR U22312 ( .A(b[453]), .B(n18665), .Z(n18666) );
  XOR U22313 ( .A(n18668), .B(n18669), .Z(n18665) );
  ANDN U22314 ( .B(n18670), .A(n614), .Z(n18668) );
  XNOR U22315 ( .A(a[452]), .B(n18671), .Z(n614) );
  IV U22316 ( .A(n18669), .Z(n18671) );
  XNOR U22317 ( .A(b[452]), .B(n18669), .Z(n18670) );
  XOR U22318 ( .A(n18672), .B(n18673), .Z(n18669) );
  ANDN U22319 ( .B(n18674), .A(n615), .Z(n18672) );
  XNOR U22320 ( .A(a[451]), .B(n18675), .Z(n615) );
  IV U22321 ( .A(n18673), .Z(n18675) );
  XNOR U22322 ( .A(b[451]), .B(n18673), .Z(n18674) );
  XOR U22323 ( .A(n18676), .B(n18677), .Z(n18673) );
  ANDN U22324 ( .B(n18678), .A(n616), .Z(n18676) );
  XNOR U22325 ( .A(a[450]), .B(n18679), .Z(n616) );
  IV U22326 ( .A(n18677), .Z(n18679) );
  XNOR U22327 ( .A(b[450]), .B(n18677), .Z(n18678) );
  XOR U22328 ( .A(n18680), .B(n18681), .Z(n18677) );
  ANDN U22329 ( .B(n18682), .A(n618), .Z(n18680) );
  XNOR U22330 ( .A(a[449]), .B(n18683), .Z(n618) );
  IV U22331 ( .A(n18681), .Z(n18683) );
  XNOR U22332 ( .A(b[449]), .B(n18681), .Z(n18682) );
  XOR U22333 ( .A(n18684), .B(n18685), .Z(n18681) );
  ANDN U22334 ( .B(n18686), .A(n619), .Z(n18684) );
  XNOR U22335 ( .A(a[448]), .B(n18687), .Z(n619) );
  IV U22336 ( .A(n18685), .Z(n18687) );
  XNOR U22337 ( .A(b[448]), .B(n18685), .Z(n18686) );
  XOR U22338 ( .A(n18688), .B(n18689), .Z(n18685) );
  ANDN U22339 ( .B(n18690), .A(n620), .Z(n18688) );
  XNOR U22340 ( .A(a[447]), .B(n18691), .Z(n620) );
  IV U22341 ( .A(n18689), .Z(n18691) );
  XNOR U22342 ( .A(b[447]), .B(n18689), .Z(n18690) );
  XOR U22343 ( .A(n18692), .B(n18693), .Z(n18689) );
  ANDN U22344 ( .B(n18694), .A(n621), .Z(n18692) );
  XNOR U22345 ( .A(a[446]), .B(n18695), .Z(n621) );
  IV U22346 ( .A(n18693), .Z(n18695) );
  XNOR U22347 ( .A(b[446]), .B(n18693), .Z(n18694) );
  XOR U22348 ( .A(n18696), .B(n18697), .Z(n18693) );
  ANDN U22349 ( .B(n18698), .A(n622), .Z(n18696) );
  XNOR U22350 ( .A(a[445]), .B(n18699), .Z(n622) );
  IV U22351 ( .A(n18697), .Z(n18699) );
  XNOR U22352 ( .A(b[445]), .B(n18697), .Z(n18698) );
  XOR U22353 ( .A(n18700), .B(n18701), .Z(n18697) );
  ANDN U22354 ( .B(n18702), .A(n623), .Z(n18700) );
  XNOR U22355 ( .A(a[444]), .B(n18703), .Z(n623) );
  IV U22356 ( .A(n18701), .Z(n18703) );
  XNOR U22357 ( .A(b[444]), .B(n18701), .Z(n18702) );
  XOR U22358 ( .A(n18704), .B(n18705), .Z(n18701) );
  ANDN U22359 ( .B(n18706), .A(n624), .Z(n18704) );
  XNOR U22360 ( .A(a[443]), .B(n18707), .Z(n624) );
  IV U22361 ( .A(n18705), .Z(n18707) );
  XNOR U22362 ( .A(b[443]), .B(n18705), .Z(n18706) );
  XOR U22363 ( .A(n18708), .B(n18709), .Z(n18705) );
  ANDN U22364 ( .B(n18710), .A(n625), .Z(n18708) );
  XNOR U22365 ( .A(a[442]), .B(n18711), .Z(n625) );
  IV U22366 ( .A(n18709), .Z(n18711) );
  XNOR U22367 ( .A(b[442]), .B(n18709), .Z(n18710) );
  XOR U22368 ( .A(n18712), .B(n18713), .Z(n18709) );
  ANDN U22369 ( .B(n18714), .A(n626), .Z(n18712) );
  XNOR U22370 ( .A(a[441]), .B(n18715), .Z(n626) );
  IV U22371 ( .A(n18713), .Z(n18715) );
  XNOR U22372 ( .A(b[441]), .B(n18713), .Z(n18714) );
  XOR U22373 ( .A(n18716), .B(n18717), .Z(n18713) );
  ANDN U22374 ( .B(n18718), .A(n627), .Z(n18716) );
  XNOR U22375 ( .A(a[440]), .B(n18719), .Z(n627) );
  IV U22376 ( .A(n18717), .Z(n18719) );
  XNOR U22377 ( .A(b[440]), .B(n18717), .Z(n18718) );
  XOR U22378 ( .A(n18720), .B(n18721), .Z(n18717) );
  ANDN U22379 ( .B(n18722), .A(n629), .Z(n18720) );
  XNOR U22380 ( .A(a[439]), .B(n18723), .Z(n629) );
  IV U22381 ( .A(n18721), .Z(n18723) );
  XNOR U22382 ( .A(b[439]), .B(n18721), .Z(n18722) );
  XOR U22383 ( .A(n18724), .B(n18725), .Z(n18721) );
  ANDN U22384 ( .B(n18726), .A(n630), .Z(n18724) );
  XNOR U22385 ( .A(a[438]), .B(n18727), .Z(n630) );
  IV U22386 ( .A(n18725), .Z(n18727) );
  XNOR U22387 ( .A(b[438]), .B(n18725), .Z(n18726) );
  XOR U22388 ( .A(n18728), .B(n18729), .Z(n18725) );
  ANDN U22389 ( .B(n18730), .A(n631), .Z(n18728) );
  XNOR U22390 ( .A(a[437]), .B(n18731), .Z(n631) );
  IV U22391 ( .A(n18729), .Z(n18731) );
  XNOR U22392 ( .A(b[437]), .B(n18729), .Z(n18730) );
  XOR U22393 ( .A(n18732), .B(n18733), .Z(n18729) );
  ANDN U22394 ( .B(n18734), .A(n632), .Z(n18732) );
  XNOR U22395 ( .A(a[436]), .B(n18735), .Z(n632) );
  IV U22396 ( .A(n18733), .Z(n18735) );
  XNOR U22397 ( .A(b[436]), .B(n18733), .Z(n18734) );
  XOR U22398 ( .A(n18736), .B(n18737), .Z(n18733) );
  ANDN U22399 ( .B(n18738), .A(n633), .Z(n18736) );
  XNOR U22400 ( .A(a[435]), .B(n18739), .Z(n633) );
  IV U22401 ( .A(n18737), .Z(n18739) );
  XNOR U22402 ( .A(b[435]), .B(n18737), .Z(n18738) );
  XOR U22403 ( .A(n18740), .B(n18741), .Z(n18737) );
  ANDN U22404 ( .B(n18742), .A(n634), .Z(n18740) );
  XNOR U22405 ( .A(a[434]), .B(n18743), .Z(n634) );
  IV U22406 ( .A(n18741), .Z(n18743) );
  XNOR U22407 ( .A(b[434]), .B(n18741), .Z(n18742) );
  XOR U22408 ( .A(n18744), .B(n18745), .Z(n18741) );
  ANDN U22409 ( .B(n18746), .A(n635), .Z(n18744) );
  XNOR U22410 ( .A(a[433]), .B(n18747), .Z(n635) );
  IV U22411 ( .A(n18745), .Z(n18747) );
  XNOR U22412 ( .A(b[433]), .B(n18745), .Z(n18746) );
  XOR U22413 ( .A(n18748), .B(n18749), .Z(n18745) );
  ANDN U22414 ( .B(n18750), .A(n636), .Z(n18748) );
  XNOR U22415 ( .A(a[432]), .B(n18751), .Z(n636) );
  IV U22416 ( .A(n18749), .Z(n18751) );
  XNOR U22417 ( .A(b[432]), .B(n18749), .Z(n18750) );
  XOR U22418 ( .A(n18752), .B(n18753), .Z(n18749) );
  ANDN U22419 ( .B(n18754), .A(n637), .Z(n18752) );
  XNOR U22420 ( .A(a[431]), .B(n18755), .Z(n637) );
  IV U22421 ( .A(n18753), .Z(n18755) );
  XNOR U22422 ( .A(b[431]), .B(n18753), .Z(n18754) );
  XOR U22423 ( .A(n18756), .B(n18757), .Z(n18753) );
  ANDN U22424 ( .B(n18758), .A(n638), .Z(n18756) );
  XNOR U22425 ( .A(a[430]), .B(n18759), .Z(n638) );
  IV U22426 ( .A(n18757), .Z(n18759) );
  XNOR U22427 ( .A(b[430]), .B(n18757), .Z(n18758) );
  XOR U22428 ( .A(n18760), .B(n18761), .Z(n18757) );
  ANDN U22429 ( .B(n18762), .A(n640), .Z(n18760) );
  XNOR U22430 ( .A(a[429]), .B(n18763), .Z(n640) );
  IV U22431 ( .A(n18761), .Z(n18763) );
  XNOR U22432 ( .A(b[429]), .B(n18761), .Z(n18762) );
  XOR U22433 ( .A(n18764), .B(n18765), .Z(n18761) );
  ANDN U22434 ( .B(n18766), .A(n641), .Z(n18764) );
  XNOR U22435 ( .A(a[428]), .B(n18767), .Z(n641) );
  IV U22436 ( .A(n18765), .Z(n18767) );
  XNOR U22437 ( .A(b[428]), .B(n18765), .Z(n18766) );
  XOR U22438 ( .A(n18768), .B(n18769), .Z(n18765) );
  ANDN U22439 ( .B(n18770), .A(n642), .Z(n18768) );
  XNOR U22440 ( .A(a[427]), .B(n18771), .Z(n642) );
  IV U22441 ( .A(n18769), .Z(n18771) );
  XNOR U22442 ( .A(b[427]), .B(n18769), .Z(n18770) );
  XOR U22443 ( .A(n18772), .B(n18773), .Z(n18769) );
  ANDN U22444 ( .B(n18774), .A(n643), .Z(n18772) );
  XNOR U22445 ( .A(a[426]), .B(n18775), .Z(n643) );
  IV U22446 ( .A(n18773), .Z(n18775) );
  XNOR U22447 ( .A(b[426]), .B(n18773), .Z(n18774) );
  XOR U22448 ( .A(n18776), .B(n18777), .Z(n18773) );
  ANDN U22449 ( .B(n18778), .A(n644), .Z(n18776) );
  XNOR U22450 ( .A(a[425]), .B(n18779), .Z(n644) );
  IV U22451 ( .A(n18777), .Z(n18779) );
  XNOR U22452 ( .A(b[425]), .B(n18777), .Z(n18778) );
  XOR U22453 ( .A(n18780), .B(n18781), .Z(n18777) );
  ANDN U22454 ( .B(n18782), .A(n645), .Z(n18780) );
  XNOR U22455 ( .A(a[424]), .B(n18783), .Z(n645) );
  IV U22456 ( .A(n18781), .Z(n18783) );
  XNOR U22457 ( .A(b[424]), .B(n18781), .Z(n18782) );
  XOR U22458 ( .A(n18784), .B(n18785), .Z(n18781) );
  ANDN U22459 ( .B(n18786), .A(n646), .Z(n18784) );
  XNOR U22460 ( .A(a[423]), .B(n18787), .Z(n646) );
  IV U22461 ( .A(n18785), .Z(n18787) );
  XNOR U22462 ( .A(b[423]), .B(n18785), .Z(n18786) );
  XOR U22463 ( .A(n18788), .B(n18789), .Z(n18785) );
  ANDN U22464 ( .B(n18790), .A(n647), .Z(n18788) );
  XNOR U22465 ( .A(a[422]), .B(n18791), .Z(n647) );
  IV U22466 ( .A(n18789), .Z(n18791) );
  XNOR U22467 ( .A(b[422]), .B(n18789), .Z(n18790) );
  XOR U22468 ( .A(n18792), .B(n18793), .Z(n18789) );
  ANDN U22469 ( .B(n18794), .A(n648), .Z(n18792) );
  XNOR U22470 ( .A(a[421]), .B(n18795), .Z(n648) );
  IV U22471 ( .A(n18793), .Z(n18795) );
  XNOR U22472 ( .A(b[421]), .B(n18793), .Z(n18794) );
  XOR U22473 ( .A(n18796), .B(n18797), .Z(n18793) );
  ANDN U22474 ( .B(n18798), .A(n649), .Z(n18796) );
  XNOR U22475 ( .A(a[420]), .B(n18799), .Z(n649) );
  IV U22476 ( .A(n18797), .Z(n18799) );
  XNOR U22477 ( .A(b[420]), .B(n18797), .Z(n18798) );
  XOR U22478 ( .A(n18800), .B(n18801), .Z(n18797) );
  ANDN U22479 ( .B(n18802), .A(n651), .Z(n18800) );
  XNOR U22480 ( .A(a[419]), .B(n18803), .Z(n651) );
  IV U22481 ( .A(n18801), .Z(n18803) );
  XNOR U22482 ( .A(b[419]), .B(n18801), .Z(n18802) );
  XOR U22483 ( .A(n18804), .B(n18805), .Z(n18801) );
  ANDN U22484 ( .B(n18806), .A(n652), .Z(n18804) );
  XNOR U22485 ( .A(a[418]), .B(n18807), .Z(n652) );
  IV U22486 ( .A(n18805), .Z(n18807) );
  XNOR U22487 ( .A(b[418]), .B(n18805), .Z(n18806) );
  XOR U22488 ( .A(n18808), .B(n18809), .Z(n18805) );
  ANDN U22489 ( .B(n18810), .A(n653), .Z(n18808) );
  XNOR U22490 ( .A(a[417]), .B(n18811), .Z(n653) );
  IV U22491 ( .A(n18809), .Z(n18811) );
  XNOR U22492 ( .A(b[417]), .B(n18809), .Z(n18810) );
  XOR U22493 ( .A(n18812), .B(n18813), .Z(n18809) );
  ANDN U22494 ( .B(n18814), .A(n654), .Z(n18812) );
  XNOR U22495 ( .A(a[416]), .B(n18815), .Z(n654) );
  IV U22496 ( .A(n18813), .Z(n18815) );
  XNOR U22497 ( .A(b[416]), .B(n18813), .Z(n18814) );
  XOR U22498 ( .A(n18816), .B(n18817), .Z(n18813) );
  ANDN U22499 ( .B(n18818), .A(n655), .Z(n18816) );
  XNOR U22500 ( .A(a[415]), .B(n18819), .Z(n655) );
  IV U22501 ( .A(n18817), .Z(n18819) );
  XNOR U22502 ( .A(b[415]), .B(n18817), .Z(n18818) );
  XOR U22503 ( .A(n18820), .B(n18821), .Z(n18817) );
  ANDN U22504 ( .B(n18822), .A(n656), .Z(n18820) );
  XNOR U22505 ( .A(a[414]), .B(n18823), .Z(n656) );
  IV U22506 ( .A(n18821), .Z(n18823) );
  XNOR U22507 ( .A(b[414]), .B(n18821), .Z(n18822) );
  XOR U22508 ( .A(n18824), .B(n18825), .Z(n18821) );
  ANDN U22509 ( .B(n18826), .A(n657), .Z(n18824) );
  XNOR U22510 ( .A(a[413]), .B(n18827), .Z(n657) );
  IV U22511 ( .A(n18825), .Z(n18827) );
  XNOR U22512 ( .A(b[413]), .B(n18825), .Z(n18826) );
  XOR U22513 ( .A(n18828), .B(n18829), .Z(n18825) );
  ANDN U22514 ( .B(n18830), .A(n658), .Z(n18828) );
  XNOR U22515 ( .A(a[412]), .B(n18831), .Z(n658) );
  IV U22516 ( .A(n18829), .Z(n18831) );
  XNOR U22517 ( .A(b[412]), .B(n18829), .Z(n18830) );
  XOR U22518 ( .A(n18832), .B(n18833), .Z(n18829) );
  ANDN U22519 ( .B(n18834), .A(n659), .Z(n18832) );
  XNOR U22520 ( .A(a[411]), .B(n18835), .Z(n659) );
  IV U22521 ( .A(n18833), .Z(n18835) );
  XNOR U22522 ( .A(b[411]), .B(n18833), .Z(n18834) );
  XOR U22523 ( .A(n18836), .B(n18837), .Z(n18833) );
  ANDN U22524 ( .B(n18838), .A(n660), .Z(n18836) );
  XNOR U22525 ( .A(a[410]), .B(n18839), .Z(n660) );
  IV U22526 ( .A(n18837), .Z(n18839) );
  XNOR U22527 ( .A(b[410]), .B(n18837), .Z(n18838) );
  XOR U22528 ( .A(n18840), .B(n18841), .Z(n18837) );
  ANDN U22529 ( .B(n18842), .A(n662), .Z(n18840) );
  XNOR U22530 ( .A(a[409]), .B(n18843), .Z(n662) );
  IV U22531 ( .A(n18841), .Z(n18843) );
  XNOR U22532 ( .A(b[409]), .B(n18841), .Z(n18842) );
  XOR U22533 ( .A(n18844), .B(n18845), .Z(n18841) );
  ANDN U22534 ( .B(n18846), .A(n692), .Z(n18844) );
  XNOR U22535 ( .A(a[408]), .B(n18847), .Z(n692) );
  IV U22536 ( .A(n18845), .Z(n18847) );
  XNOR U22537 ( .A(b[408]), .B(n18845), .Z(n18846) );
  XOR U22538 ( .A(n18848), .B(n18849), .Z(n18845) );
  ANDN U22539 ( .B(n18850), .A(n743), .Z(n18848) );
  XNOR U22540 ( .A(a[407]), .B(n18851), .Z(n743) );
  IV U22541 ( .A(n18849), .Z(n18851) );
  XNOR U22542 ( .A(b[407]), .B(n18849), .Z(n18850) );
  XOR U22543 ( .A(n18852), .B(n18853), .Z(n18849) );
  ANDN U22544 ( .B(n18854), .A(n794), .Z(n18852) );
  XNOR U22545 ( .A(a[406]), .B(n18855), .Z(n794) );
  IV U22546 ( .A(n18853), .Z(n18855) );
  XNOR U22547 ( .A(b[406]), .B(n18853), .Z(n18854) );
  XOR U22548 ( .A(n18856), .B(n18857), .Z(n18853) );
  ANDN U22549 ( .B(n18858), .A(n845), .Z(n18856) );
  XNOR U22550 ( .A(a[405]), .B(n18859), .Z(n845) );
  IV U22551 ( .A(n18857), .Z(n18859) );
  XNOR U22552 ( .A(b[405]), .B(n18857), .Z(n18858) );
  XOR U22553 ( .A(n18860), .B(n18861), .Z(n18857) );
  ANDN U22554 ( .B(n18862), .A(n896), .Z(n18860) );
  XNOR U22555 ( .A(a[404]), .B(n18863), .Z(n896) );
  IV U22556 ( .A(n18861), .Z(n18863) );
  XNOR U22557 ( .A(b[404]), .B(n18861), .Z(n18862) );
  XOR U22558 ( .A(n18864), .B(n18865), .Z(n18861) );
  ANDN U22559 ( .B(n18866), .A(n947), .Z(n18864) );
  XNOR U22560 ( .A(a[403]), .B(n18867), .Z(n947) );
  IV U22561 ( .A(n18865), .Z(n18867) );
  XNOR U22562 ( .A(b[403]), .B(n18865), .Z(n18866) );
  XOR U22563 ( .A(n18868), .B(n18869), .Z(n18865) );
  ANDN U22564 ( .B(n18870), .A(n998), .Z(n18868) );
  XNOR U22565 ( .A(a[402]), .B(n18871), .Z(n998) );
  IV U22566 ( .A(n18869), .Z(n18871) );
  XNOR U22567 ( .A(b[402]), .B(n18869), .Z(n18870) );
  XOR U22568 ( .A(n18872), .B(n18873), .Z(n18869) );
  ANDN U22569 ( .B(n18874), .A(n1049), .Z(n18872) );
  XNOR U22570 ( .A(a[401]), .B(n18875), .Z(n1049) );
  IV U22571 ( .A(n18873), .Z(n18875) );
  XNOR U22572 ( .A(b[401]), .B(n18873), .Z(n18874) );
  XOR U22573 ( .A(n18876), .B(n18877), .Z(n18873) );
  ANDN U22574 ( .B(n18878), .A(n1100), .Z(n18876) );
  XNOR U22575 ( .A(a[400]), .B(n18879), .Z(n1100) );
  IV U22576 ( .A(n18877), .Z(n18879) );
  XNOR U22577 ( .A(b[400]), .B(n18877), .Z(n18878) );
  XOR U22578 ( .A(n18880), .B(n18881), .Z(n18877) );
  ANDN U22579 ( .B(n18882), .A(n1153), .Z(n18880) );
  XNOR U22580 ( .A(a[399]), .B(n18883), .Z(n1153) );
  IV U22581 ( .A(n18881), .Z(n18883) );
  XNOR U22582 ( .A(b[399]), .B(n18881), .Z(n18882) );
  XOR U22583 ( .A(n18884), .B(n18885), .Z(n18881) );
  ANDN U22584 ( .B(n18886), .A(n1204), .Z(n18884) );
  XNOR U22585 ( .A(a[398]), .B(n18887), .Z(n1204) );
  IV U22586 ( .A(n18885), .Z(n18887) );
  XNOR U22587 ( .A(b[398]), .B(n18885), .Z(n18886) );
  XOR U22588 ( .A(n18888), .B(n18889), .Z(n18885) );
  ANDN U22589 ( .B(n18890), .A(n1255), .Z(n18888) );
  XNOR U22590 ( .A(a[397]), .B(n18891), .Z(n1255) );
  IV U22591 ( .A(n18889), .Z(n18891) );
  XNOR U22592 ( .A(b[397]), .B(n18889), .Z(n18890) );
  XOR U22593 ( .A(n18892), .B(n18893), .Z(n18889) );
  ANDN U22594 ( .B(n18894), .A(n1306), .Z(n18892) );
  XNOR U22595 ( .A(a[396]), .B(n18895), .Z(n1306) );
  IV U22596 ( .A(n18893), .Z(n18895) );
  XNOR U22597 ( .A(b[396]), .B(n18893), .Z(n18894) );
  XOR U22598 ( .A(n18896), .B(n18897), .Z(n18893) );
  ANDN U22599 ( .B(n18898), .A(n1357), .Z(n18896) );
  XNOR U22600 ( .A(a[395]), .B(n18899), .Z(n1357) );
  IV U22601 ( .A(n18897), .Z(n18899) );
  XNOR U22602 ( .A(b[395]), .B(n18897), .Z(n18898) );
  XOR U22603 ( .A(n18900), .B(n18901), .Z(n18897) );
  ANDN U22604 ( .B(n18902), .A(n1408), .Z(n18900) );
  XNOR U22605 ( .A(a[394]), .B(n18903), .Z(n1408) );
  IV U22606 ( .A(n18901), .Z(n18903) );
  XNOR U22607 ( .A(b[394]), .B(n18901), .Z(n18902) );
  XOR U22608 ( .A(n18904), .B(n18905), .Z(n18901) );
  ANDN U22609 ( .B(n18906), .A(n1459), .Z(n18904) );
  XNOR U22610 ( .A(a[393]), .B(n18907), .Z(n1459) );
  IV U22611 ( .A(n18905), .Z(n18907) );
  XNOR U22612 ( .A(b[393]), .B(n18905), .Z(n18906) );
  XOR U22613 ( .A(n18908), .B(n18909), .Z(n18905) );
  ANDN U22614 ( .B(n18910), .A(n1510), .Z(n18908) );
  XNOR U22615 ( .A(a[392]), .B(n18911), .Z(n1510) );
  IV U22616 ( .A(n18909), .Z(n18911) );
  XNOR U22617 ( .A(b[392]), .B(n18909), .Z(n18910) );
  XOR U22618 ( .A(n18912), .B(n18913), .Z(n18909) );
  ANDN U22619 ( .B(n18914), .A(n1561), .Z(n18912) );
  XNOR U22620 ( .A(a[391]), .B(n18915), .Z(n1561) );
  IV U22621 ( .A(n18913), .Z(n18915) );
  XNOR U22622 ( .A(b[391]), .B(n18913), .Z(n18914) );
  XOR U22623 ( .A(n18916), .B(n18917), .Z(n18913) );
  ANDN U22624 ( .B(n18918), .A(n1612), .Z(n18916) );
  XNOR U22625 ( .A(a[390]), .B(n18919), .Z(n1612) );
  IV U22626 ( .A(n18917), .Z(n18919) );
  XNOR U22627 ( .A(b[390]), .B(n18917), .Z(n18918) );
  XOR U22628 ( .A(n18920), .B(n18921), .Z(n18917) );
  ANDN U22629 ( .B(n18922), .A(n1664), .Z(n18920) );
  XNOR U22630 ( .A(a[389]), .B(n18923), .Z(n1664) );
  IV U22631 ( .A(n18921), .Z(n18923) );
  XNOR U22632 ( .A(b[389]), .B(n18921), .Z(n18922) );
  XOR U22633 ( .A(n18924), .B(n18925), .Z(n18921) );
  ANDN U22634 ( .B(n18926), .A(n1715), .Z(n18924) );
  XNOR U22635 ( .A(a[388]), .B(n18927), .Z(n1715) );
  IV U22636 ( .A(n18925), .Z(n18927) );
  XNOR U22637 ( .A(b[388]), .B(n18925), .Z(n18926) );
  XOR U22638 ( .A(n18928), .B(n18929), .Z(n18925) );
  ANDN U22639 ( .B(n18930), .A(n1766), .Z(n18928) );
  XNOR U22640 ( .A(a[387]), .B(n18931), .Z(n1766) );
  IV U22641 ( .A(n18929), .Z(n18931) );
  XNOR U22642 ( .A(b[387]), .B(n18929), .Z(n18930) );
  XOR U22643 ( .A(n18932), .B(n18933), .Z(n18929) );
  ANDN U22644 ( .B(n18934), .A(n1817), .Z(n18932) );
  XNOR U22645 ( .A(a[386]), .B(n18935), .Z(n1817) );
  IV U22646 ( .A(n18933), .Z(n18935) );
  XNOR U22647 ( .A(b[386]), .B(n18933), .Z(n18934) );
  XOR U22648 ( .A(n18936), .B(n18937), .Z(n18933) );
  ANDN U22649 ( .B(n18938), .A(n1868), .Z(n18936) );
  XNOR U22650 ( .A(a[385]), .B(n18939), .Z(n1868) );
  IV U22651 ( .A(n18937), .Z(n18939) );
  XNOR U22652 ( .A(b[385]), .B(n18937), .Z(n18938) );
  XOR U22653 ( .A(n18940), .B(n18941), .Z(n18937) );
  ANDN U22654 ( .B(n18942), .A(n1919), .Z(n18940) );
  XNOR U22655 ( .A(a[384]), .B(n18943), .Z(n1919) );
  IV U22656 ( .A(n18941), .Z(n18943) );
  XNOR U22657 ( .A(b[384]), .B(n18941), .Z(n18942) );
  XOR U22658 ( .A(n18944), .B(n18945), .Z(n18941) );
  ANDN U22659 ( .B(n18946), .A(n1970), .Z(n18944) );
  XNOR U22660 ( .A(a[383]), .B(n18947), .Z(n1970) );
  IV U22661 ( .A(n18945), .Z(n18947) );
  XNOR U22662 ( .A(b[383]), .B(n18945), .Z(n18946) );
  XOR U22663 ( .A(n18948), .B(n18949), .Z(n18945) );
  ANDN U22664 ( .B(n18950), .A(n2021), .Z(n18948) );
  XNOR U22665 ( .A(a[382]), .B(n18951), .Z(n2021) );
  IV U22666 ( .A(n18949), .Z(n18951) );
  XNOR U22667 ( .A(b[382]), .B(n18949), .Z(n18950) );
  XOR U22668 ( .A(n18952), .B(n18953), .Z(n18949) );
  ANDN U22669 ( .B(n18954), .A(n2072), .Z(n18952) );
  XNOR U22670 ( .A(a[381]), .B(n18955), .Z(n2072) );
  IV U22671 ( .A(n18953), .Z(n18955) );
  XNOR U22672 ( .A(b[381]), .B(n18953), .Z(n18954) );
  XOR U22673 ( .A(n18956), .B(n18957), .Z(n18953) );
  ANDN U22674 ( .B(n18958), .A(n2123), .Z(n18956) );
  XNOR U22675 ( .A(a[380]), .B(n18959), .Z(n2123) );
  IV U22676 ( .A(n18957), .Z(n18959) );
  XNOR U22677 ( .A(b[380]), .B(n18957), .Z(n18958) );
  XOR U22678 ( .A(n18960), .B(n18961), .Z(n18957) );
  ANDN U22679 ( .B(n18962), .A(n2175), .Z(n18960) );
  XNOR U22680 ( .A(a[379]), .B(n18963), .Z(n2175) );
  IV U22681 ( .A(n18961), .Z(n18963) );
  XNOR U22682 ( .A(b[379]), .B(n18961), .Z(n18962) );
  XOR U22683 ( .A(n18964), .B(n18965), .Z(n18961) );
  ANDN U22684 ( .B(n18966), .A(n2226), .Z(n18964) );
  XNOR U22685 ( .A(a[378]), .B(n18967), .Z(n2226) );
  IV U22686 ( .A(n18965), .Z(n18967) );
  XNOR U22687 ( .A(b[378]), .B(n18965), .Z(n18966) );
  XOR U22688 ( .A(n18968), .B(n18969), .Z(n18965) );
  ANDN U22689 ( .B(n18970), .A(n2277), .Z(n18968) );
  XNOR U22690 ( .A(a[377]), .B(n18971), .Z(n2277) );
  IV U22691 ( .A(n18969), .Z(n18971) );
  XNOR U22692 ( .A(b[377]), .B(n18969), .Z(n18970) );
  XOR U22693 ( .A(n18972), .B(n18973), .Z(n18969) );
  ANDN U22694 ( .B(n18974), .A(n2328), .Z(n18972) );
  XNOR U22695 ( .A(a[376]), .B(n18975), .Z(n2328) );
  IV U22696 ( .A(n18973), .Z(n18975) );
  XNOR U22697 ( .A(b[376]), .B(n18973), .Z(n18974) );
  XOR U22698 ( .A(n18976), .B(n18977), .Z(n18973) );
  ANDN U22699 ( .B(n18978), .A(n2379), .Z(n18976) );
  XNOR U22700 ( .A(a[375]), .B(n18979), .Z(n2379) );
  IV U22701 ( .A(n18977), .Z(n18979) );
  XNOR U22702 ( .A(b[375]), .B(n18977), .Z(n18978) );
  XOR U22703 ( .A(n18980), .B(n18981), .Z(n18977) );
  ANDN U22704 ( .B(n18982), .A(n2430), .Z(n18980) );
  XNOR U22705 ( .A(a[374]), .B(n18983), .Z(n2430) );
  IV U22706 ( .A(n18981), .Z(n18983) );
  XNOR U22707 ( .A(b[374]), .B(n18981), .Z(n18982) );
  XOR U22708 ( .A(n18984), .B(n18985), .Z(n18981) );
  ANDN U22709 ( .B(n18986), .A(n2481), .Z(n18984) );
  XNOR U22710 ( .A(a[373]), .B(n18987), .Z(n2481) );
  IV U22711 ( .A(n18985), .Z(n18987) );
  XNOR U22712 ( .A(b[373]), .B(n18985), .Z(n18986) );
  XOR U22713 ( .A(n18988), .B(n18989), .Z(n18985) );
  ANDN U22714 ( .B(n18990), .A(n2532), .Z(n18988) );
  XNOR U22715 ( .A(a[372]), .B(n18991), .Z(n2532) );
  IV U22716 ( .A(n18989), .Z(n18991) );
  XNOR U22717 ( .A(b[372]), .B(n18989), .Z(n18990) );
  XOR U22718 ( .A(n18992), .B(n18993), .Z(n18989) );
  ANDN U22719 ( .B(n18994), .A(n2583), .Z(n18992) );
  XNOR U22720 ( .A(a[371]), .B(n18995), .Z(n2583) );
  IV U22721 ( .A(n18993), .Z(n18995) );
  XNOR U22722 ( .A(b[371]), .B(n18993), .Z(n18994) );
  XOR U22723 ( .A(n18996), .B(n18997), .Z(n18993) );
  ANDN U22724 ( .B(n18998), .A(n2634), .Z(n18996) );
  XNOR U22725 ( .A(a[370]), .B(n18999), .Z(n2634) );
  IV U22726 ( .A(n18997), .Z(n18999) );
  XNOR U22727 ( .A(b[370]), .B(n18997), .Z(n18998) );
  XOR U22728 ( .A(n19000), .B(n19001), .Z(n18997) );
  ANDN U22729 ( .B(n19002), .A(n2686), .Z(n19000) );
  XNOR U22730 ( .A(a[369]), .B(n19003), .Z(n2686) );
  IV U22731 ( .A(n19001), .Z(n19003) );
  XNOR U22732 ( .A(b[369]), .B(n19001), .Z(n19002) );
  XOR U22733 ( .A(n19004), .B(n19005), .Z(n19001) );
  ANDN U22734 ( .B(n19006), .A(n2737), .Z(n19004) );
  XNOR U22735 ( .A(a[368]), .B(n19007), .Z(n2737) );
  IV U22736 ( .A(n19005), .Z(n19007) );
  XNOR U22737 ( .A(b[368]), .B(n19005), .Z(n19006) );
  XOR U22738 ( .A(n19008), .B(n19009), .Z(n19005) );
  ANDN U22739 ( .B(n19010), .A(n2788), .Z(n19008) );
  XNOR U22740 ( .A(a[367]), .B(n19011), .Z(n2788) );
  IV U22741 ( .A(n19009), .Z(n19011) );
  XNOR U22742 ( .A(b[367]), .B(n19009), .Z(n19010) );
  XOR U22743 ( .A(n19012), .B(n19013), .Z(n19009) );
  ANDN U22744 ( .B(n19014), .A(n2839), .Z(n19012) );
  XNOR U22745 ( .A(a[366]), .B(n19015), .Z(n2839) );
  IV U22746 ( .A(n19013), .Z(n19015) );
  XNOR U22747 ( .A(b[366]), .B(n19013), .Z(n19014) );
  XOR U22748 ( .A(n19016), .B(n19017), .Z(n19013) );
  ANDN U22749 ( .B(n19018), .A(n2890), .Z(n19016) );
  XNOR U22750 ( .A(a[365]), .B(n19019), .Z(n2890) );
  IV U22751 ( .A(n19017), .Z(n19019) );
  XNOR U22752 ( .A(b[365]), .B(n19017), .Z(n19018) );
  XOR U22753 ( .A(n19020), .B(n19021), .Z(n19017) );
  ANDN U22754 ( .B(n19022), .A(n2941), .Z(n19020) );
  XNOR U22755 ( .A(a[364]), .B(n19023), .Z(n2941) );
  IV U22756 ( .A(n19021), .Z(n19023) );
  XNOR U22757 ( .A(b[364]), .B(n19021), .Z(n19022) );
  XOR U22758 ( .A(n19024), .B(n19025), .Z(n19021) );
  ANDN U22759 ( .B(n19026), .A(n2992), .Z(n19024) );
  XNOR U22760 ( .A(a[363]), .B(n19027), .Z(n2992) );
  IV U22761 ( .A(n19025), .Z(n19027) );
  XNOR U22762 ( .A(b[363]), .B(n19025), .Z(n19026) );
  XOR U22763 ( .A(n19028), .B(n19029), .Z(n19025) );
  ANDN U22764 ( .B(n19030), .A(n3043), .Z(n19028) );
  XNOR U22765 ( .A(a[362]), .B(n19031), .Z(n3043) );
  IV U22766 ( .A(n19029), .Z(n19031) );
  XNOR U22767 ( .A(b[362]), .B(n19029), .Z(n19030) );
  XOR U22768 ( .A(n19032), .B(n19033), .Z(n19029) );
  ANDN U22769 ( .B(n19034), .A(n3094), .Z(n19032) );
  XNOR U22770 ( .A(a[361]), .B(n19035), .Z(n3094) );
  IV U22771 ( .A(n19033), .Z(n19035) );
  XNOR U22772 ( .A(b[361]), .B(n19033), .Z(n19034) );
  XOR U22773 ( .A(n19036), .B(n19037), .Z(n19033) );
  ANDN U22774 ( .B(n19038), .A(n3145), .Z(n19036) );
  XNOR U22775 ( .A(a[360]), .B(n19039), .Z(n3145) );
  IV U22776 ( .A(n19037), .Z(n19039) );
  XNOR U22777 ( .A(b[360]), .B(n19037), .Z(n19038) );
  XOR U22778 ( .A(n19040), .B(n19041), .Z(n19037) );
  ANDN U22779 ( .B(n19042), .A(n3197), .Z(n19040) );
  XNOR U22780 ( .A(a[359]), .B(n19043), .Z(n3197) );
  IV U22781 ( .A(n19041), .Z(n19043) );
  XNOR U22782 ( .A(b[359]), .B(n19041), .Z(n19042) );
  XOR U22783 ( .A(n19044), .B(n19045), .Z(n19041) );
  ANDN U22784 ( .B(n19046), .A(n3248), .Z(n19044) );
  XNOR U22785 ( .A(a[358]), .B(n19047), .Z(n3248) );
  IV U22786 ( .A(n19045), .Z(n19047) );
  XNOR U22787 ( .A(b[358]), .B(n19045), .Z(n19046) );
  XOR U22788 ( .A(n19048), .B(n19049), .Z(n19045) );
  ANDN U22789 ( .B(n19050), .A(n3299), .Z(n19048) );
  XNOR U22790 ( .A(a[357]), .B(n19051), .Z(n3299) );
  IV U22791 ( .A(n19049), .Z(n19051) );
  XNOR U22792 ( .A(b[357]), .B(n19049), .Z(n19050) );
  XOR U22793 ( .A(n19052), .B(n19053), .Z(n19049) );
  ANDN U22794 ( .B(n19054), .A(n3350), .Z(n19052) );
  XNOR U22795 ( .A(a[356]), .B(n19055), .Z(n3350) );
  IV U22796 ( .A(n19053), .Z(n19055) );
  XNOR U22797 ( .A(b[356]), .B(n19053), .Z(n19054) );
  XOR U22798 ( .A(n19056), .B(n19057), .Z(n19053) );
  ANDN U22799 ( .B(n19058), .A(n3401), .Z(n19056) );
  XNOR U22800 ( .A(a[355]), .B(n19059), .Z(n3401) );
  IV U22801 ( .A(n19057), .Z(n19059) );
  XNOR U22802 ( .A(b[355]), .B(n19057), .Z(n19058) );
  XOR U22803 ( .A(n19060), .B(n19061), .Z(n19057) );
  ANDN U22804 ( .B(n19062), .A(n3452), .Z(n19060) );
  XNOR U22805 ( .A(a[354]), .B(n19063), .Z(n3452) );
  IV U22806 ( .A(n19061), .Z(n19063) );
  XNOR U22807 ( .A(b[354]), .B(n19061), .Z(n19062) );
  XOR U22808 ( .A(n19064), .B(n19065), .Z(n19061) );
  ANDN U22809 ( .B(n19066), .A(n3503), .Z(n19064) );
  XNOR U22810 ( .A(a[353]), .B(n19067), .Z(n3503) );
  IV U22811 ( .A(n19065), .Z(n19067) );
  XNOR U22812 ( .A(b[353]), .B(n19065), .Z(n19066) );
  XOR U22813 ( .A(n19068), .B(n19069), .Z(n19065) );
  ANDN U22814 ( .B(n19070), .A(n3554), .Z(n19068) );
  XNOR U22815 ( .A(a[352]), .B(n19071), .Z(n3554) );
  IV U22816 ( .A(n19069), .Z(n19071) );
  XNOR U22817 ( .A(b[352]), .B(n19069), .Z(n19070) );
  XOR U22818 ( .A(n19072), .B(n19073), .Z(n19069) );
  ANDN U22819 ( .B(n19074), .A(n3605), .Z(n19072) );
  XNOR U22820 ( .A(a[351]), .B(n19075), .Z(n3605) );
  IV U22821 ( .A(n19073), .Z(n19075) );
  XNOR U22822 ( .A(b[351]), .B(n19073), .Z(n19074) );
  XOR U22823 ( .A(n19076), .B(n19077), .Z(n19073) );
  ANDN U22824 ( .B(n19078), .A(n3656), .Z(n19076) );
  XNOR U22825 ( .A(a[350]), .B(n19079), .Z(n3656) );
  IV U22826 ( .A(n19077), .Z(n19079) );
  XNOR U22827 ( .A(b[350]), .B(n19077), .Z(n19078) );
  XOR U22828 ( .A(n19080), .B(n19081), .Z(n19077) );
  ANDN U22829 ( .B(n19082), .A(n3708), .Z(n19080) );
  XNOR U22830 ( .A(a[349]), .B(n19083), .Z(n3708) );
  IV U22831 ( .A(n19081), .Z(n19083) );
  XNOR U22832 ( .A(b[349]), .B(n19081), .Z(n19082) );
  XOR U22833 ( .A(n19084), .B(n19085), .Z(n19081) );
  ANDN U22834 ( .B(n19086), .A(n3759), .Z(n19084) );
  XNOR U22835 ( .A(a[348]), .B(n19087), .Z(n3759) );
  IV U22836 ( .A(n19085), .Z(n19087) );
  XNOR U22837 ( .A(b[348]), .B(n19085), .Z(n19086) );
  XOR U22838 ( .A(n19088), .B(n19089), .Z(n19085) );
  ANDN U22839 ( .B(n19090), .A(n3810), .Z(n19088) );
  XNOR U22840 ( .A(a[347]), .B(n19091), .Z(n3810) );
  IV U22841 ( .A(n19089), .Z(n19091) );
  XNOR U22842 ( .A(b[347]), .B(n19089), .Z(n19090) );
  XOR U22843 ( .A(n19092), .B(n19093), .Z(n19089) );
  ANDN U22844 ( .B(n19094), .A(n3861), .Z(n19092) );
  XNOR U22845 ( .A(a[346]), .B(n19095), .Z(n3861) );
  IV U22846 ( .A(n19093), .Z(n19095) );
  XNOR U22847 ( .A(b[346]), .B(n19093), .Z(n19094) );
  XOR U22848 ( .A(n19096), .B(n19097), .Z(n19093) );
  ANDN U22849 ( .B(n19098), .A(n3912), .Z(n19096) );
  XNOR U22850 ( .A(a[345]), .B(n19099), .Z(n3912) );
  IV U22851 ( .A(n19097), .Z(n19099) );
  XNOR U22852 ( .A(b[345]), .B(n19097), .Z(n19098) );
  XOR U22853 ( .A(n19100), .B(n19101), .Z(n19097) );
  ANDN U22854 ( .B(n19102), .A(n3963), .Z(n19100) );
  XNOR U22855 ( .A(a[344]), .B(n19103), .Z(n3963) );
  IV U22856 ( .A(n19101), .Z(n19103) );
  XNOR U22857 ( .A(b[344]), .B(n19101), .Z(n19102) );
  XOR U22858 ( .A(n19104), .B(n19105), .Z(n19101) );
  ANDN U22859 ( .B(n19106), .A(n4014), .Z(n19104) );
  XNOR U22860 ( .A(a[343]), .B(n19107), .Z(n4014) );
  IV U22861 ( .A(n19105), .Z(n19107) );
  XNOR U22862 ( .A(b[343]), .B(n19105), .Z(n19106) );
  XOR U22863 ( .A(n19108), .B(n19109), .Z(n19105) );
  ANDN U22864 ( .B(n19110), .A(n4065), .Z(n19108) );
  XNOR U22865 ( .A(a[342]), .B(n19111), .Z(n4065) );
  IV U22866 ( .A(n19109), .Z(n19111) );
  XNOR U22867 ( .A(b[342]), .B(n19109), .Z(n19110) );
  XOR U22868 ( .A(n19112), .B(n19113), .Z(n19109) );
  ANDN U22869 ( .B(n19114), .A(n4116), .Z(n19112) );
  XNOR U22870 ( .A(a[341]), .B(n19115), .Z(n4116) );
  IV U22871 ( .A(n19113), .Z(n19115) );
  XNOR U22872 ( .A(b[341]), .B(n19113), .Z(n19114) );
  XOR U22873 ( .A(n19116), .B(n19117), .Z(n19113) );
  ANDN U22874 ( .B(n19118), .A(n4167), .Z(n19116) );
  XNOR U22875 ( .A(a[340]), .B(n19119), .Z(n4167) );
  IV U22876 ( .A(n19117), .Z(n19119) );
  XNOR U22877 ( .A(b[340]), .B(n19117), .Z(n19118) );
  XOR U22878 ( .A(n19120), .B(n19121), .Z(n19117) );
  ANDN U22879 ( .B(n19122), .A(n4219), .Z(n19120) );
  XNOR U22880 ( .A(a[339]), .B(n19123), .Z(n4219) );
  IV U22881 ( .A(n19121), .Z(n19123) );
  XNOR U22882 ( .A(b[339]), .B(n19121), .Z(n19122) );
  XOR U22883 ( .A(n19124), .B(n19125), .Z(n19121) );
  ANDN U22884 ( .B(n19126), .A(n4270), .Z(n19124) );
  XNOR U22885 ( .A(a[338]), .B(n19127), .Z(n4270) );
  IV U22886 ( .A(n19125), .Z(n19127) );
  XNOR U22887 ( .A(b[338]), .B(n19125), .Z(n19126) );
  XOR U22888 ( .A(n19128), .B(n19129), .Z(n19125) );
  ANDN U22889 ( .B(n19130), .A(n4321), .Z(n19128) );
  XNOR U22890 ( .A(a[337]), .B(n19131), .Z(n4321) );
  IV U22891 ( .A(n19129), .Z(n19131) );
  XNOR U22892 ( .A(b[337]), .B(n19129), .Z(n19130) );
  XOR U22893 ( .A(n19132), .B(n19133), .Z(n19129) );
  ANDN U22894 ( .B(n19134), .A(n4372), .Z(n19132) );
  XNOR U22895 ( .A(a[336]), .B(n19135), .Z(n4372) );
  IV U22896 ( .A(n19133), .Z(n19135) );
  XNOR U22897 ( .A(b[336]), .B(n19133), .Z(n19134) );
  XOR U22898 ( .A(n19136), .B(n19137), .Z(n19133) );
  ANDN U22899 ( .B(n19138), .A(n4423), .Z(n19136) );
  XNOR U22900 ( .A(a[335]), .B(n19139), .Z(n4423) );
  IV U22901 ( .A(n19137), .Z(n19139) );
  XNOR U22902 ( .A(b[335]), .B(n19137), .Z(n19138) );
  XOR U22903 ( .A(n19140), .B(n19141), .Z(n19137) );
  ANDN U22904 ( .B(n19142), .A(n4474), .Z(n19140) );
  XNOR U22905 ( .A(a[334]), .B(n19143), .Z(n4474) );
  IV U22906 ( .A(n19141), .Z(n19143) );
  XNOR U22907 ( .A(b[334]), .B(n19141), .Z(n19142) );
  XOR U22908 ( .A(n19144), .B(n19145), .Z(n19141) );
  ANDN U22909 ( .B(n19146), .A(n4525), .Z(n19144) );
  XNOR U22910 ( .A(a[333]), .B(n19147), .Z(n4525) );
  IV U22911 ( .A(n19145), .Z(n19147) );
  XNOR U22912 ( .A(b[333]), .B(n19145), .Z(n19146) );
  XOR U22913 ( .A(n19148), .B(n19149), .Z(n19145) );
  ANDN U22914 ( .B(n19150), .A(n4576), .Z(n19148) );
  XNOR U22915 ( .A(a[332]), .B(n19151), .Z(n4576) );
  IV U22916 ( .A(n19149), .Z(n19151) );
  XNOR U22917 ( .A(b[332]), .B(n19149), .Z(n19150) );
  XOR U22918 ( .A(n19152), .B(n19153), .Z(n19149) );
  ANDN U22919 ( .B(n19154), .A(n4627), .Z(n19152) );
  XNOR U22920 ( .A(a[331]), .B(n19155), .Z(n4627) );
  IV U22921 ( .A(n19153), .Z(n19155) );
  XNOR U22922 ( .A(b[331]), .B(n19153), .Z(n19154) );
  XOR U22923 ( .A(n19156), .B(n19157), .Z(n19153) );
  ANDN U22924 ( .B(n19158), .A(n4678), .Z(n19156) );
  XNOR U22925 ( .A(a[330]), .B(n19159), .Z(n4678) );
  IV U22926 ( .A(n19157), .Z(n19159) );
  XNOR U22927 ( .A(b[330]), .B(n19157), .Z(n19158) );
  XOR U22928 ( .A(n19160), .B(n19161), .Z(n19157) );
  ANDN U22929 ( .B(n19162), .A(n4730), .Z(n19160) );
  XNOR U22930 ( .A(a[329]), .B(n19163), .Z(n4730) );
  IV U22931 ( .A(n19161), .Z(n19163) );
  XNOR U22932 ( .A(b[329]), .B(n19161), .Z(n19162) );
  XOR U22933 ( .A(n19164), .B(n19165), .Z(n19161) );
  ANDN U22934 ( .B(n19166), .A(n4781), .Z(n19164) );
  XNOR U22935 ( .A(a[328]), .B(n19167), .Z(n4781) );
  IV U22936 ( .A(n19165), .Z(n19167) );
  XNOR U22937 ( .A(b[328]), .B(n19165), .Z(n19166) );
  XOR U22938 ( .A(n19168), .B(n19169), .Z(n19165) );
  ANDN U22939 ( .B(n19170), .A(n4832), .Z(n19168) );
  XNOR U22940 ( .A(a[327]), .B(n19171), .Z(n4832) );
  IV U22941 ( .A(n19169), .Z(n19171) );
  XNOR U22942 ( .A(b[327]), .B(n19169), .Z(n19170) );
  XOR U22943 ( .A(n19172), .B(n19173), .Z(n19169) );
  ANDN U22944 ( .B(n19174), .A(n4883), .Z(n19172) );
  XNOR U22945 ( .A(a[326]), .B(n19175), .Z(n4883) );
  IV U22946 ( .A(n19173), .Z(n19175) );
  XNOR U22947 ( .A(b[326]), .B(n19173), .Z(n19174) );
  XOR U22948 ( .A(n19176), .B(n19177), .Z(n19173) );
  ANDN U22949 ( .B(n19178), .A(n4934), .Z(n19176) );
  XNOR U22950 ( .A(a[325]), .B(n19179), .Z(n4934) );
  IV U22951 ( .A(n19177), .Z(n19179) );
  XNOR U22952 ( .A(b[325]), .B(n19177), .Z(n19178) );
  XOR U22953 ( .A(n19180), .B(n19181), .Z(n19177) );
  ANDN U22954 ( .B(n19182), .A(n4985), .Z(n19180) );
  XNOR U22955 ( .A(a[324]), .B(n19183), .Z(n4985) );
  IV U22956 ( .A(n19181), .Z(n19183) );
  XNOR U22957 ( .A(b[324]), .B(n19181), .Z(n19182) );
  XOR U22958 ( .A(n19184), .B(n19185), .Z(n19181) );
  ANDN U22959 ( .B(n19186), .A(n5036), .Z(n19184) );
  XNOR U22960 ( .A(a[323]), .B(n19187), .Z(n5036) );
  IV U22961 ( .A(n19185), .Z(n19187) );
  XNOR U22962 ( .A(b[323]), .B(n19185), .Z(n19186) );
  XOR U22963 ( .A(n19188), .B(n19189), .Z(n19185) );
  ANDN U22964 ( .B(n19190), .A(n5087), .Z(n19188) );
  XNOR U22965 ( .A(a[322]), .B(n19191), .Z(n5087) );
  IV U22966 ( .A(n19189), .Z(n19191) );
  XNOR U22967 ( .A(b[322]), .B(n19189), .Z(n19190) );
  XOR U22968 ( .A(n19192), .B(n19193), .Z(n19189) );
  ANDN U22969 ( .B(n19194), .A(n5138), .Z(n19192) );
  XNOR U22970 ( .A(a[321]), .B(n19195), .Z(n5138) );
  IV U22971 ( .A(n19193), .Z(n19195) );
  XNOR U22972 ( .A(b[321]), .B(n19193), .Z(n19194) );
  XOR U22973 ( .A(n19196), .B(n19197), .Z(n19193) );
  ANDN U22974 ( .B(n19198), .A(n5189), .Z(n19196) );
  XNOR U22975 ( .A(a[320]), .B(n19199), .Z(n5189) );
  IV U22976 ( .A(n19197), .Z(n19199) );
  XNOR U22977 ( .A(b[320]), .B(n19197), .Z(n19198) );
  XOR U22978 ( .A(n19200), .B(n19201), .Z(n19197) );
  ANDN U22979 ( .B(n19202), .A(n5241), .Z(n19200) );
  XNOR U22980 ( .A(a[319]), .B(n19203), .Z(n5241) );
  IV U22981 ( .A(n19201), .Z(n19203) );
  XNOR U22982 ( .A(b[319]), .B(n19201), .Z(n19202) );
  XOR U22983 ( .A(n19204), .B(n19205), .Z(n19201) );
  ANDN U22984 ( .B(n19206), .A(n5292), .Z(n19204) );
  XNOR U22985 ( .A(a[318]), .B(n19207), .Z(n5292) );
  IV U22986 ( .A(n19205), .Z(n19207) );
  XNOR U22987 ( .A(b[318]), .B(n19205), .Z(n19206) );
  XOR U22988 ( .A(n19208), .B(n19209), .Z(n19205) );
  ANDN U22989 ( .B(n19210), .A(n5343), .Z(n19208) );
  XNOR U22990 ( .A(a[317]), .B(n19211), .Z(n5343) );
  IV U22991 ( .A(n19209), .Z(n19211) );
  XNOR U22992 ( .A(b[317]), .B(n19209), .Z(n19210) );
  XOR U22993 ( .A(n19212), .B(n19213), .Z(n19209) );
  ANDN U22994 ( .B(n19214), .A(n5394), .Z(n19212) );
  XNOR U22995 ( .A(a[316]), .B(n19215), .Z(n5394) );
  IV U22996 ( .A(n19213), .Z(n19215) );
  XNOR U22997 ( .A(b[316]), .B(n19213), .Z(n19214) );
  XOR U22998 ( .A(n19216), .B(n19217), .Z(n19213) );
  ANDN U22999 ( .B(n19218), .A(n5445), .Z(n19216) );
  XNOR U23000 ( .A(a[315]), .B(n19219), .Z(n5445) );
  IV U23001 ( .A(n19217), .Z(n19219) );
  XNOR U23002 ( .A(b[315]), .B(n19217), .Z(n19218) );
  XOR U23003 ( .A(n19220), .B(n19221), .Z(n19217) );
  ANDN U23004 ( .B(n19222), .A(n5496), .Z(n19220) );
  XNOR U23005 ( .A(a[314]), .B(n19223), .Z(n5496) );
  IV U23006 ( .A(n19221), .Z(n19223) );
  XNOR U23007 ( .A(b[314]), .B(n19221), .Z(n19222) );
  XOR U23008 ( .A(n19224), .B(n19225), .Z(n19221) );
  ANDN U23009 ( .B(n19226), .A(n5547), .Z(n19224) );
  XNOR U23010 ( .A(a[313]), .B(n19227), .Z(n5547) );
  IV U23011 ( .A(n19225), .Z(n19227) );
  XNOR U23012 ( .A(b[313]), .B(n19225), .Z(n19226) );
  XOR U23013 ( .A(n19228), .B(n19229), .Z(n19225) );
  ANDN U23014 ( .B(n19230), .A(n5598), .Z(n19228) );
  XNOR U23015 ( .A(a[312]), .B(n19231), .Z(n5598) );
  IV U23016 ( .A(n19229), .Z(n19231) );
  XNOR U23017 ( .A(b[312]), .B(n19229), .Z(n19230) );
  XOR U23018 ( .A(n19232), .B(n19233), .Z(n19229) );
  ANDN U23019 ( .B(n19234), .A(n5649), .Z(n19232) );
  XNOR U23020 ( .A(a[311]), .B(n19235), .Z(n5649) );
  IV U23021 ( .A(n19233), .Z(n19235) );
  XNOR U23022 ( .A(b[311]), .B(n19233), .Z(n19234) );
  XOR U23023 ( .A(n19236), .B(n19237), .Z(n19233) );
  ANDN U23024 ( .B(n19238), .A(n5700), .Z(n19236) );
  XNOR U23025 ( .A(a[310]), .B(n19239), .Z(n5700) );
  IV U23026 ( .A(n19237), .Z(n19239) );
  XNOR U23027 ( .A(b[310]), .B(n19237), .Z(n19238) );
  XOR U23028 ( .A(n19240), .B(n19241), .Z(n19237) );
  ANDN U23029 ( .B(n19242), .A(n5752), .Z(n19240) );
  XNOR U23030 ( .A(a[309]), .B(n19243), .Z(n5752) );
  IV U23031 ( .A(n19241), .Z(n19243) );
  XNOR U23032 ( .A(b[309]), .B(n19241), .Z(n19242) );
  XOR U23033 ( .A(n19244), .B(n19245), .Z(n19241) );
  ANDN U23034 ( .B(n19246), .A(n5803), .Z(n19244) );
  XNOR U23035 ( .A(a[308]), .B(n19247), .Z(n5803) );
  IV U23036 ( .A(n19245), .Z(n19247) );
  XNOR U23037 ( .A(b[308]), .B(n19245), .Z(n19246) );
  XOR U23038 ( .A(n19248), .B(n19249), .Z(n19245) );
  ANDN U23039 ( .B(n19250), .A(n5854), .Z(n19248) );
  XNOR U23040 ( .A(a[307]), .B(n19251), .Z(n5854) );
  IV U23041 ( .A(n19249), .Z(n19251) );
  XNOR U23042 ( .A(b[307]), .B(n19249), .Z(n19250) );
  XOR U23043 ( .A(n19252), .B(n19253), .Z(n19249) );
  ANDN U23044 ( .B(n19254), .A(n5905), .Z(n19252) );
  XNOR U23045 ( .A(a[306]), .B(n19255), .Z(n5905) );
  IV U23046 ( .A(n19253), .Z(n19255) );
  XNOR U23047 ( .A(b[306]), .B(n19253), .Z(n19254) );
  XOR U23048 ( .A(n19256), .B(n19257), .Z(n19253) );
  ANDN U23049 ( .B(n19258), .A(n5956), .Z(n19256) );
  XNOR U23050 ( .A(a[305]), .B(n19259), .Z(n5956) );
  IV U23051 ( .A(n19257), .Z(n19259) );
  XNOR U23052 ( .A(b[305]), .B(n19257), .Z(n19258) );
  XOR U23053 ( .A(n19260), .B(n19261), .Z(n19257) );
  ANDN U23054 ( .B(n19262), .A(n6007), .Z(n19260) );
  XNOR U23055 ( .A(a[304]), .B(n19263), .Z(n6007) );
  IV U23056 ( .A(n19261), .Z(n19263) );
  XNOR U23057 ( .A(b[304]), .B(n19261), .Z(n19262) );
  XOR U23058 ( .A(n19264), .B(n19265), .Z(n19261) );
  ANDN U23059 ( .B(n19266), .A(n6058), .Z(n19264) );
  XNOR U23060 ( .A(a[303]), .B(n19267), .Z(n6058) );
  IV U23061 ( .A(n19265), .Z(n19267) );
  XNOR U23062 ( .A(b[303]), .B(n19265), .Z(n19266) );
  XOR U23063 ( .A(n19268), .B(n19269), .Z(n19265) );
  ANDN U23064 ( .B(n19270), .A(n6109), .Z(n19268) );
  XNOR U23065 ( .A(a[302]), .B(n19271), .Z(n6109) );
  IV U23066 ( .A(n19269), .Z(n19271) );
  XNOR U23067 ( .A(b[302]), .B(n19269), .Z(n19270) );
  XOR U23068 ( .A(n19272), .B(n19273), .Z(n19269) );
  ANDN U23069 ( .B(n19274), .A(n6160), .Z(n19272) );
  XNOR U23070 ( .A(a[301]), .B(n19275), .Z(n6160) );
  IV U23071 ( .A(n19273), .Z(n19275) );
  XNOR U23072 ( .A(b[301]), .B(n19273), .Z(n19274) );
  XOR U23073 ( .A(n19276), .B(n19277), .Z(n19273) );
  ANDN U23074 ( .B(n19278), .A(n6211), .Z(n19276) );
  XNOR U23075 ( .A(a[300]), .B(n19279), .Z(n6211) );
  IV U23076 ( .A(n19277), .Z(n19279) );
  XNOR U23077 ( .A(b[300]), .B(n19277), .Z(n19278) );
  XOR U23078 ( .A(n19280), .B(n19281), .Z(n19277) );
  ANDN U23079 ( .B(n19282), .A(n6264), .Z(n19280) );
  XNOR U23080 ( .A(a[299]), .B(n19283), .Z(n6264) );
  IV U23081 ( .A(n19281), .Z(n19283) );
  XNOR U23082 ( .A(b[299]), .B(n19281), .Z(n19282) );
  XOR U23083 ( .A(n19284), .B(n19285), .Z(n19281) );
  ANDN U23084 ( .B(n19286), .A(n6315), .Z(n19284) );
  XNOR U23085 ( .A(a[298]), .B(n19287), .Z(n6315) );
  IV U23086 ( .A(n19285), .Z(n19287) );
  XNOR U23087 ( .A(b[298]), .B(n19285), .Z(n19286) );
  XOR U23088 ( .A(n19288), .B(n19289), .Z(n19285) );
  ANDN U23089 ( .B(n19290), .A(n6366), .Z(n19288) );
  XNOR U23090 ( .A(a[297]), .B(n19291), .Z(n6366) );
  IV U23091 ( .A(n19289), .Z(n19291) );
  XNOR U23092 ( .A(b[297]), .B(n19289), .Z(n19290) );
  XOR U23093 ( .A(n19292), .B(n19293), .Z(n19289) );
  ANDN U23094 ( .B(n19294), .A(n6417), .Z(n19292) );
  XNOR U23095 ( .A(a[296]), .B(n19295), .Z(n6417) );
  IV U23096 ( .A(n19293), .Z(n19295) );
  XNOR U23097 ( .A(b[296]), .B(n19293), .Z(n19294) );
  XOR U23098 ( .A(n19296), .B(n19297), .Z(n19293) );
  ANDN U23099 ( .B(n19298), .A(n6468), .Z(n19296) );
  XNOR U23100 ( .A(a[295]), .B(n19299), .Z(n6468) );
  IV U23101 ( .A(n19297), .Z(n19299) );
  XNOR U23102 ( .A(b[295]), .B(n19297), .Z(n19298) );
  XOR U23103 ( .A(n19300), .B(n19301), .Z(n19297) );
  ANDN U23104 ( .B(n19302), .A(n6519), .Z(n19300) );
  XNOR U23105 ( .A(a[294]), .B(n19303), .Z(n6519) );
  IV U23106 ( .A(n19301), .Z(n19303) );
  XNOR U23107 ( .A(b[294]), .B(n19301), .Z(n19302) );
  XOR U23108 ( .A(n19304), .B(n19305), .Z(n19301) );
  ANDN U23109 ( .B(n19306), .A(n6570), .Z(n19304) );
  XNOR U23110 ( .A(a[293]), .B(n19307), .Z(n6570) );
  IV U23111 ( .A(n19305), .Z(n19307) );
  XNOR U23112 ( .A(b[293]), .B(n19305), .Z(n19306) );
  XOR U23113 ( .A(n19308), .B(n19309), .Z(n19305) );
  ANDN U23114 ( .B(n19310), .A(n6621), .Z(n19308) );
  XNOR U23115 ( .A(a[292]), .B(n19311), .Z(n6621) );
  IV U23116 ( .A(n19309), .Z(n19311) );
  XNOR U23117 ( .A(b[292]), .B(n19309), .Z(n19310) );
  XOR U23118 ( .A(n19312), .B(n19313), .Z(n19309) );
  ANDN U23119 ( .B(n19314), .A(n6672), .Z(n19312) );
  XNOR U23120 ( .A(a[291]), .B(n19315), .Z(n6672) );
  IV U23121 ( .A(n19313), .Z(n19315) );
  XNOR U23122 ( .A(b[291]), .B(n19313), .Z(n19314) );
  XOR U23123 ( .A(n19316), .B(n19317), .Z(n19313) );
  ANDN U23124 ( .B(n19318), .A(n6723), .Z(n19316) );
  XNOR U23125 ( .A(a[290]), .B(n19319), .Z(n6723) );
  IV U23126 ( .A(n19317), .Z(n19319) );
  XNOR U23127 ( .A(b[290]), .B(n19317), .Z(n19318) );
  XOR U23128 ( .A(n19320), .B(n19321), .Z(n19317) );
  ANDN U23129 ( .B(n19322), .A(n6775), .Z(n19320) );
  XNOR U23130 ( .A(a[289]), .B(n19323), .Z(n6775) );
  IV U23131 ( .A(n19321), .Z(n19323) );
  XNOR U23132 ( .A(b[289]), .B(n19321), .Z(n19322) );
  XOR U23133 ( .A(n19324), .B(n19325), .Z(n19321) );
  ANDN U23134 ( .B(n19326), .A(n6826), .Z(n19324) );
  XNOR U23135 ( .A(a[288]), .B(n19327), .Z(n6826) );
  IV U23136 ( .A(n19325), .Z(n19327) );
  XNOR U23137 ( .A(b[288]), .B(n19325), .Z(n19326) );
  XOR U23138 ( .A(n19328), .B(n19329), .Z(n19325) );
  ANDN U23139 ( .B(n19330), .A(n6877), .Z(n19328) );
  XNOR U23140 ( .A(a[287]), .B(n19331), .Z(n6877) );
  IV U23141 ( .A(n19329), .Z(n19331) );
  XNOR U23142 ( .A(b[287]), .B(n19329), .Z(n19330) );
  XOR U23143 ( .A(n19332), .B(n19333), .Z(n19329) );
  ANDN U23144 ( .B(n19334), .A(n6928), .Z(n19332) );
  XNOR U23145 ( .A(a[286]), .B(n19335), .Z(n6928) );
  IV U23146 ( .A(n19333), .Z(n19335) );
  XNOR U23147 ( .A(b[286]), .B(n19333), .Z(n19334) );
  XOR U23148 ( .A(n19336), .B(n19337), .Z(n19333) );
  ANDN U23149 ( .B(n19338), .A(n6979), .Z(n19336) );
  XNOR U23150 ( .A(a[285]), .B(n19339), .Z(n6979) );
  IV U23151 ( .A(n19337), .Z(n19339) );
  XNOR U23152 ( .A(b[285]), .B(n19337), .Z(n19338) );
  XOR U23153 ( .A(n19340), .B(n19341), .Z(n19337) );
  ANDN U23154 ( .B(n19342), .A(n7030), .Z(n19340) );
  XNOR U23155 ( .A(a[284]), .B(n19343), .Z(n7030) );
  IV U23156 ( .A(n19341), .Z(n19343) );
  XNOR U23157 ( .A(b[284]), .B(n19341), .Z(n19342) );
  XOR U23158 ( .A(n19344), .B(n19345), .Z(n19341) );
  ANDN U23159 ( .B(n19346), .A(n7081), .Z(n19344) );
  XNOR U23160 ( .A(a[283]), .B(n19347), .Z(n7081) );
  IV U23161 ( .A(n19345), .Z(n19347) );
  XNOR U23162 ( .A(b[283]), .B(n19345), .Z(n19346) );
  XOR U23163 ( .A(n19348), .B(n19349), .Z(n19345) );
  ANDN U23164 ( .B(n19350), .A(n7132), .Z(n19348) );
  XNOR U23165 ( .A(a[282]), .B(n19351), .Z(n7132) );
  IV U23166 ( .A(n19349), .Z(n19351) );
  XNOR U23167 ( .A(b[282]), .B(n19349), .Z(n19350) );
  XOR U23168 ( .A(n19352), .B(n19353), .Z(n19349) );
  ANDN U23169 ( .B(n19354), .A(n7183), .Z(n19352) );
  XNOR U23170 ( .A(a[281]), .B(n19355), .Z(n7183) );
  IV U23171 ( .A(n19353), .Z(n19355) );
  XNOR U23172 ( .A(b[281]), .B(n19353), .Z(n19354) );
  XOR U23173 ( .A(n19356), .B(n19357), .Z(n19353) );
  ANDN U23174 ( .B(n19358), .A(n7234), .Z(n19356) );
  XNOR U23175 ( .A(a[280]), .B(n19359), .Z(n7234) );
  IV U23176 ( .A(n19357), .Z(n19359) );
  XNOR U23177 ( .A(b[280]), .B(n19357), .Z(n19358) );
  XOR U23178 ( .A(n19360), .B(n19361), .Z(n19357) );
  ANDN U23179 ( .B(n19362), .A(n7286), .Z(n19360) );
  XNOR U23180 ( .A(a[279]), .B(n19363), .Z(n7286) );
  IV U23181 ( .A(n19361), .Z(n19363) );
  XNOR U23182 ( .A(b[279]), .B(n19361), .Z(n19362) );
  XOR U23183 ( .A(n19364), .B(n19365), .Z(n19361) );
  ANDN U23184 ( .B(n19366), .A(n7337), .Z(n19364) );
  XNOR U23185 ( .A(a[278]), .B(n19367), .Z(n7337) );
  IV U23186 ( .A(n19365), .Z(n19367) );
  XNOR U23187 ( .A(b[278]), .B(n19365), .Z(n19366) );
  XOR U23188 ( .A(n19368), .B(n19369), .Z(n19365) );
  ANDN U23189 ( .B(n19370), .A(n7388), .Z(n19368) );
  XNOR U23190 ( .A(a[277]), .B(n19371), .Z(n7388) );
  IV U23191 ( .A(n19369), .Z(n19371) );
  XNOR U23192 ( .A(b[277]), .B(n19369), .Z(n19370) );
  XOR U23193 ( .A(n19372), .B(n19373), .Z(n19369) );
  ANDN U23194 ( .B(n19374), .A(n7439), .Z(n19372) );
  XNOR U23195 ( .A(a[276]), .B(n19375), .Z(n7439) );
  IV U23196 ( .A(n19373), .Z(n19375) );
  XNOR U23197 ( .A(b[276]), .B(n19373), .Z(n19374) );
  XOR U23198 ( .A(n19376), .B(n19377), .Z(n19373) );
  ANDN U23199 ( .B(n19378), .A(n7490), .Z(n19376) );
  XNOR U23200 ( .A(a[275]), .B(n19379), .Z(n7490) );
  IV U23201 ( .A(n19377), .Z(n19379) );
  XNOR U23202 ( .A(b[275]), .B(n19377), .Z(n19378) );
  XOR U23203 ( .A(n19380), .B(n19381), .Z(n19377) );
  ANDN U23204 ( .B(n19382), .A(n7541), .Z(n19380) );
  XNOR U23205 ( .A(a[274]), .B(n19383), .Z(n7541) );
  IV U23206 ( .A(n19381), .Z(n19383) );
  XNOR U23207 ( .A(b[274]), .B(n19381), .Z(n19382) );
  XOR U23208 ( .A(n19384), .B(n19385), .Z(n19381) );
  ANDN U23209 ( .B(n19386), .A(n7592), .Z(n19384) );
  XNOR U23210 ( .A(a[273]), .B(n19387), .Z(n7592) );
  IV U23211 ( .A(n19385), .Z(n19387) );
  XNOR U23212 ( .A(b[273]), .B(n19385), .Z(n19386) );
  XOR U23213 ( .A(n19388), .B(n19389), .Z(n19385) );
  ANDN U23214 ( .B(n19390), .A(n7643), .Z(n19388) );
  XNOR U23215 ( .A(a[272]), .B(n19391), .Z(n7643) );
  IV U23216 ( .A(n19389), .Z(n19391) );
  XNOR U23217 ( .A(b[272]), .B(n19389), .Z(n19390) );
  XOR U23218 ( .A(n19392), .B(n19393), .Z(n19389) );
  ANDN U23219 ( .B(n19394), .A(n7694), .Z(n19392) );
  XNOR U23220 ( .A(a[271]), .B(n19395), .Z(n7694) );
  IV U23221 ( .A(n19393), .Z(n19395) );
  XNOR U23222 ( .A(b[271]), .B(n19393), .Z(n19394) );
  XOR U23223 ( .A(n19396), .B(n19397), .Z(n19393) );
  ANDN U23224 ( .B(n19398), .A(n7745), .Z(n19396) );
  XNOR U23225 ( .A(a[270]), .B(n19399), .Z(n7745) );
  IV U23226 ( .A(n19397), .Z(n19399) );
  XNOR U23227 ( .A(b[270]), .B(n19397), .Z(n19398) );
  XOR U23228 ( .A(n19400), .B(n19401), .Z(n19397) );
  ANDN U23229 ( .B(n19402), .A(n7797), .Z(n19400) );
  XNOR U23230 ( .A(a[269]), .B(n19403), .Z(n7797) );
  IV U23231 ( .A(n19401), .Z(n19403) );
  XNOR U23232 ( .A(b[269]), .B(n19401), .Z(n19402) );
  XOR U23233 ( .A(n19404), .B(n19405), .Z(n19401) );
  ANDN U23234 ( .B(n19406), .A(n7848), .Z(n19404) );
  XNOR U23235 ( .A(a[268]), .B(n19407), .Z(n7848) );
  IV U23236 ( .A(n19405), .Z(n19407) );
  XNOR U23237 ( .A(b[268]), .B(n19405), .Z(n19406) );
  XOR U23238 ( .A(n19408), .B(n19409), .Z(n19405) );
  ANDN U23239 ( .B(n19410), .A(n7899), .Z(n19408) );
  XNOR U23240 ( .A(a[267]), .B(n19411), .Z(n7899) );
  IV U23241 ( .A(n19409), .Z(n19411) );
  XNOR U23242 ( .A(b[267]), .B(n19409), .Z(n19410) );
  XOR U23243 ( .A(n19412), .B(n19413), .Z(n19409) );
  ANDN U23244 ( .B(n19414), .A(n7950), .Z(n19412) );
  XNOR U23245 ( .A(a[266]), .B(n19415), .Z(n7950) );
  IV U23246 ( .A(n19413), .Z(n19415) );
  XNOR U23247 ( .A(b[266]), .B(n19413), .Z(n19414) );
  XOR U23248 ( .A(n19416), .B(n19417), .Z(n19413) );
  ANDN U23249 ( .B(n19418), .A(n8001), .Z(n19416) );
  XNOR U23250 ( .A(a[265]), .B(n19419), .Z(n8001) );
  IV U23251 ( .A(n19417), .Z(n19419) );
  XNOR U23252 ( .A(b[265]), .B(n19417), .Z(n19418) );
  XOR U23253 ( .A(n19420), .B(n19421), .Z(n19417) );
  ANDN U23254 ( .B(n19422), .A(n8052), .Z(n19420) );
  XNOR U23255 ( .A(a[264]), .B(n19423), .Z(n8052) );
  IV U23256 ( .A(n19421), .Z(n19423) );
  XNOR U23257 ( .A(b[264]), .B(n19421), .Z(n19422) );
  XOR U23258 ( .A(n19424), .B(n19425), .Z(n19421) );
  ANDN U23259 ( .B(n19426), .A(n8103), .Z(n19424) );
  XNOR U23260 ( .A(a[263]), .B(n19427), .Z(n8103) );
  IV U23261 ( .A(n19425), .Z(n19427) );
  XNOR U23262 ( .A(b[263]), .B(n19425), .Z(n19426) );
  XOR U23263 ( .A(n19428), .B(n19429), .Z(n19425) );
  ANDN U23264 ( .B(n19430), .A(n8154), .Z(n19428) );
  XNOR U23265 ( .A(a[262]), .B(n19431), .Z(n8154) );
  IV U23266 ( .A(n19429), .Z(n19431) );
  XNOR U23267 ( .A(b[262]), .B(n19429), .Z(n19430) );
  XOR U23268 ( .A(n19432), .B(n19433), .Z(n19429) );
  ANDN U23269 ( .B(n19434), .A(n8205), .Z(n19432) );
  XNOR U23270 ( .A(a[261]), .B(n19435), .Z(n8205) );
  IV U23271 ( .A(n19433), .Z(n19435) );
  XNOR U23272 ( .A(b[261]), .B(n19433), .Z(n19434) );
  XOR U23273 ( .A(n19436), .B(n19437), .Z(n19433) );
  ANDN U23274 ( .B(n19438), .A(n8256), .Z(n19436) );
  XNOR U23275 ( .A(a[260]), .B(n19439), .Z(n8256) );
  IV U23276 ( .A(n19437), .Z(n19439) );
  XNOR U23277 ( .A(b[260]), .B(n19437), .Z(n19438) );
  XOR U23278 ( .A(n19440), .B(n19441), .Z(n19437) );
  ANDN U23279 ( .B(n19442), .A(n8308), .Z(n19440) );
  XNOR U23280 ( .A(a[259]), .B(n19443), .Z(n8308) );
  IV U23281 ( .A(n19441), .Z(n19443) );
  XNOR U23282 ( .A(b[259]), .B(n19441), .Z(n19442) );
  XOR U23283 ( .A(n19444), .B(n19445), .Z(n19441) );
  ANDN U23284 ( .B(n19446), .A(n8359), .Z(n19444) );
  XNOR U23285 ( .A(a[258]), .B(n19447), .Z(n8359) );
  IV U23286 ( .A(n19445), .Z(n19447) );
  XNOR U23287 ( .A(b[258]), .B(n19445), .Z(n19446) );
  XOR U23288 ( .A(n19448), .B(n19449), .Z(n19445) );
  ANDN U23289 ( .B(n19450), .A(n8410), .Z(n19448) );
  XNOR U23290 ( .A(a[257]), .B(n19451), .Z(n8410) );
  IV U23291 ( .A(n19449), .Z(n19451) );
  XNOR U23292 ( .A(b[257]), .B(n19449), .Z(n19450) );
  XOR U23293 ( .A(n19452), .B(n19453), .Z(n19449) );
  ANDN U23294 ( .B(n19454), .A(n8461), .Z(n19452) );
  XNOR U23295 ( .A(a[256]), .B(n19455), .Z(n8461) );
  IV U23296 ( .A(n19453), .Z(n19455) );
  XNOR U23297 ( .A(b[256]), .B(n19453), .Z(n19454) );
  XOR U23298 ( .A(n19456), .B(n19457), .Z(n19453) );
  ANDN U23299 ( .B(n19458), .A(n8512), .Z(n19456) );
  XNOR U23300 ( .A(a[255]), .B(n19459), .Z(n8512) );
  IV U23301 ( .A(n19457), .Z(n19459) );
  XNOR U23302 ( .A(b[255]), .B(n19457), .Z(n19458) );
  XOR U23303 ( .A(n19460), .B(n19461), .Z(n19457) );
  ANDN U23304 ( .B(n19462), .A(n8563), .Z(n19460) );
  XNOR U23305 ( .A(a[254]), .B(n19463), .Z(n8563) );
  IV U23306 ( .A(n19461), .Z(n19463) );
  XNOR U23307 ( .A(b[254]), .B(n19461), .Z(n19462) );
  XOR U23308 ( .A(n19464), .B(n19465), .Z(n19461) );
  ANDN U23309 ( .B(n19466), .A(n8614), .Z(n19464) );
  XNOR U23310 ( .A(a[253]), .B(n19467), .Z(n8614) );
  IV U23311 ( .A(n19465), .Z(n19467) );
  XNOR U23312 ( .A(b[253]), .B(n19465), .Z(n19466) );
  XOR U23313 ( .A(n19468), .B(n19469), .Z(n19465) );
  ANDN U23314 ( .B(n19470), .A(n8665), .Z(n19468) );
  XNOR U23315 ( .A(a[252]), .B(n19471), .Z(n8665) );
  IV U23316 ( .A(n19469), .Z(n19471) );
  XNOR U23317 ( .A(b[252]), .B(n19469), .Z(n19470) );
  XOR U23318 ( .A(n19472), .B(n19473), .Z(n19469) );
  ANDN U23319 ( .B(n19474), .A(n8716), .Z(n19472) );
  XNOR U23320 ( .A(a[251]), .B(n19475), .Z(n8716) );
  IV U23321 ( .A(n19473), .Z(n19475) );
  XNOR U23322 ( .A(b[251]), .B(n19473), .Z(n19474) );
  XOR U23323 ( .A(n19476), .B(n19477), .Z(n19473) );
  ANDN U23324 ( .B(n19478), .A(n8767), .Z(n19476) );
  XNOR U23325 ( .A(a[250]), .B(n19479), .Z(n8767) );
  IV U23326 ( .A(n19477), .Z(n19479) );
  XNOR U23327 ( .A(b[250]), .B(n19477), .Z(n19478) );
  XOR U23328 ( .A(n19480), .B(n19481), .Z(n19477) );
  ANDN U23329 ( .B(n19482), .A(n8819), .Z(n19480) );
  XNOR U23330 ( .A(a[249]), .B(n19483), .Z(n8819) );
  IV U23331 ( .A(n19481), .Z(n19483) );
  XNOR U23332 ( .A(b[249]), .B(n19481), .Z(n19482) );
  XOR U23333 ( .A(n19484), .B(n19485), .Z(n19481) );
  ANDN U23334 ( .B(n19486), .A(n8870), .Z(n19484) );
  XNOR U23335 ( .A(a[248]), .B(n19487), .Z(n8870) );
  IV U23336 ( .A(n19485), .Z(n19487) );
  XNOR U23337 ( .A(b[248]), .B(n19485), .Z(n19486) );
  XOR U23338 ( .A(n19488), .B(n19489), .Z(n19485) );
  ANDN U23339 ( .B(n19490), .A(n8921), .Z(n19488) );
  XNOR U23340 ( .A(a[247]), .B(n19491), .Z(n8921) );
  IV U23341 ( .A(n19489), .Z(n19491) );
  XNOR U23342 ( .A(b[247]), .B(n19489), .Z(n19490) );
  XOR U23343 ( .A(n19492), .B(n19493), .Z(n19489) );
  ANDN U23344 ( .B(n19494), .A(n8972), .Z(n19492) );
  XNOR U23345 ( .A(a[246]), .B(n19495), .Z(n8972) );
  IV U23346 ( .A(n19493), .Z(n19495) );
  XNOR U23347 ( .A(b[246]), .B(n19493), .Z(n19494) );
  XOR U23348 ( .A(n19496), .B(n19497), .Z(n19493) );
  ANDN U23349 ( .B(n19498), .A(n9023), .Z(n19496) );
  XNOR U23350 ( .A(a[245]), .B(n19499), .Z(n9023) );
  IV U23351 ( .A(n19497), .Z(n19499) );
  XNOR U23352 ( .A(b[245]), .B(n19497), .Z(n19498) );
  XOR U23353 ( .A(n19500), .B(n19501), .Z(n19497) );
  ANDN U23354 ( .B(n19502), .A(n9074), .Z(n19500) );
  XNOR U23355 ( .A(a[244]), .B(n19503), .Z(n9074) );
  IV U23356 ( .A(n19501), .Z(n19503) );
  XNOR U23357 ( .A(b[244]), .B(n19501), .Z(n19502) );
  XOR U23358 ( .A(n19504), .B(n19505), .Z(n19501) );
  ANDN U23359 ( .B(n19506), .A(n9125), .Z(n19504) );
  XNOR U23360 ( .A(a[243]), .B(n19507), .Z(n9125) );
  IV U23361 ( .A(n19505), .Z(n19507) );
  XNOR U23362 ( .A(b[243]), .B(n19505), .Z(n19506) );
  XOR U23363 ( .A(n19508), .B(n19509), .Z(n19505) );
  ANDN U23364 ( .B(n19510), .A(n9176), .Z(n19508) );
  XNOR U23365 ( .A(a[242]), .B(n19511), .Z(n9176) );
  IV U23366 ( .A(n19509), .Z(n19511) );
  XNOR U23367 ( .A(b[242]), .B(n19509), .Z(n19510) );
  XOR U23368 ( .A(n19512), .B(n19513), .Z(n19509) );
  ANDN U23369 ( .B(n19514), .A(n9227), .Z(n19512) );
  XNOR U23370 ( .A(a[241]), .B(n19515), .Z(n9227) );
  IV U23371 ( .A(n19513), .Z(n19515) );
  XNOR U23372 ( .A(b[241]), .B(n19513), .Z(n19514) );
  XOR U23373 ( .A(n19516), .B(n19517), .Z(n19513) );
  ANDN U23374 ( .B(n19518), .A(n9278), .Z(n19516) );
  XNOR U23375 ( .A(a[240]), .B(n19519), .Z(n9278) );
  IV U23376 ( .A(n19517), .Z(n19519) );
  XNOR U23377 ( .A(b[240]), .B(n19517), .Z(n19518) );
  XOR U23378 ( .A(n19520), .B(n19521), .Z(n19517) );
  ANDN U23379 ( .B(n19522), .A(n9330), .Z(n19520) );
  XNOR U23380 ( .A(a[239]), .B(n19523), .Z(n9330) );
  IV U23381 ( .A(n19521), .Z(n19523) );
  XNOR U23382 ( .A(b[239]), .B(n19521), .Z(n19522) );
  XOR U23383 ( .A(n19524), .B(n19525), .Z(n19521) );
  ANDN U23384 ( .B(n19526), .A(n9381), .Z(n19524) );
  XNOR U23385 ( .A(a[238]), .B(n19527), .Z(n9381) );
  IV U23386 ( .A(n19525), .Z(n19527) );
  XNOR U23387 ( .A(b[238]), .B(n19525), .Z(n19526) );
  XOR U23388 ( .A(n19528), .B(n19529), .Z(n19525) );
  ANDN U23389 ( .B(n19530), .A(n9432), .Z(n19528) );
  XNOR U23390 ( .A(a[237]), .B(n19531), .Z(n9432) );
  IV U23391 ( .A(n19529), .Z(n19531) );
  XNOR U23392 ( .A(b[237]), .B(n19529), .Z(n19530) );
  XOR U23393 ( .A(n19532), .B(n19533), .Z(n19529) );
  ANDN U23394 ( .B(n19534), .A(n9483), .Z(n19532) );
  XNOR U23395 ( .A(a[236]), .B(n19535), .Z(n9483) );
  IV U23396 ( .A(n19533), .Z(n19535) );
  XNOR U23397 ( .A(b[236]), .B(n19533), .Z(n19534) );
  XOR U23398 ( .A(n19536), .B(n19537), .Z(n19533) );
  ANDN U23399 ( .B(n19538), .A(n9534), .Z(n19536) );
  XNOR U23400 ( .A(a[235]), .B(n19539), .Z(n9534) );
  IV U23401 ( .A(n19537), .Z(n19539) );
  XNOR U23402 ( .A(b[235]), .B(n19537), .Z(n19538) );
  XOR U23403 ( .A(n19540), .B(n19541), .Z(n19537) );
  ANDN U23404 ( .B(n19542), .A(n9585), .Z(n19540) );
  XNOR U23405 ( .A(a[234]), .B(n19543), .Z(n9585) );
  IV U23406 ( .A(n19541), .Z(n19543) );
  XNOR U23407 ( .A(b[234]), .B(n19541), .Z(n19542) );
  XOR U23408 ( .A(n19544), .B(n19545), .Z(n19541) );
  ANDN U23409 ( .B(n19546), .A(n9636), .Z(n19544) );
  XNOR U23410 ( .A(a[233]), .B(n19547), .Z(n9636) );
  IV U23411 ( .A(n19545), .Z(n19547) );
  XNOR U23412 ( .A(b[233]), .B(n19545), .Z(n19546) );
  XOR U23413 ( .A(n19548), .B(n19549), .Z(n19545) );
  ANDN U23414 ( .B(n19550), .A(n9687), .Z(n19548) );
  XNOR U23415 ( .A(a[232]), .B(n19551), .Z(n9687) );
  IV U23416 ( .A(n19549), .Z(n19551) );
  XNOR U23417 ( .A(b[232]), .B(n19549), .Z(n19550) );
  XOR U23418 ( .A(n19552), .B(n19553), .Z(n19549) );
  ANDN U23419 ( .B(n19554), .A(n9738), .Z(n19552) );
  XNOR U23420 ( .A(a[231]), .B(n19555), .Z(n9738) );
  IV U23421 ( .A(n19553), .Z(n19555) );
  XNOR U23422 ( .A(b[231]), .B(n19553), .Z(n19554) );
  XOR U23423 ( .A(n19556), .B(n19557), .Z(n19553) );
  ANDN U23424 ( .B(n19558), .A(n9789), .Z(n19556) );
  XNOR U23425 ( .A(a[230]), .B(n19559), .Z(n9789) );
  IV U23426 ( .A(n19557), .Z(n19559) );
  XNOR U23427 ( .A(b[230]), .B(n19557), .Z(n19558) );
  XOR U23428 ( .A(n19560), .B(n19561), .Z(n19557) );
  ANDN U23429 ( .B(n19562), .A(n9841), .Z(n19560) );
  XNOR U23430 ( .A(a[229]), .B(n19563), .Z(n9841) );
  IV U23431 ( .A(n19561), .Z(n19563) );
  XNOR U23432 ( .A(b[229]), .B(n19561), .Z(n19562) );
  XOR U23433 ( .A(n19564), .B(n19565), .Z(n19561) );
  ANDN U23434 ( .B(n19566), .A(n9892), .Z(n19564) );
  XNOR U23435 ( .A(a[228]), .B(n19567), .Z(n9892) );
  IV U23436 ( .A(n19565), .Z(n19567) );
  XNOR U23437 ( .A(b[228]), .B(n19565), .Z(n19566) );
  XOR U23438 ( .A(n19568), .B(n19569), .Z(n19565) );
  ANDN U23439 ( .B(n19570), .A(n9943), .Z(n19568) );
  XNOR U23440 ( .A(a[227]), .B(n19571), .Z(n9943) );
  IV U23441 ( .A(n19569), .Z(n19571) );
  XNOR U23442 ( .A(b[227]), .B(n19569), .Z(n19570) );
  XOR U23443 ( .A(n19572), .B(n19573), .Z(n19569) );
  ANDN U23444 ( .B(n19574), .A(n9994), .Z(n19572) );
  XNOR U23445 ( .A(a[226]), .B(n19575), .Z(n9994) );
  IV U23446 ( .A(n19573), .Z(n19575) );
  XNOR U23447 ( .A(b[226]), .B(n19573), .Z(n19574) );
  XOR U23448 ( .A(n19576), .B(n19577), .Z(n19573) );
  ANDN U23449 ( .B(n19578), .A(n10045), .Z(n19576) );
  XNOR U23450 ( .A(a[225]), .B(n19579), .Z(n10045) );
  IV U23451 ( .A(n19577), .Z(n19579) );
  XNOR U23452 ( .A(b[225]), .B(n19577), .Z(n19578) );
  XOR U23453 ( .A(n19580), .B(n19581), .Z(n19577) );
  ANDN U23454 ( .B(n19582), .A(n10096), .Z(n19580) );
  XNOR U23455 ( .A(a[224]), .B(n19583), .Z(n10096) );
  IV U23456 ( .A(n19581), .Z(n19583) );
  XNOR U23457 ( .A(b[224]), .B(n19581), .Z(n19582) );
  XOR U23458 ( .A(n19584), .B(n19585), .Z(n19581) );
  ANDN U23459 ( .B(n19586), .A(n10147), .Z(n19584) );
  XNOR U23460 ( .A(a[223]), .B(n19587), .Z(n10147) );
  IV U23461 ( .A(n19585), .Z(n19587) );
  XNOR U23462 ( .A(b[223]), .B(n19585), .Z(n19586) );
  XOR U23463 ( .A(n19588), .B(n19589), .Z(n19585) );
  ANDN U23464 ( .B(n19590), .A(n10198), .Z(n19588) );
  XNOR U23465 ( .A(a[222]), .B(n19591), .Z(n10198) );
  IV U23466 ( .A(n19589), .Z(n19591) );
  XNOR U23467 ( .A(b[222]), .B(n19589), .Z(n19590) );
  XOR U23468 ( .A(n19592), .B(n19593), .Z(n19589) );
  ANDN U23469 ( .B(n19594), .A(n10249), .Z(n19592) );
  XNOR U23470 ( .A(a[221]), .B(n19595), .Z(n10249) );
  IV U23471 ( .A(n19593), .Z(n19595) );
  XNOR U23472 ( .A(b[221]), .B(n19593), .Z(n19594) );
  XOR U23473 ( .A(n19596), .B(n19597), .Z(n19593) );
  ANDN U23474 ( .B(n19598), .A(n10300), .Z(n19596) );
  XNOR U23475 ( .A(a[220]), .B(n19599), .Z(n10300) );
  IV U23476 ( .A(n19597), .Z(n19599) );
  XNOR U23477 ( .A(b[220]), .B(n19597), .Z(n19598) );
  XOR U23478 ( .A(n19600), .B(n19601), .Z(n19597) );
  ANDN U23479 ( .B(n19602), .A(n10352), .Z(n19600) );
  XNOR U23480 ( .A(a[219]), .B(n19603), .Z(n10352) );
  IV U23481 ( .A(n19601), .Z(n19603) );
  XNOR U23482 ( .A(b[219]), .B(n19601), .Z(n19602) );
  XOR U23483 ( .A(n19604), .B(n19605), .Z(n19601) );
  ANDN U23484 ( .B(n19606), .A(n10403), .Z(n19604) );
  XNOR U23485 ( .A(a[218]), .B(n19607), .Z(n10403) );
  IV U23486 ( .A(n19605), .Z(n19607) );
  XNOR U23487 ( .A(b[218]), .B(n19605), .Z(n19606) );
  XOR U23488 ( .A(n19608), .B(n19609), .Z(n19605) );
  ANDN U23489 ( .B(n19610), .A(n10454), .Z(n19608) );
  XNOR U23490 ( .A(a[217]), .B(n19611), .Z(n10454) );
  IV U23491 ( .A(n19609), .Z(n19611) );
  XNOR U23492 ( .A(b[217]), .B(n19609), .Z(n19610) );
  XOR U23493 ( .A(n19612), .B(n19613), .Z(n19609) );
  ANDN U23494 ( .B(n19614), .A(n10505), .Z(n19612) );
  XNOR U23495 ( .A(a[216]), .B(n19615), .Z(n10505) );
  IV U23496 ( .A(n19613), .Z(n19615) );
  XNOR U23497 ( .A(b[216]), .B(n19613), .Z(n19614) );
  XOR U23498 ( .A(n19616), .B(n19617), .Z(n19613) );
  ANDN U23499 ( .B(n19618), .A(n10556), .Z(n19616) );
  XNOR U23500 ( .A(a[215]), .B(n19619), .Z(n10556) );
  IV U23501 ( .A(n19617), .Z(n19619) );
  XNOR U23502 ( .A(b[215]), .B(n19617), .Z(n19618) );
  XOR U23503 ( .A(n19620), .B(n19621), .Z(n19617) );
  ANDN U23504 ( .B(n19622), .A(n10607), .Z(n19620) );
  XNOR U23505 ( .A(a[214]), .B(n19623), .Z(n10607) );
  IV U23506 ( .A(n19621), .Z(n19623) );
  XNOR U23507 ( .A(b[214]), .B(n19621), .Z(n19622) );
  XOR U23508 ( .A(n19624), .B(n19625), .Z(n19621) );
  ANDN U23509 ( .B(n19626), .A(n10658), .Z(n19624) );
  XNOR U23510 ( .A(a[213]), .B(n19627), .Z(n10658) );
  IV U23511 ( .A(n19625), .Z(n19627) );
  XNOR U23512 ( .A(b[213]), .B(n19625), .Z(n19626) );
  XOR U23513 ( .A(n19628), .B(n19629), .Z(n19625) );
  ANDN U23514 ( .B(n19630), .A(n10709), .Z(n19628) );
  XNOR U23515 ( .A(a[212]), .B(n19631), .Z(n10709) );
  IV U23516 ( .A(n19629), .Z(n19631) );
  XNOR U23517 ( .A(b[212]), .B(n19629), .Z(n19630) );
  XOR U23518 ( .A(n19632), .B(n19633), .Z(n19629) );
  ANDN U23519 ( .B(n19634), .A(n10760), .Z(n19632) );
  XNOR U23520 ( .A(a[211]), .B(n19635), .Z(n10760) );
  IV U23521 ( .A(n19633), .Z(n19635) );
  XNOR U23522 ( .A(b[211]), .B(n19633), .Z(n19634) );
  XOR U23523 ( .A(n19636), .B(n19637), .Z(n19633) );
  ANDN U23524 ( .B(n19638), .A(n10811), .Z(n19636) );
  XNOR U23525 ( .A(a[210]), .B(n19639), .Z(n10811) );
  IV U23526 ( .A(n19637), .Z(n19639) );
  XNOR U23527 ( .A(b[210]), .B(n19637), .Z(n19638) );
  XOR U23528 ( .A(n19640), .B(n19641), .Z(n19637) );
  ANDN U23529 ( .B(n19642), .A(n10863), .Z(n19640) );
  XNOR U23530 ( .A(a[209]), .B(n19643), .Z(n10863) );
  IV U23531 ( .A(n19641), .Z(n19643) );
  XNOR U23532 ( .A(b[209]), .B(n19641), .Z(n19642) );
  XOR U23533 ( .A(n19644), .B(n19645), .Z(n19641) );
  ANDN U23534 ( .B(n19646), .A(n10914), .Z(n19644) );
  XNOR U23535 ( .A(a[208]), .B(n19647), .Z(n10914) );
  IV U23536 ( .A(n19645), .Z(n19647) );
  XNOR U23537 ( .A(b[208]), .B(n19645), .Z(n19646) );
  XOR U23538 ( .A(n19648), .B(n19649), .Z(n19645) );
  ANDN U23539 ( .B(n19650), .A(n10965), .Z(n19648) );
  XNOR U23540 ( .A(a[207]), .B(n19651), .Z(n10965) );
  IV U23541 ( .A(n19649), .Z(n19651) );
  XNOR U23542 ( .A(b[207]), .B(n19649), .Z(n19650) );
  XOR U23543 ( .A(n19652), .B(n19653), .Z(n19649) );
  ANDN U23544 ( .B(n19654), .A(n11016), .Z(n19652) );
  XNOR U23545 ( .A(a[206]), .B(n19655), .Z(n11016) );
  IV U23546 ( .A(n19653), .Z(n19655) );
  XNOR U23547 ( .A(b[206]), .B(n19653), .Z(n19654) );
  XOR U23548 ( .A(n19656), .B(n19657), .Z(n19653) );
  ANDN U23549 ( .B(n19658), .A(n11067), .Z(n19656) );
  XNOR U23550 ( .A(a[205]), .B(n19659), .Z(n11067) );
  IV U23551 ( .A(n19657), .Z(n19659) );
  XNOR U23552 ( .A(b[205]), .B(n19657), .Z(n19658) );
  XOR U23553 ( .A(n19660), .B(n19661), .Z(n19657) );
  ANDN U23554 ( .B(n19662), .A(n11118), .Z(n19660) );
  XNOR U23555 ( .A(a[204]), .B(n19663), .Z(n11118) );
  IV U23556 ( .A(n19661), .Z(n19663) );
  XNOR U23557 ( .A(b[204]), .B(n19661), .Z(n19662) );
  XOR U23558 ( .A(n19664), .B(n19665), .Z(n19661) );
  ANDN U23559 ( .B(n19666), .A(n11169), .Z(n19664) );
  XNOR U23560 ( .A(a[203]), .B(n19667), .Z(n11169) );
  IV U23561 ( .A(n19665), .Z(n19667) );
  XNOR U23562 ( .A(b[203]), .B(n19665), .Z(n19666) );
  XOR U23563 ( .A(n19668), .B(n19669), .Z(n19665) );
  ANDN U23564 ( .B(n19670), .A(n11220), .Z(n19668) );
  XNOR U23565 ( .A(a[202]), .B(n19671), .Z(n11220) );
  IV U23566 ( .A(n19669), .Z(n19671) );
  XNOR U23567 ( .A(b[202]), .B(n19669), .Z(n19670) );
  XOR U23568 ( .A(n19672), .B(n19673), .Z(n19669) );
  ANDN U23569 ( .B(n19674), .A(n11271), .Z(n19672) );
  XNOR U23570 ( .A(a[201]), .B(n19675), .Z(n11271) );
  IV U23571 ( .A(n19673), .Z(n19675) );
  XNOR U23572 ( .A(b[201]), .B(n19673), .Z(n19674) );
  XOR U23573 ( .A(n19676), .B(n19677), .Z(n19673) );
  ANDN U23574 ( .B(n19678), .A(n11322), .Z(n19676) );
  XNOR U23575 ( .A(a[200]), .B(n19679), .Z(n11322) );
  IV U23576 ( .A(n19677), .Z(n19679) );
  XNOR U23577 ( .A(b[200]), .B(n19677), .Z(n19678) );
  XOR U23578 ( .A(n19680), .B(n19681), .Z(n19677) );
  ANDN U23579 ( .B(n19682), .A(n11375), .Z(n19680) );
  XNOR U23580 ( .A(a[199]), .B(n19683), .Z(n11375) );
  IV U23581 ( .A(n19681), .Z(n19683) );
  XNOR U23582 ( .A(b[199]), .B(n19681), .Z(n19682) );
  XOR U23583 ( .A(n19684), .B(n19685), .Z(n19681) );
  ANDN U23584 ( .B(n19686), .A(n11426), .Z(n19684) );
  XNOR U23585 ( .A(a[198]), .B(n19687), .Z(n11426) );
  IV U23586 ( .A(n19685), .Z(n19687) );
  XNOR U23587 ( .A(b[198]), .B(n19685), .Z(n19686) );
  XOR U23588 ( .A(n19688), .B(n19689), .Z(n19685) );
  ANDN U23589 ( .B(n19690), .A(n11477), .Z(n19688) );
  XNOR U23590 ( .A(a[197]), .B(n19691), .Z(n11477) );
  IV U23591 ( .A(n19689), .Z(n19691) );
  XNOR U23592 ( .A(b[197]), .B(n19689), .Z(n19690) );
  XOR U23593 ( .A(n19692), .B(n19693), .Z(n19689) );
  ANDN U23594 ( .B(n19694), .A(n11528), .Z(n19692) );
  XNOR U23595 ( .A(a[196]), .B(n19695), .Z(n11528) );
  IV U23596 ( .A(n19693), .Z(n19695) );
  XNOR U23597 ( .A(b[196]), .B(n19693), .Z(n19694) );
  XOR U23598 ( .A(n19696), .B(n19697), .Z(n19693) );
  ANDN U23599 ( .B(n19698), .A(n11579), .Z(n19696) );
  XNOR U23600 ( .A(a[195]), .B(n19699), .Z(n11579) );
  IV U23601 ( .A(n19697), .Z(n19699) );
  XNOR U23602 ( .A(b[195]), .B(n19697), .Z(n19698) );
  XOR U23603 ( .A(n19700), .B(n19701), .Z(n19697) );
  ANDN U23604 ( .B(n19702), .A(n11630), .Z(n19700) );
  XNOR U23605 ( .A(a[194]), .B(n19703), .Z(n11630) );
  IV U23606 ( .A(n19701), .Z(n19703) );
  XNOR U23607 ( .A(b[194]), .B(n19701), .Z(n19702) );
  XOR U23608 ( .A(n19704), .B(n19705), .Z(n19701) );
  ANDN U23609 ( .B(n19706), .A(n11681), .Z(n19704) );
  XNOR U23610 ( .A(a[193]), .B(n19707), .Z(n11681) );
  IV U23611 ( .A(n19705), .Z(n19707) );
  XNOR U23612 ( .A(b[193]), .B(n19705), .Z(n19706) );
  XOR U23613 ( .A(n19708), .B(n19709), .Z(n19705) );
  ANDN U23614 ( .B(n19710), .A(n11732), .Z(n19708) );
  XNOR U23615 ( .A(a[192]), .B(n19711), .Z(n11732) );
  IV U23616 ( .A(n19709), .Z(n19711) );
  XNOR U23617 ( .A(b[192]), .B(n19709), .Z(n19710) );
  XOR U23618 ( .A(n19712), .B(n19713), .Z(n19709) );
  ANDN U23619 ( .B(n19714), .A(n11783), .Z(n19712) );
  XNOR U23620 ( .A(a[191]), .B(n19715), .Z(n11783) );
  IV U23621 ( .A(n19713), .Z(n19715) );
  XNOR U23622 ( .A(b[191]), .B(n19713), .Z(n19714) );
  XOR U23623 ( .A(n19716), .B(n19717), .Z(n19713) );
  ANDN U23624 ( .B(n19718), .A(n11834), .Z(n19716) );
  XNOR U23625 ( .A(a[190]), .B(n19719), .Z(n11834) );
  IV U23626 ( .A(n19717), .Z(n19719) );
  XNOR U23627 ( .A(b[190]), .B(n19717), .Z(n19718) );
  XOR U23628 ( .A(n19720), .B(n19721), .Z(n19717) );
  ANDN U23629 ( .B(n19722), .A(n11886), .Z(n19720) );
  XNOR U23630 ( .A(a[189]), .B(n19723), .Z(n11886) );
  IV U23631 ( .A(n19721), .Z(n19723) );
  XNOR U23632 ( .A(b[189]), .B(n19721), .Z(n19722) );
  XOR U23633 ( .A(n19724), .B(n19725), .Z(n19721) );
  ANDN U23634 ( .B(n19726), .A(n11937), .Z(n19724) );
  XNOR U23635 ( .A(a[188]), .B(n19727), .Z(n11937) );
  IV U23636 ( .A(n19725), .Z(n19727) );
  XNOR U23637 ( .A(b[188]), .B(n19725), .Z(n19726) );
  XOR U23638 ( .A(n19728), .B(n19729), .Z(n19725) );
  ANDN U23639 ( .B(n19730), .A(n11988), .Z(n19728) );
  XNOR U23640 ( .A(a[187]), .B(n19731), .Z(n11988) );
  IV U23641 ( .A(n19729), .Z(n19731) );
  XNOR U23642 ( .A(b[187]), .B(n19729), .Z(n19730) );
  XOR U23643 ( .A(n19732), .B(n19733), .Z(n19729) );
  ANDN U23644 ( .B(n19734), .A(n12039), .Z(n19732) );
  XNOR U23645 ( .A(a[186]), .B(n19735), .Z(n12039) );
  IV U23646 ( .A(n19733), .Z(n19735) );
  XNOR U23647 ( .A(b[186]), .B(n19733), .Z(n19734) );
  XOR U23648 ( .A(n19736), .B(n19737), .Z(n19733) );
  ANDN U23649 ( .B(n19738), .A(n12090), .Z(n19736) );
  XNOR U23650 ( .A(a[185]), .B(n19739), .Z(n12090) );
  IV U23651 ( .A(n19737), .Z(n19739) );
  XNOR U23652 ( .A(b[185]), .B(n19737), .Z(n19738) );
  XOR U23653 ( .A(n19740), .B(n19741), .Z(n19737) );
  ANDN U23654 ( .B(n19742), .A(n12141), .Z(n19740) );
  XNOR U23655 ( .A(a[184]), .B(n19743), .Z(n12141) );
  IV U23656 ( .A(n19741), .Z(n19743) );
  XNOR U23657 ( .A(b[184]), .B(n19741), .Z(n19742) );
  XOR U23658 ( .A(n19744), .B(n19745), .Z(n19741) );
  ANDN U23659 ( .B(n19746), .A(n12192), .Z(n19744) );
  XNOR U23660 ( .A(a[183]), .B(n19747), .Z(n12192) );
  IV U23661 ( .A(n19745), .Z(n19747) );
  XNOR U23662 ( .A(b[183]), .B(n19745), .Z(n19746) );
  XOR U23663 ( .A(n19748), .B(n19749), .Z(n19745) );
  ANDN U23664 ( .B(n19750), .A(n12243), .Z(n19748) );
  XNOR U23665 ( .A(a[182]), .B(n19751), .Z(n12243) );
  IV U23666 ( .A(n19749), .Z(n19751) );
  XNOR U23667 ( .A(b[182]), .B(n19749), .Z(n19750) );
  XOR U23668 ( .A(n19752), .B(n19753), .Z(n19749) );
  ANDN U23669 ( .B(n19754), .A(n12294), .Z(n19752) );
  XNOR U23670 ( .A(a[181]), .B(n19755), .Z(n12294) );
  IV U23671 ( .A(n19753), .Z(n19755) );
  XNOR U23672 ( .A(b[181]), .B(n19753), .Z(n19754) );
  XOR U23673 ( .A(n19756), .B(n19757), .Z(n19753) );
  ANDN U23674 ( .B(n19758), .A(n12345), .Z(n19756) );
  XNOR U23675 ( .A(a[180]), .B(n19759), .Z(n12345) );
  IV U23676 ( .A(n19757), .Z(n19759) );
  XNOR U23677 ( .A(b[180]), .B(n19757), .Z(n19758) );
  XOR U23678 ( .A(n19760), .B(n19761), .Z(n19757) );
  ANDN U23679 ( .B(n19762), .A(n12397), .Z(n19760) );
  XNOR U23680 ( .A(a[179]), .B(n19763), .Z(n12397) );
  IV U23681 ( .A(n19761), .Z(n19763) );
  XNOR U23682 ( .A(b[179]), .B(n19761), .Z(n19762) );
  XOR U23683 ( .A(n19764), .B(n19765), .Z(n19761) );
  ANDN U23684 ( .B(n19766), .A(n12448), .Z(n19764) );
  XNOR U23685 ( .A(a[178]), .B(n19767), .Z(n12448) );
  IV U23686 ( .A(n19765), .Z(n19767) );
  XNOR U23687 ( .A(b[178]), .B(n19765), .Z(n19766) );
  XOR U23688 ( .A(n19768), .B(n19769), .Z(n19765) );
  ANDN U23689 ( .B(n19770), .A(n12499), .Z(n19768) );
  XNOR U23690 ( .A(a[177]), .B(n19771), .Z(n12499) );
  IV U23691 ( .A(n19769), .Z(n19771) );
  XNOR U23692 ( .A(b[177]), .B(n19769), .Z(n19770) );
  XOR U23693 ( .A(n19772), .B(n19773), .Z(n19769) );
  ANDN U23694 ( .B(n19774), .A(n12550), .Z(n19772) );
  XNOR U23695 ( .A(a[176]), .B(n19775), .Z(n12550) );
  IV U23696 ( .A(n19773), .Z(n19775) );
  XNOR U23697 ( .A(b[176]), .B(n19773), .Z(n19774) );
  XOR U23698 ( .A(n19776), .B(n19777), .Z(n19773) );
  ANDN U23699 ( .B(n19778), .A(n12601), .Z(n19776) );
  XNOR U23700 ( .A(a[175]), .B(n19779), .Z(n12601) );
  IV U23701 ( .A(n19777), .Z(n19779) );
  XNOR U23702 ( .A(b[175]), .B(n19777), .Z(n19778) );
  XOR U23703 ( .A(n19780), .B(n19781), .Z(n19777) );
  ANDN U23704 ( .B(n19782), .A(n12652), .Z(n19780) );
  XNOR U23705 ( .A(a[174]), .B(n19783), .Z(n12652) );
  IV U23706 ( .A(n19781), .Z(n19783) );
  XNOR U23707 ( .A(b[174]), .B(n19781), .Z(n19782) );
  XOR U23708 ( .A(n19784), .B(n19785), .Z(n19781) );
  ANDN U23709 ( .B(n19786), .A(n12703), .Z(n19784) );
  XNOR U23710 ( .A(a[173]), .B(n19787), .Z(n12703) );
  IV U23711 ( .A(n19785), .Z(n19787) );
  XNOR U23712 ( .A(b[173]), .B(n19785), .Z(n19786) );
  XOR U23713 ( .A(n19788), .B(n19789), .Z(n19785) );
  ANDN U23714 ( .B(n19790), .A(n12754), .Z(n19788) );
  XNOR U23715 ( .A(a[172]), .B(n19791), .Z(n12754) );
  IV U23716 ( .A(n19789), .Z(n19791) );
  XNOR U23717 ( .A(b[172]), .B(n19789), .Z(n19790) );
  XOR U23718 ( .A(n19792), .B(n19793), .Z(n19789) );
  ANDN U23719 ( .B(n19794), .A(n12805), .Z(n19792) );
  XNOR U23720 ( .A(a[171]), .B(n19795), .Z(n12805) );
  IV U23721 ( .A(n19793), .Z(n19795) );
  XNOR U23722 ( .A(b[171]), .B(n19793), .Z(n19794) );
  XOR U23723 ( .A(n19796), .B(n19797), .Z(n19793) );
  ANDN U23724 ( .B(n19798), .A(n12856), .Z(n19796) );
  XNOR U23725 ( .A(a[170]), .B(n19799), .Z(n12856) );
  IV U23726 ( .A(n19797), .Z(n19799) );
  XNOR U23727 ( .A(b[170]), .B(n19797), .Z(n19798) );
  XOR U23728 ( .A(n19800), .B(n19801), .Z(n19797) );
  ANDN U23729 ( .B(n19802), .A(n12908), .Z(n19800) );
  XNOR U23730 ( .A(a[169]), .B(n19803), .Z(n12908) );
  IV U23731 ( .A(n19801), .Z(n19803) );
  XNOR U23732 ( .A(b[169]), .B(n19801), .Z(n19802) );
  XOR U23733 ( .A(n19804), .B(n19805), .Z(n19801) );
  ANDN U23734 ( .B(n19806), .A(n12959), .Z(n19804) );
  XNOR U23735 ( .A(a[168]), .B(n19807), .Z(n12959) );
  IV U23736 ( .A(n19805), .Z(n19807) );
  XNOR U23737 ( .A(b[168]), .B(n19805), .Z(n19806) );
  XOR U23738 ( .A(n19808), .B(n19809), .Z(n19805) );
  ANDN U23739 ( .B(n19810), .A(n13010), .Z(n19808) );
  XNOR U23740 ( .A(a[167]), .B(n19811), .Z(n13010) );
  IV U23741 ( .A(n19809), .Z(n19811) );
  XNOR U23742 ( .A(b[167]), .B(n19809), .Z(n19810) );
  XOR U23743 ( .A(n19812), .B(n19813), .Z(n19809) );
  ANDN U23744 ( .B(n19814), .A(n13061), .Z(n19812) );
  XNOR U23745 ( .A(a[166]), .B(n19815), .Z(n13061) );
  IV U23746 ( .A(n19813), .Z(n19815) );
  XNOR U23747 ( .A(b[166]), .B(n19813), .Z(n19814) );
  XOR U23748 ( .A(n19816), .B(n19817), .Z(n19813) );
  ANDN U23749 ( .B(n19818), .A(n13112), .Z(n19816) );
  XNOR U23750 ( .A(a[165]), .B(n19819), .Z(n13112) );
  IV U23751 ( .A(n19817), .Z(n19819) );
  XNOR U23752 ( .A(b[165]), .B(n19817), .Z(n19818) );
  XOR U23753 ( .A(n19820), .B(n19821), .Z(n19817) );
  ANDN U23754 ( .B(n19822), .A(n13163), .Z(n19820) );
  XNOR U23755 ( .A(a[164]), .B(n19823), .Z(n13163) );
  IV U23756 ( .A(n19821), .Z(n19823) );
  XNOR U23757 ( .A(b[164]), .B(n19821), .Z(n19822) );
  XOR U23758 ( .A(n19824), .B(n19825), .Z(n19821) );
  ANDN U23759 ( .B(n19826), .A(n13214), .Z(n19824) );
  XNOR U23760 ( .A(a[163]), .B(n19827), .Z(n13214) );
  IV U23761 ( .A(n19825), .Z(n19827) );
  XNOR U23762 ( .A(b[163]), .B(n19825), .Z(n19826) );
  XOR U23763 ( .A(n19828), .B(n19829), .Z(n19825) );
  ANDN U23764 ( .B(n19830), .A(n13265), .Z(n19828) );
  XNOR U23765 ( .A(a[162]), .B(n19831), .Z(n13265) );
  IV U23766 ( .A(n19829), .Z(n19831) );
  XNOR U23767 ( .A(b[162]), .B(n19829), .Z(n19830) );
  XOR U23768 ( .A(n19832), .B(n19833), .Z(n19829) );
  ANDN U23769 ( .B(n19834), .A(n13316), .Z(n19832) );
  XNOR U23770 ( .A(a[161]), .B(n19835), .Z(n13316) );
  IV U23771 ( .A(n19833), .Z(n19835) );
  XNOR U23772 ( .A(b[161]), .B(n19833), .Z(n19834) );
  XOR U23773 ( .A(n19836), .B(n19837), .Z(n19833) );
  ANDN U23774 ( .B(n19838), .A(n13367), .Z(n19836) );
  XNOR U23775 ( .A(a[160]), .B(n19839), .Z(n13367) );
  IV U23776 ( .A(n19837), .Z(n19839) );
  XNOR U23777 ( .A(b[160]), .B(n19837), .Z(n19838) );
  XOR U23778 ( .A(n19840), .B(n19841), .Z(n19837) );
  ANDN U23779 ( .B(n19842), .A(n13419), .Z(n19840) );
  XNOR U23780 ( .A(a[159]), .B(n19843), .Z(n13419) );
  IV U23781 ( .A(n19841), .Z(n19843) );
  XNOR U23782 ( .A(b[159]), .B(n19841), .Z(n19842) );
  XOR U23783 ( .A(n19844), .B(n19845), .Z(n19841) );
  ANDN U23784 ( .B(n19846), .A(n13470), .Z(n19844) );
  XNOR U23785 ( .A(a[158]), .B(n19847), .Z(n13470) );
  IV U23786 ( .A(n19845), .Z(n19847) );
  XNOR U23787 ( .A(b[158]), .B(n19845), .Z(n19846) );
  XOR U23788 ( .A(n19848), .B(n19849), .Z(n19845) );
  ANDN U23789 ( .B(n19850), .A(n13521), .Z(n19848) );
  XNOR U23790 ( .A(a[157]), .B(n19851), .Z(n13521) );
  IV U23791 ( .A(n19849), .Z(n19851) );
  XNOR U23792 ( .A(b[157]), .B(n19849), .Z(n19850) );
  XOR U23793 ( .A(n19852), .B(n19853), .Z(n19849) );
  ANDN U23794 ( .B(n19854), .A(n13572), .Z(n19852) );
  XNOR U23795 ( .A(a[156]), .B(n19855), .Z(n13572) );
  IV U23796 ( .A(n19853), .Z(n19855) );
  XNOR U23797 ( .A(b[156]), .B(n19853), .Z(n19854) );
  XOR U23798 ( .A(n19856), .B(n19857), .Z(n19853) );
  ANDN U23799 ( .B(n19858), .A(n13623), .Z(n19856) );
  XNOR U23800 ( .A(a[155]), .B(n19859), .Z(n13623) );
  IV U23801 ( .A(n19857), .Z(n19859) );
  XNOR U23802 ( .A(b[155]), .B(n19857), .Z(n19858) );
  XOR U23803 ( .A(n19860), .B(n19861), .Z(n19857) );
  ANDN U23804 ( .B(n19862), .A(n13674), .Z(n19860) );
  XNOR U23805 ( .A(a[154]), .B(n19863), .Z(n13674) );
  IV U23806 ( .A(n19861), .Z(n19863) );
  XNOR U23807 ( .A(b[154]), .B(n19861), .Z(n19862) );
  XOR U23808 ( .A(n19864), .B(n19865), .Z(n19861) );
  ANDN U23809 ( .B(n19866), .A(n13725), .Z(n19864) );
  XNOR U23810 ( .A(a[153]), .B(n19867), .Z(n13725) );
  IV U23811 ( .A(n19865), .Z(n19867) );
  XNOR U23812 ( .A(b[153]), .B(n19865), .Z(n19866) );
  XOR U23813 ( .A(n19868), .B(n19869), .Z(n19865) );
  ANDN U23814 ( .B(n19870), .A(n13776), .Z(n19868) );
  XNOR U23815 ( .A(a[152]), .B(n19871), .Z(n13776) );
  IV U23816 ( .A(n19869), .Z(n19871) );
  XNOR U23817 ( .A(b[152]), .B(n19869), .Z(n19870) );
  XOR U23818 ( .A(n19872), .B(n19873), .Z(n19869) );
  ANDN U23819 ( .B(n19874), .A(n13827), .Z(n19872) );
  XNOR U23820 ( .A(a[151]), .B(n19875), .Z(n13827) );
  IV U23821 ( .A(n19873), .Z(n19875) );
  XNOR U23822 ( .A(b[151]), .B(n19873), .Z(n19874) );
  XOR U23823 ( .A(n19876), .B(n19877), .Z(n19873) );
  ANDN U23824 ( .B(n19878), .A(n13878), .Z(n19876) );
  XNOR U23825 ( .A(a[150]), .B(n19879), .Z(n13878) );
  IV U23826 ( .A(n19877), .Z(n19879) );
  XNOR U23827 ( .A(b[150]), .B(n19877), .Z(n19878) );
  XOR U23828 ( .A(n19880), .B(n19881), .Z(n19877) );
  ANDN U23829 ( .B(n19882), .A(n13930), .Z(n19880) );
  XNOR U23830 ( .A(a[149]), .B(n19883), .Z(n13930) );
  IV U23831 ( .A(n19881), .Z(n19883) );
  XNOR U23832 ( .A(b[149]), .B(n19881), .Z(n19882) );
  XOR U23833 ( .A(n19884), .B(n19885), .Z(n19881) );
  ANDN U23834 ( .B(n19886), .A(n13981), .Z(n19884) );
  XNOR U23835 ( .A(a[148]), .B(n19887), .Z(n13981) );
  IV U23836 ( .A(n19885), .Z(n19887) );
  XNOR U23837 ( .A(b[148]), .B(n19885), .Z(n19886) );
  XOR U23838 ( .A(n19888), .B(n19889), .Z(n19885) );
  ANDN U23839 ( .B(n19890), .A(n14032), .Z(n19888) );
  XNOR U23840 ( .A(a[147]), .B(n19891), .Z(n14032) );
  IV U23841 ( .A(n19889), .Z(n19891) );
  XNOR U23842 ( .A(b[147]), .B(n19889), .Z(n19890) );
  XOR U23843 ( .A(n19892), .B(n19893), .Z(n19889) );
  ANDN U23844 ( .B(n19894), .A(n14083), .Z(n19892) );
  XNOR U23845 ( .A(a[146]), .B(n19895), .Z(n14083) );
  IV U23846 ( .A(n19893), .Z(n19895) );
  XNOR U23847 ( .A(b[146]), .B(n19893), .Z(n19894) );
  XOR U23848 ( .A(n19896), .B(n19897), .Z(n19893) );
  ANDN U23849 ( .B(n19898), .A(n14134), .Z(n19896) );
  XNOR U23850 ( .A(a[145]), .B(n19899), .Z(n14134) );
  IV U23851 ( .A(n19897), .Z(n19899) );
  XNOR U23852 ( .A(b[145]), .B(n19897), .Z(n19898) );
  XOR U23853 ( .A(n19900), .B(n19901), .Z(n19897) );
  ANDN U23854 ( .B(n19902), .A(n14185), .Z(n19900) );
  XNOR U23855 ( .A(a[144]), .B(n19903), .Z(n14185) );
  IV U23856 ( .A(n19901), .Z(n19903) );
  XNOR U23857 ( .A(b[144]), .B(n19901), .Z(n19902) );
  XOR U23858 ( .A(n19904), .B(n19905), .Z(n19901) );
  ANDN U23859 ( .B(n19906), .A(n14236), .Z(n19904) );
  XNOR U23860 ( .A(a[143]), .B(n19907), .Z(n14236) );
  IV U23861 ( .A(n19905), .Z(n19907) );
  XNOR U23862 ( .A(b[143]), .B(n19905), .Z(n19906) );
  XOR U23863 ( .A(n19908), .B(n19909), .Z(n19905) );
  ANDN U23864 ( .B(n19910), .A(n14287), .Z(n19908) );
  XNOR U23865 ( .A(a[142]), .B(n19911), .Z(n14287) );
  IV U23866 ( .A(n19909), .Z(n19911) );
  XNOR U23867 ( .A(b[142]), .B(n19909), .Z(n19910) );
  XOR U23868 ( .A(n19912), .B(n19913), .Z(n19909) );
  ANDN U23869 ( .B(n19914), .A(n14338), .Z(n19912) );
  XNOR U23870 ( .A(a[141]), .B(n19915), .Z(n14338) );
  IV U23871 ( .A(n19913), .Z(n19915) );
  XNOR U23872 ( .A(b[141]), .B(n19913), .Z(n19914) );
  XOR U23873 ( .A(n19916), .B(n19917), .Z(n19913) );
  ANDN U23874 ( .B(n19918), .A(n14389), .Z(n19916) );
  XNOR U23875 ( .A(a[140]), .B(n19919), .Z(n14389) );
  IV U23876 ( .A(n19917), .Z(n19919) );
  XNOR U23877 ( .A(b[140]), .B(n19917), .Z(n19918) );
  XOR U23878 ( .A(n19920), .B(n19921), .Z(n19917) );
  ANDN U23879 ( .B(n19922), .A(n14441), .Z(n19920) );
  XNOR U23880 ( .A(a[139]), .B(n19923), .Z(n14441) );
  IV U23881 ( .A(n19921), .Z(n19923) );
  XNOR U23882 ( .A(b[139]), .B(n19921), .Z(n19922) );
  XOR U23883 ( .A(n19924), .B(n19925), .Z(n19921) );
  ANDN U23884 ( .B(n19926), .A(n14492), .Z(n19924) );
  XNOR U23885 ( .A(a[138]), .B(n19927), .Z(n14492) );
  IV U23886 ( .A(n19925), .Z(n19927) );
  XNOR U23887 ( .A(b[138]), .B(n19925), .Z(n19926) );
  XOR U23888 ( .A(n19928), .B(n19929), .Z(n19925) );
  ANDN U23889 ( .B(n19930), .A(n14543), .Z(n19928) );
  XNOR U23890 ( .A(a[137]), .B(n19931), .Z(n14543) );
  IV U23891 ( .A(n19929), .Z(n19931) );
  XNOR U23892 ( .A(b[137]), .B(n19929), .Z(n19930) );
  XOR U23893 ( .A(n19932), .B(n19933), .Z(n19929) );
  ANDN U23894 ( .B(n19934), .A(n14594), .Z(n19932) );
  XNOR U23895 ( .A(a[136]), .B(n19935), .Z(n14594) );
  IV U23896 ( .A(n19933), .Z(n19935) );
  XNOR U23897 ( .A(b[136]), .B(n19933), .Z(n19934) );
  XOR U23898 ( .A(n19936), .B(n19937), .Z(n19933) );
  ANDN U23899 ( .B(n19938), .A(n14645), .Z(n19936) );
  XNOR U23900 ( .A(a[135]), .B(n19939), .Z(n14645) );
  IV U23901 ( .A(n19937), .Z(n19939) );
  XNOR U23902 ( .A(b[135]), .B(n19937), .Z(n19938) );
  XOR U23903 ( .A(n19940), .B(n19941), .Z(n19937) );
  ANDN U23904 ( .B(n19942), .A(n14696), .Z(n19940) );
  XNOR U23905 ( .A(a[134]), .B(n19943), .Z(n14696) );
  IV U23906 ( .A(n19941), .Z(n19943) );
  XNOR U23907 ( .A(b[134]), .B(n19941), .Z(n19942) );
  XOR U23908 ( .A(n19944), .B(n19945), .Z(n19941) );
  ANDN U23909 ( .B(n19946), .A(n14747), .Z(n19944) );
  XNOR U23910 ( .A(a[133]), .B(n19947), .Z(n14747) );
  IV U23911 ( .A(n19945), .Z(n19947) );
  XNOR U23912 ( .A(b[133]), .B(n19945), .Z(n19946) );
  XOR U23913 ( .A(n19948), .B(n19949), .Z(n19945) );
  ANDN U23914 ( .B(n19950), .A(n14798), .Z(n19948) );
  XNOR U23915 ( .A(a[132]), .B(n19951), .Z(n14798) );
  IV U23916 ( .A(n19949), .Z(n19951) );
  XNOR U23917 ( .A(b[132]), .B(n19949), .Z(n19950) );
  XOR U23918 ( .A(n19952), .B(n19953), .Z(n19949) );
  ANDN U23919 ( .B(n19954), .A(n14849), .Z(n19952) );
  XNOR U23920 ( .A(a[131]), .B(n19955), .Z(n14849) );
  IV U23921 ( .A(n19953), .Z(n19955) );
  XNOR U23922 ( .A(b[131]), .B(n19953), .Z(n19954) );
  XOR U23923 ( .A(n19956), .B(n19957), .Z(n19953) );
  ANDN U23924 ( .B(n19958), .A(n14900), .Z(n19956) );
  XNOR U23925 ( .A(a[130]), .B(n19959), .Z(n14900) );
  IV U23926 ( .A(n19957), .Z(n19959) );
  XNOR U23927 ( .A(b[130]), .B(n19957), .Z(n19958) );
  XOR U23928 ( .A(n19960), .B(n19961), .Z(n19957) );
  ANDN U23929 ( .B(n19962), .A(n14952), .Z(n19960) );
  XNOR U23930 ( .A(a[129]), .B(n19963), .Z(n14952) );
  IV U23931 ( .A(n19961), .Z(n19963) );
  XNOR U23932 ( .A(b[129]), .B(n19961), .Z(n19962) );
  XOR U23933 ( .A(n19964), .B(n19965), .Z(n19961) );
  ANDN U23934 ( .B(n19966), .A(n15003), .Z(n19964) );
  XNOR U23935 ( .A(a[128]), .B(n19967), .Z(n15003) );
  IV U23936 ( .A(n19965), .Z(n19967) );
  XNOR U23937 ( .A(b[128]), .B(n19965), .Z(n19966) );
  XOR U23938 ( .A(n19968), .B(n19969), .Z(n19965) );
  ANDN U23939 ( .B(n19970), .A(n15054), .Z(n19968) );
  XNOR U23940 ( .A(a[127]), .B(n19971), .Z(n15054) );
  IV U23941 ( .A(n19969), .Z(n19971) );
  XNOR U23942 ( .A(b[127]), .B(n19969), .Z(n19970) );
  XOR U23943 ( .A(n19972), .B(n19973), .Z(n19969) );
  ANDN U23944 ( .B(n19974), .A(n15105), .Z(n19972) );
  XNOR U23945 ( .A(a[126]), .B(n19975), .Z(n15105) );
  IV U23946 ( .A(n19973), .Z(n19975) );
  XNOR U23947 ( .A(b[126]), .B(n19973), .Z(n19974) );
  XOR U23948 ( .A(n19976), .B(n19977), .Z(n19973) );
  ANDN U23949 ( .B(n19978), .A(n15156), .Z(n19976) );
  XNOR U23950 ( .A(a[125]), .B(n19979), .Z(n15156) );
  IV U23951 ( .A(n19977), .Z(n19979) );
  XNOR U23952 ( .A(b[125]), .B(n19977), .Z(n19978) );
  XOR U23953 ( .A(n19980), .B(n19981), .Z(n19977) );
  ANDN U23954 ( .B(n19982), .A(n15207), .Z(n19980) );
  XNOR U23955 ( .A(a[124]), .B(n19983), .Z(n15207) );
  IV U23956 ( .A(n19981), .Z(n19983) );
  XNOR U23957 ( .A(b[124]), .B(n19981), .Z(n19982) );
  XOR U23958 ( .A(n19984), .B(n19985), .Z(n19981) );
  ANDN U23959 ( .B(n19986), .A(n15258), .Z(n19984) );
  XNOR U23960 ( .A(a[123]), .B(n19987), .Z(n15258) );
  IV U23961 ( .A(n19985), .Z(n19987) );
  XNOR U23962 ( .A(b[123]), .B(n19985), .Z(n19986) );
  XOR U23963 ( .A(n19988), .B(n19989), .Z(n19985) );
  ANDN U23964 ( .B(n19990), .A(n15309), .Z(n19988) );
  XNOR U23965 ( .A(a[122]), .B(n19991), .Z(n15309) );
  IV U23966 ( .A(n19989), .Z(n19991) );
  XNOR U23967 ( .A(b[122]), .B(n19989), .Z(n19990) );
  XOR U23968 ( .A(n19992), .B(n19993), .Z(n19989) );
  ANDN U23969 ( .B(n19994), .A(n15360), .Z(n19992) );
  XNOR U23970 ( .A(a[121]), .B(n19995), .Z(n15360) );
  IV U23971 ( .A(n19993), .Z(n19995) );
  XNOR U23972 ( .A(b[121]), .B(n19993), .Z(n19994) );
  XOR U23973 ( .A(n19996), .B(n19997), .Z(n19993) );
  ANDN U23974 ( .B(n19998), .A(n15411), .Z(n19996) );
  XNOR U23975 ( .A(a[120]), .B(n19999), .Z(n15411) );
  IV U23976 ( .A(n19997), .Z(n19999) );
  XNOR U23977 ( .A(b[120]), .B(n19997), .Z(n19998) );
  XOR U23978 ( .A(n20000), .B(n20001), .Z(n19997) );
  ANDN U23979 ( .B(n20002), .A(n15463), .Z(n20000) );
  XNOR U23980 ( .A(a[119]), .B(n20003), .Z(n15463) );
  IV U23981 ( .A(n20001), .Z(n20003) );
  XNOR U23982 ( .A(b[119]), .B(n20001), .Z(n20002) );
  XOR U23983 ( .A(n20004), .B(n20005), .Z(n20001) );
  ANDN U23984 ( .B(n20006), .A(n15514), .Z(n20004) );
  XNOR U23985 ( .A(a[118]), .B(n20007), .Z(n15514) );
  IV U23986 ( .A(n20005), .Z(n20007) );
  XNOR U23987 ( .A(b[118]), .B(n20005), .Z(n20006) );
  XOR U23988 ( .A(n20008), .B(n20009), .Z(n20005) );
  ANDN U23989 ( .B(n20010), .A(n15565), .Z(n20008) );
  XNOR U23990 ( .A(a[117]), .B(n20011), .Z(n15565) );
  IV U23991 ( .A(n20009), .Z(n20011) );
  XNOR U23992 ( .A(b[117]), .B(n20009), .Z(n20010) );
  XOR U23993 ( .A(n20012), .B(n20013), .Z(n20009) );
  ANDN U23994 ( .B(n20014), .A(n15616), .Z(n20012) );
  XNOR U23995 ( .A(a[116]), .B(n20015), .Z(n15616) );
  IV U23996 ( .A(n20013), .Z(n20015) );
  XNOR U23997 ( .A(b[116]), .B(n20013), .Z(n20014) );
  XOR U23998 ( .A(n20016), .B(n20017), .Z(n20013) );
  ANDN U23999 ( .B(n20018), .A(n15667), .Z(n20016) );
  XNOR U24000 ( .A(a[115]), .B(n20019), .Z(n15667) );
  IV U24001 ( .A(n20017), .Z(n20019) );
  XNOR U24002 ( .A(b[115]), .B(n20017), .Z(n20018) );
  XOR U24003 ( .A(n20020), .B(n20021), .Z(n20017) );
  ANDN U24004 ( .B(n20022), .A(n15718), .Z(n20020) );
  XNOR U24005 ( .A(a[114]), .B(n20023), .Z(n15718) );
  IV U24006 ( .A(n20021), .Z(n20023) );
  XNOR U24007 ( .A(b[114]), .B(n20021), .Z(n20022) );
  XOR U24008 ( .A(n20024), .B(n20025), .Z(n20021) );
  ANDN U24009 ( .B(n20026), .A(n15769), .Z(n20024) );
  XNOR U24010 ( .A(a[113]), .B(n20027), .Z(n15769) );
  IV U24011 ( .A(n20025), .Z(n20027) );
  XNOR U24012 ( .A(b[113]), .B(n20025), .Z(n20026) );
  XOR U24013 ( .A(n20028), .B(n20029), .Z(n20025) );
  ANDN U24014 ( .B(n20030), .A(n15820), .Z(n20028) );
  XNOR U24015 ( .A(a[112]), .B(n20031), .Z(n15820) );
  IV U24016 ( .A(n20029), .Z(n20031) );
  XNOR U24017 ( .A(b[112]), .B(n20029), .Z(n20030) );
  XOR U24018 ( .A(n20032), .B(n20033), .Z(n20029) );
  ANDN U24019 ( .B(n20034), .A(n15871), .Z(n20032) );
  XNOR U24020 ( .A(a[111]), .B(n20035), .Z(n15871) );
  IV U24021 ( .A(n20033), .Z(n20035) );
  XNOR U24022 ( .A(b[111]), .B(n20033), .Z(n20034) );
  XOR U24023 ( .A(n20036), .B(n20037), .Z(n20033) );
  ANDN U24024 ( .B(n20038), .A(n15922), .Z(n20036) );
  XNOR U24025 ( .A(a[110]), .B(n20039), .Z(n15922) );
  IV U24026 ( .A(n20037), .Z(n20039) );
  XNOR U24027 ( .A(b[110]), .B(n20037), .Z(n20038) );
  XOR U24028 ( .A(n20040), .B(n20041), .Z(n20037) );
  ANDN U24029 ( .B(n20042), .A(n15974), .Z(n20040) );
  XNOR U24030 ( .A(a[109]), .B(n20043), .Z(n15974) );
  IV U24031 ( .A(n20041), .Z(n20043) );
  XNOR U24032 ( .A(b[109]), .B(n20041), .Z(n20042) );
  XOR U24033 ( .A(n20044), .B(n20045), .Z(n20041) );
  ANDN U24034 ( .B(n20046), .A(n16025), .Z(n20044) );
  XNOR U24035 ( .A(a[108]), .B(n20047), .Z(n16025) );
  IV U24036 ( .A(n20045), .Z(n20047) );
  XNOR U24037 ( .A(b[108]), .B(n20045), .Z(n20046) );
  XOR U24038 ( .A(n20048), .B(n20049), .Z(n20045) );
  ANDN U24039 ( .B(n20050), .A(n16076), .Z(n20048) );
  XNOR U24040 ( .A(a[107]), .B(n20051), .Z(n16076) );
  IV U24041 ( .A(n20049), .Z(n20051) );
  XNOR U24042 ( .A(b[107]), .B(n20049), .Z(n20050) );
  XOR U24043 ( .A(n20052), .B(n20053), .Z(n20049) );
  ANDN U24044 ( .B(n20054), .A(n16127), .Z(n20052) );
  XNOR U24045 ( .A(a[106]), .B(n20055), .Z(n16127) );
  IV U24046 ( .A(n20053), .Z(n20055) );
  XNOR U24047 ( .A(b[106]), .B(n20053), .Z(n20054) );
  XOR U24048 ( .A(n20056), .B(n20057), .Z(n20053) );
  ANDN U24049 ( .B(n20058), .A(n16178), .Z(n20056) );
  XNOR U24050 ( .A(a[105]), .B(n20059), .Z(n16178) );
  IV U24051 ( .A(n20057), .Z(n20059) );
  XNOR U24052 ( .A(b[105]), .B(n20057), .Z(n20058) );
  XOR U24053 ( .A(n20060), .B(n20061), .Z(n20057) );
  ANDN U24054 ( .B(n20062), .A(n16229), .Z(n20060) );
  XNOR U24055 ( .A(a[104]), .B(n20063), .Z(n16229) );
  IV U24056 ( .A(n20061), .Z(n20063) );
  XNOR U24057 ( .A(b[104]), .B(n20061), .Z(n20062) );
  XOR U24058 ( .A(n20064), .B(n20065), .Z(n20061) );
  ANDN U24059 ( .B(n20066), .A(n16280), .Z(n20064) );
  XNOR U24060 ( .A(a[103]), .B(n20067), .Z(n16280) );
  IV U24061 ( .A(n20065), .Z(n20067) );
  XNOR U24062 ( .A(b[103]), .B(n20065), .Z(n20066) );
  XOR U24063 ( .A(n20068), .B(n20069), .Z(n20065) );
  ANDN U24064 ( .B(n20070), .A(n16331), .Z(n20068) );
  XNOR U24065 ( .A(a[102]), .B(n20071), .Z(n16331) );
  IV U24066 ( .A(n20069), .Z(n20071) );
  XNOR U24067 ( .A(b[102]), .B(n20069), .Z(n20070) );
  XOR U24068 ( .A(n20072), .B(n20073), .Z(n20069) );
  ANDN U24069 ( .B(n20074), .A(n16382), .Z(n20072) );
  XNOR U24070 ( .A(a[101]), .B(n20075), .Z(n16382) );
  IV U24071 ( .A(n20073), .Z(n20075) );
  XNOR U24072 ( .A(b[101]), .B(n20073), .Z(n20074) );
  XOR U24073 ( .A(n20076), .B(n20077), .Z(n20073) );
  ANDN U24074 ( .B(n20078), .A(n16433), .Z(n20076) );
  XNOR U24075 ( .A(a[100]), .B(n20079), .Z(n16433) );
  IV U24076 ( .A(n20077), .Z(n20079) );
  XNOR U24077 ( .A(b[100]), .B(n20077), .Z(n20078) );
  XOR U24078 ( .A(n20080), .B(n20081), .Z(n20077) );
  ANDN U24079 ( .B(n20082), .A(n7), .Z(n20080) );
  XNOR U24080 ( .A(a[99]), .B(n20083), .Z(n7) );
  IV U24081 ( .A(n20081), .Z(n20083) );
  XNOR U24082 ( .A(b[99]), .B(n20081), .Z(n20082) );
  XOR U24083 ( .A(n20084), .B(n20085), .Z(n20081) );
  ANDN U24084 ( .B(n20086), .A(n18), .Z(n20084) );
  XNOR U24085 ( .A(a[98]), .B(n20087), .Z(n18) );
  IV U24086 ( .A(n20085), .Z(n20087) );
  XNOR U24087 ( .A(b[98]), .B(n20085), .Z(n20086) );
  XOR U24088 ( .A(n20088), .B(n20089), .Z(n20085) );
  ANDN U24089 ( .B(n20090), .A(n29), .Z(n20088) );
  XNOR U24090 ( .A(a[97]), .B(n20091), .Z(n29) );
  IV U24091 ( .A(n20089), .Z(n20091) );
  XNOR U24092 ( .A(b[97]), .B(n20089), .Z(n20090) );
  XOR U24093 ( .A(n20092), .B(n20093), .Z(n20089) );
  ANDN U24094 ( .B(n20094), .A(n40), .Z(n20092) );
  XNOR U24095 ( .A(a[96]), .B(n20095), .Z(n40) );
  IV U24096 ( .A(n20093), .Z(n20095) );
  XNOR U24097 ( .A(b[96]), .B(n20093), .Z(n20094) );
  XOR U24098 ( .A(n20096), .B(n20097), .Z(n20093) );
  ANDN U24099 ( .B(n20098), .A(n51), .Z(n20096) );
  XNOR U24100 ( .A(a[95]), .B(n20099), .Z(n51) );
  IV U24101 ( .A(n20097), .Z(n20099) );
  XNOR U24102 ( .A(b[95]), .B(n20097), .Z(n20098) );
  XOR U24103 ( .A(n20100), .B(n20101), .Z(n20097) );
  ANDN U24104 ( .B(n20102), .A(n62), .Z(n20100) );
  XNOR U24105 ( .A(a[94]), .B(n20103), .Z(n62) );
  IV U24106 ( .A(n20101), .Z(n20103) );
  XNOR U24107 ( .A(b[94]), .B(n20101), .Z(n20102) );
  XOR U24108 ( .A(n20104), .B(n20105), .Z(n20101) );
  ANDN U24109 ( .B(n20106), .A(n73), .Z(n20104) );
  XNOR U24110 ( .A(a[93]), .B(n20107), .Z(n73) );
  IV U24111 ( .A(n20105), .Z(n20107) );
  XNOR U24112 ( .A(b[93]), .B(n20105), .Z(n20106) );
  XOR U24113 ( .A(n20108), .B(n20109), .Z(n20105) );
  ANDN U24114 ( .B(n20110), .A(n84), .Z(n20108) );
  XNOR U24115 ( .A(a[92]), .B(n20111), .Z(n84) );
  IV U24116 ( .A(n20109), .Z(n20111) );
  XNOR U24117 ( .A(b[92]), .B(n20109), .Z(n20110) );
  XOR U24118 ( .A(n20112), .B(n20113), .Z(n20109) );
  ANDN U24119 ( .B(n20114), .A(n95), .Z(n20112) );
  XNOR U24120 ( .A(a[91]), .B(n20115), .Z(n95) );
  IV U24121 ( .A(n20113), .Z(n20115) );
  XNOR U24122 ( .A(b[91]), .B(n20113), .Z(n20114) );
  XOR U24123 ( .A(n20116), .B(n20117), .Z(n20113) );
  ANDN U24124 ( .B(n20118), .A(n106), .Z(n20116) );
  XNOR U24125 ( .A(a[90]), .B(n20119), .Z(n106) );
  IV U24126 ( .A(n20117), .Z(n20119) );
  XNOR U24127 ( .A(b[90]), .B(n20117), .Z(n20118) );
  XOR U24128 ( .A(n20120), .B(n20121), .Z(n20117) );
  ANDN U24129 ( .B(n20122), .A(n118), .Z(n20120) );
  XNOR U24130 ( .A(a[89]), .B(n20123), .Z(n118) );
  IV U24131 ( .A(n20121), .Z(n20123) );
  XNOR U24132 ( .A(b[89]), .B(n20121), .Z(n20122) );
  XOR U24133 ( .A(n20124), .B(n20125), .Z(n20121) );
  ANDN U24134 ( .B(n20126), .A(n129), .Z(n20124) );
  XNOR U24135 ( .A(a[88]), .B(n20127), .Z(n129) );
  IV U24136 ( .A(n20125), .Z(n20127) );
  XNOR U24137 ( .A(b[88]), .B(n20125), .Z(n20126) );
  XOR U24138 ( .A(n20128), .B(n20129), .Z(n20125) );
  ANDN U24139 ( .B(n20130), .A(n140), .Z(n20128) );
  XNOR U24140 ( .A(a[87]), .B(n20131), .Z(n140) );
  IV U24141 ( .A(n20129), .Z(n20131) );
  XNOR U24142 ( .A(b[87]), .B(n20129), .Z(n20130) );
  XOR U24143 ( .A(n20132), .B(n20133), .Z(n20129) );
  ANDN U24144 ( .B(n20134), .A(n151), .Z(n20132) );
  XNOR U24145 ( .A(a[86]), .B(n20135), .Z(n151) );
  IV U24146 ( .A(n20133), .Z(n20135) );
  XNOR U24147 ( .A(b[86]), .B(n20133), .Z(n20134) );
  XOR U24148 ( .A(n20136), .B(n20137), .Z(n20133) );
  ANDN U24149 ( .B(n20138), .A(n162), .Z(n20136) );
  XNOR U24150 ( .A(a[85]), .B(n20139), .Z(n162) );
  IV U24151 ( .A(n20137), .Z(n20139) );
  XNOR U24152 ( .A(b[85]), .B(n20137), .Z(n20138) );
  XOR U24153 ( .A(n20140), .B(n20141), .Z(n20137) );
  ANDN U24154 ( .B(n20142), .A(n173), .Z(n20140) );
  XNOR U24155 ( .A(a[84]), .B(n20143), .Z(n173) );
  IV U24156 ( .A(n20141), .Z(n20143) );
  XNOR U24157 ( .A(b[84]), .B(n20141), .Z(n20142) );
  XOR U24158 ( .A(n20144), .B(n20145), .Z(n20141) );
  ANDN U24159 ( .B(n20146), .A(n184), .Z(n20144) );
  XNOR U24160 ( .A(a[83]), .B(n20147), .Z(n184) );
  IV U24161 ( .A(n20145), .Z(n20147) );
  XNOR U24162 ( .A(b[83]), .B(n20145), .Z(n20146) );
  XOR U24163 ( .A(n20148), .B(n20149), .Z(n20145) );
  ANDN U24164 ( .B(n20150), .A(n195), .Z(n20148) );
  XNOR U24165 ( .A(a[82]), .B(n20151), .Z(n195) );
  IV U24166 ( .A(n20149), .Z(n20151) );
  XNOR U24167 ( .A(b[82]), .B(n20149), .Z(n20150) );
  XOR U24168 ( .A(n20152), .B(n20153), .Z(n20149) );
  ANDN U24169 ( .B(n20154), .A(n206), .Z(n20152) );
  XNOR U24170 ( .A(a[81]), .B(n20155), .Z(n206) );
  IV U24171 ( .A(n20153), .Z(n20155) );
  XNOR U24172 ( .A(b[81]), .B(n20153), .Z(n20154) );
  XOR U24173 ( .A(n20156), .B(n20157), .Z(n20153) );
  ANDN U24174 ( .B(n20158), .A(n217), .Z(n20156) );
  XNOR U24175 ( .A(a[80]), .B(n20159), .Z(n217) );
  IV U24176 ( .A(n20157), .Z(n20159) );
  XNOR U24177 ( .A(b[80]), .B(n20157), .Z(n20158) );
  XOR U24178 ( .A(n20160), .B(n20161), .Z(n20157) );
  ANDN U24179 ( .B(n20162), .A(n229), .Z(n20160) );
  XNOR U24180 ( .A(a[79]), .B(n20163), .Z(n229) );
  IV U24181 ( .A(n20161), .Z(n20163) );
  XNOR U24182 ( .A(b[79]), .B(n20161), .Z(n20162) );
  XOR U24183 ( .A(n20164), .B(n20165), .Z(n20161) );
  ANDN U24184 ( .B(n20166), .A(n240), .Z(n20164) );
  XNOR U24185 ( .A(a[78]), .B(n20167), .Z(n240) );
  IV U24186 ( .A(n20165), .Z(n20167) );
  XNOR U24187 ( .A(b[78]), .B(n20165), .Z(n20166) );
  XOR U24188 ( .A(n20168), .B(n20169), .Z(n20165) );
  ANDN U24189 ( .B(n20170), .A(n251), .Z(n20168) );
  XNOR U24190 ( .A(a[77]), .B(n20171), .Z(n251) );
  IV U24191 ( .A(n20169), .Z(n20171) );
  XNOR U24192 ( .A(b[77]), .B(n20169), .Z(n20170) );
  XOR U24193 ( .A(n20172), .B(n20173), .Z(n20169) );
  ANDN U24194 ( .B(n20174), .A(n262), .Z(n20172) );
  XNOR U24195 ( .A(a[76]), .B(n20175), .Z(n262) );
  IV U24196 ( .A(n20173), .Z(n20175) );
  XNOR U24197 ( .A(b[76]), .B(n20173), .Z(n20174) );
  XOR U24198 ( .A(n20176), .B(n20177), .Z(n20173) );
  ANDN U24199 ( .B(n20178), .A(n273), .Z(n20176) );
  XNOR U24200 ( .A(a[75]), .B(n20179), .Z(n273) );
  IV U24201 ( .A(n20177), .Z(n20179) );
  XNOR U24202 ( .A(b[75]), .B(n20177), .Z(n20178) );
  XOR U24203 ( .A(n20180), .B(n20181), .Z(n20177) );
  ANDN U24204 ( .B(n20182), .A(n284), .Z(n20180) );
  XNOR U24205 ( .A(a[74]), .B(n20183), .Z(n284) );
  IV U24206 ( .A(n20181), .Z(n20183) );
  XNOR U24207 ( .A(b[74]), .B(n20181), .Z(n20182) );
  XOR U24208 ( .A(n20184), .B(n20185), .Z(n20181) );
  ANDN U24209 ( .B(n20186), .A(n295), .Z(n20184) );
  XNOR U24210 ( .A(a[73]), .B(n20187), .Z(n295) );
  IV U24211 ( .A(n20185), .Z(n20187) );
  XNOR U24212 ( .A(b[73]), .B(n20185), .Z(n20186) );
  XOR U24213 ( .A(n20188), .B(n20189), .Z(n20185) );
  ANDN U24214 ( .B(n20190), .A(n306), .Z(n20188) );
  XNOR U24215 ( .A(a[72]), .B(n20191), .Z(n306) );
  IV U24216 ( .A(n20189), .Z(n20191) );
  XNOR U24217 ( .A(b[72]), .B(n20189), .Z(n20190) );
  XOR U24218 ( .A(n20192), .B(n20193), .Z(n20189) );
  ANDN U24219 ( .B(n20194), .A(n317), .Z(n20192) );
  XNOR U24220 ( .A(a[71]), .B(n20195), .Z(n317) );
  IV U24221 ( .A(n20193), .Z(n20195) );
  XNOR U24222 ( .A(b[71]), .B(n20193), .Z(n20194) );
  XOR U24223 ( .A(n20196), .B(n20197), .Z(n20193) );
  ANDN U24224 ( .B(n20198), .A(n328), .Z(n20196) );
  XNOR U24225 ( .A(a[70]), .B(n20199), .Z(n328) );
  IV U24226 ( .A(n20197), .Z(n20199) );
  XNOR U24227 ( .A(b[70]), .B(n20197), .Z(n20198) );
  XOR U24228 ( .A(n20200), .B(n20201), .Z(n20197) );
  ANDN U24229 ( .B(n20202), .A(n340), .Z(n20200) );
  XNOR U24230 ( .A(a[69]), .B(n20203), .Z(n340) );
  IV U24231 ( .A(n20201), .Z(n20203) );
  XNOR U24232 ( .A(b[69]), .B(n20201), .Z(n20202) );
  XOR U24233 ( .A(n20204), .B(n20205), .Z(n20201) );
  ANDN U24234 ( .B(n20206), .A(n351), .Z(n20204) );
  XNOR U24235 ( .A(a[68]), .B(n20207), .Z(n351) );
  IV U24236 ( .A(n20205), .Z(n20207) );
  XNOR U24237 ( .A(b[68]), .B(n20205), .Z(n20206) );
  XOR U24238 ( .A(n20208), .B(n20209), .Z(n20205) );
  ANDN U24239 ( .B(n20210), .A(n362), .Z(n20208) );
  XNOR U24240 ( .A(a[67]), .B(n20211), .Z(n362) );
  IV U24241 ( .A(n20209), .Z(n20211) );
  XNOR U24242 ( .A(b[67]), .B(n20209), .Z(n20210) );
  XOR U24243 ( .A(n20212), .B(n20213), .Z(n20209) );
  ANDN U24244 ( .B(n20214), .A(n373), .Z(n20212) );
  XNOR U24245 ( .A(a[66]), .B(n20215), .Z(n373) );
  IV U24246 ( .A(n20213), .Z(n20215) );
  XNOR U24247 ( .A(b[66]), .B(n20213), .Z(n20214) );
  XOR U24248 ( .A(n20216), .B(n20217), .Z(n20213) );
  ANDN U24249 ( .B(n20218), .A(n384), .Z(n20216) );
  XNOR U24250 ( .A(a[65]), .B(n20219), .Z(n384) );
  IV U24251 ( .A(n20217), .Z(n20219) );
  XNOR U24252 ( .A(b[65]), .B(n20217), .Z(n20218) );
  XOR U24253 ( .A(n20220), .B(n20221), .Z(n20217) );
  ANDN U24254 ( .B(n20222), .A(n395), .Z(n20220) );
  XNOR U24255 ( .A(a[64]), .B(n20223), .Z(n395) );
  IV U24256 ( .A(n20221), .Z(n20223) );
  XNOR U24257 ( .A(b[64]), .B(n20221), .Z(n20222) );
  XOR U24258 ( .A(n20224), .B(n20225), .Z(n20221) );
  ANDN U24259 ( .B(n20226), .A(n406), .Z(n20224) );
  XNOR U24260 ( .A(a[63]), .B(n20227), .Z(n406) );
  IV U24261 ( .A(n20225), .Z(n20227) );
  XNOR U24262 ( .A(b[63]), .B(n20225), .Z(n20226) );
  XOR U24263 ( .A(n20228), .B(n20229), .Z(n20225) );
  ANDN U24264 ( .B(n20230), .A(n417), .Z(n20228) );
  XNOR U24265 ( .A(a[62]), .B(n20231), .Z(n417) );
  IV U24266 ( .A(n20229), .Z(n20231) );
  XNOR U24267 ( .A(b[62]), .B(n20229), .Z(n20230) );
  XOR U24268 ( .A(n20232), .B(n20233), .Z(n20229) );
  ANDN U24269 ( .B(n20234), .A(n428), .Z(n20232) );
  XNOR U24270 ( .A(a[61]), .B(n20235), .Z(n428) );
  IV U24271 ( .A(n20233), .Z(n20235) );
  XNOR U24272 ( .A(b[61]), .B(n20233), .Z(n20234) );
  XOR U24273 ( .A(n20236), .B(n20237), .Z(n20233) );
  ANDN U24274 ( .B(n20238), .A(n439), .Z(n20236) );
  XNOR U24275 ( .A(a[60]), .B(n20239), .Z(n439) );
  IV U24276 ( .A(n20237), .Z(n20239) );
  XNOR U24277 ( .A(b[60]), .B(n20237), .Z(n20238) );
  XOR U24278 ( .A(n20240), .B(n20241), .Z(n20237) );
  ANDN U24279 ( .B(n20242), .A(n451), .Z(n20240) );
  XNOR U24280 ( .A(a[59]), .B(n20243), .Z(n451) );
  IV U24281 ( .A(n20241), .Z(n20243) );
  XNOR U24282 ( .A(b[59]), .B(n20241), .Z(n20242) );
  XOR U24283 ( .A(n20244), .B(n20245), .Z(n20241) );
  ANDN U24284 ( .B(n20246), .A(n462), .Z(n20244) );
  XNOR U24285 ( .A(a[58]), .B(n20247), .Z(n462) );
  IV U24286 ( .A(n20245), .Z(n20247) );
  XNOR U24287 ( .A(b[58]), .B(n20245), .Z(n20246) );
  XOR U24288 ( .A(n20248), .B(n20249), .Z(n20245) );
  ANDN U24289 ( .B(n20250), .A(n473), .Z(n20248) );
  XNOR U24290 ( .A(a[57]), .B(n20251), .Z(n473) );
  IV U24291 ( .A(n20249), .Z(n20251) );
  XNOR U24292 ( .A(b[57]), .B(n20249), .Z(n20250) );
  XOR U24293 ( .A(n20252), .B(n20253), .Z(n20249) );
  ANDN U24294 ( .B(n20254), .A(n484), .Z(n20252) );
  XNOR U24295 ( .A(a[56]), .B(n20255), .Z(n484) );
  IV U24296 ( .A(n20253), .Z(n20255) );
  XNOR U24297 ( .A(b[56]), .B(n20253), .Z(n20254) );
  XOR U24298 ( .A(n20256), .B(n20257), .Z(n20253) );
  ANDN U24299 ( .B(n20258), .A(n495), .Z(n20256) );
  XNOR U24300 ( .A(a[55]), .B(n20259), .Z(n495) );
  IV U24301 ( .A(n20257), .Z(n20259) );
  XNOR U24302 ( .A(b[55]), .B(n20257), .Z(n20258) );
  XOR U24303 ( .A(n20260), .B(n20261), .Z(n20257) );
  ANDN U24304 ( .B(n20262), .A(n506), .Z(n20260) );
  XNOR U24305 ( .A(a[54]), .B(n20263), .Z(n506) );
  IV U24306 ( .A(n20261), .Z(n20263) );
  XNOR U24307 ( .A(b[54]), .B(n20261), .Z(n20262) );
  XOR U24308 ( .A(n20264), .B(n20265), .Z(n20261) );
  ANDN U24309 ( .B(n20266), .A(n517), .Z(n20264) );
  XNOR U24310 ( .A(a[53]), .B(n20267), .Z(n517) );
  IV U24311 ( .A(n20265), .Z(n20267) );
  XNOR U24312 ( .A(b[53]), .B(n20265), .Z(n20266) );
  XOR U24313 ( .A(n20268), .B(n20269), .Z(n20265) );
  ANDN U24314 ( .B(n20270), .A(n528), .Z(n20268) );
  XNOR U24315 ( .A(a[52]), .B(n20271), .Z(n528) );
  IV U24316 ( .A(n20269), .Z(n20271) );
  XNOR U24317 ( .A(b[52]), .B(n20269), .Z(n20270) );
  XOR U24318 ( .A(n20272), .B(n20273), .Z(n20269) );
  ANDN U24319 ( .B(n20274), .A(n539), .Z(n20272) );
  XNOR U24320 ( .A(a[51]), .B(n20275), .Z(n539) );
  IV U24321 ( .A(n20273), .Z(n20275) );
  XNOR U24322 ( .A(b[51]), .B(n20273), .Z(n20274) );
  XOR U24323 ( .A(n20276), .B(n20277), .Z(n20273) );
  ANDN U24324 ( .B(n20278), .A(n550), .Z(n20276) );
  XNOR U24325 ( .A(a[50]), .B(n20279), .Z(n550) );
  IV U24326 ( .A(n20277), .Z(n20279) );
  XNOR U24327 ( .A(b[50]), .B(n20277), .Z(n20278) );
  XOR U24328 ( .A(n20280), .B(n20281), .Z(n20277) );
  ANDN U24329 ( .B(n20282), .A(n562), .Z(n20280) );
  XNOR U24330 ( .A(a[49]), .B(n20283), .Z(n562) );
  IV U24331 ( .A(n20281), .Z(n20283) );
  XNOR U24332 ( .A(b[49]), .B(n20281), .Z(n20282) );
  XOR U24333 ( .A(n20284), .B(n20285), .Z(n20281) );
  ANDN U24334 ( .B(n20286), .A(n573), .Z(n20284) );
  XNOR U24335 ( .A(a[48]), .B(n20287), .Z(n573) );
  IV U24336 ( .A(n20285), .Z(n20287) );
  XNOR U24337 ( .A(b[48]), .B(n20285), .Z(n20286) );
  XOR U24338 ( .A(n20288), .B(n20289), .Z(n20285) );
  ANDN U24339 ( .B(n20290), .A(n584), .Z(n20288) );
  XNOR U24340 ( .A(a[47]), .B(n20291), .Z(n584) );
  IV U24341 ( .A(n20289), .Z(n20291) );
  XNOR U24342 ( .A(b[47]), .B(n20289), .Z(n20290) );
  XOR U24343 ( .A(n20292), .B(n20293), .Z(n20289) );
  ANDN U24344 ( .B(n20294), .A(n595), .Z(n20292) );
  XNOR U24345 ( .A(a[46]), .B(n20295), .Z(n595) );
  IV U24346 ( .A(n20293), .Z(n20295) );
  XNOR U24347 ( .A(b[46]), .B(n20293), .Z(n20294) );
  XOR U24348 ( .A(n20296), .B(n20297), .Z(n20293) );
  ANDN U24349 ( .B(n20298), .A(n606), .Z(n20296) );
  XNOR U24350 ( .A(a[45]), .B(n20299), .Z(n606) );
  IV U24351 ( .A(n20297), .Z(n20299) );
  XNOR U24352 ( .A(b[45]), .B(n20297), .Z(n20298) );
  XOR U24353 ( .A(n20300), .B(n20301), .Z(n20297) );
  ANDN U24354 ( .B(n20302), .A(n617), .Z(n20300) );
  XNOR U24355 ( .A(a[44]), .B(n20303), .Z(n617) );
  IV U24356 ( .A(n20301), .Z(n20303) );
  XNOR U24357 ( .A(b[44]), .B(n20301), .Z(n20302) );
  XOR U24358 ( .A(n20304), .B(n20305), .Z(n20301) );
  ANDN U24359 ( .B(n20306), .A(n628), .Z(n20304) );
  XNOR U24360 ( .A(a[43]), .B(n20307), .Z(n628) );
  IV U24361 ( .A(n20305), .Z(n20307) );
  XNOR U24362 ( .A(b[43]), .B(n20305), .Z(n20306) );
  XOR U24363 ( .A(n20308), .B(n20309), .Z(n20305) );
  ANDN U24364 ( .B(n20310), .A(n639), .Z(n20308) );
  XNOR U24365 ( .A(a[42]), .B(n20311), .Z(n639) );
  IV U24366 ( .A(n20309), .Z(n20311) );
  XNOR U24367 ( .A(b[42]), .B(n20309), .Z(n20310) );
  XOR U24368 ( .A(n20312), .B(n20313), .Z(n20309) );
  ANDN U24369 ( .B(n20314), .A(n650), .Z(n20312) );
  XNOR U24370 ( .A(a[41]), .B(n20315), .Z(n650) );
  IV U24371 ( .A(n20313), .Z(n20315) );
  XNOR U24372 ( .A(b[41]), .B(n20313), .Z(n20314) );
  XOR U24373 ( .A(n20316), .B(n20317), .Z(n20313) );
  ANDN U24374 ( .B(n20318), .A(n661), .Z(n20316) );
  XNOR U24375 ( .A(a[40]), .B(n20319), .Z(n661) );
  IV U24376 ( .A(n20317), .Z(n20319) );
  XNOR U24377 ( .A(b[40]), .B(n20317), .Z(n20318) );
  XOR U24378 ( .A(n20320), .B(n20321), .Z(n20317) );
  ANDN U24379 ( .B(n20322), .A(n1152), .Z(n20320) );
  XNOR U24380 ( .A(a[39]), .B(n20323), .Z(n1152) );
  IV U24381 ( .A(n20321), .Z(n20323) );
  XNOR U24382 ( .A(b[39]), .B(n20321), .Z(n20322) );
  XOR U24383 ( .A(n20324), .B(n20325), .Z(n20321) );
  ANDN U24384 ( .B(n20326), .A(n1663), .Z(n20324) );
  XNOR U24385 ( .A(a[38]), .B(n20327), .Z(n1663) );
  IV U24386 ( .A(n20325), .Z(n20327) );
  XNOR U24387 ( .A(b[38]), .B(n20325), .Z(n20326) );
  XOR U24388 ( .A(n20328), .B(n20329), .Z(n20325) );
  ANDN U24389 ( .B(n20330), .A(n2174), .Z(n20328) );
  XNOR U24390 ( .A(a[37]), .B(n20331), .Z(n2174) );
  IV U24391 ( .A(n20329), .Z(n20331) );
  XNOR U24392 ( .A(b[37]), .B(n20329), .Z(n20330) );
  XOR U24393 ( .A(n20332), .B(n20333), .Z(n20329) );
  ANDN U24394 ( .B(n20334), .A(n2685), .Z(n20332) );
  XNOR U24395 ( .A(a[36]), .B(n20335), .Z(n2685) );
  IV U24396 ( .A(n20333), .Z(n20335) );
  XNOR U24397 ( .A(b[36]), .B(n20333), .Z(n20334) );
  XOR U24398 ( .A(n20336), .B(n20337), .Z(n20333) );
  ANDN U24399 ( .B(n20338), .A(n3196), .Z(n20336) );
  XNOR U24400 ( .A(a[35]), .B(n20339), .Z(n3196) );
  IV U24401 ( .A(n20337), .Z(n20339) );
  XNOR U24402 ( .A(b[35]), .B(n20337), .Z(n20338) );
  XOR U24403 ( .A(n20340), .B(n20341), .Z(n20337) );
  ANDN U24404 ( .B(n20342), .A(n3707), .Z(n20340) );
  XNOR U24405 ( .A(a[34]), .B(n20343), .Z(n3707) );
  IV U24406 ( .A(n20341), .Z(n20343) );
  XNOR U24407 ( .A(b[34]), .B(n20341), .Z(n20342) );
  XOR U24408 ( .A(n20344), .B(n20345), .Z(n20341) );
  ANDN U24409 ( .B(n20346), .A(n4218), .Z(n20344) );
  XNOR U24410 ( .A(a[33]), .B(n20347), .Z(n4218) );
  IV U24411 ( .A(n20345), .Z(n20347) );
  XNOR U24412 ( .A(b[33]), .B(n20345), .Z(n20346) );
  XOR U24413 ( .A(n20348), .B(n20349), .Z(n20345) );
  ANDN U24414 ( .B(n20350), .A(n4729), .Z(n20348) );
  XNOR U24415 ( .A(a[32]), .B(n20351), .Z(n4729) );
  IV U24416 ( .A(n20349), .Z(n20351) );
  XNOR U24417 ( .A(b[32]), .B(n20349), .Z(n20350) );
  XOR U24418 ( .A(n20352), .B(n20353), .Z(n20349) );
  ANDN U24419 ( .B(n20354), .A(n5240), .Z(n20352) );
  XNOR U24420 ( .A(a[31]), .B(n20355), .Z(n5240) );
  IV U24421 ( .A(n20353), .Z(n20355) );
  XNOR U24422 ( .A(b[31]), .B(n20353), .Z(n20354) );
  XOR U24423 ( .A(n20356), .B(n20357), .Z(n20353) );
  ANDN U24424 ( .B(n20358), .A(n5751), .Z(n20356) );
  XNOR U24425 ( .A(a[30]), .B(n20359), .Z(n5751) );
  IV U24426 ( .A(n20357), .Z(n20359) );
  XNOR U24427 ( .A(b[30]), .B(n20357), .Z(n20358) );
  XOR U24428 ( .A(n20360), .B(n20361), .Z(n20357) );
  ANDN U24429 ( .B(n20362), .A(n6263), .Z(n20360) );
  XNOR U24430 ( .A(a[29]), .B(n20363), .Z(n6263) );
  IV U24431 ( .A(n20361), .Z(n20363) );
  XNOR U24432 ( .A(b[29]), .B(n20361), .Z(n20362) );
  XOR U24433 ( .A(n20364), .B(n20365), .Z(n20361) );
  ANDN U24434 ( .B(n20366), .A(n6774), .Z(n20364) );
  XNOR U24435 ( .A(a[28]), .B(n20367), .Z(n6774) );
  IV U24436 ( .A(n20365), .Z(n20367) );
  XNOR U24437 ( .A(b[28]), .B(n20365), .Z(n20366) );
  XOR U24438 ( .A(n20368), .B(n20369), .Z(n20365) );
  ANDN U24439 ( .B(n20370), .A(n7285), .Z(n20368) );
  XNOR U24440 ( .A(a[27]), .B(n20371), .Z(n7285) );
  IV U24441 ( .A(n20369), .Z(n20371) );
  XNOR U24442 ( .A(b[27]), .B(n20369), .Z(n20370) );
  XOR U24443 ( .A(n20372), .B(n20373), .Z(n20369) );
  ANDN U24444 ( .B(n20374), .A(n7796), .Z(n20372) );
  XNOR U24445 ( .A(a[26]), .B(n20375), .Z(n7796) );
  IV U24446 ( .A(n20373), .Z(n20375) );
  XNOR U24447 ( .A(b[26]), .B(n20373), .Z(n20374) );
  XOR U24448 ( .A(n20376), .B(n20377), .Z(n20373) );
  ANDN U24449 ( .B(n20378), .A(n8307), .Z(n20376) );
  XNOR U24450 ( .A(a[25]), .B(n20379), .Z(n8307) );
  IV U24451 ( .A(n20377), .Z(n20379) );
  XNOR U24452 ( .A(b[25]), .B(n20377), .Z(n20378) );
  XOR U24453 ( .A(n20380), .B(n20381), .Z(n20377) );
  ANDN U24454 ( .B(n20382), .A(n8818), .Z(n20380) );
  XNOR U24455 ( .A(a[24]), .B(n20383), .Z(n8818) );
  IV U24456 ( .A(n20381), .Z(n20383) );
  XNOR U24457 ( .A(b[24]), .B(n20381), .Z(n20382) );
  XOR U24458 ( .A(n20384), .B(n20385), .Z(n20381) );
  ANDN U24459 ( .B(n20386), .A(n9329), .Z(n20384) );
  XNOR U24460 ( .A(a[23]), .B(n20387), .Z(n9329) );
  IV U24461 ( .A(n20385), .Z(n20387) );
  XNOR U24462 ( .A(b[23]), .B(n20385), .Z(n20386) );
  XOR U24463 ( .A(n20388), .B(n20389), .Z(n20385) );
  ANDN U24464 ( .B(n20390), .A(n9840), .Z(n20388) );
  XNOR U24465 ( .A(a[22]), .B(n20391), .Z(n9840) );
  IV U24466 ( .A(n20389), .Z(n20391) );
  XNOR U24467 ( .A(b[22]), .B(n20389), .Z(n20390) );
  XOR U24468 ( .A(n20392), .B(n20393), .Z(n20389) );
  ANDN U24469 ( .B(n20394), .A(n10351), .Z(n20392) );
  XNOR U24470 ( .A(a[21]), .B(n20395), .Z(n10351) );
  IV U24471 ( .A(n20393), .Z(n20395) );
  XNOR U24472 ( .A(b[21]), .B(n20393), .Z(n20394) );
  XOR U24473 ( .A(n20396), .B(n20397), .Z(n20393) );
  ANDN U24474 ( .B(n20398), .A(n10862), .Z(n20396) );
  XNOR U24475 ( .A(a[20]), .B(n20399), .Z(n10862) );
  IV U24476 ( .A(n20397), .Z(n20399) );
  XNOR U24477 ( .A(b[20]), .B(n20397), .Z(n20398) );
  XOR U24478 ( .A(n20400), .B(n20401), .Z(n20397) );
  ANDN U24479 ( .B(n20402), .A(n11374), .Z(n20400) );
  XNOR U24480 ( .A(a[19]), .B(n20403), .Z(n11374) );
  IV U24481 ( .A(n20401), .Z(n20403) );
  XNOR U24482 ( .A(b[19]), .B(n20401), .Z(n20402) );
  XOR U24483 ( .A(n20404), .B(n20405), .Z(n20401) );
  ANDN U24484 ( .B(n20406), .A(n11885), .Z(n20404) );
  XNOR U24485 ( .A(a[18]), .B(n20407), .Z(n11885) );
  IV U24486 ( .A(n20405), .Z(n20407) );
  XNOR U24487 ( .A(b[18]), .B(n20405), .Z(n20406) );
  XOR U24488 ( .A(n20408), .B(n20409), .Z(n20405) );
  ANDN U24489 ( .B(n20410), .A(n12396), .Z(n20408) );
  XNOR U24490 ( .A(a[17]), .B(n20411), .Z(n12396) );
  IV U24491 ( .A(n20409), .Z(n20411) );
  XNOR U24492 ( .A(b[17]), .B(n20409), .Z(n20410) );
  XOR U24493 ( .A(n20412), .B(n20413), .Z(n20409) );
  ANDN U24494 ( .B(n20414), .A(n12907), .Z(n20412) );
  XNOR U24495 ( .A(a[16]), .B(n20415), .Z(n12907) );
  IV U24496 ( .A(n20413), .Z(n20415) );
  XNOR U24497 ( .A(b[16]), .B(n20413), .Z(n20414) );
  XOR U24498 ( .A(n20416), .B(n20417), .Z(n20413) );
  ANDN U24499 ( .B(n20418), .A(n13418), .Z(n20416) );
  XNOR U24500 ( .A(a[15]), .B(n20419), .Z(n13418) );
  IV U24501 ( .A(n20417), .Z(n20419) );
  XNOR U24502 ( .A(b[15]), .B(n20417), .Z(n20418) );
  XOR U24503 ( .A(n20420), .B(n20421), .Z(n20417) );
  ANDN U24504 ( .B(n20422), .A(n13929), .Z(n20420) );
  XNOR U24505 ( .A(a[14]), .B(n20423), .Z(n13929) );
  IV U24506 ( .A(n20421), .Z(n20423) );
  XNOR U24507 ( .A(b[14]), .B(n20421), .Z(n20422) );
  XOR U24508 ( .A(n20424), .B(n20425), .Z(n20421) );
  ANDN U24509 ( .B(n20426), .A(n14440), .Z(n20424) );
  XNOR U24510 ( .A(a[13]), .B(n20427), .Z(n14440) );
  IV U24511 ( .A(n20425), .Z(n20427) );
  XNOR U24512 ( .A(b[13]), .B(n20425), .Z(n20426) );
  XOR U24513 ( .A(n20428), .B(n20429), .Z(n20425) );
  ANDN U24514 ( .B(n20430), .A(n14951), .Z(n20428) );
  XNOR U24515 ( .A(a[12]), .B(n20431), .Z(n14951) );
  IV U24516 ( .A(n20429), .Z(n20431) );
  XNOR U24517 ( .A(b[12]), .B(n20429), .Z(n20430) );
  XOR U24518 ( .A(n20432), .B(n20433), .Z(n20429) );
  ANDN U24519 ( .B(n20434), .A(n15462), .Z(n20432) );
  XNOR U24520 ( .A(a[11]), .B(n20435), .Z(n15462) );
  IV U24521 ( .A(n20433), .Z(n20435) );
  XNOR U24522 ( .A(b[11]), .B(n20433), .Z(n20434) );
  XOR U24523 ( .A(n20436), .B(n20437), .Z(n20433) );
  ANDN U24524 ( .B(n20438), .A(n15973), .Z(n20436) );
  XNOR U24525 ( .A(a[10]), .B(n20439), .Z(n15973) );
  IV U24526 ( .A(n20437), .Z(n20439) );
  XNOR U24527 ( .A(b[10]), .B(n20437), .Z(n20438) );
  XOR U24528 ( .A(n20440), .B(n20441), .Z(n20437) );
  ANDN U24529 ( .B(n20442), .A(n6), .Z(n20440) );
  XNOR U24530 ( .A(a[9]), .B(n20443), .Z(n6) );
  IV U24531 ( .A(n20441), .Z(n20443) );
  XNOR U24532 ( .A(b[9]), .B(n20441), .Z(n20442) );
  XOR U24533 ( .A(n20444), .B(n20445), .Z(n20441) );
  ANDN U24534 ( .B(n20446), .A(n117), .Z(n20444) );
  XNOR U24535 ( .A(a[8]), .B(n20447), .Z(n117) );
  IV U24536 ( .A(n20445), .Z(n20447) );
  XNOR U24537 ( .A(b[8]), .B(n20445), .Z(n20446) );
  XOR U24538 ( .A(n20448), .B(n20449), .Z(n20445) );
  ANDN U24539 ( .B(n20450), .A(n228), .Z(n20448) );
  XNOR U24540 ( .A(a[7]), .B(n20451), .Z(n228) );
  IV U24541 ( .A(n20449), .Z(n20451) );
  XNOR U24542 ( .A(b[7]), .B(n20449), .Z(n20450) );
  XOR U24543 ( .A(n20452), .B(n20453), .Z(n20449) );
  ANDN U24544 ( .B(n20454), .A(n339), .Z(n20452) );
  XNOR U24545 ( .A(a[6]), .B(n20455), .Z(n339) );
  IV U24546 ( .A(n20453), .Z(n20455) );
  XNOR U24547 ( .A(b[6]), .B(n20453), .Z(n20454) );
  XOR U24548 ( .A(n20456), .B(n20457), .Z(n20453) );
  ANDN U24549 ( .B(n20458), .A(n450), .Z(n20456) );
  XNOR U24550 ( .A(a[5]), .B(n20459), .Z(n450) );
  IV U24551 ( .A(n20457), .Z(n20459) );
  XNOR U24552 ( .A(b[5]), .B(n20457), .Z(n20458) );
  XOR U24553 ( .A(n20460), .B(n20461), .Z(n20457) );
  ANDN U24554 ( .B(n20462), .A(n561), .Z(n20460) );
  XNOR U24555 ( .A(a[4]), .B(n20463), .Z(n561) );
  IV U24556 ( .A(n20461), .Z(n20463) );
  XNOR U24557 ( .A(b[4]), .B(n20461), .Z(n20462) );
  XOR U24558 ( .A(n20464), .B(n20465), .Z(n20461) );
  ANDN U24559 ( .B(n20466), .A(n1151), .Z(n20464) );
  XNOR U24560 ( .A(a[3]), .B(n20467), .Z(n1151) );
  IV U24561 ( .A(n20465), .Z(n20467) );
  XNOR U24562 ( .A(b[3]), .B(n20465), .Z(n20466) );
  XOR U24563 ( .A(n20468), .B(n20469), .Z(n20465) );
  ANDN U24564 ( .B(n20470), .A(n6262), .Z(n20468) );
  XNOR U24565 ( .A(a[2]), .B(n20471), .Z(n6262) );
  IV U24566 ( .A(n20469), .Z(n20471) );
  XNOR U24567 ( .A(b[2]), .B(n20469), .Z(n20470) );
  XOR U24568 ( .A(n20472), .B(n20473), .Z(n20469) );
  ANDN U24569 ( .B(n20474), .A(n11373), .Z(n20472) );
  XNOR U24570 ( .A(a[1]), .B(n20475), .Z(n11373) );
  IV U24571 ( .A(n20473), .Z(n20475) );
  XNOR U24572 ( .A(b[1]), .B(n20473), .Z(n20474) );
  XOR U24573 ( .A(carry_on), .B(n20476), .Z(n20473) );
  NANDN U24574 ( .A(n20477), .B(n20478), .Z(n20476) );
  XOR U24575 ( .A(carry_on), .B(b[0]), .Z(n20478) );
  XNOR U24576 ( .A(b[0]), .B(n20477), .Z(c[0]) );
  XNOR U24577 ( .A(a[0]), .B(carry_on), .Z(n20477) );
endmodule

