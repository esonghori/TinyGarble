
module modmult_step_N256_4 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506,
         N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517,
         N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528,
         N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539,
         N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550,
         N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561,
         N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572,
         N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583,
         N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594,
         N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605,
         N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616,
         N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627,
         N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638,
         N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649,
         N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660,
         N661, N662, N663, N664, N665, N666, N667, N668, N669, N670, N671,
         N672, N673, N674, N675, N676, N677, N678, N679, N680, N681, N682,
         N683, N684, N685, N686, N687, N688, N689, N690, N691, N692, N693,
         N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704,
         N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715,
         N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726,
         N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737,
         N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770,
         N771, N772, N773, N774, N775, N776, N777, N778, N779, N780;
  wire   [257:0] z2;
  wire   [257:0] z3;

  GT_UNS_OP gt_123 ( .A(z2), .B(n), .Z(N262) );
  GEQ_UNS_OP gte_128 ( .A(z3), .B(n), .Z(N522) );
  ADD_UNS_OP add_119 ( .A({zin[256:0], 1'b0}), .B(y), .Z({N261, N260, N259, 
        N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, 
        N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, 
        N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, 
        N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, 
        N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, 
        N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, 
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
        N4}) );
  SUB_UNS_OP sub_124 ( .A(z2), .B(n), .Z({N521, N520, N519, N518, N517, N516, 
        N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, 
        N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, 
        N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, 
        N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, 
        N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, 
        N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, 
        N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, 
        N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, 
        N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, 
        N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, 
        N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, 
        N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, 
        N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, 
        N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, 
        N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, 
        N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, 
        N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, 
        N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, 
        N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, 
        N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, 
        N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264}) );
  SUB_UNS_OP sub_129_aco ( .A(z3), .B({N780, N779, N778, N777, N776, N775, 
        N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, 
        N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, 
        N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, 
        N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, 
        N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, 
        N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, 
        N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, 
        N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, 
        N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, 
        N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, 
        N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, 
        N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, 
        N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, 
        N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, 
        N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, 
        N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, 
        N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, 
        N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, 
        N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, 
        N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, 
        N534, N533, N532, N531, N530, N529, N528, N527, N526, N525}), .Z(zout)
         );
  SELECT_OP C794 ( .DATA1({N261, N260, N259, N258, N257, N256, N255, N254, 
        N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, 
        N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, 
        N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, 
        N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, 
        N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, 
        N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, 
        N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, 
        N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, 
        N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, 
        N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, 
        N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, 
        N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, 
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, 
        N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, 
        N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}), .DATA2({zin[256:0], 1'b0}), .CONTROL1(N0), .CONTROL2(N1), .Z(z2) );
  GTECH_BUF B_0 ( .A(xregN_1), .Z(N0) );
  GTECH_BUF B_1 ( .A(N3), .Z(N1) );
  SELECT_OP C795 ( .DATA1({N521, N520, N519, N518, N517, N516, N515, N514, 
        N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, 
        N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, 
        N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, 
        N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, 
        N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, 
        N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, 
        N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, 
        N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, 
        N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, 
        N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, 
        N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, 
        N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, 
        N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, 
        N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, 
        N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, 
        N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, 
        N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, 
        N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, 
        N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, 
        N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, 
        N273, N272, N271, N270, N269, N268, N267, N266, N265, N264}), .DATA2(
        z2), .CONTROL1(N2), .CONTROL2(N263), .Z(z3) );
  GTECH_BUF B_2 ( .A(N262), .Z(N2) );
  MULT_UNS_OP mult_sub_129_aco ( .A(n), .B(N522), .Z({N780, N779, N778, N777, 
        N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, 
        N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, 
        N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, 
        N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, 
        N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, 
        N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, 
        N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, 
        N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, 
        N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, 
        N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, 
        N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, 
        N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, 
        N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, 
        N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, 
        N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, 
        N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, 
        N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, 
        N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, 
        N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, 
        N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, 
        N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525}) );
  GTECH_NOT I_0 ( .A(xregN_1), .Z(N3) );
  GTECH_BUF B_3 ( .A(xregN_1) );
  GTECH_NOT I_1 ( .A(N262), .Z(N263) );
  GTECH_BUF B_4 ( .A(N262) );
  GTECH_NOT I_2 ( .A(N522), .Z(N523) );
  GTECH_BUF B_5 ( .A(N522), .Z(N524) );
  GTECH_OR2 C811 ( .A(N524), .B(N523) );
endmodule


module modmult_N256_CC256_1 ( clk, rst, start, x, y, n, o );
  input [255:0] x;
  input [255:0] y;
  input [255:0] n;
  output [255:0] o;
  input clk, rst, start;
  wire   N0, N1, \zout[0][257] , \zout[0][256] , \zin[0][257] , \zin[0][256] ,
         \zin[0][255] , \zin[0][254] , \zin[0][253] , \zin[0][252] ,
         \zin[0][251] , \zin[0][250] , \zin[0][249] , \zin[0][248] ,
         \zin[0][247] , \zin[0][246] , \zin[0][245] , \zin[0][244] ,
         \zin[0][243] , \zin[0][242] , \zin[0][241] , \zin[0][240] ,
         \zin[0][239] , \zin[0][238] , \zin[0][237] , \zin[0][236] ,
         \zin[0][235] , \zin[0][234] , \zin[0][233] , \zin[0][232] ,
         \zin[0][231] , \zin[0][230] , \zin[0][229] , \zin[0][228] ,
         \zin[0][227] , \zin[0][226] , \zin[0][225] , \zin[0][224] ,
         \zin[0][223] , \zin[0][222] , \zin[0][221] , \zin[0][220] ,
         \zin[0][219] , \zin[0][218] , \zin[0][217] , \zin[0][216] ,
         \zin[0][215] , \zin[0][214] , \zin[0][213] , \zin[0][212] ,
         \zin[0][211] , \zin[0][210] , \zin[0][209] , \zin[0][208] ,
         \zin[0][207] , \zin[0][206] , \zin[0][205] , \zin[0][204] ,
         \zin[0][203] , \zin[0][202] , \zin[0][201] , \zin[0][200] ,
         \zin[0][199] , \zin[0][198] , \zin[0][197] , \zin[0][196] ,
         \zin[0][195] , \zin[0][194] , \zin[0][193] , \zin[0][192] ,
         \zin[0][191] , \zin[0][190] , \zin[0][189] , \zin[0][188] ,
         \zin[0][187] , \zin[0][186] , \zin[0][185] , \zin[0][184] ,
         \zin[0][183] , \zin[0][182] , \zin[0][181] , \zin[0][180] ,
         \zin[0][179] , \zin[0][178] , \zin[0][177] , \zin[0][176] ,
         \zin[0][175] , \zin[0][174] , \zin[0][173] , \zin[0][172] ,
         \zin[0][171] , \zin[0][170] , \zin[0][169] , \zin[0][168] ,
         \zin[0][167] , \zin[0][166] , \zin[0][165] , \zin[0][164] ,
         \zin[0][163] , \zin[0][162] , \zin[0][161] , \zin[0][160] ,
         \zin[0][159] , \zin[0][158] , \zin[0][157] , \zin[0][156] ,
         \zin[0][155] , \zin[0][154] , \zin[0][153] , \zin[0][152] ,
         \zin[0][151] , \zin[0][150] , \zin[0][149] , \zin[0][148] ,
         \zin[0][147] , \zin[0][146] , \zin[0][145] , \zin[0][144] ,
         \zin[0][143] , \zin[0][142] , \zin[0][141] , \zin[0][140] ,
         \zin[0][139] , \zin[0][138] , \zin[0][137] , \zin[0][136] ,
         \zin[0][135] , \zin[0][134] , \zin[0][133] , \zin[0][132] ,
         \zin[0][131] , \zin[0][130] , \zin[0][129] , \zin[0][128] ,
         \zin[0][127] , \zin[0][126] , \zin[0][125] , \zin[0][124] ,
         \zin[0][123] , \zin[0][122] , \zin[0][121] , \zin[0][120] ,
         \zin[0][119] , \zin[0][118] , \zin[0][117] , \zin[0][116] ,
         \zin[0][115] , \zin[0][114] , \zin[0][113] , \zin[0][112] ,
         \zin[0][111] , \zin[0][110] , \zin[0][109] , \zin[0][108] ,
         \zin[0][107] , \zin[0][106] , \zin[0][105] , \zin[0][104] ,
         \zin[0][103] , \zin[0][102] , \zin[0][101] , \zin[0][100] ,
         \zin[0][99] , \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] ,
         \zin[0][94] , \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] ,
         \zin[0][89] , \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] ,
         \zin[0][84] , \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] ,
         \zin[0][79] , \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] ,
         \zin[0][74] , \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] ,
         \zin[0][69] , \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] ,
         \zin[0][64] , \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] ,
         \zin[0][59] , \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] ,
         \zin[0][54] , \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] ,
         \zin[0][49] , \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] ,
         \zin[0][44] , \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] ,
         \zin[0][39] , \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] ,
         \zin[0][34] , \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] ,
         \zin[0][29] , \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] ,
         \zin[0][24] , \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] ,
         \zin[0][19] , \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] ,
         \zin[0][14] , \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] ,
         \zin[0][9] , \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] ,
         \zin[0][4] , \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] , N2;
  wire   [257:0] zreg;
  wire   [255:0] xin;
  wire   [255:0] xreg;

  modmult_step_N256_4 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[255]), 
        .y(y), .n(n), .zin({\zin[0][257] , \zin[0][256] , \zin[0][255] , 
        \zin[0][254] , \zin[0][253] , \zin[0][252] , \zin[0][251] , 
        \zin[0][250] , \zin[0][249] , \zin[0][248] , \zin[0][247] , 
        \zin[0][246] , \zin[0][245] , \zin[0][244] , \zin[0][243] , 
        \zin[0][242] , \zin[0][241] , \zin[0][240] , \zin[0][239] , 
        \zin[0][238] , \zin[0][237] , \zin[0][236] , \zin[0][235] , 
        \zin[0][234] , \zin[0][233] , \zin[0][232] , \zin[0][231] , 
        \zin[0][230] , \zin[0][229] , \zin[0][228] , \zin[0][227] , 
        \zin[0][226] , \zin[0][225] , \zin[0][224] , \zin[0][223] , 
        \zin[0][222] , \zin[0][221] , \zin[0][220] , \zin[0][219] , 
        \zin[0][218] , \zin[0][217] , \zin[0][216] , \zin[0][215] , 
        \zin[0][214] , \zin[0][213] , \zin[0][212] , \zin[0][211] , 
        \zin[0][210] , \zin[0][209] , \zin[0][208] , \zin[0][207] , 
        \zin[0][206] , \zin[0][205] , \zin[0][204] , \zin[0][203] , 
        \zin[0][202] , \zin[0][201] , \zin[0][200] , \zin[0][199] , 
        \zin[0][198] , \zin[0][197] , \zin[0][196] , \zin[0][195] , 
        \zin[0][194] , \zin[0][193] , \zin[0][192] , \zin[0][191] , 
        \zin[0][190] , \zin[0][189] , \zin[0][188] , \zin[0][187] , 
        \zin[0][186] , \zin[0][185] , \zin[0][184] , \zin[0][183] , 
        \zin[0][182] , \zin[0][181] , \zin[0][180] , \zin[0][179] , 
        \zin[0][178] , \zin[0][177] , \zin[0][176] , \zin[0][175] , 
        \zin[0][174] , \zin[0][173] , \zin[0][172] , \zin[0][171] , 
        \zin[0][170] , \zin[0][169] , \zin[0][168] , \zin[0][167] , 
        \zin[0][166] , \zin[0][165] , \zin[0][164] , \zin[0][163] , 
        \zin[0][162] , \zin[0][161] , \zin[0][160] , \zin[0][159] , 
        \zin[0][158] , \zin[0][157] , \zin[0][156] , \zin[0][155] , 
        \zin[0][154] , \zin[0][153] , \zin[0][152] , \zin[0][151] , 
        \zin[0][150] , \zin[0][149] , \zin[0][148] , \zin[0][147] , 
        \zin[0][146] , \zin[0][145] , \zin[0][144] , \zin[0][143] , 
        \zin[0][142] , \zin[0][141] , \zin[0][140] , \zin[0][139] , 
        \zin[0][138] , \zin[0][137] , \zin[0][136] , \zin[0][135] , 
        \zin[0][134] , \zin[0][133] , \zin[0][132] , \zin[0][131] , 
        \zin[0][130] , \zin[0][129] , \zin[0][128] , \zin[0][127] , 
        \zin[0][126] , \zin[0][125] , \zin[0][124] , \zin[0][123] , 
        \zin[0][122] , \zin[0][121] , \zin[0][120] , \zin[0][119] , 
        \zin[0][118] , \zin[0][117] , \zin[0][116] , \zin[0][115] , 
        \zin[0][114] , \zin[0][113] , \zin[0][112] , \zin[0][111] , 
        \zin[0][110] , \zin[0][109] , \zin[0][108] , \zin[0][107] , 
        \zin[0][106] , \zin[0][105] , \zin[0][104] , \zin[0][103] , 
        \zin[0][102] , \zin[0][101] , \zin[0][100] , \zin[0][99] , 
        \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] , 
        \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] , 
        \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] , 
        \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] , 
        \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] , 
        \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] , 
        \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] , 
        \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] , 
        \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] , 
        \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] , 
        \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] , 
        \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] , 
        \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] , 
        \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] , 
        \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] , 
        \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] , 
        \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] , 
        \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] , 
        \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] , 
        \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] }), .zout({
        \zout[0][257] , \zout[0][256] , o}) );
  \**SEQGEN**  \zreg_reg[257]  ( .clear(rst), .preset(1'b0), .next_state(
        \zout[0][257] ), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        zreg[257]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[256]  ( .clear(rst), .preset(1'b0), .next_state(
        \zout[0][256] ), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        zreg[256]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[255]  ( .clear(rst), .preset(1'b0), .next_state(
        o[255]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[255]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[254]  ( .clear(rst), .preset(1'b0), .next_state(
        o[254]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[254]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[253]  ( .clear(rst), .preset(1'b0), .next_state(
        o[253]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[253]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[252]  ( .clear(rst), .preset(1'b0), .next_state(
        o[252]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[252]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[251]  ( .clear(rst), .preset(1'b0), .next_state(
        o[251]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[251]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[250]  ( .clear(rst), .preset(1'b0), .next_state(
        o[250]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[250]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[249]  ( .clear(rst), .preset(1'b0), .next_state(
        o[249]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[249]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[248]  ( .clear(rst), .preset(1'b0), .next_state(
        o[248]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[248]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[247]  ( .clear(rst), .preset(1'b0), .next_state(
        o[247]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[247]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[246]  ( .clear(rst), .preset(1'b0), .next_state(
        o[246]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[246]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[245]  ( .clear(rst), .preset(1'b0), .next_state(
        o[245]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[245]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[244]  ( .clear(rst), .preset(1'b0), .next_state(
        o[244]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[244]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[243]  ( .clear(rst), .preset(1'b0), .next_state(
        o[243]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[243]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[242]  ( .clear(rst), .preset(1'b0), .next_state(
        o[242]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[242]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[241]  ( .clear(rst), .preset(1'b0), .next_state(
        o[241]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[241]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[240]  ( .clear(rst), .preset(1'b0), .next_state(
        o[240]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[240]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[239]  ( .clear(rst), .preset(1'b0), .next_state(
        o[239]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[239]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[238]  ( .clear(rst), .preset(1'b0), .next_state(
        o[238]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[238]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[237]  ( .clear(rst), .preset(1'b0), .next_state(
        o[237]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[237]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[236]  ( .clear(rst), .preset(1'b0), .next_state(
        o[236]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[236]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[235]  ( .clear(rst), .preset(1'b0), .next_state(
        o[235]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[235]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[234]  ( .clear(rst), .preset(1'b0), .next_state(
        o[234]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[234]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[233]  ( .clear(rst), .preset(1'b0), .next_state(
        o[233]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[233]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[232]  ( .clear(rst), .preset(1'b0), .next_state(
        o[232]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[232]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[231]  ( .clear(rst), .preset(1'b0), .next_state(
        o[231]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[231]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[230]  ( .clear(rst), .preset(1'b0), .next_state(
        o[230]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[230]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[229]  ( .clear(rst), .preset(1'b0), .next_state(
        o[229]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[229]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[228]  ( .clear(rst), .preset(1'b0), .next_state(
        o[228]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[228]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[227]  ( .clear(rst), .preset(1'b0), .next_state(
        o[227]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[227]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[226]  ( .clear(rst), .preset(1'b0), .next_state(
        o[226]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[226]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[225]  ( .clear(rst), .preset(1'b0), .next_state(
        o[225]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[225]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[224]  ( .clear(rst), .preset(1'b0), .next_state(
        o[224]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[224]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[223]  ( .clear(rst), .preset(1'b0), .next_state(
        o[223]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[223]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[222]  ( .clear(rst), .preset(1'b0), .next_state(
        o[222]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[222]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[221]  ( .clear(rst), .preset(1'b0), .next_state(
        o[221]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[221]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[220]  ( .clear(rst), .preset(1'b0), .next_state(
        o[220]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[220]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[219]  ( .clear(rst), .preset(1'b0), .next_state(
        o[219]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[219]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[218]  ( .clear(rst), .preset(1'b0), .next_state(
        o[218]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[218]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[217]  ( .clear(rst), .preset(1'b0), .next_state(
        o[217]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[217]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[216]  ( .clear(rst), .preset(1'b0), .next_state(
        o[216]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[216]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[215]  ( .clear(rst), .preset(1'b0), .next_state(
        o[215]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[215]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[214]  ( .clear(rst), .preset(1'b0), .next_state(
        o[214]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[214]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[213]  ( .clear(rst), .preset(1'b0), .next_state(
        o[213]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[213]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[212]  ( .clear(rst), .preset(1'b0), .next_state(
        o[212]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[212]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[211]  ( .clear(rst), .preset(1'b0), .next_state(
        o[211]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[211]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[210]  ( .clear(rst), .preset(1'b0), .next_state(
        o[210]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[210]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[209]  ( .clear(rst), .preset(1'b0), .next_state(
        o[209]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[209]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[208]  ( .clear(rst), .preset(1'b0), .next_state(
        o[208]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[208]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[207]  ( .clear(rst), .preset(1'b0), .next_state(
        o[207]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[207]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[206]  ( .clear(rst), .preset(1'b0), .next_state(
        o[206]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[206]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[205]  ( .clear(rst), .preset(1'b0), .next_state(
        o[205]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[205]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[204]  ( .clear(rst), .preset(1'b0), .next_state(
        o[204]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[204]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[203]  ( .clear(rst), .preset(1'b0), .next_state(
        o[203]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[203]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[202]  ( .clear(rst), .preset(1'b0), .next_state(
        o[202]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[202]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[201]  ( .clear(rst), .preset(1'b0), .next_state(
        o[201]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[201]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[200]  ( .clear(rst), .preset(1'b0), .next_state(
        o[200]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[200]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[199]  ( .clear(rst), .preset(1'b0), .next_state(
        o[199]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[199]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[198]  ( .clear(rst), .preset(1'b0), .next_state(
        o[198]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[198]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[197]  ( .clear(rst), .preset(1'b0), .next_state(
        o[197]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[197]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[196]  ( .clear(rst), .preset(1'b0), .next_state(
        o[196]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[196]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[195]  ( .clear(rst), .preset(1'b0), .next_state(
        o[195]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[195]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[194]  ( .clear(rst), .preset(1'b0), .next_state(
        o[194]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[194]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[193]  ( .clear(rst), .preset(1'b0), .next_state(
        o[193]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[193]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[192]  ( .clear(rst), .preset(1'b0), .next_state(
        o[192]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[192]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[191]  ( .clear(rst), .preset(1'b0), .next_state(
        o[191]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[191]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[190]  ( .clear(rst), .preset(1'b0), .next_state(
        o[190]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[190]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[189]  ( .clear(rst), .preset(1'b0), .next_state(
        o[189]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[189]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[188]  ( .clear(rst), .preset(1'b0), .next_state(
        o[188]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[188]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[187]  ( .clear(rst), .preset(1'b0), .next_state(
        o[187]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[187]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[186]  ( .clear(rst), .preset(1'b0), .next_state(
        o[186]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[186]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[185]  ( .clear(rst), .preset(1'b0), .next_state(
        o[185]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[185]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[184]  ( .clear(rst), .preset(1'b0), .next_state(
        o[184]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[184]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[183]  ( .clear(rst), .preset(1'b0), .next_state(
        o[183]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[183]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[182]  ( .clear(rst), .preset(1'b0), .next_state(
        o[182]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[182]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[181]  ( .clear(rst), .preset(1'b0), .next_state(
        o[181]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[181]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[180]  ( .clear(rst), .preset(1'b0), .next_state(
        o[180]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[180]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[179]  ( .clear(rst), .preset(1'b0), .next_state(
        o[179]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[179]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[178]  ( .clear(rst), .preset(1'b0), .next_state(
        o[178]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[178]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[177]  ( .clear(rst), .preset(1'b0), .next_state(
        o[177]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[177]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[176]  ( .clear(rst), .preset(1'b0), .next_state(
        o[176]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[176]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[175]  ( .clear(rst), .preset(1'b0), .next_state(
        o[175]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[175]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[174]  ( .clear(rst), .preset(1'b0), .next_state(
        o[174]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[174]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[173]  ( .clear(rst), .preset(1'b0), .next_state(
        o[173]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[173]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[172]  ( .clear(rst), .preset(1'b0), .next_state(
        o[172]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[172]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[171]  ( .clear(rst), .preset(1'b0), .next_state(
        o[171]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[171]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[170]  ( .clear(rst), .preset(1'b0), .next_state(
        o[170]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[170]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[169]  ( .clear(rst), .preset(1'b0), .next_state(
        o[169]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[169]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[168]  ( .clear(rst), .preset(1'b0), .next_state(
        o[168]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[168]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[167]  ( .clear(rst), .preset(1'b0), .next_state(
        o[167]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[167]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[166]  ( .clear(rst), .preset(1'b0), .next_state(
        o[166]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[166]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[165]  ( .clear(rst), .preset(1'b0), .next_state(
        o[165]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[165]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[164]  ( .clear(rst), .preset(1'b0), .next_state(
        o[164]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[164]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[163]  ( .clear(rst), .preset(1'b0), .next_state(
        o[163]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[163]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[162]  ( .clear(rst), .preset(1'b0), .next_state(
        o[162]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[162]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[161]  ( .clear(rst), .preset(1'b0), .next_state(
        o[161]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[161]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[160]  ( .clear(rst), .preset(1'b0), .next_state(
        o[160]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[160]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[159]  ( .clear(rst), .preset(1'b0), .next_state(
        o[159]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[159]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[158]  ( .clear(rst), .preset(1'b0), .next_state(
        o[158]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[158]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[157]  ( .clear(rst), .preset(1'b0), .next_state(
        o[157]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[157]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[156]  ( .clear(rst), .preset(1'b0), .next_state(
        o[156]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[156]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[155]  ( .clear(rst), .preset(1'b0), .next_state(
        o[155]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[155]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[154]  ( .clear(rst), .preset(1'b0), .next_state(
        o[154]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[154]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[153]  ( .clear(rst), .preset(1'b0), .next_state(
        o[153]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[153]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[152]  ( .clear(rst), .preset(1'b0), .next_state(
        o[152]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[152]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[151]  ( .clear(rst), .preset(1'b0), .next_state(
        o[151]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[151]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[150]  ( .clear(rst), .preset(1'b0), .next_state(
        o[150]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[150]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[149]  ( .clear(rst), .preset(1'b0), .next_state(
        o[149]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[149]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[148]  ( .clear(rst), .preset(1'b0), .next_state(
        o[148]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[148]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[147]  ( .clear(rst), .preset(1'b0), .next_state(
        o[147]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[147]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[146]  ( .clear(rst), .preset(1'b0), .next_state(
        o[146]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[146]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[145]  ( .clear(rst), .preset(1'b0), .next_state(
        o[145]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[145]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[144]  ( .clear(rst), .preset(1'b0), .next_state(
        o[144]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[144]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[143]  ( .clear(rst), .preset(1'b0), .next_state(
        o[143]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[143]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[142]  ( .clear(rst), .preset(1'b0), .next_state(
        o[142]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[142]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[141]  ( .clear(rst), .preset(1'b0), .next_state(
        o[141]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[141]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[140]  ( .clear(rst), .preset(1'b0), .next_state(
        o[140]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[140]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[139]  ( .clear(rst), .preset(1'b0), .next_state(
        o[139]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[139]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[138]  ( .clear(rst), .preset(1'b0), .next_state(
        o[138]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[138]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[137]  ( .clear(rst), .preset(1'b0), .next_state(
        o[137]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[137]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[136]  ( .clear(rst), .preset(1'b0), .next_state(
        o[136]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[136]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[135]  ( .clear(rst), .preset(1'b0), .next_state(
        o[135]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[135]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[134]  ( .clear(rst), .preset(1'b0), .next_state(
        o[134]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[134]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[133]  ( .clear(rst), .preset(1'b0), .next_state(
        o[133]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[133]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[132]  ( .clear(rst), .preset(1'b0), .next_state(
        o[132]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[132]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[131]  ( .clear(rst), .preset(1'b0), .next_state(
        o[131]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[131]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[130]  ( .clear(rst), .preset(1'b0), .next_state(
        o[130]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[130]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[129]  ( .clear(rst), .preset(1'b0), .next_state(
        o[129]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[129]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[128]  ( .clear(rst), .preset(1'b0), .next_state(
        o[128]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[128]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[127]  ( .clear(rst), .preset(1'b0), .next_state(
        o[127]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[127]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[126]  ( .clear(rst), .preset(1'b0), .next_state(
        o[126]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[126]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[125]  ( .clear(rst), .preset(1'b0), .next_state(
        o[125]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[125]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[124]  ( .clear(rst), .preset(1'b0), .next_state(
        o[124]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[124]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[123]  ( .clear(rst), .preset(1'b0), .next_state(
        o[123]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[123]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[122]  ( .clear(rst), .preset(1'b0), .next_state(
        o[122]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[122]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[121]  ( .clear(rst), .preset(1'b0), .next_state(
        o[121]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[121]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[120]  ( .clear(rst), .preset(1'b0), .next_state(
        o[120]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[120]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[119]  ( .clear(rst), .preset(1'b0), .next_state(
        o[119]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[119]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[118]  ( .clear(rst), .preset(1'b0), .next_state(
        o[118]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[118]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[117]  ( .clear(rst), .preset(1'b0), .next_state(
        o[117]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[117]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[116]  ( .clear(rst), .preset(1'b0), .next_state(
        o[116]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[116]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[115]  ( .clear(rst), .preset(1'b0), .next_state(
        o[115]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[115]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[114]  ( .clear(rst), .preset(1'b0), .next_state(
        o[114]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[114]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[113]  ( .clear(rst), .preset(1'b0), .next_state(
        o[113]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[113]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[112]  ( .clear(rst), .preset(1'b0), .next_state(
        o[112]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[112]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[111]  ( .clear(rst), .preset(1'b0), .next_state(
        o[111]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[111]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[110]  ( .clear(rst), .preset(1'b0), .next_state(
        o[110]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[110]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[109]  ( .clear(rst), .preset(1'b0), .next_state(
        o[109]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[109]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[108]  ( .clear(rst), .preset(1'b0), .next_state(
        o[108]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[108]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[107]  ( .clear(rst), .preset(1'b0), .next_state(
        o[107]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[107]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[106]  ( .clear(rst), .preset(1'b0), .next_state(
        o[106]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[106]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[105]  ( .clear(rst), .preset(1'b0), .next_state(
        o[105]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[105]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[104]  ( .clear(rst), .preset(1'b0), .next_state(
        o[104]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[104]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[103]  ( .clear(rst), .preset(1'b0), .next_state(
        o[103]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[103]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[102]  ( .clear(rst), .preset(1'b0), .next_state(
        o[102]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[102]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[101]  ( .clear(rst), .preset(1'b0), .next_state(
        o[101]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[101]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[100]  ( .clear(rst), .preset(1'b0), .next_state(
        o[100]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[100]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \zreg_reg[99]  ( .clear(rst), .preset(1'b0), .next_state(o[99]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[99]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[98]  ( .clear(rst), .preset(1'b0), .next_state(o[98]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[98]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[97]  ( .clear(rst), .preset(1'b0), .next_state(o[97]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[97]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[96]  ( .clear(rst), .preset(1'b0), .next_state(o[96]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[96]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[95]  ( .clear(rst), .preset(1'b0), .next_state(o[95]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[95]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[94]  ( .clear(rst), .preset(1'b0), .next_state(o[94]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[94]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[93]  ( .clear(rst), .preset(1'b0), .next_state(o[93]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[93]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[92]  ( .clear(rst), .preset(1'b0), .next_state(o[92]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[92]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[91]  ( .clear(rst), .preset(1'b0), .next_state(o[91]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[91]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[90]  ( .clear(rst), .preset(1'b0), .next_state(o[90]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[90]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[89]  ( .clear(rst), .preset(1'b0), .next_state(o[89]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[89]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[88]  ( .clear(rst), .preset(1'b0), .next_state(o[88]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[88]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[87]  ( .clear(rst), .preset(1'b0), .next_state(o[87]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[87]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[86]  ( .clear(rst), .preset(1'b0), .next_state(o[86]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[86]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[85]  ( .clear(rst), .preset(1'b0), .next_state(o[85]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[85]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[84]  ( .clear(rst), .preset(1'b0), .next_state(o[84]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[84]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[83]  ( .clear(rst), .preset(1'b0), .next_state(o[83]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[83]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[82]  ( .clear(rst), .preset(1'b0), .next_state(o[82]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[82]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[81]  ( .clear(rst), .preset(1'b0), .next_state(o[81]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[80]  ( .clear(rst), .preset(1'b0), .next_state(o[80]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[79]  ( .clear(rst), .preset(1'b0), .next_state(o[79]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[78]  ( .clear(rst), .preset(1'b0), .next_state(o[78]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[77]  ( .clear(rst), .preset(1'b0), .next_state(o[77]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[76]  ( .clear(rst), .preset(1'b0), .next_state(o[76]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[75]  ( .clear(rst), .preset(1'b0), .next_state(o[75]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[74]  ( .clear(rst), .preset(1'b0), .next_state(o[74]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[73]  ( .clear(rst), .preset(1'b0), .next_state(o[73]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[72]  ( .clear(rst), .preset(1'b0), .next_state(o[72]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[71]  ( .clear(rst), .preset(1'b0), .next_state(o[71]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[70]  ( .clear(rst), .preset(1'b0), .next_state(o[70]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[69]  ( .clear(rst), .preset(1'b0), .next_state(o[69]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[68]  ( .clear(rst), .preset(1'b0), .next_state(o[68]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[67]  ( .clear(rst), .preset(1'b0), .next_state(o[67]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[66]  ( .clear(rst), .preset(1'b0), .next_state(o[66]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[65]  ( .clear(rst), .preset(1'b0), .next_state(o[65]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[64]  ( .clear(rst), .preset(1'b0), .next_state(o[64]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[63]  ( .clear(rst), .preset(1'b0), .next_state(o[63]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[62]  ( .clear(rst), .preset(1'b0), .next_state(o[62]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[61]  ( .clear(rst), .preset(1'b0), .next_state(o[61]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[60]  ( .clear(rst), .preset(1'b0), .next_state(o[60]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[59]  ( .clear(rst), .preset(1'b0), .next_state(o[59]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[58]  ( .clear(rst), .preset(1'b0), .next_state(o[58]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[57]  ( .clear(rst), .preset(1'b0), .next_state(o[57]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[56]  ( .clear(rst), .preset(1'b0), .next_state(o[56]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[55]  ( .clear(rst), .preset(1'b0), .next_state(o[55]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[54]  ( .clear(rst), .preset(1'b0), .next_state(o[54]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[53]  ( .clear(rst), .preset(1'b0), .next_state(o[53]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[52]  ( .clear(rst), .preset(1'b0), .next_state(o[52]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[51]  ( .clear(rst), .preset(1'b0), .next_state(o[51]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[50]  ( .clear(rst), .preset(1'b0), .next_state(o[50]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[49]  ( .clear(rst), .preset(1'b0), .next_state(o[49]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[48]  ( .clear(rst), .preset(1'b0), .next_state(o[48]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[47]  ( .clear(rst), .preset(1'b0), .next_state(o[47]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[46]  ( .clear(rst), .preset(1'b0), .next_state(o[46]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[45]  ( .clear(rst), .preset(1'b0), .next_state(o[45]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[44]  ( .clear(rst), .preset(1'b0), .next_state(o[44]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[43]  ( .clear(rst), .preset(1'b0), .next_state(o[43]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[42]  ( .clear(rst), .preset(1'b0), .next_state(o[42]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[41]  ( .clear(rst), .preset(1'b0), .next_state(o[41]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[40]  ( .clear(rst), .preset(1'b0), .next_state(o[40]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[39]  ( .clear(rst), .preset(1'b0), .next_state(o[39]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[38]  ( .clear(rst), .preset(1'b0), .next_state(o[38]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[37]  ( .clear(rst), .preset(1'b0), .next_state(o[37]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[36]  ( .clear(rst), .preset(1'b0), .next_state(o[36]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[35]  ( .clear(rst), .preset(1'b0), .next_state(o[35]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[34]  ( .clear(rst), .preset(1'b0), .next_state(o[34]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[33]  ( .clear(rst), .preset(1'b0), .next_state(o[33]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[32]  ( .clear(rst), .preset(1'b0), .next_state(o[32]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[31]  ( .clear(rst), .preset(1'b0), .next_state(o[31]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[30]  ( .clear(rst), .preset(1'b0), .next_state(o[30]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[29]  ( .clear(rst), .preset(1'b0), .next_state(o[29]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[28]  ( .clear(rst), .preset(1'b0), .next_state(o[28]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[27]  ( .clear(rst), .preset(1'b0), .next_state(o[27]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[26]  ( .clear(rst), .preset(1'b0), .next_state(o[26]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[25]  ( .clear(rst), .preset(1'b0), .next_state(o[25]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[24]  ( .clear(rst), .preset(1'b0), .next_state(o[24]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[23]  ( .clear(rst), .preset(1'b0), .next_state(o[23]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[22]  ( .clear(rst), .preset(1'b0), .next_state(o[22]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[21]  ( .clear(rst), .preset(1'b0), .next_state(o[21]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[20]  ( .clear(rst), .preset(1'b0), .next_state(o[20]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[19]  ( .clear(rst), .preset(1'b0), .next_state(o[19]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[18]  ( .clear(rst), .preset(1'b0), .next_state(o[18]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[17]  ( .clear(rst), .preset(1'b0), .next_state(o[17]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[16]  ( .clear(rst), .preset(1'b0), .next_state(o[16]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[15]  ( .clear(rst), .preset(1'b0), .next_state(o[15]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[14]  ( .clear(rst), .preset(1'b0), .next_state(o[14]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[13]  ( .clear(rst), .preset(1'b0), .next_state(o[13]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[12]  ( .clear(rst), .preset(1'b0), .next_state(o[12]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[11]  ( .clear(rst), .preset(1'b0), .next_state(o[11]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[10]  ( .clear(rst), .preset(1'b0), .next_state(o[10]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[9]  ( .clear(rst), .preset(1'b0), .next_state(o[9]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[8]  ( .clear(rst), .preset(1'b0), .next_state(o[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[7]  ( .clear(rst), .preset(1'b0), .next_state(o[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[6]  ( .clear(rst), .preset(1'b0), .next_state(o[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[5]  ( .clear(rst), .preset(1'b0), .next_state(o[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[4]  ( .clear(rst), .preset(1'b0), .next_state(o[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[3]  ( .clear(rst), .preset(1'b0), .next_state(o[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[2]  ( .clear(rst), .preset(1'b0), .next_state(o[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[1]  ( .clear(rst), .preset(1'b0), .next_state(o[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \zreg_reg[0]  ( .clear(rst), .preset(1'b0), .next_state(o[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(zreg[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[255]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[254]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[255]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[254]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[253]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[254]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[253]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[252]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[253]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[252]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[251]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[252]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[251]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[250]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[251]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[250]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[249]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[250]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[249]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[248]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[249]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[248]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[247]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[248]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[247]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[246]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[247]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[246]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[245]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[246]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[245]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[244]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[245]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[244]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[243]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[244]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[243]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[242]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[243]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[242]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[241]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[242]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[241]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[240]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[241]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[240]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[239]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[240]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[239]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[238]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[239]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[238]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[237]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[238]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[237]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[236]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[237]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[236]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[235]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[236]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[235]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[234]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[235]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[234]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[233]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[234]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[233]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[232]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[233]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[232]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[231]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[232]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[231]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[230]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[231]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[230]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[229]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[230]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[229]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[228]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[229]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[228]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[227]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[228]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[227]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[226]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[227]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[226]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[225]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[226]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[225]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[224]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[225]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[224]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[223]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[224]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[223]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[222]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[223]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[222]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[221]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[222]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[221]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[220]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[221]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[220]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[219]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[220]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[219]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[218]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[219]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[218]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[217]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[218]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[217]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[216]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[217]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[216]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[215]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[216]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[215]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[214]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[215]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[214]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[213]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[214]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[213]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[212]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[213]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[212]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[211]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[212]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[211]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[210]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[211]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[210]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[209]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[210]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[209]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[208]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[209]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[208]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[207]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[208]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[207]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[206]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[207]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[206]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[205]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[206]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[205]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[204]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[205]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[204]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[203]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[204]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[203]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[202]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[203]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[202]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[201]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[202]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[201]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[200]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[201]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[200]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[199]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[200]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[199]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[198]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[199]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[198]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[197]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[198]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[197]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[196]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[197]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[196]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[195]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[196]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[195]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[194]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[195]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[194]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[193]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[194]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[193]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[192]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[193]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[192]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[191]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[192]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[191]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[190]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[191]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[190]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[189]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[190]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[189]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[188]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[189]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[188]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[187]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[188]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[187]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[186]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[187]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[186]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[185]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[186]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[185]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[184]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[185]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[184]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[183]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[184]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[183]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[182]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[183]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[182]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[181]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[182]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[181]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[180]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[181]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[180]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[179]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[180]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[179]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[178]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[179]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[178]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[177]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[178]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[177]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[176]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[177]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[176]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[175]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[176]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[175]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[174]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[175]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[174]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[173]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[174]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[173]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[172]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[173]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[172]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[171]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[172]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[171]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[170]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[171]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[170]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[169]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[170]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[169]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[168]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[169]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[168]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[167]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[168]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[167]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[166]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[167]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[166]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[165]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[166]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[165]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[164]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[165]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[164]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[163]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[164]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[163]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[162]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[163]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[162]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[161]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[162]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[161]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[160]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[161]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[160]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[159]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[160]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[159]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[158]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[159]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[158]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[157]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[158]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[157]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[156]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[157]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[156]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[155]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[156]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[155]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[154]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[155]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[154]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[153]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[154]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[153]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[152]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[153]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[152]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[151]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[152]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[151]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[150]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[151]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[150]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[149]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[150]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[149]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[148]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[149]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[148]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[147]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[148]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[147]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[146]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[147]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[146]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[145]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[146]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[145]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[144]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[145]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[144]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[143]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[144]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[143]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[142]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[143]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[142]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[141]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[142]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[141]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[140]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[141]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[140]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[139]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[140]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[139]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[138]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[139]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[138]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[137]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[138]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[137]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[136]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[137]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[136]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[135]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[136]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[135]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[134]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[135]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[134]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[133]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[134]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[133]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[132]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[133]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[132]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[131]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[132]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[131]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[130]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[131]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[130]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[129]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[130]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[129]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[128]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[129]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[128]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[127]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[128]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[127]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[126]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[127]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[126]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[125]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[126]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[125]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[124]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[125]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[124]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[123]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[124]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[123]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[122]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[123]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[122]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[121]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[122]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[121]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[120]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[121]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[120]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[119]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[120]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[119]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[118]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[119]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[118]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[117]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[118]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[117]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[116]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[117]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[116]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[115]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[116]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[115]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[114]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[115]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[114]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[113]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[114]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[113]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[112]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[113]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[112]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[111]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[112]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[111]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[110]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[111]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[110]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[109]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[110]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[109]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[108]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[109]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[108]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[107]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[108]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[107]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[106]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[107]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[106]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[105]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[106]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[105]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[104]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[105]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[104]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[103]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[104]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[103]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[102]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[103]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[102]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[101]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[102]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[101]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[100]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[101]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[100]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[99]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        xreg[100]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[99]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[98]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[99]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[98]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[97]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[98]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[97]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[96]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[97]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[96]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[95]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[96]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[95]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[94]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[95]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[94]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[93]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[94]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[93]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[92]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[93]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[92]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[91]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[92]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[91]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[90]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[91]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[90]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[89]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[90]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[89]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[88]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[89]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[88]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[87]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[88]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[87]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[86]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[87]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[86]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[85]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[86]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[85]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[84]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[85]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[84]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[83]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[84]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[83]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[82]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[83]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[82]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[81]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[82]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[81]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[80]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[81]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[80]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[79]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[80]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[79]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[78]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[79]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[78]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[77]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[78]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[77]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[76]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[77]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[76]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[75]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[76]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[75]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[74]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[75]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[74]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[73]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[74]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[73]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[72]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[73]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[72]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[71]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[72]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[71]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[70]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[71]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[70]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[69]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[70]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[69]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[68]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[69]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[68]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[67]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[68]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[67]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[66]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[67]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[66]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[65]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[66]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[65]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[64]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[65]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[64]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[63]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[64]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[63]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[62]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[63]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[62]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[61]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[62]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[61]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[60]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[61]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[60]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[59]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[60]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[59]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[58]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[59]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[58]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[57]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[58]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[57]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[56]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[57]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[56]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[55]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[56]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[55]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[54]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[55]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[54]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[53]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[54]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[53]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[52]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[53]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[52]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[51]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[52]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[51]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[50]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[51]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[50]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[49]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[50]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[49]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[48]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[49]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[48]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[47]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[48]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[47]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[46]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[47]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[46]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[45]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[46]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[45]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[44]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[45]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[44]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[43]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[44]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[43]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[42]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[43]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[42]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[42]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[41]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[41]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[40]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[40]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[39]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[39]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[38]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[38]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[37]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[37]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[36]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[36]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[35]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[35]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[34]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[34]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[33]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[33]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[32]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[32]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[31]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[30]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[29]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[28]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[27]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[26]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[25]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[24]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[23]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[22]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[21]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[20]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[19]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[18]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[17]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[16]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[15]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[14]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[13]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[12]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[11]  ( .clear(rst), .preset(1'b0), .next_state(
        xin[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(
        1'b1) );
  \**SEQGEN**  \xreg_reg[10]  ( .clear(rst), .preset(1'b0), .next_state(xin[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[10]), .synch_clear(
        1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), .synch_enable(1'b1)
         );
  \**SEQGEN**  \xreg_reg[9]  ( .clear(rst), .preset(1'b0), .next_state(xin[8]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[8]  ( .clear(rst), .preset(1'b0), .next_state(xin[7]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[7]  ( .clear(rst), .preset(1'b0), .next_state(xin[6]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[6]  ( .clear(rst), .preset(1'b0), .next_state(xin[5]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[5]  ( .clear(rst), .preset(1'b0), .next_state(xin[4]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[4]  ( .clear(rst), .preset(1'b0), .next_state(xin[3]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[3]  ( .clear(rst), .preset(1'b0), .next_state(xin[2]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[2]  ( .clear(rst), .preset(1'b0), .next_state(xin[1]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[1]  ( .clear(rst), .preset(1'b0), .next_state(xin[0]), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \xreg_reg[0]  ( .clear(rst), .preset(1'b0), .next_state(1'b0), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(xreg[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  SELECT_OP C1562 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .DATA2(
        zreg), .CONTROL1(N0), .CONTROL2(N1), .Z({\zin[0][257] , \zin[0][256] , 
        \zin[0][255] , \zin[0][254] , \zin[0][253] , \zin[0][252] , 
        \zin[0][251] , \zin[0][250] , \zin[0][249] , \zin[0][248] , 
        \zin[0][247] , \zin[0][246] , \zin[0][245] , \zin[0][244] , 
        \zin[0][243] , \zin[0][242] , \zin[0][241] , \zin[0][240] , 
        \zin[0][239] , \zin[0][238] , \zin[0][237] , \zin[0][236] , 
        \zin[0][235] , \zin[0][234] , \zin[0][233] , \zin[0][232] , 
        \zin[0][231] , \zin[0][230] , \zin[0][229] , \zin[0][228] , 
        \zin[0][227] , \zin[0][226] , \zin[0][225] , \zin[0][224] , 
        \zin[0][223] , \zin[0][222] , \zin[0][221] , \zin[0][220] , 
        \zin[0][219] , \zin[0][218] , \zin[0][217] , \zin[0][216] , 
        \zin[0][215] , \zin[0][214] , \zin[0][213] , \zin[0][212] , 
        \zin[0][211] , \zin[0][210] , \zin[0][209] , \zin[0][208] , 
        \zin[0][207] , \zin[0][206] , \zin[0][205] , \zin[0][204] , 
        \zin[0][203] , \zin[0][202] , \zin[0][201] , \zin[0][200] , 
        \zin[0][199] , \zin[0][198] , \zin[0][197] , \zin[0][196] , 
        \zin[0][195] , \zin[0][194] , \zin[0][193] , \zin[0][192] , 
        \zin[0][191] , \zin[0][190] , \zin[0][189] , \zin[0][188] , 
        \zin[0][187] , \zin[0][186] , \zin[0][185] , \zin[0][184] , 
        \zin[0][183] , \zin[0][182] , \zin[0][181] , \zin[0][180] , 
        \zin[0][179] , \zin[0][178] , \zin[0][177] , \zin[0][176] , 
        \zin[0][175] , \zin[0][174] , \zin[0][173] , \zin[0][172] , 
        \zin[0][171] , \zin[0][170] , \zin[0][169] , \zin[0][168] , 
        \zin[0][167] , \zin[0][166] , \zin[0][165] , \zin[0][164] , 
        \zin[0][163] , \zin[0][162] , \zin[0][161] , \zin[0][160] , 
        \zin[0][159] , \zin[0][158] , \zin[0][157] , \zin[0][156] , 
        \zin[0][155] , \zin[0][154] , \zin[0][153] , \zin[0][152] , 
        \zin[0][151] , \zin[0][150] , \zin[0][149] , \zin[0][148] , 
        \zin[0][147] , \zin[0][146] , \zin[0][145] , \zin[0][144] , 
        \zin[0][143] , \zin[0][142] , \zin[0][141] , \zin[0][140] , 
        \zin[0][139] , \zin[0][138] , \zin[0][137] , \zin[0][136] , 
        \zin[0][135] , \zin[0][134] , \zin[0][133] , \zin[0][132] , 
        \zin[0][131] , \zin[0][130] , \zin[0][129] , \zin[0][128] , 
        \zin[0][127] , \zin[0][126] , \zin[0][125] , \zin[0][124] , 
        \zin[0][123] , \zin[0][122] , \zin[0][121] , \zin[0][120] , 
        \zin[0][119] , \zin[0][118] , \zin[0][117] , \zin[0][116] , 
        \zin[0][115] , \zin[0][114] , \zin[0][113] , \zin[0][112] , 
        \zin[0][111] , \zin[0][110] , \zin[0][109] , \zin[0][108] , 
        \zin[0][107] , \zin[0][106] , \zin[0][105] , \zin[0][104] , 
        \zin[0][103] , \zin[0][102] , \zin[0][101] , \zin[0][100] , 
        \zin[0][99] , \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] , 
        \zin[0][94] , \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] , 
        \zin[0][89] , \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] , 
        \zin[0][84] , \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] , 
        \zin[0][79] , \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] , 
        \zin[0][74] , \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] , 
        \zin[0][69] , \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] , 
        \zin[0][64] , \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] , 
        \zin[0][59] , \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] , 
        \zin[0][54] , \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] , 
        \zin[0][49] , \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] , 
        \zin[0][44] , \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] , 
        \zin[0][39] , \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] , 
        \zin[0][34] , \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] , 
        \zin[0][29] , \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] , 
        \zin[0][24] , \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] , 
        \zin[0][19] , \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] , 
        \zin[0][14] , \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] , 
        \zin[0][9] , \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] , 
        \zin[0][4] , \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] }) );
  GTECH_BUF B_0 ( .A(start), .Z(N0) );
  GTECH_BUF B_1 ( .A(N2), .Z(N1) );
  SELECT_OP C1563 ( .DATA1(x), .DATA2(xreg), .CONTROL1(N0), .CONTROL2(N1), .Z(
        xin) );
  GTECH_NOT I_0 ( .A(start), .Z(N2) );
endmodule


module modexp_2N_NN_N256_CC131072 ( clk, rst, m, e, n, c );
  input [255:0] m;
  input [255:0] e;
  input [255:0] n;
  output [255:0] c;
  input clk, rst;
  wire   N0, N1, N2, N3, N4, init, N5, N6, mul_pow, N7, first_one, N8, N9, N10,
         N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370,
         N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458,
         N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491,
         N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502,
         N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540;
  wire   [255:0] start_in;
  wire   [255:0] start_reg;
  wire   [255:0] ein;
  wire   [255:0] ereg;
  wire   [255:0] o;
  wire   [255:0] creg;
  wire   [255:0] x;
  wire   [255:0] y;

  \**SEQGEN**  first_one_reg ( .clear(rst), .preset(1'b0), .next_state(1'b1), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(first_one), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N532) );
  \**SEQGEN**  init_reg ( .clear(rst), .preset(1'b0), .next_state(1'b1), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(init), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(1'b1) );
  \**SEQGEN**  \ereg_reg[255]  ( .clear(rst), .preset(1'b0), .next_state(N272), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[255]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[254]  ( .clear(rst), .preset(1'b0), .next_state(N271), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[254]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[253]  ( .clear(rst), .preset(1'b0), .next_state(N270), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[253]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[252]  ( .clear(rst), .preset(1'b0), .next_state(N269), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[252]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[251]  ( .clear(rst), .preset(1'b0), .next_state(N268), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[251]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[250]  ( .clear(rst), .preset(1'b0), .next_state(N267), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[250]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[249]  ( .clear(rst), .preset(1'b0), .next_state(N266), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[249]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[248]  ( .clear(rst), .preset(1'b0), .next_state(N265), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[248]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[247]  ( .clear(rst), .preset(1'b0), .next_state(N264), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[247]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[246]  ( .clear(rst), .preset(1'b0), .next_state(N263), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[246]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[245]  ( .clear(rst), .preset(1'b0), .next_state(N262), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[245]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[244]  ( .clear(rst), .preset(1'b0), .next_state(N261), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[244]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[243]  ( .clear(rst), .preset(1'b0), .next_state(N260), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[243]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[242]  ( .clear(rst), .preset(1'b0), .next_state(N259), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[242]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[241]  ( .clear(rst), .preset(1'b0), .next_state(N258), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[241]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[240]  ( .clear(rst), .preset(1'b0), .next_state(N257), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[240]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[239]  ( .clear(rst), .preset(1'b0), .next_state(N256), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[239]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[238]  ( .clear(rst), .preset(1'b0), .next_state(N255), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[238]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[237]  ( .clear(rst), .preset(1'b0), .next_state(N254), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[237]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[236]  ( .clear(rst), .preset(1'b0), .next_state(N253), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[236]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[235]  ( .clear(rst), .preset(1'b0), .next_state(N252), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[235]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[234]  ( .clear(rst), .preset(1'b0), .next_state(N251), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[234]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[233]  ( .clear(rst), .preset(1'b0), .next_state(N250), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[233]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[232]  ( .clear(rst), .preset(1'b0), .next_state(N249), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[232]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[231]  ( .clear(rst), .preset(1'b0), .next_state(N248), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[231]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[230]  ( .clear(rst), .preset(1'b0), .next_state(N247), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[230]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[229]  ( .clear(rst), .preset(1'b0), .next_state(N246), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[229]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[228]  ( .clear(rst), .preset(1'b0), .next_state(N245), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[228]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[227]  ( .clear(rst), .preset(1'b0), .next_state(N244), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[227]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[226]  ( .clear(rst), .preset(1'b0), .next_state(N243), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[226]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[225]  ( .clear(rst), .preset(1'b0), .next_state(N242), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[225]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[224]  ( .clear(rst), .preset(1'b0), .next_state(N241), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[224]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[223]  ( .clear(rst), .preset(1'b0), .next_state(N240), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[223]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[222]  ( .clear(rst), .preset(1'b0), .next_state(N239), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[222]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[221]  ( .clear(rst), .preset(1'b0), .next_state(N238), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[221]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[220]  ( .clear(rst), .preset(1'b0), .next_state(N237), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[220]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[219]  ( .clear(rst), .preset(1'b0), .next_state(N236), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[219]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[218]  ( .clear(rst), .preset(1'b0), .next_state(N235), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[218]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[217]  ( .clear(rst), .preset(1'b0), .next_state(N234), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[217]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[216]  ( .clear(rst), .preset(1'b0), .next_state(N233), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[216]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[215]  ( .clear(rst), .preset(1'b0), .next_state(N232), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[215]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[214]  ( .clear(rst), .preset(1'b0), .next_state(N231), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[214]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[213]  ( .clear(rst), .preset(1'b0), .next_state(N230), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[213]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[212]  ( .clear(rst), .preset(1'b0), .next_state(N229), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[212]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[211]  ( .clear(rst), .preset(1'b0), .next_state(N228), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[211]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[210]  ( .clear(rst), .preset(1'b0), .next_state(N227), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[210]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[209]  ( .clear(rst), .preset(1'b0), .next_state(N226), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[209]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[208]  ( .clear(rst), .preset(1'b0), .next_state(N225), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[208]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[207]  ( .clear(rst), .preset(1'b0), .next_state(N224), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[207]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[206]  ( .clear(rst), .preset(1'b0), .next_state(N223), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[206]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[205]  ( .clear(rst), .preset(1'b0), .next_state(N222), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[205]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[204]  ( .clear(rst), .preset(1'b0), .next_state(N221), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[204]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[203]  ( .clear(rst), .preset(1'b0), .next_state(N220), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[203]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[202]  ( .clear(rst), .preset(1'b0), .next_state(N219), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[202]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[201]  ( .clear(rst), .preset(1'b0), .next_state(N218), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[201]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[200]  ( .clear(rst), .preset(1'b0), .next_state(N217), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[200]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[199]  ( .clear(rst), .preset(1'b0), .next_state(N216), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[199]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[198]  ( .clear(rst), .preset(1'b0), .next_state(N215), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[198]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N214) );
  \**SEQGEN**  \ereg_reg[197]  ( .clear(rst), .preset(1'b0), .next_state(N213), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[197]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[196]  ( .clear(rst), .preset(1'b0), .next_state(N212), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[196]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[195]  ( .clear(rst), .preset(1'b0), .next_state(N211), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[195]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[194]  ( .clear(rst), .preset(1'b0), .next_state(N210), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[194]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[193]  ( .clear(rst), .preset(1'b0), .next_state(N209), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[193]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[192]  ( .clear(rst), .preset(1'b0), .next_state(N208), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[192]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[191]  ( .clear(rst), .preset(1'b0), .next_state(N207), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[191]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[190]  ( .clear(rst), .preset(1'b0), .next_state(N206), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[190]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[189]  ( .clear(rst), .preset(1'b0), .next_state(N205), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[189]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[188]  ( .clear(rst), .preset(1'b0), .next_state(N204), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[188]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[187]  ( .clear(rst), .preset(1'b0), .next_state(N203), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[187]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[186]  ( .clear(rst), .preset(1'b0), .next_state(N202), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[186]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[185]  ( .clear(rst), .preset(1'b0), .next_state(N201), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[185]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[184]  ( .clear(rst), .preset(1'b0), .next_state(N200), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[184]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[183]  ( .clear(rst), .preset(1'b0), .next_state(N199), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[183]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[182]  ( .clear(rst), .preset(1'b0), .next_state(N198), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[182]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[181]  ( .clear(rst), .preset(1'b0), .next_state(N197), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[181]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[180]  ( .clear(rst), .preset(1'b0), .next_state(N196), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[180]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[179]  ( .clear(rst), .preset(1'b0), .next_state(N195), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[179]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[178]  ( .clear(rst), .preset(1'b0), .next_state(N194), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[178]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[177]  ( .clear(rst), .preset(1'b0), .next_state(N193), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[177]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[176]  ( .clear(rst), .preset(1'b0), .next_state(N192), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[176]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[175]  ( .clear(rst), .preset(1'b0), .next_state(N191), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[175]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[174]  ( .clear(rst), .preset(1'b0), .next_state(N190), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[174]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[173]  ( .clear(rst), .preset(1'b0), .next_state(N189), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[173]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[172]  ( .clear(rst), .preset(1'b0), .next_state(N188), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[172]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[171]  ( .clear(rst), .preset(1'b0), .next_state(N187), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[171]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[170]  ( .clear(rst), .preset(1'b0), .next_state(N186), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[170]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[169]  ( .clear(rst), .preset(1'b0), .next_state(N185), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[169]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[168]  ( .clear(rst), .preset(1'b0), .next_state(N184), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[168]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[167]  ( .clear(rst), .preset(1'b0), .next_state(N183), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[167]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[166]  ( .clear(rst), .preset(1'b0), .next_state(N182), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[166]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[165]  ( .clear(rst), .preset(1'b0), .next_state(N181), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[165]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[164]  ( .clear(rst), .preset(1'b0), .next_state(N180), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[164]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[163]  ( .clear(rst), .preset(1'b0), .next_state(N179), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[163]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[162]  ( .clear(rst), .preset(1'b0), .next_state(N178), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[162]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[161]  ( .clear(rst), .preset(1'b0), .next_state(N177), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[161]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[160]  ( .clear(rst), .preset(1'b0), .next_state(N176), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[160]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[159]  ( .clear(rst), .preset(1'b0), .next_state(N175), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[159]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[158]  ( .clear(rst), .preset(1'b0), .next_state(N174), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[158]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[157]  ( .clear(rst), .preset(1'b0), .next_state(N173), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[157]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[156]  ( .clear(rst), .preset(1'b0), .next_state(N172), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[156]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[155]  ( .clear(rst), .preset(1'b0), .next_state(N171), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[155]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[154]  ( .clear(rst), .preset(1'b0), .next_state(N170), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[154]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[153]  ( .clear(rst), .preset(1'b0), .next_state(N169), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[153]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[152]  ( .clear(rst), .preset(1'b0), .next_state(N168), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[152]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[151]  ( .clear(rst), .preset(1'b0), .next_state(N167), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[151]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[150]  ( .clear(rst), .preset(1'b0), .next_state(N166), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[150]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[149]  ( .clear(rst), .preset(1'b0), .next_state(N165), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[149]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[148]  ( .clear(rst), .preset(1'b0), .next_state(N164), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[148]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[147]  ( .clear(rst), .preset(1'b0), .next_state(N163), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[147]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[146]  ( .clear(rst), .preset(1'b0), .next_state(N162), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[146]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[145]  ( .clear(rst), .preset(1'b0), .next_state(N161), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[145]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[144]  ( .clear(rst), .preset(1'b0), .next_state(N160), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[144]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[143]  ( .clear(rst), .preset(1'b0), .next_state(N159), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[143]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[142]  ( .clear(rst), .preset(1'b0), .next_state(N158), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[142]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[141]  ( .clear(rst), .preset(1'b0), .next_state(N157), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[141]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[140]  ( .clear(rst), .preset(1'b0), .next_state(N156), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[140]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[139]  ( .clear(rst), .preset(1'b0), .next_state(N155), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[139]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[138]  ( .clear(rst), .preset(1'b0), .next_state(N154), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[138]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[137]  ( .clear(rst), .preset(1'b0), .next_state(N153), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[137]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[136]  ( .clear(rst), .preset(1'b0), .next_state(N152), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[136]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[135]  ( .clear(rst), .preset(1'b0), .next_state(N151), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[135]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[134]  ( .clear(rst), .preset(1'b0), .next_state(N150), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[134]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[133]  ( .clear(rst), .preset(1'b0), .next_state(N149), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[133]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[132]  ( .clear(rst), .preset(1'b0), .next_state(N148), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[132]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[131]  ( .clear(rst), .preset(1'b0), .next_state(N147), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[131]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[130]  ( .clear(rst), .preset(1'b0), .next_state(N146), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[130]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[129]  ( .clear(rst), .preset(1'b0), .next_state(N145), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[129]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[128]  ( .clear(rst), .preset(1'b0), .next_state(N144), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[128]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[127]  ( .clear(rst), .preset(1'b0), .next_state(N143), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[127]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[126]  ( .clear(rst), .preset(1'b0), .next_state(N142), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[126]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[125]  ( .clear(rst), .preset(1'b0), .next_state(N141), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[125]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[124]  ( .clear(rst), .preset(1'b0), .next_state(N140), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[124]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[123]  ( .clear(rst), .preset(1'b0), .next_state(N139), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[123]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[122]  ( .clear(rst), .preset(1'b0), .next_state(N138), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[122]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[121]  ( .clear(rst), .preset(1'b0), .next_state(N137), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[121]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[120]  ( .clear(rst), .preset(1'b0), .next_state(N136), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[120]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[119]  ( .clear(rst), .preset(1'b0), .next_state(N135), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[119]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[118]  ( .clear(rst), .preset(1'b0), .next_state(N134), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[118]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[117]  ( .clear(rst), .preset(1'b0), .next_state(N133), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[117]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[116]  ( .clear(rst), .preset(1'b0), .next_state(N132), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[116]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[115]  ( .clear(rst), .preset(1'b0), .next_state(N131), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[115]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[114]  ( .clear(rst), .preset(1'b0), .next_state(N130), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[114]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[113]  ( .clear(rst), .preset(1'b0), .next_state(N129), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[113]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[112]  ( .clear(rst), .preset(1'b0), .next_state(N128), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[112]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[111]  ( .clear(rst), .preset(1'b0), .next_state(N127), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[111]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[110]  ( .clear(rst), .preset(1'b0), .next_state(N126), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[110]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[109]  ( .clear(rst), .preset(1'b0), .next_state(N125), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[109]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[108]  ( .clear(rst), .preset(1'b0), .next_state(N124), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[108]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[107]  ( .clear(rst), .preset(1'b0), .next_state(N123), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[107]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[106]  ( .clear(rst), .preset(1'b0), .next_state(N122), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[106]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[105]  ( .clear(rst), .preset(1'b0), .next_state(N121), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[105]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[104]  ( .clear(rst), .preset(1'b0), .next_state(N120), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[104]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[103]  ( .clear(rst), .preset(1'b0), .next_state(N119), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[103]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[102]  ( .clear(rst), .preset(1'b0), .next_state(N118), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[102]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[101]  ( .clear(rst), .preset(1'b0), .next_state(N117), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[101]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[100]  ( .clear(rst), .preset(1'b0), .next_state(N116), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[100]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[99]  ( .clear(rst), .preset(1'b0), .next_state(N115), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[99]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N114) );
  \**SEQGEN**  \ereg_reg[98]  ( .clear(rst), .preset(1'b0), .next_state(N113), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[98]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[97]  ( .clear(rst), .preset(1'b0), .next_state(N112), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[97]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[96]  ( .clear(rst), .preset(1'b0), .next_state(N111), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[96]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[95]  ( .clear(rst), .preset(1'b0), .next_state(N110), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[95]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[94]  ( .clear(rst), .preset(1'b0), .next_state(N109), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[94]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[93]  ( .clear(rst), .preset(1'b0), .next_state(N108), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[93]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[92]  ( .clear(rst), .preset(1'b0), .next_state(N107), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[92]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[91]  ( .clear(rst), .preset(1'b0), .next_state(N106), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[91]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[90]  ( .clear(rst), .preset(1'b0), .next_state(N105), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[90]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[89]  ( .clear(rst), .preset(1'b0), .next_state(N104), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[89]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[88]  ( .clear(rst), .preset(1'b0), .next_state(N103), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[88]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[87]  ( .clear(rst), .preset(1'b0), .next_state(N102), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[87]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[86]  ( .clear(rst), .preset(1'b0), .next_state(N101), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[86]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[85]  ( .clear(rst), .preset(1'b0), .next_state(N100), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[85]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[84]  ( .clear(rst), .preset(1'b0), .next_state(N99), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[84]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[83]  ( .clear(rst), .preset(1'b0), .next_state(N98), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[83]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[82]  ( .clear(rst), .preset(1'b0), .next_state(N97), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[82]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[81]  ( .clear(rst), .preset(1'b0), .next_state(N96), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[80]  ( .clear(rst), .preset(1'b0), .next_state(N95), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[79]  ( .clear(rst), .preset(1'b0), .next_state(N94), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[78]  ( .clear(rst), .preset(1'b0), .next_state(N93), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[77]  ( .clear(rst), .preset(1'b0), .next_state(N92), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[76]  ( .clear(rst), .preset(1'b0), .next_state(N91), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[75]  ( .clear(rst), .preset(1'b0), .next_state(N90), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[74]  ( .clear(rst), .preset(1'b0), .next_state(N89), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[73]  ( .clear(rst), .preset(1'b0), .next_state(N88), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[72]  ( .clear(rst), .preset(1'b0), .next_state(N87), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[71]  ( .clear(rst), .preset(1'b0), .next_state(N86), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[70]  ( .clear(rst), .preset(1'b0), .next_state(N85), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[69]  ( .clear(rst), .preset(1'b0), .next_state(N84), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[68]  ( .clear(rst), .preset(1'b0), .next_state(N83), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[67]  ( .clear(rst), .preset(1'b0), .next_state(N82), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[66]  ( .clear(rst), .preset(1'b0), .next_state(N81), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[65]  ( .clear(rst), .preset(1'b0), .next_state(N80), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[64]  ( .clear(rst), .preset(1'b0), .next_state(N79), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[63]  ( .clear(rst), .preset(1'b0), .next_state(N78), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[62]  ( .clear(rst), .preset(1'b0), .next_state(N77), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[61]  ( .clear(rst), .preset(1'b0), .next_state(N76), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[60]  ( .clear(rst), .preset(1'b0), .next_state(N75), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[59]  ( .clear(rst), .preset(1'b0), .next_state(N74), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[58]  ( .clear(rst), .preset(1'b0), .next_state(N73), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[57]  ( .clear(rst), .preset(1'b0), .next_state(N72), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[56]  ( .clear(rst), .preset(1'b0), .next_state(N71), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[55]  ( .clear(rst), .preset(1'b0), .next_state(N70), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[54]  ( .clear(rst), .preset(1'b0), .next_state(N69), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[53]  ( .clear(rst), .preset(1'b0), .next_state(N68), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[52]  ( .clear(rst), .preset(1'b0), .next_state(N67), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[51]  ( .clear(rst), .preset(1'b0), .next_state(N66), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[50]  ( .clear(rst), .preset(1'b0), .next_state(N65), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[49]  ( .clear(rst), .preset(1'b0), .next_state(N64), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[48]  ( .clear(rst), .preset(1'b0), .next_state(N63), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[47]  ( .clear(rst), .preset(1'b0), .next_state(N62), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[46]  ( .clear(rst), .preset(1'b0), .next_state(N61), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[45]  ( .clear(rst), .preset(1'b0), .next_state(N60), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[44]  ( .clear(rst), .preset(1'b0), .next_state(N59), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[43]  ( .clear(rst), .preset(1'b0), .next_state(N58), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[42]  ( .clear(rst), .preset(1'b0), .next_state(N57), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[41]  ( .clear(rst), .preset(1'b0), .next_state(N56), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[40]  ( .clear(rst), .preset(1'b0), .next_state(N55), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[39]  ( .clear(rst), .preset(1'b0), .next_state(N54), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[38]  ( .clear(rst), .preset(1'b0), .next_state(N53), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[37]  ( .clear(rst), .preset(1'b0), .next_state(N52), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[36]  ( .clear(rst), .preset(1'b0), .next_state(N51), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[35]  ( .clear(rst), .preset(1'b0), .next_state(N50), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[34]  ( .clear(rst), .preset(1'b0), .next_state(N49), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[33]  ( .clear(rst), .preset(1'b0), .next_state(N48), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[32]  ( .clear(rst), .preset(1'b0), .next_state(N47), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[31]  ( .clear(rst), .preset(1'b0), .next_state(N46), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[30]  ( .clear(rst), .preset(1'b0), .next_state(N45), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[29]  ( .clear(rst), .preset(1'b0), .next_state(N44), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[28]  ( .clear(rst), .preset(1'b0), .next_state(N43), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[27]  ( .clear(rst), .preset(1'b0), .next_state(N42), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[26]  ( .clear(rst), .preset(1'b0), .next_state(N41), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[25]  ( .clear(rst), .preset(1'b0), .next_state(N40), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[24]  ( .clear(rst), .preset(1'b0), .next_state(N39), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[23]  ( .clear(rst), .preset(1'b0), .next_state(N38), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[22]  ( .clear(rst), .preset(1'b0), .next_state(N37), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[21]  ( .clear(rst), .preset(1'b0), .next_state(N36), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[20]  ( .clear(rst), .preset(1'b0), .next_state(N35), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[19]  ( .clear(rst), .preset(1'b0), .next_state(N34), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[18]  ( .clear(rst), .preset(1'b0), .next_state(N33), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[17]  ( .clear(rst), .preset(1'b0), .next_state(N32), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[16]  ( .clear(rst), .preset(1'b0), .next_state(N31), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[15]  ( .clear(rst), .preset(1'b0), .next_state(N30), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[14]  ( .clear(rst), .preset(1'b0), .next_state(N29), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[13]  ( .clear(rst), .preset(1'b0), .next_state(N28), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[12]  ( .clear(rst), .preset(1'b0), .next_state(N27), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[11]  ( .clear(rst), .preset(1'b0), .next_state(N26), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[10]  ( .clear(rst), .preset(1'b0), .next_state(N25), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[9]  ( .clear(rst), .preset(1'b0), .next_state(N24), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[8]  ( .clear(rst), .preset(1'b0), .next_state(N23), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[7]  ( .clear(rst), .preset(1'b0), .next_state(N22), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[6]  ( .clear(rst), .preset(1'b0), .next_state(N21), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[5]  ( .clear(rst), .preset(1'b0), .next_state(N20), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[4]  ( .clear(rst), .preset(1'b0), .next_state(N19), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[3]  ( .clear(rst), .preset(1'b0), .next_state(N18), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[2]  ( .clear(rst), .preset(1'b0), .next_state(N17), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[1]  ( .clear(rst), .preset(1'b0), .next_state(N16), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  \ereg_reg[0]  ( .clear(rst), .preset(1'b0), .next_state(N15), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(ereg[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N14) );
  \**SEQGEN**  mul_pow_reg ( .clear(rst), .preset(1'b0), .next_state(N7), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(mul_pow), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(start_in[255]) );
  \**SEQGEN**  \creg_reg[255]  ( .clear(rst), .preset(1'b0), .next_state(N531), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[255]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[254]  ( .clear(rst), .preset(1'b0), .next_state(N530), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[254]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[253]  ( .clear(rst), .preset(1'b0), .next_state(N529), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[253]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[252]  ( .clear(rst), .preset(1'b0), .next_state(N528), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[252]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[251]  ( .clear(rst), .preset(1'b0), .next_state(N527), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[251]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[250]  ( .clear(rst), .preset(1'b0), .next_state(N526), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[250]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[249]  ( .clear(rst), .preset(1'b0), .next_state(N525), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[249]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[248]  ( .clear(rst), .preset(1'b0), .next_state(N524), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[248]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[247]  ( .clear(rst), .preset(1'b0), .next_state(N523), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[247]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[246]  ( .clear(rst), .preset(1'b0), .next_state(N522), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[246]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[245]  ( .clear(rst), .preset(1'b0), .next_state(N521), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[245]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[244]  ( .clear(rst), .preset(1'b0), .next_state(N520), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[244]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[243]  ( .clear(rst), .preset(1'b0), .next_state(N519), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[243]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[242]  ( .clear(rst), .preset(1'b0), .next_state(N518), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[242]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[241]  ( .clear(rst), .preset(1'b0), .next_state(N517), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[241]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[240]  ( .clear(rst), .preset(1'b0), .next_state(N516), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[240]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[239]  ( .clear(rst), .preset(1'b0), .next_state(N515), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[239]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[238]  ( .clear(rst), .preset(1'b0), .next_state(N514), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[238]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[237]  ( .clear(rst), .preset(1'b0), .next_state(N513), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[237]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[236]  ( .clear(rst), .preset(1'b0), .next_state(N512), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[236]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[235]  ( .clear(rst), .preset(1'b0), .next_state(N511), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[235]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[234]  ( .clear(rst), .preset(1'b0), .next_state(N510), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[234]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[233]  ( .clear(rst), .preset(1'b0), .next_state(N509), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[233]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[232]  ( .clear(rst), .preset(1'b0), .next_state(N508), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[232]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[231]  ( .clear(rst), .preset(1'b0), .next_state(N507), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[231]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[230]  ( .clear(rst), .preset(1'b0), .next_state(N506), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[230]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[229]  ( .clear(rst), .preset(1'b0), .next_state(N505), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[229]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[228]  ( .clear(rst), .preset(1'b0), .next_state(N504), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[228]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[227]  ( .clear(rst), .preset(1'b0), .next_state(N503), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[227]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[226]  ( .clear(rst), .preset(1'b0), .next_state(N502), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[226]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[225]  ( .clear(rst), .preset(1'b0), .next_state(N501), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[225]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[224]  ( .clear(rst), .preset(1'b0), .next_state(N500), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[224]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[223]  ( .clear(rst), .preset(1'b0), .next_state(N499), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[223]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[222]  ( .clear(rst), .preset(1'b0), .next_state(N498), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[222]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[221]  ( .clear(rst), .preset(1'b0), .next_state(N497), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[221]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[220]  ( .clear(rst), .preset(1'b0), .next_state(N496), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[220]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[219]  ( .clear(rst), .preset(1'b0), .next_state(N495), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[219]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[218]  ( .clear(rst), .preset(1'b0), .next_state(N494), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[218]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[217]  ( .clear(rst), .preset(1'b0), .next_state(N493), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[217]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[216]  ( .clear(rst), .preset(1'b0), .next_state(N492), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[216]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[215]  ( .clear(rst), .preset(1'b0), .next_state(N491), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[215]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[214]  ( .clear(rst), .preset(1'b0), .next_state(N490), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[214]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[213]  ( .clear(rst), .preset(1'b0), .next_state(N489), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[213]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[212]  ( .clear(rst), .preset(1'b0), .next_state(N488), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[212]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[211]  ( .clear(rst), .preset(1'b0), .next_state(N487), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[211]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[210]  ( .clear(rst), .preset(1'b0), .next_state(N486), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[210]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[209]  ( .clear(rst), .preset(1'b0), .next_state(N485), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[209]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[208]  ( .clear(rst), .preset(1'b0), .next_state(N484), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[208]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[207]  ( .clear(rst), .preset(1'b0), .next_state(N483), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[207]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[206]  ( .clear(rst), .preset(1'b0), .next_state(N482), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[206]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[205]  ( .clear(rst), .preset(1'b0), .next_state(N481), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[205]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[204]  ( .clear(rst), .preset(1'b0), .next_state(N480), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[204]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[203]  ( .clear(rst), .preset(1'b0), .next_state(N479), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[203]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[202]  ( .clear(rst), .preset(1'b0), .next_state(N478), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[202]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[201]  ( .clear(rst), .preset(1'b0), .next_state(N477), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[201]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[200]  ( .clear(rst), .preset(1'b0), .next_state(N476), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[200]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[199]  ( .clear(rst), .preset(1'b0), .next_state(N475), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[199]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[198]  ( .clear(rst), .preset(1'b0), .next_state(N474), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[198]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N473) );
  \**SEQGEN**  \creg_reg[197]  ( .clear(rst), .preset(1'b0), .next_state(N472), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[197]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[196]  ( .clear(rst), .preset(1'b0), .next_state(N471), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[196]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[195]  ( .clear(rst), .preset(1'b0), .next_state(N470), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[195]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[194]  ( .clear(rst), .preset(1'b0), .next_state(N469), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[194]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[193]  ( .clear(rst), .preset(1'b0), .next_state(N468), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[193]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[192]  ( .clear(rst), .preset(1'b0), .next_state(N467), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[192]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[191]  ( .clear(rst), .preset(1'b0), .next_state(N466), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[191]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[190]  ( .clear(rst), .preset(1'b0), .next_state(N465), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[190]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[189]  ( .clear(rst), .preset(1'b0), .next_state(N464), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[189]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[188]  ( .clear(rst), .preset(1'b0), .next_state(N463), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[188]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[187]  ( .clear(rst), .preset(1'b0), .next_state(N462), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[187]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[186]  ( .clear(rst), .preset(1'b0), .next_state(N461), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[186]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[185]  ( .clear(rst), .preset(1'b0), .next_state(N460), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[185]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[184]  ( .clear(rst), .preset(1'b0), .next_state(N459), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[184]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[183]  ( .clear(rst), .preset(1'b0), .next_state(N458), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[183]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[182]  ( .clear(rst), .preset(1'b0), .next_state(N457), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[182]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[181]  ( .clear(rst), .preset(1'b0), .next_state(N456), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[181]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[180]  ( .clear(rst), .preset(1'b0), .next_state(N455), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[180]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[179]  ( .clear(rst), .preset(1'b0), .next_state(N454), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[179]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[178]  ( .clear(rst), .preset(1'b0), .next_state(N453), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[178]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[177]  ( .clear(rst), .preset(1'b0), .next_state(N452), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[177]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[176]  ( .clear(rst), .preset(1'b0), .next_state(N451), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[176]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[175]  ( .clear(rst), .preset(1'b0), .next_state(N450), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[175]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[174]  ( .clear(rst), .preset(1'b0), .next_state(N449), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[174]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[173]  ( .clear(rst), .preset(1'b0), .next_state(N448), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[173]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[172]  ( .clear(rst), .preset(1'b0), .next_state(N447), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[172]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[171]  ( .clear(rst), .preset(1'b0), .next_state(N446), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[171]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[170]  ( .clear(rst), .preset(1'b0), .next_state(N445), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[170]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[169]  ( .clear(rst), .preset(1'b0), .next_state(N444), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[169]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[168]  ( .clear(rst), .preset(1'b0), .next_state(N443), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[168]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[167]  ( .clear(rst), .preset(1'b0), .next_state(N442), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[167]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[166]  ( .clear(rst), .preset(1'b0), .next_state(N441), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[166]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[165]  ( .clear(rst), .preset(1'b0), .next_state(N440), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[165]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[164]  ( .clear(rst), .preset(1'b0), .next_state(N439), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[164]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[163]  ( .clear(rst), .preset(1'b0), .next_state(N438), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[163]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[162]  ( .clear(rst), .preset(1'b0), .next_state(N437), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[162]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[161]  ( .clear(rst), .preset(1'b0), .next_state(N436), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[161]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[160]  ( .clear(rst), .preset(1'b0), .next_state(N435), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[160]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[159]  ( .clear(rst), .preset(1'b0), .next_state(N434), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[159]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[158]  ( .clear(rst), .preset(1'b0), .next_state(N433), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[158]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[157]  ( .clear(rst), .preset(1'b0), .next_state(N432), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[157]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[156]  ( .clear(rst), .preset(1'b0), .next_state(N431), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[156]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[155]  ( .clear(rst), .preset(1'b0), .next_state(N430), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[155]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[154]  ( .clear(rst), .preset(1'b0), .next_state(N429), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[154]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[153]  ( .clear(rst), .preset(1'b0), .next_state(N428), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[153]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[152]  ( .clear(rst), .preset(1'b0), .next_state(N427), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[152]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[151]  ( .clear(rst), .preset(1'b0), .next_state(N426), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[151]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[150]  ( .clear(rst), .preset(1'b0), .next_state(N425), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[150]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[149]  ( .clear(rst), .preset(1'b0), .next_state(N424), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[149]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[148]  ( .clear(rst), .preset(1'b0), .next_state(N423), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[148]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[147]  ( .clear(rst), .preset(1'b0), .next_state(N422), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[147]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[146]  ( .clear(rst), .preset(1'b0), .next_state(N421), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[146]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[145]  ( .clear(rst), .preset(1'b0), .next_state(N420), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[145]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[144]  ( .clear(rst), .preset(1'b0), .next_state(N419), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[144]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[143]  ( .clear(rst), .preset(1'b0), .next_state(N418), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[143]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[142]  ( .clear(rst), .preset(1'b0), .next_state(N417), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[142]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[141]  ( .clear(rst), .preset(1'b0), .next_state(N416), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[141]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[140]  ( .clear(rst), .preset(1'b0), .next_state(N415), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[140]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[139]  ( .clear(rst), .preset(1'b0), .next_state(N414), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[139]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[138]  ( .clear(rst), .preset(1'b0), .next_state(N413), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[138]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[137]  ( .clear(rst), .preset(1'b0), .next_state(N412), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[137]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[136]  ( .clear(rst), .preset(1'b0), .next_state(N411), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[136]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[135]  ( .clear(rst), .preset(1'b0), .next_state(N410), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[135]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[134]  ( .clear(rst), .preset(1'b0), .next_state(N409), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[134]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[133]  ( .clear(rst), .preset(1'b0), .next_state(N408), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[133]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[132]  ( .clear(rst), .preset(1'b0), .next_state(N407), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[132]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[131]  ( .clear(rst), .preset(1'b0), .next_state(N406), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[131]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[130]  ( .clear(rst), .preset(1'b0), .next_state(N405), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[130]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[129]  ( .clear(rst), .preset(1'b0), .next_state(N404), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[129]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[128]  ( .clear(rst), .preset(1'b0), .next_state(N403), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[128]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[127]  ( .clear(rst), .preset(1'b0), .next_state(N402), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[127]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[126]  ( .clear(rst), .preset(1'b0), .next_state(N401), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[126]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[125]  ( .clear(rst), .preset(1'b0), .next_state(N400), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[125]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[124]  ( .clear(rst), .preset(1'b0), .next_state(N399), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[124]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[123]  ( .clear(rst), .preset(1'b0), .next_state(N398), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[123]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[122]  ( .clear(rst), .preset(1'b0), .next_state(N397), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[122]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[121]  ( .clear(rst), .preset(1'b0), .next_state(N396), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[121]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[120]  ( .clear(rst), .preset(1'b0), .next_state(N395), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[120]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[119]  ( .clear(rst), .preset(1'b0), .next_state(N394), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[119]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[118]  ( .clear(rst), .preset(1'b0), .next_state(N393), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[118]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[117]  ( .clear(rst), .preset(1'b0), .next_state(N392), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[117]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[116]  ( .clear(rst), .preset(1'b0), .next_state(N391), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[116]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[115]  ( .clear(rst), .preset(1'b0), .next_state(N390), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[115]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[114]  ( .clear(rst), .preset(1'b0), .next_state(N389), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[114]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[113]  ( .clear(rst), .preset(1'b0), .next_state(N388), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[113]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[112]  ( .clear(rst), .preset(1'b0), .next_state(N387), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[112]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[111]  ( .clear(rst), .preset(1'b0), .next_state(N386), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[111]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[110]  ( .clear(rst), .preset(1'b0), .next_state(N385), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[110]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[109]  ( .clear(rst), .preset(1'b0), .next_state(N384), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[109]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[108]  ( .clear(rst), .preset(1'b0), .next_state(N383), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[108]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[107]  ( .clear(rst), .preset(1'b0), .next_state(N382), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[107]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[106]  ( .clear(rst), .preset(1'b0), .next_state(N381), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[106]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[105]  ( .clear(rst), .preset(1'b0), .next_state(N380), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[105]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[104]  ( .clear(rst), .preset(1'b0), .next_state(N379), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[104]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[103]  ( .clear(rst), .preset(1'b0), .next_state(N378), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[103]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[102]  ( .clear(rst), .preset(1'b0), .next_state(N377), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[102]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[101]  ( .clear(rst), .preset(1'b0), .next_state(N376), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[101]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[100]  ( .clear(rst), .preset(1'b0), .next_state(N375), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[100]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[99]  ( .clear(rst), .preset(1'b0), .next_state(N374), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[99]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N373) );
  \**SEQGEN**  \creg_reg[98]  ( .clear(rst), .preset(1'b0), .next_state(N372), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[98]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[97]  ( .clear(rst), .preset(1'b0), .next_state(N371), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[97]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[96]  ( .clear(rst), .preset(1'b0), .next_state(N370), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[96]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[95]  ( .clear(rst), .preset(1'b0), .next_state(N369), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[95]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[94]  ( .clear(rst), .preset(1'b0), .next_state(N368), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[94]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[93]  ( .clear(rst), .preset(1'b0), .next_state(N367), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[93]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[92]  ( .clear(rst), .preset(1'b0), .next_state(N366), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[92]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[91]  ( .clear(rst), .preset(1'b0), .next_state(N365), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[91]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[90]  ( .clear(rst), .preset(1'b0), .next_state(N364), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[90]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[89]  ( .clear(rst), .preset(1'b0), .next_state(N363), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[89]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[88]  ( .clear(rst), .preset(1'b0), .next_state(N362), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[88]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[87]  ( .clear(rst), .preset(1'b0), .next_state(N361), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[87]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[86]  ( .clear(rst), .preset(1'b0), .next_state(N360), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[86]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[85]  ( .clear(rst), .preset(1'b0), .next_state(N359), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[85]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[84]  ( .clear(rst), .preset(1'b0), .next_state(N358), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[84]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[83]  ( .clear(rst), .preset(1'b0), .next_state(N357), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[83]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[82]  ( .clear(rst), .preset(1'b0), .next_state(N356), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[82]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[81]  ( .clear(rst), .preset(1'b0), .next_state(N355), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[81]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[80]  ( .clear(rst), .preset(1'b0), .next_state(N354), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[80]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[79]  ( .clear(rst), .preset(1'b0), .next_state(N353), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[79]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[78]  ( .clear(rst), .preset(1'b0), .next_state(N352), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[78]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[77]  ( .clear(rst), .preset(1'b0), .next_state(N351), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[77]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[76]  ( .clear(rst), .preset(1'b0), .next_state(N350), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[76]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[75]  ( .clear(rst), .preset(1'b0), .next_state(N349), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[75]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[74]  ( .clear(rst), .preset(1'b0), .next_state(N348), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[74]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[73]  ( .clear(rst), .preset(1'b0), .next_state(N347), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[73]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[72]  ( .clear(rst), .preset(1'b0), .next_state(N346), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[72]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[71]  ( .clear(rst), .preset(1'b0), .next_state(N345), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[71]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[70]  ( .clear(rst), .preset(1'b0), .next_state(N344), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[70]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[69]  ( .clear(rst), .preset(1'b0), .next_state(N343), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[69]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[68]  ( .clear(rst), .preset(1'b0), .next_state(N342), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[68]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[67]  ( .clear(rst), .preset(1'b0), .next_state(N341), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[67]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[66]  ( .clear(rst), .preset(1'b0), .next_state(N340), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[66]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[65]  ( .clear(rst), .preset(1'b0), .next_state(N339), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[65]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[64]  ( .clear(rst), .preset(1'b0), .next_state(N338), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[64]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[63]  ( .clear(rst), .preset(1'b0), .next_state(N337), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[63]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[62]  ( .clear(rst), .preset(1'b0), .next_state(N336), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[62]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[61]  ( .clear(rst), .preset(1'b0), .next_state(N335), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[61]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[60]  ( .clear(rst), .preset(1'b0), .next_state(N334), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[60]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[59]  ( .clear(rst), .preset(1'b0), .next_state(N333), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[59]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[58]  ( .clear(rst), .preset(1'b0), .next_state(N332), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[58]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[57]  ( .clear(rst), .preset(1'b0), .next_state(N331), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[57]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[56]  ( .clear(rst), .preset(1'b0), .next_state(N330), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[56]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[55]  ( .clear(rst), .preset(1'b0), .next_state(N329), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[55]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[54]  ( .clear(rst), .preset(1'b0), .next_state(N328), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[54]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[53]  ( .clear(rst), .preset(1'b0), .next_state(N327), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[53]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[52]  ( .clear(rst), .preset(1'b0), .next_state(N326), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[52]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[51]  ( .clear(rst), .preset(1'b0), .next_state(N325), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[51]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[50]  ( .clear(rst), .preset(1'b0), .next_state(N324), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[50]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[49]  ( .clear(rst), .preset(1'b0), .next_state(N323), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[49]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[48]  ( .clear(rst), .preset(1'b0), .next_state(N322), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[48]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[47]  ( .clear(rst), .preset(1'b0), .next_state(N321), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[47]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[46]  ( .clear(rst), .preset(1'b0), .next_state(N320), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[46]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[45]  ( .clear(rst), .preset(1'b0), .next_state(N319), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[45]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[44]  ( .clear(rst), .preset(1'b0), .next_state(N318), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[44]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[43]  ( .clear(rst), .preset(1'b0), .next_state(N317), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[43]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[42]  ( .clear(rst), .preset(1'b0), .next_state(N316), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[42]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[41]  ( .clear(rst), .preset(1'b0), .next_state(N315), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[41]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[40]  ( .clear(rst), .preset(1'b0), .next_state(N314), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[40]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[39]  ( .clear(rst), .preset(1'b0), .next_state(N313), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[39]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[38]  ( .clear(rst), .preset(1'b0), .next_state(N312), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[38]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[37]  ( .clear(rst), .preset(1'b0), .next_state(N311), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[37]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[36]  ( .clear(rst), .preset(1'b0), .next_state(N310), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[36]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[35]  ( .clear(rst), .preset(1'b0), .next_state(N309), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[35]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[34]  ( .clear(rst), .preset(1'b0), .next_state(N308), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[34]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[33]  ( .clear(rst), .preset(1'b0), .next_state(N307), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[33]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[32]  ( .clear(rst), .preset(1'b0), .next_state(N306), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[32]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[31]  ( .clear(rst), .preset(1'b0), .next_state(N305), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[31]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[30]  ( .clear(rst), .preset(1'b0), .next_state(N304), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[30]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[29]  ( .clear(rst), .preset(1'b0), .next_state(N303), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[29]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[28]  ( .clear(rst), .preset(1'b0), .next_state(N302), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[28]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[27]  ( .clear(rst), .preset(1'b0), .next_state(N301), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[27]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[26]  ( .clear(rst), .preset(1'b0), .next_state(N300), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[26]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[25]  ( .clear(rst), .preset(1'b0), .next_state(N299), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[25]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[24]  ( .clear(rst), .preset(1'b0), .next_state(N298), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[24]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[23]  ( .clear(rst), .preset(1'b0), .next_state(N297), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[23]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[22]  ( .clear(rst), .preset(1'b0), .next_state(N296), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[22]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[21]  ( .clear(rst), .preset(1'b0), .next_state(N295), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[21]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[20]  ( .clear(rst), .preset(1'b0), .next_state(N294), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[20]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[19]  ( .clear(rst), .preset(1'b0), .next_state(N293), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[19]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[18]  ( .clear(rst), .preset(1'b0), .next_state(N292), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[18]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[17]  ( .clear(rst), .preset(1'b0), .next_state(N291), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[17]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[16]  ( .clear(rst), .preset(1'b0), .next_state(N290), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[16]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[15]  ( .clear(rst), .preset(1'b0), .next_state(N289), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[15]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[14]  ( .clear(rst), .preset(1'b0), .next_state(N288), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[14]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[13]  ( .clear(rst), .preset(1'b0), .next_state(N287), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[13]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[12]  ( .clear(rst), .preset(1'b0), .next_state(N286), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[12]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[11]  ( .clear(rst), .preset(1'b0), .next_state(N285), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[11]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[10]  ( .clear(rst), .preset(1'b0), .next_state(N284), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[10]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[9]  ( .clear(rst), .preset(1'b0), .next_state(N283), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[9]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[8]  ( .clear(rst), .preset(1'b0), .next_state(N282), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[8]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[7]  ( .clear(rst), .preset(1'b0), .next_state(N281), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[7]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[6]  ( .clear(rst), .preset(1'b0), .next_state(N280), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[6]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[5]  ( .clear(rst), .preset(1'b0), .next_state(N279), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[5]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[4]  ( .clear(rst), .preset(1'b0), .next_state(N278), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[4]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[3]  ( .clear(rst), .preset(1'b0), .next_state(N277), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[3]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[2]  ( .clear(rst), .preset(1'b0), .next_state(N276), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[2]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[1]  ( .clear(rst), .preset(1'b0), .next_state(N275), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[1]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \creg_reg[0]  ( .clear(rst), .preset(1'b0), .next_state(N274), 
        .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(creg[0]), 
        .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(1'b0), 
        .synch_enable(N273) );
  \**SEQGEN**  \start_reg_reg[255]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[254]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[255]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[254]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[253]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[254]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[253]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[252]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[253]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[252]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[251]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[252]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[251]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[250]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[251]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[250]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[249]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[250]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[249]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[248]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[249]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[248]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[247]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[248]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[247]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[246]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[247]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[246]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[245]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[246]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[245]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[244]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[245]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[244]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[243]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[244]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[243]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[242]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[243]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[242]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[241]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[242]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[241]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[240]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[241]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[240]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[239]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[240]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[239]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[238]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[239]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[238]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[237]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[238]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[237]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[236]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[237]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[236]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[235]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[236]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[235]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[234]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[235]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[234]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[233]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[234]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[233]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[232]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[233]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[232]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[231]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[232]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[231]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[230]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[231]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[230]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[229]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[230]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[229]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[228]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[229]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[228]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[227]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[228]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[227]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[226]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[227]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[226]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[225]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[226]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[225]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[224]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[225]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[224]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[223]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[224]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[223]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[222]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[223]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[222]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[221]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[222]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[221]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[220]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[221]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[220]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[219]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[220]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[219]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[218]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[219]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[218]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[217]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[218]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[217]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[216]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[217]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[216]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[215]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[216]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[215]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[214]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[215]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[214]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[213]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[214]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[213]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[212]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[213]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[212]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[211]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[212]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[211]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[210]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[211]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[210]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[209]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[210]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[209]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[208]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[209]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[208]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[207]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[208]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[207]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[206]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[207]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[206]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[205]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[206]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[205]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[204]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[205]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[204]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[203]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[204]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[203]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[202]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[203]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[202]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[201]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[202]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[201]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[200]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[201]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[200]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[199]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[200]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[199]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[198]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[199]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[198]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[197]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[198]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[197]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[196]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[197]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[196]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[195]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[196]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[195]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[194]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[195]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[194]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[193]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[194]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[193]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[192]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[193]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[192]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[191]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[192]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[191]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[190]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[191]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[190]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[189]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[190]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[189]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[188]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[189]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[188]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[187]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[188]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[187]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[186]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[187]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[186]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[185]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[186]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[185]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[184]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[185]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[184]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[183]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[184]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[183]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[182]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[183]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[182]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[181]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[182]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[181]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[180]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[181]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[180]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[179]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[180]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[179]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[178]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[179]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[178]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[177]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[178]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[177]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[176]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[177]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[176]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[175]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[176]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[175]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[174]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[175]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[174]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[173]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[174]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[173]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[172]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[173]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[172]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[171]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[172]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[171]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[170]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[171]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[170]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[169]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[170]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[169]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[168]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[169]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[168]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[167]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[168]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[167]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[166]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[167]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[166]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[165]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[166]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[165]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[164]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[165]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[164]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[163]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[164]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[163]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[162]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[163]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[162]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[161]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[162]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[161]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[160]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[161]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[160]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[159]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[160]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[159]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[158]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[159]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[158]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[157]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[158]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[157]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[156]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[157]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[156]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[155]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[156]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[155]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[154]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[155]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[154]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[153]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[154]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[153]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[152]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[153]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[152]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[151]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[152]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[151]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[150]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[151]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[150]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[149]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[150]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[149]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[148]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[149]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[148]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[147]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[148]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[147]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[146]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[147]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[146]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[145]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[146]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[145]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[144]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[145]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[144]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[143]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[144]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[143]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[142]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[143]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[142]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[141]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[142]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[141]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[140]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[141]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[140]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[139]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[140]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[139]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[138]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[139]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[138]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[137]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[138]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[137]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[136]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[137]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[136]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[135]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[136]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[135]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[134]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[135]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[134]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[133]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[134]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[133]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[132]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[133]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[132]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[131]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[132]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[131]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[130]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[131]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[130]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[129]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[130]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[129]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[128]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[129]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[128]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[127]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[128]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[127]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[126]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[127]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[126]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[125]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[126]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[125]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[124]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[125]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[124]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[123]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[124]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[123]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[122]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[123]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[122]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[121]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[122]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[121]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[120]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[121]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[120]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[119]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[120]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[119]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[118]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[119]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[118]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[117]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[118]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[117]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[116]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[117]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[116]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[115]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[116]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[115]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[114]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[115]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[114]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[113]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[114]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[113]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[112]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[113]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[112]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[111]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[112]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[111]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[110]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[111]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[110]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[109]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[110]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[109]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[108]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[109]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[108]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[107]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[108]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[107]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[106]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[107]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[106]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[105]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[106]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[105]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[104]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[105]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[104]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[103]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[104]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[103]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[102]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[103]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[102]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[101]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[102]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[101]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[100]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[101]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[100]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[99]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[100]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[99]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[98]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[99]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[98]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[97]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[98]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[97]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[96]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[97]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[96]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[95]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[96]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[95]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[94]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[95]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[94]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[93]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[94]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[93]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[92]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[93]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[92]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[91]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[92]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[91]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[90]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[91]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[90]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[89]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[90]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[89]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[88]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[89]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[88]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[87]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[88]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[87]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[86]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[87]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[86]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[85]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[86]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[85]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[84]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[85]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[84]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[83]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[84]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[83]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[82]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[83]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[82]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[81]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[82]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[81]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[80]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[81]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[80]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[79]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[80]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[79]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[78]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[79]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[78]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[77]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[78]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[77]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[76]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[77]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[76]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[75]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[76]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[75]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[74]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[75]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[74]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[73]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[74]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[73]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[72]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[73]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[72]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[71]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[72]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[71]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[70]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[71]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[70]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[69]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[70]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[69]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[68]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[69]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[68]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[67]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[68]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[67]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[66]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[67]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[66]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[65]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[66]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[65]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[64]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[65]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[64]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[63]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[64]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[63]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[62]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[63]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[62]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[61]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[62]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[61]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[60]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[61]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[60]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[59]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[60]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[59]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[58]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[59]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[58]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[57]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[58]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[57]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[56]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[57]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[56]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[55]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[56]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[55]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[54]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[55]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[54]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[53]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[54]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[53]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[52]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[53]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[52]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[51]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[52]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[51]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[50]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[51]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[50]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[49]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[50]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[49]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[48]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[49]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[48]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[47]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[48]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[47]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[46]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[47]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[46]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[45]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[46]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[45]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[44]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[45]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[44]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[43]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[44]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[43]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[42]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[43]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[42]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[41]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[42]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[41]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[40]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[41]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[40]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[39]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[40]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[39]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[38]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[39]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[38]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[37]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[38]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[37]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[36]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[37]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[36]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[35]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[36]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[35]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[34]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[35]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[34]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[33]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[34]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[33]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[32]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[33]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[32]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[32]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[31]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[31]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[30]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[30]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[29]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[29]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[28]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[28]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[27]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[27]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[26]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[26]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[25]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[25]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[24]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[24]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[23]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[23]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[22]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[22]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[21]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[21]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[20]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[20]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[19]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[19]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[18]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[18]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[17]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[17]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[16]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[16]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[15]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[15]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[14]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[14]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[13]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[13]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[12]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[12]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[11]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[11]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[10]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[10]), .synch_clear(1'b0), .synch_preset(1'b0), 
        .synch_toggle(1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[9]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[8]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[7]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[6]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[5]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[4]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[3]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[2]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[1]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \start_reg_reg[0]  ( .clear(rst), .preset(1'b0), .next_state(
        start_in[255]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        start_reg[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  modmult_N256_CC256_1 modmult_1 ( .clk(clk), .rst(rst), .start(start_in[0]), 
        .x(x), .y(y), .n(n), .o(o) );
  GTECH_OR2 C4972 ( .A(mul_pow), .B(N535), .Z(N538) );
  GTECH_OR2 C5484 ( .A(N5), .B(N9), .Z(N539) );
  GTECH_OR2 C5486 ( .A(N11), .B(N12), .Z(N13) );
  SELECT_OP C5998 ( .DATA1(start_reg), .DATA2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), 
        .CONTROL1(N0), .CONTROL2(N1), .Z(start_in) );
  GTECH_BUF B_0 ( .A(init), .Z(N0) );
  GTECH_BUF B_1 ( .A(N5), .Z(N1) );
  SELECT_OP C5999 ( .DATA1(ereg), .DATA2(e), .CONTROL1(N0), .CONTROL2(N1), .Z(
        ein) );
  SELECT_OP C6000 ( .DATA1(o), .DATA2(creg), .CONTROL1(N2), .CONTROL2(N6), .Z(
        c) );
  GTECH_BUF B_2 ( .A(ein[255]), .Z(N2) );
  SELECT_OP C6001 ( .DATA1({1'b1, 1'b1, 1'b1}), .DATA2({mul_pow, mul_pow, 
        mul_pow}), .DATA3({1'b0, 1'b0, 1'b0}), .CONTROL1(N1), .CONTROL2(N533), 
        .CONTROL3(N9), .Z({N214, N114, N14}) );
  SELECT_OP C6002 ( .DATA1(e), .DATA2({ein[254:0], 1'b0}), .CONTROL1(N1), 
        .CONTROL2(N533), .Z({N272, N271, N270, N269, N268, N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, 
        N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, 
        N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, 
        N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, 
        N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, 
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, 
        N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, 
        N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, 
        N119, N118, N117, N116, N115, N113, N112, N111, N110, N109, N108, N107, 
        N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, 
        N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, 
        N23, N22, N21, N20, N19, N18, N17, N16, N15}) );
  SELECT_OP C6003 ( .DATA1({1'b1, 1'b1, 1'b1}), .DATA2({N13, N13, N13}), 
        .DATA3({1'b0, 1'b0, 1'b0}), .CONTROL1(N1), .CONTROL2(N533), .CONTROL3(
        N9), .Z({N473, N373, N273}) );
  SELECT_OP C6004 ( .DATA1(m), .DATA2(o), .CONTROL1(N1), .CONTROL2(N533), .Z({
        N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, 
        N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, 
        N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, 
        N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, 
        N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N472, N471, 
        N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, 
        N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, 
        N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, 
        N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, 
        N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, 
        N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, 
        N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, 
        N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, 
        N374, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, 
        N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, 
        N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, 
        N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, 
        N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, 
        N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, 
        N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, 
        N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, 
        N277, N276, N275, N274}) );
  SELECT_OP C6005 ( .DATA1(1'b0), .DATA2(N10), .CONTROL1(N3), .CONTROL2(N533), 
        .Z(N532) );
  GTECH_BUF B_3 ( .A(N539), .Z(N3) );
  SELECT_OP C6006 ( .DATA1(creg), .DATA2(m), .CONTROL1(N0), .CONTROL2(N1), .Z(
        x) );
  SELECT_OP C6007 ( .DATA1(m), .DATA2(creg), .CONTROL1(N4), .CONTROL2(N537), 
        .Z(y) );
  GTECH_BUF B_4 ( .A(N538), .Z(N4) );
  GTECH_NOT I_0 ( .A(init), .Z(N5) );
  GTECH_NOT I_1 ( .A(ein[255]), .Z(N6) );
  GTECH_NOT I_2 ( .A(mul_pow), .Z(N7) );
  GTECH_OR2 C6023 ( .A(start_in[255]), .B(N5), .Z(N8) );
  GTECH_NOT I_3 ( .A(N8), .Z(N9) );
  GTECH_AND2 C6025 ( .A(ein[255]), .B(mul_pow), .Z(N10) );
  GTECH_AND2 C6027 ( .A(N540), .B(mul_pow), .Z(N11) );
  GTECH_AND2 C6028 ( .A(first_one), .B(ein[255]), .Z(N540) );
  GTECH_AND2 C6029 ( .A(first_one), .B(N7), .Z(N12) );
  GTECH_AND2 C6036 ( .A(start_in[255]), .B(init), .Z(N533) );
  GTECH_OR2 C6042 ( .A(init), .B(mul_pow), .Z(N534) );
  GTECH_NOT I_4 ( .A(N534), .Z(N535) );
  GTECH_NOT I_5 ( .A(mul_pow), .Z(N536) );
  GTECH_AND2 C6045 ( .A(init), .B(N536), .Z(N537) );
endmodule

