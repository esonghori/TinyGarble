
module mult_N1024_CC1024 ( clk, rst, g_input, e_input, o );
  input [1023:0] g_input;
  input [0:0] e_input;
  output [2047:0] o;
  input clk, rst;
  wire   \add_42/carry[2047] , \add_42/carry[2046] , \add_42/carry[2045] ,
         \add_42/carry[2044] , \add_42/carry[2043] , \add_42/carry[2042] ,
         \add_42/carry[2041] , \add_42/carry[2040] , \add_42/carry[2039] ,
         \add_42/carry[2038] , \add_42/carry[2037] , \add_42/carry[2036] ,
         \add_42/carry[2035] , \add_42/carry[2034] , \add_42/carry[2033] ,
         \add_42/carry[2032] , \add_42/carry[2031] , \add_42/carry[2030] ,
         \add_42/carry[2029] , \add_42/carry[2028] , \add_42/carry[2027] ,
         \add_42/carry[2026] , \add_42/carry[2025] , \add_42/carry[2024] ,
         \add_42/carry[2023] , \add_42/carry[2022] , \add_42/carry[2021] ,
         \add_42/carry[2020] , \add_42/carry[2019] , \add_42/carry[2018] ,
         \add_42/carry[2017] , \add_42/carry[2016] , \add_42/carry[2015] ,
         \add_42/carry[2014] , \add_42/carry[2013] , \add_42/carry[2012] ,
         \add_42/carry[2011] , \add_42/carry[2010] , \add_42/carry[2009] ,
         \add_42/carry[2008] , \add_42/carry[2007] , \add_42/carry[2006] ,
         \add_42/carry[2005] , \add_42/carry[2004] , \add_42/carry[2003] ,
         \add_42/carry[2002] , \add_42/carry[2001] , \add_42/carry[2000] ,
         \add_42/carry[1999] , \add_42/carry[1998] , \add_42/carry[1997] ,
         \add_42/carry[1996] , \add_42/carry[1995] , \add_42/carry[1994] ,
         \add_42/carry[1993] , \add_42/carry[1992] , \add_42/carry[1991] ,
         \add_42/carry[1990] , \add_42/carry[1989] , \add_42/carry[1988] ,
         \add_42/carry[1987] , \add_42/carry[1986] , \add_42/carry[1985] ,
         \add_42/carry[1984] , \add_42/carry[1983] , \add_42/carry[1982] ,
         \add_42/carry[1981] , \add_42/carry[1980] , \add_42/carry[1979] ,
         \add_42/carry[1978] , \add_42/carry[1977] , \add_42/carry[1976] ,
         \add_42/carry[1975] , \add_42/carry[1974] , \add_42/carry[1973] ,
         \add_42/carry[1972] , \add_42/carry[1971] , \add_42/carry[1970] ,
         \add_42/carry[1969] , \add_42/carry[1968] , \add_42/carry[1967] ,
         \add_42/carry[1966] , \add_42/carry[1965] , \add_42/carry[1964] ,
         \add_42/carry[1963] , \add_42/carry[1962] , \add_42/carry[1961] ,
         \add_42/carry[1960] , \add_42/carry[1959] , \add_42/carry[1958] ,
         \add_42/carry[1957] , \add_42/carry[1956] , \add_42/carry[1955] ,
         \add_42/carry[1954] , \add_42/carry[1953] , \add_42/carry[1952] ,
         \add_42/carry[1951] , \add_42/carry[1950] , \add_42/carry[1949] ,
         \add_42/carry[1948] , \add_42/carry[1947] , \add_42/carry[1946] ,
         \add_42/carry[1945] , \add_42/carry[1944] , \add_42/carry[1943] ,
         \add_42/carry[1942] , \add_42/carry[1941] , \add_42/carry[1940] ,
         \add_42/carry[1939] , \add_42/carry[1938] , \add_42/carry[1937] ,
         \add_42/carry[1936] , \add_42/carry[1935] , \add_42/carry[1934] ,
         \add_42/carry[1933] , \add_42/carry[1932] , \add_42/carry[1931] ,
         \add_42/carry[1930] , \add_42/carry[1929] , \add_42/carry[1928] ,
         \add_42/carry[1927] , \add_42/carry[1926] , \add_42/carry[1925] ,
         \add_42/carry[1924] , \add_42/carry[1923] , \add_42/carry[1922] ,
         \add_42/carry[1921] , \add_42/carry[1920] , \add_42/carry[1919] ,
         \add_42/carry[1918] , \add_42/carry[1917] , \add_42/carry[1916] ,
         \add_42/carry[1915] , \add_42/carry[1914] , \add_42/carry[1913] ,
         \add_42/carry[1912] , \add_42/carry[1911] , \add_42/carry[1910] ,
         \add_42/carry[1909] , \add_42/carry[1908] , \add_42/carry[1907] ,
         \add_42/carry[1906] , \add_42/carry[1905] , \add_42/carry[1904] ,
         \add_42/carry[1903] , \add_42/carry[1902] , \add_42/carry[1901] ,
         \add_42/carry[1900] , \add_42/carry[1899] , \add_42/carry[1898] ,
         \add_42/carry[1897] , \add_42/carry[1896] , \add_42/carry[1895] ,
         \add_42/carry[1894] , \add_42/carry[1893] , \add_42/carry[1892] ,
         \add_42/carry[1891] , \add_42/carry[1890] , \add_42/carry[1889] ,
         \add_42/carry[1888] , \add_42/carry[1887] , \add_42/carry[1886] ,
         \add_42/carry[1885] , \add_42/carry[1884] , \add_42/carry[1883] ,
         \add_42/carry[1882] , \add_42/carry[1881] , \add_42/carry[1880] ,
         \add_42/carry[1879] , \add_42/carry[1878] , \add_42/carry[1877] ,
         \add_42/carry[1876] , \add_42/carry[1875] , \add_42/carry[1874] ,
         \add_42/carry[1873] , \add_42/carry[1872] , \add_42/carry[1871] ,
         \add_42/carry[1870] , \add_42/carry[1869] , \add_42/carry[1868] ,
         \add_42/carry[1867] , \add_42/carry[1866] , \add_42/carry[1865] ,
         \add_42/carry[1864] , \add_42/carry[1863] , \add_42/carry[1862] ,
         \add_42/carry[1861] , \add_42/carry[1860] , \add_42/carry[1859] ,
         \add_42/carry[1858] , \add_42/carry[1857] , \add_42/carry[1856] ,
         \add_42/carry[1855] , \add_42/carry[1854] , \add_42/carry[1853] ,
         \add_42/carry[1852] , \add_42/carry[1851] , \add_42/carry[1850] ,
         \add_42/carry[1849] , \add_42/carry[1848] , \add_42/carry[1847] ,
         \add_42/carry[1846] , \add_42/carry[1845] , \add_42/carry[1844] ,
         \add_42/carry[1843] , \add_42/carry[1842] , \add_42/carry[1841] ,
         \add_42/carry[1840] , \add_42/carry[1839] , \add_42/carry[1838] ,
         \add_42/carry[1837] , \add_42/carry[1836] , \add_42/carry[1835] ,
         \add_42/carry[1834] , \add_42/carry[1833] , \add_42/carry[1832] ,
         \add_42/carry[1831] , \add_42/carry[1830] , \add_42/carry[1829] ,
         \add_42/carry[1828] , \add_42/carry[1827] , \add_42/carry[1826] ,
         \add_42/carry[1825] , \add_42/carry[1824] , \add_42/carry[1823] ,
         \add_42/carry[1822] , \add_42/carry[1821] , \add_42/carry[1820] ,
         \add_42/carry[1819] , \add_42/carry[1818] , \add_42/carry[1817] ,
         \add_42/carry[1816] , \add_42/carry[1815] , \add_42/carry[1814] ,
         \add_42/carry[1813] , \add_42/carry[1812] , \add_42/carry[1811] ,
         \add_42/carry[1810] , \add_42/carry[1809] , \add_42/carry[1808] ,
         \add_42/carry[1807] , \add_42/carry[1806] , \add_42/carry[1805] ,
         \add_42/carry[1804] , \add_42/carry[1803] , \add_42/carry[1802] ,
         \add_42/carry[1801] , \add_42/carry[1800] , \add_42/carry[1799] ,
         \add_42/carry[1798] , \add_42/carry[1797] , \add_42/carry[1796] ,
         \add_42/carry[1795] , \add_42/carry[1794] , \add_42/carry[1793] ,
         \add_42/carry[1792] , \add_42/carry[1791] , \add_42/carry[1790] ,
         \add_42/carry[1789] , \add_42/carry[1788] , \add_42/carry[1787] ,
         \add_42/carry[1786] , \add_42/carry[1785] , \add_42/carry[1784] ,
         \add_42/carry[1783] , \add_42/carry[1782] , \add_42/carry[1781] ,
         \add_42/carry[1780] , \add_42/carry[1779] , \add_42/carry[1778] ,
         \add_42/carry[1777] , \add_42/carry[1776] , \add_42/carry[1775] ,
         \add_42/carry[1774] , \add_42/carry[1773] , \add_42/carry[1772] ,
         \add_42/carry[1771] , \add_42/carry[1770] , \add_42/carry[1769] ,
         \add_42/carry[1768] , \add_42/carry[1767] , \add_42/carry[1766] ,
         \add_42/carry[1765] , \add_42/carry[1764] , \add_42/carry[1763] ,
         \add_42/carry[1762] , \add_42/carry[1761] , \add_42/carry[1760] ,
         \add_42/carry[1759] , \add_42/carry[1758] , \add_42/carry[1757] ,
         \add_42/carry[1756] , \add_42/carry[1755] , \add_42/carry[1754] ,
         \add_42/carry[1753] , \add_42/carry[1752] , \add_42/carry[1751] ,
         \add_42/carry[1750] , \add_42/carry[1749] , \add_42/carry[1748] ,
         \add_42/carry[1747] , \add_42/carry[1746] , \add_42/carry[1745] ,
         \add_42/carry[1744] , \add_42/carry[1743] , \add_42/carry[1742] ,
         \add_42/carry[1741] , \add_42/carry[1740] , \add_42/carry[1739] ,
         \add_42/carry[1738] , \add_42/carry[1737] , \add_42/carry[1736] ,
         \add_42/carry[1735] , \add_42/carry[1734] , \add_42/carry[1733] ,
         \add_42/carry[1732] , \add_42/carry[1731] , \add_42/carry[1730] ,
         \add_42/carry[1729] , \add_42/carry[1728] , \add_42/carry[1727] ,
         \add_42/carry[1726] , \add_42/carry[1725] , \add_42/carry[1724] ,
         \add_42/carry[1723] , \add_42/carry[1722] , \add_42/carry[1721] ,
         \add_42/carry[1720] , \add_42/carry[1719] , \add_42/carry[1718] ,
         \add_42/carry[1717] , \add_42/carry[1716] , \add_42/carry[1715] ,
         \add_42/carry[1714] , \add_42/carry[1713] , \add_42/carry[1712] ,
         \add_42/carry[1711] , \add_42/carry[1710] , \add_42/carry[1709] ,
         \add_42/carry[1708] , \add_42/carry[1707] , \add_42/carry[1706] ,
         \add_42/carry[1705] , \add_42/carry[1704] , \add_42/carry[1703] ,
         \add_42/carry[1702] , \add_42/carry[1701] , \add_42/carry[1700] ,
         \add_42/carry[1699] , \add_42/carry[1698] , \add_42/carry[1697] ,
         \add_42/carry[1696] , \add_42/carry[1695] , \add_42/carry[1694] ,
         \add_42/carry[1693] , \add_42/carry[1692] , \add_42/carry[1691] ,
         \add_42/carry[1690] , \add_42/carry[1689] , \add_42/carry[1688] ,
         \add_42/carry[1687] , \add_42/carry[1686] , \add_42/carry[1685] ,
         \add_42/carry[1684] , \add_42/carry[1683] , \add_42/carry[1682] ,
         \add_42/carry[1681] , \add_42/carry[1680] , \add_42/carry[1679] ,
         \add_42/carry[1678] , \add_42/carry[1677] , \add_42/carry[1676] ,
         \add_42/carry[1675] , \add_42/carry[1674] , \add_42/carry[1673] ,
         \add_42/carry[1672] , \add_42/carry[1671] , \add_42/carry[1670] ,
         \add_42/carry[1669] , \add_42/carry[1668] , \add_42/carry[1667] ,
         \add_42/carry[1666] , \add_42/carry[1665] , \add_42/carry[1664] ,
         \add_42/carry[1663] , \add_42/carry[1662] , \add_42/carry[1661] ,
         \add_42/carry[1660] , \add_42/carry[1659] , \add_42/carry[1658] ,
         \add_42/carry[1657] , \add_42/carry[1656] , \add_42/carry[1655] ,
         \add_42/carry[1654] , \add_42/carry[1653] , \add_42/carry[1652] ,
         \add_42/carry[1651] , \add_42/carry[1650] , \add_42/carry[1649] ,
         \add_42/carry[1648] , \add_42/carry[1647] , \add_42/carry[1646] ,
         \add_42/carry[1645] , \add_42/carry[1644] , \add_42/carry[1643] ,
         \add_42/carry[1642] , \add_42/carry[1641] , \add_42/carry[1640] ,
         \add_42/carry[1639] , \add_42/carry[1638] , \add_42/carry[1637] ,
         \add_42/carry[1636] , \add_42/carry[1635] , \add_42/carry[1634] ,
         \add_42/carry[1633] , \add_42/carry[1632] , \add_42/carry[1631] ,
         \add_42/carry[1630] , \add_42/carry[1629] , \add_42/carry[1628] ,
         \add_42/carry[1627] , \add_42/carry[1626] , \add_42/carry[1625] ,
         \add_42/carry[1624] , \add_42/carry[1623] , \add_42/carry[1622] ,
         \add_42/carry[1621] , \add_42/carry[1620] , \add_42/carry[1619] ,
         \add_42/carry[1618] , \add_42/carry[1617] , \add_42/carry[1616] ,
         \add_42/carry[1615] , \add_42/carry[1614] , \add_42/carry[1613] ,
         \add_42/carry[1612] , \add_42/carry[1611] , \add_42/carry[1610] ,
         \add_42/carry[1609] , \add_42/carry[1608] , \add_42/carry[1607] ,
         \add_42/carry[1606] , \add_42/carry[1605] , \add_42/carry[1604] ,
         \add_42/carry[1603] , \add_42/carry[1602] , \add_42/carry[1601] ,
         \add_42/carry[1600] , \add_42/carry[1599] , \add_42/carry[1598] ,
         \add_42/carry[1597] , \add_42/carry[1596] , \add_42/carry[1595] ,
         \add_42/carry[1594] , \add_42/carry[1593] , \add_42/carry[1592] ,
         \add_42/carry[1591] , \add_42/carry[1590] , \add_42/carry[1589] ,
         \add_42/carry[1588] , \add_42/carry[1587] , \add_42/carry[1586] ,
         \add_42/carry[1585] , \add_42/carry[1584] , \add_42/carry[1583] ,
         \add_42/carry[1582] , \add_42/carry[1581] , \add_42/carry[1580] ,
         \add_42/carry[1579] , \add_42/carry[1578] , \add_42/carry[1577] ,
         \add_42/carry[1576] , \add_42/carry[1575] , \add_42/carry[1574] ,
         \add_42/carry[1573] , \add_42/carry[1572] , \add_42/carry[1571] ,
         \add_42/carry[1570] , \add_42/carry[1569] , \add_42/carry[1568] ,
         \add_42/carry[1567] , \add_42/carry[1566] , \add_42/carry[1565] ,
         \add_42/carry[1564] , \add_42/carry[1563] , \add_42/carry[1562] ,
         \add_42/carry[1561] , \add_42/carry[1560] , \add_42/carry[1559] ,
         \add_42/carry[1558] , \add_42/carry[1557] , \add_42/carry[1556] ,
         \add_42/carry[1555] , \add_42/carry[1554] , \add_42/carry[1553] ,
         \add_42/carry[1552] , \add_42/carry[1551] , \add_42/carry[1550] ,
         \add_42/carry[1549] , \add_42/carry[1548] , \add_42/carry[1547] ,
         \add_42/carry[1546] , \add_42/carry[1545] , \add_42/carry[1544] ,
         \add_42/carry[1543] , \add_42/carry[1542] , \add_42/carry[1541] ,
         \add_42/carry[1540] , \add_42/carry[1539] , \add_42/carry[1538] ,
         \add_42/carry[1537] , \add_42/carry[1536] , \add_42/carry[1535] ,
         \add_42/carry[1534] , \add_42/carry[1533] , \add_42/carry[1532] ,
         \add_42/carry[1531] , \add_42/carry[1530] , \add_42/carry[1529] ,
         \add_42/carry[1528] , \add_42/carry[1527] , \add_42/carry[1526] ,
         \add_42/carry[1525] , \add_42/carry[1524] , \add_42/carry[1523] ,
         \add_42/carry[1522] , \add_42/carry[1521] , \add_42/carry[1520] ,
         \add_42/carry[1519] , \add_42/carry[1518] , \add_42/carry[1517] ,
         \add_42/carry[1516] , \add_42/carry[1515] , \add_42/carry[1514] ,
         \add_42/carry[1513] , \add_42/carry[1512] , \add_42/carry[1511] ,
         \add_42/carry[1510] , \add_42/carry[1509] , \add_42/carry[1508] ,
         \add_42/carry[1507] , \add_42/carry[1506] , \add_42/carry[1505] ,
         \add_42/carry[1504] , \add_42/carry[1503] , \add_42/carry[1502] ,
         \add_42/carry[1501] , \add_42/carry[1500] , \add_42/carry[1499] ,
         \add_42/carry[1498] , \add_42/carry[1497] , \add_42/carry[1496] ,
         \add_42/carry[1495] , \add_42/carry[1494] , \add_42/carry[1493] ,
         \add_42/carry[1492] , \add_42/carry[1491] , \add_42/carry[1490] ,
         \add_42/carry[1489] , \add_42/carry[1488] , \add_42/carry[1487] ,
         \add_42/carry[1486] , \add_42/carry[1485] , \add_42/carry[1484] ,
         \add_42/carry[1483] , \add_42/carry[1482] , \add_42/carry[1481] ,
         \add_42/carry[1480] , \add_42/carry[1479] , \add_42/carry[1478] ,
         \add_42/carry[1477] , \add_42/carry[1476] , \add_42/carry[1475] ,
         \add_42/carry[1474] , \add_42/carry[1473] , \add_42/carry[1472] ,
         \add_42/carry[1471] , \add_42/carry[1470] , \add_42/carry[1469] ,
         \add_42/carry[1468] , \add_42/carry[1467] , \add_42/carry[1466] ,
         \add_42/carry[1465] , \add_42/carry[1464] , \add_42/carry[1463] ,
         \add_42/carry[1462] , \add_42/carry[1461] , \add_42/carry[1460] ,
         \add_42/carry[1459] , \add_42/carry[1458] , \add_42/carry[1457] ,
         \add_42/carry[1456] , \add_42/carry[1455] , \add_42/carry[1454] ,
         \add_42/carry[1453] , \add_42/carry[1452] , \add_42/carry[1451] ,
         \add_42/carry[1450] , \add_42/carry[1449] , \add_42/carry[1448] ,
         \add_42/carry[1447] , \add_42/carry[1446] , \add_42/carry[1445] ,
         \add_42/carry[1444] , \add_42/carry[1443] , \add_42/carry[1442] ,
         \add_42/carry[1441] , \add_42/carry[1440] , \add_42/carry[1439] ,
         \add_42/carry[1438] , \add_42/carry[1437] , \add_42/carry[1436] ,
         \add_42/carry[1435] , \add_42/carry[1434] , \add_42/carry[1433] ,
         \add_42/carry[1432] , \add_42/carry[1431] , \add_42/carry[1430] ,
         \add_42/carry[1429] , \add_42/carry[1428] , \add_42/carry[1427] ,
         \add_42/carry[1426] , \add_42/carry[1425] , \add_42/carry[1424] ,
         \add_42/carry[1423] , \add_42/carry[1422] , \add_42/carry[1421] ,
         \add_42/carry[1420] , \add_42/carry[1419] , \add_42/carry[1418] ,
         \add_42/carry[1417] , \add_42/carry[1416] , \add_42/carry[1415] ,
         \add_42/carry[1414] , \add_42/carry[1413] , \add_42/carry[1412] ,
         \add_42/carry[1411] , \add_42/carry[1410] , \add_42/carry[1409] ,
         \add_42/carry[1408] , \add_42/carry[1407] , \add_42/carry[1406] ,
         \add_42/carry[1405] , \add_42/carry[1404] , \add_42/carry[1403] ,
         \add_42/carry[1402] , \add_42/carry[1401] , \add_42/carry[1400] ,
         \add_42/carry[1399] , \add_42/carry[1398] , \add_42/carry[1397] ,
         \add_42/carry[1396] , \add_42/carry[1395] , \add_42/carry[1394] ,
         \add_42/carry[1393] , \add_42/carry[1392] , \add_42/carry[1391] ,
         \add_42/carry[1390] , \add_42/carry[1389] , \add_42/carry[1388] ,
         \add_42/carry[1387] , \add_42/carry[1386] , \add_42/carry[1385] ,
         \add_42/carry[1384] , \add_42/carry[1383] , \add_42/carry[1382] ,
         \add_42/carry[1381] , \add_42/carry[1380] , \add_42/carry[1379] ,
         \add_42/carry[1378] , \add_42/carry[1377] , \add_42/carry[1376] ,
         \add_42/carry[1375] , \add_42/carry[1374] , \add_42/carry[1373] ,
         \add_42/carry[1372] , \add_42/carry[1371] , \add_42/carry[1370] ,
         \add_42/carry[1369] , \add_42/carry[1368] , \add_42/carry[1367] ,
         \add_42/carry[1366] , \add_42/carry[1365] , \add_42/carry[1364] ,
         \add_42/carry[1363] , \add_42/carry[1362] , \add_42/carry[1361] ,
         \add_42/carry[1360] , \add_42/carry[1359] , \add_42/carry[1358] ,
         \add_42/carry[1357] , \add_42/carry[1356] , \add_42/carry[1355] ,
         \add_42/carry[1354] , \add_42/carry[1353] , \add_42/carry[1352] ,
         \add_42/carry[1351] , \add_42/carry[1350] , \add_42/carry[1349] ,
         \add_42/carry[1348] , \add_42/carry[1347] , \add_42/carry[1346] ,
         \add_42/carry[1345] , \add_42/carry[1344] , \add_42/carry[1343] ,
         \add_42/carry[1342] , \add_42/carry[1341] , \add_42/carry[1340] ,
         \add_42/carry[1339] , \add_42/carry[1338] , \add_42/carry[1337] ,
         \add_42/carry[1336] , \add_42/carry[1335] , \add_42/carry[1334] ,
         \add_42/carry[1333] , \add_42/carry[1332] , \add_42/carry[1331] ,
         \add_42/carry[1330] , \add_42/carry[1329] , \add_42/carry[1328] ,
         \add_42/carry[1327] , \add_42/carry[1326] , \add_42/carry[1325] ,
         \add_42/carry[1324] , \add_42/carry[1323] , \add_42/carry[1322] ,
         \add_42/carry[1321] , \add_42/carry[1320] , \add_42/carry[1319] ,
         \add_42/carry[1318] , \add_42/carry[1317] , \add_42/carry[1316] ,
         \add_42/carry[1315] , \add_42/carry[1314] , \add_42/carry[1313] ,
         \add_42/carry[1312] , \add_42/carry[1311] , \add_42/carry[1310] ,
         \add_42/carry[1309] , \add_42/carry[1308] , \add_42/carry[1307] ,
         \add_42/carry[1306] , \add_42/carry[1305] , \add_42/carry[1304] ,
         \add_42/carry[1303] , \add_42/carry[1302] , \add_42/carry[1301] ,
         \add_42/carry[1300] , \add_42/carry[1299] , \add_42/carry[1298] ,
         \add_42/carry[1297] , \add_42/carry[1296] , \add_42/carry[1295] ,
         \add_42/carry[1294] , \add_42/carry[1293] , \add_42/carry[1292] ,
         \add_42/carry[1291] , \add_42/carry[1290] , \add_42/carry[1289] ,
         \add_42/carry[1288] , \add_42/carry[1287] , \add_42/carry[1286] ,
         \add_42/carry[1285] , \add_42/carry[1284] , \add_42/carry[1283] ,
         \add_42/carry[1282] , \add_42/carry[1281] , \add_42/carry[1280] ,
         \add_42/carry[1279] , \add_42/carry[1278] , \add_42/carry[1277] ,
         \add_42/carry[1276] , \add_42/carry[1275] , \add_42/carry[1274] ,
         \add_42/carry[1273] , \add_42/carry[1272] , \add_42/carry[1271] ,
         \add_42/carry[1270] , \add_42/carry[1269] , \add_42/carry[1268] ,
         \add_42/carry[1267] , \add_42/carry[1266] , \add_42/carry[1265] ,
         \add_42/carry[1264] , \add_42/carry[1263] , \add_42/carry[1262] ,
         \add_42/carry[1261] , \add_42/carry[1260] , \add_42/carry[1259] ,
         \add_42/carry[1258] , \add_42/carry[1257] , \add_42/carry[1256] ,
         \add_42/carry[1255] , \add_42/carry[1254] , \add_42/carry[1253] ,
         \add_42/carry[1252] , \add_42/carry[1251] , \add_42/carry[1250] ,
         \add_42/carry[1249] , \add_42/carry[1248] , \add_42/carry[1247] ,
         \add_42/carry[1246] , \add_42/carry[1245] , \add_42/carry[1244] ,
         \add_42/carry[1243] , \add_42/carry[1242] , \add_42/carry[1241] ,
         \add_42/carry[1240] , \add_42/carry[1239] , \add_42/carry[1238] ,
         \add_42/carry[1237] , \add_42/carry[1236] , \add_42/carry[1235] ,
         \add_42/carry[1234] , \add_42/carry[1233] , \add_42/carry[1232] ,
         \add_42/carry[1231] , \add_42/carry[1230] , \add_42/carry[1229] ,
         \add_42/carry[1228] , \add_42/carry[1227] , \add_42/carry[1226] ,
         \add_42/carry[1225] , \add_42/carry[1224] , \add_42/carry[1223] ,
         \add_42/carry[1222] , \add_42/carry[1221] , \add_42/carry[1220] ,
         \add_42/carry[1219] , \add_42/carry[1218] , \add_42/carry[1217] ,
         \add_42/carry[1216] , \add_42/carry[1215] , \add_42/carry[1214] ,
         \add_42/carry[1213] , \add_42/carry[1212] , \add_42/carry[1211] ,
         \add_42/carry[1210] , \add_42/carry[1209] , \add_42/carry[1208] ,
         \add_42/carry[1207] , \add_42/carry[1206] , \add_42/carry[1205] ,
         \add_42/carry[1204] , \add_42/carry[1203] , \add_42/carry[1202] ,
         \add_42/carry[1201] , \add_42/carry[1200] , \add_42/carry[1199] ,
         \add_42/carry[1198] , \add_42/carry[1197] , \add_42/carry[1196] ,
         \add_42/carry[1195] , \add_42/carry[1194] , \add_42/carry[1193] ,
         \add_42/carry[1192] , \add_42/carry[1191] , \add_42/carry[1190] ,
         \add_42/carry[1189] , \add_42/carry[1188] , \add_42/carry[1187] ,
         \add_42/carry[1186] , \add_42/carry[1185] , \add_42/carry[1184] ,
         \add_42/carry[1183] , \add_42/carry[1182] , \add_42/carry[1181] ,
         \add_42/carry[1180] , \add_42/carry[1179] , \add_42/carry[1178] ,
         \add_42/carry[1177] , \add_42/carry[1176] , \add_42/carry[1175] ,
         \add_42/carry[1174] , \add_42/carry[1173] , \add_42/carry[1172] ,
         \add_42/carry[1171] , \add_42/carry[1170] , \add_42/carry[1169] ,
         \add_42/carry[1168] , \add_42/carry[1167] , \add_42/carry[1166] ,
         \add_42/carry[1165] , \add_42/carry[1164] , \add_42/carry[1163] ,
         \add_42/carry[1162] , \add_42/carry[1161] , \add_42/carry[1160] ,
         \add_42/carry[1159] , \add_42/carry[1158] , \add_42/carry[1157] ,
         \add_42/carry[1156] , \add_42/carry[1155] , \add_42/carry[1154] ,
         \add_42/carry[1153] , \add_42/carry[1152] , \add_42/carry[1151] ,
         \add_42/carry[1150] , \add_42/carry[1149] , \add_42/carry[1148] ,
         \add_42/carry[1147] , \add_42/carry[1146] , \add_42/carry[1145] ,
         \add_42/carry[1144] , \add_42/carry[1143] , \add_42/carry[1142] ,
         \add_42/carry[1141] , \add_42/carry[1140] , \add_42/carry[1139] ,
         \add_42/carry[1138] , \add_42/carry[1137] , \add_42/carry[1136] ,
         \add_42/carry[1135] , \add_42/carry[1134] , \add_42/carry[1133] ,
         \add_42/carry[1132] , \add_42/carry[1131] , \add_42/carry[1130] ,
         \add_42/carry[1129] , \add_42/carry[1128] , \add_42/carry[1127] ,
         \add_42/carry[1126] , \add_42/carry[1125] , \add_42/carry[1124] ,
         \add_42/carry[1123] , \add_42/carry[1122] , \add_42/carry[1121] ,
         \add_42/carry[1120] , \add_42/carry[1119] , \add_42/carry[1118] ,
         \add_42/carry[1117] , \add_42/carry[1116] , \add_42/carry[1115] ,
         \add_42/carry[1114] , \add_42/carry[1113] , \add_42/carry[1112] ,
         \add_42/carry[1111] , \add_42/carry[1110] , \add_42/carry[1109] ,
         \add_42/carry[1108] , \add_42/carry[1107] , \add_42/carry[1106] ,
         \add_42/carry[1105] , \add_42/carry[1104] , \add_42/carry[1103] ,
         \add_42/carry[1102] , \add_42/carry[1101] , \add_42/carry[1100] ,
         \add_42/carry[1099] , \add_42/carry[1098] , \add_42/carry[1097] ,
         \add_42/carry[1096] , \add_42/carry[1095] , \add_42/carry[1094] ,
         \add_42/carry[1093] , \add_42/carry[1092] , \add_42/carry[1091] ,
         \add_42/carry[1090] , \add_42/carry[1089] , \add_42/carry[1088] ,
         \add_42/carry[1087] , \add_42/carry[1086] , \add_42/carry[1085] ,
         \add_42/carry[1084] , \add_42/carry[1083] , \add_42/carry[1082] ,
         \add_42/carry[1081] , \add_42/carry[1080] , \add_42/carry[1079] ,
         \add_42/carry[1078] , \add_42/carry[1077] , \add_42/carry[1076] ,
         \add_42/carry[1075] , \add_42/carry[1074] , \add_42/carry[1073] ,
         \add_42/carry[1072] , \add_42/carry[1071] , \add_42/carry[1070] ,
         \add_42/carry[1069] , \add_42/carry[1068] , \add_42/carry[1067] ,
         \add_42/carry[1066] , \add_42/carry[1065] , \add_42/carry[1064] ,
         \add_42/carry[1063] , \add_42/carry[1062] , \add_42/carry[1061] ,
         \add_42/carry[1060] , \add_42/carry[1059] , \add_42/carry[1058] ,
         \add_42/carry[1057] , \add_42/carry[1056] , \add_42/carry[1055] ,
         \add_42/carry[1054] , \add_42/carry[1053] , \add_42/carry[1052] ,
         \add_42/carry[1051] , \add_42/carry[1050] , \add_42/carry[1049] ,
         \add_42/carry[1048] , \add_42/carry[1047] , \add_42/carry[1046] ,
         \add_42/carry[1045] , \add_42/carry[1044] , \add_42/carry[1043] ,
         \add_42/carry[1042] , \add_42/carry[1041] , \add_42/carry[1040] ,
         \add_42/carry[1039] , \add_42/carry[1038] , \add_42/carry[1037] ,
         \add_42/carry[1036] , \add_42/carry[1035] , \add_42/carry[1034] ,
         \add_42/carry[1033] , \add_42/carry[1032] , \add_42/carry[1031] ,
         \add_42/carry[1030] , \add_42/carry[1029] , \add_42/carry[1028] ,
         \add_42/carry[1027] , \add_42/carry[1026] , \add_42/carry[1025] ,
         \add_42/carry[1024] , n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073;
  wire   [2047:0] sreg;
  assign o[1022] = sreg[1022];
  assign o[1021] = sreg[1021];
  assign o[1020] = sreg[1020];
  assign o[1019] = sreg[1019];
  assign o[1018] = sreg[1018];
  assign o[1017] = sreg[1017];
  assign o[1016] = sreg[1016];
  assign o[1015] = sreg[1015];
  assign o[1014] = sreg[1014];
  assign o[1013] = sreg[1013];
  assign o[1012] = sreg[1012];
  assign o[1011] = sreg[1011];
  assign o[1010] = sreg[1010];
  assign o[1009] = sreg[1009];
  assign o[1008] = sreg[1008];
  assign o[1007] = sreg[1007];
  assign o[1006] = sreg[1006];
  assign o[1005] = sreg[1005];
  assign o[1004] = sreg[1004];
  assign o[1003] = sreg[1003];
  assign o[1002] = sreg[1002];
  assign o[1001] = sreg[1001];
  assign o[1000] = sreg[1000];
  assign o[999] = sreg[999];
  assign o[998] = sreg[998];
  assign o[997] = sreg[997];
  assign o[996] = sreg[996];
  assign o[995] = sreg[995];
  assign o[994] = sreg[994];
  assign o[993] = sreg[993];
  assign o[992] = sreg[992];
  assign o[991] = sreg[991];
  assign o[990] = sreg[990];
  assign o[989] = sreg[989];
  assign o[988] = sreg[988];
  assign o[987] = sreg[987];
  assign o[986] = sreg[986];
  assign o[985] = sreg[985];
  assign o[984] = sreg[984];
  assign o[983] = sreg[983];
  assign o[982] = sreg[982];
  assign o[981] = sreg[981];
  assign o[980] = sreg[980];
  assign o[979] = sreg[979];
  assign o[978] = sreg[978];
  assign o[977] = sreg[977];
  assign o[976] = sreg[976];
  assign o[975] = sreg[975];
  assign o[974] = sreg[974];
  assign o[973] = sreg[973];
  assign o[972] = sreg[972];
  assign o[971] = sreg[971];
  assign o[970] = sreg[970];
  assign o[969] = sreg[969];
  assign o[968] = sreg[968];
  assign o[967] = sreg[967];
  assign o[966] = sreg[966];
  assign o[965] = sreg[965];
  assign o[964] = sreg[964];
  assign o[963] = sreg[963];
  assign o[962] = sreg[962];
  assign o[961] = sreg[961];
  assign o[960] = sreg[960];
  assign o[959] = sreg[959];
  assign o[958] = sreg[958];
  assign o[957] = sreg[957];
  assign o[956] = sreg[956];
  assign o[955] = sreg[955];
  assign o[954] = sreg[954];
  assign o[953] = sreg[953];
  assign o[952] = sreg[952];
  assign o[951] = sreg[951];
  assign o[950] = sreg[950];
  assign o[949] = sreg[949];
  assign o[948] = sreg[948];
  assign o[947] = sreg[947];
  assign o[946] = sreg[946];
  assign o[945] = sreg[945];
  assign o[944] = sreg[944];
  assign o[943] = sreg[943];
  assign o[942] = sreg[942];
  assign o[941] = sreg[941];
  assign o[940] = sreg[940];
  assign o[939] = sreg[939];
  assign o[938] = sreg[938];
  assign o[937] = sreg[937];
  assign o[936] = sreg[936];
  assign o[935] = sreg[935];
  assign o[934] = sreg[934];
  assign o[933] = sreg[933];
  assign o[932] = sreg[932];
  assign o[931] = sreg[931];
  assign o[930] = sreg[930];
  assign o[929] = sreg[929];
  assign o[928] = sreg[928];
  assign o[927] = sreg[927];
  assign o[926] = sreg[926];
  assign o[925] = sreg[925];
  assign o[924] = sreg[924];
  assign o[923] = sreg[923];
  assign o[922] = sreg[922];
  assign o[921] = sreg[921];
  assign o[920] = sreg[920];
  assign o[919] = sreg[919];
  assign o[918] = sreg[918];
  assign o[917] = sreg[917];
  assign o[916] = sreg[916];
  assign o[915] = sreg[915];
  assign o[914] = sreg[914];
  assign o[913] = sreg[913];
  assign o[912] = sreg[912];
  assign o[911] = sreg[911];
  assign o[910] = sreg[910];
  assign o[909] = sreg[909];
  assign o[908] = sreg[908];
  assign o[907] = sreg[907];
  assign o[906] = sreg[906];
  assign o[905] = sreg[905];
  assign o[904] = sreg[904];
  assign o[903] = sreg[903];
  assign o[902] = sreg[902];
  assign o[901] = sreg[901];
  assign o[900] = sreg[900];
  assign o[899] = sreg[899];
  assign o[898] = sreg[898];
  assign o[897] = sreg[897];
  assign o[896] = sreg[896];
  assign o[895] = sreg[895];
  assign o[894] = sreg[894];
  assign o[893] = sreg[893];
  assign o[892] = sreg[892];
  assign o[891] = sreg[891];
  assign o[890] = sreg[890];
  assign o[889] = sreg[889];
  assign o[888] = sreg[888];
  assign o[887] = sreg[887];
  assign o[886] = sreg[886];
  assign o[885] = sreg[885];
  assign o[884] = sreg[884];
  assign o[883] = sreg[883];
  assign o[882] = sreg[882];
  assign o[881] = sreg[881];
  assign o[880] = sreg[880];
  assign o[879] = sreg[879];
  assign o[878] = sreg[878];
  assign o[877] = sreg[877];
  assign o[876] = sreg[876];
  assign o[875] = sreg[875];
  assign o[874] = sreg[874];
  assign o[873] = sreg[873];
  assign o[872] = sreg[872];
  assign o[871] = sreg[871];
  assign o[870] = sreg[870];
  assign o[869] = sreg[869];
  assign o[868] = sreg[868];
  assign o[867] = sreg[867];
  assign o[866] = sreg[866];
  assign o[865] = sreg[865];
  assign o[864] = sreg[864];
  assign o[863] = sreg[863];
  assign o[862] = sreg[862];
  assign o[861] = sreg[861];
  assign o[860] = sreg[860];
  assign o[859] = sreg[859];
  assign o[858] = sreg[858];
  assign o[857] = sreg[857];
  assign o[856] = sreg[856];
  assign o[855] = sreg[855];
  assign o[854] = sreg[854];
  assign o[853] = sreg[853];
  assign o[852] = sreg[852];
  assign o[851] = sreg[851];
  assign o[850] = sreg[850];
  assign o[849] = sreg[849];
  assign o[848] = sreg[848];
  assign o[847] = sreg[847];
  assign o[846] = sreg[846];
  assign o[845] = sreg[845];
  assign o[844] = sreg[844];
  assign o[843] = sreg[843];
  assign o[842] = sreg[842];
  assign o[841] = sreg[841];
  assign o[840] = sreg[840];
  assign o[839] = sreg[839];
  assign o[838] = sreg[838];
  assign o[837] = sreg[837];
  assign o[836] = sreg[836];
  assign o[835] = sreg[835];
  assign o[834] = sreg[834];
  assign o[833] = sreg[833];
  assign o[832] = sreg[832];
  assign o[831] = sreg[831];
  assign o[830] = sreg[830];
  assign o[829] = sreg[829];
  assign o[828] = sreg[828];
  assign o[827] = sreg[827];
  assign o[826] = sreg[826];
  assign o[825] = sreg[825];
  assign o[824] = sreg[824];
  assign o[823] = sreg[823];
  assign o[822] = sreg[822];
  assign o[821] = sreg[821];
  assign o[820] = sreg[820];
  assign o[819] = sreg[819];
  assign o[818] = sreg[818];
  assign o[817] = sreg[817];
  assign o[816] = sreg[816];
  assign o[815] = sreg[815];
  assign o[814] = sreg[814];
  assign o[813] = sreg[813];
  assign o[812] = sreg[812];
  assign o[811] = sreg[811];
  assign o[810] = sreg[810];
  assign o[809] = sreg[809];
  assign o[808] = sreg[808];
  assign o[807] = sreg[807];
  assign o[806] = sreg[806];
  assign o[805] = sreg[805];
  assign o[804] = sreg[804];
  assign o[803] = sreg[803];
  assign o[802] = sreg[802];
  assign o[801] = sreg[801];
  assign o[800] = sreg[800];
  assign o[799] = sreg[799];
  assign o[798] = sreg[798];
  assign o[797] = sreg[797];
  assign o[796] = sreg[796];
  assign o[795] = sreg[795];
  assign o[794] = sreg[794];
  assign o[793] = sreg[793];
  assign o[792] = sreg[792];
  assign o[791] = sreg[791];
  assign o[790] = sreg[790];
  assign o[789] = sreg[789];
  assign o[788] = sreg[788];
  assign o[787] = sreg[787];
  assign o[786] = sreg[786];
  assign o[785] = sreg[785];
  assign o[784] = sreg[784];
  assign o[783] = sreg[783];
  assign o[782] = sreg[782];
  assign o[781] = sreg[781];
  assign o[780] = sreg[780];
  assign o[779] = sreg[779];
  assign o[778] = sreg[778];
  assign o[777] = sreg[777];
  assign o[776] = sreg[776];
  assign o[775] = sreg[775];
  assign o[774] = sreg[774];
  assign o[773] = sreg[773];
  assign o[772] = sreg[772];
  assign o[771] = sreg[771];
  assign o[770] = sreg[770];
  assign o[769] = sreg[769];
  assign o[768] = sreg[768];
  assign o[767] = sreg[767];
  assign o[766] = sreg[766];
  assign o[765] = sreg[765];
  assign o[764] = sreg[764];
  assign o[763] = sreg[763];
  assign o[762] = sreg[762];
  assign o[761] = sreg[761];
  assign o[760] = sreg[760];
  assign o[759] = sreg[759];
  assign o[758] = sreg[758];
  assign o[757] = sreg[757];
  assign o[756] = sreg[756];
  assign o[755] = sreg[755];
  assign o[754] = sreg[754];
  assign o[753] = sreg[753];
  assign o[752] = sreg[752];
  assign o[751] = sreg[751];
  assign o[750] = sreg[750];
  assign o[749] = sreg[749];
  assign o[748] = sreg[748];
  assign o[747] = sreg[747];
  assign o[746] = sreg[746];
  assign o[745] = sreg[745];
  assign o[744] = sreg[744];
  assign o[743] = sreg[743];
  assign o[742] = sreg[742];
  assign o[741] = sreg[741];
  assign o[740] = sreg[740];
  assign o[739] = sreg[739];
  assign o[738] = sreg[738];
  assign o[737] = sreg[737];
  assign o[736] = sreg[736];
  assign o[735] = sreg[735];
  assign o[734] = sreg[734];
  assign o[733] = sreg[733];
  assign o[732] = sreg[732];
  assign o[731] = sreg[731];
  assign o[730] = sreg[730];
  assign o[729] = sreg[729];
  assign o[728] = sreg[728];
  assign o[727] = sreg[727];
  assign o[726] = sreg[726];
  assign o[725] = sreg[725];
  assign o[724] = sreg[724];
  assign o[723] = sreg[723];
  assign o[722] = sreg[722];
  assign o[721] = sreg[721];
  assign o[720] = sreg[720];
  assign o[719] = sreg[719];
  assign o[718] = sreg[718];
  assign o[717] = sreg[717];
  assign o[716] = sreg[716];
  assign o[715] = sreg[715];
  assign o[714] = sreg[714];
  assign o[713] = sreg[713];
  assign o[712] = sreg[712];
  assign o[711] = sreg[711];
  assign o[710] = sreg[710];
  assign o[709] = sreg[709];
  assign o[708] = sreg[708];
  assign o[707] = sreg[707];
  assign o[706] = sreg[706];
  assign o[705] = sreg[705];
  assign o[704] = sreg[704];
  assign o[703] = sreg[703];
  assign o[702] = sreg[702];
  assign o[701] = sreg[701];
  assign o[700] = sreg[700];
  assign o[699] = sreg[699];
  assign o[698] = sreg[698];
  assign o[697] = sreg[697];
  assign o[696] = sreg[696];
  assign o[695] = sreg[695];
  assign o[694] = sreg[694];
  assign o[693] = sreg[693];
  assign o[692] = sreg[692];
  assign o[691] = sreg[691];
  assign o[690] = sreg[690];
  assign o[689] = sreg[689];
  assign o[688] = sreg[688];
  assign o[687] = sreg[687];
  assign o[686] = sreg[686];
  assign o[685] = sreg[685];
  assign o[684] = sreg[684];
  assign o[683] = sreg[683];
  assign o[682] = sreg[682];
  assign o[681] = sreg[681];
  assign o[680] = sreg[680];
  assign o[679] = sreg[679];
  assign o[678] = sreg[678];
  assign o[677] = sreg[677];
  assign o[676] = sreg[676];
  assign o[675] = sreg[675];
  assign o[674] = sreg[674];
  assign o[673] = sreg[673];
  assign o[672] = sreg[672];
  assign o[671] = sreg[671];
  assign o[670] = sreg[670];
  assign o[669] = sreg[669];
  assign o[668] = sreg[668];
  assign o[667] = sreg[667];
  assign o[666] = sreg[666];
  assign o[665] = sreg[665];
  assign o[664] = sreg[664];
  assign o[663] = sreg[663];
  assign o[662] = sreg[662];
  assign o[661] = sreg[661];
  assign o[660] = sreg[660];
  assign o[659] = sreg[659];
  assign o[658] = sreg[658];
  assign o[657] = sreg[657];
  assign o[656] = sreg[656];
  assign o[655] = sreg[655];
  assign o[654] = sreg[654];
  assign o[653] = sreg[653];
  assign o[652] = sreg[652];
  assign o[651] = sreg[651];
  assign o[650] = sreg[650];
  assign o[649] = sreg[649];
  assign o[648] = sreg[648];
  assign o[647] = sreg[647];
  assign o[646] = sreg[646];
  assign o[645] = sreg[645];
  assign o[644] = sreg[644];
  assign o[643] = sreg[643];
  assign o[642] = sreg[642];
  assign o[641] = sreg[641];
  assign o[640] = sreg[640];
  assign o[639] = sreg[639];
  assign o[638] = sreg[638];
  assign o[637] = sreg[637];
  assign o[636] = sreg[636];
  assign o[635] = sreg[635];
  assign o[634] = sreg[634];
  assign o[633] = sreg[633];
  assign o[632] = sreg[632];
  assign o[631] = sreg[631];
  assign o[630] = sreg[630];
  assign o[629] = sreg[629];
  assign o[628] = sreg[628];
  assign o[627] = sreg[627];
  assign o[626] = sreg[626];
  assign o[625] = sreg[625];
  assign o[624] = sreg[624];
  assign o[623] = sreg[623];
  assign o[622] = sreg[622];
  assign o[621] = sreg[621];
  assign o[620] = sreg[620];
  assign o[619] = sreg[619];
  assign o[618] = sreg[618];
  assign o[617] = sreg[617];
  assign o[616] = sreg[616];
  assign o[615] = sreg[615];
  assign o[614] = sreg[614];
  assign o[613] = sreg[613];
  assign o[612] = sreg[612];
  assign o[611] = sreg[611];
  assign o[610] = sreg[610];
  assign o[609] = sreg[609];
  assign o[608] = sreg[608];
  assign o[607] = sreg[607];
  assign o[606] = sreg[606];
  assign o[605] = sreg[605];
  assign o[604] = sreg[604];
  assign o[603] = sreg[603];
  assign o[602] = sreg[602];
  assign o[601] = sreg[601];
  assign o[600] = sreg[600];
  assign o[599] = sreg[599];
  assign o[598] = sreg[598];
  assign o[597] = sreg[597];
  assign o[596] = sreg[596];
  assign o[595] = sreg[595];
  assign o[594] = sreg[594];
  assign o[593] = sreg[593];
  assign o[592] = sreg[592];
  assign o[591] = sreg[591];
  assign o[590] = sreg[590];
  assign o[589] = sreg[589];
  assign o[588] = sreg[588];
  assign o[587] = sreg[587];
  assign o[586] = sreg[586];
  assign o[585] = sreg[585];
  assign o[584] = sreg[584];
  assign o[583] = sreg[583];
  assign o[582] = sreg[582];
  assign o[581] = sreg[581];
  assign o[580] = sreg[580];
  assign o[579] = sreg[579];
  assign o[578] = sreg[578];
  assign o[577] = sreg[577];
  assign o[576] = sreg[576];
  assign o[575] = sreg[575];
  assign o[574] = sreg[574];
  assign o[573] = sreg[573];
  assign o[572] = sreg[572];
  assign o[571] = sreg[571];
  assign o[570] = sreg[570];
  assign o[569] = sreg[569];
  assign o[568] = sreg[568];
  assign o[567] = sreg[567];
  assign o[566] = sreg[566];
  assign o[565] = sreg[565];
  assign o[564] = sreg[564];
  assign o[563] = sreg[563];
  assign o[562] = sreg[562];
  assign o[561] = sreg[561];
  assign o[560] = sreg[560];
  assign o[559] = sreg[559];
  assign o[558] = sreg[558];
  assign o[557] = sreg[557];
  assign o[556] = sreg[556];
  assign o[555] = sreg[555];
  assign o[554] = sreg[554];
  assign o[553] = sreg[553];
  assign o[552] = sreg[552];
  assign o[551] = sreg[551];
  assign o[550] = sreg[550];
  assign o[549] = sreg[549];
  assign o[548] = sreg[548];
  assign o[547] = sreg[547];
  assign o[546] = sreg[546];
  assign o[545] = sreg[545];
  assign o[544] = sreg[544];
  assign o[543] = sreg[543];
  assign o[542] = sreg[542];
  assign o[541] = sreg[541];
  assign o[540] = sreg[540];
  assign o[539] = sreg[539];
  assign o[538] = sreg[538];
  assign o[537] = sreg[537];
  assign o[536] = sreg[536];
  assign o[535] = sreg[535];
  assign o[534] = sreg[534];
  assign o[533] = sreg[533];
  assign o[532] = sreg[532];
  assign o[531] = sreg[531];
  assign o[530] = sreg[530];
  assign o[529] = sreg[529];
  assign o[528] = sreg[528];
  assign o[527] = sreg[527];
  assign o[526] = sreg[526];
  assign o[525] = sreg[525];
  assign o[524] = sreg[524];
  assign o[523] = sreg[523];
  assign o[522] = sreg[522];
  assign o[521] = sreg[521];
  assign o[520] = sreg[520];
  assign o[519] = sreg[519];
  assign o[518] = sreg[518];
  assign o[517] = sreg[517];
  assign o[516] = sreg[516];
  assign o[515] = sreg[515];
  assign o[514] = sreg[514];
  assign o[513] = sreg[513];
  assign o[512] = sreg[512];
  assign o[511] = sreg[511];
  assign o[510] = sreg[510];
  assign o[509] = sreg[509];
  assign o[508] = sreg[508];
  assign o[507] = sreg[507];
  assign o[506] = sreg[506];
  assign o[505] = sreg[505];
  assign o[504] = sreg[504];
  assign o[503] = sreg[503];
  assign o[502] = sreg[502];
  assign o[501] = sreg[501];
  assign o[500] = sreg[500];
  assign o[499] = sreg[499];
  assign o[498] = sreg[498];
  assign o[497] = sreg[497];
  assign o[496] = sreg[496];
  assign o[495] = sreg[495];
  assign o[494] = sreg[494];
  assign o[493] = sreg[493];
  assign o[492] = sreg[492];
  assign o[491] = sreg[491];
  assign o[490] = sreg[490];
  assign o[489] = sreg[489];
  assign o[488] = sreg[488];
  assign o[487] = sreg[487];
  assign o[486] = sreg[486];
  assign o[485] = sreg[485];
  assign o[484] = sreg[484];
  assign o[483] = sreg[483];
  assign o[482] = sreg[482];
  assign o[481] = sreg[481];
  assign o[480] = sreg[480];
  assign o[479] = sreg[479];
  assign o[478] = sreg[478];
  assign o[477] = sreg[477];
  assign o[476] = sreg[476];
  assign o[475] = sreg[475];
  assign o[474] = sreg[474];
  assign o[473] = sreg[473];
  assign o[472] = sreg[472];
  assign o[471] = sreg[471];
  assign o[470] = sreg[470];
  assign o[469] = sreg[469];
  assign o[468] = sreg[468];
  assign o[467] = sreg[467];
  assign o[466] = sreg[466];
  assign o[465] = sreg[465];
  assign o[464] = sreg[464];
  assign o[463] = sreg[463];
  assign o[462] = sreg[462];
  assign o[461] = sreg[461];
  assign o[460] = sreg[460];
  assign o[459] = sreg[459];
  assign o[458] = sreg[458];
  assign o[457] = sreg[457];
  assign o[456] = sreg[456];
  assign o[455] = sreg[455];
  assign o[454] = sreg[454];
  assign o[453] = sreg[453];
  assign o[452] = sreg[452];
  assign o[451] = sreg[451];
  assign o[450] = sreg[450];
  assign o[449] = sreg[449];
  assign o[448] = sreg[448];
  assign o[447] = sreg[447];
  assign o[446] = sreg[446];
  assign o[445] = sreg[445];
  assign o[444] = sreg[444];
  assign o[443] = sreg[443];
  assign o[442] = sreg[442];
  assign o[441] = sreg[441];
  assign o[440] = sreg[440];
  assign o[439] = sreg[439];
  assign o[438] = sreg[438];
  assign o[437] = sreg[437];
  assign o[436] = sreg[436];
  assign o[435] = sreg[435];
  assign o[434] = sreg[434];
  assign o[433] = sreg[433];
  assign o[432] = sreg[432];
  assign o[431] = sreg[431];
  assign o[430] = sreg[430];
  assign o[429] = sreg[429];
  assign o[428] = sreg[428];
  assign o[427] = sreg[427];
  assign o[426] = sreg[426];
  assign o[425] = sreg[425];
  assign o[424] = sreg[424];
  assign o[423] = sreg[423];
  assign o[422] = sreg[422];
  assign o[421] = sreg[421];
  assign o[420] = sreg[420];
  assign o[419] = sreg[419];
  assign o[418] = sreg[418];
  assign o[417] = sreg[417];
  assign o[416] = sreg[416];
  assign o[415] = sreg[415];
  assign o[414] = sreg[414];
  assign o[413] = sreg[413];
  assign o[412] = sreg[412];
  assign o[411] = sreg[411];
  assign o[410] = sreg[410];
  assign o[409] = sreg[409];
  assign o[408] = sreg[408];
  assign o[407] = sreg[407];
  assign o[406] = sreg[406];
  assign o[405] = sreg[405];
  assign o[404] = sreg[404];
  assign o[403] = sreg[403];
  assign o[402] = sreg[402];
  assign o[401] = sreg[401];
  assign o[400] = sreg[400];
  assign o[399] = sreg[399];
  assign o[398] = sreg[398];
  assign o[397] = sreg[397];
  assign o[396] = sreg[396];
  assign o[395] = sreg[395];
  assign o[394] = sreg[394];
  assign o[393] = sreg[393];
  assign o[392] = sreg[392];
  assign o[391] = sreg[391];
  assign o[390] = sreg[390];
  assign o[389] = sreg[389];
  assign o[388] = sreg[388];
  assign o[387] = sreg[387];
  assign o[386] = sreg[386];
  assign o[385] = sreg[385];
  assign o[384] = sreg[384];
  assign o[383] = sreg[383];
  assign o[382] = sreg[382];
  assign o[381] = sreg[381];
  assign o[380] = sreg[380];
  assign o[379] = sreg[379];
  assign o[378] = sreg[378];
  assign o[377] = sreg[377];
  assign o[376] = sreg[376];
  assign o[375] = sreg[375];
  assign o[374] = sreg[374];
  assign o[373] = sreg[373];
  assign o[372] = sreg[372];
  assign o[371] = sreg[371];
  assign o[370] = sreg[370];
  assign o[369] = sreg[369];
  assign o[368] = sreg[368];
  assign o[367] = sreg[367];
  assign o[366] = sreg[366];
  assign o[365] = sreg[365];
  assign o[364] = sreg[364];
  assign o[363] = sreg[363];
  assign o[362] = sreg[362];
  assign o[361] = sreg[361];
  assign o[360] = sreg[360];
  assign o[359] = sreg[359];
  assign o[358] = sreg[358];
  assign o[357] = sreg[357];
  assign o[356] = sreg[356];
  assign o[355] = sreg[355];
  assign o[354] = sreg[354];
  assign o[353] = sreg[353];
  assign o[352] = sreg[352];
  assign o[351] = sreg[351];
  assign o[350] = sreg[350];
  assign o[349] = sreg[349];
  assign o[348] = sreg[348];
  assign o[347] = sreg[347];
  assign o[346] = sreg[346];
  assign o[345] = sreg[345];
  assign o[344] = sreg[344];
  assign o[343] = sreg[343];
  assign o[342] = sreg[342];
  assign o[341] = sreg[341];
  assign o[340] = sreg[340];
  assign o[339] = sreg[339];
  assign o[338] = sreg[338];
  assign o[337] = sreg[337];
  assign o[336] = sreg[336];
  assign o[335] = sreg[335];
  assign o[334] = sreg[334];
  assign o[333] = sreg[333];
  assign o[332] = sreg[332];
  assign o[331] = sreg[331];
  assign o[330] = sreg[330];
  assign o[329] = sreg[329];
  assign o[328] = sreg[328];
  assign o[327] = sreg[327];
  assign o[326] = sreg[326];
  assign o[325] = sreg[325];
  assign o[324] = sreg[324];
  assign o[323] = sreg[323];
  assign o[322] = sreg[322];
  assign o[321] = sreg[321];
  assign o[320] = sreg[320];
  assign o[319] = sreg[319];
  assign o[318] = sreg[318];
  assign o[317] = sreg[317];
  assign o[316] = sreg[316];
  assign o[315] = sreg[315];
  assign o[314] = sreg[314];
  assign o[313] = sreg[313];
  assign o[312] = sreg[312];
  assign o[311] = sreg[311];
  assign o[310] = sreg[310];
  assign o[309] = sreg[309];
  assign o[308] = sreg[308];
  assign o[307] = sreg[307];
  assign o[306] = sreg[306];
  assign o[305] = sreg[305];
  assign o[304] = sreg[304];
  assign o[303] = sreg[303];
  assign o[302] = sreg[302];
  assign o[301] = sreg[301];
  assign o[300] = sreg[300];
  assign o[299] = sreg[299];
  assign o[298] = sreg[298];
  assign o[297] = sreg[297];
  assign o[296] = sreg[296];
  assign o[295] = sreg[295];
  assign o[294] = sreg[294];
  assign o[293] = sreg[293];
  assign o[292] = sreg[292];
  assign o[291] = sreg[291];
  assign o[290] = sreg[290];
  assign o[289] = sreg[289];
  assign o[288] = sreg[288];
  assign o[287] = sreg[287];
  assign o[286] = sreg[286];
  assign o[285] = sreg[285];
  assign o[284] = sreg[284];
  assign o[283] = sreg[283];
  assign o[282] = sreg[282];
  assign o[281] = sreg[281];
  assign o[280] = sreg[280];
  assign o[279] = sreg[279];
  assign o[278] = sreg[278];
  assign o[277] = sreg[277];
  assign o[276] = sreg[276];
  assign o[275] = sreg[275];
  assign o[274] = sreg[274];
  assign o[273] = sreg[273];
  assign o[272] = sreg[272];
  assign o[271] = sreg[271];
  assign o[270] = sreg[270];
  assign o[269] = sreg[269];
  assign o[268] = sreg[268];
  assign o[267] = sreg[267];
  assign o[266] = sreg[266];
  assign o[265] = sreg[265];
  assign o[264] = sreg[264];
  assign o[263] = sreg[263];
  assign o[262] = sreg[262];
  assign o[261] = sreg[261];
  assign o[260] = sreg[260];
  assign o[259] = sreg[259];
  assign o[258] = sreg[258];
  assign o[257] = sreg[257];
  assign o[256] = sreg[256];
  assign o[255] = sreg[255];
  assign o[254] = sreg[254];
  assign o[253] = sreg[253];
  assign o[252] = sreg[252];
  assign o[251] = sreg[251];
  assign o[250] = sreg[250];
  assign o[249] = sreg[249];
  assign o[248] = sreg[248];
  assign o[247] = sreg[247];
  assign o[246] = sreg[246];
  assign o[245] = sreg[245];
  assign o[244] = sreg[244];
  assign o[243] = sreg[243];
  assign o[242] = sreg[242];
  assign o[241] = sreg[241];
  assign o[240] = sreg[240];
  assign o[239] = sreg[239];
  assign o[238] = sreg[238];
  assign o[237] = sreg[237];
  assign o[236] = sreg[236];
  assign o[235] = sreg[235];
  assign o[234] = sreg[234];
  assign o[233] = sreg[233];
  assign o[232] = sreg[232];
  assign o[231] = sreg[231];
  assign o[230] = sreg[230];
  assign o[229] = sreg[229];
  assign o[228] = sreg[228];
  assign o[227] = sreg[227];
  assign o[226] = sreg[226];
  assign o[225] = sreg[225];
  assign o[224] = sreg[224];
  assign o[223] = sreg[223];
  assign o[222] = sreg[222];
  assign o[221] = sreg[221];
  assign o[220] = sreg[220];
  assign o[219] = sreg[219];
  assign o[218] = sreg[218];
  assign o[217] = sreg[217];
  assign o[216] = sreg[216];
  assign o[215] = sreg[215];
  assign o[214] = sreg[214];
  assign o[213] = sreg[213];
  assign o[212] = sreg[212];
  assign o[211] = sreg[211];
  assign o[210] = sreg[210];
  assign o[209] = sreg[209];
  assign o[208] = sreg[208];
  assign o[207] = sreg[207];
  assign o[206] = sreg[206];
  assign o[205] = sreg[205];
  assign o[204] = sreg[204];
  assign o[203] = sreg[203];
  assign o[202] = sreg[202];
  assign o[201] = sreg[201];
  assign o[200] = sreg[200];
  assign o[199] = sreg[199];
  assign o[198] = sreg[198];
  assign o[197] = sreg[197];
  assign o[196] = sreg[196];
  assign o[195] = sreg[195];
  assign o[194] = sreg[194];
  assign o[193] = sreg[193];
  assign o[192] = sreg[192];
  assign o[191] = sreg[191];
  assign o[190] = sreg[190];
  assign o[189] = sreg[189];
  assign o[188] = sreg[188];
  assign o[187] = sreg[187];
  assign o[186] = sreg[186];
  assign o[185] = sreg[185];
  assign o[184] = sreg[184];
  assign o[183] = sreg[183];
  assign o[182] = sreg[182];
  assign o[181] = sreg[181];
  assign o[180] = sreg[180];
  assign o[179] = sreg[179];
  assign o[178] = sreg[178];
  assign o[177] = sreg[177];
  assign o[176] = sreg[176];
  assign o[175] = sreg[175];
  assign o[174] = sreg[174];
  assign o[173] = sreg[173];
  assign o[172] = sreg[172];
  assign o[171] = sreg[171];
  assign o[170] = sreg[170];
  assign o[169] = sreg[169];
  assign o[168] = sreg[168];
  assign o[167] = sreg[167];
  assign o[166] = sreg[166];
  assign o[165] = sreg[165];
  assign o[164] = sreg[164];
  assign o[163] = sreg[163];
  assign o[162] = sreg[162];
  assign o[161] = sreg[161];
  assign o[160] = sreg[160];
  assign o[159] = sreg[159];
  assign o[158] = sreg[158];
  assign o[157] = sreg[157];
  assign o[156] = sreg[156];
  assign o[155] = sreg[155];
  assign o[154] = sreg[154];
  assign o[153] = sreg[153];
  assign o[152] = sreg[152];
  assign o[151] = sreg[151];
  assign o[150] = sreg[150];
  assign o[149] = sreg[149];
  assign o[148] = sreg[148];
  assign o[147] = sreg[147];
  assign o[146] = sreg[146];
  assign o[145] = sreg[145];
  assign o[144] = sreg[144];
  assign o[143] = sreg[143];
  assign o[142] = sreg[142];
  assign o[141] = sreg[141];
  assign o[140] = sreg[140];
  assign o[139] = sreg[139];
  assign o[138] = sreg[138];
  assign o[137] = sreg[137];
  assign o[136] = sreg[136];
  assign o[135] = sreg[135];
  assign o[134] = sreg[134];
  assign o[133] = sreg[133];
  assign o[132] = sreg[132];
  assign o[131] = sreg[131];
  assign o[130] = sreg[130];
  assign o[129] = sreg[129];
  assign o[128] = sreg[128];
  assign o[127] = sreg[127];
  assign o[126] = sreg[126];
  assign o[125] = sreg[125];
  assign o[124] = sreg[124];
  assign o[123] = sreg[123];
  assign o[122] = sreg[122];
  assign o[121] = sreg[121];
  assign o[120] = sreg[120];
  assign o[119] = sreg[119];
  assign o[118] = sreg[118];
  assign o[117] = sreg[117];
  assign o[116] = sreg[116];
  assign o[115] = sreg[115];
  assign o[114] = sreg[114];
  assign o[113] = sreg[113];
  assign o[112] = sreg[112];
  assign o[111] = sreg[111];
  assign o[110] = sreg[110];
  assign o[109] = sreg[109];
  assign o[108] = sreg[108];
  assign o[107] = sreg[107];
  assign o[106] = sreg[106];
  assign o[105] = sreg[105];
  assign o[104] = sreg[104];
  assign o[103] = sreg[103];
  assign o[102] = sreg[102];
  assign o[101] = sreg[101];
  assign o[100] = sreg[100];
  assign o[99] = sreg[99];
  assign o[98] = sreg[98];
  assign o[97] = sreg[97];
  assign o[96] = sreg[96];
  assign o[95] = sreg[95];
  assign o[94] = sreg[94];
  assign o[93] = sreg[93];
  assign o[92] = sreg[92];
  assign o[91] = sreg[91];
  assign o[90] = sreg[90];
  assign o[89] = sreg[89];
  assign o[88] = sreg[88];
  assign o[87] = sreg[87];
  assign o[86] = sreg[86];
  assign o[85] = sreg[85];
  assign o[84] = sreg[84];
  assign o[83] = sreg[83];
  assign o[82] = sreg[82];
  assign o[81] = sreg[81];
  assign o[80] = sreg[80];
  assign o[79] = sreg[79];
  assign o[78] = sreg[78];
  assign o[77] = sreg[77];
  assign o[76] = sreg[76];
  assign o[75] = sreg[75];
  assign o[74] = sreg[74];
  assign o[73] = sreg[73];
  assign o[72] = sreg[72];
  assign o[71] = sreg[71];
  assign o[70] = sreg[70];
  assign o[69] = sreg[69];
  assign o[68] = sreg[68];
  assign o[67] = sreg[67];
  assign o[66] = sreg[66];
  assign o[65] = sreg[65];
  assign o[64] = sreg[64];
  assign o[63] = sreg[63];
  assign o[62] = sreg[62];
  assign o[61] = sreg[61];
  assign o[60] = sreg[60];
  assign o[59] = sreg[59];
  assign o[58] = sreg[58];
  assign o[57] = sreg[57];
  assign o[56] = sreg[56];
  assign o[55] = sreg[55];
  assign o[54] = sreg[54];
  assign o[53] = sreg[53];
  assign o[52] = sreg[52];
  assign o[51] = sreg[51];
  assign o[50] = sreg[50];
  assign o[49] = sreg[49];
  assign o[48] = sreg[48];
  assign o[47] = sreg[47];
  assign o[46] = sreg[46];
  assign o[45] = sreg[45];
  assign o[44] = sreg[44];
  assign o[43] = sreg[43];
  assign o[42] = sreg[42];
  assign o[41] = sreg[41];
  assign o[40] = sreg[40];
  assign o[39] = sreg[39];
  assign o[38] = sreg[38];
  assign o[37] = sreg[37];
  assign o[36] = sreg[36];
  assign o[35] = sreg[35];
  assign o[34] = sreg[34];
  assign o[33] = sreg[33];
  assign o[32] = sreg[32];
  assign o[31] = sreg[31];
  assign o[30] = sreg[30];
  assign o[29] = sreg[29];
  assign o[28] = sreg[28];
  assign o[27] = sreg[27];
  assign o[26] = sreg[26];
  assign o[25] = sreg[25];
  assign o[24] = sreg[24];
  assign o[23] = sreg[23];
  assign o[22] = sreg[22];
  assign o[21] = sreg[21];
  assign o[20] = sreg[20];
  assign o[19] = sreg[19];
  assign o[18] = sreg[18];
  assign o[17] = sreg[17];
  assign o[16] = sreg[16];
  assign o[15] = sreg[15];
  assign o[14] = sreg[14];
  assign o[13] = sreg[13];
  assign o[12] = sreg[12];
  assign o[11] = sreg[11];
  assign o[10] = sreg[10];
  assign o[9] = sreg[9];
  assign o[8] = sreg[8];
  assign o[7] = sreg[7];
  assign o[6] = sreg[6];
  assign o[5] = sreg[5];
  assign o[4] = sreg[4];
  assign o[3] = sreg[3];
  assign o[2] = sreg[2];
  assign o[1] = sreg[1];
  assign o[2047] = \add_42/carry[2047] ;

  DFF \sreg_reg[0]  ( .D(sreg[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[0]) );
  DFF \sreg_reg[1]  ( .D(sreg[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[1])
         );
  DFF \sreg_reg[2]  ( .D(sreg[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[2])
         );
  DFF \sreg_reg[3]  ( .D(sreg[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[3])
         );
  DFF \sreg_reg[4]  ( .D(sreg[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[4])
         );
  DFF \sreg_reg[5]  ( .D(sreg[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[5])
         );
  DFF \sreg_reg[6]  ( .D(sreg[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[6])
         );
  DFF \sreg_reg[7]  ( .D(sreg[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[7])
         );
  DFF \sreg_reg[8]  ( .D(sreg[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[8])
         );
  DFF \sreg_reg[9]  ( .D(sreg[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(sreg[9]) );
  DFF \sreg_reg[10]  ( .D(sreg[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[10]) );
  DFF \sreg_reg[11]  ( .D(sreg[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[11]) );
  DFF \sreg_reg[12]  ( .D(sreg[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[12]) );
  DFF \sreg_reg[13]  ( .D(sreg[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[13]) );
  DFF \sreg_reg[14]  ( .D(sreg[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[14]) );
  DFF \sreg_reg[15]  ( .D(sreg[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[15]) );
  DFF \sreg_reg[16]  ( .D(sreg[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[16]) );
  DFF \sreg_reg[17]  ( .D(sreg[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[17]) );
  DFF \sreg_reg[18]  ( .D(sreg[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[18]) );
  DFF \sreg_reg[19]  ( .D(sreg[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[19]) );
  DFF \sreg_reg[20]  ( .D(sreg[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[20]) );
  DFF \sreg_reg[21]  ( .D(sreg[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[21]) );
  DFF \sreg_reg[22]  ( .D(sreg[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[22]) );
  DFF \sreg_reg[23]  ( .D(sreg[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[23]) );
  DFF \sreg_reg[24]  ( .D(sreg[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[24]) );
  DFF \sreg_reg[25]  ( .D(sreg[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[25]) );
  DFF \sreg_reg[26]  ( .D(sreg[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[26]) );
  DFF \sreg_reg[27]  ( .D(sreg[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[27]) );
  DFF \sreg_reg[28]  ( .D(sreg[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[28]) );
  DFF \sreg_reg[29]  ( .D(sreg[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[29]) );
  DFF \sreg_reg[30]  ( .D(sreg[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[30]) );
  DFF \sreg_reg[31]  ( .D(sreg[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[31]) );
  DFF \sreg_reg[32]  ( .D(sreg[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[32]) );
  DFF \sreg_reg[33]  ( .D(sreg[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[33]) );
  DFF \sreg_reg[34]  ( .D(sreg[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[34]) );
  DFF \sreg_reg[35]  ( .D(sreg[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[35]) );
  DFF \sreg_reg[36]  ( .D(sreg[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[36]) );
  DFF \sreg_reg[37]  ( .D(sreg[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[37]) );
  DFF \sreg_reg[38]  ( .D(sreg[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[38]) );
  DFF \sreg_reg[39]  ( .D(sreg[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[39]) );
  DFF \sreg_reg[40]  ( .D(sreg[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[40]) );
  DFF \sreg_reg[41]  ( .D(sreg[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[41]) );
  DFF \sreg_reg[42]  ( .D(sreg[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[42]) );
  DFF \sreg_reg[43]  ( .D(sreg[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[43]) );
  DFF \sreg_reg[44]  ( .D(sreg[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[44]) );
  DFF \sreg_reg[45]  ( .D(sreg[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[45]) );
  DFF \sreg_reg[46]  ( .D(sreg[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[46]) );
  DFF \sreg_reg[47]  ( .D(sreg[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[47]) );
  DFF \sreg_reg[48]  ( .D(sreg[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[48]) );
  DFF \sreg_reg[49]  ( .D(sreg[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[49]) );
  DFF \sreg_reg[50]  ( .D(sreg[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[50]) );
  DFF \sreg_reg[51]  ( .D(sreg[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[51]) );
  DFF \sreg_reg[52]  ( .D(sreg[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[52]) );
  DFF \sreg_reg[53]  ( .D(sreg[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[53]) );
  DFF \sreg_reg[54]  ( .D(sreg[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[54]) );
  DFF \sreg_reg[55]  ( .D(sreg[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[55]) );
  DFF \sreg_reg[56]  ( .D(sreg[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[56]) );
  DFF \sreg_reg[57]  ( .D(sreg[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[57]) );
  DFF \sreg_reg[58]  ( .D(sreg[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[58]) );
  DFF \sreg_reg[59]  ( .D(sreg[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[59]) );
  DFF \sreg_reg[60]  ( .D(sreg[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[60]) );
  DFF \sreg_reg[61]  ( .D(sreg[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[61]) );
  DFF \sreg_reg[62]  ( .D(sreg[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[62]) );
  DFF \sreg_reg[63]  ( .D(sreg[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[63]) );
  DFF \sreg_reg[64]  ( .D(sreg[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[64]) );
  DFF \sreg_reg[65]  ( .D(sreg[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[65]) );
  DFF \sreg_reg[66]  ( .D(sreg[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[66]) );
  DFF \sreg_reg[67]  ( .D(sreg[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[67]) );
  DFF \sreg_reg[68]  ( .D(sreg[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[68]) );
  DFF \sreg_reg[69]  ( .D(sreg[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[69]) );
  DFF \sreg_reg[70]  ( .D(sreg[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[70]) );
  DFF \sreg_reg[71]  ( .D(sreg[72]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[71]) );
  DFF \sreg_reg[72]  ( .D(sreg[73]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[72]) );
  DFF \sreg_reg[73]  ( .D(sreg[74]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[73]) );
  DFF \sreg_reg[74]  ( .D(sreg[75]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[74]) );
  DFF \sreg_reg[75]  ( .D(sreg[76]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[75]) );
  DFF \sreg_reg[76]  ( .D(sreg[77]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[76]) );
  DFF \sreg_reg[77]  ( .D(sreg[78]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[77]) );
  DFF \sreg_reg[78]  ( .D(sreg[79]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[78]) );
  DFF \sreg_reg[79]  ( .D(sreg[80]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[79]) );
  DFF \sreg_reg[80]  ( .D(sreg[81]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[80]) );
  DFF \sreg_reg[81]  ( .D(sreg[82]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[81]) );
  DFF \sreg_reg[82]  ( .D(sreg[83]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[82]) );
  DFF \sreg_reg[83]  ( .D(sreg[84]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[83]) );
  DFF \sreg_reg[84]  ( .D(sreg[85]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[84]) );
  DFF \sreg_reg[85]  ( .D(sreg[86]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[85]) );
  DFF \sreg_reg[86]  ( .D(sreg[87]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[86]) );
  DFF \sreg_reg[87]  ( .D(sreg[88]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[87]) );
  DFF \sreg_reg[88]  ( .D(sreg[89]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[88]) );
  DFF \sreg_reg[89]  ( .D(sreg[90]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[89]) );
  DFF \sreg_reg[90]  ( .D(sreg[91]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[90]) );
  DFF \sreg_reg[91]  ( .D(sreg[92]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[91]) );
  DFF \sreg_reg[92]  ( .D(sreg[93]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[92]) );
  DFF \sreg_reg[93]  ( .D(sreg[94]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[93]) );
  DFF \sreg_reg[94]  ( .D(sreg[95]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[94]) );
  DFF \sreg_reg[95]  ( .D(sreg[96]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[95]) );
  DFF \sreg_reg[96]  ( .D(sreg[97]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[96]) );
  DFF \sreg_reg[97]  ( .D(sreg[98]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[97]) );
  DFF \sreg_reg[98]  ( .D(sreg[99]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[98]) );
  DFF \sreg_reg[99]  ( .D(sreg[100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[99]) );
  DFF \sreg_reg[100]  ( .D(sreg[101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[100]) );
  DFF \sreg_reg[101]  ( .D(sreg[102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[101]) );
  DFF \sreg_reg[102]  ( .D(sreg[103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[102]) );
  DFF \sreg_reg[103]  ( .D(sreg[104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[103]) );
  DFF \sreg_reg[104]  ( .D(sreg[105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[104]) );
  DFF \sreg_reg[105]  ( .D(sreg[106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[105]) );
  DFF \sreg_reg[106]  ( .D(sreg[107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[106]) );
  DFF \sreg_reg[107]  ( .D(sreg[108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[107]) );
  DFF \sreg_reg[108]  ( .D(sreg[109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[108]) );
  DFF \sreg_reg[109]  ( .D(sreg[110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[109]) );
  DFF \sreg_reg[110]  ( .D(sreg[111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[110]) );
  DFF \sreg_reg[111]  ( .D(sreg[112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[111]) );
  DFF \sreg_reg[112]  ( .D(sreg[113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[112]) );
  DFF \sreg_reg[113]  ( .D(sreg[114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[113]) );
  DFF \sreg_reg[114]  ( .D(sreg[115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[114]) );
  DFF \sreg_reg[115]  ( .D(sreg[116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[115]) );
  DFF \sreg_reg[116]  ( .D(sreg[117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[116]) );
  DFF \sreg_reg[117]  ( .D(sreg[118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[117]) );
  DFF \sreg_reg[118]  ( .D(sreg[119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[118]) );
  DFF \sreg_reg[119]  ( .D(sreg[120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[119]) );
  DFF \sreg_reg[120]  ( .D(sreg[121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[120]) );
  DFF \sreg_reg[121]  ( .D(sreg[122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[121]) );
  DFF \sreg_reg[122]  ( .D(sreg[123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[122]) );
  DFF \sreg_reg[123]  ( .D(sreg[124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[123]) );
  DFF \sreg_reg[124]  ( .D(sreg[125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[124]) );
  DFF \sreg_reg[125]  ( .D(sreg[126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[125]) );
  DFF \sreg_reg[126]  ( .D(sreg[127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[126]) );
  DFF \sreg_reg[127]  ( .D(sreg[128]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[127]) );
  DFF \sreg_reg[128]  ( .D(sreg[129]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[128]) );
  DFF \sreg_reg[129]  ( .D(sreg[130]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[129]) );
  DFF \sreg_reg[130]  ( .D(sreg[131]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[130]) );
  DFF \sreg_reg[131]  ( .D(sreg[132]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[131]) );
  DFF \sreg_reg[132]  ( .D(sreg[133]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[132]) );
  DFF \sreg_reg[133]  ( .D(sreg[134]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[133]) );
  DFF \sreg_reg[134]  ( .D(sreg[135]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[134]) );
  DFF \sreg_reg[135]  ( .D(sreg[136]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[135]) );
  DFF \sreg_reg[136]  ( .D(sreg[137]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[136]) );
  DFF \sreg_reg[137]  ( .D(sreg[138]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[137]) );
  DFF \sreg_reg[138]  ( .D(sreg[139]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[138]) );
  DFF \sreg_reg[139]  ( .D(sreg[140]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[139]) );
  DFF \sreg_reg[140]  ( .D(sreg[141]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[140]) );
  DFF \sreg_reg[141]  ( .D(sreg[142]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[141]) );
  DFF \sreg_reg[142]  ( .D(sreg[143]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[142]) );
  DFF \sreg_reg[143]  ( .D(sreg[144]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[143]) );
  DFF \sreg_reg[144]  ( .D(sreg[145]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[144]) );
  DFF \sreg_reg[145]  ( .D(sreg[146]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[145]) );
  DFF \sreg_reg[146]  ( .D(sreg[147]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[146]) );
  DFF \sreg_reg[147]  ( .D(sreg[148]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[147]) );
  DFF \sreg_reg[148]  ( .D(sreg[149]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[148]) );
  DFF \sreg_reg[149]  ( .D(sreg[150]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[149]) );
  DFF \sreg_reg[150]  ( .D(sreg[151]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[150]) );
  DFF \sreg_reg[151]  ( .D(sreg[152]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[151]) );
  DFF \sreg_reg[152]  ( .D(sreg[153]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[152]) );
  DFF \sreg_reg[153]  ( .D(sreg[154]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[153]) );
  DFF \sreg_reg[154]  ( .D(sreg[155]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[154]) );
  DFF \sreg_reg[155]  ( .D(sreg[156]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[155]) );
  DFF \sreg_reg[156]  ( .D(sreg[157]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[156]) );
  DFF \sreg_reg[157]  ( .D(sreg[158]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[157]) );
  DFF \sreg_reg[158]  ( .D(sreg[159]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[158]) );
  DFF \sreg_reg[159]  ( .D(sreg[160]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[159]) );
  DFF \sreg_reg[160]  ( .D(sreg[161]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[160]) );
  DFF \sreg_reg[161]  ( .D(sreg[162]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[161]) );
  DFF \sreg_reg[162]  ( .D(sreg[163]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[162]) );
  DFF \sreg_reg[163]  ( .D(sreg[164]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[163]) );
  DFF \sreg_reg[164]  ( .D(sreg[165]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[164]) );
  DFF \sreg_reg[165]  ( .D(sreg[166]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[165]) );
  DFF \sreg_reg[166]  ( .D(sreg[167]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[166]) );
  DFF \sreg_reg[167]  ( .D(sreg[168]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[167]) );
  DFF \sreg_reg[168]  ( .D(sreg[169]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[168]) );
  DFF \sreg_reg[169]  ( .D(sreg[170]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[169]) );
  DFF \sreg_reg[170]  ( .D(sreg[171]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[170]) );
  DFF \sreg_reg[171]  ( .D(sreg[172]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[171]) );
  DFF \sreg_reg[172]  ( .D(sreg[173]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[172]) );
  DFF \sreg_reg[173]  ( .D(sreg[174]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[173]) );
  DFF \sreg_reg[174]  ( .D(sreg[175]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[174]) );
  DFF \sreg_reg[175]  ( .D(sreg[176]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[175]) );
  DFF \sreg_reg[176]  ( .D(sreg[177]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[176]) );
  DFF \sreg_reg[177]  ( .D(sreg[178]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[177]) );
  DFF \sreg_reg[178]  ( .D(sreg[179]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[178]) );
  DFF \sreg_reg[179]  ( .D(sreg[180]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[179]) );
  DFF \sreg_reg[180]  ( .D(sreg[181]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[180]) );
  DFF \sreg_reg[181]  ( .D(sreg[182]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[181]) );
  DFF \sreg_reg[182]  ( .D(sreg[183]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[182]) );
  DFF \sreg_reg[183]  ( .D(sreg[184]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[183]) );
  DFF \sreg_reg[184]  ( .D(sreg[185]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[184]) );
  DFF \sreg_reg[185]  ( .D(sreg[186]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[185]) );
  DFF \sreg_reg[186]  ( .D(sreg[187]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[186]) );
  DFF \sreg_reg[187]  ( .D(sreg[188]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[187]) );
  DFF \sreg_reg[188]  ( .D(sreg[189]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[188]) );
  DFF \sreg_reg[189]  ( .D(sreg[190]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[189]) );
  DFF \sreg_reg[190]  ( .D(sreg[191]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[190]) );
  DFF \sreg_reg[191]  ( .D(sreg[192]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[191]) );
  DFF \sreg_reg[192]  ( .D(sreg[193]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[192]) );
  DFF \sreg_reg[193]  ( .D(sreg[194]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[193]) );
  DFF \sreg_reg[194]  ( .D(sreg[195]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[194]) );
  DFF \sreg_reg[195]  ( .D(sreg[196]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[195]) );
  DFF \sreg_reg[196]  ( .D(sreg[197]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[196]) );
  DFF \sreg_reg[197]  ( .D(sreg[198]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[197]) );
  DFF \sreg_reg[198]  ( .D(sreg[199]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[198]) );
  DFF \sreg_reg[199]  ( .D(sreg[200]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[199]) );
  DFF \sreg_reg[200]  ( .D(sreg[201]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[200]) );
  DFF \sreg_reg[201]  ( .D(sreg[202]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[201]) );
  DFF \sreg_reg[202]  ( .D(sreg[203]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[202]) );
  DFF \sreg_reg[203]  ( .D(sreg[204]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[203]) );
  DFF \sreg_reg[204]  ( .D(sreg[205]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[204]) );
  DFF \sreg_reg[205]  ( .D(sreg[206]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[205]) );
  DFF \sreg_reg[206]  ( .D(sreg[207]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[206]) );
  DFF \sreg_reg[207]  ( .D(sreg[208]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[207]) );
  DFF \sreg_reg[208]  ( .D(sreg[209]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[208]) );
  DFF \sreg_reg[209]  ( .D(sreg[210]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[209]) );
  DFF \sreg_reg[210]  ( .D(sreg[211]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[210]) );
  DFF \sreg_reg[211]  ( .D(sreg[212]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[211]) );
  DFF \sreg_reg[212]  ( .D(sreg[213]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[212]) );
  DFF \sreg_reg[213]  ( .D(sreg[214]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[213]) );
  DFF \sreg_reg[214]  ( .D(sreg[215]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[214]) );
  DFF \sreg_reg[215]  ( .D(sreg[216]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[215]) );
  DFF \sreg_reg[216]  ( .D(sreg[217]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[216]) );
  DFF \sreg_reg[217]  ( .D(sreg[218]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[217]) );
  DFF \sreg_reg[218]  ( .D(sreg[219]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[218]) );
  DFF \sreg_reg[219]  ( .D(sreg[220]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[219]) );
  DFF \sreg_reg[220]  ( .D(sreg[221]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[220]) );
  DFF \sreg_reg[221]  ( .D(sreg[222]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[221]) );
  DFF \sreg_reg[222]  ( .D(sreg[223]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[222]) );
  DFF \sreg_reg[223]  ( .D(sreg[224]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[223]) );
  DFF \sreg_reg[224]  ( .D(sreg[225]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[224]) );
  DFF \sreg_reg[225]  ( .D(sreg[226]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[225]) );
  DFF \sreg_reg[226]  ( .D(sreg[227]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[226]) );
  DFF \sreg_reg[227]  ( .D(sreg[228]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[227]) );
  DFF \sreg_reg[228]  ( .D(sreg[229]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[228]) );
  DFF \sreg_reg[229]  ( .D(sreg[230]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[229]) );
  DFF \sreg_reg[230]  ( .D(sreg[231]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[230]) );
  DFF \sreg_reg[231]  ( .D(sreg[232]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[231]) );
  DFF \sreg_reg[232]  ( .D(sreg[233]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[232]) );
  DFF \sreg_reg[233]  ( .D(sreg[234]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[233]) );
  DFF \sreg_reg[234]  ( .D(sreg[235]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[234]) );
  DFF \sreg_reg[235]  ( .D(sreg[236]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[235]) );
  DFF \sreg_reg[236]  ( .D(sreg[237]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[236]) );
  DFF \sreg_reg[237]  ( .D(sreg[238]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[237]) );
  DFF \sreg_reg[238]  ( .D(sreg[239]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[238]) );
  DFF \sreg_reg[239]  ( .D(sreg[240]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[239]) );
  DFF \sreg_reg[240]  ( .D(sreg[241]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[240]) );
  DFF \sreg_reg[241]  ( .D(sreg[242]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[241]) );
  DFF \sreg_reg[242]  ( .D(sreg[243]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[242]) );
  DFF \sreg_reg[243]  ( .D(sreg[244]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[243]) );
  DFF \sreg_reg[244]  ( .D(sreg[245]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[244]) );
  DFF \sreg_reg[245]  ( .D(sreg[246]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[245]) );
  DFF \sreg_reg[246]  ( .D(sreg[247]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[246]) );
  DFF \sreg_reg[247]  ( .D(sreg[248]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[247]) );
  DFF \sreg_reg[248]  ( .D(sreg[249]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[248]) );
  DFF \sreg_reg[249]  ( .D(sreg[250]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[249]) );
  DFF \sreg_reg[250]  ( .D(sreg[251]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[250]) );
  DFF \sreg_reg[251]  ( .D(sreg[252]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[251]) );
  DFF \sreg_reg[252]  ( .D(sreg[253]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[252]) );
  DFF \sreg_reg[253]  ( .D(sreg[254]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[253]) );
  DFF \sreg_reg[254]  ( .D(sreg[255]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[254]) );
  DFF \sreg_reg[255]  ( .D(sreg[256]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[255]) );
  DFF \sreg_reg[256]  ( .D(sreg[257]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[256]) );
  DFF \sreg_reg[257]  ( .D(sreg[258]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[257]) );
  DFF \sreg_reg[258]  ( .D(sreg[259]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[258]) );
  DFF \sreg_reg[259]  ( .D(sreg[260]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[259]) );
  DFF \sreg_reg[260]  ( .D(sreg[261]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[260]) );
  DFF \sreg_reg[261]  ( .D(sreg[262]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[261]) );
  DFF \sreg_reg[262]  ( .D(sreg[263]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[262]) );
  DFF \sreg_reg[263]  ( .D(sreg[264]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[263]) );
  DFF \sreg_reg[264]  ( .D(sreg[265]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[264]) );
  DFF \sreg_reg[265]  ( .D(sreg[266]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[265]) );
  DFF \sreg_reg[266]  ( .D(sreg[267]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[266]) );
  DFF \sreg_reg[267]  ( .D(sreg[268]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[267]) );
  DFF \sreg_reg[268]  ( .D(sreg[269]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[268]) );
  DFF \sreg_reg[269]  ( .D(sreg[270]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[269]) );
  DFF \sreg_reg[270]  ( .D(sreg[271]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[270]) );
  DFF \sreg_reg[271]  ( .D(sreg[272]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[271]) );
  DFF \sreg_reg[272]  ( .D(sreg[273]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[272]) );
  DFF \sreg_reg[273]  ( .D(sreg[274]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[273]) );
  DFF \sreg_reg[274]  ( .D(sreg[275]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[274]) );
  DFF \sreg_reg[275]  ( .D(sreg[276]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[275]) );
  DFF \sreg_reg[276]  ( .D(sreg[277]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[276]) );
  DFF \sreg_reg[277]  ( .D(sreg[278]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[277]) );
  DFF \sreg_reg[278]  ( .D(sreg[279]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[278]) );
  DFF \sreg_reg[279]  ( .D(sreg[280]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[279]) );
  DFF \sreg_reg[280]  ( .D(sreg[281]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[280]) );
  DFF \sreg_reg[281]  ( .D(sreg[282]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[281]) );
  DFF \sreg_reg[282]  ( .D(sreg[283]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[282]) );
  DFF \sreg_reg[283]  ( .D(sreg[284]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[283]) );
  DFF \sreg_reg[284]  ( .D(sreg[285]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[284]) );
  DFF \sreg_reg[285]  ( .D(sreg[286]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[285]) );
  DFF \sreg_reg[286]  ( .D(sreg[287]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[286]) );
  DFF \sreg_reg[287]  ( .D(sreg[288]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[287]) );
  DFF \sreg_reg[288]  ( .D(sreg[289]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[288]) );
  DFF \sreg_reg[289]  ( .D(sreg[290]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[289]) );
  DFF \sreg_reg[290]  ( .D(sreg[291]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[290]) );
  DFF \sreg_reg[291]  ( .D(sreg[292]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[291]) );
  DFF \sreg_reg[292]  ( .D(sreg[293]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[292]) );
  DFF \sreg_reg[293]  ( .D(sreg[294]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[293]) );
  DFF \sreg_reg[294]  ( .D(sreg[295]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[294]) );
  DFF \sreg_reg[295]  ( .D(sreg[296]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[295]) );
  DFF \sreg_reg[296]  ( .D(sreg[297]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[296]) );
  DFF \sreg_reg[297]  ( .D(sreg[298]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[297]) );
  DFF \sreg_reg[298]  ( .D(sreg[299]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[298]) );
  DFF \sreg_reg[299]  ( .D(sreg[300]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[299]) );
  DFF \sreg_reg[300]  ( .D(sreg[301]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[300]) );
  DFF \sreg_reg[301]  ( .D(sreg[302]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[301]) );
  DFF \sreg_reg[302]  ( .D(sreg[303]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[302]) );
  DFF \sreg_reg[303]  ( .D(sreg[304]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[303]) );
  DFF \sreg_reg[304]  ( .D(sreg[305]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[304]) );
  DFF \sreg_reg[305]  ( .D(sreg[306]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[305]) );
  DFF \sreg_reg[306]  ( .D(sreg[307]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[306]) );
  DFF \sreg_reg[307]  ( .D(sreg[308]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[307]) );
  DFF \sreg_reg[308]  ( .D(sreg[309]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[308]) );
  DFF \sreg_reg[309]  ( .D(sreg[310]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[309]) );
  DFF \sreg_reg[310]  ( .D(sreg[311]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[310]) );
  DFF \sreg_reg[311]  ( .D(sreg[312]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[311]) );
  DFF \sreg_reg[312]  ( .D(sreg[313]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[312]) );
  DFF \sreg_reg[313]  ( .D(sreg[314]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[313]) );
  DFF \sreg_reg[314]  ( .D(sreg[315]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[314]) );
  DFF \sreg_reg[315]  ( .D(sreg[316]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[315]) );
  DFF \sreg_reg[316]  ( .D(sreg[317]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[316]) );
  DFF \sreg_reg[317]  ( .D(sreg[318]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[317]) );
  DFF \sreg_reg[318]  ( .D(sreg[319]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[318]) );
  DFF \sreg_reg[319]  ( .D(sreg[320]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[319]) );
  DFF \sreg_reg[320]  ( .D(sreg[321]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[320]) );
  DFF \sreg_reg[321]  ( .D(sreg[322]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[321]) );
  DFF \sreg_reg[322]  ( .D(sreg[323]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[322]) );
  DFF \sreg_reg[323]  ( .D(sreg[324]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[323]) );
  DFF \sreg_reg[324]  ( .D(sreg[325]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[324]) );
  DFF \sreg_reg[325]  ( .D(sreg[326]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[325]) );
  DFF \sreg_reg[326]  ( .D(sreg[327]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[326]) );
  DFF \sreg_reg[327]  ( .D(sreg[328]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[327]) );
  DFF \sreg_reg[328]  ( .D(sreg[329]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[328]) );
  DFF \sreg_reg[329]  ( .D(sreg[330]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[329]) );
  DFF \sreg_reg[330]  ( .D(sreg[331]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[330]) );
  DFF \sreg_reg[331]  ( .D(sreg[332]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[331]) );
  DFF \sreg_reg[332]  ( .D(sreg[333]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[332]) );
  DFF \sreg_reg[333]  ( .D(sreg[334]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[333]) );
  DFF \sreg_reg[334]  ( .D(sreg[335]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[334]) );
  DFF \sreg_reg[335]  ( .D(sreg[336]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[335]) );
  DFF \sreg_reg[336]  ( .D(sreg[337]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[336]) );
  DFF \sreg_reg[337]  ( .D(sreg[338]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[337]) );
  DFF \sreg_reg[338]  ( .D(sreg[339]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[338]) );
  DFF \sreg_reg[339]  ( .D(sreg[340]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[339]) );
  DFF \sreg_reg[340]  ( .D(sreg[341]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[340]) );
  DFF \sreg_reg[341]  ( .D(sreg[342]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[341]) );
  DFF \sreg_reg[342]  ( .D(sreg[343]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[342]) );
  DFF \sreg_reg[343]  ( .D(sreg[344]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[343]) );
  DFF \sreg_reg[344]  ( .D(sreg[345]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[344]) );
  DFF \sreg_reg[345]  ( .D(sreg[346]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[345]) );
  DFF \sreg_reg[346]  ( .D(sreg[347]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[346]) );
  DFF \sreg_reg[347]  ( .D(sreg[348]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[347]) );
  DFF \sreg_reg[348]  ( .D(sreg[349]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[348]) );
  DFF \sreg_reg[349]  ( .D(sreg[350]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[349]) );
  DFF \sreg_reg[350]  ( .D(sreg[351]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[350]) );
  DFF \sreg_reg[351]  ( .D(sreg[352]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[351]) );
  DFF \sreg_reg[352]  ( .D(sreg[353]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[352]) );
  DFF \sreg_reg[353]  ( .D(sreg[354]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[353]) );
  DFF \sreg_reg[354]  ( .D(sreg[355]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[354]) );
  DFF \sreg_reg[355]  ( .D(sreg[356]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[355]) );
  DFF \sreg_reg[356]  ( .D(sreg[357]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[356]) );
  DFF \sreg_reg[357]  ( .D(sreg[358]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[357]) );
  DFF \sreg_reg[358]  ( .D(sreg[359]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[358]) );
  DFF \sreg_reg[359]  ( .D(sreg[360]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[359]) );
  DFF \sreg_reg[360]  ( .D(sreg[361]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[360]) );
  DFF \sreg_reg[361]  ( .D(sreg[362]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[361]) );
  DFF \sreg_reg[362]  ( .D(sreg[363]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[362]) );
  DFF \sreg_reg[363]  ( .D(sreg[364]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[363]) );
  DFF \sreg_reg[364]  ( .D(sreg[365]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[364]) );
  DFF \sreg_reg[365]  ( .D(sreg[366]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[365]) );
  DFF \sreg_reg[366]  ( .D(sreg[367]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[366]) );
  DFF \sreg_reg[367]  ( .D(sreg[368]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[367]) );
  DFF \sreg_reg[368]  ( .D(sreg[369]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[368]) );
  DFF \sreg_reg[369]  ( .D(sreg[370]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[369]) );
  DFF \sreg_reg[370]  ( .D(sreg[371]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[370]) );
  DFF \sreg_reg[371]  ( .D(sreg[372]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[371]) );
  DFF \sreg_reg[372]  ( .D(sreg[373]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[372]) );
  DFF \sreg_reg[373]  ( .D(sreg[374]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[373]) );
  DFF \sreg_reg[374]  ( .D(sreg[375]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[374]) );
  DFF \sreg_reg[375]  ( .D(sreg[376]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[375]) );
  DFF \sreg_reg[376]  ( .D(sreg[377]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[376]) );
  DFF \sreg_reg[377]  ( .D(sreg[378]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[377]) );
  DFF \sreg_reg[378]  ( .D(sreg[379]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[378]) );
  DFF \sreg_reg[379]  ( .D(sreg[380]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[379]) );
  DFF \sreg_reg[380]  ( .D(sreg[381]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[380]) );
  DFF \sreg_reg[381]  ( .D(sreg[382]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[381]) );
  DFF \sreg_reg[382]  ( .D(sreg[383]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[382]) );
  DFF \sreg_reg[383]  ( .D(sreg[384]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[383]) );
  DFF \sreg_reg[384]  ( .D(sreg[385]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[384]) );
  DFF \sreg_reg[385]  ( .D(sreg[386]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[385]) );
  DFF \sreg_reg[386]  ( .D(sreg[387]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[386]) );
  DFF \sreg_reg[387]  ( .D(sreg[388]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[387]) );
  DFF \sreg_reg[388]  ( .D(sreg[389]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[388]) );
  DFF \sreg_reg[389]  ( .D(sreg[390]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[389]) );
  DFF \sreg_reg[390]  ( .D(sreg[391]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[390]) );
  DFF \sreg_reg[391]  ( .D(sreg[392]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[391]) );
  DFF \sreg_reg[392]  ( .D(sreg[393]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[392]) );
  DFF \sreg_reg[393]  ( .D(sreg[394]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[393]) );
  DFF \sreg_reg[394]  ( .D(sreg[395]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[394]) );
  DFF \sreg_reg[395]  ( .D(sreg[396]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[395]) );
  DFF \sreg_reg[396]  ( .D(sreg[397]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[396]) );
  DFF \sreg_reg[397]  ( .D(sreg[398]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[397]) );
  DFF \sreg_reg[398]  ( .D(sreg[399]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[398]) );
  DFF \sreg_reg[399]  ( .D(sreg[400]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[399]) );
  DFF \sreg_reg[400]  ( .D(sreg[401]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[400]) );
  DFF \sreg_reg[401]  ( .D(sreg[402]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[401]) );
  DFF \sreg_reg[402]  ( .D(sreg[403]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[402]) );
  DFF \sreg_reg[403]  ( .D(sreg[404]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[403]) );
  DFF \sreg_reg[404]  ( .D(sreg[405]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[404]) );
  DFF \sreg_reg[405]  ( .D(sreg[406]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[405]) );
  DFF \sreg_reg[406]  ( .D(sreg[407]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[406]) );
  DFF \sreg_reg[407]  ( .D(sreg[408]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[407]) );
  DFF \sreg_reg[408]  ( .D(sreg[409]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[408]) );
  DFF \sreg_reg[409]  ( .D(sreg[410]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[409]) );
  DFF \sreg_reg[410]  ( .D(sreg[411]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[410]) );
  DFF \sreg_reg[411]  ( .D(sreg[412]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[411]) );
  DFF \sreg_reg[412]  ( .D(sreg[413]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[412]) );
  DFF \sreg_reg[413]  ( .D(sreg[414]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[413]) );
  DFF \sreg_reg[414]  ( .D(sreg[415]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[414]) );
  DFF \sreg_reg[415]  ( .D(sreg[416]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[415]) );
  DFF \sreg_reg[416]  ( .D(sreg[417]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[416]) );
  DFF \sreg_reg[417]  ( .D(sreg[418]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[417]) );
  DFF \sreg_reg[418]  ( .D(sreg[419]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[418]) );
  DFF \sreg_reg[419]  ( .D(sreg[420]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[419]) );
  DFF \sreg_reg[420]  ( .D(sreg[421]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[420]) );
  DFF \sreg_reg[421]  ( .D(sreg[422]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[421]) );
  DFF \sreg_reg[422]  ( .D(sreg[423]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[422]) );
  DFF \sreg_reg[423]  ( .D(sreg[424]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[423]) );
  DFF \sreg_reg[424]  ( .D(sreg[425]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[424]) );
  DFF \sreg_reg[425]  ( .D(sreg[426]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[425]) );
  DFF \sreg_reg[426]  ( .D(sreg[427]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[426]) );
  DFF \sreg_reg[427]  ( .D(sreg[428]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[427]) );
  DFF \sreg_reg[428]  ( .D(sreg[429]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[428]) );
  DFF \sreg_reg[429]  ( .D(sreg[430]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[429]) );
  DFF \sreg_reg[430]  ( .D(sreg[431]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[430]) );
  DFF \sreg_reg[431]  ( .D(sreg[432]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[431]) );
  DFF \sreg_reg[432]  ( .D(sreg[433]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[432]) );
  DFF \sreg_reg[433]  ( .D(sreg[434]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[433]) );
  DFF \sreg_reg[434]  ( .D(sreg[435]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[434]) );
  DFF \sreg_reg[435]  ( .D(sreg[436]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[435]) );
  DFF \sreg_reg[436]  ( .D(sreg[437]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[436]) );
  DFF \sreg_reg[437]  ( .D(sreg[438]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[437]) );
  DFF \sreg_reg[438]  ( .D(sreg[439]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[438]) );
  DFF \sreg_reg[439]  ( .D(sreg[440]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[439]) );
  DFF \sreg_reg[440]  ( .D(sreg[441]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[440]) );
  DFF \sreg_reg[441]  ( .D(sreg[442]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[441]) );
  DFF \sreg_reg[442]  ( .D(sreg[443]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[442]) );
  DFF \sreg_reg[443]  ( .D(sreg[444]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[443]) );
  DFF \sreg_reg[444]  ( .D(sreg[445]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[444]) );
  DFF \sreg_reg[445]  ( .D(sreg[446]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[445]) );
  DFF \sreg_reg[446]  ( .D(sreg[447]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[446]) );
  DFF \sreg_reg[447]  ( .D(sreg[448]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[447]) );
  DFF \sreg_reg[448]  ( .D(sreg[449]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[448]) );
  DFF \sreg_reg[449]  ( .D(sreg[450]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[449]) );
  DFF \sreg_reg[450]  ( .D(sreg[451]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[450]) );
  DFF \sreg_reg[451]  ( .D(sreg[452]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[451]) );
  DFF \sreg_reg[452]  ( .D(sreg[453]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[452]) );
  DFF \sreg_reg[453]  ( .D(sreg[454]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[453]) );
  DFF \sreg_reg[454]  ( .D(sreg[455]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[454]) );
  DFF \sreg_reg[455]  ( .D(sreg[456]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[455]) );
  DFF \sreg_reg[456]  ( .D(sreg[457]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[456]) );
  DFF \sreg_reg[457]  ( .D(sreg[458]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[457]) );
  DFF \sreg_reg[458]  ( .D(sreg[459]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[458]) );
  DFF \sreg_reg[459]  ( .D(sreg[460]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[459]) );
  DFF \sreg_reg[460]  ( .D(sreg[461]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[460]) );
  DFF \sreg_reg[461]  ( .D(sreg[462]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[461]) );
  DFF \sreg_reg[462]  ( .D(sreg[463]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[462]) );
  DFF \sreg_reg[463]  ( .D(sreg[464]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[463]) );
  DFF \sreg_reg[464]  ( .D(sreg[465]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[464]) );
  DFF \sreg_reg[465]  ( .D(sreg[466]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[465]) );
  DFF \sreg_reg[466]  ( .D(sreg[467]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[466]) );
  DFF \sreg_reg[467]  ( .D(sreg[468]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[467]) );
  DFF \sreg_reg[468]  ( .D(sreg[469]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[468]) );
  DFF \sreg_reg[469]  ( .D(sreg[470]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[469]) );
  DFF \sreg_reg[470]  ( .D(sreg[471]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[470]) );
  DFF \sreg_reg[471]  ( .D(sreg[472]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[471]) );
  DFF \sreg_reg[472]  ( .D(sreg[473]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[472]) );
  DFF \sreg_reg[473]  ( .D(sreg[474]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[473]) );
  DFF \sreg_reg[474]  ( .D(sreg[475]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[474]) );
  DFF \sreg_reg[475]  ( .D(sreg[476]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[475]) );
  DFF \sreg_reg[476]  ( .D(sreg[477]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[476]) );
  DFF \sreg_reg[477]  ( .D(sreg[478]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[477]) );
  DFF \sreg_reg[478]  ( .D(sreg[479]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[478]) );
  DFF \sreg_reg[479]  ( .D(sreg[480]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[479]) );
  DFF \sreg_reg[480]  ( .D(sreg[481]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[480]) );
  DFF \sreg_reg[481]  ( .D(sreg[482]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[481]) );
  DFF \sreg_reg[482]  ( .D(sreg[483]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[482]) );
  DFF \sreg_reg[483]  ( .D(sreg[484]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[483]) );
  DFF \sreg_reg[484]  ( .D(sreg[485]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[484]) );
  DFF \sreg_reg[485]  ( .D(sreg[486]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[485]) );
  DFF \sreg_reg[486]  ( .D(sreg[487]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[486]) );
  DFF \sreg_reg[487]  ( .D(sreg[488]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[487]) );
  DFF \sreg_reg[488]  ( .D(sreg[489]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[488]) );
  DFF \sreg_reg[489]  ( .D(sreg[490]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[489]) );
  DFF \sreg_reg[490]  ( .D(sreg[491]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[490]) );
  DFF \sreg_reg[491]  ( .D(sreg[492]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[491]) );
  DFF \sreg_reg[492]  ( .D(sreg[493]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[492]) );
  DFF \sreg_reg[493]  ( .D(sreg[494]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[493]) );
  DFF \sreg_reg[494]  ( .D(sreg[495]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[494]) );
  DFF \sreg_reg[495]  ( .D(sreg[496]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[495]) );
  DFF \sreg_reg[496]  ( .D(sreg[497]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[496]) );
  DFF \sreg_reg[497]  ( .D(sreg[498]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[497]) );
  DFF \sreg_reg[498]  ( .D(sreg[499]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[498]) );
  DFF \sreg_reg[499]  ( .D(sreg[500]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[499]) );
  DFF \sreg_reg[500]  ( .D(sreg[501]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[500]) );
  DFF \sreg_reg[501]  ( .D(sreg[502]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[501]) );
  DFF \sreg_reg[502]  ( .D(sreg[503]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[502]) );
  DFF \sreg_reg[503]  ( .D(sreg[504]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[503]) );
  DFF \sreg_reg[504]  ( .D(sreg[505]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[504]) );
  DFF \sreg_reg[505]  ( .D(sreg[506]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[505]) );
  DFF \sreg_reg[506]  ( .D(sreg[507]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[506]) );
  DFF \sreg_reg[507]  ( .D(sreg[508]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[507]) );
  DFF \sreg_reg[508]  ( .D(sreg[509]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[508]) );
  DFF \sreg_reg[509]  ( .D(sreg[510]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[509]) );
  DFF \sreg_reg[510]  ( .D(sreg[511]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[510]) );
  DFF \sreg_reg[511]  ( .D(sreg[512]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[511]) );
  DFF \sreg_reg[512]  ( .D(sreg[513]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[512]) );
  DFF \sreg_reg[513]  ( .D(sreg[514]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[513]) );
  DFF \sreg_reg[514]  ( .D(sreg[515]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[514]) );
  DFF \sreg_reg[515]  ( .D(sreg[516]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[515]) );
  DFF \sreg_reg[516]  ( .D(sreg[517]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[516]) );
  DFF \sreg_reg[517]  ( .D(sreg[518]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[517]) );
  DFF \sreg_reg[518]  ( .D(sreg[519]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[518]) );
  DFF \sreg_reg[519]  ( .D(sreg[520]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[519]) );
  DFF \sreg_reg[520]  ( .D(sreg[521]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[520]) );
  DFF \sreg_reg[521]  ( .D(sreg[522]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[521]) );
  DFF \sreg_reg[522]  ( .D(sreg[523]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[522]) );
  DFF \sreg_reg[523]  ( .D(sreg[524]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[523]) );
  DFF \sreg_reg[524]  ( .D(sreg[525]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[524]) );
  DFF \sreg_reg[525]  ( .D(sreg[526]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[525]) );
  DFF \sreg_reg[526]  ( .D(sreg[527]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[526]) );
  DFF \sreg_reg[527]  ( .D(sreg[528]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[527]) );
  DFF \sreg_reg[528]  ( .D(sreg[529]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[528]) );
  DFF \sreg_reg[529]  ( .D(sreg[530]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[529]) );
  DFF \sreg_reg[530]  ( .D(sreg[531]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[530]) );
  DFF \sreg_reg[531]  ( .D(sreg[532]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[531]) );
  DFF \sreg_reg[532]  ( .D(sreg[533]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[532]) );
  DFF \sreg_reg[533]  ( .D(sreg[534]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[533]) );
  DFF \sreg_reg[534]  ( .D(sreg[535]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[534]) );
  DFF \sreg_reg[535]  ( .D(sreg[536]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[535]) );
  DFF \sreg_reg[536]  ( .D(sreg[537]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[536]) );
  DFF \sreg_reg[537]  ( .D(sreg[538]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[537]) );
  DFF \sreg_reg[538]  ( .D(sreg[539]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[538]) );
  DFF \sreg_reg[539]  ( .D(sreg[540]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[539]) );
  DFF \sreg_reg[540]  ( .D(sreg[541]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[540]) );
  DFF \sreg_reg[541]  ( .D(sreg[542]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[541]) );
  DFF \sreg_reg[542]  ( .D(sreg[543]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[542]) );
  DFF \sreg_reg[543]  ( .D(sreg[544]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[543]) );
  DFF \sreg_reg[544]  ( .D(sreg[545]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[544]) );
  DFF \sreg_reg[545]  ( .D(sreg[546]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[545]) );
  DFF \sreg_reg[546]  ( .D(sreg[547]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[546]) );
  DFF \sreg_reg[547]  ( .D(sreg[548]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[547]) );
  DFF \sreg_reg[548]  ( .D(sreg[549]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[548]) );
  DFF \sreg_reg[549]  ( .D(sreg[550]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[549]) );
  DFF \sreg_reg[550]  ( .D(sreg[551]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[550]) );
  DFF \sreg_reg[551]  ( .D(sreg[552]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[551]) );
  DFF \sreg_reg[552]  ( .D(sreg[553]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[552]) );
  DFF \sreg_reg[553]  ( .D(sreg[554]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[553]) );
  DFF \sreg_reg[554]  ( .D(sreg[555]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[554]) );
  DFF \sreg_reg[555]  ( .D(sreg[556]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[555]) );
  DFF \sreg_reg[556]  ( .D(sreg[557]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[556]) );
  DFF \sreg_reg[557]  ( .D(sreg[558]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[557]) );
  DFF \sreg_reg[558]  ( .D(sreg[559]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[558]) );
  DFF \sreg_reg[559]  ( .D(sreg[560]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[559]) );
  DFF \sreg_reg[560]  ( .D(sreg[561]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[560]) );
  DFF \sreg_reg[561]  ( .D(sreg[562]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[561]) );
  DFF \sreg_reg[562]  ( .D(sreg[563]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[562]) );
  DFF \sreg_reg[563]  ( .D(sreg[564]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[563]) );
  DFF \sreg_reg[564]  ( .D(sreg[565]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[564]) );
  DFF \sreg_reg[565]  ( .D(sreg[566]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[565]) );
  DFF \sreg_reg[566]  ( .D(sreg[567]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[566]) );
  DFF \sreg_reg[567]  ( .D(sreg[568]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[567]) );
  DFF \sreg_reg[568]  ( .D(sreg[569]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[568]) );
  DFF \sreg_reg[569]  ( .D(sreg[570]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[569]) );
  DFF \sreg_reg[570]  ( .D(sreg[571]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[570]) );
  DFF \sreg_reg[571]  ( .D(sreg[572]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[571]) );
  DFF \sreg_reg[572]  ( .D(sreg[573]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[572]) );
  DFF \sreg_reg[573]  ( .D(sreg[574]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[573]) );
  DFF \sreg_reg[574]  ( .D(sreg[575]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[574]) );
  DFF \sreg_reg[575]  ( .D(sreg[576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[575]) );
  DFF \sreg_reg[576]  ( .D(sreg[577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[576]) );
  DFF \sreg_reg[577]  ( .D(sreg[578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[577]) );
  DFF \sreg_reg[578]  ( .D(sreg[579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[578]) );
  DFF \sreg_reg[579]  ( .D(sreg[580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[579]) );
  DFF \sreg_reg[580]  ( .D(sreg[581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[580]) );
  DFF \sreg_reg[581]  ( .D(sreg[582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[581]) );
  DFF \sreg_reg[582]  ( .D(sreg[583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[582]) );
  DFF \sreg_reg[583]  ( .D(sreg[584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[583]) );
  DFF \sreg_reg[584]  ( .D(sreg[585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[584]) );
  DFF \sreg_reg[585]  ( .D(sreg[586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[585]) );
  DFF \sreg_reg[586]  ( .D(sreg[587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[586]) );
  DFF \sreg_reg[587]  ( .D(sreg[588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[587]) );
  DFF \sreg_reg[588]  ( .D(sreg[589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[588]) );
  DFF \sreg_reg[589]  ( .D(sreg[590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[589]) );
  DFF \sreg_reg[590]  ( .D(sreg[591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[590]) );
  DFF \sreg_reg[591]  ( .D(sreg[592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[591]) );
  DFF \sreg_reg[592]  ( .D(sreg[593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[592]) );
  DFF \sreg_reg[593]  ( .D(sreg[594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[593]) );
  DFF \sreg_reg[594]  ( .D(sreg[595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[594]) );
  DFF \sreg_reg[595]  ( .D(sreg[596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[595]) );
  DFF \sreg_reg[596]  ( .D(sreg[597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[596]) );
  DFF \sreg_reg[597]  ( .D(sreg[598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[597]) );
  DFF \sreg_reg[598]  ( .D(sreg[599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[598]) );
  DFF \sreg_reg[599]  ( .D(sreg[600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[599]) );
  DFF \sreg_reg[600]  ( .D(sreg[601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[600]) );
  DFF \sreg_reg[601]  ( .D(sreg[602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[601]) );
  DFF \sreg_reg[602]  ( .D(sreg[603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[602]) );
  DFF \sreg_reg[603]  ( .D(sreg[604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[603]) );
  DFF \sreg_reg[604]  ( .D(sreg[605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[604]) );
  DFF \sreg_reg[605]  ( .D(sreg[606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[605]) );
  DFF \sreg_reg[606]  ( .D(sreg[607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[606]) );
  DFF \sreg_reg[607]  ( .D(sreg[608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[607]) );
  DFF \sreg_reg[608]  ( .D(sreg[609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[608]) );
  DFF \sreg_reg[609]  ( .D(sreg[610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[609]) );
  DFF \sreg_reg[610]  ( .D(sreg[611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[610]) );
  DFF \sreg_reg[611]  ( .D(sreg[612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[611]) );
  DFF \sreg_reg[612]  ( .D(sreg[613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[612]) );
  DFF \sreg_reg[613]  ( .D(sreg[614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[613]) );
  DFF \sreg_reg[614]  ( .D(sreg[615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[614]) );
  DFF \sreg_reg[615]  ( .D(sreg[616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[615]) );
  DFF \sreg_reg[616]  ( .D(sreg[617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[616]) );
  DFF \sreg_reg[617]  ( .D(sreg[618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[617]) );
  DFF \sreg_reg[618]  ( .D(sreg[619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[618]) );
  DFF \sreg_reg[619]  ( .D(sreg[620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[619]) );
  DFF \sreg_reg[620]  ( .D(sreg[621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[620]) );
  DFF \sreg_reg[621]  ( .D(sreg[622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[621]) );
  DFF \sreg_reg[622]  ( .D(sreg[623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[622]) );
  DFF \sreg_reg[623]  ( .D(sreg[624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[623]) );
  DFF \sreg_reg[624]  ( .D(sreg[625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[624]) );
  DFF \sreg_reg[625]  ( .D(sreg[626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[625]) );
  DFF \sreg_reg[626]  ( .D(sreg[627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[626]) );
  DFF \sreg_reg[627]  ( .D(sreg[628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[627]) );
  DFF \sreg_reg[628]  ( .D(sreg[629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[628]) );
  DFF \sreg_reg[629]  ( .D(sreg[630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[629]) );
  DFF \sreg_reg[630]  ( .D(sreg[631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[630]) );
  DFF \sreg_reg[631]  ( .D(sreg[632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[631]) );
  DFF \sreg_reg[632]  ( .D(sreg[633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[632]) );
  DFF \sreg_reg[633]  ( .D(sreg[634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[633]) );
  DFF \sreg_reg[634]  ( .D(sreg[635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[634]) );
  DFF \sreg_reg[635]  ( .D(sreg[636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[635]) );
  DFF \sreg_reg[636]  ( .D(sreg[637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[636]) );
  DFF \sreg_reg[637]  ( .D(sreg[638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[637]) );
  DFF \sreg_reg[638]  ( .D(sreg[639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[638]) );
  DFF \sreg_reg[639]  ( .D(sreg[640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[639]) );
  DFF \sreg_reg[640]  ( .D(sreg[641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[640]) );
  DFF \sreg_reg[641]  ( .D(sreg[642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[641]) );
  DFF \sreg_reg[642]  ( .D(sreg[643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[642]) );
  DFF \sreg_reg[643]  ( .D(sreg[644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[643]) );
  DFF \sreg_reg[644]  ( .D(sreg[645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[644]) );
  DFF \sreg_reg[645]  ( .D(sreg[646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[645]) );
  DFF \sreg_reg[646]  ( .D(sreg[647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[646]) );
  DFF \sreg_reg[647]  ( .D(sreg[648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[647]) );
  DFF \sreg_reg[648]  ( .D(sreg[649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[648]) );
  DFF \sreg_reg[649]  ( .D(sreg[650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[649]) );
  DFF \sreg_reg[650]  ( .D(sreg[651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[650]) );
  DFF \sreg_reg[651]  ( .D(sreg[652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[651]) );
  DFF \sreg_reg[652]  ( .D(sreg[653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[652]) );
  DFF \sreg_reg[653]  ( .D(sreg[654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[653]) );
  DFF \sreg_reg[654]  ( .D(sreg[655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[654]) );
  DFF \sreg_reg[655]  ( .D(sreg[656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[655]) );
  DFF \sreg_reg[656]  ( .D(sreg[657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[656]) );
  DFF \sreg_reg[657]  ( .D(sreg[658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[657]) );
  DFF \sreg_reg[658]  ( .D(sreg[659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[658]) );
  DFF \sreg_reg[659]  ( .D(sreg[660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[659]) );
  DFF \sreg_reg[660]  ( .D(sreg[661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[660]) );
  DFF \sreg_reg[661]  ( .D(sreg[662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[661]) );
  DFF \sreg_reg[662]  ( .D(sreg[663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[662]) );
  DFF \sreg_reg[663]  ( .D(sreg[664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[663]) );
  DFF \sreg_reg[664]  ( .D(sreg[665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[664]) );
  DFF \sreg_reg[665]  ( .D(sreg[666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[665]) );
  DFF \sreg_reg[666]  ( .D(sreg[667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[666]) );
  DFF \sreg_reg[667]  ( .D(sreg[668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[667]) );
  DFF \sreg_reg[668]  ( .D(sreg[669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[668]) );
  DFF \sreg_reg[669]  ( .D(sreg[670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[669]) );
  DFF \sreg_reg[670]  ( .D(sreg[671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[670]) );
  DFF \sreg_reg[671]  ( .D(sreg[672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[671]) );
  DFF \sreg_reg[672]  ( .D(sreg[673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[672]) );
  DFF \sreg_reg[673]  ( .D(sreg[674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[673]) );
  DFF \sreg_reg[674]  ( .D(sreg[675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[674]) );
  DFF \sreg_reg[675]  ( .D(sreg[676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[675]) );
  DFF \sreg_reg[676]  ( .D(sreg[677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[676]) );
  DFF \sreg_reg[677]  ( .D(sreg[678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[677]) );
  DFF \sreg_reg[678]  ( .D(sreg[679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[678]) );
  DFF \sreg_reg[679]  ( .D(sreg[680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[679]) );
  DFF \sreg_reg[680]  ( .D(sreg[681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[680]) );
  DFF \sreg_reg[681]  ( .D(sreg[682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[681]) );
  DFF \sreg_reg[682]  ( .D(sreg[683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[682]) );
  DFF \sreg_reg[683]  ( .D(sreg[684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[683]) );
  DFF \sreg_reg[684]  ( .D(sreg[685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[684]) );
  DFF \sreg_reg[685]  ( .D(sreg[686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[685]) );
  DFF \sreg_reg[686]  ( .D(sreg[687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[686]) );
  DFF \sreg_reg[687]  ( .D(sreg[688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[687]) );
  DFF \sreg_reg[688]  ( .D(sreg[689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[688]) );
  DFF \sreg_reg[689]  ( .D(sreg[690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[689]) );
  DFF \sreg_reg[690]  ( .D(sreg[691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[690]) );
  DFF \sreg_reg[691]  ( .D(sreg[692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[691]) );
  DFF \sreg_reg[692]  ( .D(sreg[693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[692]) );
  DFF \sreg_reg[693]  ( .D(sreg[694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[693]) );
  DFF \sreg_reg[694]  ( .D(sreg[695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[694]) );
  DFF \sreg_reg[695]  ( .D(sreg[696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[695]) );
  DFF \sreg_reg[696]  ( .D(sreg[697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[696]) );
  DFF \sreg_reg[697]  ( .D(sreg[698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[697]) );
  DFF \sreg_reg[698]  ( .D(sreg[699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[698]) );
  DFF \sreg_reg[699]  ( .D(sreg[700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[699]) );
  DFF \sreg_reg[700]  ( .D(sreg[701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[700]) );
  DFF \sreg_reg[701]  ( .D(sreg[702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[701]) );
  DFF \sreg_reg[702]  ( .D(sreg[703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[702]) );
  DFF \sreg_reg[703]  ( .D(sreg[704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[703]) );
  DFF \sreg_reg[704]  ( .D(sreg[705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[704]) );
  DFF \sreg_reg[705]  ( .D(sreg[706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[705]) );
  DFF \sreg_reg[706]  ( .D(sreg[707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[706]) );
  DFF \sreg_reg[707]  ( .D(sreg[708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[707]) );
  DFF \sreg_reg[708]  ( .D(sreg[709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[708]) );
  DFF \sreg_reg[709]  ( .D(sreg[710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[709]) );
  DFF \sreg_reg[710]  ( .D(sreg[711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[710]) );
  DFF \sreg_reg[711]  ( .D(sreg[712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[711]) );
  DFF \sreg_reg[712]  ( .D(sreg[713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[712]) );
  DFF \sreg_reg[713]  ( .D(sreg[714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[713]) );
  DFF \sreg_reg[714]  ( .D(sreg[715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[714]) );
  DFF \sreg_reg[715]  ( .D(sreg[716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[715]) );
  DFF \sreg_reg[716]  ( .D(sreg[717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[716]) );
  DFF \sreg_reg[717]  ( .D(sreg[718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[717]) );
  DFF \sreg_reg[718]  ( .D(sreg[719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[718]) );
  DFF \sreg_reg[719]  ( .D(sreg[720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[719]) );
  DFF \sreg_reg[720]  ( .D(sreg[721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[720]) );
  DFF \sreg_reg[721]  ( .D(sreg[722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[721]) );
  DFF \sreg_reg[722]  ( .D(sreg[723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[722]) );
  DFF \sreg_reg[723]  ( .D(sreg[724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[723]) );
  DFF \sreg_reg[724]  ( .D(sreg[725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[724]) );
  DFF \sreg_reg[725]  ( .D(sreg[726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[725]) );
  DFF \sreg_reg[726]  ( .D(sreg[727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[726]) );
  DFF \sreg_reg[727]  ( .D(sreg[728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[727]) );
  DFF \sreg_reg[728]  ( .D(sreg[729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[728]) );
  DFF \sreg_reg[729]  ( .D(sreg[730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[729]) );
  DFF \sreg_reg[730]  ( .D(sreg[731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[730]) );
  DFF \sreg_reg[731]  ( .D(sreg[732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[731]) );
  DFF \sreg_reg[732]  ( .D(sreg[733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[732]) );
  DFF \sreg_reg[733]  ( .D(sreg[734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[733]) );
  DFF \sreg_reg[734]  ( .D(sreg[735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[734]) );
  DFF \sreg_reg[735]  ( .D(sreg[736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[735]) );
  DFF \sreg_reg[736]  ( .D(sreg[737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[736]) );
  DFF \sreg_reg[737]  ( .D(sreg[738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[737]) );
  DFF \sreg_reg[738]  ( .D(sreg[739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[738]) );
  DFF \sreg_reg[739]  ( .D(sreg[740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[739]) );
  DFF \sreg_reg[740]  ( .D(sreg[741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[740]) );
  DFF \sreg_reg[741]  ( .D(sreg[742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[741]) );
  DFF \sreg_reg[742]  ( .D(sreg[743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[742]) );
  DFF \sreg_reg[743]  ( .D(sreg[744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[743]) );
  DFF \sreg_reg[744]  ( .D(sreg[745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[744]) );
  DFF \sreg_reg[745]  ( .D(sreg[746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[745]) );
  DFF \sreg_reg[746]  ( .D(sreg[747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[746]) );
  DFF \sreg_reg[747]  ( .D(sreg[748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[747]) );
  DFF \sreg_reg[748]  ( .D(sreg[749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[748]) );
  DFF \sreg_reg[749]  ( .D(sreg[750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[749]) );
  DFF \sreg_reg[750]  ( .D(sreg[751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[750]) );
  DFF \sreg_reg[751]  ( .D(sreg[752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[751]) );
  DFF \sreg_reg[752]  ( .D(sreg[753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[752]) );
  DFF \sreg_reg[753]  ( .D(sreg[754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[753]) );
  DFF \sreg_reg[754]  ( .D(sreg[755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[754]) );
  DFF \sreg_reg[755]  ( .D(sreg[756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[755]) );
  DFF \sreg_reg[756]  ( .D(sreg[757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[756]) );
  DFF \sreg_reg[757]  ( .D(sreg[758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[757]) );
  DFF \sreg_reg[758]  ( .D(sreg[759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[758]) );
  DFF \sreg_reg[759]  ( .D(sreg[760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[759]) );
  DFF \sreg_reg[760]  ( .D(sreg[761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[760]) );
  DFF \sreg_reg[761]  ( .D(sreg[762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[761]) );
  DFF \sreg_reg[762]  ( .D(sreg[763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[762]) );
  DFF \sreg_reg[763]  ( .D(sreg[764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[763]) );
  DFF \sreg_reg[764]  ( .D(sreg[765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[764]) );
  DFF \sreg_reg[765]  ( .D(sreg[766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[765]) );
  DFF \sreg_reg[766]  ( .D(sreg[767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[766]) );
  DFF \sreg_reg[767]  ( .D(sreg[768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[767]) );
  DFF \sreg_reg[768]  ( .D(sreg[769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[768]) );
  DFF \sreg_reg[769]  ( .D(sreg[770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[769]) );
  DFF \sreg_reg[770]  ( .D(sreg[771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[770]) );
  DFF \sreg_reg[771]  ( .D(sreg[772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[771]) );
  DFF \sreg_reg[772]  ( .D(sreg[773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[772]) );
  DFF \sreg_reg[773]  ( .D(sreg[774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[773]) );
  DFF \sreg_reg[774]  ( .D(sreg[775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[774]) );
  DFF \sreg_reg[775]  ( .D(sreg[776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[775]) );
  DFF \sreg_reg[776]  ( .D(sreg[777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[776]) );
  DFF \sreg_reg[777]  ( .D(sreg[778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[777]) );
  DFF \sreg_reg[778]  ( .D(sreg[779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[778]) );
  DFF \sreg_reg[779]  ( .D(sreg[780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[779]) );
  DFF \sreg_reg[780]  ( .D(sreg[781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[780]) );
  DFF \sreg_reg[781]  ( .D(sreg[782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[781]) );
  DFF \sreg_reg[782]  ( .D(sreg[783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[782]) );
  DFF \sreg_reg[783]  ( .D(sreg[784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[783]) );
  DFF \sreg_reg[784]  ( .D(sreg[785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[784]) );
  DFF \sreg_reg[785]  ( .D(sreg[786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[785]) );
  DFF \sreg_reg[786]  ( .D(sreg[787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[786]) );
  DFF \sreg_reg[787]  ( .D(sreg[788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[787]) );
  DFF \sreg_reg[788]  ( .D(sreg[789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[788]) );
  DFF \sreg_reg[789]  ( .D(sreg[790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[789]) );
  DFF \sreg_reg[790]  ( .D(sreg[791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[790]) );
  DFF \sreg_reg[791]  ( .D(sreg[792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[791]) );
  DFF \sreg_reg[792]  ( .D(sreg[793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[792]) );
  DFF \sreg_reg[793]  ( .D(sreg[794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[793]) );
  DFF \sreg_reg[794]  ( .D(sreg[795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[794]) );
  DFF \sreg_reg[795]  ( .D(sreg[796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[795]) );
  DFF \sreg_reg[796]  ( .D(sreg[797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[796]) );
  DFF \sreg_reg[797]  ( .D(sreg[798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[797]) );
  DFF \sreg_reg[798]  ( .D(sreg[799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[798]) );
  DFF \sreg_reg[799]  ( .D(sreg[800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[799]) );
  DFF \sreg_reg[800]  ( .D(sreg[801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[800]) );
  DFF \sreg_reg[801]  ( .D(sreg[802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[801]) );
  DFF \sreg_reg[802]  ( .D(sreg[803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[802]) );
  DFF \sreg_reg[803]  ( .D(sreg[804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[803]) );
  DFF \sreg_reg[804]  ( .D(sreg[805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[804]) );
  DFF \sreg_reg[805]  ( .D(sreg[806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[805]) );
  DFF \sreg_reg[806]  ( .D(sreg[807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[806]) );
  DFF \sreg_reg[807]  ( .D(sreg[808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[807]) );
  DFF \sreg_reg[808]  ( .D(sreg[809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[808]) );
  DFF \sreg_reg[809]  ( .D(sreg[810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[809]) );
  DFF \sreg_reg[810]  ( .D(sreg[811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[810]) );
  DFF \sreg_reg[811]  ( .D(sreg[812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[811]) );
  DFF \sreg_reg[812]  ( .D(sreg[813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[812]) );
  DFF \sreg_reg[813]  ( .D(sreg[814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[813]) );
  DFF \sreg_reg[814]  ( .D(sreg[815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[814]) );
  DFF \sreg_reg[815]  ( .D(sreg[816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[815]) );
  DFF \sreg_reg[816]  ( .D(sreg[817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[816]) );
  DFF \sreg_reg[817]  ( .D(sreg[818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[817]) );
  DFF \sreg_reg[818]  ( .D(sreg[819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[818]) );
  DFF \sreg_reg[819]  ( .D(sreg[820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[819]) );
  DFF \sreg_reg[820]  ( .D(sreg[821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[820]) );
  DFF \sreg_reg[821]  ( .D(sreg[822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[821]) );
  DFF \sreg_reg[822]  ( .D(sreg[823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[822]) );
  DFF \sreg_reg[823]  ( .D(sreg[824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[823]) );
  DFF \sreg_reg[824]  ( .D(sreg[825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[824]) );
  DFF \sreg_reg[825]  ( .D(sreg[826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[825]) );
  DFF \sreg_reg[826]  ( .D(sreg[827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[826]) );
  DFF \sreg_reg[827]  ( .D(sreg[828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[827]) );
  DFF \sreg_reg[828]  ( .D(sreg[829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[828]) );
  DFF \sreg_reg[829]  ( .D(sreg[830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[829]) );
  DFF \sreg_reg[830]  ( .D(sreg[831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[830]) );
  DFF \sreg_reg[831]  ( .D(sreg[832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[831]) );
  DFF \sreg_reg[832]  ( .D(sreg[833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[832]) );
  DFF \sreg_reg[833]  ( .D(sreg[834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[833]) );
  DFF \sreg_reg[834]  ( .D(sreg[835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[834]) );
  DFF \sreg_reg[835]  ( .D(sreg[836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[835]) );
  DFF \sreg_reg[836]  ( .D(sreg[837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[836]) );
  DFF \sreg_reg[837]  ( .D(sreg[838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[837]) );
  DFF \sreg_reg[838]  ( .D(sreg[839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[838]) );
  DFF \sreg_reg[839]  ( .D(sreg[840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[839]) );
  DFF \sreg_reg[840]  ( .D(sreg[841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[840]) );
  DFF \sreg_reg[841]  ( .D(sreg[842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[841]) );
  DFF \sreg_reg[842]  ( .D(sreg[843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[842]) );
  DFF \sreg_reg[843]  ( .D(sreg[844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[843]) );
  DFF \sreg_reg[844]  ( .D(sreg[845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[844]) );
  DFF \sreg_reg[845]  ( .D(sreg[846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[845]) );
  DFF \sreg_reg[846]  ( .D(sreg[847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[846]) );
  DFF \sreg_reg[847]  ( .D(sreg[848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[847]) );
  DFF \sreg_reg[848]  ( .D(sreg[849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[848]) );
  DFF \sreg_reg[849]  ( .D(sreg[850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[849]) );
  DFF \sreg_reg[850]  ( .D(sreg[851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[850]) );
  DFF \sreg_reg[851]  ( .D(sreg[852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[851]) );
  DFF \sreg_reg[852]  ( .D(sreg[853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[852]) );
  DFF \sreg_reg[853]  ( .D(sreg[854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[853]) );
  DFF \sreg_reg[854]  ( .D(sreg[855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[854]) );
  DFF \sreg_reg[855]  ( .D(sreg[856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[855]) );
  DFF \sreg_reg[856]  ( .D(sreg[857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[856]) );
  DFF \sreg_reg[857]  ( .D(sreg[858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[857]) );
  DFF \sreg_reg[858]  ( .D(sreg[859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[858]) );
  DFF \sreg_reg[859]  ( .D(sreg[860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[859]) );
  DFF \sreg_reg[860]  ( .D(sreg[861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[860]) );
  DFF \sreg_reg[861]  ( .D(sreg[862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[861]) );
  DFF \sreg_reg[862]  ( .D(sreg[863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[862]) );
  DFF \sreg_reg[863]  ( .D(sreg[864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[863]) );
  DFF \sreg_reg[864]  ( .D(sreg[865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[864]) );
  DFF \sreg_reg[865]  ( .D(sreg[866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[865]) );
  DFF \sreg_reg[866]  ( .D(sreg[867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[866]) );
  DFF \sreg_reg[867]  ( .D(sreg[868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[867]) );
  DFF \sreg_reg[868]  ( .D(sreg[869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[868]) );
  DFF \sreg_reg[869]  ( .D(sreg[870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[869]) );
  DFF \sreg_reg[870]  ( .D(sreg[871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[870]) );
  DFF \sreg_reg[871]  ( .D(sreg[872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[871]) );
  DFF \sreg_reg[872]  ( .D(sreg[873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[872]) );
  DFF \sreg_reg[873]  ( .D(sreg[874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[873]) );
  DFF \sreg_reg[874]  ( .D(sreg[875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[874]) );
  DFF \sreg_reg[875]  ( .D(sreg[876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[875]) );
  DFF \sreg_reg[876]  ( .D(sreg[877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[876]) );
  DFF \sreg_reg[877]  ( .D(sreg[878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[877]) );
  DFF \sreg_reg[878]  ( .D(sreg[879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[878]) );
  DFF \sreg_reg[879]  ( .D(sreg[880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[879]) );
  DFF \sreg_reg[880]  ( .D(sreg[881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[880]) );
  DFF \sreg_reg[881]  ( .D(sreg[882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[881]) );
  DFF \sreg_reg[882]  ( .D(sreg[883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[882]) );
  DFF \sreg_reg[883]  ( .D(sreg[884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[883]) );
  DFF \sreg_reg[884]  ( .D(sreg[885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[884]) );
  DFF \sreg_reg[885]  ( .D(sreg[886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[885]) );
  DFF \sreg_reg[886]  ( .D(sreg[887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[886]) );
  DFF \sreg_reg[887]  ( .D(sreg[888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[887]) );
  DFF \sreg_reg[888]  ( .D(sreg[889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[888]) );
  DFF \sreg_reg[889]  ( .D(sreg[890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[889]) );
  DFF \sreg_reg[890]  ( .D(sreg[891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[890]) );
  DFF \sreg_reg[891]  ( .D(sreg[892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[891]) );
  DFF \sreg_reg[892]  ( .D(sreg[893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[892]) );
  DFF \sreg_reg[893]  ( .D(sreg[894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[893]) );
  DFF \sreg_reg[894]  ( .D(sreg[895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[894]) );
  DFF \sreg_reg[895]  ( .D(sreg[896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[895]) );
  DFF \sreg_reg[896]  ( .D(sreg[897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[896]) );
  DFF \sreg_reg[897]  ( .D(sreg[898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[897]) );
  DFF \sreg_reg[898]  ( .D(sreg[899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[898]) );
  DFF \sreg_reg[899]  ( .D(sreg[900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[899]) );
  DFF \sreg_reg[900]  ( .D(sreg[901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[900]) );
  DFF \sreg_reg[901]  ( .D(sreg[902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[901]) );
  DFF \sreg_reg[902]  ( .D(sreg[903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[902]) );
  DFF \sreg_reg[903]  ( .D(sreg[904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[903]) );
  DFF \sreg_reg[904]  ( .D(sreg[905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[904]) );
  DFF \sreg_reg[905]  ( .D(sreg[906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[905]) );
  DFF \sreg_reg[906]  ( .D(sreg[907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[906]) );
  DFF \sreg_reg[907]  ( .D(sreg[908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[907]) );
  DFF \sreg_reg[908]  ( .D(sreg[909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[908]) );
  DFF \sreg_reg[909]  ( .D(sreg[910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[909]) );
  DFF \sreg_reg[910]  ( .D(sreg[911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[910]) );
  DFF \sreg_reg[911]  ( .D(sreg[912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[911]) );
  DFF \sreg_reg[912]  ( .D(sreg[913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[912]) );
  DFF \sreg_reg[913]  ( .D(sreg[914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[913]) );
  DFF \sreg_reg[914]  ( .D(sreg[915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[914]) );
  DFF \sreg_reg[915]  ( .D(sreg[916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[915]) );
  DFF \sreg_reg[916]  ( .D(sreg[917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[916]) );
  DFF \sreg_reg[917]  ( .D(sreg[918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[917]) );
  DFF \sreg_reg[918]  ( .D(sreg[919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[918]) );
  DFF \sreg_reg[919]  ( .D(sreg[920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[919]) );
  DFF \sreg_reg[920]  ( .D(sreg[921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[920]) );
  DFF \sreg_reg[921]  ( .D(sreg[922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[921]) );
  DFF \sreg_reg[922]  ( .D(sreg[923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[922]) );
  DFF \sreg_reg[923]  ( .D(sreg[924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[923]) );
  DFF \sreg_reg[924]  ( .D(sreg[925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[924]) );
  DFF \sreg_reg[925]  ( .D(sreg[926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[925]) );
  DFF \sreg_reg[926]  ( .D(sreg[927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[926]) );
  DFF \sreg_reg[927]  ( .D(sreg[928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[927]) );
  DFF \sreg_reg[928]  ( .D(sreg[929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[928]) );
  DFF \sreg_reg[929]  ( .D(sreg[930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[929]) );
  DFF \sreg_reg[930]  ( .D(sreg[931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[930]) );
  DFF \sreg_reg[931]  ( .D(sreg[932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[931]) );
  DFF \sreg_reg[932]  ( .D(sreg[933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[932]) );
  DFF \sreg_reg[933]  ( .D(sreg[934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[933]) );
  DFF \sreg_reg[934]  ( .D(sreg[935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[934]) );
  DFF \sreg_reg[935]  ( .D(sreg[936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[935]) );
  DFF \sreg_reg[936]  ( .D(sreg[937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[936]) );
  DFF \sreg_reg[937]  ( .D(sreg[938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[937]) );
  DFF \sreg_reg[938]  ( .D(sreg[939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[938]) );
  DFF \sreg_reg[939]  ( .D(sreg[940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[939]) );
  DFF \sreg_reg[940]  ( .D(sreg[941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[940]) );
  DFF \sreg_reg[941]  ( .D(sreg[942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[941]) );
  DFF \sreg_reg[942]  ( .D(sreg[943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[942]) );
  DFF \sreg_reg[943]  ( .D(sreg[944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[943]) );
  DFF \sreg_reg[944]  ( .D(sreg[945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[944]) );
  DFF \sreg_reg[945]  ( .D(sreg[946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[945]) );
  DFF \sreg_reg[946]  ( .D(sreg[947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[946]) );
  DFF \sreg_reg[947]  ( .D(sreg[948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[947]) );
  DFF \sreg_reg[948]  ( .D(sreg[949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[948]) );
  DFF \sreg_reg[949]  ( .D(sreg[950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[949]) );
  DFF \sreg_reg[950]  ( .D(sreg[951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[950]) );
  DFF \sreg_reg[951]  ( .D(sreg[952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[951]) );
  DFF \sreg_reg[952]  ( .D(sreg[953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[952]) );
  DFF \sreg_reg[953]  ( .D(sreg[954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[953]) );
  DFF \sreg_reg[954]  ( .D(sreg[955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[954]) );
  DFF \sreg_reg[955]  ( .D(sreg[956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[955]) );
  DFF \sreg_reg[956]  ( .D(sreg[957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[956]) );
  DFF \sreg_reg[957]  ( .D(sreg[958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[957]) );
  DFF \sreg_reg[958]  ( .D(sreg[959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[958]) );
  DFF \sreg_reg[959]  ( .D(sreg[960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[959]) );
  DFF \sreg_reg[960]  ( .D(sreg[961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[960]) );
  DFF \sreg_reg[961]  ( .D(sreg[962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[961]) );
  DFF \sreg_reg[962]  ( .D(sreg[963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[962]) );
  DFF \sreg_reg[963]  ( .D(sreg[964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[963]) );
  DFF \sreg_reg[964]  ( .D(sreg[965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[964]) );
  DFF \sreg_reg[965]  ( .D(sreg[966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[965]) );
  DFF \sreg_reg[966]  ( .D(sreg[967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[966]) );
  DFF \sreg_reg[967]  ( .D(sreg[968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[967]) );
  DFF \sreg_reg[968]  ( .D(sreg[969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[968]) );
  DFF \sreg_reg[969]  ( .D(sreg[970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[969]) );
  DFF \sreg_reg[970]  ( .D(sreg[971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[970]) );
  DFF \sreg_reg[971]  ( .D(sreg[972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[971]) );
  DFF \sreg_reg[972]  ( .D(sreg[973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[972]) );
  DFF \sreg_reg[973]  ( .D(sreg[974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[973]) );
  DFF \sreg_reg[974]  ( .D(sreg[975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[974]) );
  DFF \sreg_reg[975]  ( .D(sreg[976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[975]) );
  DFF \sreg_reg[976]  ( .D(sreg[977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[976]) );
  DFF \sreg_reg[977]  ( .D(sreg[978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[977]) );
  DFF \sreg_reg[978]  ( .D(sreg[979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[978]) );
  DFF \sreg_reg[979]  ( .D(sreg[980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[979]) );
  DFF \sreg_reg[980]  ( .D(sreg[981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[980]) );
  DFF \sreg_reg[981]  ( .D(sreg[982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[981]) );
  DFF \sreg_reg[982]  ( .D(sreg[983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[982]) );
  DFF \sreg_reg[983]  ( .D(sreg[984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[983]) );
  DFF \sreg_reg[984]  ( .D(sreg[985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[984]) );
  DFF \sreg_reg[985]  ( .D(sreg[986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[985]) );
  DFF \sreg_reg[986]  ( .D(sreg[987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[986]) );
  DFF \sreg_reg[987]  ( .D(sreg[988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[987]) );
  DFF \sreg_reg[988]  ( .D(sreg[989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[988]) );
  DFF \sreg_reg[989]  ( .D(sreg[990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[989]) );
  DFF \sreg_reg[990]  ( .D(sreg[991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[990]) );
  DFF \sreg_reg[991]  ( .D(sreg[992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[991]) );
  DFF \sreg_reg[992]  ( .D(sreg[993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[992]) );
  DFF \sreg_reg[993]  ( .D(sreg[994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[993]) );
  DFF \sreg_reg[994]  ( .D(sreg[995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[994]) );
  DFF \sreg_reg[995]  ( .D(sreg[996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[995]) );
  DFF \sreg_reg[996]  ( .D(sreg[997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[996]) );
  DFF \sreg_reg[997]  ( .D(sreg[998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[997]) );
  DFF \sreg_reg[998]  ( .D(sreg[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[998]) );
  DFF \sreg_reg[999]  ( .D(sreg[1000]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[999]) );
  DFF \sreg_reg[1000]  ( .D(sreg[1001]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1000]) );
  DFF \sreg_reg[1001]  ( .D(sreg[1002]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1001]) );
  DFF \sreg_reg[1002]  ( .D(sreg[1003]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1002]) );
  DFF \sreg_reg[1003]  ( .D(sreg[1004]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1003]) );
  DFF \sreg_reg[1004]  ( .D(sreg[1005]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1004]) );
  DFF \sreg_reg[1005]  ( .D(sreg[1006]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1005]) );
  DFF \sreg_reg[1006]  ( .D(sreg[1007]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1006]) );
  DFF \sreg_reg[1007]  ( .D(sreg[1008]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1007]) );
  DFF \sreg_reg[1008]  ( .D(sreg[1009]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1008]) );
  DFF \sreg_reg[1009]  ( .D(sreg[1010]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1009]) );
  DFF \sreg_reg[1010]  ( .D(sreg[1011]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1010]) );
  DFF \sreg_reg[1011]  ( .D(sreg[1012]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1011]) );
  DFF \sreg_reg[1012]  ( .D(sreg[1013]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1012]) );
  DFF \sreg_reg[1013]  ( .D(sreg[1014]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1013]) );
  DFF \sreg_reg[1014]  ( .D(sreg[1015]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1014]) );
  DFF \sreg_reg[1015]  ( .D(sreg[1016]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1015]) );
  DFF \sreg_reg[1016]  ( .D(sreg[1017]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1016]) );
  DFF \sreg_reg[1017]  ( .D(sreg[1018]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1017]) );
  DFF \sreg_reg[1018]  ( .D(sreg[1019]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1018]) );
  DFF \sreg_reg[1019]  ( .D(sreg[1020]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1019]) );
  DFF \sreg_reg[1020]  ( .D(sreg[1021]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1020]) );
  DFF \sreg_reg[1021]  ( .D(sreg[1022]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1021]) );
  DFF \sreg_reg[1022]  ( .D(o[1023]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1022]) );
  DFF \sreg_reg[1023]  ( .D(o[1024]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1023]) );
  DFF \sreg_reg[1024]  ( .D(o[1025]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1024]) );
  DFF \sreg_reg[1025]  ( .D(o[1026]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1025]) );
  DFF \sreg_reg[1026]  ( .D(o[1027]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1026]) );
  DFF \sreg_reg[1027]  ( .D(o[1028]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1027]) );
  DFF \sreg_reg[1028]  ( .D(o[1029]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1028]) );
  DFF \sreg_reg[1029]  ( .D(o[1030]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1029]) );
  DFF \sreg_reg[1030]  ( .D(o[1031]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1030]) );
  DFF \sreg_reg[1031]  ( .D(o[1032]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1031]) );
  DFF \sreg_reg[1032]  ( .D(o[1033]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1032]) );
  DFF \sreg_reg[1033]  ( .D(o[1034]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1033]) );
  DFF \sreg_reg[1034]  ( .D(o[1035]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1034]) );
  DFF \sreg_reg[1035]  ( .D(o[1036]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1035]) );
  DFF \sreg_reg[1036]  ( .D(o[1037]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1036]) );
  DFF \sreg_reg[1037]  ( .D(o[1038]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1037]) );
  DFF \sreg_reg[1038]  ( .D(o[1039]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1038]) );
  DFF \sreg_reg[1039]  ( .D(o[1040]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1039]) );
  DFF \sreg_reg[1040]  ( .D(o[1041]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1040]) );
  DFF \sreg_reg[1041]  ( .D(o[1042]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1041]) );
  DFF \sreg_reg[1042]  ( .D(o[1043]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1042]) );
  DFF \sreg_reg[1043]  ( .D(o[1044]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1043]) );
  DFF \sreg_reg[1044]  ( .D(o[1045]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1044]) );
  DFF \sreg_reg[1045]  ( .D(o[1046]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1045]) );
  DFF \sreg_reg[1046]  ( .D(o[1047]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1046]) );
  DFF \sreg_reg[1047]  ( .D(o[1048]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1047]) );
  DFF \sreg_reg[1048]  ( .D(o[1049]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1048]) );
  DFF \sreg_reg[1049]  ( .D(o[1050]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1049]) );
  DFF \sreg_reg[1050]  ( .D(o[1051]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1050]) );
  DFF \sreg_reg[1051]  ( .D(o[1052]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1051]) );
  DFF \sreg_reg[1052]  ( .D(o[1053]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1052]) );
  DFF \sreg_reg[1053]  ( .D(o[1054]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1053]) );
  DFF \sreg_reg[1054]  ( .D(o[1055]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1054]) );
  DFF \sreg_reg[1055]  ( .D(o[1056]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1055]) );
  DFF \sreg_reg[1056]  ( .D(o[1057]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1056]) );
  DFF \sreg_reg[1057]  ( .D(o[1058]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1057]) );
  DFF \sreg_reg[1058]  ( .D(o[1059]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1058]) );
  DFF \sreg_reg[1059]  ( .D(o[1060]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1059]) );
  DFF \sreg_reg[1060]  ( .D(o[1061]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1060]) );
  DFF \sreg_reg[1061]  ( .D(o[1062]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1061]) );
  DFF \sreg_reg[1062]  ( .D(o[1063]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1062]) );
  DFF \sreg_reg[1063]  ( .D(o[1064]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1063]) );
  DFF \sreg_reg[1064]  ( .D(o[1065]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1064]) );
  DFF \sreg_reg[1065]  ( .D(o[1066]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1065]) );
  DFF \sreg_reg[1066]  ( .D(o[1067]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1066]) );
  DFF \sreg_reg[1067]  ( .D(o[1068]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1067]) );
  DFF \sreg_reg[1068]  ( .D(o[1069]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1068]) );
  DFF \sreg_reg[1069]  ( .D(o[1070]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1069]) );
  DFF \sreg_reg[1070]  ( .D(o[1071]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1070]) );
  DFF \sreg_reg[1071]  ( .D(o[1072]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1071]) );
  DFF \sreg_reg[1072]  ( .D(o[1073]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1072]) );
  DFF \sreg_reg[1073]  ( .D(o[1074]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1073]) );
  DFF \sreg_reg[1074]  ( .D(o[1075]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1074]) );
  DFF \sreg_reg[1075]  ( .D(o[1076]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1075]) );
  DFF \sreg_reg[1076]  ( .D(o[1077]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1076]) );
  DFF \sreg_reg[1077]  ( .D(o[1078]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1077]) );
  DFF \sreg_reg[1078]  ( .D(o[1079]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1078]) );
  DFF \sreg_reg[1079]  ( .D(o[1080]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1079]) );
  DFF \sreg_reg[1080]  ( .D(o[1081]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1080]) );
  DFF \sreg_reg[1081]  ( .D(o[1082]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1081]) );
  DFF \sreg_reg[1082]  ( .D(o[1083]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1082]) );
  DFF \sreg_reg[1083]  ( .D(o[1084]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1083]) );
  DFF \sreg_reg[1084]  ( .D(o[1085]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1084]) );
  DFF \sreg_reg[1085]  ( .D(o[1086]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1085]) );
  DFF \sreg_reg[1086]  ( .D(o[1087]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1086]) );
  DFF \sreg_reg[1087]  ( .D(o[1088]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1087]) );
  DFF \sreg_reg[1088]  ( .D(o[1089]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1088]) );
  DFF \sreg_reg[1089]  ( .D(o[1090]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1089]) );
  DFF \sreg_reg[1090]  ( .D(o[1091]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1090]) );
  DFF \sreg_reg[1091]  ( .D(o[1092]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1091]) );
  DFF \sreg_reg[1092]  ( .D(o[1093]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1092]) );
  DFF \sreg_reg[1093]  ( .D(o[1094]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1093]) );
  DFF \sreg_reg[1094]  ( .D(o[1095]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1094]) );
  DFF \sreg_reg[1095]  ( .D(o[1096]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1095]) );
  DFF \sreg_reg[1096]  ( .D(o[1097]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1096]) );
  DFF \sreg_reg[1097]  ( .D(o[1098]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1097]) );
  DFF \sreg_reg[1098]  ( .D(o[1099]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1098]) );
  DFF \sreg_reg[1099]  ( .D(o[1100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1099]) );
  DFF \sreg_reg[1100]  ( .D(o[1101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1100]) );
  DFF \sreg_reg[1101]  ( .D(o[1102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1101]) );
  DFF \sreg_reg[1102]  ( .D(o[1103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1102]) );
  DFF \sreg_reg[1103]  ( .D(o[1104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1103]) );
  DFF \sreg_reg[1104]  ( .D(o[1105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1104]) );
  DFF \sreg_reg[1105]  ( .D(o[1106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1105]) );
  DFF \sreg_reg[1106]  ( .D(o[1107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1106]) );
  DFF \sreg_reg[1107]  ( .D(o[1108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1107]) );
  DFF \sreg_reg[1108]  ( .D(o[1109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1108]) );
  DFF \sreg_reg[1109]  ( .D(o[1110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1109]) );
  DFF \sreg_reg[1110]  ( .D(o[1111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1110]) );
  DFF \sreg_reg[1111]  ( .D(o[1112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1111]) );
  DFF \sreg_reg[1112]  ( .D(o[1113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1112]) );
  DFF \sreg_reg[1113]  ( .D(o[1114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1113]) );
  DFF \sreg_reg[1114]  ( .D(o[1115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1114]) );
  DFF \sreg_reg[1115]  ( .D(o[1116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1115]) );
  DFF \sreg_reg[1116]  ( .D(o[1117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1116]) );
  DFF \sreg_reg[1117]  ( .D(o[1118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1117]) );
  DFF \sreg_reg[1118]  ( .D(o[1119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1118]) );
  DFF \sreg_reg[1119]  ( .D(o[1120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1119]) );
  DFF \sreg_reg[1120]  ( .D(o[1121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1120]) );
  DFF \sreg_reg[1121]  ( .D(o[1122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1121]) );
  DFF \sreg_reg[1122]  ( .D(o[1123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1122]) );
  DFF \sreg_reg[1123]  ( .D(o[1124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1123]) );
  DFF \sreg_reg[1124]  ( .D(o[1125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1124]) );
  DFF \sreg_reg[1125]  ( .D(o[1126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1125]) );
  DFF \sreg_reg[1126]  ( .D(o[1127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1126]) );
  DFF \sreg_reg[1127]  ( .D(o[1128]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1127]) );
  DFF \sreg_reg[1128]  ( .D(o[1129]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1128]) );
  DFF \sreg_reg[1129]  ( .D(o[1130]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1129]) );
  DFF \sreg_reg[1130]  ( .D(o[1131]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1130]) );
  DFF \sreg_reg[1131]  ( .D(o[1132]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1131]) );
  DFF \sreg_reg[1132]  ( .D(o[1133]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1132]) );
  DFF \sreg_reg[1133]  ( .D(o[1134]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1133]) );
  DFF \sreg_reg[1134]  ( .D(o[1135]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1134]) );
  DFF \sreg_reg[1135]  ( .D(o[1136]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1135]) );
  DFF \sreg_reg[1136]  ( .D(o[1137]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1136]) );
  DFF \sreg_reg[1137]  ( .D(o[1138]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1137]) );
  DFF \sreg_reg[1138]  ( .D(o[1139]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1138]) );
  DFF \sreg_reg[1139]  ( .D(o[1140]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1139]) );
  DFF \sreg_reg[1140]  ( .D(o[1141]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1140]) );
  DFF \sreg_reg[1141]  ( .D(o[1142]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1141]) );
  DFF \sreg_reg[1142]  ( .D(o[1143]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1142]) );
  DFF \sreg_reg[1143]  ( .D(o[1144]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1143]) );
  DFF \sreg_reg[1144]  ( .D(o[1145]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1144]) );
  DFF \sreg_reg[1145]  ( .D(o[1146]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1145]) );
  DFF \sreg_reg[1146]  ( .D(o[1147]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1146]) );
  DFF \sreg_reg[1147]  ( .D(o[1148]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1147]) );
  DFF \sreg_reg[1148]  ( .D(o[1149]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1148]) );
  DFF \sreg_reg[1149]  ( .D(o[1150]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1149]) );
  DFF \sreg_reg[1150]  ( .D(o[1151]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1150]) );
  DFF \sreg_reg[1151]  ( .D(o[1152]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1151]) );
  DFF \sreg_reg[1152]  ( .D(o[1153]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1152]) );
  DFF \sreg_reg[1153]  ( .D(o[1154]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1153]) );
  DFF \sreg_reg[1154]  ( .D(o[1155]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1154]) );
  DFF \sreg_reg[1155]  ( .D(o[1156]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1155]) );
  DFF \sreg_reg[1156]  ( .D(o[1157]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1156]) );
  DFF \sreg_reg[1157]  ( .D(o[1158]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1157]) );
  DFF \sreg_reg[1158]  ( .D(o[1159]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1158]) );
  DFF \sreg_reg[1159]  ( .D(o[1160]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1159]) );
  DFF \sreg_reg[1160]  ( .D(o[1161]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1160]) );
  DFF \sreg_reg[1161]  ( .D(o[1162]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1161]) );
  DFF \sreg_reg[1162]  ( .D(o[1163]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1162]) );
  DFF \sreg_reg[1163]  ( .D(o[1164]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1163]) );
  DFF \sreg_reg[1164]  ( .D(o[1165]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1164]) );
  DFF \sreg_reg[1165]  ( .D(o[1166]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1165]) );
  DFF \sreg_reg[1166]  ( .D(o[1167]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1166]) );
  DFF \sreg_reg[1167]  ( .D(o[1168]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1167]) );
  DFF \sreg_reg[1168]  ( .D(o[1169]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1168]) );
  DFF \sreg_reg[1169]  ( .D(o[1170]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1169]) );
  DFF \sreg_reg[1170]  ( .D(o[1171]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1170]) );
  DFF \sreg_reg[1171]  ( .D(o[1172]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1171]) );
  DFF \sreg_reg[1172]  ( .D(o[1173]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1172]) );
  DFF \sreg_reg[1173]  ( .D(o[1174]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1173]) );
  DFF \sreg_reg[1174]  ( .D(o[1175]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1174]) );
  DFF \sreg_reg[1175]  ( .D(o[1176]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1175]) );
  DFF \sreg_reg[1176]  ( .D(o[1177]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1176]) );
  DFF \sreg_reg[1177]  ( .D(o[1178]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1177]) );
  DFF \sreg_reg[1178]  ( .D(o[1179]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1178]) );
  DFF \sreg_reg[1179]  ( .D(o[1180]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1179]) );
  DFF \sreg_reg[1180]  ( .D(o[1181]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1180]) );
  DFF \sreg_reg[1181]  ( .D(o[1182]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1181]) );
  DFF \sreg_reg[1182]  ( .D(o[1183]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1182]) );
  DFF \sreg_reg[1183]  ( .D(o[1184]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1183]) );
  DFF \sreg_reg[1184]  ( .D(o[1185]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1184]) );
  DFF \sreg_reg[1185]  ( .D(o[1186]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1185]) );
  DFF \sreg_reg[1186]  ( .D(o[1187]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1186]) );
  DFF \sreg_reg[1187]  ( .D(o[1188]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1187]) );
  DFF \sreg_reg[1188]  ( .D(o[1189]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1188]) );
  DFF \sreg_reg[1189]  ( .D(o[1190]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1189]) );
  DFF \sreg_reg[1190]  ( .D(o[1191]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1190]) );
  DFF \sreg_reg[1191]  ( .D(o[1192]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1191]) );
  DFF \sreg_reg[1192]  ( .D(o[1193]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1192]) );
  DFF \sreg_reg[1193]  ( .D(o[1194]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1193]) );
  DFF \sreg_reg[1194]  ( .D(o[1195]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1194]) );
  DFF \sreg_reg[1195]  ( .D(o[1196]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1195]) );
  DFF \sreg_reg[1196]  ( .D(o[1197]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1196]) );
  DFF \sreg_reg[1197]  ( .D(o[1198]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1197]) );
  DFF \sreg_reg[1198]  ( .D(o[1199]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1198]) );
  DFF \sreg_reg[1199]  ( .D(o[1200]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1199]) );
  DFF \sreg_reg[1200]  ( .D(o[1201]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1200]) );
  DFF \sreg_reg[1201]  ( .D(o[1202]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1201]) );
  DFF \sreg_reg[1202]  ( .D(o[1203]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1202]) );
  DFF \sreg_reg[1203]  ( .D(o[1204]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1203]) );
  DFF \sreg_reg[1204]  ( .D(o[1205]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1204]) );
  DFF \sreg_reg[1205]  ( .D(o[1206]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1205]) );
  DFF \sreg_reg[1206]  ( .D(o[1207]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1206]) );
  DFF \sreg_reg[1207]  ( .D(o[1208]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1207]) );
  DFF \sreg_reg[1208]  ( .D(o[1209]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1208]) );
  DFF \sreg_reg[1209]  ( .D(o[1210]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1209]) );
  DFF \sreg_reg[1210]  ( .D(o[1211]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1210]) );
  DFF \sreg_reg[1211]  ( .D(o[1212]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1211]) );
  DFF \sreg_reg[1212]  ( .D(o[1213]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1212]) );
  DFF \sreg_reg[1213]  ( .D(o[1214]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1213]) );
  DFF \sreg_reg[1214]  ( .D(o[1215]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1214]) );
  DFF \sreg_reg[1215]  ( .D(o[1216]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1215]) );
  DFF \sreg_reg[1216]  ( .D(o[1217]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1216]) );
  DFF \sreg_reg[1217]  ( .D(o[1218]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1217]) );
  DFF \sreg_reg[1218]  ( .D(o[1219]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1218]) );
  DFF \sreg_reg[1219]  ( .D(o[1220]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1219]) );
  DFF \sreg_reg[1220]  ( .D(o[1221]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1220]) );
  DFF \sreg_reg[1221]  ( .D(o[1222]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1221]) );
  DFF \sreg_reg[1222]  ( .D(o[1223]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1222]) );
  DFF \sreg_reg[1223]  ( .D(o[1224]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1223]) );
  DFF \sreg_reg[1224]  ( .D(o[1225]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1224]) );
  DFF \sreg_reg[1225]  ( .D(o[1226]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1225]) );
  DFF \sreg_reg[1226]  ( .D(o[1227]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1226]) );
  DFF \sreg_reg[1227]  ( .D(o[1228]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1227]) );
  DFF \sreg_reg[1228]  ( .D(o[1229]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1228]) );
  DFF \sreg_reg[1229]  ( .D(o[1230]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1229]) );
  DFF \sreg_reg[1230]  ( .D(o[1231]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1230]) );
  DFF \sreg_reg[1231]  ( .D(o[1232]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1231]) );
  DFF \sreg_reg[1232]  ( .D(o[1233]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1232]) );
  DFF \sreg_reg[1233]  ( .D(o[1234]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1233]) );
  DFF \sreg_reg[1234]  ( .D(o[1235]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1234]) );
  DFF \sreg_reg[1235]  ( .D(o[1236]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1235]) );
  DFF \sreg_reg[1236]  ( .D(o[1237]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1236]) );
  DFF \sreg_reg[1237]  ( .D(o[1238]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1237]) );
  DFF \sreg_reg[1238]  ( .D(o[1239]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1238]) );
  DFF \sreg_reg[1239]  ( .D(o[1240]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1239]) );
  DFF \sreg_reg[1240]  ( .D(o[1241]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1240]) );
  DFF \sreg_reg[1241]  ( .D(o[1242]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1241]) );
  DFF \sreg_reg[1242]  ( .D(o[1243]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1242]) );
  DFF \sreg_reg[1243]  ( .D(o[1244]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1243]) );
  DFF \sreg_reg[1244]  ( .D(o[1245]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1244]) );
  DFF \sreg_reg[1245]  ( .D(o[1246]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1245]) );
  DFF \sreg_reg[1246]  ( .D(o[1247]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1246]) );
  DFF \sreg_reg[1247]  ( .D(o[1248]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1247]) );
  DFF \sreg_reg[1248]  ( .D(o[1249]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1248]) );
  DFF \sreg_reg[1249]  ( .D(o[1250]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1249]) );
  DFF \sreg_reg[1250]  ( .D(o[1251]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1250]) );
  DFF \sreg_reg[1251]  ( .D(o[1252]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1251]) );
  DFF \sreg_reg[1252]  ( .D(o[1253]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1252]) );
  DFF \sreg_reg[1253]  ( .D(o[1254]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1253]) );
  DFF \sreg_reg[1254]  ( .D(o[1255]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1254]) );
  DFF \sreg_reg[1255]  ( .D(o[1256]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1255]) );
  DFF \sreg_reg[1256]  ( .D(o[1257]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1256]) );
  DFF \sreg_reg[1257]  ( .D(o[1258]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1257]) );
  DFF \sreg_reg[1258]  ( .D(o[1259]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1258]) );
  DFF \sreg_reg[1259]  ( .D(o[1260]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1259]) );
  DFF \sreg_reg[1260]  ( .D(o[1261]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1260]) );
  DFF \sreg_reg[1261]  ( .D(o[1262]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1261]) );
  DFF \sreg_reg[1262]  ( .D(o[1263]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1262]) );
  DFF \sreg_reg[1263]  ( .D(o[1264]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1263]) );
  DFF \sreg_reg[1264]  ( .D(o[1265]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1264]) );
  DFF \sreg_reg[1265]  ( .D(o[1266]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1265]) );
  DFF \sreg_reg[1266]  ( .D(o[1267]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1266]) );
  DFF \sreg_reg[1267]  ( .D(o[1268]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1267]) );
  DFF \sreg_reg[1268]  ( .D(o[1269]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1268]) );
  DFF \sreg_reg[1269]  ( .D(o[1270]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1269]) );
  DFF \sreg_reg[1270]  ( .D(o[1271]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1270]) );
  DFF \sreg_reg[1271]  ( .D(o[1272]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1271]) );
  DFF \sreg_reg[1272]  ( .D(o[1273]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1272]) );
  DFF \sreg_reg[1273]  ( .D(o[1274]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1273]) );
  DFF \sreg_reg[1274]  ( .D(o[1275]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1274]) );
  DFF \sreg_reg[1275]  ( .D(o[1276]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1275]) );
  DFF \sreg_reg[1276]  ( .D(o[1277]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1276]) );
  DFF \sreg_reg[1277]  ( .D(o[1278]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1277]) );
  DFF \sreg_reg[1278]  ( .D(o[1279]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1278]) );
  DFF \sreg_reg[1279]  ( .D(o[1280]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1279]) );
  DFF \sreg_reg[1280]  ( .D(o[1281]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1280]) );
  DFF \sreg_reg[1281]  ( .D(o[1282]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1281]) );
  DFF \sreg_reg[1282]  ( .D(o[1283]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1282]) );
  DFF \sreg_reg[1283]  ( .D(o[1284]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1283]) );
  DFF \sreg_reg[1284]  ( .D(o[1285]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1284]) );
  DFF \sreg_reg[1285]  ( .D(o[1286]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1285]) );
  DFF \sreg_reg[1286]  ( .D(o[1287]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1286]) );
  DFF \sreg_reg[1287]  ( .D(o[1288]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1287]) );
  DFF \sreg_reg[1288]  ( .D(o[1289]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1288]) );
  DFF \sreg_reg[1289]  ( .D(o[1290]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1289]) );
  DFF \sreg_reg[1290]  ( .D(o[1291]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1290]) );
  DFF \sreg_reg[1291]  ( .D(o[1292]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1291]) );
  DFF \sreg_reg[1292]  ( .D(o[1293]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1292]) );
  DFF \sreg_reg[1293]  ( .D(o[1294]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1293]) );
  DFF \sreg_reg[1294]  ( .D(o[1295]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1294]) );
  DFF \sreg_reg[1295]  ( .D(o[1296]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1295]) );
  DFF \sreg_reg[1296]  ( .D(o[1297]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1296]) );
  DFF \sreg_reg[1297]  ( .D(o[1298]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1297]) );
  DFF \sreg_reg[1298]  ( .D(o[1299]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1298]) );
  DFF \sreg_reg[1299]  ( .D(o[1300]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1299]) );
  DFF \sreg_reg[1300]  ( .D(o[1301]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1300]) );
  DFF \sreg_reg[1301]  ( .D(o[1302]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1301]) );
  DFF \sreg_reg[1302]  ( .D(o[1303]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1302]) );
  DFF \sreg_reg[1303]  ( .D(o[1304]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1303]) );
  DFF \sreg_reg[1304]  ( .D(o[1305]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1304]) );
  DFF \sreg_reg[1305]  ( .D(o[1306]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1305]) );
  DFF \sreg_reg[1306]  ( .D(o[1307]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1306]) );
  DFF \sreg_reg[1307]  ( .D(o[1308]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1307]) );
  DFF \sreg_reg[1308]  ( .D(o[1309]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1308]) );
  DFF \sreg_reg[1309]  ( .D(o[1310]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1309]) );
  DFF \sreg_reg[1310]  ( .D(o[1311]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1310]) );
  DFF \sreg_reg[1311]  ( .D(o[1312]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1311]) );
  DFF \sreg_reg[1312]  ( .D(o[1313]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1312]) );
  DFF \sreg_reg[1313]  ( .D(o[1314]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1313]) );
  DFF \sreg_reg[1314]  ( .D(o[1315]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1314]) );
  DFF \sreg_reg[1315]  ( .D(o[1316]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1315]) );
  DFF \sreg_reg[1316]  ( .D(o[1317]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1316]) );
  DFF \sreg_reg[1317]  ( .D(o[1318]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1317]) );
  DFF \sreg_reg[1318]  ( .D(o[1319]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1318]) );
  DFF \sreg_reg[1319]  ( .D(o[1320]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1319]) );
  DFF \sreg_reg[1320]  ( .D(o[1321]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1320]) );
  DFF \sreg_reg[1321]  ( .D(o[1322]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1321]) );
  DFF \sreg_reg[1322]  ( .D(o[1323]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1322]) );
  DFF \sreg_reg[1323]  ( .D(o[1324]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1323]) );
  DFF \sreg_reg[1324]  ( .D(o[1325]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1324]) );
  DFF \sreg_reg[1325]  ( .D(o[1326]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1325]) );
  DFF \sreg_reg[1326]  ( .D(o[1327]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1326]) );
  DFF \sreg_reg[1327]  ( .D(o[1328]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1327]) );
  DFF \sreg_reg[1328]  ( .D(o[1329]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1328]) );
  DFF \sreg_reg[1329]  ( .D(o[1330]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1329]) );
  DFF \sreg_reg[1330]  ( .D(o[1331]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1330]) );
  DFF \sreg_reg[1331]  ( .D(o[1332]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1331]) );
  DFF \sreg_reg[1332]  ( .D(o[1333]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1332]) );
  DFF \sreg_reg[1333]  ( .D(o[1334]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1333]) );
  DFF \sreg_reg[1334]  ( .D(o[1335]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1334]) );
  DFF \sreg_reg[1335]  ( .D(o[1336]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1335]) );
  DFF \sreg_reg[1336]  ( .D(o[1337]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1336]) );
  DFF \sreg_reg[1337]  ( .D(o[1338]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1337]) );
  DFF \sreg_reg[1338]  ( .D(o[1339]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1338]) );
  DFF \sreg_reg[1339]  ( .D(o[1340]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1339]) );
  DFF \sreg_reg[1340]  ( .D(o[1341]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1340]) );
  DFF \sreg_reg[1341]  ( .D(o[1342]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1341]) );
  DFF \sreg_reg[1342]  ( .D(o[1343]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1342]) );
  DFF \sreg_reg[1343]  ( .D(o[1344]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1343]) );
  DFF \sreg_reg[1344]  ( .D(o[1345]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1344]) );
  DFF \sreg_reg[1345]  ( .D(o[1346]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1345]) );
  DFF \sreg_reg[1346]  ( .D(o[1347]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1346]) );
  DFF \sreg_reg[1347]  ( .D(o[1348]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1347]) );
  DFF \sreg_reg[1348]  ( .D(o[1349]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1348]) );
  DFF \sreg_reg[1349]  ( .D(o[1350]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1349]) );
  DFF \sreg_reg[1350]  ( .D(o[1351]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1350]) );
  DFF \sreg_reg[1351]  ( .D(o[1352]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1351]) );
  DFF \sreg_reg[1352]  ( .D(o[1353]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1352]) );
  DFF \sreg_reg[1353]  ( .D(o[1354]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1353]) );
  DFF \sreg_reg[1354]  ( .D(o[1355]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1354]) );
  DFF \sreg_reg[1355]  ( .D(o[1356]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1355]) );
  DFF \sreg_reg[1356]  ( .D(o[1357]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1356]) );
  DFF \sreg_reg[1357]  ( .D(o[1358]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1357]) );
  DFF \sreg_reg[1358]  ( .D(o[1359]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1358]) );
  DFF \sreg_reg[1359]  ( .D(o[1360]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1359]) );
  DFF \sreg_reg[1360]  ( .D(o[1361]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1360]) );
  DFF \sreg_reg[1361]  ( .D(o[1362]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1361]) );
  DFF \sreg_reg[1362]  ( .D(o[1363]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1362]) );
  DFF \sreg_reg[1363]  ( .D(o[1364]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1363]) );
  DFF \sreg_reg[1364]  ( .D(o[1365]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1364]) );
  DFF \sreg_reg[1365]  ( .D(o[1366]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1365]) );
  DFF \sreg_reg[1366]  ( .D(o[1367]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1366]) );
  DFF \sreg_reg[1367]  ( .D(o[1368]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1367]) );
  DFF \sreg_reg[1368]  ( .D(o[1369]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1368]) );
  DFF \sreg_reg[1369]  ( .D(o[1370]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1369]) );
  DFF \sreg_reg[1370]  ( .D(o[1371]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1370]) );
  DFF \sreg_reg[1371]  ( .D(o[1372]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1371]) );
  DFF \sreg_reg[1372]  ( .D(o[1373]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1372]) );
  DFF \sreg_reg[1373]  ( .D(o[1374]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1373]) );
  DFF \sreg_reg[1374]  ( .D(o[1375]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1374]) );
  DFF \sreg_reg[1375]  ( .D(o[1376]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1375]) );
  DFF \sreg_reg[1376]  ( .D(o[1377]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1376]) );
  DFF \sreg_reg[1377]  ( .D(o[1378]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1377]) );
  DFF \sreg_reg[1378]  ( .D(o[1379]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1378]) );
  DFF \sreg_reg[1379]  ( .D(o[1380]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1379]) );
  DFF \sreg_reg[1380]  ( .D(o[1381]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1380]) );
  DFF \sreg_reg[1381]  ( .D(o[1382]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1381]) );
  DFF \sreg_reg[1382]  ( .D(o[1383]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1382]) );
  DFF \sreg_reg[1383]  ( .D(o[1384]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1383]) );
  DFF \sreg_reg[1384]  ( .D(o[1385]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1384]) );
  DFF \sreg_reg[1385]  ( .D(o[1386]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1385]) );
  DFF \sreg_reg[1386]  ( .D(o[1387]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1386]) );
  DFF \sreg_reg[1387]  ( .D(o[1388]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1387]) );
  DFF \sreg_reg[1388]  ( .D(o[1389]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1388]) );
  DFF \sreg_reg[1389]  ( .D(o[1390]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1389]) );
  DFF \sreg_reg[1390]  ( .D(o[1391]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1390]) );
  DFF \sreg_reg[1391]  ( .D(o[1392]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1391]) );
  DFF \sreg_reg[1392]  ( .D(o[1393]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1392]) );
  DFF \sreg_reg[1393]  ( .D(o[1394]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1393]) );
  DFF \sreg_reg[1394]  ( .D(o[1395]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1394]) );
  DFF \sreg_reg[1395]  ( .D(o[1396]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1395]) );
  DFF \sreg_reg[1396]  ( .D(o[1397]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1396]) );
  DFF \sreg_reg[1397]  ( .D(o[1398]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1397]) );
  DFF \sreg_reg[1398]  ( .D(o[1399]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1398]) );
  DFF \sreg_reg[1399]  ( .D(o[1400]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1399]) );
  DFF \sreg_reg[1400]  ( .D(o[1401]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1400]) );
  DFF \sreg_reg[1401]  ( .D(o[1402]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1401]) );
  DFF \sreg_reg[1402]  ( .D(o[1403]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1402]) );
  DFF \sreg_reg[1403]  ( .D(o[1404]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1403]) );
  DFF \sreg_reg[1404]  ( .D(o[1405]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1404]) );
  DFF \sreg_reg[1405]  ( .D(o[1406]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1405]) );
  DFF \sreg_reg[1406]  ( .D(o[1407]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1406]) );
  DFF \sreg_reg[1407]  ( .D(o[1408]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1407]) );
  DFF \sreg_reg[1408]  ( .D(o[1409]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1408]) );
  DFF \sreg_reg[1409]  ( .D(o[1410]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1409]) );
  DFF \sreg_reg[1410]  ( .D(o[1411]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1410]) );
  DFF \sreg_reg[1411]  ( .D(o[1412]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1411]) );
  DFF \sreg_reg[1412]  ( .D(o[1413]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1412]) );
  DFF \sreg_reg[1413]  ( .D(o[1414]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1413]) );
  DFF \sreg_reg[1414]  ( .D(o[1415]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1414]) );
  DFF \sreg_reg[1415]  ( .D(o[1416]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1415]) );
  DFF \sreg_reg[1416]  ( .D(o[1417]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1416]) );
  DFF \sreg_reg[1417]  ( .D(o[1418]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1417]) );
  DFF \sreg_reg[1418]  ( .D(o[1419]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1418]) );
  DFF \sreg_reg[1419]  ( .D(o[1420]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1419]) );
  DFF \sreg_reg[1420]  ( .D(o[1421]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1420]) );
  DFF \sreg_reg[1421]  ( .D(o[1422]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1421]) );
  DFF \sreg_reg[1422]  ( .D(o[1423]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1422]) );
  DFF \sreg_reg[1423]  ( .D(o[1424]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1423]) );
  DFF \sreg_reg[1424]  ( .D(o[1425]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1424]) );
  DFF \sreg_reg[1425]  ( .D(o[1426]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1425]) );
  DFF \sreg_reg[1426]  ( .D(o[1427]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1426]) );
  DFF \sreg_reg[1427]  ( .D(o[1428]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1427]) );
  DFF \sreg_reg[1428]  ( .D(o[1429]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1428]) );
  DFF \sreg_reg[1429]  ( .D(o[1430]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1429]) );
  DFF \sreg_reg[1430]  ( .D(o[1431]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1430]) );
  DFF \sreg_reg[1431]  ( .D(o[1432]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1431]) );
  DFF \sreg_reg[1432]  ( .D(o[1433]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1432]) );
  DFF \sreg_reg[1433]  ( .D(o[1434]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1433]) );
  DFF \sreg_reg[1434]  ( .D(o[1435]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1434]) );
  DFF \sreg_reg[1435]  ( .D(o[1436]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1435]) );
  DFF \sreg_reg[1436]  ( .D(o[1437]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1436]) );
  DFF \sreg_reg[1437]  ( .D(o[1438]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1437]) );
  DFF \sreg_reg[1438]  ( .D(o[1439]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1438]) );
  DFF \sreg_reg[1439]  ( .D(o[1440]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1439]) );
  DFF \sreg_reg[1440]  ( .D(o[1441]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1440]) );
  DFF \sreg_reg[1441]  ( .D(o[1442]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1441]) );
  DFF \sreg_reg[1442]  ( .D(o[1443]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1442]) );
  DFF \sreg_reg[1443]  ( .D(o[1444]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1443]) );
  DFF \sreg_reg[1444]  ( .D(o[1445]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1444]) );
  DFF \sreg_reg[1445]  ( .D(o[1446]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1445]) );
  DFF \sreg_reg[1446]  ( .D(o[1447]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1446]) );
  DFF \sreg_reg[1447]  ( .D(o[1448]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1447]) );
  DFF \sreg_reg[1448]  ( .D(o[1449]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1448]) );
  DFF \sreg_reg[1449]  ( .D(o[1450]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1449]) );
  DFF \sreg_reg[1450]  ( .D(o[1451]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1450]) );
  DFF \sreg_reg[1451]  ( .D(o[1452]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1451]) );
  DFF \sreg_reg[1452]  ( .D(o[1453]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1452]) );
  DFF \sreg_reg[1453]  ( .D(o[1454]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1453]) );
  DFF \sreg_reg[1454]  ( .D(o[1455]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1454]) );
  DFF \sreg_reg[1455]  ( .D(o[1456]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1455]) );
  DFF \sreg_reg[1456]  ( .D(o[1457]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1456]) );
  DFF \sreg_reg[1457]  ( .D(o[1458]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1457]) );
  DFF \sreg_reg[1458]  ( .D(o[1459]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1458]) );
  DFF \sreg_reg[1459]  ( .D(o[1460]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1459]) );
  DFF \sreg_reg[1460]  ( .D(o[1461]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1460]) );
  DFF \sreg_reg[1461]  ( .D(o[1462]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1461]) );
  DFF \sreg_reg[1462]  ( .D(o[1463]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1462]) );
  DFF \sreg_reg[1463]  ( .D(o[1464]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1463]) );
  DFF \sreg_reg[1464]  ( .D(o[1465]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1464]) );
  DFF \sreg_reg[1465]  ( .D(o[1466]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1465]) );
  DFF \sreg_reg[1466]  ( .D(o[1467]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1466]) );
  DFF \sreg_reg[1467]  ( .D(o[1468]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1467]) );
  DFF \sreg_reg[1468]  ( .D(o[1469]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1468]) );
  DFF \sreg_reg[1469]  ( .D(o[1470]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1469]) );
  DFF \sreg_reg[1470]  ( .D(o[1471]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1470]) );
  DFF \sreg_reg[1471]  ( .D(o[1472]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1471]) );
  DFF \sreg_reg[1472]  ( .D(o[1473]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1472]) );
  DFF \sreg_reg[1473]  ( .D(o[1474]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1473]) );
  DFF \sreg_reg[1474]  ( .D(o[1475]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1474]) );
  DFF \sreg_reg[1475]  ( .D(o[1476]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1475]) );
  DFF \sreg_reg[1476]  ( .D(o[1477]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1476]) );
  DFF \sreg_reg[1477]  ( .D(o[1478]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1477]) );
  DFF \sreg_reg[1478]  ( .D(o[1479]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1478]) );
  DFF \sreg_reg[1479]  ( .D(o[1480]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1479]) );
  DFF \sreg_reg[1480]  ( .D(o[1481]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1480]) );
  DFF \sreg_reg[1481]  ( .D(o[1482]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1481]) );
  DFF \sreg_reg[1482]  ( .D(o[1483]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1482]) );
  DFF \sreg_reg[1483]  ( .D(o[1484]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1483]) );
  DFF \sreg_reg[1484]  ( .D(o[1485]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1484]) );
  DFF \sreg_reg[1485]  ( .D(o[1486]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1485]) );
  DFF \sreg_reg[1486]  ( .D(o[1487]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1486]) );
  DFF \sreg_reg[1487]  ( .D(o[1488]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1487]) );
  DFF \sreg_reg[1488]  ( .D(o[1489]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1488]) );
  DFF \sreg_reg[1489]  ( .D(o[1490]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1489]) );
  DFF \sreg_reg[1490]  ( .D(o[1491]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1490]) );
  DFF \sreg_reg[1491]  ( .D(o[1492]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1491]) );
  DFF \sreg_reg[1492]  ( .D(o[1493]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1492]) );
  DFF \sreg_reg[1493]  ( .D(o[1494]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1493]) );
  DFF \sreg_reg[1494]  ( .D(o[1495]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1494]) );
  DFF \sreg_reg[1495]  ( .D(o[1496]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1495]) );
  DFF \sreg_reg[1496]  ( .D(o[1497]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1496]) );
  DFF \sreg_reg[1497]  ( .D(o[1498]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1497]) );
  DFF \sreg_reg[1498]  ( .D(o[1499]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1498]) );
  DFF \sreg_reg[1499]  ( .D(o[1500]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1499]) );
  DFF \sreg_reg[1500]  ( .D(o[1501]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1500]) );
  DFF \sreg_reg[1501]  ( .D(o[1502]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1501]) );
  DFF \sreg_reg[1502]  ( .D(o[1503]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1502]) );
  DFF \sreg_reg[1503]  ( .D(o[1504]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1503]) );
  DFF \sreg_reg[1504]  ( .D(o[1505]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1504]) );
  DFF \sreg_reg[1505]  ( .D(o[1506]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1505]) );
  DFF \sreg_reg[1506]  ( .D(o[1507]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1506]) );
  DFF \sreg_reg[1507]  ( .D(o[1508]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1507]) );
  DFF \sreg_reg[1508]  ( .D(o[1509]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1508]) );
  DFF \sreg_reg[1509]  ( .D(o[1510]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1509]) );
  DFF \sreg_reg[1510]  ( .D(o[1511]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1510]) );
  DFF \sreg_reg[1511]  ( .D(o[1512]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1511]) );
  DFF \sreg_reg[1512]  ( .D(o[1513]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1512]) );
  DFF \sreg_reg[1513]  ( .D(o[1514]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1513]) );
  DFF \sreg_reg[1514]  ( .D(o[1515]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1514]) );
  DFF \sreg_reg[1515]  ( .D(o[1516]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1515]) );
  DFF \sreg_reg[1516]  ( .D(o[1517]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1516]) );
  DFF \sreg_reg[1517]  ( .D(o[1518]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1517]) );
  DFF \sreg_reg[1518]  ( .D(o[1519]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1518]) );
  DFF \sreg_reg[1519]  ( .D(o[1520]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1519]) );
  DFF \sreg_reg[1520]  ( .D(o[1521]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1520]) );
  DFF \sreg_reg[1521]  ( .D(o[1522]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1521]) );
  DFF \sreg_reg[1522]  ( .D(o[1523]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1522]) );
  DFF \sreg_reg[1523]  ( .D(o[1524]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1523]) );
  DFF \sreg_reg[1524]  ( .D(o[1525]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1524]) );
  DFF \sreg_reg[1525]  ( .D(o[1526]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1525]) );
  DFF \sreg_reg[1526]  ( .D(o[1527]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1526]) );
  DFF \sreg_reg[1527]  ( .D(o[1528]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1527]) );
  DFF \sreg_reg[1528]  ( .D(o[1529]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1528]) );
  DFF \sreg_reg[1529]  ( .D(o[1530]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1529]) );
  DFF \sreg_reg[1530]  ( .D(o[1531]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1530]) );
  DFF \sreg_reg[1531]  ( .D(o[1532]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1531]) );
  DFF \sreg_reg[1532]  ( .D(o[1533]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1532]) );
  DFF \sreg_reg[1533]  ( .D(o[1534]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1533]) );
  DFF \sreg_reg[1534]  ( .D(o[1535]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1534]) );
  DFF \sreg_reg[1535]  ( .D(o[1536]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1535]) );
  DFF \sreg_reg[1536]  ( .D(o[1537]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1536]) );
  DFF \sreg_reg[1537]  ( .D(o[1538]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1537]) );
  DFF \sreg_reg[1538]  ( .D(o[1539]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1538]) );
  DFF \sreg_reg[1539]  ( .D(o[1540]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1539]) );
  DFF \sreg_reg[1540]  ( .D(o[1541]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1540]) );
  DFF \sreg_reg[1541]  ( .D(o[1542]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1541]) );
  DFF \sreg_reg[1542]  ( .D(o[1543]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1542]) );
  DFF \sreg_reg[1543]  ( .D(o[1544]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1543]) );
  DFF \sreg_reg[1544]  ( .D(o[1545]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1544]) );
  DFF \sreg_reg[1545]  ( .D(o[1546]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1545]) );
  DFF \sreg_reg[1546]  ( .D(o[1547]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1546]) );
  DFF \sreg_reg[1547]  ( .D(o[1548]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1547]) );
  DFF \sreg_reg[1548]  ( .D(o[1549]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1548]) );
  DFF \sreg_reg[1549]  ( .D(o[1550]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1549]) );
  DFF \sreg_reg[1550]  ( .D(o[1551]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1550]) );
  DFF \sreg_reg[1551]  ( .D(o[1552]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1551]) );
  DFF \sreg_reg[1552]  ( .D(o[1553]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1552]) );
  DFF \sreg_reg[1553]  ( .D(o[1554]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1553]) );
  DFF \sreg_reg[1554]  ( .D(o[1555]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1554]) );
  DFF \sreg_reg[1555]  ( .D(o[1556]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1555]) );
  DFF \sreg_reg[1556]  ( .D(o[1557]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1556]) );
  DFF \sreg_reg[1557]  ( .D(o[1558]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1557]) );
  DFF \sreg_reg[1558]  ( .D(o[1559]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1558]) );
  DFF \sreg_reg[1559]  ( .D(o[1560]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1559]) );
  DFF \sreg_reg[1560]  ( .D(o[1561]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1560]) );
  DFF \sreg_reg[1561]  ( .D(o[1562]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1561]) );
  DFF \sreg_reg[1562]  ( .D(o[1563]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1562]) );
  DFF \sreg_reg[1563]  ( .D(o[1564]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1563]) );
  DFF \sreg_reg[1564]  ( .D(o[1565]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1564]) );
  DFF \sreg_reg[1565]  ( .D(o[1566]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1565]) );
  DFF \sreg_reg[1566]  ( .D(o[1567]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1566]) );
  DFF \sreg_reg[1567]  ( .D(o[1568]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1567]) );
  DFF \sreg_reg[1568]  ( .D(o[1569]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1568]) );
  DFF \sreg_reg[1569]  ( .D(o[1570]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1569]) );
  DFF \sreg_reg[1570]  ( .D(o[1571]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1570]) );
  DFF \sreg_reg[1571]  ( .D(o[1572]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1571]) );
  DFF \sreg_reg[1572]  ( .D(o[1573]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1572]) );
  DFF \sreg_reg[1573]  ( .D(o[1574]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1573]) );
  DFF \sreg_reg[1574]  ( .D(o[1575]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1574]) );
  DFF \sreg_reg[1575]  ( .D(o[1576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1575]) );
  DFF \sreg_reg[1576]  ( .D(o[1577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1576]) );
  DFF \sreg_reg[1577]  ( .D(o[1578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1577]) );
  DFF \sreg_reg[1578]  ( .D(o[1579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1578]) );
  DFF \sreg_reg[1579]  ( .D(o[1580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1579]) );
  DFF \sreg_reg[1580]  ( .D(o[1581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1580]) );
  DFF \sreg_reg[1581]  ( .D(o[1582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1581]) );
  DFF \sreg_reg[1582]  ( .D(o[1583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1582]) );
  DFF \sreg_reg[1583]  ( .D(o[1584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1583]) );
  DFF \sreg_reg[1584]  ( .D(o[1585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1584]) );
  DFF \sreg_reg[1585]  ( .D(o[1586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1585]) );
  DFF \sreg_reg[1586]  ( .D(o[1587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1586]) );
  DFF \sreg_reg[1587]  ( .D(o[1588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1587]) );
  DFF \sreg_reg[1588]  ( .D(o[1589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1588]) );
  DFF \sreg_reg[1589]  ( .D(o[1590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1589]) );
  DFF \sreg_reg[1590]  ( .D(o[1591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1590]) );
  DFF \sreg_reg[1591]  ( .D(o[1592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1591]) );
  DFF \sreg_reg[1592]  ( .D(o[1593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1592]) );
  DFF \sreg_reg[1593]  ( .D(o[1594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1593]) );
  DFF \sreg_reg[1594]  ( .D(o[1595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1594]) );
  DFF \sreg_reg[1595]  ( .D(o[1596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1595]) );
  DFF \sreg_reg[1596]  ( .D(o[1597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1596]) );
  DFF \sreg_reg[1597]  ( .D(o[1598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1597]) );
  DFF \sreg_reg[1598]  ( .D(o[1599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1598]) );
  DFF \sreg_reg[1599]  ( .D(o[1600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1599]) );
  DFF \sreg_reg[1600]  ( .D(o[1601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1600]) );
  DFF \sreg_reg[1601]  ( .D(o[1602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1601]) );
  DFF \sreg_reg[1602]  ( .D(o[1603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1602]) );
  DFF \sreg_reg[1603]  ( .D(o[1604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1603]) );
  DFF \sreg_reg[1604]  ( .D(o[1605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1604]) );
  DFF \sreg_reg[1605]  ( .D(o[1606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1605]) );
  DFF \sreg_reg[1606]  ( .D(o[1607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1606]) );
  DFF \sreg_reg[1607]  ( .D(o[1608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1607]) );
  DFF \sreg_reg[1608]  ( .D(o[1609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1608]) );
  DFF \sreg_reg[1609]  ( .D(o[1610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1609]) );
  DFF \sreg_reg[1610]  ( .D(o[1611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1610]) );
  DFF \sreg_reg[1611]  ( .D(o[1612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1611]) );
  DFF \sreg_reg[1612]  ( .D(o[1613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1612]) );
  DFF \sreg_reg[1613]  ( .D(o[1614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1613]) );
  DFF \sreg_reg[1614]  ( .D(o[1615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1614]) );
  DFF \sreg_reg[1615]  ( .D(o[1616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1615]) );
  DFF \sreg_reg[1616]  ( .D(o[1617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1616]) );
  DFF \sreg_reg[1617]  ( .D(o[1618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1617]) );
  DFF \sreg_reg[1618]  ( .D(o[1619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1618]) );
  DFF \sreg_reg[1619]  ( .D(o[1620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1619]) );
  DFF \sreg_reg[1620]  ( .D(o[1621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1620]) );
  DFF \sreg_reg[1621]  ( .D(o[1622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1621]) );
  DFF \sreg_reg[1622]  ( .D(o[1623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1622]) );
  DFF \sreg_reg[1623]  ( .D(o[1624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1623]) );
  DFF \sreg_reg[1624]  ( .D(o[1625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1624]) );
  DFF \sreg_reg[1625]  ( .D(o[1626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1625]) );
  DFF \sreg_reg[1626]  ( .D(o[1627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1626]) );
  DFF \sreg_reg[1627]  ( .D(o[1628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1627]) );
  DFF \sreg_reg[1628]  ( .D(o[1629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1628]) );
  DFF \sreg_reg[1629]  ( .D(o[1630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1629]) );
  DFF \sreg_reg[1630]  ( .D(o[1631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1630]) );
  DFF \sreg_reg[1631]  ( .D(o[1632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1631]) );
  DFF \sreg_reg[1632]  ( .D(o[1633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1632]) );
  DFF \sreg_reg[1633]  ( .D(o[1634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1633]) );
  DFF \sreg_reg[1634]  ( .D(o[1635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1634]) );
  DFF \sreg_reg[1635]  ( .D(o[1636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1635]) );
  DFF \sreg_reg[1636]  ( .D(o[1637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1636]) );
  DFF \sreg_reg[1637]  ( .D(o[1638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1637]) );
  DFF \sreg_reg[1638]  ( .D(o[1639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1638]) );
  DFF \sreg_reg[1639]  ( .D(o[1640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1639]) );
  DFF \sreg_reg[1640]  ( .D(o[1641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1640]) );
  DFF \sreg_reg[1641]  ( .D(o[1642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1641]) );
  DFF \sreg_reg[1642]  ( .D(o[1643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1642]) );
  DFF \sreg_reg[1643]  ( .D(o[1644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1643]) );
  DFF \sreg_reg[1644]  ( .D(o[1645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1644]) );
  DFF \sreg_reg[1645]  ( .D(o[1646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1645]) );
  DFF \sreg_reg[1646]  ( .D(o[1647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1646]) );
  DFF \sreg_reg[1647]  ( .D(o[1648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1647]) );
  DFF \sreg_reg[1648]  ( .D(o[1649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1648]) );
  DFF \sreg_reg[1649]  ( .D(o[1650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1649]) );
  DFF \sreg_reg[1650]  ( .D(o[1651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1650]) );
  DFF \sreg_reg[1651]  ( .D(o[1652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1651]) );
  DFF \sreg_reg[1652]  ( .D(o[1653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1652]) );
  DFF \sreg_reg[1653]  ( .D(o[1654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1653]) );
  DFF \sreg_reg[1654]  ( .D(o[1655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1654]) );
  DFF \sreg_reg[1655]  ( .D(o[1656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1655]) );
  DFF \sreg_reg[1656]  ( .D(o[1657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1656]) );
  DFF \sreg_reg[1657]  ( .D(o[1658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1657]) );
  DFF \sreg_reg[1658]  ( .D(o[1659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1658]) );
  DFF \sreg_reg[1659]  ( .D(o[1660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1659]) );
  DFF \sreg_reg[1660]  ( .D(o[1661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1660]) );
  DFF \sreg_reg[1661]  ( .D(o[1662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1661]) );
  DFF \sreg_reg[1662]  ( .D(o[1663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1662]) );
  DFF \sreg_reg[1663]  ( .D(o[1664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1663]) );
  DFF \sreg_reg[1664]  ( .D(o[1665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1664]) );
  DFF \sreg_reg[1665]  ( .D(o[1666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1665]) );
  DFF \sreg_reg[1666]  ( .D(o[1667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1666]) );
  DFF \sreg_reg[1667]  ( .D(o[1668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1667]) );
  DFF \sreg_reg[1668]  ( .D(o[1669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1668]) );
  DFF \sreg_reg[1669]  ( .D(o[1670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1669]) );
  DFF \sreg_reg[1670]  ( .D(o[1671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1670]) );
  DFF \sreg_reg[1671]  ( .D(o[1672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1671]) );
  DFF \sreg_reg[1672]  ( .D(o[1673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1672]) );
  DFF \sreg_reg[1673]  ( .D(o[1674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1673]) );
  DFF \sreg_reg[1674]  ( .D(o[1675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1674]) );
  DFF \sreg_reg[1675]  ( .D(o[1676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1675]) );
  DFF \sreg_reg[1676]  ( .D(o[1677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1676]) );
  DFF \sreg_reg[1677]  ( .D(o[1678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1677]) );
  DFF \sreg_reg[1678]  ( .D(o[1679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1678]) );
  DFF \sreg_reg[1679]  ( .D(o[1680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1679]) );
  DFF \sreg_reg[1680]  ( .D(o[1681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1680]) );
  DFF \sreg_reg[1681]  ( .D(o[1682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1681]) );
  DFF \sreg_reg[1682]  ( .D(o[1683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1682]) );
  DFF \sreg_reg[1683]  ( .D(o[1684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1683]) );
  DFF \sreg_reg[1684]  ( .D(o[1685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1684]) );
  DFF \sreg_reg[1685]  ( .D(o[1686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1685]) );
  DFF \sreg_reg[1686]  ( .D(o[1687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1686]) );
  DFF \sreg_reg[1687]  ( .D(o[1688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1687]) );
  DFF \sreg_reg[1688]  ( .D(o[1689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1688]) );
  DFF \sreg_reg[1689]  ( .D(o[1690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1689]) );
  DFF \sreg_reg[1690]  ( .D(o[1691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1690]) );
  DFF \sreg_reg[1691]  ( .D(o[1692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1691]) );
  DFF \sreg_reg[1692]  ( .D(o[1693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1692]) );
  DFF \sreg_reg[1693]  ( .D(o[1694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1693]) );
  DFF \sreg_reg[1694]  ( .D(o[1695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1694]) );
  DFF \sreg_reg[1695]  ( .D(o[1696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1695]) );
  DFF \sreg_reg[1696]  ( .D(o[1697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1696]) );
  DFF \sreg_reg[1697]  ( .D(o[1698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1697]) );
  DFF \sreg_reg[1698]  ( .D(o[1699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1698]) );
  DFF \sreg_reg[1699]  ( .D(o[1700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1699]) );
  DFF \sreg_reg[1700]  ( .D(o[1701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1700]) );
  DFF \sreg_reg[1701]  ( .D(o[1702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1701]) );
  DFF \sreg_reg[1702]  ( .D(o[1703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1702]) );
  DFF \sreg_reg[1703]  ( .D(o[1704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1703]) );
  DFF \sreg_reg[1704]  ( .D(o[1705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1704]) );
  DFF \sreg_reg[1705]  ( .D(o[1706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1705]) );
  DFF \sreg_reg[1706]  ( .D(o[1707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1706]) );
  DFF \sreg_reg[1707]  ( .D(o[1708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1707]) );
  DFF \sreg_reg[1708]  ( .D(o[1709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1708]) );
  DFF \sreg_reg[1709]  ( .D(o[1710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1709]) );
  DFF \sreg_reg[1710]  ( .D(o[1711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1710]) );
  DFF \sreg_reg[1711]  ( .D(o[1712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1711]) );
  DFF \sreg_reg[1712]  ( .D(o[1713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1712]) );
  DFF \sreg_reg[1713]  ( .D(o[1714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1713]) );
  DFF \sreg_reg[1714]  ( .D(o[1715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1714]) );
  DFF \sreg_reg[1715]  ( .D(o[1716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1715]) );
  DFF \sreg_reg[1716]  ( .D(o[1717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1716]) );
  DFF \sreg_reg[1717]  ( .D(o[1718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1717]) );
  DFF \sreg_reg[1718]  ( .D(o[1719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1718]) );
  DFF \sreg_reg[1719]  ( .D(o[1720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1719]) );
  DFF \sreg_reg[1720]  ( .D(o[1721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1720]) );
  DFF \sreg_reg[1721]  ( .D(o[1722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1721]) );
  DFF \sreg_reg[1722]  ( .D(o[1723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1722]) );
  DFF \sreg_reg[1723]  ( .D(o[1724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1723]) );
  DFF \sreg_reg[1724]  ( .D(o[1725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1724]) );
  DFF \sreg_reg[1725]  ( .D(o[1726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1725]) );
  DFF \sreg_reg[1726]  ( .D(o[1727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1726]) );
  DFF \sreg_reg[1727]  ( .D(o[1728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1727]) );
  DFF \sreg_reg[1728]  ( .D(o[1729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1728]) );
  DFF \sreg_reg[1729]  ( .D(o[1730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1729]) );
  DFF \sreg_reg[1730]  ( .D(o[1731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1730]) );
  DFF \sreg_reg[1731]  ( .D(o[1732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1731]) );
  DFF \sreg_reg[1732]  ( .D(o[1733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1732]) );
  DFF \sreg_reg[1733]  ( .D(o[1734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1733]) );
  DFF \sreg_reg[1734]  ( .D(o[1735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1734]) );
  DFF \sreg_reg[1735]  ( .D(o[1736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1735]) );
  DFF \sreg_reg[1736]  ( .D(o[1737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1736]) );
  DFF \sreg_reg[1737]  ( .D(o[1738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1737]) );
  DFF \sreg_reg[1738]  ( .D(o[1739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1738]) );
  DFF \sreg_reg[1739]  ( .D(o[1740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1739]) );
  DFF \sreg_reg[1740]  ( .D(o[1741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1740]) );
  DFF \sreg_reg[1741]  ( .D(o[1742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1741]) );
  DFF \sreg_reg[1742]  ( .D(o[1743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1742]) );
  DFF \sreg_reg[1743]  ( .D(o[1744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1743]) );
  DFF \sreg_reg[1744]  ( .D(o[1745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1744]) );
  DFF \sreg_reg[1745]  ( .D(o[1746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1745]) );
  DFF \sreg_reg[1746]  ( .D(o[1747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1746]) );
  DFF \sreg_reg[1747]  ( .D(o[1748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1747]) );
  DFF \sreg_reg[1748]  ( .D(o[1749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1748]) );
  DFF \sreg_reg[1749]  ( .D(o[1750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1749]) );
  DFF \sreg_reg[1750]  ( .D(o[1751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1750]) );
  DFF \sreg_reg[1751]  ( .D(o[1752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1751]) );
  DFF \sreg_reg[1752]  ( .D(o[1753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1752]) );
  DFF \sreg_reg[1753]  ( .D(o[1754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1753]) );
  DFF \sreg_reg[1754]  ( .D(o[1755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1754]) );
  DFF \sreg_reg[1755]  ( .D(o[1756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1755]) );
  DFF \sreg_reg[1756]  ( .D(o[1757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1756]) );
  DFF \sreg_reg[1757]  ( .D(o[1758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1757]) );
  DFF \sreg_reg[1758]  ( .D(o[1759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1758]) );
  DFF \sreg_reg[1759]  ( .D(o[1760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1759]) );
  DFF \sreg_reg[1760]  ( .D(o[1761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1760]) );
  DFF \sreg_reg[1761]  ( .D(o[1762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1761]) );
  DFF \sreg_reg[1762]  ( .D(o[1763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1762]) );
  DFF \sreg_reg[1763]  ( .D(o[1764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1763]) );
  DFF \sreg_reg[1764]  ( .D(o[1765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1764]) );
  DFF \sreg_reg[1765]  ( .D(o[1766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1765]) );
  DFF \sreg_reg[1766]  ( .D(o[1767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1766]) );
  DFF \sreg_reg[1767]  ( .D(o[1768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1767]) );
  DFF \sreg_reg[1768]  ( .D(o[1769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1768]) );
  DFF \sreg_reg[1769]  ( .D(o[1770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1769]) );
  DFF \sreg_reg[1770]  ( .D(o[1771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1770]) );
  DFF \sreg_reg[1771]  ( .D(o[1772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1771]) );
  DFF \sreg_reg[1772]  ( .D(o[1773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1772]) );
  DFF \sreg_reg[1773]  ( .D(o[1774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1773]) );
  DFF \sreg_reg[1774]  ( .D(o[1775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1774]) );
  DFF \sreg_reg[1775]  ( .D(o[1776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1775]) );
  DFF \sreg_reg[1776]  ( .D(o[1777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1776]) );
  DFF \sreg_reg[1777]  ( .D(o[1778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1777]) );
  DFF \sreg_reg[1778]  ( .D(o[1779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1778]) );
  DFF \sreg_reg[1779]  ( .D(o[1780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1779]) );
  DFF \sreg_reg[1780]  ( .D(o[1781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1780]) );
  DFF \sreg_reg[1781]  ( .D(o[1782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1781]) );
  DFF \sreg_reg[1782]  ( .D(o[1783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1782]) );
  DFF \sreg_reg[1783]  ( .D(o[1784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1783]) );
  DFF \sreg_reg[1784]  ( .D(o[1785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1784]) );
  DFF \sreg_reg[1785]  ( .D(o[1786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1785]) );
  DFF \sreg_reg[1786]  ( .D(o[1787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1786]) );
  DFF \sreg_reg[1787]  ( .D(o[1788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1787]) );
  DFF \sreg_reg[1788]  ( .D(o[1789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1788]) );
  DFF \sreg_reg[1789]  ( .D(o[1790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1789]) );
  DFF \sreg_reg[1790]  ( .D(o[1791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1790]) );
  DFF \sreg_reg[1791]  ( .D(o[1792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1791]) );
  DFF \sreg_reg[1792]  ( .D(o[1793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1792]) );
  DFF \sreg_reg[1793]  ( .D(o[1794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1793]) );
  DFF \sreg_reg[1794]  ( .D(o[1795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1794]) );
  DFF \sreg_reg[1795]  ( .D(o[1796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1795]) );
  DFF \sreg_reg[1796]  ( .D(o[1797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1796]) );
  DFF \sreg_reg[1797]  ( .D(o[1798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1797]) );
  DFF \sreg_reg[1798]  ( .D(o[1799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1798]) );
  DFF \sreg_reg[1799]  ( .D(o[1800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1799]) );
  DFF \sreg_reg[1800]  ( .D(o[1801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1800]) );
  DFF \sreg_reg[1801]  ( .D(o[1802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1801]) );
  DFF \sreg_reg[1802]  ( .D(o[1803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1802]) );
  DFF \sreg_reg[1803]  ( .D(o[1804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1803]) );
  DFF \sreg_reg[1804]  ( .D(o[1805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1804]) );
  DFF \sreg_reg[1805]  ( .D(o[1806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1805]) );
  DFF \sreg_reg[1806]  ( .D(o[1807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1806]) );
  DFF \sreg_reg[1807]  ( .D(o[1808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1807]) );
  DFF \sreg_reg[1808]  ( .D(o[1809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1808]) );
  DFF \sreg_reg[1809]  ( .D(o[1810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1809]) );
  DFF \sreg_reg[1810]  ( .D(o[1811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1810]) );
  DFF \sreg_reg[1811]  ( .D(o[1812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1811]) );
  DFF \sreg_reg[1812]  ( .D(o[1813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1812]) );
  DFF \sreg_reg[1813]  ( .D(o[1814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1813]) );
  DFF \sreg_reg[1814]  ( .D(o[1815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1814]) );
  DFF \sreg_reg[1815]  ( .D(o[1816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1815]) );
  DFF \sreg_reg[1816]  ( .D(o[1817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1816]) );
  DFF \sreg_reg[1817]  ( .D(o[1818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1817]) );
  DFF \sreg_reg[1818]  ( .D(o[1819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1818]) );
  DFF \sreg_reg[1819]  ( .D(o[1820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1819]) );
  DFF \sreg_reg[1820]  ( .D(o[1821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1820]) );
  DFF \sreg_reg[1821]  ( .D(o[1822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1821]) );
  DFF \sreg_reg[1822]  ( .D(o[1823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1822]) );
  DFF \sreg_reg[1823]  ( .D(o[1824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1823]) );
  DFF \sreg_reg[1824]  ( .D(o[1825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1824]) );
  DFF \sreg_reg[1825]  ( .D(o[1826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1825]) );
  DFF \sreg_reg[1826]  ( .D(o[1827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1826]) );
  DFF \sreg_reg[1827]  ( .D(o[1828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1827]) );
  DFF \sreg_reg[1828]  ( .D(o[1829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1828]) );
  DFF \sreg_reg[1829]  ( .D(o[1830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1829]) );
  DFF \sreg_reg[1830]  ( .D(o[1831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1830]) );
  DFF \sreg_reg[1831]  ( .D(o[1832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1831]) );
  DFF \sreg_reg[1832]  ( .D(o[1833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1832]) );
  DFF \sreg_reg[1833]  ( .D(o[1834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1833]) );
  DFF \sreg_reg[1834]  ( .D(o[1835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1834]) );
  DFF \sreg_reg[1835]  ( .D(o[1836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1835]) );
  DFF \sreg_reg[1836]  ( .D(o[1837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1836]) );
  DFF \sreg_reg[1837]  ( .D(o[1838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1837]) );
  DFF \sreg_reg[1838]  ( .D(o[1839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1838]) );
  DFF \sreg_reg[1839]  ( .D(o[1840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1839]) );
  DFF \sreg_reg[1840]  ( .D(o[1841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1840]) );
  DFF \sreg_reg[1841]  ( .D(o[1842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1841]) );
  DFF \sreg_reg[1842]  ( .D(o[1843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1842]) );
  DFF \sreg_reg[1843]  ( .D(o[1844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1843]) );
  DFF \sreg_reg[1844]  ( .D(o[1845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1844]) );
  DFF \sreg_reg[1845]  ( .D(o[1846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1845]) );
  DFF \sreg_reg[1846]  ( .D(o[1847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1846]) );
  DFF \sreg_reg[1847]  ( .D(o[1848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1847]) );
  DFF \sreg_reg[1848]  ( .D(o[1849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1848]) );
  DFF \sreg_reg[1849]  ( .D(o[1850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1849]) );
  DFF \sreg_reg[1850]  ( .D(o[1851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1850]) );
  DFF \sreg_reg[1851]  ( .D(o[1852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1851]) );
  DFF \sreg_reg[1852]  ( .D(o[1853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1852]) );
  DFF \sreg_reg[1853]  ( .D(o[1854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1853]) );
  DFF \sreg_reg[1854]  ( .D(o[1855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1854]) );
  DFF \sreg_reg[1855]  ( .D(o[1856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1855]) );
  DFF \sreg_reg[1856]  ( .D(o[1857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1856]) );
  DFF \sreg_reg[1857]  ( .D(o[1858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1857]) );
  DFF \sreg_reg[1858]  ( .D(o[1859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1858]) );
  DFF \sreg_reg[1859]  ( .D(o[1860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1859]) );
  DFF \sreg_reg[1860]  ( .D(o[1861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1860]) );
  DFF \sreg_reg[1861]  ( .D(o[1862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1861]) );
  DFF \sreg_reg[1862]  ( .D(o[1863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1862]) );
  DFF \sreg_reg[1863]  ( .D(o[1864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1863]) );
  DFF \sreg_reg[1864]  ( .D(o[1865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1864]) );
  DFF \sreg_reg[1865]  ( .D(o[1866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1865]) );
  DFF \sreg_reg[1866]  ( .D(o[1867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1866]) );
  DFF \sreg_reg[1867]  ( .D(o[1868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1867]) );
  DFF \sreg_reg[1868]  ( .D(o[1869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1868]) );
  DFF \sreg_reg[1869]  ( .D(o[1870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1869]) );
  DFF \sreg_reg[1870]  ( .D(o[1871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1870]) );
  DFF \sreg_reg[1871]  ( .D(o[1872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1871]) );
  DFF \sreg_reg[1872]  ( .D(o[1873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1872]) );
  DFF \sreg_reg[1873]  ( .D(o[1874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1873]) );
  DFF \sreg_reg[1874]  ( .D(o[1875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1874]) );
  DFF \sreg_reg[1875]  ( .D(o[1876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1875]) );
  DFF \sreg_reg[1876]  ( .D(o[1877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1876]) );
  DFF \sreg_reg[1877]  ( .D(o[1878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1877]) );
  DFF \sreg_reg[1878]  ( .D(o[1879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1878]) );
  DFF \sreg_reg[1879]  ( .D(o[1880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1879]) );
  DFF \sreg_reg[1880]  ( .D(o[1881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1880]) );
  DFF \sreg_reg[1881]  ( .D(o[1882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1881]) );
  DFF \sreg_reg[1882]  ( .D(o[1883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1882]) );
  DFF \sreg_reg[1883]  ( .D(o[1884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1883]) );
  DFF \sreg_reg[1884]  ( .D(o[1885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1884]) );
  DFF \sreg_reg[1885]  ( .D(o[1886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1885]) );
  DFF \sreg_reg[1886]  ( .D(o[1887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1886]) );
  DFF \sreg_reg[1887]  ( .D(o[1888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1887]) );
  DFF \sreg_reg[1888]  ( .D(o[1889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1888]) );
  DFF \sreg_reg[1889]  ( .D(o[1890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1889]) );
  DFF \sreg_reg[1890]  ( .D(o[1891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1890]) );
  DFF \sreg_reg[1891]  ( .D(o[1892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1891]) );
  DFF \sreg_reg[1892]  ( .D(o[1893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1892]) );
  DFF \sreg_reg[1893]  ( .D(o[1894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1893]) );
  DFF \sreg_reg[1894]  ( .D(o[1895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1894]) );
  DFF \sreg_reg[1895]  ( .D(o[1896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1895]) );
  DFF \sreg_reg[1896]  ( .D(o[1897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1896]) );
  DFF \sreg_reg[1897]  ( .D(o[1898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1897]) );
  DFF \sreg_reg[1898]  ( .D(o[1899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1898]) );
  DFF \sreg_reg[1899]  ( .D(o[1900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1899]) );
  DFF \sreg_reg[1900]  ( .D(o[1901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1900]) );
  DFF \sreg_reg[1901]  ( .D(o[1902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1901]) );
  DFF \sreg_reg[1902]  ( .D(o[1903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1902]) );
  DFF \sreg_reg[1903]  ( .D(o[1904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1903]) );
  DFF \sreg_reg[1904]  ( .D(o[1905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1904]) );
  DFF \sreg_reg[1905]  ( .D(o[1906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1905]) );
  DFF \sreg_reg[1906]  ( .D(o[1907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1906]) );
  DFF \sreg_reg[1907]  ( .D(o[1908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1907]) );
  DFF \sreg_reg[1908]  ( .D(o[1909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1908]) );
  DFF \sreg_reg[1909]  ( .D(o[1910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1909]) );
  DFF \sreg_reg[1910]  ( .D(o[1911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1910]) );
  DFF \sreg_reg[1911]  ( .D(o[1912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1911]) );
  DFF \sreg_reg[1912]  ( .D(o[1913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1912]) );
  DFF \sreg_reg[1913]  ( .D(o[1914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1913]) );
  DFF \sreg_reg[1914]  ( .D(o[1915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1914]) );
  DFF \sreg_reg[1915]  ( .D(o[1916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1915]) );
  DFF \sreg_reg[1916]  ( .D(o[1917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1916]) );
  DFF \sreg_reg[1917]  ( .D(o[1918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1917]) );
  DFF \sreg_reg[1918]  ( .D(o[1919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1918]) );
  DFF \sreg_reg[1919]  ( .D(o[1920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1919]) );
  DFF \sreg_reg[1920]  ( .D(o[1921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1920]) );
  DFF \sreg_reg[1921]  ( .D(o[1922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1921]) );
  DFF \sreg_reg[1922]  ( .D(o[1923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1922]) );
  DFF \sreg_reg[1923]  ( .D(o[1924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1923]) );
  DFF \sreg_reg[1924]  ( .D(o[1925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1924]) );
  DFF \sreg_reg[1925]  ( .D(o[1926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1925]) );
  DFF \sreg_reg[1926]  ( .D(o[1927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1926]) );
  DFF \sreg_reg[1927]  ( .D(o[1928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1927]) );
  DFF \sreg_reg[1928]  ( .D(o[1929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1928]) );
  DFF \sreg_reg[1929]  ( .D(o[1930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1929]) );
  DFF \sreg_reg[1930]  ( .D(o[1931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1930]) );
  DFF \sreg_reg[1931]  ( .D(o[1932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1931]) );
  DFF \sreg_reg[1932]  ( .D(o[1933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1932]) );
  DFF \sreg_reg[1933]  ( .D(o[1934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1933]) );
  DFF \sreg_reg[1934]  ( .D(o[1935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1934]) );
  DFF \sreg_reg[1935]  ( .D(o[1936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1935]) );
  DFF \sreg_reg[1936]  ( .D(o[1937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1936]) );
  DFF \sreg_reg[1937]  ( .D(o[1938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1937]) );
  DFF \sreg_reg[1938]  ( .D(o[1939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1938]) );
  DFF \sreg_reg[1939]  ( .D(o[1940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1939]) );
  DFF \sreg_reg[1940]  ( .D(o[1941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1940]) );
  DFF \sreg_reg[1941]  ( .D(o[1942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1941]) );
  DFF \sreg_reg[1942]  ( .D(o[1943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1942]) );
  DFF \sreg_reg[1943]  ( .D(o[1944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1943]) );
  DFF \sreg_reg[1944]  ( .D(o[1945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1944]) );
  DFF \sreg_reg[1945]  ( .D(o[1946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1945]) );
  DFF \sreg_reg[1946]  ( .D(o[1947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1946]) );
  DFF \sreg_reg[1947]  ( .D(o[1948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1947]) );
  DFF \sreg_reg[1948]  ( .D(o[1949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1948]) );
  DFF \sreg_reg[1949]  ( .D(o[1950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1949]) );
  DFF \sreg_reg[1950]  ( .D(o[1951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1950]) );
  DFF \sreg_reg[1951]  ( .D(o[1952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1951]) );
  DFF \sreg_reg[1952]  ( .D(o[1953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1952]) );
  DFF \sreg_reg[1953]  ( .D(o[1954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1953]) );
  DFF \sreg_reg[1954]  ( .D(o[1955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1954]) );
  DFF \sreg_reg[1955]  ( .D(o[1956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1955]) );
  DFF \sreg_reg[1956]  ( .D(o[1957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1956]) );
  DFF \sreg_reg[1957]  ( .D(o[1958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1957]) );
  DFF \sreg_reg[1958]  ( .D(o[1959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1958]) );
  DFF \sreg_reg[1959]  ( .D(o[1960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1959]) );
  DFF \sreg_reg[1960]  ( .D(o[1961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1960]) );
  DFF \sreg_reg[1961]  ( .D(o[1962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1961]) );
  DFF \sreg_reg[1962]  ( .D(o[1963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1962]) );
  DFF \sreg_reg[1963]  ( .D(o[1964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1963]) );
  DFF \sreg_reg[1964]  ( .D(o[1965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1964]) );
  DFF \sreg_reg[1965]  ( .D(o[1966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1965]) );
  DFF \sreg_reg[1966]  ( .D(o[1967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1966]) );
  DFF \sreg_reg[1967]  ( .D(o[1968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1967]) );
  DFF \sreg_reg[1968]  ( .D(o[1969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1968]) );
  DFF \sreg_reg[1969]  ( .D(o[1970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1969]) );
  DFF \sreg_reg[1970]  ( .D(o[1971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1970]) );
  DFF \sreg_reg[1971]  ( .D(o[1972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1971]) );
  DFF \sreg_reg[1972]  ( .D(o[1973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1972]) );
  DFF \sreg_reg[1973]  ( .D(o[1974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1973]) );
  DFF \sreg_reg[1974]  ( .D(o[1975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1974]) );
  DFF \sreg_reg[1975]  ( .D(o[1976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1975]) );
  DFF \sreg_reg[1976]  ( .D(o[1977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1976]) );
  DFF \sreg_reg[1977]  ( .D(o[1978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1977]) );
  DFF \sreg_reg[1978]  ( .D(o[1979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1978]) );
  DFF \sreg_reg[1979]  ( .D(o[1980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1979]) );
  DFF \sreg_reg[1980]  ( .D(o[1981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1980]) );
  DFF \sreg_reg[1981]  ( .D(o[1982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1981]) );
  DFF \sreg_reg[1982]  ( .D(o[1983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1982]) );
  DFF \sreg_reg[1983]  ( .D(o[1984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1983]) );
  DFF \sreg_reg[1984]  ( .D(o[1985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1984]) );
  DFF \sreg_reg[1985]  ( .D(o[1986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1985]) );
  DFF \sreg_reg[1986]  ( .D(o[1987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1986]) );
  DFF \sreg_reg[1987]  ( .D(o[1988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1987]) );
  DFF \sreg_reg[1988]  ( .D(o[1989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1988]) );
  DFF \sreg_reg[1989]  ( .D(o[1990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1989]) );
  DFF \sreg_reg[1990]  ( .D(o[1991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1990]) );
  DFF \sreg_reg[1991]  ( .D(o[1992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1991]) );
  DFF \sreg_reg[1992]  ( .D(o[1993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1992]) );
  DFF \sreg_reg[1993]  ( .D(o[1994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1993]) );
  DFF \sreg_reg[1994]  ( .D(o[1995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1994]) );
  DFF \sreg_reg[1995]  ( .D(o[1996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1995]) );
  DFF \sreg_reg[1996]  ( .D(o[1997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1996]) );
  DFF \sreg_reg[1997]  ( .D(o[1998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1997]) );
  DFF \sreg_reg[1998]  ( .D(o[1999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1998]) );
  DFF \sreg_reg[1999]  ( .D(o[2000]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1999]) );
  DFF \sreg_reg[2000]  ( .D(o[2001]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2000]) );
  DFF \sreg_reg[2001]  ( .D(o[2002]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2001]) );
  DFF \sreg_reg[2002]  ( .D(o[2003]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2002]) );
  DFF \sreg_reg[2003]  ( .D(o[2004]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2003]) );
  DFF \sreg_reg[2004]  ( .D(o[2005]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2004]) );
  DFF \sreg_reg[2005]  ( .D(o[2006]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2005]) );
  DFF \sreg_reg[2006]  ( .D(o[2007]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2006]) );
  DFF \sreg_reg[2007]  ( .D(o[2008]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2007]) );
  DFF \sreg_reg[2008]  ( .D(o[2009]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2008]) );
  DFF \sreg_reg[2009]  ( .D(o[2010]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2009]) );
  DFF \sreg_reg[2010]  ( .D(o[2011]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2010]) );
  DFF \sreg_reg[2011]  ( .D(o[2012]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2011]) );
  DFF \sreg_reg[2012]  ( .D(o[2013]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2012]) );
  DFF \sreg_reg[2013]  ( .D(o[2014]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2013]) );
  DFF \sreg_reg[2014]  ( .D(o[2015]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2014]) );
  DFF \sreg_reg[2015]  ( .D(o[2016]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2015]) );
  DFF \sreg_reg[2016]  ( .D(o[2017]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2016]) );
  DFF \sreg_reg[2017]  ( .D(o[2018]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2017]) );
  DFF \sreg_reg[2018]  ( .D(o[2019]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2018]) );
  DFF \sreg_reg[2019]  ( .D(o[2020]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2019]) );
  DFF \sreg_reg[2020]  ( .D(o[2021]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2020]) );
  DFF \sreg_reg[2021]  ( .D(o[2022]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2021]) );
  DFF \sreg_reg[2022]  ( .D(o[2023]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2022]) );
  DFF \sreg_reg[2023]  ( .D(o[2024]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2023]) );
  DFF \sreg_reg[2024]  ( .D(o[2025]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2024]) );
  DFF \sreg_reg[2025]  ( .D(o[2026]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2025]) );
  DFF \sreg_reg[2026]  ( .D(o[2027]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2026]) );
  DFF \sreg_reg[2027]  ( .D(o[2028]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2027]) );
  DFF \sreg_reg[2028]  ( .D(o[2029]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2028]) );
  DFF \sreg_reg[2029]  ( .D(o[2030]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2029]) );
  DFF \sreg_reg[2030]  ( .D(o[2031]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2030]) );
  DFF \sreg_reg[2031]  ( .D(o[2032]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2031]) );
  DFF \sreg_reg[2032]  ( .D(o[2033]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2032]) );
  DFF \sreg_reg[2033]  ( .D(o[2034]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2033]) );
  DFF \sreg_reg[2034]  ( .D(o[2035]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2034]) );
  DFF \sreg_reg[2035]  ( .D(o[2036]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2035]) );
  DFF \sreg_reg[2036]  ( .D(o[2037]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2036]) );
  DFF \sreg_reg[2037]  ( .D(o[2038]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2037]) );
  DFF \sreg_reg[2038]  ( .D(o[2039]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2038]) );
  DFF \sreg_reg[2039]  ( .D(o[2040]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2039]) );
  DFF \sreg_reg[2040]  ( .D(o[2041]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2040]) );
  DFF \sreg_reg[2041]  ( .D(o[2042]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2041]) );
  DFF \sreg_reg[2042]  ( .D(o[2043]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2042]) );
  DFF \sreg_reg[2043]  ( .D(o[2044]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2043]) );
  DFF \sreg_reg[2044]  ( .D(o[2045]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2044]) );
  DFF \sreg_reg[2045]  ( .D(o[2046]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2045]) );
  DFF \sreg_reg[2046]  ( .D(\add_42/carry[2047] ), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(sreg[2046]) );
  FADDER \add_42/U1_1024  ( .CIN(sreg[1024]), .IN0(n3072), .IN1(
        \add_42/carry[1024] ), .COUT(\add_42/carry[1025] ), .SUM(o[1024]) );
  FADDER \add_42/U1_1025  ( .CIN(sreg[1025]), .IN0(n3071), .IN1(
        \add_42/carry[1025] ), .COUT(\add_42/carry[1026] ), .SUM(o[1025]) );
  FADDER \add_42/U1_1026  ( .CIN(sreg[1026]), .IN0(n3070), .IN1(
        \add_42/carry[1026] ), .COUT(\add_42/carry[1027] ), .SUM(o[1026]) );
  FADDER \add_42/U1_1027  ( .CIN(sreg[1027]), .IN0(n3069), .IN1(
        \add_42/carry[1027] ), .COUT(\add_42/carry[1028] ), .SUM(o[1027]) );
  FADDER \add_42/U1_1028  ( .CIN(sreg[1028]), .IN0(n3068), .IN1(
        \add_42/carry[1028] ), .COUT(\add_42/carry[1029] ), .SUM(o[1028]) );
  FADDER \add_42/U1_1029  ( .CIN(sreg[1029]), .IN0(n3067), .IN1(
        \add_42/carry[1029] ), .COUT(\add_42/carry[1030] ), .SUM(o[1029]) );
  FADDER \add_42/U1_1030  ( .CIN(sreg[1030]), .IN0(n3066), .IN1(
        \add_42/carry[1030] ), .COUT(\add_42/carry[1031] ), .SUM(o[1030]) );
  FADDER \add_42/U1_1031  ( .CIN(sreg[1031]), .IN0(n3065), .IN1(
        \add_42/carry[1031] ), .COUT(\add_42/carry[1032] ), .SUM(o[1031]) );
  FADDER \add_42/U1_1032  ( .CIN(sreg[1032]), .IN0(n3064), .IN1(
        \add_42/carry[1032] ), .COUT(\add_42/carry[1033] ), .SUM(o[1032]) );
  FADDER \add_42/U1_1033  ( .CIN(sreg[1033]), .IN0(n3063), .IN1(
        \add_42/carry[1033] ), .COUT(\add_42/carry[1034] ), .SUM(o[1033]) );
  FADDER \add_42/U1_1034  ( .CIN(sreg[1034]), .IN0(n3062), .IN1(
        \add_42/carry[1034] ), .COUT(\add_42/carry[1035] ), .SUM(o[1034]) );
  FADDER \add_42/U1_1035  ( .CIN(sreg[1035]), .IN0(n3061), .IN1(
        \add_42/carry[1035] ), .COUT(\add_42/carry[1036] ), .SUM(o[1035]) );
  FADDER \add_42/U1_1036  ( .CIN(sreg[1036]), .IN0(n3060), .IN1(
        \add_42/carry[1036] ), .COUT(\add_42/carry[1037] ), .SUM(o[1036]) );
  FADDER \add_42/U1_1037  ( .CIN(sreg[1037]), .IN0(n3059), .IN1(
        \add_42/carry[1037] ), .COUT(\add_42/carry[1038] ), .SUM(o[1037]) );
  FADDER \add_42/U1_1038  ( .CIN(sreg[1038]), .IN0(n3058), .IN1(
        \add_42/carry[1038] ), .COUT(\add_42/carry[1039] ), .SUM(o[1038]) );
  FADDER \add_42/U1_1039  ( .CIN(sreg[1039]), .IN0(n3057), .IN1(
        \add_42/carry[1039] ), .COUT(\add_42/carry[1040] ), .SUM(o[1039]) );
  FADDER \add_42/U1_1040  ( .CIN(sreg[1040]), .IN0(n3056), .IN1(
        \add_42/carry[1040] ), .COUT(\add_42/carry[1041] ), .SUM(o[1040]) );
  FADDER \add_42/U1_1041  ( .CIN(sreg[1041]), .IN0(n3055), .IN1(
        \add_42/carry[1041] ), .COUT(\add_42/carry[1042] ), .SUM(o[1041]) );
  FADDER \add_42/U1_1042  ( .CIN(sreg[1042]), .IN0(n3054), .IN1(
        \add_42/carry[1042] ), .COUT(\add_42/carry[1043] ), .SUM(o[1042]) );
  FADDER \add_42/U1_1043  ( .CIN(sreg[1043]), .IN0(n3053), .IN1(
        \add_42/carry[1043] ), .COUT(\add_42/carry[1044] ), .SUM(o[1043]) );
  FADDER \add_42/U1_1044  ( .CIN(sreg[1044]), .IN0(n3052), .IN1(
        \add_42/carry[1044] ), .COUT(\add_42/carry[1045] ), .SUM(o[1044]) );
  FADDER \add_42/U1_1045  ( .CIN(sreg[1045]), .IN0(n3051), .IN1(
        \add_42/carry[1045] ), .COUT(\add_42/carry[1046] ), .SUM(o[1045]) );
  FADDER \add_42/U1_1046  ( .CIN(sreg[1046]), .IN0(n3050), .IN1(
        \add_42/carry[1046] ), .COUT(\add_42/carry[1047] ), .SUM(o[1046]) );
  FADDER \add_42/U1_1047  ( .CIN(sreg[1047]), .IN0(n3049), .IN1(
        \add_42/carry[1047] ), .COUT(\add_42/carry[1048] ), .SUM(o[1047]) );
  FADDER \add_42/U1_1048  ( .CIN(sreg[1048]), .IN0(n3048), .IN1(
        \add_42/carry[1048] ), .COUT(\add_42/carry[1049] ), .SUM(o[1048]) );
  FADDER \add_42/U1_1049  ( .CIN(sreg[1049]), .IN0(n3047), .IN1(
        \add_42/carry[1049] ), .COUT(\add_42/carry[1050] ), .SUM(o[1049]) );
  FADDER \add_42/U1_1050  ( .CIN(sreg[1050]), .IN0(n3046), .IN1(
        \add_42/carry[1050] ), .COUT(\add_42/carry[1051] ), .SUM(o[1050]) );
  FADDER \add_42/U1_1051  ( .CIN(sreg[1051]), .IN0(n3045), .IN1(
        \add_42/carry[1051] ), .COUT(\add_42/carry[1052] ), .SUM(o[1051]) );
  FADDER \add_42/U1_1052  ( .CIN(sreg[1052]), .IN0(n3044), .IN1(
        \add_42/carry[1052] ), .COUT(\add_42/carry[1053] ), .SUM(o[1052]) );
  FADDER \add_42/U1_1053  ( .CIN(sreg[1053]), .IN0(n3043), .IN1(
        \add_42/carry[1053] ), .COUT(\add_42/carry[1054] ), .SUM(o[1053]) );
  FADDER \add_42/U1_1054  ( .CIN(sreg[1054]), .IN0(n3042), .IN1(
        \add_42/carry[1054] ), .COUT(\add_42/carry[1055] ), .SUM(o[1054]) );
  FADDER \add_42/U1_1055  ( .CIN(sreg[1055]), .IN0(n3041), .IN1(
        \add_42/carry[1055] ), .COUT(\add_42/carry[1056] ), .SUM(o[1055]) );
  FADDER \add_42/U1_1056  ( .CIN(sreg[1056]), .IN0(n3040), .IN1(
        \add_42/carry[1056] ), .COUT(\add_42/carry[1057] ), .SUM(o[1056]) );
  FADDER \add_42/U1_1057  ( .CIN(sreg[1057]), .IN0(n3039), .IN1(
        \add_42/carry[1057] ), .COUT(\add_42/carry[1058] ), .SUM(o[1057]) );
  FADDER \add_42/U1_1058  ( .CIN(sreg[1058]), .IN0(n3038), .IN1(
        \add_42/carry[1058] ), .COUT(\add_42/carry[1059] ), .SUM(o[1058]) );
  FADDER \add_42/U1_1059  ( .CIN(sreg[1059]), .IN0(n3037), .IN1(
        \add_42/carry[1059] ), .COUT(\add_42/carry[1060] ), .SUM(o[1059]) );
  FADDER \add_42/U1_1060  ( .CIN(sreg[1060]), .IN0(n3036), .IN1(
        \add_42/carry[1060] ), .COUT(\add_42/carry[1061] ), .SUM(o[1060]) );
  FADDER \add_42/U1_1061  ( .CIN(sreg[1061]), .IN0(n3035), .IN1(
        \add_42/carry[1061] ), .COUT(\add_42/carry[1062] ), .SUM(o[1061]) );
  FADDER \add_42/U1_1062  ( .CIN(sreg[1062]), .IN0(n3034), .IN1(
        \add_42/carry[1062] ), .COUT(\add_42/carry[1063] ), .SUM(o[1062]) );
  FADDER \add_42/U1_1063  ( .CIN(sreg[1063]), .IN0(n3033), .IN1(
        \add_42/carry[1063] ), .COUT(\add_42/carry[1064] ), .SUM(o[1063]) );
  FADDER \add_42/U1_1064  ( .CIN(sreg[1064]), .IN0(n3032), .IN1(
        \add_42/carry[1064] ), .COUT(\add_42/carry[1065] ), .SUM(o[1064]) );
  FADDER \add_42/U1_1065  ( .CIN(sreg[1065]), .IN0(n3031), .IN1(
        \add_42/carry[1065] ), .COUT(\add_42/carry[1066] ), .SUM(o[1065]) );
  FADDER \add_42/U1_1066  ( .CIN(sreg[1066]), .IN0(n3030), .IN1(
        \add_42/carry[1066] ), .COUT(\add_42/carry[1067] ), .SUM(o[1066]) );
  FADDER \add_42/U1_1067  ( .CIN(sreg[1067]), .IN0(n3029), .IN1(
        \add_42/carry[1067] ), .COUT(\add_42/carry[1068] ), .SUM(o[1067]) );
  FADDER \add_42/U1_1068  ( .CIN(sreg[1068]), .IN0(n3028), .IN1(
        \add_42/carry[1068] ), .COUT(\add_42/carry[1069] ), .SUM(o[1068]) );
  FADDER \add_42/U1_1069  ( .CIN(sreg[1069]), .IN0(n3027), .IN1(
        \add_42/carry[1069] ), .COUT(\add_42/carry[1070] ), .SUM(o[1069]) );
  FADDER \add_42/U1_1070  ( .CIN(sreg[1070]), .IN0(n3026), .IN1(
        \add_42/carry[1070] ), .COUT(\add_42/carry[1071] ), .SUM(o[1070]) );
  FADDER \add_42/U1_1071  ( .CIN(sreg[1071]), .IN0(n3025), .IN1(
        \add_42/carry[1071] ), .COUT(\add_42/carry[1072] ), .SUM(o[1071]) );
  FADDER \add_42/U1_1072  ( .CIN(sreg[1072]), .IN0(n3024), .IN1(
        \add_42/carry[1072] ), .COUT(\add_42/carry[1073] ), .SUM(o[1072]) );
  FADDER \add_42/U1_1073  ( .CIN(sreg[1073]), .IN0(n3023), .IN1(
        \add_42/carry[1073] ), .COUT(\add_42/carry[1074] ), .SUM(o[1073]) );
  FADDER \add_42/U1_1074  ( .CIN(sreg[1074]), .IN0(n3022), .IN1(
        \add_42/carry[1074] ), .COUT(\add_42/carry[1075] ), .SUM(o[1074]) );
  FADDER \add_42/U1_1075  ( .CIN(sreg[1075]), .IN0(n3021), .IN1(
        \add_42/carry[1075] ), .COUT(\add_42/carry[1076] ), .SUM(o[1075]) );
  FADDER \add_42/U1_1076  ( .CIN(sreg[1076]), .IN0(n3020), .IN1(
        \add_42/carry[1076] ), .COUT(\add_42/carry[1077] ), .SUM(o[1076]) );
  FADDER \add_42/U1_1077  ( .CIN(sreg[1077]), .IN0(n3019), .IN1(
        \add_42/carry[1077] ), .COUT(\add_42/carry[1078] ), .SUM(o[1077]) );
  FADDER \add_42/U1_1078  ( .CIN(sreg[1078]), .IN0(n3018), .IN1(
        \add_42/carry[1078] ), .COUT(\add_42/carry[1079] ), .SUM(o[1078]) );
  FADDER \add_42/U1_1079  ( .CIN(sreg[1079]), .IN0(n3017), .IN1(
        \add_42/carry[1079] ), .COUT(\add_42/carry[1080] ), .SUM(o[1079]) );
  FADDER \add_42/U1_1080  ( .CIN(sreg[1080]), .IN0(n3016), .IN1(
        \add_42/carry[1080] ), .COUT(\add_42/carry[1081] ), .SUM(o[1080]) );
  FADDER \add_42/U1_1081  ( .CIN(sreg[1081]), .IN0(n3015), .IN1(
        \add_42/carry[1081] ), .COUT(\add_42/carry[1082] ), .SUM(o[1081]) );
  FADDER \add_42/U1_1082  ( .CIN(sreg[1082]), .IN0(n3014), .IN1(
        \add_42/carry[1082] ), .COUT(\add_42/carry[1083] ), .SUM(o[1082]) );
  FADDER \add_42/U1_1083  ( .CIN(sreg[1083]), .IN0(n3013), .IN1(
        \add_42/carry[1083] ), .COUT(\add_42/carry[1084] ), .SUM(o[1083]) );
  FADDER \add_42/U1_1084  ( .CIN(sreg[1084]), .IN0(n3012), .IN1(
        \add_42/carry[1084] ), .COUT(\add_42/carry[1085] ), .SUM(o[1084]) );
  FADDER \add_42/U1_1085  ( .CIN(sreg[1085]), .IN0(n3011), .IN1(
        \add_42/carry[1085] ), .COUT(\add_42/carry[1086] ), .SUM(o[1085]) );
  FADDER \add_42/U1_1086  ( .CIN(sreg[1086]), .IN0(n3010), .IN1(
        \add_42/carry[1086] ), .COUT(\add_42/carry[1087] ), .SUM(o[1086]) );
  FADDER \add_42/U1_1087  ( .CIN(sreg[1087]), .IN0(n3009), .IN1(
        \add_42/carry[1087] ), .COUT(\add_42/carry[1088] ), .SUM(o[1087]) );
  FADDER \add_42/U1_1088  ( .CIN(sreg[1088]), .IN0(n3008), .IN1(
        \add_42/carry[1088] ), .COUT(\add_42/carry[1089] ), .SUM(o[1088]) );
  FADDER \add_42/U1_1089  ( .CIN(sreg[1089]), .IN0(n3007), .IN1(
        \add_42/carry[1089] ), .COUT(\add_42/carry[1090] ), .SUM(o[1089]) );
  FADDER \add_42/U1_1090  ( .CIN(sreg[1090]), .IN0(n3006), .IN1(
        \add_42/carry[1090] ), .COUT(\add_42/carry[1091] ), .SUM(o[1090]) );
  FADDER \add_42/U1_1091  ( .CIN(sreg[1091]), .IN0(n3005), .IN1(
        \add_42/carry[1091] ), .COUT(\add_42/carry[1092] ), .SUM(o[1091]) );
  FADDER \add_42/U1_1092  ( .CIN(sreg[1092]), .IN0(n3004), .IN1(
        \add_42/carry[1092] ), .COUT(\add_42/carry[1093] ), .SUM(o[1092]) );
  FADDER \add_42/U1_1093  ( .CIN(sreg[1093]), .IN0(n3003), .IN1(
        \add_42/carry[1093] ), .COUT(\add_42/carry[1094] ), .SUM(o[1093]) );
  FADDER \add_42/U1_1094  ( .CIN(sreg[1094]), .IN0(n3002), .IN1(
        \add_42/carry[1094] ), .COUT(\add_42/carry[1095] ), .SUM(o[1094]) );
  FADDER \add_42/U1_1095  ( .CIN(sreg[1095]), .IN0(n3001), .IN1(
        \add_42/carry[1095] ), .COUT(\add_42/carry[1096] ), .SUM(o[1095]) );
  FADDER \add_42/U1_1096  ( .CIN(sreg[1096]), .IN0(n3000), .IN1(
        \add_42/carry[1096] ), .COUT(\add_42/carry[1097] ), .SUM(o[1096]) );
  FADDER \add_42/U1_1097  ( .CIN(sreg[1097]), .IN0(n2999), .IN1(
        \add_42/carry[1097] ), .COUT(\add_42/carry[1098] ), .SUM(o[1097]) );
  FADDER \add_42/U1_1098  ( .CIN(sreg[1098]), .IN0(n2998), .IN1(
        \add_42/carry[1098] ), .COUT(\add_42/carry[1099] ), .SUM(o[1098]) );
  FADDER \add_42/U1_1099  ( .CIN(sreg[1099]), .IN0(n2997), .IN1(
        \add_42/carry[1099] ), .COUT(\add_42/carry[1100] ), .SUM(o[1099]) );
  FADDER \add_42/U1_1100  ( .CIN(sreg[1100]), .IN0(n2996), .IN1(
        \add_42/carry[1100] ), .COUT(\add_42/carry[1101] ), .SUM(o[1100]) );
  FADDER \add_42/U1_1101  ( .CIN(sreg[1101]), .IN0(n2995), .IN1(
        \add_42/carry[1101] ), .COUT(\add_42/carry[1102] ), .SUM(o[1101]) );
  FADDER \add_42/U1_1102  ( .CIN(sreg[1102]), .IN0(n2994), .IN1(
        \add_42/carry[1102] ), .COUT(\add_42/carry[1103] ), .SUM(o[1102]) );
  FADDER \add_42/U1_1103  ( .CIN(sreg[1103]), .IN0(n2993), .IN1(
        \add_42/carry[1103] ), .COUT(\add_42/carry[1104] ), .SUM(o[1103]) );
  FADDER \add_42/U1_1104  ( .CIN(sreg[1104]), .IN0(n2992), .IN1(
        \add_42/carry[1104] ), .COUT(\add_42/carry[1105] ), .SUM(o[1104]) );
  FADDER \add_42/U1_1105  ( .CIN(sreg[1105]), .IN0(n2991), .IN1(
        \add_42/carry[1105] ), .COUT(\add_42/carry[1106] ), .SUM(o[1105]) );
  FADDER \add_42/U1_1106  ( .CIN(sreg[1106]), .IN0(n2990), .IN1(
        \add_42/carry[1106] ), .COUT(\add_42/carry[1107] ), .SUM(o[1106]) );
  FADDER \add_42/U1_1107  ( .CIN(sreg[1107]), .IN0(n2989), .IN1(
        \add_42/carry[1107] ), .COUT(\add_42/carry[1108] ), .SUM(o[1107]) );
  FADDER \add_42/U1_1108  ( .CIN(sreg[1108]), .IN0(n2988), .IN1(
        \add_42/carry[1108] ), .COUT(\add_42/carry[1109] ), .SUM(o[1108]) );
  FADDER \add_42/U1_1109  ( .CIN(sreg[1109]), .IN0(n2987), .IN1(
        \add_42/carry[1109] ), .COUT(\add_42/carry[1110] ), .SUM(o[1109]) );
  FADDER \add_42/U1_1110  ( .CIN(sreg[1110]), .IN0(n2986), .IN1(
        \add_42/carry[1110] ), .COUT(\add_42/carry[1111] ), .SUM(o[1110]) );
  FADDER \add_42/U1_1111  ( .CIN(sreg[1111]), .IN0(n2985), .IN1(
        \add_42/carry[1111] ), .COUT(\add_42/carry[1112] ), .SUM(o[1111]) );
  FADDER \add_42/U1_1112  ( .CIN(sreg[1112]), .IN0(n2984), .IN1(
        \add_42/carry[1112] ), .COUT(\add_42/carry[1113] ), .SUM(o[1112]) );
  FADDER \add_42/U1_1113  ( .CIN(sreg[1113]), .IN0(n2983), .IN1(
        \add_42/carry[1113] ), .COUT(\add_42/carry[1114] ), .SUM(o[1113]) );
  FADDER \add_42/U1_1114  ( .CIN(sreg[1114]), .IN0(n2982), .IN1(
        \add_42/carry[1114] ), .COUT(\add_42/carry[1115] ), .SUM(o[1114]) );
  FADDER \add_42/U1_1115  ( .CIN(sreg[1115]), .IN0(n2981), .IN1(
        \add_42/carry[1115] ), .COUT(\add_42/carry[1116] ), .SUM(o[1115]) );
  FADDER \add_42/U1_1116  ( .CIN(sreg[1116]), .IN0(n2980), .IN1(
        \add_42/carry[1116] ), .COUT(\add_42/carry[1117] ), .SUM(o[1116]) );
  FADDER \add_42/U1_1117  ( .CIN(sreg[1117]), .IN0(n2979), .IN1(
        \add_42/carry[1117] ), .COUT(\add_42/carry[1118] ), .SUM(o[1117]) );
  FADDER \add_42/U1_1118  ( .CIN(sreg[1118]), .IN0(n2978), .IN1(
        \add_42/carry[1118] ), .COUT(\add_42/carry[1119] ), .SUM(o[1118]) );
  FADDER \add_42/U1_1119  ( .CIN(sreg[1119]), .IN0(n2977), .IN1(
        \add_42/carry[1119] ), .COUT(\add_42/carry[1120] ), .SUM(o[1119]) );
  FADDER \add_42/U1_1120  ( .CIN(sreg[1120]), .IN0(n2976), .IN1(
        \add_42/carry[1120] ), .COUT(\add_42/carry[1121] ), .SUM(o[1120]) );
  FADDER \add_42/U1_1121  ( .CIN(sreg[1121]), .IN0(n2975), .IN1(
        \add_42/carry[1121] ), .COUT(\add_42/carry[1122] ), .SUM(o[1121]) );
  FADDER \add_42/U1_1122  ( .CIN(sreg[1122]), .IN0(n2974), .IN1(
        \add_42/carry[1122] ), .COUT(\add_42/carry[1123] ), .SUM(o[1122]) );
  FADDER \add_42/U1_1123  ( .CIN(sreg[1123]), .IN0(n2973), .IN1(
        \add_42/carry[1123] ), .COUT(\add_42/carry[1124] ), .SUM(o[1123]) );
  FADDER \add_42/U1_1124  ( .CIN(sreg[1124]), .IN0(n2972), .IN1(
        \add_42/carry[1124] ), .COUT(\add_42/carry[1125] ), .SUM(o[1124]) );
  FADDER \add_42/U1_1125  ( .CIN(sreg[1125]), .IN0(n2971), .IN1(
        \add_42/carry[1125] ), .COUT(\add_42/carry[1126] ), .SUM(o[1125]) );
  FADDER \add_42/U1_1126  ( .CIN(sreg[1126]), .IN0(n2970), .IN1(
        \add_42/carry[1126] ), .COUT(\add_42/carry[1127] ), .SUM(o[1126]) );
  FADDER \add_42/U1_1127  ( .CIN(sreg[1127]), .IN0(n2969), .IN1(
        \add_42/carry[1127] ), .COUT(\add_42/carry[1128] ), .SUM(o[1127]) );
  FADDER \add_42/U1_1128  ( .CIN(sreg[1128]), .IN0(n2968), .IN1(
        \add_42/carry[1128] ), .COUT(\add_42/carry[1129] ), .SUM(o[1128]) );
  FADDER \add_42/U1_1129  ( .CIN(sreg[1129]), .IN0(n2967), .IN1(
        \add_42/carry[1129] ), .COUT(\add_42/carry[1130] ), .SUM(o[1129]) );
  FADDER \add_42/U1_1130  ( .CIN(sreg[1130]), .IN0(n2966), .IN1(
        \add_42/carry[1130] ), .COUT(\add_42/carry[1131] ), .SUM(o[1130]) );
  FADDER \add_42/U1_1131  ( .CIN(sreg[1131]), .IN0(n2965), .IN1(
        \add_42/carry[1131] ), .COUT(\add_42/carry[1132] ), .SUM(o[1131]) );
  FADDER \add_42/U1_1132  ( .CIN(sreg[1132]), .IN0(n2964), .IN1(
        \add_42/carry[1132] ), .COUT(\add_42/carry[1133] ), .SUM(o[1132]) );
  FADDER \add_42/U1_1133  ( .CIN(sreg[1133]), .IN0(n2963), .IN1(
        \add_42/carry[1133] ), .COUT(\add_42/carry[1134] ), .SUM(o[1133]) );
  FADDER \add_42/U1_1134  ( .CIN(sreg[1134]), .IN0(n2962), .IN1(
        \add_42/carry[1134] ), .COUT(\add_42/carry[1135] ), .SUM(o[1134]) );
  FADDER \add_42/U1_1135  ( .CIN(sreg[1135]), .IN0(n2961), .IN1(
        \add_42/carry[1135] ), .COUT(\add_42/carry[1136] ), .SUM(o[1135]) );
  FADDER \add_42/U1_1136  ( .CIN(sreg[1136]), .IN0(n2960), .IN1(
        \add_42/carry[1136] ), .COUT(\add_42/carry[1137] ), .SUM(o[1136]) );
  FADDER \add_42/U1_1137  ( .CIN(sreg[1137]), .IN0(n2959), .IN1(
        \add_42/carry[1137] ), .COUT(\add_42/carry[1138] ), .SUM(o[1137]) );
  FADDER \add_42/U1_1138  ( .CIN(sreg[1138]), .IN0(n2958), .IN1(
        \add_42/carry[1138] ), .COUT(\add_42/carry[1139] ), .SUM(o[1138]) );
  FADDER \add_42/U1_1139  ( .CIN(sreg[1139]), .IN0(n2957), .IN1(
        \add_42/carry[1139] ), .COUT(\add_42/carry[1140] ), .SUM(o[1139]) );
  FADDER \add_42/U1_1140  ( .CIN(sreg[1140]), .IN0(n2956), .IN1(
        \add_42/carry[1140] ), .COUT(\add_42/carry[1141] ), .SUM(o[1140]) );
  FADDER \add_42/U1_1141  ( .CIN(sreg[1141]), .IN0(n2955), .IN1(
        \add_42/carry[1141] ), .COUT(\add_42/carry[1142] ), .SUM(o[1141]) );
  FADDER \add_42/U1_1142  ( .CIN(sreg[1142]), .IN0(n2954), .IN1(
        \add_42/carry[1142] ), .COUT(\add_42/carry[1143] ), .SUM(o[1142]) );
  FADDER \add_42/U1_1143  ( .CIN(sreg[1143]), .IN0(n2953), .IN1(
        \add_42/carry[1143] ), .COUT(\add_42/carry[1144] ), .SUM(o[1143]) );
  FADDER \add_42/U1_1144  ( .CIN(sreg[1144]), .IN0(n2952), .IN1(
        \add_42/carry[1144] ), .COUT(\add_42/carry[1145] ), .SUM(o[1144]) );
  FADDER \add_42/U1_1145  ( .CIN(sreg[1145]), .IN0(n2951), .IN1(
        \add_42/carry[1145] ), .COUT(\add_42/carry[1146] ), .SUM(o[1145]) );
  FADDER \add_42/U1_1146  ( .CIN(sreg[1146]), .IN0(n2950), .IN1(
        \add_42/carry[1146] ), .COUT(\add_42/carry[1147] ), .SUM(o[1146]) );
  FADDER \add_42/U1_1147  ( .CIN(sreg[1147]), .IN0(n2949), .IN1(
        \add_42/carry[1147] ), .COUT(\add_42/carry[1148] ), .SUM(o[1147]) );
  FADDER \add_42/U1_1148  ( .CIN(sreg[1148]), .IN0(n2948), .IN1(
        \add_42/carry[1148] ), .COUT(\add_42/carry[1149] ), .SUM(o[1148]) );
  FADDER \add_42/U1_1149  ( .CIN(sreg[1149]), .IN0(n2947), .IN1(
        \add_42/carry[1149] ), .COUT(\add_42/carry[1150] ), .SUM(o[1149]) );
  FADDER \add_42/U1_1150  ( .CIN(sreg[1150]), .IN0(n2946), .IN1(
        \add_42/carry[1150] ), .COUT(\add_42/carry[1151] ), .SUM(o[1150]) );
  FADDER \add_42/U1_1151  ( .CIN(sreg[1151]), .IN0(n2945), .IN1(
        \add_42/carry[1151] ), .COUT(\add_42/carry[1152] ), .SUM(o[1151]) );
  FADDER \add_42/U1_1152  ( .CIN(sreg[1152]), .IN0(n2944), .IN1(
        \add_42/carry[1152] ), .COUT(\add_42/carry[1153] ), .SUM(o[1152]) );
  FADDER \add_42/U1_1153  ( .CIN(sreg[1153]), .IN0(n2943), .IN1(
        \add_42/carry[1153] ), .COUT(\add_42/carry[1154] ), .SUM(o[1153]) );
  FADDER \add_42/U1_1154  ( .CIN(sreg[1154]), .IN0(n2942), .IN1(
        \add_42/carry[1154] ), .COUT(\add_42/carry[1155] ), .SUM(o[1154]) );
  FADDER \add_42/U1_1155  ( .CIN(sreg[1155]), .IN0(n2941), .IN1(
        \add_42/carry[1155] ), .COUT(\add_42/carry[1156] ), .SUM(o[1155]) );
  FADDER \add_42/U1_1156  ( .CIN(sreg[1156]), .IN0(n2940), .IN1(
        \add_42/carry[1156] ), .COUT(\add_42/carry[1157] ), .SUM(o[1156]) );
  FADDER \add_42/U1_1157  ( .CIN(sreg[1157]), .IN0(n2939), .IN1(
        \add_42/carry[1157] ), .COUT(\add_42/carry[1158] ), .SUM(o[1157]) );
  FADDER \add_42/U1_1158  ( .CIN(sreg[1158]), .IN0(n2938), .IN1(
        \add_42/carry[1158] ), .COUT(\add_42/carry[1159] ), .SUM(o[1158]) );
  FADDER \add_42/U1_1159  ( .CIN(sreg[1159]), .IN0(n2937), .IN1(
        \add_42/carry[1159] ), .COUT(\add_42/carry[1160] ), .SUM(o[1159]) );
  FADDER \add_42/U1_1160  ( .CIN(sreg[1160]), .IN0(n2936), .IN1(
        \add_42/carry[1160] ), .COUT(\add_42/carry[1161] ), .SUM(o[1160]) );
  FADDER \add_42/U1_1161  ( .CIN(sreg[1161]), .IN0(n2935), .IN1(
        \add_42/carry[1161] ), .COUT(\add_42/carry[1162] ), .SUM(o[1161]) );
  FADDER \add_42/U1_1162  ( .CIN(sreg[1162]), .IN0(n2934), .IN1(
        \add_42/carry[1162] ), .COUT(\add_42/carry[1163] ), .SUM(o[1162]) );
  FADDER \add_42/U1_1163  ( .CIN(sreg[1163]), .IN0(n2933), .IN1(
        \add_42/carry[1163] ), .COUT(\add_42/carry[1164] ), .SUM(o[1163]) );
  FADDER \add_42/U1_1164  ( .CIN(sreg[1164]), .IN0(n2932), .IN1(
        \add_42/carry[1164] ), .COUT(\add_42/carry[1165] ), .SUM(o[1164]) );
  FADDER \add_42/U1_1165  ( .CIN(sreg[1165]), .IN0(n2931), .IN1(
        \add_42/carry[1165] ), .COUT(\add_42/carry[1166] ), .SUM(o[1165]) );
  FADDER \add_42/U1_1166  ( .CIN(sreg[1166]), .IN0(n2930), .IN1(
        \add_42/carry[1166] ), .COUT(\add_42/carry[1167] ), .SUM(o[1166]) );
  FADDER \add_42/U1_1167  ( .CIN(sreg[1167]), .IN0(n2929), .IN1(
        \add_42/carry[1167] ), .COUT(\add_42/carry[1168] ), .SUM(o[1167]) );
  FADDER \add_42/U1_1168  ( .CIN(sreg[1168]), .IN0(n2928), .IN1(
        \add_42/carry[1168] ), .COUT(\add_42/carry[1169] ), .SUM(o[1168]) );
  FADDER \add_42/U1_1169  ( .CIN(sreg[1169]), .IN0(n2927), .IN1(
        \add_42/carry[1169] ), .COUT(\add_42/carry[1170] ), .SUM(o[1169]) );
  FADDER \add_42/U1_1170  ( .CIN(sreg[1170]), .IN0(n2926), .IN1(
        \add_42/carry[1170] ), .COUT(\add_42/carry[1171] ), .SUM(o[1170]) );
  FADDER \add_42/U1_1171  ( .CIN(sreg[1171]), .IN0(n2925), .IN1(
        \add_42/carry[1171] ), .COUT(\add_42/carry[1172] ), .SUM(o[1171]) );
  FADDER \add_42/U1_1172  ( .CIN(sreg[1172]), .IN0(n2924), .IN1(
        \add_42/carry[1172] ), .COUT(\add_42/carry[1173] ), .SUM(o[1172]) );
  FADDER \add_42/U1_1173  ( .CIN(sreg[1173]), .IN0(n2923), .IN1(
        \add_42/carry[1173] ), .COUT(\add_42/carry[1174] ), .SUM(o[1173]) );
  FADDER \add_42/U1_1174  ( .CIN(sreg[1174]), .IN0(n2922), .IN1(
        \add_42/carry[1174] ), .COUT(\add_42/carry[1175] ), .SUM(o[1174]) );
  FADDER \add_42/U1_1175  ( .CIN(sreg[1175]), .IN0(n2921), .IN1(
        \add_42/carry[1175] ), .COUT(\add_42/carry[1176] ), .SUM(o[1175]) );
  FADDER \add_42/U1_1176  ( .CIN(sreg[1176]), .IN0(n2920), .IN1(
        \add_42/carry[1176] ), .COUT(\add_42/carry[1177] ), .SUM(o[1176]) );
  FADDER \add_42/U1_1177  ( .CIN(sreg[1177]), .IN0(n2919), .IN1(
        \add_42/carry[1177] ), .COUT(\add_42/carry[1178] ), .SUM(o[1177]) );
  FADDER \add_42/U1_1178  ( .CIN(sreg[1178]), .IN0(n2918), .IN1(
        \add_42/carry[1178] ), .COUT(\add_42/carry[1179] ), .SUM(o[1178]) );
  FADDER \add_42/U1_1179  ( .CIN(sreg[1179]), .IN0(n2917), .IN1(
        \add_42/carry[1179] ), .COUT(\add_42/carry[1180] ), .SUM(o[1179]) );
  FADDER \add_42/U1_1180  ( .CIN(sreg[1180]), .IN0(n2916), .IN1(
        \add_42/carry[1180] ), .COUT(\add_42/carry[1181] ), .SUM(o[1180]) );
  FADDER \add_42/U1_1181  ( .CIN(sreg[1181]), .IN0(n2915), .IN1(
        \add_42/carry[1181] ), .COUT(\add_42/carry[1182] ), .SUM(o[1181]) );
  FADDER \add_42/U1_1182  ( .CIN(sreg[1182]), .IN0(n2914), .IN1(
        \add_42/carry[1182] ), .COUT(\add_42/carry[1183] ), .SUM(o[1182]) );
  FADDER \add_42/U1_1183  ( .CIN(sreg[1183]), .IN0(n2913), .IN1(
        \add_42/carry[1183] ), .COUT(\add_42/carry[1184] ), .SUM(o[1183]) );
  FADDER \add_42/U1_1184  ( .CIN(sreg[1184]), .IN0(n2912), .IN1(
        \add_42/carry[1184] ), .COUT(\add_42/carry[1185] ), .SUM(o[1184]) );
  FADDER \add_42/U1_1185  ( .CIN(sreg[1185]), .IN0(n2911), .IN1(
        \add_42/carry[1185] ), .COUT(\add_42/carry[1186] ), .SUM(o[1185]) );
  FADDER \add_42/U1_1186  ( .CIN(sreg[1186]), .IN0(n2910), .IN1(
        \add_42/carry[1186] ), .COUT(\add_42/carry[1187] ), .SUM(o[1186]) );
  FADDER \add_42/U1_1187  ( .CIN(sreg[1187]), .IN0(n2909), .IN1(
        \add_42/carry[1187] ), .COUT(\add_42/carry[1188] ), .SUM(o[1187]) );
  FADDER \add_42/U1_1188  ( .CIN(sreg[1188]), .IN0(n2908), .IN1(
        \add_42/carry[1188] ), .COUT(\add_42/carry[1189] ), .SUM(o[1188]) );
  FADDER \add_42/U1_1189  ( .CIN(sreg[1189]), .IN0(n2907), .IN1(
        \add_42/carry[1189] ), .COUT(\add_42/carry[1190] ), .SUM(o[1189]) );
  FADDER \add_42/U1_1190  ( .CIN(sreg[1190]), .IN0(n2906), .IN1(
        \add_42/carry[1190] ), .COUT(\add_42/carry[1191] ), .SUM(o[1190]) );
  FADDER \add_42/U1_1191  ( .CIN(sreg[1191]), .IN0(n2905), .IN1(
        \add_42/carry[1191] ), .COUT(\add_42/carry[1192] ), .SUM(o[1191]) );
  FADDER \add_42/U1_1192  ( .CIN(sreg[1192]), .IN0(n2904), .IN1(
        \add_42/carry[1192] ), .COUT(\add_42/carry[1193] ), .SUM(o[1192]) );
  FADDER \add_42/U1_1193  ( .CIN(sreg[1193]), .IN0(n2903), .IN1(
        \add_42/carry[1193] ), .COUT(\add_42/carry[1194] ), .SUM(o[1193]) );
  FADDER \add_42/U1_1194  ( .CIN(sreg[1194]), .IN0(n2902), .IN1(
        \add_42/carry[1194] ), .COUT(\add_42/carry[1195] ), .SUM(o[1194]) );
  FADDER \add_42/U1_1195  ( .CIN(sreg[1195]), .IN0(n2901), .IN1(
        \add_42/carry[1195] ), .COUT(\add_42/carry[1196] ), .SUM(o[1195]) );
  FADDER \add_42/U1_1196  ( .CIN(sreg[1196]), .IN0(n2900), .IN1(
        \add_42/carry[1196] ), .COUT(\add_42/carry[1197] ), .SUM(o[1196]) );
  FADDER \add_42/U1_1197  ( .CIN(sreg[1197]), .IN0(n2899), .IN1(
        \add_42/carry[1197] ), .COUT(\add_42/carry[1198] ), .SUM(o[1197]) );
  FADDER \add_42/U1_1198  ( .CIN(sreg[1198]), .IN0(n2898), .IN1(
        \add_42/carry[1198] ), .COUT(\add_42/carry[1199] ), .SUM(o[1198]) );
  FADDER \add_42/U1_1199  ( .CIN(sreg[1199]), .IN0(n2897), .IN1(
        \add_42/carry[1199] ), .COUT(\add_42/carry[1200] ), .SUM(o[1199]) );
  FADDER \add_42/U1_1200  ( .CIN(sreg[1200]), .IN0(n2896), .IN1(
        \add_42/carry[1200] ), .COUT(\add_42/carry[1201] ), .SUM(o[1200]) );
  FADDER \add_42/U1_1201  ( .CIN(sreg[1201]), .IN0(n2895), .IN1(
        \add_42/carry[1201] ), .COUT(\add_42/carry[1202] ), .SUM(o[1201]) );
  FADDER \add_42/U1_1202  ( .CIN(sreg[1202]), .IN0(n2894), .IN1(
        \add_42/carry[1202] ), .COUT(\add_42/carry[1203] ), .SUM(o[1202]) );
  FADDER \add_42/U1_1203  ( .CIN(sreg[1203]), .IN0(n2893), .IN1(
        \add_42/carry[1203] ), .COUT(\add_42/carry[1204] ), .SUM(o[1203]) );
  FADDER \add_42/U1_1204  ( .CIN(sreg[1204]), .IN0(n2892), .IN1(
        \add_42/carry[1204] ), .COUT(\add_42/carry[1205] ), .SUM(o[1204]) );
  FADDER \add_42/U1_1205  ( .CIN(sreg[1205]), .IN0(n2891), .IN1(
        \add_42/carry[1205] ), .COUT(\add_42/carry[1206] ), .SUM(o[1205]) );
  FADDER \add_42/U1_1206  ( .CIN(sreg[1206]), .IN0(n2890), .IN1(
        \add_42/carry[1206] ), .COUT(\add_42/carry[1207] ), .SUM(o[1206]) );
  FADDER \add_42/U1_1207  ( .CIN(sreg[1207]), .IN0(n2889), .IN1(
        \add_42/carry[1207] ), .COUT(\add_42/carry[1208] ), .SUM(o[1207]) );
  FADDER \add_42/U1_1208  ( .CIN(sreg[1208]), .IN0(n2888), .IN1(
        \add_42/carry[1208] ), .COUT(\add_42/carry[1209] ), .SUM(o[1208]) );
  FADDER \add_42/U1_1209  ( .CIN(sreg[1209]), .IN0(n2887), .IN1(
        \add_42/carry[1209] ), .COUT(\add_42/carry[1210] ), .SUM(o[1209]) );
  FADDER \add_42/U1_1210  ( .CIN(sreg[1210]), .IN0(n2886), .IN1(
        \add_42/carry[1210] ), .COUT(\add_42/carry[1211] ), .SUM(o[1210]) );
  FADDER \add_42/U1_1211  ( .CIN(sreg[1211]), .IN0(n2885), .IN1(
        \add_42/carry[1211] ), .COUT(\add_42/carry[1212] ), .SUM(o[1211]) );
  FADDER \add_42/U1_1212  ( .CIN(sreg[1212]), .IN0(n2884), .IN1(
        \add_42/carry[1212] ), .COUT(\add_42/carry[1213] ), .SUM(o[1212]) );
  FADDER \add_42/U1_1213  ( .CIN(sreg[1213]), .IN0(n2883), .IN1(
        \add_42/carry[1213] ), .COUT(\add_42/carry[1214] ), .SUM(o[1213]) );
  FADDER \add_42/U1_1214  ( .CIN(sreg[1214]), .IN0(n2882), .IN1(
        \add_42/carry[1214] ), .COUT(\add_42/carry[1215] ), .SUM(o[1214]) );
  FADDER \add_42/U1_1215  ( .CIN(sreg[1215]), .IN0(n2881), .IN1(
        \add_42/carry[1215] ), .COUT(\add_42/carry[1216] ), .SUM(o[1215]) );
  FADDER \add_42/U1_1216  ( .CIN(sreg[1216]), .IN0(n2880), .IN1(
        \add_42/carry[1216] ), .COUT(\add_42/carry[1217] ), .SUM(o[1216]) );
  FADDER \add_42/U1_1217  ( .CIN(sreg[1217]), .IN0(n2879), .IN1(
        \add_42/carry[1217] ), .COUT(\add_42/carry[1218] ), .SUM(o[1217]) );
  FADDER \add_42/U1_1218  ( .CIN(sreg[1218]), .IN0(n2878), .IN1(
        \add_42/carry[1218] ), .COUT(\add_42/carry[1219] ), .SUM(o[1218]) );
  FADDER \add_42/U1_1219  ( .CIN(sreg[1219]), .IN0(n2877), .IN1(
        \add_42/carry[1219] ), .COUT(\add_42/carry[1220] ), .SUM(o[1219]) );
  FADDER \add_42/U1_1220  ( .CIN(sreg[1220]), .IN0(n2876), .IN1(
        \add_42/carry[1220] ), .COUT(\add_42/carry[1221] ), .SUM(o[1220]) );
  FADDER \add_42/U1_1221  ( .CIN(sreg[1221]), .IN0(n2875), .IN1(
        \add_42/carry[1221] ), .COUT(\add_42/carry[1222] ), .SUM(o[1221]) );
  FADDER \add_42/U1_1222  ( .CIN(sreg[1222]), .IN0(n2874), .IN1(
        \add_42/carry[1222] ), .COUT(\add_42/carry[1223] ), .SUM(o[1222]) );
  FADDER \add_42/U1_1223  ( .CIN(sreg[1223]), .IN0(n2873), .IN1(
        \add_42/carry[1223] ), .COUT(\add_42/carry[1224] ), .SUM(o[1223]) );
  FADDER \add_42/U1_1224  ( .CIN(sreg[1224]), .IN0(n2872), .IN1(
        \add_42/carry[1224] ), .COUT(\add_42/carry[1225] ), .SUM(o[1224]) );
  FADDER \add_42/U1_1225  ( .CIN(sreg[1225]), .IN0(n2871), .IN1(
        \add_42/carry[1225] ), .COUT(\add_42/carry[1226] ), .SUM(o[1225]) );
  FADDER \add_42/U1_1226  ( .CIN(sreg[1226]), .IN0(n2870), .IN1(
        \add_42/carry[1226] ), .COUT(\add_42/carry[1227] ), .SUM(o[1226]) );
  FADDER \add_42/U1_1227  ( .CIN(sreg[1227]), .IN0(n2869), .IN1(
        \add_42/carry[1227] ), .COUT(\add_42/carry[1228] ), .SUM(o[1227]) );
  FADDER \add_42/U1_1228  ( .CIN(sreg[1228]), .IN0(n2868), .IN1(
        \add_42/carry[1228] ), .COUT(\add_42/carry[1229] ), .SUM(o[1228]) );
  FADDER \add_42/U1_1229  ( .CIN(sreg[1229]), .IN0(n2867), .IN1(
        \add_42/carry[1229] ), .COUT(\add_42/carry[1230] ), .SUM(o[1229]) );
  FADDER \add_42/U1_1230  ( .CIN(sreg[1230]), .IN0(n2866), .IN1(
        \add_42/carry[1230] ), .COUT(\add_42/carry[1231] ), .SUM(o[1230]) );
  FADDER \add_42/U1_1231  ( .CIN(sreg[1231]), .IN0(n2865), .IN1(
        \add_42/carry[1231] ), .COUT(\add_42/carry[1232] ), .SUM(o[1231]) );
  FADDER \add_42/U1_1232  ( .CIN(sreg[1232]), .IN0(n2864), .IN1(
        \add_42/carry[1232] ), .COUT(\add_42/carry[1233] ), .SUM(o[1232]) );
  FADDER \add_42/U1_1233  ( .CIN(sreg[1233]), .IN0(n2863), .IN1(
        \add_42/carry[1233] ), .COUT(\add_42/carry[1234] ), .SUM(o[1233]) );
  FADDER \add_42/U1_1234  ( .CIN(sreg[1234]), .IN0(n2862), .IN1(
        \add_42/carry[1234] ), .COUT(\add_42/carry[1235] ), .SUM(o[1234]) );
  FADDER \add_42/U1_1235  ( .CIN(sreg[1235]), .IN0(n2861), .IN1(
        \add_42/carry[1235] ), .COUT(\add_42/carry[1236] ), .SUM(o[1235]) );
  FADDER \add_42/U1_1236  ( .CIN(sreg[1236]), .IN0(n2860), .IN1(
        \add_42/carry[1236] ), .COUT(\add_42/carry[1237] ), .SUM(o[1236]) );
  FADDER \add_42/U1_1237  ( .CIN(sreg[1237]), .IN0(n2859), .IN1(
        \add_42/carry[1237] ), .COUT(\add_42/carry[1238] ), .SUM(o[1237]) );
  FADDER \add_42/U1_1238  ( .CIN(sreg[1238]), .IN0(n2858), .IN1(
        \add_42/carry[1238] ), .COUT(\add_42/carry[1239] ), .SUM(o[1238]) );
  FADDER \add_42/U1_1239  ( .CIN(sreg[1239]), .IN0(n2857), .IN1(
        \add_42/carry[1239] ), .COUT(\add_42/carry[1240] ), .SUM(o[1239]) );
  FADDER \add_42/U1_1240  ( .CIN(sreg[1240]), .IN0(n2856), .IN1(
        \add_42/carry[1240] ), .COUT(\add_42/carry[1241] ), .SUM(o[1240]) );
  FADDER \add_42/U1_1241  ( .CIN(sreg[1241]), .IN0(n2855), .IN1(
        \add_42/carry[1241] ), .COUT(\add_42/carry[1242] ), .SUM(o[1241]) );
  FADDER \add_42/U1_1242  ( .CIN(sreg[1242]), .IN0(n2854), .IN1(
        \add_42/carry[1242] ), .COUT(\add_42/carry[1243] ), .SUM(o[1242]) );
  FADDER \add_42/U1_1243  ( .CIN(sreg[1243]), .IN0(n2853), .IN1(
        \add_42/carry[1243] ), .COUT(\add_42/carry[1244] ), .SUM(o[1243]) );
  FADDER \add_42/U1_1244  ( .CIN(sreg[1244]), .IN0(n2852), .IN1(
        \add_42/carry[1244] ), .COUT(\add_42/carry[1245] ), .SUM(o[1244]) );
  FADDER \add_42/U1_1245  ( .CIN(sreg[1245]), .IN0(n2851), .IN1(
        \add_42/carry[1245] ), .COUT(\add_42/carry[1246] ), .SUM(o[1245]) );
  FADDER \add_42/U1_1246  ( .CIN(sreg[1246]), .IN0(n2850), .IN1(
        \add_42/carry[1246] ), .COUT(\add_42/carry[1247] ), .SUM(o[1246]) );
  FADDER \add_42/U1_1247  ( .CIN(sreg[1247]), .IN0(n2849), .IN1(
        \add_42/carry[1247] ), .COUT(\add_42/carry[1248] ), .SUM(o[1247]) );
  FADDER \add_42/U1_1248  ( .CIN(sreg[1248]), .IN0(n2848), .IN1(
        \add_42/carry[1248] ), .COUT(\add_42/carry[1249] ), .SUM(o[1248]) );
  FADDER \add_42/U1_1249  ( .CIN(sreg[1249]), .IN0(n2847), .IN1(
        \add_42/carry[1249] ), .COUT(\add_42/carry[1250] ), .SUM(o[1249]) );
  FADDER \add_42/U1_1250  ( .CIN(sreg[1250]), .IN0(n2846), .IN1(
        \add_42/carry[1250] ), .COUT(\add_42/carry[1251] ), .SUM(o[1250]) );
  FADDER \add_42/U1_1251  ( .CIN(sreg[1251]), .IN0(n2845), .IN1(
        \add_42/carry[1251] ), .COUT(\add_42/carry[1252] ), .SUM(o[1251]) );
  FADDER \add_42/U1_1252  ( .CIN(sreg[1252]), .IN0(n2844), .IN1(
        \add_42/carry[1252] ), .COUT(\add_42/carry[1253] ), .SUM(o[1252]) );
  FADDER \add_42/U1_1253  ( .CIN(sreg[1253]), .IN0(n2843), .IN1(
        \add_42/carry[1253] ), .COUT(\add_42/carry[1254] ), .SUM(o[1253]) );
  FADDER \add_42/U1_1254  ( .CIN(sreg[1254]), .IN0(n2842), .IN1(
        \add_42/carry[1254] ), .COUT(\add_42/carry[1255] ), .SUM(o[1254]) );
  FADDER \add_42/U1_1255  ( .CIN(sreg[1255]), .IN0(n2841), .IN1(
        \add_42/carry[1255] ), .COUT(\add_42/carry[1256] ), .SUM(o[1255]) );
  FADDER \add_42/U1_1256  ( .CIN(sreg[1256]), .IN0(n2840), .IN1(
        \add_42/carry[1256] ), .COUT(\add_42/carry[1257] ), .SUM(o[1256]) );
  FADDER \add_42/U1_1257  ( .CIN(sreg[1257]), .IN0(n2839), .IN1(
        \add_42/carry[1257] ), .COUT(\add_42/carry[1258] ), .SUM(o[1257]) );
  FADDER \add_42/U1_1258  ( .CIN(sreg[1258]), .IN0(n2838), .IN1(
        \add_42/carry[1258] ), .COUT(\add_42/carry[1259] ), .SUM(o[1258]) );
  FADDER \add_42/U1_1259  ( .CIN(sreg[1259]), .IN0(n2837), .IN1(
        \add_42/carry[1259] ), .COUT(\add_42/carry[1260] ), .SUM(o[1259]) );
  FADDER \add_42/U1_1260  ( .CIN(sreg[1260]), .IN0(n2836), .IN1(
        \add_42/carry[1260] ), .COUT(\add_42/carry[1261] ), .SUM(o[1260]) );
  FADDER \add_42/U1_1261  ( .CIN(sreg[1261]), .IN0(n2835), .IN1(
        \add_42/carry[1261] ), .COUT(\add_42/carry[1262] ), .SUM(o[1261]) );
  FADDER \add_42/U1_1262  ( .CIN(sreg[1262]), .IN0(n2834), .IN1(
        \add_42/carry[1262] ), .COUT(\add_42/carry[1263] ), .SUM(o[1262]) );
  FADDER \add_42/U1_1263  ( .CIN(sreg[1263]), .IN0(n2833), .IN1(
        \add_42/carry[1263] ), .COUT(\add_42/carry[1264] ), .SUM(o[1263]) );
  FADDER \add_42/U1_1264  ( .CIN(sreg[1264]), .IN0(n2832), .IN1(
        \add_42/carry[1264] ), .COUT(\add_42/carry[1265] ), .SUM(o[1264]) );
  FADDER \add_42/U1_1265  ( .CIN(sreg[1265]), .IN0(n2831), .IN1(
        \add_42/carry[1265] ), .COUT(\add_42/carry[1266] ), .SUM(o[1265]) );
  FADDER \add_42/U1_1266  ( .CIN(sreg[1266]), .IN0(n2830), .IN1(
        \add_42/carry[1266] ), .COUT(\add_42/carry[1267] ), .SUM(o[1266]) );
  FADDER \add_42/U1_1267  ( .CIN(sreg[1267]), .IN0(n2829), .IN1(
        \add_42/carry[1267] ), .COUT(\add_42/carry[1268] ), .SUM(o[1267]) );
  FADDER \add_42/U1_1268  ( .CIN(sreg[1268]), .IN0(n2828), .IN1(
        \add_42/carry[1268] ), .COUT(\add_42/carry[1269] ), .SUM(o[1268]) );
  FADDER \add_42/U1_1269  ( .CIN(sreg[1269]), .IN0(n2827), .IN1(
        \add_42/carry[1269] ), .COUT(\add_42/carry[1270] ), .SUM(o[1269]) );
  FADDER \add_42/U1_1270  ( .CIN(sreg[1270]), .IN0(n2826), .IN1(
        \add_42/carry[1270] ), .COUT(\add_42/carry[1271] ), .SUM(o[1270]) );
  FADDER \add_42/U1_1271  ( .CIN(sreg[1271]), .IN0(n2825), .IN1(
        \add_42/carry[1271] ), .COUT(\add_42/carry[1272] ), .SUM(o[1271]) );
  FADDER \add_42/U1_1272  ( .CIN(sreg[1272]), .IN0(n2824), .IN1(
        \add_42/carry[1272] ), .COUT(\add_42/carry[1273] ), .SUM(o[1272]) );
  FADDER \add_42/U1_1273  ( .CIN(sreg[1273]), .IN0(n2823), .IN1(
        \add_42/carry[1273] ), .COUT(\add_42/carry[1274] ), .SUM(o[1273]) );
  FADDER \add_42/U1_1274  ( .CIN(sreg[1274]), .IN0(n2822), .IN1(
        \add_42/carry[1274] ), .COUT(\add_42/carry[1275] ), .SUM(o[1274]) );
  FADDER \add_42/U1_1275  ( .CIN(sreg[1275]), .IN0(n2821), .IN1(
        \add_42/carry[1275] ), .COUT(\add_42/carry[1276] ), .SUM(o[1275]) );
  FADDER \add_42/U1_1276  ( .CIN(sreg[1276]), .IN0(n2820), .IN1(
        \add_42/carry[1276] ), .COUT(\add_42/carry[1277] ), .SUM(o[1276]) );
  FADDER \add_42/U1_1277  ( .CIN(sreg[1277]), .IN0(n2819), .IN1(
        \add_42/carry[1277] ), .COUT(\add_42/carry[1278] ), .SUM(o[1277]) );
  FADDER \add_42/U1_1278  ( .CIN(sreg[1278]), .IN0(n2818), .IN1(
        \add_42/carry[1278] ), .COUT(\add_42/carry[1279] ), .SUM(o[1278]) );
  FADDER \add_42/U1_1279  ( .CIN(sreg[1279]), .IN0(n2817), .IN1(
        \add_42/carry[1279] ), .COUT(\add_42/carry[1280] ), .SUM(o[1279]) );
  FADDER \add_42/U1_1280  ( .CIN(sreg[1280]), .IN0(n2816), .IN1(
        \add_42/carry[1280] ), .COUT(\add_42/carry[1281] ), .SUM(o[1280]) );
  FADDER \add_42/U1_1281  ( .CIN(sreg[1281]), .IN0(n2815), .IN1(
        \add_42/carry[1281] ), .COUT(\add_42/carry[1282] ), .SUM(o[1281]) );
  FADDER \add_42/U1_1282  ( .CIN(sreg[1282]), .IN0(n2814), .IN1(
        \add_42/carry[1282] ), .COUT(\add_42/carry[1283] ), .SUM(o[1282]) );
  FADDER \add_42/U1_1283  ( .CIN(sreg[1283]), .IN0(n2813), .IN1(
        \add_42/carry[1283] ), .COUT(\add_42/carry[1284] ), .SUM(o[1283]) );
  FADDER \add_42/U1_1284  ( .CIN(sreg[1284]), .IN0(n2812), .IN1(
        \add_42/carry[1284] ), .COUT(\add_42/carry[1285] ), .SUM(o[1284]) );
  FADDER \add_42/U1_1285  ( .CIN(sreg[1285]), .IN0(n2811), .IN1(
        \add_42/carry[1285] ), .COUT(\add_42/carry[1286] ), .SUM(o[1285]) );
  FADDER \add_42/U1_1286  ( .CIN(sreg[1286]), .IN0(n2810), .IN1(
        \add_42/carry[1286] ), .COUT(\add_42/carry[1287] ), .SUM(o[1286]) );
  FADDER \add_42/U1_1287  ( .CIN(sreg[1287]), .IN0(n2809), .IN1(
        \add_42/carry[1287] ), .COUT(\add_42/carry[1288] ), .SUM(o[1287]) );
  FADDER \add_42/U1_1288  ( .CIN(sreg[1288]), .IN0(n2808), .IN1(
        \add_42/carry[1288] ), .COUT(\add_42/carry[1289] ), .SUM(o[1288]) );
  FADDER \add_42/U1_1289  ( .CIN(sreg[1289]), .IN0(n2807), .IN1(
        \add_42/carry[1289] ), .COUT(\add_42/carry[1290] ), .SUM(o[1289]) );
  FADDER \add_42/U1_1290  ( .CIN(sreg[1290]), .IN0(n2806), .IN1(
        \add_42/carry[1290] ), .COUT(\add_42/carry[1291] ), .SUM(o[1290]) );
  FADDER \add_42/U1_1291  ( .CIN(sreg[1291]), .IN0(n2805), .IN1(
        \add_42/carry[1291] ), .COUT(\add_42/carry[1292] ), .SUM(o[1291]) );
  FADDER \add_42/U1_1292  ( .CIN(sreg[1292]), .IN0(n2804), .IN1(
        \add_42/carry[1292] ), .COUT(\add_42/carry[1293] ), .SUM(o[1292]) );
  FADDER \add_42/U1_1293  ( .CIN(sreg[1293]), .IN0(n2803), .IN1(
        \add_42/carry[1293] ), .COUT(\add_42/carry[1294] ), .SUM(o[1293]) );
  FADDER \add_42/U1_1294  ( .CIN(sreg[1294]), .IN0(n2802), .IN1(
        \add_42/carry[1294] ), .COUT(\add_42/carry[1295] ), .SUM(o[1294]) );
  FADDER \add_42/U1_1295  ( .CIN(sreg[1295]), .IN0(n2801), .IN1(
        \add_42/carry[1295] ), .COUT(\add_42/carry[1296] ), .SUM(o[1295]) );
  FADDER \add_42/U1_1296  ( .CIN(sreg[1296]), .IN0(n2800), .IN1(
        \add_42/carry[1296] ), .COUT(\add_42/carry[1297] ), .SUM(o[1296]) );
  FADDER \add_42/U1_1297  ( .CIN(sreg[1297]), .IN0(n2799), .IN1(
        \add_42/carry[1297] ), .COUT(\add_42/carry[1298] ), .SUM(o[1297]) );
  FADDER \add_42/U1_1298  ( .CIN(sreg[1298]), .IN0(n2798), .IN1(
        \add_42/carry[1298] ), .COUT(\add_42/carry[1299] ), .SUM(o[1298]) );
  FADDER \add_42/U1_1299  ( .CIN(sreg[1299]), .IN0(n2797), .IN1(
        \add_42/carry[1299] ), .COUT(\add_42/carry[1300] ), .SUM(o[1299]) );
  FADDER \add_42/U1_1300  ( .CIN(sreg[1300]), .IN0(n2796), .IN1(
        \add_42/carry[1300] ), .COUT(\add_42/carry[1301] ), .SUM(o[1300]) );
  FADDER \add_42/U1_1301  ( .CIN(sreg[1301]), .IN0(n2795), .IN1(
        \add_42/carry[1301] ), .COUT(\add_42/carry[1302] ), .SUM(o[1301]) );
  FADDER \add_42/U1_1302  ( .CIN(sreg[1302]), .IN0(n2794), .IN1(
        \add_42/carry[1302] ), .COUT(\add_42/carry[1303] ), .SUM(o[1302]) );
  FADDER \add_42/U1_1303  ( .CIN(sreg[1303]), .IN0(n2793), .IN1(
        \add_42/carry[1303] ), .COUT(\add_42/carry[1304] ), .SUM(o[1303]) );
  FADDER \add_42/U1_1304  ( .CIN(sreg[1304]), .IN0(n2792), .IN1(
        \add_42/carry[1304] ), .COUT(\add_42/carry[1305] ), .SUM(o[1304]) );
  FADDER \add_42/U1_1305  ( .CIN(sreg[1305]), .IN0(n2791), .IN1(
        \add_42/carry[1305] ), .COUT(\add_42/carry[1306] ), .SUM(o[1305]) );
  FADDER \add_42/U1_1306  ( .CIN(sreg[1306]), .IN0(n2790), .IN1(
        \add_42/carry[1306] ), .COUT(\add_42/carry[1307] ), .SUM(o[1306]) );
  FADDER \add_42/U1_1307  ( .CIN(sreg[1307]), .IN0(n2789), .IN1(
        \add_42/carry[1307] ), .COUT(\add_42/carry[1308] ), .SUM(o[1307]) );
  FADDER \add_42/U1_1308  ( .CIN(sreg[1308]), .IN0(n2788), .IN1(
        \add_42/carry[1308] ), .COUT(\add_42/carry[1309] ), .SUM(o[1308]) );
  FADDER \add_42/U1_1309  ( .CIN(sreg[1309]), .IN0(n2787), .IN1(
        \add_42/carry[1309] ), .COUT(\add_42/carry[1310] ), .SUM(o[1309]) );
  FADDER \add_42/U1_1310  ( .CIN(sreg[1310]), .IN0(n2786), .IN1(
        \add_42/carry[1310] ), .COUT(\add_42/carry[1311] ), .SUM(o[1310]) );
  FADDER \add_42/U1_1311  ( .CIN(sreg[1311]), .IN0(n2785), .IN1(
        \add_42/carry[1311] ), .COUT(\add_42/carry[1312] ), .SUM(o[1311]) );
  FADDER \add_42/U1_1312  ( .CIN(sreg[1312]), .IN0(n2784), .IN1(
        \add_42/carry[1312] ), .COUT(\add_42/carry[1313] ), .SUM(o[1312]) );
  FADDER \add_42/U1_1313  ( .CIN(sreg[1313]), .IN0(n2783), .IN1(
        \add_42/carry[1313] ), .COUT(\add_42/carry[1314] ), .SUM(o[1313]) );
  FADDER \add_42/U1_1314  ( .CIN(sreg[1314]), .IN0(n2782), .IN1(
        \add_42/carry[1314] ), .COUT(\add_42/carry[1315] ), .SUM(o[1314]) );
  FADDER \add_42/U1_1315  ( .CIN(sreg[1315]), .IN0(n2781), .IN1(
        \add_42/carry[1315] ), .COUT(\add_42/carry[1316] ), .SUM(o[1315]) );
  FADDER \add_42/U1_1316  ( .CIN(sreg[1316]), .IN0(n2780), .IN1(
        \add_42/carry[1316] ), .COUT(\add_42/carry[1317] ), .SUM(o[1316]) );
  FADDER \add_42/U1_1317  ( .CIN(sreg[1317]), .IN0(n2779), .IN1(
        \add_42/carry[1317] ), .COUT(\add_42/carry[1318] ), .SUM(o[1317]) );
  FADDER \add_42/U1_1318  ( .CIN(sreg[1318]), .IN0(n2778), .IN1(
        \add_42/carry[1318] ), .COUT(\add_42/carry[1319] ), .SUM(o[1318]) );
  FADDER \add_42/U1_1319  ( .CIN(sreg[1319]), .IN0(n2777), .IN1(
        \add_42/carry[1319] ), .COUT(\add_42/carry[1320] ), .SUM(o[1319]) );
  FADDER \add_42/U1_1320  ( .CIN(sreg[1320]), .IN0(n2776), .IN1(
        \add_42/carry[1320] ), .COUT(\add_42/carry[1321] ), .SUM(o[1320]) );
  FADDER \add_42/U1_1321  ( .CIN(sreg[1321]), .IN0(n2775), .IN1(
        \add_42/carry[1321] ), .COUT(\add_42/carry[1322] ), .SUM(o[1321]) );
  FADDER \add_42/U1_1322  ( .CIN(sreg[1322]), .IN0(n2774), .IN1(
        \add_42/carry[1322] ), .COUT(\add_42/carry[1323] ), .SUM(o[1322]) );
  FADDER \add_42/U1_1323  ( .CIN(sreg[1323]), .IN0(n2773), .IN1(
        \add_42/carry[1323] ), .COUT(\add_42/carry[1324] ), .SUM(o[1323]) );
  FADDER \add_42/U1_1324  ( .CIN(sreg[1324]), .IN0(n2772), .IN1(
        \add_42/carry[1324] ), .COUT(\add_42/carry[1325] ), .SUM(o[1324]) );
  FADDER \add_42/U1_1325  ( .CIN(sreg[1325]), .IN0(n2771), .IN1(
        \add_42/carry[1325] ), .COUT(\add_42/carry[1326] ), .SUM(o[1325]) );
  FADDER \add_42/U1_1326  ( .CIN(sreg[1326]), .IN0(n2770), .IN1(
        \add_42/carry[1326] ), .COUT(\add_42/carry[1327] ), .SUM(o[1326]) );
  FADDER \add_42/U1_1327  ( .CIN(sreg[1327]), .IN0(n2769), .IN1(
        \add_42/carry[1327] ), .COUT(\add_42/carry[1328] ), .SUM(o[1327]) );
  FADDER \add_42/U1_1328  ( .CIN(sreg[1328]), .IN0(n2768), .IN1(
        \add_42/carry[1328] ), .COUT(\add_42/carry[1329] ), .SUM(o[1328]) );
  FADDER \add_42/U1_1329  ( .CIN(sreg[1329]), .IN0(n2767), .IN1(
        \add_42/carry[1329] ), .COUT(\add_42/carry[1330] ), .SUM(o[1329]) );
  FADDER \add_42/U1_1330  ( .CIN(sreg[1330]), .IN0(n2766), .IN1(
        \add_42/carry[1330] ), .COUT(\add_42/carry[1331] ), .SUM(o[1330]) );
  FADDER \add_42/U1_1331  ( .CIN(sreg[1331]), .IN0(n2765), .IN1(
        \add_42/carry[1331] ), .COUT(\add_42/carry[1332] ), .SUM(o[1331]) );
  FADDER \add_42/U1_1332  ( .CIN(sreg[1332]), .IN0(n2764), .IN1(
        \add_42/carry[1332] ), .COUT(\add_42/carry[1333] ), .SUM(o[1332]) );
  FADDER \add_42/U1_1333  ( .CIN(sreg[1333]), .IN0(n2763), .IN1(
        \add_42/carry[1333] ), .COUT(\add_42/carry[1334] ), .SUM(o[1333]) );
  FADDER \add_42/U1_1334  ( .CIN(sreg[1334]), .IN0(n2762), .IN1(
        \add_42/carry[1334] ), .COUT(\add_42/carry[1335] ), .SUM(o[1334]) );
  FADDER \add_42/U1_1335  ( .CIN(sreg[1335]), .IN0(n2761), .IN1(
        \add_42/carry[1335] ), .COUT(\add_42/carry[1336] ), .SUM(o[1335]) );
  FADDER \add_42/U1_1336  ( .CIN(sreg[1336]), .IN0(n2760), .IN1(
        \add_42/carry[1336] ), .COUT(\add_42/carry[1337] ), .SUM(o[1336]) );
  FADDER \add_42/U1_1337  ( .CIN(sreg[1337]), .IN0(n2759), .IN1(
        \add_42/carry[1337] ), .COUT(\add_42/carry[1338] ), .SUM(o[1337]) );
  FADDER \add_42/U1_1338  ( .CIN(sreg[1338]), .IN0(n2758), .IN1(
        \add_42/carry[1338] ), .COUT(\add_42/carry[1339] ), .SUM(o[1338]) );
  FADDER \add_42/U1_1339  ( .CIN(sreg[1339]), .IN0(n2757), .IN1(
        \add_42/carry[1339] ), .COUT(\add_42/carry[1340] ), .SUM(o[1339]) );
  FADDER \add_42/U1_1340  ( .CIN(sreg[1340]), .IN0(n2756), .IN1(
        \add_42/carry[1340] ), .COUT(\add_42/carry[1341] ), .SUM(o[1340]) );
  FADDER \add_42/U1_1341  ( .CIN(sreg[1341]), .IN0(n2755), .IN1(
        \add_42/carry[1341] ), .COUT(\add_42/carry[1342] ), .SUM(o[1341]) );
  FADDER \add_42/U1_1342  ( .CIN(sreg[1342]), .IN0(n2754), .IN1(
        \add_42/carry[1342] ), .COUT(\add_42/carry[1343] ), .SUM(o[1342]) );
  FADDER \add_42/U1_1343  ( .CIN(sreg[1343]), .IN0(n2753), .IN1(
        \add_42/carry[1343] ), .COUT(\add_42/carry[1344] ), .SUM(o[1343]) );
  FADDER \add_42/U1_1344  ( .CIN(sreg[1344]), .IN0(n2752), .IN1(
        \add_42/carry[1344] ), .COUT(\add_42/carry[1345] ), .SUM(o[1344]) );
  FADDER \add_42/U1_1345  ( .CIN(sreg[1345]), .IN0(n2751), .IN1(
        \add_42/carry[1345] ), .COUT(\add_42/carry[1346] ), .SUM(o[1345]) );
  FADDER \add_42/U1_1346  ( .CIN(sreg[1346]), .IN0(n2750), .IN1(
        \add_42/carry[1346] ), .COUT(\add_42/carry[1347] ), .SUM(o[1346]) );
  FADDER \add_42/U1_1347  ( .CIN(sreg[1347]), .IN0(n2749), .IN1(
        \add_42/carry[1347] ), .COUT(\add_42/carry[1348] ), .SUM(o[1347]) );
  FADDER \add_42/U1_1348  ( .CIN(sreg[1348]), .IN0(n2748), .IN1(
        \add_42/carry[1348] ), .COUT(\add_42/carry[1349] ), .SUM(o[1348]) );
  FADDER \add_42/U1_1349  ( .CIN(sreg[1349]), .IN0(n2747), .IN1(
        \add_42/carry[1349] ), .COUT(\add_42/carry[1350] ), .SUM(o[1349]) );
  FADDER \add_42/U1_1350  ( .CIN(sreg[1350]), .IN0(n2746), .IN1(
        \add_42/carry[1350] ), .COUT(\add_42/carry[1351] ), .SUM(o[1350]) );
  FADDER \add_42/U1_1351  ( .CIN(sreg[1351]), .IN0(n2745), .IN1(
        \add_42/carry[1351] ), .COUT(\add_42/carry[1352] ), .SUM(o[1351]) );
  FADDER \add_42/U1_1352  ( .CIN(sreg[1352]), .IN0(n2744), .IN1(
        \add_42/carry[1352] ), .COUT(\add_42/carry[1353] ), .SUM(o[1352]) );
  FADDER \add_42/U1_1353  ( .CIN(sreg[1353]), .IN0(n2743), .IN1(
        \add_42/carry[1353] ), .COUT(\add_42/carry[1354] ), .SUM(o[1353]) );
  FADDER \add_42/U1_1354  ( .CIN(sreg[1354]), .IN0(n2742), .IN1(
        \add_42/carry[1354] ), .COUT(\add_42/carry[1355] ), .SUM(o[1354]) );
  FADDER \add_42/U1_1355  ( .CIN(sreg[1355]), .IN0(n2741), .IN1(
        \add_42/carry[1355] ), .COUT(\add_42/carry[1356] ), .SUM(o[1355]) );
  FADDER \add_42/U1_1356  ( .CIN(sreg[1356]), .IN0(n2740), .IN1(
        \add_42/carry[1356] ), .COUT(\add_42/carry[1357] ), .SUM(o[1356]) );
  FADDER \add_42/U1_1357  ( .CIN(sreg[1357]), .IN0(n2739), .IN1(
        \add_42/carry[1357] ), .COUT(\add_42/carry[1358] ), .SUM(o[1357]) );
  FADDER \add_42/U1_1358  ( .CIN(sreg[1358]), .IN0(n2738), .IN1(
        \add_42/carry[1358] ), .COUT(\add_42/carry[1359] ), .SUM(o[1358]) );
  FADDER \add_42/U1_1359  ( .CIN(sreg[1359]), .IN0(n2737), .IN1(
        \add_42/carry[1359] ), .COUT(\add_42/carry[1360] ), .SUM(o[1359]) );
  FADDER \add_42/U1_1360  ( .CIN(sreg[1360]), .IN0(n2736), .IN1(
        \add_42/carry[1360] ), .COUT(\add_42/carry[1361] ), .SUM(o[1360]) );
  FADDER \add_42/U1_1361  ( .CIN(sreg[1361]), .IN0(n2735), .IN1(
        \add_42/carry[1361] ), .COUT(\add_42/carry[1362] ), .SUM(o[1361]) );
  FADDER \add_42/U1_1362  ( .CIN(sreg[1362]), .IN0(n2734), .IN1(
        \add_42/carry[1362] ), .COUT(\add_42/carry[1363] ), .SUM(o[1362]) );
  FADDER \add_42/U1_1363  ( .CIN(sreg[1363]), .IN0(n2733), .IN1(
        \add_42/carry[1363] ), .COUT(\add_42/carry[1364] ), .SUM(o[1363]) );
  FADDER \add_42/U1_1364  ( .CIN(sreg[1364]), .IN0(n2732), .IN1(
        \add_42/carry[1364] ), .COUT(\add_42/carry[1365] ), .SUM(o[1364]) );
  FADDER \add_42/U1_1365  ( .CIN(sreg[1365]), .IN0(n2731), .IN1(
        \add_42/carry[1365] ), .COUT(\add_42/carry[1366] ), .SUM(o[1365]) );
  FADDER \add_42/U1_1366  ( .CIN(sreg[1366]), .IN0(n2730), .IN1(
        \add_42/carry[1366] ), .COUT(\add_42/carry[1367] ), .SUM(o[1366]) );
  FADDER \add_42/U1_1367  ( .CIN(sreg[1367]), .IN0(n2729), .IN1(
        \add_42/carry[1367] ), .COUT(\add_42/carry[1368] ), .SUM(o[1367]) );
  FADDER \add_42/U1_1368  ( .CIN(sreg[1368]), .IN0(n2728), .IN1(
        \add_42/carry[1368] ), .COUT(\add_42/carry[1369] ), .SUM(o[1368]) );
  FADDER \add_42/U1_1369  ( .CIN(sreg[1369]), .IN0(n2727), .IN1(
        \add_42/carry[1369] ), .COUT(\add_42/carry[1370] ), .SUM(o[1369]) );
  FADDER \add_42/U1_1370  ( .CIN(sreg[1370]), .IN0(n2726), .IN1(
        \add_42/carry[1370] ), .COUT(\add_42/carry[1371] ), .SUM(o[1370]) );
  FADDER \add_42/U1_1371  ( .CIN(sreg[1371]), .IN0(n2725), .IN1(
        \add_42/carry[1371] ), .COUT(\add_42/carry[1372] ), .SUM(o[1371]) );
  FADDER \add_42/U1_1372  ( .CIN(sreg[1372]), .IN0(n2724), .IN1(
        \add_42/carry[1372] ), .COUT(\add_42/carry[1373] ), .SUM(o[1372]) );
  FADDER \add_42/U1_1373  ( .CIN(sreg[1373]), .IN0(n2723), .IN1(
        \add_42/carry[1373] ), .COUT(\add_42/carry[1374] ), .SUM(o[1373]) );
  FADDER \add_42/U1_1374  ( .CIN(sreg[1374]), .IN0(n2722), .IN1(
        \add_42/carry[1374] ), .COUT(\add_42/carry[1375] ), .SUM(o[1374]) );
  FADDER \add_42/U1_1375  ( .CIN(sreg[1375]), .IN0(n2721), .IN1(
        \add_42/carry[1375] ), .COUT(\add_42/carry[1376] ), .SUM(o[1375]) );
  FADDER \add_42/U1_1376  ( .CIN(sreg[1376]), .IN0(n2720), .IN1(
        \add_42/carry[1376] ), .COUT(\add_42/carry[1377] ), .SUM(o[1376]) );
  FADDER \add_42/U1_1377  ( .CIN(sreg[1377]), .IN0(n2719), .IN1(
        \add_42/carry[1377] ), .COUT(\add_42/carry[1378] ), .SUM(o[1377]) );
  FADDER \add_42/U1_1378  ( .CIN(sreg[1378]), .IN0(n2718), .IN1(
        \add_42/carry[1378] ), .COUT(\add_42/carry[1379] ), .SUM(o[1378]) );
  FADDER \add_42/U1_1379  ( .CIN(sreg[1379]), .IN0(n2717), .IN1(
        \add_42/carry[1379] ), .COUT(\add_42/carry[1380] ), .SUM(o[1379]) );
  FADDER \add_42/U1_1380  ( .CIN(sreg[1380]), .IN0(n2716), .IN1(
        \add_42/carry[1380] ), .COUT(\add_42/carry[1381] ), .SUM(o[1380]) );
  FADDER \add_42/U1_1381  ( .CIN(sreg[1381]), .IN0(n2715), .IN1(
        \add_42/carry[1381] ), .COUT(\add_42/carry[1382] ), .SUM(o[1381]) );
  FADDER \add_42/U1_1382  ( .CIN(sreg[1382]), .IN0(n2714), .IN1(
        \add_42/carry[1382] ), .COUT(\add_42/carry[1383] ), .SUM(o[1382]) );
  FADDER \add_42/U1_1383  ( .CIN(sreg[1383]), .IN0(n2713), .IN1(
        \add_42/carry[1383] ), .COUT(\add_42/carry[1384] ), .SUM(o[1383]) );
  FADDER \add_42/U1_1384  ( .CIN(sreg[1384]), .IN0(n2712), .IN1(
        \add_42/carry[1384] ), .COUT(\add_42/carry[1385] ), .SUM(o[1384]) );
  FADDER \add_42/U1_1385  ( .CIN(sreg[1385]), .IN0(n2711), .IN1(
        \add_42/carry[1385] ), .COUT(\add_42/carry[1386] ), .SUM(o[1385]) );
  FADDER \add_42/U1_1386  ( .CIN(sreg[1386]), .IN0(n2710), .IN1(
        \add_42/carry[1386] ), .COUT(\add_42/carry[1387] ), .SUM(o[1386]) );
  FADDER \add_42/U1_1387  ( .CIN(sreg[1387]), .IN0(n2709), .IN1(
        \add_42/carry[1387] ), .COUT(\add_42/carry[1388] ), .SUM(o[1387]) );
  FADDER \add_42/U1_1388  ( .CIN(sreg[1388]), .IN0(n2708), .IN1(
        \add_42/carry[1388] ), .COUT(\add_42/carry[1389] ), .SUM(o[1388]) );
  FADDER \add_42/U1_1389  ( .CIN(sreg[1389]), .IN0(n2707), .IN1(
        \add_42/carry[1389] ), .COUT(\add_42/carry[1390] ), .SUM(o[1389]) );
  FADDER \add_42/U1_1390  ( .CIN(sreg[1390]), .IN0(n2706), .IN1(
        \add_42/carry[1390] ), .COUT(\add_42/carry[1391] ), .SUM(o[1390]) );
  FADDER \add_42/U1_1391  ( .CIN(sreg[1391]), .IN0(n2705), .IN1(
        \add_42/carry[1391] ), .COUT(\add_42/carry[1392] ), .SUM(o[1391]) );
  FADDER \add_42/U1_1392  ( .CIN(sreg[1392]), .IN0(n2704), .IN1(
        \add_42/carry[1392] ), .COUT(\add_42/carry[1393] ), .SUM(o[1392]) );
  FADDER \add_42/U1_1393  ( .CIN(sreg[1393]), .IN0(n2703), .IN1(
        \add_42/carry[1393] ), .COUT(\add_42/carry[1394] ), .SUM(o[1393]) );
  FADDER \add_42/U1_1394  ( .CIN(sreg[1394]), .IN0(n2702), .IN1(
        \add_42/carry[1394] ), .COUT(\add_42/carry[1395] ), .SUM(o[1394]) );
  FADDER \add_42/U1_1395  ( .CIN(sreg[1395]), .IN0(n2701), .IN1(
        \add_42/carry[1395] ), .COUT(\add_42/carry[1396] ), .SUM(o[1395]) );
  FADDER \add_42/U1_1396  ( .CIN(sreg[1396]), .IN0(n2700), .IN1(
        \add_42/carry[1396] ), .COUT(\add_42/carry[1397] ), .SUM(o[1396]) );
  FADDER \add_42/U1_1397  ( .CIN(sreg[1397]), .IN0(n2699), .IN1(
        \add_42/carry[1397] ), .COUT(\add_42/carry[1398] ), .SUM(o[1397]) );
  FADDER \add_42/U1_1398  ( .CIN(sreg[1398]), .IN0(n2698), .IN1(
        \add_42/carry[1398] ), .COUT(\add_42/carry[1399] ), .SUM(o[1398]) );
  FADDER \add_42/U1_1399  ( .CIN(sreg[1399]), .IN0(n2697), .IN1(
        \add_42/carry[1399] ), .COUT(\add_42/carry[1400] ), .SUM(o[1399]) );
  FADDER \add_42/U1_1400  ( .CIN(sreg[1400]), .IN0(n2696), .IN1(
        \add_42/carry[1400] ), .COUT(\add_42/carry[1401] ), .SUM(o[1400]) );
  FADDER \add_42/U1_1401  ( .CIN(sreg[1401]), .IN0(n2695), .IN1(
        \add_42/carry[1401] ), .COUT(\add_42/carry[1402] ), .SUM(o[1401]) );
  FADDER \add_42/U1_1402  ( .CIN(sreg[1402]), .IN0(n2694), .IN1(
        \add_42/carry[1402] ), .COUT(\add_42/carry[1403] ), .SUM(o[1402]) );
  FADDER \add_42/U1_1403  ( .CIN(sreg[1403]), .IN0(n2693), .IN1(
        \add_42/carry[1403] ), .COUT(\add_42/carry[1404] ), .SUM(o[1403]) );
  FADDER \add_42/U1_1404  ( .CIN(sreg[1404]), .IN0(n2692), .IN1(
        \add_42/carry[1404] ), .COUT(\add_42/carry[1405] ), .SUM(o[1404]) );
  FADDER \add_42/U1_1405  ( .CIN(sreg[1405]), .IN0(n2691), .IN1(
        \add_42/carry[1405] ), .COUT(\add_42/carry[1406] ), .SUM(o[1405]) );
  FADDER \add_42/U1_1406  ( .CIN(sreg[1406]), .IN0(n2690), .IN1(
        \add_42/carry[1406] ), .COUT(\add_42/carry[1407] ), .SUM(o[1406]) );
  FADDER \add_42/U1_1407  ( .CIN(sreg[1407]), .IN0(n2689), .IN1(
        \add_42/carry[1407] ), .COUT(\add_42/carry[1408] ), .SUM(o[1407]) );
  FADDER \add_42/U1_1408  ( .CIN(sreg[1408]), .IN0(n2688), .IN1(
        \add_42/carry[1408] ), .COUT(\add_42/carry[1409] ), .SUM(o[1408]) );
  FADDER \add_42/U1_1409  ( .CIN(sreg[1409]), .IN0(n2687), .IN1(
        \add_42/carry[1409] ), .COUT(\add_42/carry[1410] ), .SUM(o[1409]) );
  FADDER \add_42/U1_1410  ( .CIN(sreg[1410]), .IN0(n2686), .IN1(
        \add_42/carry[1410] ), .COUT(\add_42/carry[1411] ), .SUM(o[1410]) );
  FADDER \add_42/U1_1411  ( .CIN(sreg[1411]), .IN0(n2685), .IN1(
        \add_42/carry[1411] ), .COUT(\add_42/carry[1412] ), .SUM(o[1411]) );
  FADDER \add_42/U1_1412  ( .CIN(sreg[1412]), .IN0(n2684), .IN1(
        \add_42/carry[1412] ), .COUT(\add_42/carry[1413] ), .SUM(o[1412]) );
  FADDER \add_42/U1_1413  ( .CIN(sreg[1413]), .IN0(n2683), .IN1(
        \add_42/carry[1413] ), .COUT(\add_42/carry[1414] ), .SUM(o[1413]) );
  FADDER \add_42/U1_1414  ( .CIN(sreg[1414]), .IN0(n2682), .IN1(
        \add_42/carry[1414] ), .COUT(\add_42/carry[1415] ), .SUM(o[1414]) );
  FADDER \add_42/U1_1415  ( .CIN(sreg[1415]), .IN0(n2681), .IN1(
        \add_42/carry[1415] ), .COUT(\add_42/carry[1416] ), .SUM(o[1415]) );
  FADDER \add_42/U1_1416  ( .CIN(sreg[1416]), .IN0(n2680), .IN1(
        \add_42/carry[1416] ), .COUT(\add_42/carry[1417] ), .SUM(o[1416]) );
  FADDER \add_42/U1_1417  ( .CIN(sreg[1417]), .IN0(n2679), .IN1(
        \add_42/carry[1417] ), .COUT(\add_42/carry[1418] ), .SUM(o[1417]) );
  FADDER \add_42/U1_1418  ( .CIN(sreg[1418]), .IN0(n2678), .IN1(
        \add_42/carry[1418] ), .COUT(\add_42/carry[1419] ), .SUM(o[1418]) );
  FADDER \add_42/U1_1419  ( .CIN(sreg[1419]), .IN0(n2677), .IN1(
        \add_42/carry[1419] ), .COUT(\add_42/carry[1420] ), .SUM(o[1419]) );
  FADDER \add_42/U1_1420  ( .CIN(sreg[1420]), .IN0(n2676), .IN1(
        \add_42/carry[1420] ), .COUT(\add_42/carry[1421] ), .SUM(o[1420]) );
  FADDER \add_42/U1_1421  ( .CIN(sreg[1421]), .IN0(n2675), .IN1(
        \add_42/carry[1421] ), .COUT(\add_42/carry[1422] ), .SUM(o[1421]) );
  FADDER \add_42/U1_1422  ( .CIN(sreg[1422]), .IN0(n2674), .IN1(
        \add_42/carry[1422] ), .COUT(\add_42/carry[1423] ), .SUM(o[1422]) );
  FADDER \add_42/U1_1423  ( .CIN(sreg[1423]), .IN0(n2673), .IN1(
        \add_42/carry[1423] ), .COUT(\add_42/carry[1424] ), .SUM(o[1423]) );
  FADDER \add_42/U1_1424  ( .CIN(sreg[1424]), .IN0(n2672), .IN1(
        \add_42/carry[1424] ), .COUT(\add_42/carry[1425] ), .SUM(o[1424]) );
  FADDER \add_42/U1_1425  ( .CIN(sreg[1425]), .IN0(n2671), .IN1(
        \add_42/carry[1425] ), .COUT(\add_42/carry[1426] ), .SUM(o[1425]) );
  FADDER \add_42/U1_1426  ( .CIN(sreg[1426]), .IN0(n2670), .IN1(
        \add_42/carry[1426] ), .COUT(\add_42/carry[1427] ), .SUM(o[1426]) );
  FADDER \add_42/U1_1427  ( .CIN(sreg[1427]), .IN0(n2669), .IN1(
        \add_42/carry[1427] ), .COUT(\add_42/carry[1428] ), .SUM(o[1427]) );
  FADDER \add_42/U1_1428  ( .CIN(sreg[1428]), .IN0(n2668), .IN1(
        \add_42/carry[1428] ), .COUT(\add_42/carry[1429] ), .SUM(o[1428]) );
  FADDER \add_42/U1_1429  ( .CIN(sreg[1429]), .IN0(n2667), .IN1(
        \add_42/carry[1429] ), .COUT(\add_42/carry[1430] ), .SUM(o[1429]) );
  FADDER \add_42/U1_1430  ( .CIN(sreg[1430]), .IN0(n2666), .IN1(
        \add_42/carry[1430] ), .COUT(\add_42/carry[1431] ), .SUM(o[1430]) );
  FADDER \add_42/U1_1431  ( .CIN(sreg[1431]), .IN0(n2665), .IN1(
        \add_42/carry[1431] ), .COUT(\add_42/carry[1432] ), .SUM(o[1431]) );
  FADDER \add_42/U1_1432  ( .CIN(sreg[1432]), .IN0(n2664), .IN1(
        \add_42/carry[1432] ), .COUT(\add_42/carry[1433] ), .SUM(o[1432]) );
  FADDER \add_42/U1_1433  ( .CIN(sreg[1433]), .IN0(n2663), .IN1(
        \add_42/carry[1433] ), .COUT(\add_42/carry[1434] ), .SUM(o[1433]) );
  FADDER \add_42/U1_1434  ( .CIN(sreg[1434]), .IN0(n2662), .IN1(
        \add_42/carry[1434] ), .COUT(\add_42/carry[1435] ), .SUM(o[1434]) );
  FADDER \add_42/U1_1435  ( .CIN(sreg[1435]), .IN0(n2661), .IN1(
        \add_42/carry[1435] ), .COUT(\add_42/carry[1436] ), .SUM(o[1435]) );
  FADDER \add_42/U1_1436  ( .CIN(sreg[1436]), .IN0(n2660), .IN1(
        \add_42/carry[1436] ), .COUT(\add_42/carry[1437] ), .SUM(o[1436]) );
  FADDER \add_42/U1_1437  ( .CIN(sreg[1437]), .IN0(n2659), .IN1(
        \add_42/carry[1437] ), .COUT(\add_42/carry[1438] ), .SUM(o[1437]) );
  FADDER \add_42/U1_1438  ( .CIN(sreg[1438]), .IN0(n2658), .IN1(
        \add_42/carry[1438] ), .COUT(\add_42/carry[1439] ), .SUM(o[1438]) );
  FADDER \add_42/U1_1439  ( .CIN(sreg[1439]), .IN0(n2657), .IN1(
        \add_42/carry[1439] ), .COUT(\add_42/carry[1440] ), .SUM(o[1439]) );
  FADDER \add_42/U1_1440  ( .CIN(sreg[1440]), .IN0(n2656), .IN1(
        \add_42/carry[1440] ), .COUT(\add_42/carry[1441] ), .SUM(o[1440]) );
  FADDER \add_42/U1_1441  ( .CIN(sreg[1441]), .IN0(n2655), .IN1(
        \add_42/carry[1441] ), .COUT(\add_42/carry[1442] ), .SUM(o[1441]) );
  FADDER \add_42/U1_1442  ( .CIN(sreg[1442]), .IN0(n2654), .IN1(
        \add_42/carry[1442] ), .COUT(\add_42/carry[1443] ), .SUM(o[1442]) );
  FADDER \add_42/U1_1443  ( .CIN(sreg[1443]), .IN0(n2653), .IN1(
        \add_42/carry[1443] ), .COUT(\add_42/carry[1444] ), .SUM(o[1443]) );
  FADDER \add_42/U1_1444  ( .CIN(sreg[1444]), .IN0(n2652), .IN1(
        \add_42/carry[1444] ), .COUT(\add_42/carry[1445] ), .SUM(o[1444]) );
  FADDER \add_42/U1_1445  ( .CIN(sreg[1445]), .IN0(n2651), .IN1(
        \add_42/carry[1445] ), .COUT(\add_42/carry[1446] ), .SUM(o[1445]) );
  FADDER \add_42/U1_1446  ( .CIN(sreg[1446]), .IN0(n2650), .IN1(
        \add_42/carry[1446] ), .COUT(\add_42/carry[1447] ), .SUM(o[1446]) );
  FADDER \add_42/U1_1447  ( .CIN(sreg[1447]), .IN0(n2649), .IN1(
        \add_42/carry[1447] ), .COUT(\add_42/carry[1448] ), .SUM(o[1447]) );
  FADDER \add_42/U1_1448  ( .CIN(sreg[1448]), .IN0(n2648), .IN1(
        \add_42/carry[1448] ), .COUT(\add_42/carry[1449] ), .SUM(o[1448]) );
  FADDER \add_42/U1_1449  ( .CIN(sreg[1449]), .IN0(n2647), .IN1(
        \add_42/carry[1449] ), .COUT(\add_42/carry[1450] ), .SUM(o[1449]) );
  FADDER \add_42/U1_1450  ( .CIN(sreg[1450]), .IN0(n2646), .IN1(
        \add_42/carry[1450] ), .COUT(\add_42/carry[1451] ), .SUM(o[1450]) );
  FADDER \add_42/U1_1451  ( .CIN(sreg[1451]), .IN0(n2645), .IN1(
        \add_42/carry[1451] ), .COUT(\add_42/carry[1452] ), .SUM(o[1451]) );
  FADDER \add_42/U1_1452  ( .CIN(sreg[1452]), .IN0(n2644), .IN1(
        \add_42/carry[1452] ), .COUT(\add_42/carry[1453] ), .SUM(o[1452]) );
  FADDER \add_42/U1_1453  ( .CIN(sreg[1453]), .IN0(n2643), .IN1(
        \add_42/carry[1453] ), .COUT(\add_42/carry[1454] ), .SUM(o[1453]) );
  FADDER \add_42/U1_1454  ( .CIN(sreg[1454]), .IN0(n2642), .IN1(
        \add_42/carry[1454] ), .COUT(\add_42/carry[1455] ), .SUM(o[1454]) );
  FADDER \add_42/U1_1455  ( .CIN(sreg[1455]), .IN0(n2641), .IN1(
        \add_42/carry[1455] ), .COUT(\add_42/carry[1456] ), .SUM(o[1455]) );
  FADDER \add_42/U1_1456  ( .CIN(sreg[1456]), .IN0(n2640), .IN1(
        \add_42/carry[1456] ), .COUT(\add_42/carry[1457] ), .SUM(o[1456]) );
  FADDER \add_42/U1_1457  ( .CIN(sreg[1457]), .IN0(n2639), .IN1(
        \add_42/carry[1457] ), .COUT(\add_42/carry[1458] ), .SUM(o[1457]) );
  FADDER \add_42/U1_1458  ( .CIN(sreg[1458]), .IN0(n2638), .IN1(
        \add_42/carry[1458] ), .COUT(\add_42/carry[1459] ), .SUM(o[1458]) );
  FADDER \add_42/U1_1459  ( .CIN(sreg[1459]), .IN0(n2637), .IN1(
        \add_42/carry[1459] ), .COUT(\add_42/carry[1460] ), .SUM(o[1459]) );
  FADDER \add_42/U1_1460  ( .CIN(sreg[1460]), .IN0(n2636), .IN1(
        \add_42/carry[1460] ), .COUT(\add_42/carry[1461] ), .SUM(o[1460]) );
  FADDER \add_42/U1_1461  ( .CIN(sreg[1461]), .IN0(n2635), .IN1(
        \add_42/carry[1461] ), .COUT(\add_42/carry[1462] ), .SUM(o[1461]) );
  FADDER \add_42/U1_1462  ( .CIN(sreg[1462]), .IN0(n2634), .IN1(
        \add_42/carry[1462] ), .COUT(\add_42/carry[1463] ), .SUM(o[1462]) );
  FADDER \add_42/U1_1463  ( .CIN(sreg[1463]), .IN0(n2633), .IN1(
        \add_42/carry[1463] ), .COUT(\add_42/carry[1464] ), .SUM(o[1463]) );
  FADDER \add_42/U1_1464  ( .CIN(sreg[1464]), .IN0(n2632), .IN1(
        \add_42/carry[1464] ), .COUT(\add_42/carry[1465] ), .SUM(o[1464]) );
  FADDER \add_42/U1_1465  ( .CIN(sreg[1465]), .IN0(n2631), .IN1(
        \add_42/carry[1465] ), .COUT(\add_42/carry[1466] ), .SUM(o[1465]) );
  FADDER \add_42/U1_1466  ( .CIN(sreg[1466]), .IN0(n2630), .IN1(
        \add_42/carry[1466] ), .COUT(\add_42/carry[1467] ), .SUM(o[1466]) );
  FADDER \add_42/U1_1467  ( .CIN(sreg[1467]), .IN0(n2629), .IN1(
        \add_42/carry[1467] ), .COUT(\add_42/carry[1468] ), .SUM(o[1467]) );
  FADDER \add_42/U1_1468  ( .CIN(sreg[1468]), .IN0(n2628), .IN1(
        \add_42/carry[1468] ), .COUT(\add_42/carry[1469] ), .SUM(o[1468]) );
  FADDER \add_42/U1_1469  ( .CIN(sreg[1469]), .IN0(n2627), .IN1(
        \add_42/carry[1469] ), .COUT(\add_42/carry[1470] ), .SUM(o[1469]) );
  FADDER \add_42/U1_1470  ( .CIN(sreg[1470]), .IN0(n2626), .IN1(
        \add_42/carry[1470] ), .COUT(\add_42/carry[1471] ), .SUM(o[1470]) );
  FADDER \add_42/U1_1471  ( .CIN(sreg[1471]), .IN0(n2625), .IN1(
        \add_42/carry[1471] ), .COUT(\add_42/carry[1472] ), .SUM(o[1471]) );
  FADDER \add_42/U1_1472  ( .CIN(sreg[1472]), .IN0(n2624), .IN1(
        \add_42/carry[1472] ), .COUT(\add_42/carry[1473] ), .SUM(o[1472]) );
  FADDER \add_42/U1_1473  ( .CIN(sreg[1473]), .IN0(n2623), .IN1(
        \add_42/carry[1473] ), .COUT(\add_42/carry[1474] ), .SUM(o[1473]) );
  FADDER \add_42/U1_1474  ( .CIN(sreg[1474]), .IN0(n2622), .IN1(
        \add_42/carry[1474] ), .COUT(\add_42/carry[1475] ), .SUM(o[1474]) );
  FADDER \add_42/U1_1475  ( .CIN(sreg[1475]), .IN0(n2621), .IN1(
        \add_42/carry[1475] ), .COUT(\add_42/carry[1476] ), .SUM(o[1475]) );
  FADDER \add_42/U1_1476  ( .CIN(sreg[1476]), .IN0(n2620), .IN1(
        \add_42/carry[1476] ), .COUT(\add_42/carry[1477] ), .SUM(o[1476]) );
  FADDER \add_42/U1_1477  ( .CIN(sreg[1477]), .IN0(n2619), .IN1(
        \add_42/carry[1477] ), .COUT(\add_42/carry[1478] ), .SUM(o[1477]) );
  FADDER \add_42/U1_1478  ( .CIN(sreg[1478]), .IN0(n2618), .IN1(
        \add_42/carry[1478] ), .COUT(\add_42/carry[1479] ), .SUM(o[1478]) );
  FADDER \add_42/U1_1479  ( .CIN(sreg[1479]), .IN0(n2617), .IN1(
        \add_42/carry[1479] ), .COUT(\add_42/carry[1480] ), .SUM(o[1479]) );
  FADDER \add_42/U1_1480  ( .CIN(sreg[1480]), .IN0(n2616), .IN1(
        \add_42/carry[1480] ), .COUT(\add_42/carry[1481] ), .SUM(o[1480]) );
  FADDER \add_42/U1_1481  ( .CIN(sreg[1481]), .IN0(n2615), .IN1(
        \add_42/carry[1481] ), .COUT(\add_42/carry[1482] ), .SUM(o[1481]) );
  FADDER \add_42/U1_1482  ( .CIN(sreg[1482]), .IN0(n2614), .IN1(
        \add_42/carry[1482] ), .COUT(\add_42/carry[1483] ), .SUM(o[1482]) );
  FADDER \add_42/U1_1483  ( .CIN(sreg[1483]), .IN0(n2613), .IN1(
        \add_42/carry[1483] ), .COUT(\add_42/carry[1484] ), .SUM(o[1483]) );
  FADDER \add_42/U1_1484  ( .CIN(sreg[1484]), .IN0(n2612), .IN1(
        \add_42/carry[1484] ), .COUT(\add_42/carry[1485] ), .SUM(o[1484]) );
  FADDER \add_42/U1_1485  ( .CIN(sreg[1485]), .IN0(n2611), .IN1(
        \add_42/carry[1485] ), .COUT(\add_42/carry[1486] ), .SUM(o[1485]) );
  FADDER \add_42/U1_1486  ( .CIN(sreg[1486]), .IN0(n2610), .IN1(
        \add_42/carry[1486] ), .COUT(\add_42/carry[1487] ), .SUM(o[1486]) );
  FADDER \add_42/U1_1487  ( .CIN(sreg[1487]), .IN0(n2609), .IN1(
        \add_42/carry[1487] ), .COUT(\add_42/carry[1488] ), .SUM(o[1487]) );
  FADDER \add_42/U1_1488  ( .CIN(sreg[1488]), .IN0(n2608), .IN1(
        \add_42/carry[1488] ), .COUT(\add_42/carry[1489] ), .SUM(o[1488]) );
  FADDER \add_42/U1_1489  ( .CIN(sreg[1489]), .IN0(n2607), .IN1(
        \add_42/carry[1489] ), .COUT(\add_42/carry[1490] ), .SUM(o[1489]) );
  FADDER \add_42/U1_1490  ( .CIN(sreg[1490]), .IN0(n2606), .IN1(
        \add_42/carry[1490] ), .COUT(\add_42/carry[1491] ), .SUM(o[1490]) );
  FADDER \add_42/U1_1491  ( .CIN(sreg[1491]), .IN0(n2605), .IN1(
        \add_42/carry[1491] ), .COUT(\add_42/carry[1492] ), .SUM(o[1491]) );
  FADDER \add_42/U1_1492  ( .CIN(sreg[1492]), .IN0(n2604), .IN1(
        \add_42/carry[1492] ), .COUT(\add_42/carry[1493] ), .SUM(o[1492]) );
  FADDER \add_42/U1_1493  ( .CIN(sreg[1493]), .IN0(n2603), .IN1(
        \add_42/carry[1493] ), .COUT(\add_42/carry[1494] ), .SUM(o[1493]) );
  FADDER \add_42/U1_1494  ( .CIN(sreg[1494]), .IN0(n2602), .IN1(
        \add_42/carry[1494] ), .COUT(\add_42/carry[1495] ), .SUM(o[1494]) );
  FADDER \add_42/U1_1495  ( .CIN(sreg[1495]), .IN0(n2601), .IN1(
        \add_42/carry[1495] ), .COUT(\add_42/carry[1496] ), .SUM(o[1495]) );
  FADDER \add_42/U1_1496  ( .CIN(sreg[1496]), .IN0(n2600), .IN1(
        \add_42/carry[1496] ), .COUT(\add_42/carry[1497] ), .SUM(o[1496]) );
  FADDER \add_42/U1_1497  ( .CIN(sreg[1497]), .IN0(n2599), .IN1(
        \add_42/carry[1497] ), .COUT(\add_42/carry[1498] ), .SUM(o[1497]) );
  FADDER \add_42/U1_1498  ( .CIN(sreg[1498]), .IN0(n2598), .IN1(
        \add_42/carry[1498] ), .COUT(\add_42/carry[1499] ), .SUM(o[1498]) );
  FADDER \add_42/U1_1499  ( .CIN(sreg[1499]), .IN0(n2597), .IN1(
        \add_42/carry[1499] ), .COUT(\add_42/carry[1500] ), .SUM(o[1499]) );
  FADDER \add_42/U1_1500  ( .CIN(sreg[1500]), .IN0(n2596), .IN1(
        \add_42/carry[1500] ), .COUT(\add_42/carry[1501] ), .SUM(o[1500]) );
  FADDER \add_42/U1_1501  ( .CIN(sreg[1501]), .IN0(n2595), .IN1(
        \add_42/carry[1501] ), .COUT(\add_42/carry[1502] ), .SUM(o[1501]) );
  FADDER \add_42/U1_1502  ( .CIN(sreg[1502]), .IN0(n2594), .IN1(
        \add_42/carry[1502] ), .COUT(\add_42/carry[1503] ), .SUM(o[1502]) );
  FADDER \add_42/U1_1503  ( .CIN(sreg[1503]), .IN0(n2593), .IN1(
        \add_42/carry[1503] ), .COUT(\add_42/carry[1504] ), .SUM(o[1503]) );
  FADDER \add_42/U1_1504  ( .CIN(sreg[1504]), .IN0(n2592), .IN1(
        \add_42/carry[1504] ), .COUT(\add_42/carry[1505] ), .SUM(o[1504]) );
  FADDER \add_42/U1_1505  ( .CIN(sreg[1505]), .IN0(n2591), .IN1(
        \add_42/carry[1505] ), .COUT(\add_42/carry[1506] ), .SUM(o[1505]) );
  FADDER \add_42/U1_1506  ( .CIN(sreg[1506]), .IN0(n2590), .IN1(
        \add_42/carry[1506] ), .COUT(\add_42/carry[1507] ), .SUM(o[1506]) );
  FADDER \add_42/U1_1507  ( .CIN(sreg[1507]), .IN0(n2589), .IN1(
        \add_42/carry[1507] ), .COUT(\add_42/carry[1508] ), .SUM(o[1507]) );
  FADDER \add_42/U1_1508  ( .CIN(sreg[1508]), .IN0(n2588), .IN1(
        \add_42/carry[1508] ), .COUT(\add_42/carry[1509] ), .SUM(o[1508]) );
  FADDER \add_42/U1_1509  ( .CIN(sreg[1509]), .IN0(n2587), .IN1(
        \add_42/carry[1509] ), .COUT(\add_42/carry[1510] ), .SUM(o[1509]) );
  FADDER \add_42/U1_1510  ( .CIN(sreg[1510]), .IN0(n2586), .IN1(
        \add_42/carry[1510] ), .COUT(\add_42/carry[1511] ), .SUM(o[1510]) );
  FADDER \add_42/U1_1511  ( .CIN(sreg[1511]), .IN0(n2585), .IN1(
        \add_42/carry[1511] ), .COUT(\add_42/carry[1512] ), .SUM(o[1511]) );
  FADDER \add_42/U1_1512  ( .CIN(sreg[1512]), .IN0(n2584), .IN1(
        \add_42/carry[1512] ), .COUT(\add_42/carry[1513] ), .SUM(o[1512]) );
  FADDER \add_42/U1_1513  ( .CIN(sreg[1513]), .IN0(n2583), .IN1(
        \add_42/carry[1513] ), .COUT(\add_42/carry[1514] ), .SUM(o[1513]) );
  FADDER \add_42/U1_1514  ( .CIN(sreg[1514]), .IN0(n2582), .IN1(
        \add_42/carry[1514] ), .COUT(\add_42/carry[1515] ), .SUM(o[1514]) );
  FADDER \add_42/U1_1515  ( .CIN(sreg[1515]), .IN0(n2581), .IN1(
        \add_42/carry[1515] ), .COUT(\add_42/carry[1516] ), .SUM(o[1515]) );
  FADDER \add_42/U1_1516  ( .CIN(sreg[1516]), .IN0(n2580), .IN1(
        \add_42/carry[1516] ), .COUT(\add_42/carry[1517] ), .SUM(o[1516]) );
  FADDER \add_42/U1_1517  ( .CIN(sreg[1517]), .IN0(n2579), .IN1(
        \add_42/carry[1517] ), .COUT(\add_42/carry[1518] ), .SUM(o[1517]) );
  FADDER \add_42/U1_1518  ( .CIN(sreg[1518]), .IN0(n2578), .IN1(
        \add_42/carry[1518] ), .COUT(\add_42/carry[1519] ), .SUM(o[1518]) );
  FADDER \add_42/U1_1519  ( .CIN(sreg[1519]), .IN0(n2577), .IN1(
        \add_42/carry[1519] ), .COUT(\add_42/carry[1520] ), .SUM(o[1519]) );
  FADDER \add_42/U1_1520  ( .CIN(sreg[1520]), .IN0(n2576), .IN1(
        \add_42/carry[1520] ), .COUT(\add_42/carry[1521] ), .SUM(o[1520]) );
  FADDER \add_42/U1_1521  ( .CIN(sreg[1521]), .IN0(n2575), .IN1(
        \add_42/carry[1521] ), .COUT(\add_42/carry[1522] ), .SUM(o[1521]) );
  FADDER \add_42/U1_1522  ( .CIN(sreg[1522]), .IN0(n2574), .IN1(
        \add_42/carry[1522] ), .COUT(\add_42/carry[1523] ), .SUM(o[1522]) );
  FADDER \add_42/U1_1523  ( .CIN(sreg[1523]), .IN0(n2573), .IN1(
        \add_42/carry[1523] ), .COUT(\add_42/carry[1524] ), .SUM(o[1523]) );
  FADDER \add_42/U1_1524  ( .CIN(sreg[1524]), .IN0(n2572), .IN1(
        \add_42/carry[1524] ), .COUT(\add_42/carry[1525] ), .SUM(o[1524]) );
  FADDER \add_42/U1_1525  ( .CIN(sreg[1525]), .IN0(n2571), .IN1(
        \add_42/carry[1525] ), .COUT(\add_42/carry[1526] ), .SUM(o[1525]) );
  FADDER \add_42/U1_1526  ( .CIN(sreg[1526]), .IN0(n2570), .IN1(
        \add_42/carry[1526] ), .COUT(\add_42/carry[1527] ), .SUM(o[1526]) );
  FADDER \add_42/U1_1527  ( .CIN(sreg[1527]), .IN0(n2569), .IN1(
        \add_42/carry[1527] ), .COUT(\add_42/carry[1528] ), .SUM(o[1527]) );
  FADDER \add_42/U1_1528  ( .CIN(sreg[1528]), .IN0(n2568), .IN1(
        \add_42/carry[1528] ), .COUT(\add_42/carry[1529] ), .SUM(o[1528]) );
  FADDER \add_42/U1_1529  ( .CIN(sreg[1529]), .IN0(n2567), .IN1(
        \add_42/carry[1529] ), .COUT(\add_42/carry[1530] ), .SUM(o[1529]) );
  FADDER \add_42/U1_1530  ( .CIN(sreg[1530]), .IN0(n2566), .IN1(
        \add_42/carry[1530] ), .COUT(\add_42/carry[1531] ), .SUM(o[1530]) );
  FADDER \add_42/U1_1531  ( .CIN(sreg[1531]), .IN0(n2565), .IN1(
        \add_42/carry[1531] ), .COUT(\add_42/carry[1532] ), .SUM(o[1531]) );
  FADDER \add_42/U1_1532  ( .CIN(sreg[1532]), .IN0(n2564), .IN1(
        \add_42/carry[1532] ), .COUT(\add_42/carry[1533] ), .SUM(o[1532]) );
  FADDER \add_42/U1_1533  ( .CIN(sreg[1533]), .IN0(n2563), .IN1(
        \add_42/carry[1533] ), .COUT(\add_42/carry[1534] ), .SUM(o[1533]) );
  FADDER \add_42/U1_1534  ( .CIN(sreg[1534]), .IN0(n2562), .IN1(
        \add_42/carry[1534] ), .COUT(\add_42/carry[1535] ), .SUM(o[1534]) );
  FADDER \add_42/U1_1535  ( .CIN(sreg[1535]), .IN0(n2561), .IN1(
        \add_42/carry[1535] ), .COUT(\add_42/carry[1536] ), .SUM(o[1535]) );
  FADDER \add_42/U1_1536  ( .CIN(sreg[1536]), .IN0(n2560), .IN1(
        \add_42/carry[1536] ), .COUT(\add_42/carry[1537] ), .SUM(o[1536]) );
  FADDER \add_42/U1_1537  ( .CIN(sreg[1537]), .IN0(n2559), .IN1(
        \add_42/carry[1537] ), .COUT(\add_42/carry[1538] ), .SUM(o[1537]) );
  FADDER \add_42/U1_1538  ( .CIN(sreg[1538]), .IN0(n2558), .IN1(
        \add_42/carry[1538] ), .COUT(\add_42/carry[1539] ), .SUM(o[1538]) );
  FADDER \add_42/U1_1539  ( .CIN(sreg[1539]), .IN0(n2557), .IN1(
        \add_42/carry[1539] ), .COUT(\add_42/carry[1540] ), .SUM(o[1539]) );
  FADDER \add_42/U1_1540  ( .CIN(sreg[1540]), .IN0(n2556), .IN1(
        \add_42/carry[1540] ), .COUT(\add_42/carry[1541] ), .SUM(o[1540]) );
  FADDER \add_42/U1_1541  ( .CIN(sreg[1541]), .IN0(n2555), .IN1(
        \add_42/carry[1541] ), .COUT(\add_42/carry[1542] ), .SUM(o[1541]) );
  FADDER \add_42/U1_1542  ( .CIN(sreg[1542]), .IN0(n2554), .IN1(
        \add_42/carry[1542] ), .COUT(\add_42/carry[1543] ), .SUM(o[1542]) );
  FADDER \add_42/U1_1543  ( .CIN(sreg[1543]), .IN0(n2553), .IN1(
        \add_42/carry[1543] ), .COUT(\add_42/carry[1544] ), .SUM(o[1543]) );
  FADDER \add_42/U1_1544  ( .CIN(sreg[1544]), .IN0(n2552), .IN1(
        \add_42/carry[1544] ), .COUT(\add_42/carry[1545] ), .SUM(o[1544]) );
  FADDER \add_42/U1_1545  ( .CIN(sreg[1545]), .IN0(n2551), .IN1(
        \add_42/carry[1545] ), .COUT(\add_42/carry[1546] ), .SUM(o[1545]) );
  FADDER \add_42/U1_1546  ( .CIN(sreg[1546]), .IN0(n2550), .IN1(
        \add_42/carry[1546] ), .COUT(\add_42/carry[1547] ), .SUM(o[1546]) );
  FADDER \add_42/U1_1547  ( .CIN(sreg[1547]), .IN0(n2549), .IN1(
        \add_42/carry[1547] ), .COUT(\add_42/carry[1548] ), .SUM(o[1547]) );
  FADDER \add_42/U1_1548  ( .CIN(sreg[1548]), .IN0(n2548), .IN1(
        \add_42/carry[1548] ), .COUT(\add_42/carry[1549] ), .SUM(o[1548]) );
  FADDER \add_42/U1_1549  ( .CIN(sreg[1549]), .IN0(n2547), .IN1(
        \add_42/carry[1549] ), .COUT(\add_42/carry[1550] ), .SUM(o[1549]) );
  FADDER \add_42/U1_1550  ( .CIN(sreg[1550]), .IN0(n2546), .IN1(
        \add_42/carry[1550] ), .COUT(\add_42/carry[1551] ), .SUM(o[1550]) );
  FADDER \add_42/U1_1551  ( .CIN(sreg[1551]), .IN0(n2545), .IN1(
        \add_42/carry[1551] ), .COUT(\add_42/carry[1552] ), .SUM(o[1551]) );
  FADDER \add_42/U1_1552  ( .CIN(sreg[1552]), .IN0(n2544), .IN1(
        \add_42/carry[1552] ), .COUT(\add_42/carry[1553] ), .SUM(o[1552]) );
  FADDER \add_42/U1_1553  ( .CIN(sreg[1553]), .IN0(n2543), .IN1(
        \add_42/carry[1553] ), .COUT(\add_42/carry[1554] ), .SUM(o[1553]) );
  FADDER \add_42/U1_1554  ( .CIN(sreg[1554]), .IN0(n2542), .IN1(
        \add_42/carry[1554] ), .COUT(\add_42/carry[1555] ), .SUM(o[1554]) );
  FADDER \add_42/U1_1555  ( .CIN(sreg[1555]), .IN0(n2541), .IN1(
        \add_42/carry[1555] ), .COUT(\add_42/carry[1556] ), .SUM(o[1555]) );
  FADDER \add_42/U1_1556  ( .CIN(sreg[1556]), .IN0(n2540), .IN1(
        \add_42/carry[1556] ), .COUT(\add_42/carry[1557] ), .SUM(o[1556]) );
  FADDER \add_42/U1_1557  ( .CIN(sreg[1557]), .IN0(n2539), .IN1(
        \add_42/carry[1557] ), .COUT(\add_42/carry[1558] ), .SUM(o[1557]) );
  FADDER \add_42/U1_1558  ( .CIN(sreg[1558]), .IN0(n2538), .IN1(
        \add_42/carry[1558] ), .COUT(\add_42/carry[1559] ), .SUM(o[1558]) );
  FADDER \add_42/U1_1559  ( .CIN(sreg[1559]), .IN0(n2537), .IN1(
        \add_42/carry[1559] ), .COUT(\add_42/carry[1560] ), .SUM(o[1559]) );
  FADDER \add_42/U1_1560  ( .CIN(sreg[1560]), .IN0(n2536), .IN1(
        \add_42/carry[1560] ), .COUT(\add_42/carry[1561] ), .SUM(o[1560]) );
  FADDER \add_42/U1_1561  ( .CIN(sreg[1561]), .IN0(n2535), .IN1(
        \add_42/carry[1561] ), .COUT(\add_42/carry[1562] ), .SUM(o[1561]) );
  FADDER \add_42/U1_1562  ( .CIN(sreg[1562]), .IN0(n2534), .IN1(
        \add_42/carry[1562] ), .COUT(\add_42/carry[1563] ), .SUM(o[1562]) );
  FADDER \add_42/U1_1563  ( .CIN(sreg[1563]), .IN0(n2533), .IN1(
        \add_42/carry[1563] ), .COUT(\add_42/carry[1564] ), .SUM(o[1563]) );
  FADDER \add_42/U1_1564  ( .CIN(sreg[1564]), .IN0(n2532), .IN1(
        \add_42/carry[1564] ), .COUT(\add_42/carry[1565] ), .SUM(o[1564]) );
  FADDER \add_42/U1_1565  ( .CIN(sreg[1565]), .IN0(n2531), .IN1(
        \add_42/carry[1565] ), .COUT(\add_42/carry[1566] ), .SUM(o[1565]) );
  FADDER \add_42/U1_1566  ( .CIN(sreg[1566]), .IN0(n2530), .IN1(
        \add_42/carry[1566] ), .COUT(\add_42/carry[1567] ), .SUM(o[1566]) );
  FADDER \add_42/U1_1567  ( .CIN(sreg[1567]), .IN0(n2529), .IN1(
        \add_42/carry[1567] ), .COUT(\add_42/carry[1568] ), .SUM(o[1567]) );
  FADDER \add_42/U1_1568  ( .CIN(sreg[1568]), .IN0(n2528), .IN1(
        \add_42/carry[1568] ), .COUT(\add_42/carry[1569] ), .SUM(o[1568]) );
  FADDER \add_42/U1_1569  ( .CIN(sreg[1569]), .IN0(n2527), .IN1(
        \add_42/carry[1569] ), .COUT(\add_42/carry[1570] ), .SUM(o[1569]) );
  FADDER \add_42/U1_1570  ( .CIN(sreg[1570]), .IN0(n2526), .IN1(
        \add_42/carry[1570] ), .COUT(\add_42/carry[1571] ), .SUM(o[1570]) );
  FADDER \add_42/U1_1571  ( .CIN(sreg[1571]), .IN0(n2525), .IN1(
        \add_42/carry[1571] ), .COUT(\add_42/carry[1572] ), .SUM(o[1571]) );
  FADDER \add_42/U1_1572  ( .CIN(sreg[1572]), .IN0(n2524), .IN1(
        \add_42/carry[1572] ), .COUT(\add_42/carry[1573] ), .SUM(o[1572]) );
  FADDER \add_42/U1_1573  ( .CIN(sreg[1573]), .IN0(n2523), .IN1(
        \add_42/carry[1573] ), .COUT(\add_42/carry[1574] ), .SUM(o[1573]) );
  FADDER \add_42/U1_1574  ( .CIN(sreg[1574]), .IN0(n2522), .IN1(
        \add_42/carry[1574] ), .COUT(\add_42/carry[1575] ), .SUM(o[1574]) );
  FADDER \add_42/U1_1575  ( .CIN(sreg[1575]), .IN0(n2521), .IN1(
        \add_42/carry[1575] ), .COUT(\add_42/carry[1576] ), .SUM(o[1575]) );
  FADDER \add_42/U1_1576  ( .CIN(sreg[1576]), .IN0(n2520), .IN1(
        \add_42/carry[1576] ), .COUT(\add_42/carry[1577] ), .SUM(o[1576]) );
  FADDER \add_42/U1_1577  ( .CIN(sreg[1577]), .IN0(n2519), .IN1(
        \add_42/carry[1577] ), .COUT(\add_42/carry[1578] ), .SUM(o[1577]) );
  FADDER \add_42/U1_1578  ( .CIN(sreg[1578]), .IN0(n2518), .IN1(
        \add_42/carry[1578] ), .COUT(\add_42/carry[1579] ), .SUM(o[1578]) );
  FADDER \add_42/U1_1579  ( .CIN(sreg[1579]), .IN0(n2517), .IN1(
        \add_42/carry[1579] ), .COUT(\add_42/carry[1580] ), .SUM(o[1579]) );
  FADDER \add_42/U1_1580  ( .CIN(sreg[1580]), .IN0(n2516), .IN1(
        \add_42/carry[1580] ), .COUT(\add_42/carry[1581] ), .SUM(o[1580]) );
  FADDER \add_42/U1_1581  ( .CIN(sreg[1581]), .IN0(n2515), .IN1(
        \add_42/carry[1581] ), .COUT(\add_42/carry[1582] ), .SUM(o[1581]) );
  FADDER \add_42/U1_1582  ( .CIN(sreg[1582]), .IN0(n2514), .IN1(
        \add_42/carry[1582] ), .COUT(\add_42/carry[1583] ), .SUM(o[1582]) );
  FADDER \add_42/U1_1583  ( .CIN(sreg[1583]), .IN0(n2513), .IN1(
        \add_42/carry[1583] ), .COUT(\add_42/carry[1584] ), .SUM(o[1583]) );
  FADDER \add_42/U1_1584  ( .CIN(sreg[1584]), .IN0(n2512), .IN1(
        \add_42/carry[1584] ), .COUT(\add_42/carry[1585] ), .SUM(o[1584]) );
  FADDER \add_42/U1_1585  ( .CIN(sreg[1585]), .IN0(n2511), .IN1(
        \add_42/carry[1585] ), .COUT(\add_42/carry[1586] ), .SUM(o[1585]) );
  FADDER \add_42/U1_1586  ( .CIN(sreg[1586]), .IN0(n2510), .IN1(
        \add_42/carry[1586] ), .COUT(\add_42/carry[1587] ), .SUM(o[1586]) );
  FADDER \add_42/U1_1587  ( .CIN(sreg[1587]), .IN0(n2509), .IN1(
        \add_42/carry[1587] ), .COUT(\add_42/carry[1588] ), .SUM(o[1587]) );
  FADDER \add_42/U1_1588  ( .CIN(sreg[1588]), .IN0(n2508), .IN1(
        \add_42/carry[1588] ), .COUT(\add_42/carry[1589] ), .SUM(o[1588]) );
  FADDER \add_42/U1_1589  ( .CIN(sreg[1589]), .IN0(n2507), .IN1(
        \add_42/carry[1589] ), .COUT(\add_42/carry[1590] ), .SUM(o[1589]) );
  FADDER \add_42/U1_1590  ( .CIN(sreg[1590]), .IN0(n2506), .IN1(
        \add_42/carry[1590] ), .COUT(\add_42/carry[1591] ), .SUM(o[1590]) );
  FADDER \add_42/U1_1591  ( .CIN(sreg[1591]), .IN0(n2505), .IN1(
        \add_42/carry[1591] ), .COUT(\add_42/carry[1592] ), .SUM(o[1591]) );
  FADDER \add_42/U1_1592  ( .CIN(sreg[1592]), .IN0(n2504), .IN1(
        \add_42/carry[1592] ), .COUT(\add_42/carry[1593] ), .SUM(o[1592]) );
  FADDER \add_42/U1_1593  ( .CIN(sreg[1593]), .IN0(n2503), .IN1(
        \add_42/carry[1593] ), .COUT(\add_42/carry[1594] ), .SUM(o[1593]) );
  FADDER \add_42/U1_1594  ( .CIN(sreg[1594]), .IN0(n2502), .IN1(
        \add_42/carry[1594] ), .COUT(\add_42/carry[1595] ), .SUM(o[1594]) );
  FADDER \add_42/U1_1595  ( .CIN(sreg[1595]), .IN0(n2501), .IN1(
        \add_42/carry[1595] ), .COUT(\add_42/carry[1596] ), .SUM(o[1595]) );
  FADDER \add_42/U1_1596  ( .CIN(sreg[1596]), .IN0(n2500), .IN1(
        \add_42/carry[1596] ), .COUT(\add_42/carry[1597] ), .SUM(o[1596]) );
  FADDER \add_42/U1_1597  ( .CIN(sreg[1597]), .IN0(n2499), .IN1(
        \add_42/carry[1597] ), .COUT(\add_42/carry[1598] ), .SUM(o[1597]) );
  FADDER \add_42/U1_1598  ( .CIN(sreg[1598]), .IN0(n2498), .IN1(
        \add_42/carry[1598] ), .COUT(\add_42/carry[1599] ), .SUM(o[1598]) );
  FADDER \add_42/U1_1599  ( .CIN(sreg[1599]), .IN0(n2497), .IN1(
        \add_42/carry[1599] ), .COUT(\add_42/carry[1600] ), .SUM(o[1599]) );
  FADDER \add_42/U1_1600  ( .CIN(sreg[1600]), .IN0(n2496), .IN1(
        \add_42/carry[1600] ), .COUT(\add_42/carry[1601] ), .SUM(o[1600]) );
  FADDER \add_42/U1_1601  ( .CIN(sreg[1601]), .IN0(n2495), .IN1(
        \add_42/carry[1601] ), .COUT(\add_42/carry[1602] ), .SUM(o[1601]) );
  FADDER \add_42/U1_1602  ( .CIN(sreg[1602]), .IN0(n2494), .IN1(
        \add_42/carry[1602] ), .COUT(\add_42/carry[1603] ), .SUM(o[1602]) );
  FADDER \add_42/U1_1603  ( .CIN(sreg[1603]), .IN0(n2493), .IN1(
        \add_42/carry[1603] ), .COUT(\add_42/carry[1604] ), .SUM(o[1603]) );
  FADDER \add_42/U1_1604  ( .CIN(sreg[1604]), .IN0(n2492), .IN1(
        \add_42/carry[1604] ), .COUT(\add_42/carry[1605] ), .SUM(o[1604]) );
  FADDER \add_42/U1_1605  ( .CIN(sreg[1605]), .IN0(n2491), .IN1(
        \add_42/carry[1605] ), .COUT(\add_42/carry[1606] ), .SUM(o[1605]) );
  FADDER \add_42/U1_1606  ( .CIN(sreg[1606]), .IN0(n2490), .IN1(
        \add_42/carry[1606] ), .COUT(\add_42/carry[1607] ), .SUM(o[1606]) );
  FADDER \add_42/U1_1607  ( .CIN(sreg[1607]), .IN0(n2489), .IN1(
        \add_42/carry[1607] ), .COUT(\add_42/carry[1608] ), .SUM(o[1607]) );
  FADDER \add_42/U1_1608  ( .CIN(sreg[1608]), .IN0(n2488), .IN1(
        \add_42/carry[1608] ), .COUT(\add_42/carry[1609] ), .SUM(o[1608]) );
  FADDER \add_42/U1_1609  ( .CIN(sreg[1609]), .IN0(n2487), .IN1(
        \add_42/carry[1609] ), .COUT(\add_42/carry[1610] ), .SUM(o[1609]) );
  FADDER \add_42/U1_1610  ( .CIN(sreg[1610]), .IN0(n2486), .IN1(
        \add_42/carry[1610] ), .COUT(\add_42/carry[1611] ), .SUM(o[1610]) );
  FADDER \add_42/U1_1611  ( .CIN(sreg[1611]), .IN0(n2485), .IN1(
        \add_42/carry[1611] ), .COUT(\add_42/carry[1612] ), .SUM(o[1611]) );
  FADDER \add_42/U1_1612  ( .CIN(sreg[1612]), .IN0(n2484), .IN1(
        \add_42/carry[1612] ), .COUT(\add_42/carry[1613] ), .SUM(o[1612]) );
  FADDER \add_42/U1_1613  ( .CIN(sreg[1613]), .IN0(n2483), .IN1(
        \add_42/carry[1613] ), .COUT(\add_42/carry[1614] ), .SUM(o[1613]) );
  FADDER \add_42/U1_1614  ( .CIN(sreg[1614]), .IN0(n2482), .IN1(
        \add_42/carry[1614] ), .COUT(\add_42/carry[1615] ), .SUM(o[1614]) );
  FADDER \add_42/U1_1615  ( .CIN(sreg[1615]), .IN0(n2481), .IN1(
        \add_42/carry[1615] ), .COUT(\add_42/carry[1616] ), .SUM(o[1615]) );
  FADDER \add_42/U1_1616  ( .CIN(sreg[1616]), .IN0(n2480), .IN1(
        \add_42/carry[1616] ), .COUT(\add_42/carry[1617] ), .SUM(o[1616]) );
  FADDER \add_42/U1_1617  ( .CIN(sreg[1617]), .IN0(n2479), .IN1(
        \add_42/carry[1617] ), .COUT(\add_42/carry[1618] ), .SUM(o[1617]) );
  FADDER \add_42/U1_1618  ( .CIN(sreg[1618]), .IN0(n2478), .IN1(
        \add_42/carry[1618] ), .COUT(\add_42/carry[1619] ), .SUM(o[1618]) );
  FADDER \add_42/U1_1619  ( .CIN(sreg[1619]), .IN0(n2477), .IN1(
        \add_42/carry[1619] ), .COUT(\add_42/carry[1620] ), .SUM(o[1619]) );
  FADDER \add_42/U1_1620  ( .CIN(sreg[1620]), .IN0(n2476), .IN1(
        \add_42/carry[1620] ), .COUT(\add_42/carry[1621] ), .SUM(o[1620]) );
  FADDER \add_42/U1_1621  ( .CIN(sreg[1621]), .IN0(n2475), .IN1(
        \add_42/carry[1621] ), .COUT(\add_42/carry[1622] ), .SUM(o[1621]) );
  FADDER \add_42/U1_1622  ( .CIN(sreg[1622]), .IN0(n2474), .IN1(
        \add_42/carry[1622] ), .COUT(\add_42/carry[1623] ), .SUM(o[1622]) );
  FADDER \add_42/U1_1623  ( .CIN(sreg[1623]), .IN0(n2473), .IN1(
        \add_42/carry[1623] ), .COUT(\add_42/carry[1624] ), .SUM(o[1623]) );
  FADDER \add_42/U1_1624  ( .CIN(sreg[1624]), .IN0(n2472), .IN1(
        \add_42/carry[1624] ), .COUT(\add_42/carry[1625] ), .SUM(o[1624]) );
  FADDER \add_42/U1_1625  ( .CIN(sreg[1625]), .IN0(n2471), .IN1(
        \add_42/carry[1625] ), .COUT(\add_42/carry[1626] ), .SUM(o[1625]) );
  FADDER \add_42/U1_1626  ( .CIN(sreg[1626]), .IN0(n2470), .IN1(
        \add_42/carry[1626] ), .COUT(\add_42/carry[1627] ), .SUM(o[1626]) );
  FADDER \add_42/U1_1627  ( .CIN(sreg[1627]), .IN0(n2469), .IN1(
        \add_42/carry[1627] ), .COUT(\add_42/carry[1628] ), .SUM(o[1627]) );
  FADDER \add_42/U1_1628  ( .CIN(sreg[1628]), .IN0(n2468), .IN1(
        \add_42/carry[1628] ), .COUT(\add_42/carry[1629] ), .SUM(o[1628]) );
  FADDER \add_42/U1_1629  ( .CIN(sreg[1629]), .IN0(n2467), .IN1(
        \add_42/carry[1629] ), .COUT(\add_42/carry[1630] ), .SUM(o[1629]) );
  FADDER \add_42/U1_1630  ( .CIN(sreg[1630]), .IN0(n2466), .IN1(
        \add_42/carry[1630] ), .COUT(\add_42/carry[1631] ), .SUM(o[1630]) );
  FADDER \add_42/U1_1631  ( .CIN(sreg[1631]), .IN0(n2465), .IN1(
        \add_42/carry[1631] ), .COUT(\add_42/carry[1632] ), .SUM(o[1631]) );
  FADDER \add_42/U1_1632  ( .CIN(sreg[1632]), .IN0(n2464), .IN1(
        \add_42/carry[1632] ), .COUT(\add_42/carry[1633] ), .SUM(o[1632]) );
  FADDER \add_42/U1_1633  ( .CIN(sreg[1633]), .IN0(n2463), .IN1(
        \add_42/carry[1633] ), .COUT(\add_42/carry[1634] ), .SUM(o[1633]) );
  FADDER \add_42/U1_1634  ( .CIN(sreg[1634]), .IN0(n2462), .IN1(
        \add_42/carry[1634] ), .COUT(\add_42/carry[1635] ), .SUM(o[1634]) );
  FADDER \add_42/U1_1635  ( .CIN(sreg[1635]), .IN0(n2461), .IN1(
        \add_42/carry[1635] ), .COUT(\add_42/carry[1636] ), .SUM(o[1635]) );
  FADDER \add_42/U1_1636  ( .CIN(sreg[1636]), .IN0(n2460), .IN1(
        \add_42/carry[1636] ), .COUT(\add_42/carry[1637] ), .SUM(o[1636]) );
  FADDER \add_42/U1_1637  ( .CIN(sreg[1637]), .IN0(n2459), .IN1(
        \add_42/carry[1637] ), .COUT(\add_42/carry[1638] ), .SUM(o[1637]) );
  FADDER \add_42/U1_1638  ( .CIN(sreg[1638]), .IN0(n2458), .IN1(
        \add_42/carry[1638] ), .COUT(\add_42/carry[1639] ), .SUM(o[1638]) );
  FADDER \add_42/U1_1639  ( .CIN(sreg[1639]), .IN0(n2457), .IN1(
        \add_42/carry[1639] ), .COUT(\add_42/carry[1640] ), .SUM(o[1639]) );
  FADDER \add_42/U1_1640  ( .CIN(sreg[1640]), .IN0(n2456), .IN1(
        \add_42/carry[1640] ), .COUT(\add_42/carry[1641] ), .SUM(o[1640]) );
  FADDER \add_42/U1_1641  ( .CIN(sreg[1641]), .IN0(n2455), .IN1(
        \add_42/carry[1641] ), .COUT(\add_42/carry[1642] ), .SUM(o[1641]) );
  FADDER \add_42/U1_1642  ( .CIN(sreg[1642]), .IN0(n2454), .IN1(
        \add_42/carry[1642] ), .COUT(\add_42/carry[1643] ), .SUM(o[1642]) );
  FADDER \add_42/U1_1643  ( .CIN(sreg[1643]), .IN0(n2453), .IN1(
        \add_42/carry[1643] ), .COUT(\add_42/carry[1644] ), .SUM(o[1643]) );
  FADDER \add_42/U1_1644  ( .CIN(sreg[1644]), .IN0(n2452), .IN1(
        \add_42/carry[1644] ), .COUT(\add_42/carry[1645] ), .SUM(o[1644]) );
  FADDER \add_42/U1_1645  ( .CIN(sreg[1645]), .IN0(n2451), .IN1(
        \add_42/carry[1645] ), .COUT(\add_42/carry[1646] ), .SUM(o[1645]) );
  FADDER \add_42/U1_1646  ( .CIN(sreg[1646]), .IN0(n2450), .IN1(
        \add_42/carry[1646] ), .COUT(\add_42/carry[1647] ), .SUM(o[1646]) );
  FADDER \add_42/U1_1647  ( .CIN(sreg[1647]), .IN0(n2449), .IN1(
        \add_42/carry[1647] ), .COUT(\add_42/carry[1648] ), .SUM(o[1647]) );
  FADDER \add_42/U1_1648  ( .CIN(sreg[1648]), .IN0(n2448), .IN1(
        \add_42/carry[1648] ), .COUT(\add_42/carry[1649] ), .SUM(o[1648]) );
  FADDER \add_42/U1_1649  ( .CIN(sreg[1649]), .IN0(n2447), .IN1(
        \add_42/carry[1649] ), .COUT(\add_42/carry[1650] ), .SUM(o[1649]) );
  FADDER \add_42/U1_1650  ( .CIN(sreg[1650]), .IN0(n2446), .IN1(
        \add_42/carry[1650] ), .COUT(\add_42/carry[1651] ), .SUM(o[1650]) );
  FADDER \add_42/U1_1651  ( .CIN(sreg[1651]), .IN0(n2445), .IN1(
        \add_42/carry[1651] ), .COUT(\add_42/carry[1652] ), .SUM(o[1651]) );
  FADDER \add_42/U1_1652  ( .CIN(sreg[1652]), .IN0(n2444), .IN1(
        \add_42/carry[1652] ), .COUT(\add_42/carry[1653] ), .SUM(o[1652]) );
  FADDER \add_42/U1_1653  ( .CIN(sreg[1653]), .IN0(n2443), .IN1(
        \add_42/carry[1653] ), .COUT(\add_42/carry[1654] ), .SUM(o[1653]) );
  FADDER \add_42/U1_1654  ( .CIN(sreg[1654]), .IN0(n2442), .IN1(
        \add_42/carry[1654] ), .COUT(\add_42/carry[1655] ), .SUM(o[1654]) );
  FADDER \add_42/U1_1655  ( .CIN(sreg[1655]), .IN0(n2441), .IN1(
        \add_42/carry[1655] ), .COUT(\add_42/carry[1656] ), .SUM(o[1655]) );
  FADDER \add_42/U1_1656  ( .CIN(sreg[1656]), .IN0(n2440), .IN1(
        \add_42/carry[1656] ), .COUT(\add_42/carry[1657] ), .SUM(o[1656]) );
  FADDER \add_42/U1_1657  ( .CIN(sreg[1657]), .IN0(n2439), .IN1(
        \add_42/carry[1657] ), .COUT(\add_42/carry[1658] ), .SUM(o[1657]) );
  FADDER \add_42/U1_1658  ( .CIN(sreg[1658]), .IN0(n2438), .IN1(
        \add_42/carry[1658] ), .COUT(\add_42/carry[1659] ), .SUM(o[1658]) );
  FADDER \add_42/U1_1659  ( .CIN(sreg[1659]), .IN0(n2437), .IN1(
        \add_42/carry[1659] ), .COUT(\add_42/carry[1660] ), .SUM(o[1659]) );
  FADDER \add_42/U1_1660  ( .CIN(sreg[1660]), .IN0(n2436), .IN1(
        \add_42/carry[1660] ), .COUT(\add_42/carry[1661] ), .SUM(o[1660]) );
  FADDER \add_42/U1_1661  ( .CIN(sreg[1661]), .IN0(n2435), .IN1(
        \add_42/carry[1661] ), .COUT(\add_42/carry[1662] ), .SUM(o[1661]) );
  FADDER \add_42/U1_1662  ( .CIN(sreg[1662]), .IN0(n2434), .IN1(
        \add_42/carry[1662] ), .COUT(\add_42/carry[1663] ), .SUM(o[1662]) );
  FADDER \add_42/U1_1663  ( .CIN(sreg[1663]), .IN0(n2433), .IN1(
        \add_42/carry[1663] ), .COUT(\add_42/carry[1664] ), .SUM(o[1663]) );
  FADDER \add_42/U1_1664  ( .CIN(sreg[1664]), .IN0(n2432), .IN1(
        \add_42/carry[1664] ), .COUT(\add_42/carry[1665] ), .SUM(o[1664]) );
  FADDER \add_42/U1_1665  ( .CIN(sreg[1665]), .IN0(n2431), .IN1(
        \add_42/carry[1665] ), .COUT(\add_42/carry[1666] ), .SUM(o[1665]) );
  FADDER \add_42/U1_1666  ( .CIN(sreg[1666]), .IN0(n2430), .IN1(
        \add_42/carry[1666] ), .COUT(\add_42/carry[1667] ), .SUM(o[1666]) );
  FADDER \add_42/U1_1667  ( .CIN(sreg[1667]), .IN0(n2429), .IN1(
        \add_42/carry[1667] ), .COUT(\add_42/carry[1668] ), .SUM(o[1667]) );
  FADDER \add_42/U1_1668  ( .CIN(sreg[1668]), .IN0(n2428), .IN1(
        \add_42/carry[1668] ), .COUT(\add_42/carry[1669] ), .SUM(o[1668]) );
  FADDER \add_42/U1_1669  ( .CIN(sreg[1669]), .IN0(n2427), .IN1(
        \add_42/carry[1669] ), .COUT(\add_42/carry[1670] ), .SUM(o[1669]) );
  FADDER \add_42/U1_1670  ( .CIN(sreg[1670]), .IN0(n2426), .IN1(
        \add_42/carry[1670] ), .COUT(\add_42/carry[1671] ), .SUM(o[1670]) );
  FADDER \add_42/U1_1671  ( .CIN(sreg[1671]), .IN0(n2425), .IN1(
        \add_42/carry[1671] ), .COUT(\add_42/carry[1672] ), .SUM(o[1671]) );
  FADDER \add_42/U1_1672  ( .CIN(sreg[1672]), .IN0(n2424), .IN1(
        \add_42/carry[1672] ), .COUT(\add_42/carry[1673] ), .SUM(o[1672]) );
  FADDER \add_42/U1_1673  ( .CIN(sreg[1673]), .IN0(n2423), .IN1(
        \add_42/carry[1673] ), .COUT(\add_42/carry[1674] ), .SUM(o[1673]) );
  FADDER \add_42/U1_1674  ( .CIN(sreg[1674]), .IN0(n2422), .IN1(
        \add_42/carry[1674] ), .COUT(\add_42/carry[1675] ), .SUM(o[1674]) );
  FADDER \add_42/U1_1675  ( .CIN(sreg[1675]), .IN0(n2421), .IN1(
        \add_42/carry[1675] ), .COUT(\add_42/carry[1676] ), .SUM(o[1675]) );
  FADDER \add_42/U1_1676  ( .CIN(sreg[1676]), .IN0(n2420), .IN1(
        \add_42/carry[1676] ), .COUT(\add_42/carry[1677] ), .SUM(o[1676]) );
  FADDER \add_42/U1_1677  ( .CIN(sreg[1677]), .IN0(n2419), .IN1(
        \add_42/carry[1677] ), .COUT(\add_42/carry[1678] ), .SUM(o[1677]) );
  FADDER \add_42/U1_1678  ( .CIN(sreg[1678]), .IN0(n2418), .IN1(
        \add_42/carry[1678] ), .COUT(\add_42/carry[1679] ), .SUM(o[1678]) );
  FADDER \add_42/U1_1679  ( .CIN(sreg[1679]), .IN0(n2417), .IN1(
        \add_42/carry[1679] ), .COUT(\add_42/carry[1680] ), .SUM(o[1679]) );
  FADDER \add_42/U1_1680  ( .CIN(sreg[1680]), .IN0(n2416), .IN1(
        \add_42/carry[1680] ), .COUT(\add_42/carry[1681] ), .SUM(o[1680]) );
  FADDER \add_42/U1_1681  ( .CIN(sreg[1681]), .IN0(n2415), .IN1(
        \add_42/carry[1681] ), .COUT(\add_42/carry[1682] ), .SUM(o[1681]) );
  FADDER \add_42/U1_1682  ( .CIN(sreg[1682]), .IN0(n2414), .IN1(
        \add_42/carry[1682] ), .COUT(\add_42/carry[1683] ), .SUM(o[1682]) );
  FADDER \add_42/U1_1683  ( .CIN(sreg[1683]), .IN0(n2413), .IN1(
        \add_42/carry[1683] ), .COUT(\add_42/carry[1684] ), .SUM(o[1683]) );
  FADDER \add_42/U1_1684  ( .CIN(sreg[1684]), .IN0(n2412), .IN1(
        \add_42/carry[1684] ), .COUT(\add_42/carry[1685] ), .SUM(o[1684]) );
  FADDER \add_42/U1_1685  ( .CIN(sreg[1685]), .IN0(n2411), .IN1(
        \add_42/carry[1685] ), .COUT(\add_42/carry[1686] ), .SUM(o[1685]) );
  FADDER \add_42/U1_1686  ( .CIN(sreg[1686]), .IN0(n2410), .IN1(
        \add_42/carry[1686] ), .COUT(\add_42/carry[1687] ), .SUM(o[1686]) );
  FADDER \add_42/U1_1687  ( .CIN(sreg[1687]), .IN0(n2409), .IN1(
        \add_42/carry[1687] ), .COUT(\add_42/carry[1688] ), .SUM(o[1687]) );
  FADDER \add_42/U1_1688  ( .CIN(sreg[1688]), .IN0(n2408), .IN1(
        \add_42/carry[1688] ), .COUT(\add_42/carry[1689] ), .SUM(o[1688]) );
  FADDER \add_42/U1_1689  ( .CIN(sreg[1689]), .IN0(n2407), .IN1(
        \add_42/carry[1689] ), .COUT(\add_42/carry[1690] ), .SUM(o[1689]) );
  FADDER \add_42/U1_1690  ( .CIN(sreg[1690]), .IN0(n2406), .IN1(
        \add_42/carry[1690] ), .COUT(\add_42/carry[1691] ), .SUM(o[1690]) );
  FADDER \add_42/U1_1691  ( .CIN(sreg[1691]), .IN0(n2405), .IN1(
        \add_42/carry[1691] ), .COUT(\add_42/carry[1692] ), .SUM(o[1691]) );
  FADDER \add_42/U1_1692  ( .CIN(sreg[1692]), .IN0(n2404), .IN1(
        \add_42/carry[1692] ), .COUT(\add_42/carry[1693] ), .SUM(o[1692]) );
  FADDER \add_42/U1_1693  ( .CIN(sreg[1693]), .IN0(n2403), .IN1(
        \add_42/carry[1693] ), .COUT(\add_42/carry[1694] ), .SUM(o[1693]) );
  FADDER \add_42/U1_1694  ( .CIN(sreg[1694]), .IN0(n2402), .IN1(
        \add_42/carry[1694] ), .COUT(\add_42/carry[1695] ), .SUM(o[1694]) );
  FADDER \add_42/U1_1695  ( .CIN(sreg[1695]), .IN0(n2401), .IN1(
        \add_42/carry[1695] ), .COUT(\add_42/carry[1696] ), .SUM(o[1695]) );
  FADDER \add_42/U1_1696  ( .CIN(sreg[1696]), .IN0(n2400), .IN1(
        \add_42/carry[1696] ), .COUT(\add_42/carry[1697] ), .SUM(o[1696]) );
  FADDER \add_42/U1_1697  ( .CIN(sreg[1697]), .IN0(n2399), .IN1(
        \add_42/carry[1697] ), .COUT(\add_42/carry[1698] ), .SUM(o[1697]) );
  FADDER \add_42/U1_1698  ( .CIN(sreg[1698]), .IN0(n2398), .IN1(
        \add_42/carry[1698] ), .COUT(\add_42/carry[1699] ), .SUM(o[1698]) );
  FADDER \add_42/U1_1699  ( .CIN(sreg[1699]), .IN0(n2397), .IN1(
        \add_42/carry[1699] ), .COUT(\add_42/carry[1700] ), .SUM(o[1699]) );
  FADDER \add_42/U1_1700  ( .CIN(sreg[1700]), .IN0(n2396), .IN1(
        \add_42/carry[1700] ), .COUT(\add_42/carry[1701] ), .SUM(o[1700]) );
  FADDER \add_42/U1_1701  ( .CIN(sreg[1701]), .IN0(n2395), .IN1(
        \add_42/carry[1701] ), .COUT(\add_42/carry[1702] ), .SUM(o[1701]) );
  FADDER \add_42/U1_1702  ( .CIN(sreg[1702]), .IN0(n2394), .IN1(
        \add_42/carry[1702] ), .COUT(\add_42/carry[1703] ), .SUM(o[1702]) );
  FADDER \add_42/U1_1703  ( .CIN(sreg[1703]), .IN0(n2393), .IN1(
        \add_42/carry[1703] ), .COUT(\add_42/carry[1704] ), .SUM(o[1703]) );
  FADDER \add_42/U1_1704  ( .CIN(sreg[1704]), .IN0(n2392), .IN1(
        \add_42/carry[1704] ), .COUT(\add_42/carry[1705] ), .SUM(o[1704]) );
  FADDER \add_42/U1_1705  ( .CIN(sreg[1705]), .IN0(n2391), .IN1(
        \add_42/carry[1705] ), .COUT(\add_42/carry[1706] ), .SUM(o[1705]) );
  FADDER \add_42/U1_1706  ( .CIN(sreg[1706]), .IN0(n2390), .IN1(
        \add_42/carry[1706] ), .COUT(\add_42/carry[1707] ), .SUM(o[1706]) );
  FADDER \add_42/U1_1707  ( .CIN(sreg[1707]), .IN0(n2389), .IN1(
        \add_42/carry[1707] ), .COUT(\add_42/carry[1708] ), .SUM(o[1707]) );
  FADDER \add_42/U1_1708  ( .CIN(sreg[1708]), .IN0(n2388), .IN1(
        \add_42/carry[1708] ), .COUT(\add_42/carry[1709] ), .SUM(o[1708]) );
  FADDER \add_42/U1_1709  ( .CIN(sreg[1709]), .IN0(n2387), .IN1(
        \add_42/carry[1709] ), .COUT(\add_42/carry[1710] ), .SUM(o[1709]) );
  FADDER \add_42/U1_1710  ( .CIN(sreg[1710]), .IN0(n2386), .IN1(
        \add_42/carry[1710] ), .COUT(\add_42/carry[1711] ), .SUM(o[1710]) );
  FADDER \add_42/U1_1711  ( .CIN(sreg[1711]), .IN0(n2385), .IN1(
        \add_42/carry[1711] ), .COUT(\add_42/carry[1712] ), .SUM(o[1711]) );
  FADDER \add_42/U1_1712  ( .CIN(sreg[1712]), .IN0(n2384), .IN1(
        \add_42/carry[1712] ), .COUT(\add_42/carry[1713] ), .SUM(o[1712]) );
  FADDER \add_42/U1_1713  ( .CIN(sreg[1713]), .IN0(n2383), .IN1(
        \add_42/carry[1713] ), .COUT(\add_42/carry[1714] ), .SUM(o[1713]) );
  FADDER \add_42/U1_1714  ( .CIN(sreg[1714]), .IN0(n2382), .IN1(
        \add_42/carry[1714] ), .COUT(\add_42/carry[1715] ), .SUM(o[1714]) );
  FADDER \add_42/U1_1715  ( .CIN(sreg[1715]), .IN0(n2381), .IN1(
        \add_42/carry[1715] ), .COUT(\add_42/carry[1716] ), .SUM(o[1715]) );
  FADDER \add_42/U1_1716  ( .CIN(sreg[1716]), .IN0(n2380), .IN1(
        \add_42/carry[1716] ), .COUT(\add_42/carry[1717] ), .SUM(o[1716]) );
  FADDER \add_42/U1_1717  ( .CIN(sreg[1717]), .IN0(n2379), .IN1(
        \add_42/carry[1717] ), .COUT(\add_42/carry[1718] ), .SUM(o[1717]) );
  FADDER \add_42/U1_1718  ( .CIN(sreg[1718]), .IN0(n2378), .IN1(
        \add_42/carry[1718] ), .COUT(\add_42/carry[1719] ), .SUM(o[1718]) );
  FADDER \add_42/U1_1719  ( .CIN(sreg[1719]), .IN0(n2377), .IN1(
        \add_42/carry[1719] ), .COUT(\add_42/carry[1720] ), .SUM(o[1719]) );
  FADDER \add_42/U1_1720  ( .CIN(sreg[1720]), .IN0(n2376), .IN1(
        \add_42/carry[1720] ), .COUT(\add_42/carry[1721] ), .SUM(o[1720]) );
  FADDER \add_42/U1_1721  ( .CIN(sreg[1721]), .IN0(n2375), .IN1(
        \add_42/carry[1721] ), .COUT(\add_42/carry[1722] ), .SUM(o[1721]) );
  FADDER \add_42/U1_1722  ( .CIN(sreg[1722]), .IN0(n2374), .IN1(
        \add_42/carry[1722] ), .COUT(\add_42/carry[1723] ), .SUM(o[1722]) );
  FADDER \add_42/U1_1723  ( .CIN(sreg[1723]), .IN0(n2373), .IN1(
        \add_42/carry[1723] ), .COUT(\add_42/carry[1724] ), .SUM(o[1723]) );
  FADDER \add_42/U1_1724  ( .CIN(sreg[1724]), .IN0(n2372), .IN1(
        \add_42/carry[1724] ), .COUT(\add_42/carry[1725] ), .SUM(o[1724]) );
  FADDER \add_42/U1_1725  ( .CIN(sreg[1725]), .IN0(n2371), .IN1(
        \add_42/carry[1725] ), .COUT(\add_42/carry[1726] ), .SUM(o[1725]) );
  FADDER \add_42/U1_1726  ( .CIN(sreg[1726]), .IN0(n2370), .IN1(
        \add_42/carry[1726] ), .COUT(\add_42/carry[1727] ), .SUM(o[1726]) );
  FADDER \add_42/U1_1727  ( .CIN(sreg[1727]), .IN0(n2369), .IN1(
        \add_42/carry[1727] ), .COUT(\add_42/carry[1728] ), .SUM(o[1727]) );
  FADDER \add_42/U1_1728  ( .CIN(sreg[1728]), .IN0(n2368), .IN1(
        \add_42/carry[1728] ), .COUT(\add_42/carry[1729] ), .SUM(o[1728]) );
  FADDER \add_42/U1_1729  ( .CIN(sreg[1729]), .IN0(n2367), .IN1(
        \add_42/carry[1729] ), .COUT(\add_42/carry[1730] ), .SUM(o[1729]) );
  FADDER \add_42/U1_1730  ( .CIN(sreg[1730]), .IN0(n2366), .IN1(
        \add_42/carry[1730] ), .COUT(\add_42/carry[1731] ), .SUM(o[1730]) );
  FADDER \add_42/U1_1731  ( .CIN(sreg[1731]), .IN0(n2365), .IN1(
        \add_42/carry[1731] ), .COUT(\add_42/carry[1732] ), .SUM(o[1731]) );
  FADDER \add_42/U1_1732  ( .CIN(sreg[1732]), .IN0(n2364), .IN1(
        \add_42/carry[1732] ), .COUT(\add_42/carry[1733] ), .SUM(o[1732]) );
  FADDER \add_42/U1_1733  ( .CIN(sreg[1733]), .IN0(n2363), .IN1(
        \add_42/carry[1733] ), .COUT(\add_42/carry[1734] ), .SUM(o[1733]) );
  FADDER \add_42/U1_1734  ( .CIN(sreg[1734]), .IN0(n2362), .IN1(
        \add_42/carry[1734] ), .COUT(\add_42/carry[1735] ), .SUM(o[1734]) );
  FADDER \add_42/U1_1735  ( .CIN(sreg[1735]), .IN0(n2361), .IN1(
        \add_42/carry[1735] ), .COUT(\add_42/carry[1736] ), .SUM(o[1735]) );
  FADDER \add_42/U1_1736  ( .CIN(sreg[1736]), .IN0(n2360), .IN1(
        \add_42/carry[1736] ), .COUT(\add_42/carry[1737] ), .SUM(o[1736]) );
  FADDER \add_42/U1_1737  ( .CIN(sreg[1737]), .IN0(n2359), .IN1(
        \add_42/carry[1737] ), .COUT(\add_42/carry[1738] ), .SUM(o[1737]) );
  FADDER \add_42/U1_1738  ( .CIN(sreg[1738]), .IN0(n2358), .IN1(
        \add_42/carry[1738] ), .COUT(\add_42/carry[1739] ), .SUM(o[1738]) );
  FADDER \add_42/U1_1739  ( .CIN(sreg[1739]), .IN0(n2357), .IN1(
        \add_42/carry[1739] ), .COUT(\add_42/carry[1740] ), .SUM(o[1739]) );
  FADDER \add_42/U1_1740  ( .CIN(sreg[1740]), .IN0(n2356), .IN1(
        \add_42/carry[1740] ), .COUT(\add_42/carry[1741] ), .SUM(o[1740]) );
  FADDER \add_42/U1_1741  ( .CIN(sreg[1741]), .IN0(n2355), .IN1(
        \add_42/carry[1741] ), .COUT(\add_42/carry[1742] ), .SUM(o[1741]) );
  FADDER \add_42/U1_1742  ( .CIN(sreg[1742]), .IN0(n2354), .IN1(
        \add_42/carry[1742] ), .COUT(\add_42/carry[1743] ), .SUM(o[1742]) );
  FADDER \add_42/U1_1743  ( .CIN(sreg[1743]), .IN0(n2353), .IN1(
        \add_42/carry[1743] ), .COUT(\add_42/carry[1744] ), .SUM(o[1743]) );
  FADDER \add_42/U1_1744  ( .CIN(sreg[1744]), .IN0(n2352), .IN1(
        \add_42/carry[1744] ), .COUT(\add_42/carry[1745] ), .SUM(o[1744]) );
  FADDER \add_42/U1_1745  ( .CIN(sreg[1745]), .IN0(n2351), .IN1(
        \add_42/carry[1745] ), .COUT(\add_42/carry[1746] ), .SUM(o[1745]) );
  FADDER \add_42/U1_1746  ( .CIN(sreg[1746]), .IN0(n2350), .IN1(
        \add_42/carry[1746] ), .COUT(\add_42/carry[1747] ), .SUM(o[1746]) );
  FADDER \add_42/U1_1747  ( .CIN(sreg[1747]), .IN0(n2349), .IN1(
        \add_42/carry[1747] ), .COUT(\add_42/carry[1748] ), .SUM(o[1747]) );
  FADDER \add_42/U1_1748  ( .CIN(sreg[1748]), .IN0(n2348), .IN1(
        \add_42/carry[1748] ), .COUT(\add_42/carry[1749] ), .SUM(o[1748]) );
  FADDER \add_42/U1_1749  ( .CIN(sreg[1749]), .IN0(n2347), .IN1(
        \add_42/carry[1749] ), .COUT(\add_42/carry[1750] ), .SUM(o[1749]) );
  FADDER \add_42/U1_1750  ( .CIN(sreg[1750]), .IN0(n2346), .IN1(
        \add_42/carry[1750] ), .COUT(\add_42/carry[1751] ), .SUM(o[1750]) );
  FADDER \add_42/U1_1751  ( .CIN(sreg[1751]), .IN0(n2345), .IN1(
        \add_42/carry[1751] ), .COUT(\add_42/carry[1752] ), .SUM(o[1751]) );
  FADDER \add_42/U1_1752  ( .CIN(sreg[1752]), .IN0(n2344), .IN1(
        \add_42/carry[1752] ), .COUT(\add_42/carry[1753] ), .SUM(o[1752]) );
  FADDER \add_42/U1_1753  ( .CIN(sreg[1753]), .IN0(n2343), .IN1(
        \add_42/carry[1753] ), .COUT(\add_42/carry[1754] ), .SUM(o[1753]) );
  FADDER \add_42/U1_1754  ( .CIN(sreg[1754]), .IN0(n2342), .IN1(
        \add_42/carry[1754] ), .COUT(\add_42/carry[1755] ), .SUM(o[1754]) );
  FADDER \add_42/U1_1755  ( .CIN(sreg[1755]), .IN0(n2341), .IN1(
        \add_42/carry[1755] ), .COUT(\add_42/carry[1756] ), .SUM(o[1755]) );
  FADDER \add_42/U1_1756  ( .CIN(sreg[1756]), .IN0(n2340), .IN1(
        \add_42/carry[1756] ), .COUT(\add_42/carry[1757] ), .SUM(o[1756]) );
  FADDER \add_42/U1_1757  ( .CIN(sreg[1757]), .IN0(n2339), .IN1(
        \add_42/carry[1757] ), .COUT(\add_42/carry[1758] ), .SUM(o[1757]) );
  FADDER \add_42/U1_1758  ( .CIN(sreg[1758]), .IN0(n2338), .IN1(
        \add_42/carry[1758] ), .COUT(\add_42/carry[1759] ), .SUM(o[1758]) );
  FADDER \add_42/U1_1759  ( .CIN(sreg[1759]), .IN0(n2337), .IN1(
        \add_42/carry[1759] ), .COUT(\add_42/carry[1760] ), .SUM(o[1759]) );
  FADDER \add_42/U1_1760  ( .CIN(sreg[1760]), .IN0(n2336), .IN1(
        \add_42/carry[1760] ), .COUT(\add_42/carry[1761] ), .SUM(o[1760]) );
  FADDER \add_42/U1_1761  ( .CIN(sreg[1761]), .IN0(n2335), .IN1(
        \add_42/carry[1761] ), .COUT(\add_42/carry[1762] ), .SUM(o[1761]) );
  FADDER \add_42/U1_1762  ( .CIN(sreg[1762]), .IN0(n2334), .IN1(
        \add_42/carry[1762] ), .COUT(\add_42/carry[1763] ), .SUM(o[1762]) );
  FADDER \add_42/U1_1763  ( .CIN(sreg[1763]), .IN0(n2333), .IN1(
        \add_42/carry[1763] ), .COUT(\add_42/carry[1764] ), .SUM(o[1763]) );
  FADDER \add_42/U1_1764  ( .CIN(sreg[1764]), .IN0(n2332), .IN1(
        \add_42/carry[1764] ), .COUT(\add_42/carry[1765] ), .SUM(o[1764]) );
  FADDER \add_42/U1_1765  ( .CIN(sreg[1765]), .IN0(n2331), .IN1(
        \add_42/carry[1765] ), .COUT(\add_42/carry[1766] ), .SUM(o[1765]) );
  FADDER \add_42/U1_1766  ( .CIN(sreg[1766]), .IN0(n2330), .IN1(
        \add_42/carry[1766] ), .COUT(\add_42/carry[1767] ), .SUM(o[1766]) );
  FADDER \add_42/U1_1767  ( .CIN(sreg[1767]), .IN0(n2329), .IN1(
        \add_42/carry[1767] ), .COUT(\add_42/carry[1768] ), .SUM(o[1767]) );
  FADDER \add_42/U1_1768  ( .CIN(sreg[1768]), .IN0(n2328), .IN1(
        \add_42/carry[1768] ), .COUT(\add_42/carry[1769] ), .SUM(o[1768]) );
  FADDER \add_42/U1_1769  ( .CIN(sreg[1769]), .IN0(n2327), .IN1(
        \add_42/carry[1769] ), .COUT(\add_42/carry[1770] ), .SUM(o[1769]) );
  FADDER \add_42/U1_1770  ( .CIN(sreg[1770]), .IN0(n2326), .IN1(
        \add_42/carry[1770] ), .COUT(\add_42/carry[1771] ), .SUM(o[1770]) );
  FADDER \add_42/U1_1771  ( .CIN(sreg[1771]), .IN0(n2325), .IN1(
        \add_42/carry[1771] ), .COUT(\add_42/carry[1772] ), .SUM(o[1771]) );
  FADDER \add_42/U1_1772  ( .CIN(sreg[1772]), .IN0(n2324), .IN1(
        \add_42/carry[1772] ), .COUT(\add_42/carry[1773] ), .SUM(o[1772]) );
  FADDER \add_42/U1_1773  ( .CIN(sreg[1773]), .IN0(n2323), .IN1(
        \add_42/carry[1773] ), .COUT(\add_42/carry[1774] ), .SUM(o[1773]) );
  FADDER \add_42/U1_1774  ( .CIN(sreg[1774]), .IN0(n2322), .IN1(
        \add_42/carry[1774] ), .COUT(\add_42/carry[1775] ), .SUM(o[1774]) );
  FADDER \add_42/U1_1775  ( .CIN(sreg[1775]), .IN0(n2321), .IN1(
        \add_42/carry[1775] ), .COUT(\add_42/carry[1776] ), .SUM(o[1775]) );
  FADDER \add_42/U1_1776  ( .CIN(sreg[1776]), .IN0(n2320), .IN1(
        \add_42/carry[1776] ), .COUT(\add_42/carry[1777] ), .SUM(o[1776]) );
  FADDER \add_42/U1_1777  ( .CIN(sreg[1777]), .IN0(n2319), .IN1(
        \add_42/carry[1777] ), .COUT(\add_42/carry[1778] ), .SUM(o[1777]) );
  FADDER \add_42/U1_1778  ( .CIN(sreg[1778]), .IN0(n2318), .IN1(
        \add_42/carry[1778] ), .COUT(\add_42/carry[1779] ), .SUM(o[1778]) );
  FADDER \add_42/U1_1779  ( .CIN(sreg[1779]), .IN0(n2317), .IN1(
        \add_42/carry[1779] ), .COUT(\add_42/carry[1780] ), .SUM(o[1779]) );
  FADDER \add_42/U1_1780  ( .CIN(sreg[1780]), .IN0(n2316), .IN1(
        \add_42/carry[1780] ), .COUT(\add_42/carry[1781] ), .SUM(o[1780]) );
  FADDER \add_42/U1_1781  ( .CIN(sreg[1781]), .IN0(n2315), .IN1(
        \add_42/carry[1781] ), .COUT(\add_42/carry[1782] ), .SUM(o[1781]) );
  FADDER \add_42/U1_1782  ( .CIN(sreg[1782]), .IN0(n2314), .IN1(
        \add_42/carry[1782] ), .COUT(\add_42/carry[1783] ), .SUM(o[1782]) );
  FADDER \add_42/U1_1783  ( .CIN(sreg[1783]), .IN0(n2313), .IN1(
        \add_42/carry[1783] ), .COUT(\add_42/carry[1784] ), .SUM(o[1783]) );
  FADDER \add_42/U1_1784  ( .CIN(sreg[1784]), .IN0(n2312), .IN1(
        \add_42/carry[1784] ), .COUT(\add_42/carry[1785] ), .SUM(o[1784]) );
  FADDER \add_42/U1_1785  ( .CIN(sreg[1785]), .IN0(n2311), .IN1(
        \add_42/carry[1785] ), .COUT(\add_42/carry[1786] ), .SUM(o[1785]) );
  FADDER \add_42/U1_1786  ( .CIN(sreg[1786]), .IN0(n2310), .IN1(
        \add_42/carry[1786] ), .COUT(\add_42/carry[1787] ), .SUM(o[1786]) );
  FADDER \add_42/U1_1787  ( .CIN(sreg[1787]), .IN0(n2309), .IN1(
        \add_42/carry[1787] ), .COUT(\add_42/carry[1788] ), .SUM(o[1787]) );
  FADDER \add_42/U1_1788  ( .CIN(sreg[1788]), .IN0(n2308), .IN1(
        \add_42/carry[1788] ), .COUT(\add_42/carry[1789] ), .SUM(o[1788]) );
  FADDER \add_42/U1_1789  ( .CIN(sreg[1789]), .IN0(n2307), .IN1(
        \add_42/carry[1789] ), .COUT(\add_42/carry[1790] ), .SUM(o[1789]) );
  FADDER \add_42/U1_1790  ( .CIN(sreg[1790]), .IN0(n2306), .IN1(
        \add_42/carry[1790] ), .COUT(\add_42/carry[1791] ), .SUM(o[1790]) );
  FADDER \add_42/U1_1791  ( .CIN(sreg[1791]), .IN0(n2305), .IN1(
        \add_42/carry[1791] ), .COUT(\add_42/carry[1792] ), .SUM(o[1791]) );
  FADDER \add_42/U1_1792  ( .CIN(sreg[1792]), .IN0(n2304), .IN1(
        \add_42/carry[1792] ), .COUT(\add_42/carry[1793] ), .SUM(o[1792]) );
  FADDER \add_42/U1_1793  ( .CIN(sreg[1793]), .IN0(n2303), .IN1(
        \add_42/carry[1793] ), .COUT(\add_42/carry[1794] ), .SUM(o[1793]) );
  FADDER \add_42/U1_1794  ( .CIN(sreg[1794]), .IN0(n2302), .IN1(
        \add_42/carry[1794] ), .COUT(\add_42/carry[1795] ), .SUM(o[1794]) );
  FADDER \add_42/U1_1795  ( .CIN(sreg[1795]), .IN0(n2301), .IN1(
        \add_42/carry[1795] ), .COUT(\add_42/carry[1796] ), .SUM(o[1795]) );
  FADDER \add_42/U1_1796  ( .CIN(sreg[1796]), .IN0(n2300), .IN1(
        \add_42/carry[1796] ), .COUT(\add_42/carry[1797] ), .SUM(o[1796]) );
  FADDER \add_42/U1_1797  ( .CIN(sreg[1797]), .IN0(n2299), .IN1(
        \add_42/carry[1797] ), .COUT(\add_42/carry[1798] ), .SUM(o[1797]) );
  FADDER \add_42/U1_1798  ( .CIN(sreg[1798]), .IN0(n2298), .IN1(
        \add_42/carry[1798] ), .COUT(\add_42/carry[1799] ), .SUM(o[1798]) );
  FADDER \add_42/U1_1799  ( .CIN(sreg[1799]), .IN0(n2297), .IN1(
        \add_42/carry[1799] ), .COUT(\add_42/carry[1800] ), .SUM(o[1799]) );
  FADDER \add_42/U1_1800  ( .CIN(sreg[1800]), .IN0(n2296), .IN1(
        \add_42/carry[1800] ), .COUT(\add_42/carry[1801] ), .SUM(o[1800]) );
  FADDER \add_42/U1_1801  ( .CIN(sreg[1801]), .IN0(n2295), .IN1(
        \add_42/carry[1801] ), .COUT(\add_42/carry[1802] ), .SUM(o[1801]) );
  FADDER \add_42/U1_1802  ( .CIN(sreg[1802]), .IN0(n2294), .IN1(
        \add_42/carry[1802] ), .COUT(\add_42/carry[1803] ), .SUM(o[1802]) );
  FADDER \add_42/U1_1803  ( .CIN(sreg[1803]), .IN0(n2293), .IN1(
        \add_42/carry[1803] ), .COUT(\add_42/carry[1804] ), .SUM(o[1803]) );
  FADDER \add_42/U1_1804  ( .CIN(sreg[1804]), .IN0(n2292), .IN1(
        \add_42/carry[1804] ), .COUT(\add_42/carry[1805] ), .SUM(o[1804]) );
  FADDER \add_42/U1_1805  ( .CIN(sreg[1805]), .IN0(n2291), .IN1(
        \add_42/carry[1805] ), .COUT(\add_42/carry[1806] ), .SUM(o[1805]) );
  FADDER \add_42/U1_1806  ( .CIN(sreg[1806]), .IN0(n2290), .IN1(
        \add_42/carry[1806] ), .COUT(\add_42/carry[1807] ), .SUM(o[1806]) );
  FADDER \add_42/U1_1807  ( .CIN(sreg[1807]), .IN0(n2289), .IN1(
        \add_42/carry[1807] ), .COUT(\add_42/carry[1808] ), .SUM(o[1807]) );
  FADDER \add_42/U1_1808  ( .CIN(sreg[1808]), .IN0(n2288), .IN1(
        \add_42/carry[1808] ), .COUT(\add_42/carry[1809] ), .SUM(o[1808]) );
  FADDER \add_42/U1_1809  ( .CIN(sreg[1809]), .IN0(n2287), .IN1(
        \add_42/carry[1809] ), .COUT(\add_42/carry[1810] ), .SUM(o[1809]) );
  FADDER \add_42/U1_1810  ( .CIN(sreg[1810]), .IN0(n2286), .IN1(
        \add_42/carry[1810] ), .COUT(\add_42/carry[1811] ), .SUM(o[1810]) );
  FADDER \add_42/U1_1811  ( .CIN(sreg[1811]), .IN0(n2285), .IN1(
        \add_42/carry[1811] ), .COUT(\add_42/carry[1812] ), .SUM(o[1811]) );
  FADDER \add_42/U1_1812  ( .CIN(sreg[1812]), .IN0(n2284), .IN1(
        \add_42/carry[1812] ), .COUT(\add_42/carry[1813] ), .SUM(o[1812]) );
  FADDER \add_42/U1_1813  ( .CIN(sreg[1813]), .IN0(n2283), .IN1(
        \add_42/carry[1813] ), .COUT(\add_42/carry[1814] ), .SUM(o[1813]) );
  FADDER \add_42/U1_1814  ( .CIN(sreg[1814]), .IN0(n2282), .IN1(
        \add_42/carry[1814] ), .COUT(\add_42/carry[1815] ), .SUM(o[1814]) );
  FADDER \add_42/U1_1815  ( .CIN(sreg[1815]), .IN0(n2281), .IN1(
        \add_42/carry[1815] ), .COUT(\add_42/carry[1816] ), .SUM(o[1815]) );
  FADDER \add_42/U1_1816  ( .CIN(sreg[1816]), .IN0(n2280), .IN1(
        \add_42/carry[1816] ), .COUT(\add_42/carry[1817] ), .SUM(o[1816]) );
  FADDER \add_42/U1_1817  ( .CIN(sreg[1817]), .IN0(n2279), .IN1(
        \add_42/carry[1817] ), .COUT(\add_42/carry[1818] ), .SUM(o[1817]) );
  FADDER \add_42/U1_1818  ( .CIN(sreg[1818]), .IN0(n2278), .IN1(
        \add_42/carry[1818] ), .COUT(\add_42/carry[1819] ), .SUM(o[1818]) );
  FADDER \add_42/U1_1819  ( .CIN(sreg[1819]), .IN0(n2277), .IN1(
        \add_42/carry[1819] ), .COUT(\add_42/carry[1820] ), .SUM(o[1819]) );
  FADDER \add_42/U1_1820  ( .CIN(sreg[1820]), .IN0(n2276), .IN1(
        \add_42/carry[1820] ), .COUT(\add_42/carry[1821] ), .SUM(o[1820]) );
  FADDER \add_42/U1_1821  ( .CIN(sreg[1821]), .IN0(n2275), .IN1(
        \add_42/carry[1821] ), .COUT(\add_42/carry[1822] ), .SUM(o[1821]) );
  FADDER \add_42/U1_1822  ( .CIN(sreg[1822]), .IN0(n2274), .IN1(
        \add_42/carry[1822] ), .COUT(\add_42/carry[1823] ), .SUM(o[1822]) );
  FADDER \add_42/U1_1823  ( .CIN(sreg[1823]), .IN0(n2273), .IN1(
        \add_42/carry[1823] ), .COUT(\add_42/carry[1824] ), .SUM(o[1823]) );
  FADDER \add_42/U1_1824  ( .CIN(sreg[1824]), .IN0(n2272), .IN1(
        \add_42/carry[1824] ), .COUT(\add_42/carry[1825] ), .SUM(o[1824]) );
  FADDER \add_42/U1_1825  ( .CIN(sreg[1825]), .IN0(n2271), .IN1(
        \add_42/carry[1825] ), .COUT(\add_42/carry[1826] ), .SUM(o[1825]) );
  FADDER \add_42/U1_1826  ( .CIN(sreg[1826]), .IN0(n2270), .IN1(
        \add_42/carry[1826] ), .COUT(\add_42/carry[1827] ), .SUM(o[1826]) );
  FADDER \add_42/U1_1827  ( .CIN(sreg[1827]), .IN0(n2269), .IN1(
        \add_42/carry[1827] ), .COUT(\add_42/carry[1828] ), .SUM(o[1827]) );
  FADDER \add_42/U1_1828  ( .CIN(sreg[1828]), .IN0(n2268), .IN1(
        \add_42/carry[1828] ), .COUT(\add_42/carry[1829] ), .SUM(o[1828]) );
  FADDER \add_42/U1_1829  ( .CIN(sreg[1829]), .IN0(n2267), .IN1(
        \add_42/carry[1829] ), .COUT(\add_42/carry[1830] ), .SUM(o[1829]) );
  FADDER \add_42/U1_1830  ( .CIN(sreg[1830]), .IN0(n2266), .IN1(
        \add_42/carry[1830] ), .COUT(\add_42/carry[1831] ), .SUM(o[1830]) );
  FADDER \add_42/U1_1831  ( .CIN(sreg[1831]), .IN0(n2265), .IN1(
        \add_42/carry[1831] ), .COUT(\add_42/carry[1832] ), .SUM(o[1831]) );
  FADDER \add_42/U1_1832  ( .CIN(sreg[1832]), .IN0(n2264), .IN1(
        \add_42/carry[1832] ), .COUT(\add_42/carry[1833] ), .SUM(o[1832]) );
  FADDER \add_42/U1_1833  ( .CIN(sreg[1833]), .IN0(n2263), .IN1(
        \add_42/carry[1833] ), .COUT(\add_42/carry[1834] ), .SUM(o[1833]) );
  FADDER \add_42/U1_1834  ( .CIN(sreg[1834]), .IN0(n2262), .IN1(
        \add_42/carry[1834] ), .COUT(\add_42/carry[1835] ), .SUM(o[1834]) );
  FADDER \add_42/U1_1835  ( .CIN(sreg[1835]), .IN0(n2261), .IN1(
        \add_42/carry[1835] ), .COUT(\add_42/carry[1836] ), .SUM(o[1835]) );
  FADDER \add_42/U1_1836  ( .CIN(sreg[1836]), .IN0(n2260), .IN1(
        \add_42/carry[1836] ), .COUT(\add_42/carry[1837] ), .SUM(o[1836]) );
  FADDER \add_42/U1_1837  ( .CIN(sreg[1837]), .IN0(n2259), .IN1(
        \add_42/carry[1837] ), .COUT(\add_42/carry[1838] ), .SUM(o[1837]) );
  FADDER \add_42/U1_1838  ( .CIN(sreg[1838]), .IN0(n2258), .IN1(
        \add_42/carry[1838] ), .COUT(\add_42/carry[1839] ), .SUM(o[1838]) );
  FADDER \add_42/U1_1839  ( .CIN(sreg[1839]), .IN0(n2257), .IN1(
        \add_42/carry[1839] ), .COUT(\add_42/carry[1840] ), .SUM(o[1839]) );
  FADDER \add_42/U1_1840  ( .CIN(sreg[1840]), .IN0(n2256), .IN1(
        \add_42/carry[1840] ), .COUT(\add_42/carry[1841] ), .SUM(o[1840]) );
  FADDER \add_42/U1_1841  ( .CIN(sreg[1841]), .IN0(n2255), .IN1(
        \add_42/carry[1841] ), .COUT(\add_42/carry[1842] ), .SUM(o[1841]) );
  FADDER \add_42/U1_1842  ( .CIN(sreg[1842]), .IN0(n2254), .IN1(
        \add_42/carry[1842] ), .COUT(\add_42/carry[1843] ), .SUM(o[1842]) );
  FADDER \add_42/U1_1843  ( .CIN(sreg[1843]), .IN0(n2253), .IN1(
        \add_42/carry[1843] ), .COUT(\add_42/carry[1844] ), .SUM(o[1843]) );
  FADDER \add_42/U1_1844  ( .CIN(sreg[1844]), .IN0(n2252), .IN1(
        \add_42/carry[1844] ), .COUT(\add_42/carry[1845] ), .SUM(o[1844]) );
  FADDER \add_42/U1_1845  ( .CIN(sreg[1845]), .IN0(n2251), .IN1(
        \add_42/carry[1845] ), .COUT(\add_42/carry[1846] ), .SUM(o[1845]) );
  FADDER \add_42/U1_1846  ( .CIN(sreg[1846]), .IN0(n2250), .IN1(
        \add_42/carry[1846] ), .COUT(\add_42/carry[1847] ), .SUM(o[1846]) );
  FADDER \add_42/U1_1847  ( .CIN(sreg[1847]), .IN0(n2249), .IN1(
        \add_42/carry[1847] ), .COUT(\add_42/carry[1848] ), .SUM(o[1847]) );
  FADDER \add_42/U1_1848  ( .CIN(sreg[1848]), .IN0(n2248), .IN1(
        \add_42/carry[1848] ), .COUT(\add_42/carry[1849] ), .SUM(o[1848]) );
  FADDER \add_42/U1_1849  ( .CIN(sreg[1849]), .IN0(n2247), .IN1(
        \add_42/carry[1849] ), .COUT(\add_42/carry[1850] ), .SUM(o[1849]) );
  FADDER \add_42/U1_1850  ( .CIN(sreg[1850]), .IN0(n2246), .IN1(
        \add_42/carry[1850] ), .COUT(\add_42/carry[1851] ), .SUM(o[1850]) );
  FADDER \add_42/U1_1851  ( .CIN(sreg[1851]), .IN0(n2245), .IN1(
        \add_42/carry[1851] ), .COUT(\add_42/carry[1852] ), .SUM(o[1851]) );
  FADDER \add_42/U1_1852  ( .CIN(sreg[1852]), .IN0(n2244), .IN1(
        \add_42/carry[1852] ), .COUT(\add_42/carry[1853] ), .SUM(o[1852]) );
  FADDER \add_42/U1_1853  ( .CIN(sreg[1853]), .IN0(n2243), .IN1(
        \add_42/carry[1853] ), .COUT(\add_42/carry[1854] ), .SUM(o[1853]) );
  FADDER \add_42/U1_1854  ( .CIN(sreg[1854]), .IN0(n2242), .IN1(
        \add_42/carry[1854] ), .COUT(\add_42/carry[1855] ), .SUM(o[1854]) );
  FADDER \add_42/U1_1855  ( .CIN(sreg[1855]), .IN0(n2241), .IN1(
        \add_42/carry[1855] ), .COUT(\add_42/carry[1856] ), .SUM(o[1855]) );
  FADDER \add_42/U1_1856  ( .CIN(sreg[1856]), .IN0(n2240), .IN1(
        \add_42/carry[1856] ), .COUT(\add_42/carry[1857] ), .SUM(o[1856]) );
  FADDER \add_42/U1_1857  ( .CIN(sreg[1857]), .IN0(n2239), .IN1(
        \add_42/carry[1857] ), .COUT(\add_42/carry[1858] ), .SUM(o[1857]) );
  FADDER \add_42/U1_1858  ( .CIN(sreg[1858]), .IN0(n2238), .IN1(
        \add_42/carry[1858] ), .COUT(\add_42/carry[1859] ), .SUM(o[1858]) );
  FADDER \add_42/U1_1859  ( .CIN(sreg[1859]), .IN0(n2237), .IN1(
        \add_42/carry[1859] ), .COUT(\add_42/carry[1860] ), .SUM(o[1859]) );
  FADDER \add_42/U1_1860  ( .CIN(sreg[1860]), .IN0(n2236), .IN1(
        \add_42/carry[1860] ), .COUT(\add_42/carry[1861] ), .SUM(o[1860]) );
  FADDER \add_42/U1_1861  ( .CIN(sreg[1861]), .IN0(n2235), .IN1(
        \add_42/carry[1861] ), .COUT(\add_42/carry[1862] ), .SUM(o[1861]) );
  FADDER \add_42/U1_1862  ( .CIN(sreg[1862]), .IN0(n2234), .IN1(
        \add_42/carry[1862] ), .COUT(\add_42/carry[1863] ), .SUM(o[1862]) );
  FADDER \add_42/U1_1863  ( .CIN(sreg[1863]), .IN0(n2233), .IN1(
        \add_42/carry[1863] ), .COUT(\add_42/carry[1864] ), .SUM(o[1863]) );
  FADDER \add_42/U1_1864  ( .CIN(sreg[1864]), .IN0(n2232), .IN1(
        \add_42/carry[1864] ), .COUT(\add_42/carry[1865] ), .SUM(o[1864]) );
  FADDER \add_42/U1_1865  ( .CIN(sreg[1865]), .IN0(n2231), .IN1(
        \add_42/carry[1865] ), .COUT(\add_42/carry[1866] ), .SUM(o[1865]) );
  FADDER \add_42/U1_1866  ( .CIN(sreg[1866]), .IN0(n2230), .IN1(
        \add_42/carry[1866] ), .COUT(\add_42/carry[1867] ), .SUM(o[1866]) );
  FADDER \add_42/U1_1867  ( .CIN(sreg[1867]), .IN0(n2229), .IN1(
        \add_42/carry[1867] ), .COUT(\add_42/carry[1868] ), .SUM(o[1867]) );
  FADDER \add_42/U1_1868  ( .CIN(sreg[1868]), .IN0(n2228), .IN1(
        \add_42/carry[1868] ), .COUT(\add_42/carry[1869] ), .SUM(o[1868]) );
  FADDER \add_42/U1_1869  ( .CIN(sreg[1869]), .IN0(n2227), .IN1(
        \add_42/carry[1869] ), .COUT(\add_42/carry[1870] ), .SUM(o[1869]) );
  FADDER \add_42/U1_1870  ( .CIN(sreg[1870]), .IN0(n2226), .IN1(
        \add_42/carry[1870] ), .COUT(\add_42/carry[1871] ), .SUM(o[1870]) );
  FADDER \add_42/U1_1871  ( .CIN(sreg[1871]), .IN0(n2225), .IN1(
        \add_42/carry[1871] ), .COUT(\add_42/carry[1872] ), .SUM(o[1871]) );
  FADDER \add_42/U1_1872  ( .CIN(sreg[1872]), .IN0(n2224), .IN1(
        \add_42/carry[1872] ), .COUT(\add_42/carry[1873] ), .SUM(o[1872]) );
  FADDER \add_42/U1_1873  ( .CIN(sreg[1873]), .IN0(n2223), .IN1(
        \add_42/carry[1873] ), .COUT(\add_42/carry[1874] ), .SUM(o[1873]) );
  FADDER \add_42/U1_1874  ( .CIN(sreg[1874]), .IN0(n2222), .IN1(
        \add_42/carry[1874] ), .COUT(\add_42/carry[1875] ), .SUM(o[1874]) );
  FADDER \add_42/U1_1875  ( .CIN(sreg[1875]), .IN0(n2221), .IN1(
        \add_42/carry[1875] ), .COUT(\add_42/carry[1876] ), .SUM(o[1875]) );
  FADDER \add_42/U1_1876  ( .CIN(sreg[1876]), .IN0(n2220), .IN1(
        \add_42/carry[1876] ), .COUT(\add_42/carry[1877] ), .SUM(o[1876]) );
  FADDER \add_42/U1_1877  ( .CIN(sreg[1877]), .IN0(n2219), .IN1(
        \add_42/carry[1877] ), .COUT(\add_42/carry[1878] ), .SUM(o[1877]) );
  FADDER \add_42/U1_1878  ( .CIN(sreg[1878]), .IN0(n2218), .IN1(
        \add_42/carry[1878] ), .COUT(\add_42/carry[1879] ), .SUM(o[1878]) );
  FADDER \add_42/U1_1879  ( .CIN(sreg[1879]), .IN0(n2217), .IN1(
        \add_42/carry[1879] ), .COUT(\add_42/carry[1880] ), .SUM(o[1879]) );
  FADDER \add_42/U1_1880  ( .CIN(sreg[1880]), .IN0(n2216), .IN1(
        \add_42/carry[1880] ), .COUT(\add_42/carry[1881] ), .SUM(o[1880]) );
  FADDER \add_42/U1_1881  ( .CIN(sreg[1881]), .IN0(n2215), .IN1(
        \add_42/carry[1881] ), .COUT(\add_42/carry[1882] ), .SUM(o[1881]) );
  FADDER \add_42/U1_1882  ( .CIN(sreg[1882]), .IN0(n2214), .IN1(
        \add_42/carry[1882] ), .COUT(\add_42/carry[1883] ), .SUM(o[1882]) );
  FADDER \add_42/U1_1883  ( .CIN(sreg[1883]), .IN0(n2213), .IN1(
        \add_42/carry[1883] ), .COUT(\add_42/carry[1884] ), .SUM(o[1883]) );
  FADDER \add_42/U1_1884  ( .CIN(sreg[1884]), .IN0(n2212), .IN1(
        \add_42/carry[1884] ), .COUT(\add_42/carry[1885] ), .SUM(o[1884]) );
  FADDER \add_42/U1_1885  ( .CIN(sreg[1885]), .IN0(n2211), .IN1(
        \add_42/carry[1885] ), .COUT(\add_42/carry[1886] ), .SUM(o[1885]) );
  FADDER \add_42/U1_1886  ( .CIN(sreg[1886]), .IN0(n2210), .IN1(
        \add_42/carry[1886] ), .COUT(\add_42/carry[1887] ), .SUM(o[1886]) );
  FADDER \add_42/U1_1887  ( .CIN(sreg[1887]), .IN0(n2209), .IN1(
        \add_42/carry[1887] ), .COUT(\add_42/carry[1888] ), .SUM(o[1887]) );
  FADDER \add_42/U1_1888  ( .CIN(sreg[1888]), .IN0(n2208), .IN1(
        \add_42/carry[1888] ), .COUT(\add_42/carry[1889] ), .SUM(o[1888]) );
  FADDER \add_42/U1_1889  ( .CIN(sreg[1889]), .IN0(n2207), .IN1(
        \add_42/carry[1889] ), .COUT(\add_42/carry[1890] ), .SUM(o[1889]) );
  FADDER \add_42/U1_1890  ( .CIN(sreg[1890]), .IN0(n2206), .IN1(
        \add_42/carry[1890] ), .COUT(\add_42/carry[1891] ), .SUM(o[1890]) );
  FADDER \add_42/U1_1891  ( .CIN(sreg[1891]), .IN0(n2205), .IN1(
        \add_42/carry[1891] ), .COUT(\add_42/carry[1892] ), .SUM(o[1891]) );
  FADDER \add_42/U1_1892  ( .CIN(sreg[1892]), .IN0(n2204), .IN1(
        \add_42/carry[1892] ), .COUT(\add_42/carry[1893] ), .SUM(o[1892]) );
  FADDER \add_42/U1_1893  ( .CIN(sreg[1893]), .IN0(n2203), .IN1(
        \add_42/carry[1893] ), .COUT(\add_42/carry[1894] ), .SUM(o[1893]) );
  FADDER \add_42/U1_1894  ( .CIN(sreg[1894]), .IN0(n2202), .IN1(
        \add_42/carry[1894] ), .COUT(\add_42/carry[1895] ), .SUM(o[1894]) );
  FADDER \add_42/U1_1895  ( .CIN(sreg[1895]), .IN0(n2201), .IN1(
        \add_42/carry[1895] ), .COUT(\add_42/carry[1896] ), .SUM(o[1895]) );
  FADDER \add_42/U1_1896  ( .CIN(sreg[1896]), .IN0(n2200), .IN1(
        \add_42/carry[1896] ), .COUT(\add_42/carry[1897] ), .SUM(o[1896]) );
  FADDER \add_42/U1_1897  ( .CIN(sreg[1897]), .IN0(n2199), .IN1(
        \add_42/carry[1897] ), .COUT(\add_42/carry[1898] ), .SUM(o[1897]) );
  FADDER \add_42/U1_1898  ( .CIN(sreg[1898]), .IN0(n2198), .IN1(
        \add_42/carry[1898] ), .COUT(\add_42/carry[1899] ), .SUM(o[1898]) );
  FADDER \add_42/U1_1899  ( .CIN(sreg[1899]), .IN0(n2197), .IN1(
        \add_42/carry[1899] ), .COUT(\add_42/carry[1900] ), .SUM(o[1899]) );
  FADDER \add_42/U1_1900  ( .CIN(sreg[1900]), .IN0(n2196), .IN1(
        \add_42/carry[1900] ), .COUT(\add_42/carry[1901] ), .SUM(o[1900]) );
  FADDER \add_42/U1_1901  ( .CIN(sreg[1901]), .IN0(n2195), .IN1(
        \add_42/carry[1901] ), .COUT(\add_42/carry[1902] ), .SUM(o[1901]) );
  FADDER \add_42/U1_1902  ( .CIN(sreg[1902]), .IN0(n2194), .IN1(
        \add_42/carry[1902] ), .COUT(\add_42/carry[1903] ), .SUM(o[1902]) );
  FADDER \add_42/U1_1903  ( .CIN(sreg[1903]), .IN0(n2193), .IN1(
        \add_42/carry[1903] ), .COUT(\add_42/carry[1904] ), .SUM(o[1903]) );
  FADDER \add_42/U1_1904  ( .CIN(sreg[1904]), .IN0(n2192), .IN1(
        \add_42/carry[1904] ), .COUT(\add_42/carry[1905] ), .SUM(o[1904]) );
  FADDER \add_42/U1_1905  ( .CIN(sreg[1905]), .IN0(n2191), .IN1(
        \add_42/carry[1905] ), .COUT(\add_42/carry[1906] ), .SUM(o[1905]) );
  FADDER \add_42/U1_1906  ( .CIN(sreg[1906]), .IN0(n2190), .IN1(
        \add_42/carry[1906] ), .COUT(\add_42/carry[1907] ), .SUM(o[1906]) );
  FADDER \add_42/U1_1907  ( .CIN(sreg[1907]), .IN0(n2189), .IN1(
        \add_42/carry[1907] ), .COUT(\add_42/carry[1908] ), .SUM(o[1907]) );
  FADDER \add_42/U1_1908  ( .CIN(sreg[1908]), .IN0(n2188), .IN1(
        \add_42/carry[1908] ), .COUT(\add_42/carry[1909] ), .SUM(o[1908]) );
  FADDER \add_42/U1_1909  ( .CIN(sreg[1909]), .IN0(n2187), .IN1(
        \add_42/carry[1909] ), .COUT(\add_42/carry[1910] ), .SUM(o[1909]) );
  FADDER \add_42/U1_1910  ( .CIN(sreg[1910]), .IN0(n2186), .IN1(
        \add_42/carry[1910] ), .COUT(\add_42/carry[1911] ), .SUM(o[1910]) );
  FADDER \add_42/U1_1911  ( .CIN(sreg[1911]), .IN0(n2185), .IN1(
        \add_42/carry[1911] ), .COUT(\add_42/carry[1912] ), .SUM(o[1911]) );
  FADDER \add_42/U1_1912  ( .CIN(sreg[1912]), .IN0(n2184), .IN1(
        \add_42/carry[1912] ), .COUT(\add_42/carry[1913] ), .SUM(o[1912]) );
  FADDER \add_42/U1_1913  ( .CIN(sreg[1913]), .IN0(n2183), .IN1(
        \add_42/carry[1913] ), .COUT(\add_42/carry[1914] ), .SUM(o[1913]) );
  FADDER \add_42/U1_1914  ( .CIN(sreg[1914]), .IN0(n2182), .IN1(
        \add_42/carry[1914] ), .COUT(\add_42/carry[1915] ), .SUM(o[1914]) );
  FADDER \add_42/U1_1915  ( .CIN(sreg[1915]), .IN0(n2181), .IN1(
        \add_42/carry[1915] ), .COUT(\add_42/carry[1916] ), .SUM(o[1915]) );
  FADDER \add_42/U1_1916  ( .CIN(sreg[1916]), .IN0(n2180), .IN1(
        \add_42/carry[1916] ), .COUT(\add_42/carry[1917] ), .SUM(o[1916]) );
  FADDER \add_42/U1_1917  ( .CIN(sreg[1917]), .IN0(n2179), .IN1(
        \add_42/carry[1917] ), .COUT(\add_42/carry[1918] ), .SUM(o[1917]) );
  FADDER \add_42/U1_1918  ( .CIN(sreg[1918]), .IN0(n2178), .IN1(
        \add_42/carry[1918] ), .COUT(\add_42/carry[1919] ), .SUM(o[1918]) );
  FADDER \add_42/U1_1919  ( .CIN(sreg[1919]), .IN0(n2177), .IN1(
        \add_42/carry[1919] ), .COUT(\add_42/carry[1920] ), .SUM(o[1919]) );
  FADDER \add_42/U1_1920  ( .CIN(sreg[1920]), .IN0(n2176), .IN1(
        \add_42/carry[1920] ), .COUT(\add_42/carry[1921] ), .SUM(o[1920]) );
  FADDER \add_42/U1_1921  ( .CIN(sreg[1921]), .IN0(n2175), .IN1(
        \add_42/carry[1921] ), .COUT(\add_42/carry[1922] ), .SUM(o[1921]) );
  FADDER \add_42/U1_1922  ( .CIN(sreg[1922]), .IN0(n2174), .IN1(
        \add_42/carry[1922] ), .COUT(\add_42/carry[1923] ), .SUM(o[1922]) );
  FADDER \add_42/U1_1923  ( .CIN(sreg[1923]), .IN0(n2173), .IN1(
        \add_42/carry[1923] ), .COUT(\add_42/carry[1924] ), .SUM(o[1923]) );
  FADDER \add_42/U1_1924  ( .CIN(sreg[1924]), .IN0(n2172), .IN1(
        \add_42/carry[1924] ), .COUT(\add_42/carry[1925] ), .SUM(o[1924]) );
  FADDER \add_42/U1_1925  ( .CIN(sreg[1925]), .IN0(n2171), .IN1(
        \add_42/carry[1925] ), .COUT(\add_42/carry[1926] ), .SUM(o[1925]) );
  FADDER \add_42/U1_1926  ( .CIN(sreg[1926]), .IN0(n2170), .IN1(
        \add_42/carry[1926] ), .COUT(\add_42/carry[1927] ), .SUM(o[1926]) );
  FADDER \add_42/U1_1927  ( .CIN(sreg[1927]), .IN0(n2169), .IN1(
        \add_42/carry[1927] ), .COUT(\add_42/carry[1928] ), .SUM(o[1927]) );
  FADDER \add_42/U1_1928  ( .CIN(sreg[1928]), .IN0(n2168), .IN1(
        \add_42/carry[1928] ), .COUT(\add_42/carry[1929] ), .SUM(o[1928]) );
  FADDER \add_42/U1_1929  ( .CIN(sreg[1929]), .IN0(n2167), .IN1(
        \add_42/carry[1929] ), .COUT(\add_42/carry[1930] ), .SUM(o[1929]) );
  FADDER \add_42/U1_1930  ( .CIN(sreg[1930]), .IN0(n2166), .IN1(
        \add_42/carry[1930] ), .COUT(\add_42/carry[1931] ), .SUM(o[1930]) );
  FADDER \add_42/U1_1931  ( .CIN(sreg[1931]), .IN0(n2165), .IN1(
        \add_42/carry[1931] ), .COUT(\add_42/carry[1932] ), .SUM(o[1931]) );
  FADDER \add_42/U1_1932  ( .CIN(sreg[1932]), .IN0(n2164), .IN1(
        \add_42/carry[1932] ), .COUT(\add_42/carry[1933] ), .SUM(o[1932]) );
  FADDER \add_42/U1_1933  ( .CIN(sreg[1933]), .IN0(n2163), .IN1(
        \add_42/carry[1933] ), .COUT(\add_42/carry[1934] ), .SUM(o[1933]) );
  FADDER \add_42/U1_1934  ( .CIN(sreg[1934]), .IN0(n2162), .IN1(
        \add_42/carry[1934] ), .COUT(\add_42/carry[1935] ), .SUM(o[1934]) );
  FADDER \add_42/U1_1935  ( .CIN(sreg[1935]), .IN0(n2161), .IN1(
        \add_42/carry[1935] ), .COUT(\add_42/carry[1936] ), .SUM(o[1935]) );
  FADDER \add_42/U1_1936  ( .CIN(sreg[1936]), .IN0(n2160), .IN1(
        \add_42/carry[1936] ), .COUT(\add_42/carry[1937] ), .SUM(o[1936]) );
  FADDER \add_42/U1_1937  ( .CIN(sreg[1937]), .IN0(n2159), .IN1(
        \add_42/carry[1937] ), .COUT(\add_42/carry[1938] ), .SUM(o[1937]) );
  FADDER \add_42/U1_1938  ( .CIN(sreg[1938]), .IN0(n2158), .IN1(
        \add_42/carry[1938] ), .COUT(\add_42/carry[1939] ), .SUM(o[1938]) );
  FADDER \add_42/U1_1939  ( .CIN(sreg[1939]), .IN0(n2157), .IN1(
        \add_42/carry[1939] ), .COUT(\add_42/carry[1940] ), .SUM(o[1939]) );
  FADDER \add_42/U1_1940  ( .CIN(sreg[1940]), .IN0(n2156), .IN1(
        \add_42/carry[1940] ), .COUT(\add_42/carry[1941] ), .SUM(o[1940]) );
  FADDER \add_42/U1_1941  ( .CIN(sreg[1941]), .IN0(n2155), .IN1(
        \add_42/carry[1941] ), .COUT(\add_42/carry[1942] ), .SUM(o[1941]) );
  FADDER \add_42/U1_1942  ( .CIN(sreg[1942]), .IN0(n2154), .IN1(
        \add_42/carry[1942] ), .COUT(\add_42/carry[1943] ), .SUM(o[1942]) );
  FADDER \add_42/U1_1943  ( .CIN(sreg[1943]), .IN0(n2153), .IN1(
        \add_42/carry[1943] ), .COUT(\add_42/carry[1944] ), .SUM(o[1943]) );
  FADDER \add_42/U1_1944  ( .CIN(sreg[1944]), .IN0(n2152), .IN1(
        \add_42/carry[1944] ), .COUT(\add_42/carry[1945] ), .SUM(o[1944]) );
  FADDER \add_42/U1_1945  ( .CIN(sreg[1945]), .IN0(n2151), .IN1(
        \add_42/carry[1945] ), .COUT(\add_42/carry[1946] ), .SUM(o[1945]) );
  FADDER \add_42/U1_1946  ( .CIN(sreg[1946]), .IN0(n2150), .IN1(
        \add_42/carry[1946] ), .COUT(\add_42/carry[1947] ), .SUM(o[1946]) );
  FADDER \add_42/U1_1947  ( .CIN(sreg[1947]), .IN0(n2149), .IN1(
        \add_42/carry[1947] ), .COUT(\add_42/carry[1948] ), .SUM(o[1947]) );
  FADDER \add_42/U1_1948  ( .CIN(sreg[1948]), .IN0(n2148), .IN1(
        \add_42/carry[1948] ), .COUT(\add_42/carry[1949] ), .SUM(o[1948]) );
  FADDER \add_42/U1_1949  ( .CIN(sreg[1949]), .IN0(n2147), .IN1(
        \add_42/carry[1949] ), .COUT(\add_42/carry[1950] ), .SUM(o[1949]) );
  FADDER \add_42/U1_1950  ( .CIN(sreg[1950]), .IN0(n2146), .IN1(
        \add_42/carry[1950] ), .COUT(\add_42/carry[1951] ), .SUM(o[1950]) );
  FADDER \add_42/U1_1951  ( .CIN(sreg[1951]), .IN0(n2145), .IN1(
        \add_42/carry[1951] ), .COUT(\add_42/carry[1952] ), .SUM(o[1951]) );
  FADDER \add_42/U1_1952  ( .CIN(sreg[1952]), .IN0(n2144), .IN1(
        \add_42/carry[1952] ), .COUT(\add_42/carry[1953] ), .SUM(o[1952]) );
  FADDER \add_42/U1_1953  ( .CIN(sreg[1953]), .IN0(n2143), .IN1(
        \add_42/carry[1953] ), .COUT(\add_42/carry[1954] ), .SUM(o[1953]) );
  FADDER \add_42/U1_1954  ( .CIN(sreg[1954]), .IN0(n2142), .IN1(
        \add_42/carry[1954] ), .COUT(\add_42/carry[1955] ), .SUM(o[1954]) );
  FADDER \add_42/U1_1955  ( .CIN(sreg[1955]), .IN0(n2141), .IN1(
        \add_42/carry[1955] ), .COUT(\add_42/carry[1956] ), .SUM(o[1955]) );
  FADDER \add_42/U1_1956  ( .CIN(sreg[1956]), .IN0(n2140), .IN1(
        \add_42/carry[1956] ), .COUT(\add_42/carry[1957] ), .SUM(o[1956]) );
  FADDER \add_42/U1_1957  ( .CIN(sreg[1957]), .IN0(n2139), .IN1(
        \add_42/carry[1957] ), .COUT(\add_42/carry[1958] ), .SUM(o[1957]) );
  FADDER \add_42/U1_1958  ( .CIN(sreg[1958]), .IN0(n2138), .IN1(
        \add_42/carry[1958] ), .COUT(\add_42/carry[1959] ), .SUM(o[1958]) );
  FADDER \add_42/U1_1959  ( .CIN(sreg[1959]), .IN0(n2137), .IN1(
        \add_42/carry[1959] ), .COUT(\add_42/carry[1960] ), .SUM(o[1959]) );
  FADDER \add_42/U1_1960  ( .CIN(sreg[1960]), .IN0(n2136), .IN1(
        \add_42/carry[1960] ), .COUT(\add_42/carry[1961] ), .SUM(o[1960]) );
  FADDER \add_42/U1_1961  ( .CIN(sreg[1961]), .IN0(n2135), .IN1(
        \add_42/carry[1961] ), .COUT(\add_42/carry[1962] ), .SUM(o[1961]) );
  FADDER \add_42/U1_1962  ( .CIN(sreg[1962]), .IN0(n2134), .IN1(
        \add_42/carry[1962] ), .COUT(\add_42/carry[1963] ), .SUM(o[1962]) );
  FADDER \add_42/U1_1963  ( .CIN(sreg[1963]), .IN0(n2133), .IN1(
        \add_42/carry[1963] ), .COUT(\add_42/carry[1964] ), .SUM(o[1963]) );
  FADDER \add_42/U1_1964  ( .CIN(sreg[1964]), .IN0(n2132), .IN1(
        \add_42/carry[1964] ), .COUT(\add_42/carry[1965] ), .SUM(o[1964]) );
  FADDER \add_42/U1_1965  ( .CIN(sreg[1965]), .IN0(n2131), .IN1(
        \add_42/carry[1965] ), .COUT(\add_42/carry[1966] ), .SUM(o[1965]) );
  FADDER \add_42/U1_1966  ( .CIN(sreg[1966]), .IN0(n2130), .IN1(
        \add_42/carry[1966] ), .COUT(\add_42/carry[1967] ), .SUM(o[1966]) );
  FADDER \add_42/U1_1967  ( .CIN(sreg[1967]), .IN0(n2129), .IN1(
        \add_42/carry[1967] ), .COUT(\add_42/carry[1968] ), .SUM(o[1967]) );
  FADDER \add_42/U1_1968  ( .CIN(sreg[1968]), .IN0(n2128), .IN1(
        \add_42/carry[1968] ), .COUT(\add_42/carry[1969] ), .SUM(o[1968]) );
  FADDER \add_42/U1_1969  ( .CIN(sreg[1969]), .IN0(n2127), .IN1(
        \add_42/carry[1969] ), .COUT(\add_42/carry[1970] ), .SUM(o[1969]) );
  FADDER \add_42/U1_1970  ( .CIN(sreg[1970]), .IN0(n2126), .IN1(
        \add_42/carry[1970] ), .COUT(\add_42/carry[1971] ), .SUM(o[1970]) );
  FADDER \add_42/U1_1971  ( .CIN(sreg[1971]), .IN0(n2125), .IN1(
        \add_42/carry[1971] ), .COUT(\add_42/carry[1972] ), .SUM(o[1971]) );
  FADDER \add_42/U1_1972  ( .CIN(sreg[1972]), .IN0(n2124), .IN1(
        \add_42/carry[1972] ), .COUT(\add_42/carry[1973] ), .SUM(o[1972]) );
  FADDER \add_42/U1_1973  ( .CIN(sreg[1973]), .IN0(n2123), .IN1(
        \add_42/carry[1973] ), .COUT(\add_42/carry[1974] ), .SUM(o[1973]) );
  FADDER \add_42/U1_1974  ( .CIN(sreg[1974]), .IN0(n2122), .IN1(
        \add_42/carry[1974] ), .COUT(\add_42/carry[1975] ), .SUM(o[1974]) );
  FADDER \add_42/U1_1975  ( .CIN(sreg[1975]), .IN0(n2121), .IN1(
        \add_42/carry[1975] ), .COUT(\add_42/carry[1976] ), .SUM(o[1975]) );
  FADDER \add_42/U1_1976  ( .CIN(sreg[1976]), .IN0(n2120), .IN1(
        \add_42/carry[1976] ), .COUT(\add_42/carry[1977] ), .SUM(o[1976]) );
  FADDER \add_42/U1_1977  ( .CIN(sreg[1977]), .IN0(n2119), .IN1(
        \add_42/carry[1977] ), .COUT(\add_42/carry[1978] ), .SUM(o[1977]) );
  FADDER \add_42/U1_1978  ( .CIN(sreg[1978]), .IN0(n2118), .IN1(
        \add_42/carry[1978] ), .COUT(\add_42/carry[1979] ), .SUM(o[1978]) );
  FADDER \add_42/U1_1979  ( .CIN(sreg[1979]), .IN0(n2117), .IN1(
        \add_42/carry[1979] ), .COUT(\add_42/carry[1980] ), .SUM(o[1979]) );
  FADDER \add_42/U1_1980  ( .CIN(sreg[1980]), .IN0(n2116), .IN1(
        \add_42/carry[1980] ), .COUT(\add_42/carry[1981] ), .SUM(o[1980]) );
  FADDER \add_42/U1_1981  ( .CIN(sreg[1981]), .IN0(n2115), .IN1(
        \add_42/carry[1981] ), .COUT(\add_42/carry[1982] ), .SUM(o[1981]) );
  FADDER \add_42/U1_1982  ( .CIN(sreg[1982]), .IN0(n2114), .IN1(
        \add_42/carry[1982] ), .COUT(\add_42/carry[1983] ), .SUM(o[1982]) );
  FADDER \add_42/U1_1983  ( .CIN(sreg[1983]), .IN0(n2113), .IN1(
        \add_42/carry[1983] ), .COUT(\add_42/carry[1984] ), .SUM(o[1983]) );
  FADDER \add_42/U1_1984  ( .CIN(sreg[1984]), .IN0(n2112), .IN1(
        \add_42/carry[1984] ), .COUT(\add_42/carry[1985] ), .SUM(o[1984]) );
  FADDER \add_42/U1_1985  ( .CIN(sreg[1985]), .IN0(n2111), .IN1(
        \add_42/carry[1985] ), .COUT(\add_42/carry[1986] ), .SUM(o[1985]) );
  FADDER \add_42/U1_1986  ( .CIN(sreg[1986]), .IN0(n2110), .IN1(
        \add_42/carry[1986] ), .COUT(\add_42/carry[1987] ), .SUM(o[1986]) );
  FADDER \add_42/U1_1987  ( .CIN(sreg[1987]), .IN0(n2109), .IN1(
        \add_42/carry[1987] ), .COUT(\add_42/carry[1988] ), .SUM(o[1987]) );
  FADDER \add_42/U1_1988  ( .CIN(sreg[1988]), .IN0(n2108), .IN1(
        \add_42/carry[1988] ), .COUT(\add_42/carry[1989] ), .SUM(o[1988]) );
  FADDER \add_42/U1_1989  ( .CIN(sreg[1989]), .IN0(n2107), .IN1(
        \add_42/carry[1989] ), .COUT(\add_42/carry[1990] ), .SUM(o[1989]) );
  FADDER \add_42/U1_1990  ( .CIN(sreg[1990]), .IN0(n2106), .IN1(
        \add_42/carry[1990] ), .COUT(\add_42/carry[1991] ), .SUM(o[1990]) );
  FADDER \add_42/U1_1991  ( .CIN(sreg[1991]), .IN0(n2105), .IN1(
        \add_42/carry[1991] ), .COUT(\add_42/carry[1992] ), .SUM(o[1991]) );
  FADDER \add_42/U1_1992  ( .CIN(sreg[1992]), .IN0(n2104), .IN1(
        \add_42/carry[1992] ), .COUT(\add_42/carry[1993] ), .SUM(o[1992]) );
  FADDER \add_42/U1_1993  ( .CIN(sreg[1993]), .IN0(n2103), .IN1(
        \add_42/carry[1993] ), .COUT(\add_42/carry[1994] ), .SUM(o[1993]) );
  FADDER \add_42/U1_1994  ( .CIN(sreg[1994]), .IN0(n2102), .IN1(
        \add_42/carry[1994] ), .COUT(\add_42/carry[1995] ), .SUM(o[1994]) );
  FADDER \add_42/U1_1995  ( .CIN(sreg[1995]), .IN0(n2101), .IN1(
        \add_42/carry[1995] ), .COUT(\add_42/carry[1996] ), .SUM(o[1995]) );
  FADDER \add_42/U1_1996  ( .CIN(sreg[1996]), .IN0(n2100), .IN1(
        \add_42/carry[1996] ), .COUT(\add_42/carry[1997] ), .SUM(o[1996]) );
  FADDER \add_42/U1_1997  ( .CIN(sreg[1997]), .IN0(n2099), .IN1(
        \add_42/carry[1997] ), .COUT(\add_42/carry[1998] ), .SUM(o[1997]) );
  FADDER \add_42/U1_1998  ( .CIN(sreg[1998]), .IN0(n2098), .IN1(
        \add_42/carry[1998] ), .COUT(\add_42/carry[1999] ), .SUM(o[1998]) );
  FADDER \add_42/U1_1999  ( .CIN(sreg[1999]), .IN0(n2097), .IN1(
        \add_42/carry[1999] ), .COUT(\add_42/carry[2000] ), .SUM(o[1999]) );
  FADDER \add_42/U1_2000  ( .CIN(sreg[2000]), .IN0(n2096), .IN1(
        \add_42/carry[2000] ), .COUT(\add_42/carry[2001] ), .SUM(o[2000]) );
  FADDER \add_42/U1_2001  ( .CIN(sreg[2001]), .IN0(n2095), .IN1(
        \add_42/carry[2001] ), .COUT(\add_42/carry[2002] ), .SUM(o[2001]) );
  FADDER \add_42/U1_2002  ( .CIN(sreg[2002]), .IN0(n2094), .IN1(
        \add_42/carry[2002] ), .COUT(\add_42/carry[2003] ), .SUM(o[2002]) );
  FADDER \add_42/U1_2003  ( .CIN(sreg[2003]), .IN0(n2093), .IN1(
        \add_42/carry[2003] ), .COUT(\add_42/carry[2004] ), .SUM(o[2003]) );
  FADDER \add_42/U1_2004  ( .CIN(sreg[2004]), .IN0(n2092), .IN1(
        \add_42/carry[2004] ), .COUT(\add_42/carry[2005] ), .SUM(o[2004]) );
  FADDER \add_42/U1_2005  ( .CIN(sreg[2005]), .IN0(n2091), .IN1(
        \add_42/carry[2005] ), .COUT(\add_42/carry[2006] ), .SUM(o[2005]) );
  FADDER \add_42/U1_2006  ( .CIN(sreg[2006]), .IN0(n2090), .IN1(
        \add_42/carry[2006] ), .COUT(\add_42/carry[2007] ), .SUM(o[2006]) );
  FADDER \add_42/U1_2007  ( .CIN(sreg[2007]), .IN0(n2089), .IN1(
        \add_42/carry[2007] ), .COUT(\add_42/carry[2008] ), .SUM(o[2007]) );
  FADDER \add_42/U1_2008  ( .CIN(sreg[2008]), .IN0(n2088), .IN1(
        \add_42/carry[2008] ), .COUT(\add_42/carry[2009] ), .SUM(o[2008]) );
  FADDER \add_42/U1_2009  ( .CIN(sreg[2009]), .IN0(n2087), .IN1(
        \add_42/carry[2009] ), .COUT(\add_42/carry[2010] ), .SUM(o[2009]) );
  FADDER \add_42/U1_2010  ( .CIN(sreg[2010]), .IN0(n2086), .IN1(
        \add_42/carry[2010] ), .COUT(\add_42/carry[2011] ), .SUM(o[2010]) );
  FADDER \add_42/U1_2011  ( .CIN(sreg[2011]), .IN0(n2085), .IN1(
        \add_42/carry[2011] ), .COUT(\add_42/carry[2012] ), .SUM(o[2011]) );
  FADDER \add_42/U1_2012  ( .CIN(sreg[2012]), .IN0(n2084), .IN1(
        \add_42/carry[2012] ), .COUT(\add_42/carry[2013] ), .SUM(o[2012]) );
  FADDER \add_42/U1_2013  ( .CIN(sreg[2013]), .IN0(n2083), .IN1(
        \add_42/carry[2013] ), .COUT(\add_42/carry[2014] ), .SUM(o[2013]) );
  FADDER \add_42/U1_2014  ( .CIN(sreg[2014]), .IN0(n2082), .IN1(
        \add_42/carry[2014] ), .COUT(\add_42/carry[2015] ), .SUM(o[2014]) );
  FADDER \add_42/U1_2015  ( .CIN(sreg[2015]), .IN0(n2081), .IN1(
        \add_42/carry[2015] ), .COUT(\add_42/carry[2016] ), .SUM(o[2015]) );
  FADDER \add_42/U1_2016  ( .CIN(sreg[2016]), .IN0(n2080), .IN1(
        \add_42/carry[2016] ), .COUT(\add_42/carry[2017] ), .SUM(o[2016]) );
  FADDER \add_42/U1_2017  ( .CIN(sreg[2017]), .IN0(n2079), .IN1(
        \add_42/carry[2017] ), .COUT(\add_42/carry[2018] ), .SUM(o[2017]) );
  FADDER \add_42/U1_2018  ( .CIN(sreg[2018]), .IN0(n2078), .IN1(
        \add_42/carry[2018] ), .COUT(\add_42/carry[2019] ), .SUM(o[2018]) );
  FADDER \add_42/U1_2019  ( .CIN(sreg[2019]), .IN0(n2077), .IN1(
        \add_42/carry[2019] ), .COUT(\add_42/carry[2020] ), .SUM(o[2019]) );
  FADDER \add_42/U1_2020  ( .CIN(sreg[2020]), .IN0(n2076), .IN1(
        \add_42/carry[2020] ), .COUT(\add_42/carry[2021] ), .SUM(o[2020]) );
  FADDER \add_42/U1_2021  ( .CIN(sreg[2021]), .IN0(n2075), .IN1(
        \add_42/carry[2021] ), .COUT(\add_42/carry[2022] ), .SUM(o[2021]) );
  FADDER \add_42/U1_2022  ( .CIN(sreg[2022]), .IN0(n2074), .IN1(
        \add_42/carry[2022] ), .COUT(\add_42/carry[2023] ), .SUM(o[2022]) );
  FADDER \add_42/U1_2023  ( .CIN(sreg[2023]), .IN0(n2073), .IN1(
        \add_42/carry[2023] ), .COUT(\add_42/carry[2024] ), .SUM(o[2023]) );
  FADDER \add_42/U1_2024  ( .CIN(sreg[2024]), .IN0(n2072), .IN1(
        \add_42/carry[2024] ), .COUT(\add_42/carry[2025] ), .SUM(o[2024]) );
  FADDER \add_42/U1_2025  ( .CIN(sreg[2025]), .IN0(n2071), .IN1(
        \add_42/carry[2025] ), .COUT(\add_42/carry[2026] ), .SUM(o[2025]) );
  FADDER \add_42/U1_2026  ( .CIN(sreg[2026]), .IN0(n2070), .IN1(
        \add_42/carry[2026] ), .COUT(\add_42/carry[2027] ), .SUM(o[2026]) );
  FADDER \add_42/U1_2027  ( .CIN(sreg[2027]), .IN0(n2069), .IN1(
        \add_42/carry[2027] ), .COUT(\add_42/carry[2028] ), .SUM(o[2027]) );
  FADDER \add_42/U1_2028  ( .CIN(sreg[2028]), .IN0(n2068), .IN1(
        \add_42/carry[2028] ), .COUT(\add_42/carry[2029] ), .SUM(o[2028]) );
  FADDER \add_42/U1_2029  ( .CIN(sreg[2029]), .IN0(n2067), .IN1(
        \add_42/carry[2029] ), .COUT(\add_42/carry[2030] ), .SUM(o[2029]) );
  FADDER \add_42/U1_2030  ( .CIN(sreg[2030]), .IN0(n2066), .IN1(
        \add_42/carry[2030] ), .COUT(\add_42/carry[2031] ), .SUM(o[2030]) );
  FADDER \add_42/U1_2031  ( .CIN(sreg[2031]), .IN0(n2065), .IN1(
        \add_42/carry[2031] ), .COUT(\add_42/carry[2032] ), .SUM(o[2031]) );
  FADDER \add_42/U1_2032  ( .CIN(sreg[2032]), .IN0(n2064), .IN1(
        \add_42/carry[2032] ), .COUT(\add_42/carry[2033] ), .SUM(o[2032]) );
  FADDER \add_42/U1_2033  ( .CIN(sreg[2033]), .IN0(n2063), .IN1(
        \add_42/carry[2033] ), .COUT(\add_42/carry[2034] ), .SUM(o[2033]) );
  FADDER \add_42/U1_2034  ( .CIN(sreg[2034]), .IN0(n2062), .IN1(
        \add_42/carry[2034] ), .COUT(\add_42/carry[2035] ), .SUM(o[2034]) );
  FADDER \add_42/U1_2035  ( .CIN(sreg[2035]), .IN0(n2061), .IN1(
        \add_42/carry[2035] ), .COUT(\add_42/carry[2036] ), .SUM(o[2035]) );
  FADDER \add_42/U1_2036  ( .CIN(sreg[2036]), .IN0(n2060), .IN1(
        \add_42/carry[2036] ), .COUT(\add_42/carry[2037] ), .SUM(o[2036]) );
  FADDER \add_42/U1_2037  ( .CIN(sreg[2037]), .IN0(n2059), .IN1(
        \add_42/carry[2037] ), .COUT(\add_42/carry[2038] ), .SUM(o[2037]) );
  FADDER \add_42/U1_2038  ( .CIN(sreg[2038]), .IN0(n2058), .IN1(
        \add_42/carry[2038] ), .COUT(\add_42/carry[2039] ), .SUM(o[2038]) );
  FADDER \add_42/U1_2039  ( .CIN(sreg[2039]), .IN0(n2057), .IN1(
        \add_42/carry[2039] ), .COUT(\add_42/carry[2040] ), .SUM(o[2039]) );
  FADDER \add_42/U1_2040  ( .CIN(sreg[2040]), .IN0(n2056), .IN1(
        \add_42/carry[2040] ), .COUT(\add_42/carry[2041] ), .SUM(o[2040]) );
  FADDER \add_42/U1_2041  ( .CIN(sreg[2041]), .IN0(n2055), .IN1(
        \add_42/carry[2041] ), .COUT(\add_42/carry[2042] ), .SUM(o[2041]) );
  FADDER \add_42/U1_2042  ( .CIN(sreg[2042]), .IN0(n2054), .IN1(
        \add_42/carry[2042] ), .COUT(\add_42/carry[2043] ), .SUM(o[2042]) );
  FADDER \add_42/U1_2043  ( .CIN(sreg[2043]), .IN0(n2053), .IN1(
        \add_42/carry[2043] ), .COUT(\add_42/carry[2044] ), .SUM(o[2043]) );
  FADDER \add_42/U1_2044  ( .CIN(sreg[2044]), .IN0(n2052), .IN1(
        \add_42/carry[2044] ), .COUT(\add_42/carry[2045] ), .SUM(o[2044]) );
  FADDER \add_42/U1_2045  ( .CIN(sreg[2045]), .IN0(n2051), .IN1(
        \add_42/carry[2045] ), .COUT(\add_42/carry[2046] ), .SUM(o[2045]) );
  FADDER \add_42/U1_2046  ( .CIN(sreg[2046]), .IN0(n2050), .IN1(
        \add_42/carry[2046] ), .COUT(\add_42/carry[2047] ), .SUM(o[2046]) );
  AND U2053 ( .A(sreg[1023]), .B(n3073), .Z(\add_42/carry[1024] ) );
  XOR U2054 ( .A(n3073), .B(sreg[1023]), .Z(o[1023]) );
  AND U2055 ( .A(g_input[1023]), .B(e_input[0]), .Z(n2050) );
  AND U2056 ( .A(g_input[1022]), .B(e_input[0]), .Z(n2051) );
  AND U2057 ( .A(g_input[1021]), .B(e_input[0]), .Z(n2052) );
  AND U2058 ( .A(g_input[1020]), .B(e_input[0]), .Z(n2053) );
  AND U2059 ( .A(g_input[1019]), .B(e_input[0]), .Z(n2054) );
  AND U2060 ( .A(g_input[1018]), .B(e_input[0]), .Z(n2055) );
  AND U2061 ( .A(g_input[1017]), .B(e_input[0]), .Z(n2056) );
  AND U2062 ( .A(g_input[1016]), .B(e_input[0]), .Z(n2057) );
  AND U2063 ( .A(g_input[1015]), .B(e_input[0]), .Z(n2058) );
  AND U2064 ( .A(g_input[1014]), .B(e_input[0]), .Z(n2059) );
  AND U2065 ( .A(g_input[1013]), .B(e_input[0]), .Z(n2060) );
  AND U2066 ( .A(g_input[1012]), .B(e_input[0]), .Z(n2061) );
  AND U2067 ( .A(g_input[1011]), .B(e_input[0]), .Z(n2062) );
  AND U2068 ( .A(g_input[1010]), .B(e_input[0]), .Z(n2063) );
  AND U2069 ( .A(g_input[1009]), .B(e_input[0]), .Z(n2064) );
  AND U2070 ( .A(g_input[1008]), .B(e_input[0]), .Z(n2065) );
  AND U2071 ( .A(g_input[1007]), .B(e_input[0]), .Z(n2066) );
  AND U2072 ( .A(g_input[1006]), .B(e_input[0]), .Z(n2067) );
  AND U2073 ( .A(g_input[1005]), .B(e_input[0]), .Z(n2068) );
  AND U2074 ( .A(g_input[1004]), .B(e_input[0]), .Z(n2069) );
  AND U2075 ( .A(g_input[1003]), .B(e_input[0]), .Z(n2070) );
  AND U2076 ( .A(g_input[1002]), .B(e_input[0]), .Z(n2071) );
  AND U2077 ( .A(g_input[1001]), .B(e_input[0]), .Z(n2072) );
  AND U2078 ( .A(g_input[1000]), .B(e_input[0]), .Z(n2073) );
  AND U2079 ( .A(g_input[999]), .B(e_input[0]), .Z(n2074) );
  AND U2080 ( .A(g_input[998]), .B(e_input[0]), .Z(n2075) );
  AND U2081 ( .A(g_input[997]), .B(e_input[0]), .Z(n2076) );
  AND U2082 ( .A(g_input[996]), .B(e_input[0]), .Z(n2077) );
  AND U2083 ( .A(g_input[995]), .B(e_input[0]), .Z(n2078) );
  AND U2084 ( .A(g_input[994]), .B(e_input[0]), .Z(n2079) );
  AND U2085 ( .A(g_input[993]), .B(e_input[0]), .Z(n2080) );
  AND U2086 ( .A(g_input[992]), .B(e_input[0]), .Z(n2081) );
  AND U2087 ( .A(g_input[991]), .B(e_input[0]), .Z(n2082) );
  AND U2088 ( .A(g_input[990]), .B(e_input[0]), .Z(n2083) );
  AND U2089 ( .A(g_input[989]), .B(e_input[0]), .Z(n2084) );
  AND U2090 ( .A(g_input[988]), .B(e_input[0]), .Z(n2085) );
  AND U2091 ( .A(g_input[987]), .B(e_input[0]), .Z(n2086) );
  AND U2092 ( .A(g_input[986]), .B(e_input[0]), .Z(n2087) );
  AND U2093 ( .A(g_input[985]), .B(e_input[0]), .Z(n2088) );
  AND U2094 ( .A(g_input[984]), .B(e_input[0]), .Z(n2089) );
  AND U2095 ( .A(g_input[983]), .B(e_input[0]), .Z(n2090) );
  AND U2096 ( .A(g_input[982]), .B(e_input[0]), .Z(n2091) );
  AND U2097 ( .A(g_input[981]), .B(e_input[0]), .Z(n2092) );
  AND U2098 ( .A(g_input[980]), .B(e_input[0]), .Z(n2093) );
  AND U2099 ( .A(g_input[979]), .B(e_input[0]), .Z(n2094) );
  AND U2100 ( .A(g_input[978]), .B(e_input[0]), .Z(n2095) );
  AND U2101 ( .A(g_input[977]), .B(e_input[0]), .Z(n2096) );
  AND U2102 ( .A(g_input[976]), .B(e_input[0]), .Z(n2097) );
  AND U2103 ( .A(g_input[975]), .B(e_input[0]), .Z(n2098) );
  AND U2104 ( .A(g_input[974]), .B(e_input[0]), .Z(n2099) );
  AND U2105 ( .A(g_input[973]), .B(e_input[0]), .Z(n2100) );
  AND U2106 ( .A(g_input[972]), .B(e_input[0]), .Z(n2101) );
  AND U2107 ( .A(g_input[971]), .B(e_input[0]), .Z(n2102) );
  AND U2108 ( .A(g_input[970]), .B(e_input[0]), .Z(n2103) );
  AND U2109 ( .A(g_input[969]), .B(e_input[0]), .Z(n2104) );
  AND U2110 ( .A(g_input[968]), .B(e_input[0]), .Z(n2105) );
  AND U2111 ( .A(g_input[967]), .B(e_input[0]), .Z(n2106) );
  AND U2112 ( .A(g_input[966]), .B(e_input[0]), .Z(n2107) );
  AND U2113 ( .A(g_input[965]), .B(e_input[0]), .Z(n2108) );
  AND U2114 ( .A(g_input[964]), .B(e_input[0]), .Z(n2109) );
  AND U2115 ( .A(g_input[963]), .B(e_input[0]), .Z(n2110) );
  AND U2116 ( .A(g_input[962]), .B(e_input[0]), .Z(n2111) );
  AND U2117 ( .A(g_input[961]), .B(e_input[0]), .Z(n2112) );
  AND U2118 ( .A(g_input[960]), .B(e_input[0]), .Z(n2113) );
  AND U2119 ( .A(g_input[959]), .B(e_input[0]), .Z(n2114) );
  AND U2120 ( .A(g_input[958]), .B(e_input[0]), .Z(n2115) );
  AND U2121 ( .A(g_input[957]), .B(e_input[0]), .Z(n2116) );
  AND U2122 ( .A(g_input[956]), .B(e_input[0]), .Z(n2117) );
  AND U2123 ( .A(g_input[955]), .B(e_input[0]), .Z(n2118) );
  AND U2124 ( .A(g_input[954]), .B(e_input[0]), .Z(n2119) );
  AND U2125 ( .A(g_input[953]), .B(e_input[0]), .Z(n2120) );
  AND U2126 ( .A(g_input[952]), .B(e_input[0]), .Z(n2121) );
  AND U2127 ( .A(g_input[951]), .B(e_input[0]), .Z(n2122) );
  AND U2128 ( .A(g_input[950]), .B(e_input[0]), .Z(n2123) );
  AND U2129 ( .A(g_input[949]), .B(e_input[0]), .Z(n2124) );
  AND U2130 ( .A(g_input[948]), .B(e_input[0]), .Z(n2125) );
  AND U2131 ( .A(g_input[947]), .B(e_input[0]), .Z(n2126) );
  AND U2132 ( .A(g_input[946]), .B(e_input[0]), .Z(n2127) );
  AND U2133 ( .A(g_input[945]), .B(e_input[0]), .Z(n2128) );
  AND U2134 ( .A(g_input[944]), .B(e_input[0]), .Z(n2129) );
  AND U2135 ( .A(g_input[943]), .B(e_input[0]), .Z(n2130) );
  AND U2136 ( .A(g_input[942]), .B(e_input[0]), .Z(n2131) );
  AND U2137 ( .A(g_input[941]), .B(e_input[0]), .Z(n2132) );
  AND U2138 ( .A(g_input[940]), .B(e_input[0]), .Z(n2133) );
  AND U2139 ( .A(g_input[939]), .B(e_input[0]), .Z(n2134) );
  AND U2140 ( .A(g_input[938]), .B(e_input[0]), .Z(n2135) );
  AND U2141 ( .A(g_input[937]), .B(e_input[0]), .Z(n2136) );
  AND U2142 ( .A(g_input[936]), .B(e_input[0]), .Z(n2137) );
  AND U2143 ( .A(g_input[935]), .B(e_input[0]), .Z(n2138) );
  AND U2144 ( .A(g_input[934]), .B(e_input[0]), .Z(n2139) );
  AND U2145 ( .A(g_input[933]), .B(e_input[0]), .Z(n2140) );
  AND U2146 ( .A(g_input[932]), .B(e_input[0]), .Z(n2141) );
  AND U2147 ( .A(g_input[931]), .B(e_input[0]), .Z(n2142) );
  AND U2148 ( .A(g_input[930]), .B(e_input[0]), .Z(n2143) );
  AND U2149 ( .A(g_input[929]), .B(e_input[0]), .Z(n2144) );
  AND U2150 ( .A(g_input[928]), .B(e_input[0]), .Z(n2145) );
  AND U2151 ( .A(g_input[927]), .B(e_input[0]), .Z(n2146) );
  AND U2152 ( .A(g_input[926]), .B(e_input[0]), .Z(n2147) );
  AND U2153 ( .A(g_input[925]), .B(e_input[0]), .Z(n2148) );
  AND U2154 ( .A(g_input[924]), .B(e_input[0]), .Z(n2149) );
  AND U2155 ( .A(g_input[923]), .B(e_input[0]), .Z(n2150) );
  AND U2156 ( .A(g_input[922]), .B(e_input[0]), .Z(n2151) );
  AND U2157 ( .A(g_input[921]), .B(e_input[0]), .Z(n2152) );
  AND U2158 ( .A(g_input[920]), .B(e_input[0]), .Z(n2153) );
  AND U2159 ( .A(g_input[919]), .B(e_input[0]), .Z(n2154) );
  AND U2160 ( .A(g_input[918]), .B(e_input[0]), .Z(n2155) );
  AND U2161 ( .A(g_input[917]), .B(e_input[0]), .Z(n2156) );
  AND U2162 ( .A(g_input[916]), .B(e_input[0]), .Z(n2157) );
  AND U2163 ( .A(g_input[915]), .B(e_input[0]), .Z(n2158) );
  AND U2164 ( .A(g_input[914]), .B(e_input[0]), .Z(n2159) );
  AND U2165 ( .A(g_input[913]), .B(e_input[0]), .Z(n2160) );
  AND U2166 ( .A(g_input[912]), .B(e_input[0]), .Z(n2161) );
  AND U2167 ( .A(g_input[911]), .B(e_input[0]), .Z(n2162) );
  AND U2168 ( .A(g_input[910]), .B(e_input[0]), .Z(n2163) );
  AND U2169 ( .A(g_input[909]), .B(e_input[0]), .Z(n2164) );
  AND U2170 ( .A(g_input[908]), .B(e_input[0]), .Z(n2165) );
  AND U2171 ( .A(g_input[907]), .B(e_input[0]), .Z(n2166) );
  AND U2172 ( .A(g_input[906]), .B(e_input[0]), .Z(n2167) );
  AND U2173 ( .A(g_input[905]), .B(e_input[0]), .Z(n2168) );
  AND U2174 ( .A(g_input[904]), .B(e_input[0]), .Z(n2169) );
  AND U2175 ( .A(g_input[903]), .B(e_input[0]), .Z(n2170) );
  AND U2176 ( .A(g_input[902]), .B(e_input[0]), .Z(n2171) );
  AND U2177 ( .A(g_input[901]), .B(e_input[0]), .Z(n2172) );
  AND U2178 ( .A(g_input[900]), .B(e_input[0]), .Z(n2173) );
  AND U2179 ( .A(g_input[899]), .B(e_input[0]), .Z(n2174) );
  AND U2180 ( .A(g_input[898]), .B(e_input[0]), .Z(n2175) );
  AND U2181 ( .A(g_input[897]), .B(e_input[0]), .Z(n2176) );
  AND U2182 ( .A(g_input[896]), .B(e_input[0]), .Z(n2177) );
  AND U2183 ( .A(g_input[895]), .B(e_input[0]), .Z(n2178) );
  AND U2184 ( .A(g_input[894]), .B(e_input[0]), .Z(n2179) );
  AND U2185 ( .A(g_input[893]), .B(e_input[0]), .Z(n2180) );
  AND U2186 ( .A(g_input[892]), .B(e_input[0]), .Z(n2181) );
  AND U2187 ( .A(g_input[891]), .B(e_input[0]), .Z(n2182) );
  AND U2188 ( .A(g_input[890]), .B(e_input[0]), .Z(n2183) );
  AND U2189 ( .A(g_input[889]), .B(e_input[0]), .Z(n2184) );
  AND U2190 ( .A(g_input[888]), .B(e_input[0]), .Z(n2185) );
  AND U2191 ( .A(g_input[887]), .B(e_input[0]), .Z(n2186) );
  AND U2192 ( .A(g_input[886]), .B(e_input[0]), .Z(n2187) );
  AND U2193 ( .A(g_input[885]), .B(e_input[0]), .Z(n2188) );
  AND U2194 ( .A(g_input[884]), .B(e_input[0]), .Z(n2189) );
  AND U2195 ( .A(g_input[883]), .B(e_input[0]), .Z(n2190) );
  AND U2196 ( .A(g_input[882]), .B(e_input[0]), .Z(n2191) );
  AND U2197 ( .A(g_input[881]), .B(e_input[0]), .Z(n2192) );
  AND U2198 ( .A(g_input[880]), .B(e_input[0]), .Z(n2193) );
  AND U2199 ( .A(g_input[879]), .B(e_input[0]), .Z(n2194) );
  AND U2200 ( .A(g_input[878]), .B(e_input[0]), .Z(n2195) );
  AND U2201 ( .A(g_input[877]), .B(e_input[0]), .Z(n2196) );
  AND U2202 ( .A(g_input[876]), .B(e_input[0]), .Z(n2197) );
  AND U2203 ( .A(g_input[875]), .B(e_input[0]), .Z(n2198) );
  AND U2204 ( .A(g_input[874]), .B(e_input[0]), .Z(n2199) );
  AND U2205 ( .A(g_input[873]), .B(e_input[0]), .Z(n2200) );
  AND U2206 ( .A(g_input[872]), .B(e_input[0]), .Z(n2201) );
  AND U2207 ( .A(g_input[871]), .B(e_input[0]), .Z(n2202) );
  AND U2208 ( .A(g_input[870]), .B(e_input[0]), .Z(n2203) );
  AND U2209 ( .A(g_input[869]), .B(e_input[0]), .Z(n2204) );
  AND U2210 ( .A(g_input[868]), .B(e_input[0]), .Z(n2205) );
  AND U2211 ( .A(g_input[867]), .B(e_input[0]), .Z(n2206) );
  AND U2212 ( .A(g_input[866]), .B(e_input[0]), .Z(n2207) );
  AND U2213 ( .A(g_input[865]), .B(e_input[0]), .Z(n2208) );
  AND U2214 ( .A(g_input[864]), .B(e_input[0]), .Z(n2209) );
  AND U2215 ( .A(g_input[863]), .B(e_input[0]), .Z(n2210) );
  AND U2216 ( .A(g_input[862]), .B(e_input[0]), .Z(n2211) );
  AND U2217 ( .A(g_input[861]), .B(e_input[0]), .Z(n2212) );
  AND U2218 ( .A(g_input[860]), .B(e_input[0]), .Z(n2213) );
  AND U2219 ( .A(g_input[859]), .B(e_input[0]), .Z(n2214) );
  AND U2220 ( .A(g_input[858]), .B(e_input[0]), .Z(n2215) );
  AND U2221 ( .A(g_input[857]), .B(e_input[0]), .Z(n2216) );
  AND U2222 ( .A(g_input[856]), .B(e_input[0]), .Z(n2217) );
  AND U2223 ( .A(g_input[855]), .B(e_input[0]), .Z(n2218) );
  AND U2224 ( .A(g_input[854]), .B(e_input[0]), .Z(n2219) );
  AND U2225 ( .A(g_input[853]), .B(e_input[0]), .Z(n2220) );
  AND U2226 ( .A(g_input[852]), .B(e_input[0]), .Z(n2221) );
  AND U2227 ( .A(g_input[851]), .B(e_input[0]), .Z(n2222) );
  AND U2228 ( .A(g_input[850]), .B(e_input[0]), .Z(n2223) );
  AND U2229 ( .A(g_input[849]), .B(e_input[0]), .Z(n2224) );
  AND U2230 ( .A(g_input[848]), .B(e_input[0]), .Z(n2225) );
  AND U2231 ( .A(g_input[847]), .B(e_input[0]), .Z(n2226) );
  AND U2232 ( .A(g_input[846]), .B(e_input[0]), .Z(n2227) );
  AND U2233 ( .A(g_input[845]), .B(e_input[0]), .Z(n2228) );
  AND U2234 ( .A(g_input[844]), .B(e_input[0]), .Z(n2229) );
  AND U2235 ( .A(g_input[843]), .B(e_input[0]), .Z(n2230) );
  AND U2236 ( .A(g_input[842]), .B(e_input[0]), .Z(n2231) );
  AND U2237 ( .A(g_input[841]), .B(e_input[0]), .Z(n2232) );
  AND U2238 ( .A(g_input[840]), .B(e_input[0]), .Z(n2233) );
  AND U2239 ( .A(g_input[839]), .B(e_input[0]), .Z(n2234) );
  AND U2240 ( .A(g_input[838]), .B(e_input[0]), .Z(n2235) );
  AND U2241 ( .A(g_input[837]), .B(e_input[0]), .Z(n2236) );
  AND U2242 ( .A(g_input[836]), .B(e_input[0]), .Z(n2237) );
  AND U2243 ( .A(g_input[835]), .B(e_input[0]), .Z(n2238) );
  AND U2244 ( .A(g_input[834]), .B(e_input[0]), .Z(n2239) );
  AND U2245 ( .A(g_input[833]), .B(e_input[0]), .Z(n2240) );
  AND U2246 ( .A(g_input[832]), .B(e_input[0]), .Z(n2241) );
  AND U2247 ( .A(g_input[831]), .B(e_input[0]), .Z(n2242) );
  AND U2248 ( .A(g_input[830]), .B(e_input[0]), .Z(n2243) );
  AND U2249 ( .A(g_input[829]), .B(e_input[0]), .Z(n2244) );
  AND U2250 ( .A(g_input[828]), .B(e_input[0]), .Z(n2245) );
  AND U2251 ( .A(g_input[827]), .B(e_input[0]), .Z(n2246) );
  AND U2252 ( .A(g_input[826]), .B(e_input[0]), .Z(n2247) );
  AND U2253 ( .A(g_input[825]), .B(e_input[0]), .Z(n2248) );
  AND U2254 ( .A(g_input[824]), .B(e_input[0]), .Z(n2249) );
  AND U2255 ( .A(g_input[823]), .B(e_input[0]), .Z(n2250) );
  AND U2256 ( .A(g_input[822]), .B(e_input[0]), .Z(n2251) );
  AND U2257 ( .A(g_input[821]), .B(e_input[0]), .Z(n2252) );
  AND U2258 ( .A(g_input[820]), .B(e_input[0]), .Z(n2253) );
  AND U2259 ( .A(g_input[819]), .B(e_input[0]), .Z(n2254) );
  AND U2260 ( .A(g_input[818]), .B(e_input[0]), .Z(n2255) );
  AND U2261 ( .A(g_input[817]), .B(e_input[0]), .Z(n2256) );
  AND U2262 ( .A(g_input[816]), .B(e_input[0]), .Z(n2257) );
  AND U2263 ( .A(g_input[815]), .B(e_input[0]), .Z(n2258) );
  AND U2264 ( .A(g_input[814]), .B(e_input[0]), .Z(n2259) );
  AND U2265 ( .A(g_input[813]), .B(e_input[0]), .Z(n2260) );
  AND U2266 ( .A(g_input[812]), .B(e_input[0]), .Z(n2261) );
  AND U2267 ( .A(g_input[811]), .B(e_input[0]), .Z(n2262) );
  AND U2268 ( .A(g_input[810]), .B(e_input[0]), .Z(n2263) );
  AND U2269 ( .A(g_input[809]), .B(e_input[0]), .Z(n2264) );
  AND U2270 ( .A(g_input[808]), .B(e_input[0]), .Z(n2265) );
  AND U2271 ( .A(g_input[807]), .B(e_input[0]), .Z(n2266) );
  AND U2272 ( .A(g_input[806]), .B(e_input[0]), .Z(n2267) );
  AND U2273 ( .A(g_input[805]), .B(e_input[0]), .Z(n2268) );
  AND U2274 ( .A(g_input[804]), .B(e_input[0]), .Z(n2269) );
  AND U2275 ( .A(g_input[803]), .B(e_input[0]), .Z(n2270) );
  AND U2276 ( .A(g_input[802]), .B(e_input[0]), .Z(n2271) );
  AND U2277 ( .A(g_input[801]), .B(e_input[0]), .Z(n2272) );
  AND U2278 ( .A(g_input[800]), .B(e_input[0]), .Z(n2273) );
  AND U2279 ( .A(g_input[799]), .B(e_input[0]), .Z(n2274) );
  AND U2280 ( .A(g_input[798]), .B(e_input[0]), .Z(n2275) );
  AND U2281 ( .A(g_input[797]), .B(e_input[0]), .Z(n2276) );
  AND U2282 ( .A(g_input[796]), .B(e_input[0]), .Z(n2277) );
  AND U2283 ( .A(g_input[795]), .B(e_input[0]), .Z(n2278) );
  AND U2284 ( .A(g_input[794]), .B(e_input[0]), .Z(n2279) );
  AND U2285 ( .A(g_input[793]), .B(e_input[0]), .Z(n2280) );
  AND U2286 ( .A(g_input[792]), .B(e_input[0]), .Z(n2281) );
  AND U2287 ( .A(g_input[791]), .B(e_input[0]), .Z(n2282) );
  AND U2288 ( .A(g_input[790]), .B(e_input[0]), .Z(n2283) );
  AND U2289 ( .A(g_input[789]), .B(e_input[0]), .Z(n2284) );
  AND U2290 ( .A(g_input[788]), .B(e_input[0]), .Z(n2285) );
  AND U2291 ( .A(g_input[787]), .B(e_input[0]), .Z(n2286) );
  AND U2292 ( .A(g_input[786]), .B(e_input[0]), .Z(n2287) );
  AND U2293 ( .A(g_input[785]), .B(e_input[0]), .Z(n2288) );
  AND U2294 ( .A(g_input[784]), .B(e_input[0]), .Z(n2289) );
  AND U2295 ( .A(g_input[783]), .B(e_input[0]), .Z(n2290) );
  AND U2296 ( .A(g_input[782]), .B(e_input[0]), .Z(n2291) );
  AND U2297 ( .A(g_input[781]), .B(e_input[0]), .Z(n2292) );
  AND U2298 ( .A(g_input[780]), .B(e_input[0]), .Z(n2293) );
  AND U2299 ( .A(g_input[779]), .B(e_input[0]), .Z(n2294) );
  AND U2300 ( .A(g_input[778]), .B(e_input[0]), .Z(n2295) );
  AND U2301 ( .A(g_input[777]), .B(e_input[0]), .Z(n2296) );
  AND U2302 ( .A(g_input[776]), .B(e_input[0]), .Z(n2297) );
  AND U2303 ( .A(g_input[775]), .B(e_input[0]), .Z(n2298) );
  AND U2304 ( .A(g_input[774]), .B(e_input[0]), .Z(n2299) );
  AND U2305 ( .A(g_input[773]), .B(e_input[0]), .Z(n2300) );
  AND U2306 ( .A(g_input[772]), .B(e_input[0]), .Z(n2301) );
  AND U2307 ( .A(g_input[771]), .B(e_input[0]), .Z(n2302) );
  AND U2308 ( .A(g_input[770]), .B(e_input[0]), .Z(n2303) );
  AND U2309 ( .A(g_input[769]), .B(e_input[0]), .Z(n2304) );
  AND U2310 ( .A(g_input[768]), .B(e_input[0]), .Z(n2305) );
  AND U2311 ( .A(g_input[767]), .B(e_input[0]), .Z(n2306) );
  AND U2312 ( .A(g_input[766]), .B(e_input[0]), .Z(n2307) );
  AND U2313 ( .A(g_input[765]), .B(e_input[0]), .Z(n2308) );
  AND U2314 ( .A(g_input[764]), .B(e_input[0]), .Z(n2309) );
  AND U2315 ( .A(g_input[763]), .B(e_input[0]), .Z(n2310) );
  AND U2316 ( .A(g_input[762]), .B(e_input[0]), .Z(n2311) );
  AND U2317 ( .A(g_input[761]), .B(e_input[0]), .Z(n2312) );
  AND U2318 ( .A(g_input[760]), .B(e_input[0]), .Z(n2313) );
  AND U2319 ( .A(g_input[759]), .B(e_input[0]), .Z(n2314) );
  AND U2320 ( .A(g_input[758]), .B(e_input[0]), .Z(n2315) );
  AND U2321 ( .A(g_input[757]), .B(e_input[0]), .Z(n2316) );
  AND U2322 ( .A(g_input[756]), .B(e_input[0]), .Z(n2317) );
  AND U2323 ( .A(g_input[755]), .B(e_input[0]), .Z(n2318) );
  AND U2324 ( .A(g_input[754]), .B(e_input[0]), .Z(n2319) );
  AND U2325 ( .A(g_input[753]), .B(e_input[0]), .Z(n2320) );
  AND U2326 ( .A(g_input[752]), .B(e_input[0]), .Z(n2321) );
  AND U2327 ( .A(g_input[751]), .B(e_input[0]), .Z(n2322) );
  AND U2328 ( .A(g_input[750]), .B(e_input[0]), .Z(n2323) );
  AND U2329 ( .A(g_input[749]), .B(e_input[0]), .Z(n2324) );
  AND U2330 ( .A(g_input[748]), .B(e_input[0]), .Z(n2325) );
  AND U2331 ( .A(g_input[747]), .B(e_input[0]), .Z(n2326) );
  AND U2332 ( .A(g_input[746]), .B(e_input[0]), .Z(n2327) );
  AND U2333 ( .A(g_input[745]), .B(e_input[0]), .Z(n2328) );
  AND U2334 ( .A(g_input[744]), .B(e_input[0]), .Z(n2329) );
  AND U2335 ( .A(g_input[743]), .B(e_input[0]), .Z(n2330) );
  AND U2336 ( .A(g_input[742]), .B(e_input[0]), .Z(n2331) );
  AND U2337 ( .A(g_input[741]), .B(e_input[0]), .Z(n2332) );
  AND U2338 ( .A(g_input[740]), .B(e_input[0]), .Z(n2333) );
  AND U2339 ( .A(g_input[739]), .B(e_input[0]), .Z(n2334) );
  AND U2340 ( .A(g_input[738]), .B(e_input[0]), .Z(n2335) );
  AND U2341 ( .A(g_input[737]), .B(e_input[0]), .Z(n2336) );
  AND U2342 ( .A(g_input[736]), .B(e_input[0]), .Z(n2337) );
  AND U2343 ( .A(g_input[735]), .B(e_input[0]), .Z(n2338) );
  AND U2344 ( .A(g_input[734]), .B(e_input[0]), .Z(n2339) );
  AND U2345 ( .A(g_input[733]), .B(e_input[0]), .Z(n2340) );
  AND U2346 ( .A(g_input[732]), .B(e_input[0]), .Z(n2341) );
  AND U2347 ( .A(g_input[731]), .B(e_input[0]), .Z(n2342) );
  AND U2348 ( .A(g_input[730]), .B(e_input[0]), .Z(n2343) );
  AND U2349 ( .A(g_input[729]), .B(e_input[0]), .Z(n2344) );
  AND U2350 ( .A(g_input[728]), .B(e_input[0]), .Z(n2345) );
  AND U2351 ( .A(g_input[727]), .B(e_input[0]), .Z(n2346) );
  AND U2352 ( .A(g_input[726]), .B(e_input[0]), .Z(n2347) );
  AND U2353 ( .A(g_input[725]), .B(e_input[0]), .Z(n2348) );
  AND U2354 ( .A(g_input[724]), .B(e_input[0]), .Z(n2349) );
  AND U2355 ( .A(g_input[723]), .B(e_input[0]), .Z(n2350) );
  AND U2356 ( .A(g_input[722]), .B(e_input[0]), .Z(n2351) );
  AND U2357 ( .A(g_input[721]), .B(e_input[0]), .Z(n2352) );
  AND U2358 ( .A(g_input[720]), .B(e_input[0]), .Z(n2353) );
  AND U2359 ( .A(g_input[719]), .B(e_input[0]), .Z(n2354) );
  AND U2360 ( .A(g_input[718]), .B(e_input[0]), .Z(n2355) );
  AND U2361 ( .A(g_input[717]), .B(e_input[0]), .Z(n2356) );
  AND U2362 ( .A(g_input[716]), .B(e_input[0]), .Z(n2357) );
  AND U2363 ( .A(g_input[715]), .B(e_input[0]), .Z(n2358) );
  AND U2364 ( .A(g_input[714]), .B(e_input[0]), .Z(n2359) );
  AND U2365 ( .A(g_input[713]), .B(e_input[0]), .Z(n2360) );
  AND U2366 ( .A(g_input[712]), .B(e_input[0]), .Z(n2361) );
  AND U2367 ( .A(g_input[711]), .B(e_input[0]), .Z(n2362) );
  AND U2368 ( .A(g_input[710]), .B(e_input[0]), .Z(n2363) );
  AND U2369 ( .A(g_input[709]), .B(e_input[0]), .Z(n2364) );
  AND U2370 ( .A(g_input[708]), .B(e_input[0]), .Z(n2365) );
  AND U2371 ( .A(g_input[707]), .B(e_input[0]), .Z(n2366) );
  AND U2372 ( .A(g_input[706]), .B(e_input[0]), .Z(n2367) );
  AND U2373 ( .A(g_input[705]), .B(e_input[0]), .Z(n2368) );
  AND U2374 ( .A(g_input[704]), .B(e_input[0]), .Z(n2369) );
  AND U2375 ( .A(g_input[703]), .B(e_input[0]), .Z(n2370) );
  AND U2376 ( .A(g_input[702]), .B(e_input[0]), .Z(n2371) );
  AND U2377 ( .A(g_input[701]), .B(e_input[0]), .Z(n2372) );
  AND U2378 ( .A(g_input[700]), .B(e_input[0]), .Z(n2373) );
  AND U2379 ( .A(g_input[699]), .B(e_input[0]), .Z(n2374) );
  AND U2380 ( .A(g_input[698]), .B(e_input[0]), .Z(n2375) );
  AND U2381 ( .A(g_input[697]), .B(e_input[0]), .Z(n2376) );
  AND U2382 ( .A(g_input[696]), .B(e_input[0]), .Z(n2377) );
  AND U2383 ( .A(g_input[695]), .B(e_input[0]), .Z(n2378) );
  AND U2384 ( .A(g_input[694]), .B(e_input[0]), .Z(n2379) );
  AND U2385 ( .A(g_input[693]), .B(e_input[0]), .Z(n2380) );
  AND U2386 ( .A(g_input[692]), .B(e_input[0]), .Z(n2381) );
  AND U2387 ( .A(g_input[691]), .B(e_input[0]), .Z(n2382) );
  AND U2388 ( .A(g_input[690]), .B(e_input[0]), .Z(n2383) );
  AND U2389 ( .A(g_input[689]), .B(e_input[0]), .Z(n2384) );
  AND U2390 ( .A(g_input[688]), .B(e_input[0]), .Z(n2385) );
  AND U2391 ( .A(g_input[687]), .B(e_input[0]), .Z(n2386) );
  AND U2392 ( .A(g_input[686]), .B(e_input[0]), .Z(n2387) );
  AND U2393 ( .A(g_input[685]), .B(e_input[0]), .Z(n2388) );
  AND U2394 ( .A(g_input[684]), .B(e_input[0]), .Z(n2389) );
  AND U2395 ( .A(g_input[683]), .B(e_input[0]), .Z(n2390) );
  AND U2396 ( .A(g_input[682]), .B(e_input[0]), .Z(n2391) );
  AND U2397 ( .A(g_input[681]), .B(e_input[0]), .Z(n2392) );
  AND U2398 ( .A(g_input[680]), .B(e_input[0]), .Z(n2393) );
  AND U2399 ( .A(g_input[679]), .B(e_input[0]), .Z(n2394) );
  AND U2400 ( .A(g_input[678]), .B(e_input[0]), .Z(n2395) );
  AND U2401 ( .A(g_input[677]), .B(e_input[0]), .Z(n2396) );
  AND U2402 ( .A(g_input[676]), .B(e_input[0]), .Z(n2397) );
  AND U2403 ( .A(g_input[675]), .B(e_input[0]), .Z(n2398) );
  AND U2404 ( .A(g_input[674]), .B(e_input[0]), .Z(n2399) );
  AND U2405 ( .A(g_input[673]), .B(e_input[0]), .Z(n2400) );
  AND U2406 ( .A(g_input[672]), .B(e_input[0]), .Z(n2401) );
  AND U2407 ( .A(g_input[671]), .B(e_input[0]), .Z(n2402) );
  AND U2408 ( .A(g_input[670]), .B(e_input[0]), .Z(n2403) );
  AND U2409 ( .A(g_input[669]), .B(e_input[0]), .Z(n2404) );
  AND U2410 ( .A(g_input[668]), .B(e_input[0]), .Z(n2405) );
  AND U2411 ( .A(g_input[667]), .B(e_input[0]), .Z(n2406) );
  AND U2412 ( .A(g_input[666]), .B(e_input[0]), .Z(n2407) );
  AND U2413 ( .A(g_input[665]), .B(e_input[0]), .Z(n2408) );
  AND U2414 ( .A(g_input[664]), .B(e_input[0]), .Z(n2409) );
  AND U2415 ( .A(g_input[663]), .B(e_input[0]), .Z(n2410) );
  AND U2416 ( .A(g_input[662]), .B(e_input[0]), .Z(n2411) );
  AND U2417 ( .A(g_input[661]), .B(e_input[0]), .Z(n2412) );
  AND U2418 ( .A(g_input[660]), .B(e_input[0]), .Z(n2413) );
  AND U2419 ( .A(g_input[659]), .B(e_input[0]), .Z(n2414) );
  AND U2420 ( .A(g_input[658]), .B(e_input[0]), .Z(n2415) );
  AND U2421 ( .A(g_input[657]), .B(e_input[0]), .Z(n2416) );
  AND U2422 ( .A(g_input[656]), .B(e_input[0]), .Z(n2417) );
  AND U2423 ( .A(g_input[655]), .B(e_input[0]), .Z(n2418) );
  AND U2424 ( .A(g_input[654]), .B(e_input[0]), .Z(n2419) );
  AND U2425 ( .A(g_input[653]), .B(e_input[0]), .Z(n2420) );
  AND U2426 ( .A(g_input[652]), .B(e_input[0]), .Z(n2421) );
  AND U2427 ( .A(g_input[651]), .B(e_input[0]), .Z(n2422) );
  AND U2428 ( .A(g_input[650]), .B(e_input[0]), .Z(n2423) );
  AND U2429 ( .A(g_input[649]), .B(e_input[0]), .Z(n2424) );
  AND U2430 ( .A(g_input[648]), .B(e_input[0]), .Z(n2425) );
  AND U2431 ( .A(g_input[647]), .B(e_input[0]), .Z(n2426) );
  AND U2432 ( .A(g_input[646]), .B(e_input[0]), .Z(n2427) );
  AND U2433 ( .A(g_input[645]), .B(e_input[0]), .Z(n2428) );
  AND U2434 ( .A(g_input[644]), .B(e_input[0]), .Z(n2429) );
  AND U2435 ( .A(g_input[643]), .B(e_input[0]), .Z(n2430) );
  AND U2436 ( .A(g_input[642]), .B(e_input[0]), .Z(n2431) );
  AND U2437 ( .A(g_input[641]), .B(e_input[0]), .Z(n2432) );
  AND U2438 ( .A(g_input[640]), .B(e_input[0]), .Z(n2433) );
  AND U2439 ( .A(g_input[639]), .B(e_input[0]), .Z(n2434) );
  AND U2440 ( .A(g_input[638]), .B(e_input[0]), .Z(n2435) );
  AND U2441 ( .A(g_input[637]), .B(e_input[0]), .Z(n2436) );
  AND U2442 ( .A(g_input[636]), .B(e_input[0]), .Z(n2437) );
  AND U2443 ( .A(g_input[635]), .B(e_input[0]), .Z(n2438) );
  AND U2444 ( .A(g_input[634]), .B(e_input[0]), .Z(n2439) );
  AND U2445 ( .A(g_input[633]), .B(e_input[0]), .Z(n2440) );
  AND U2446 ( .A(g_input[632]), .B(e_input[0]), .Z(n2441) );
  AND U2447 ( .A(g_input[631]), .B(e_input[0]), .Z(n2442) );
  AND U2448 ( .A(g_input[630]), .B(e_input[0]), .Z(n2443) );
  AND U2449 ( .A(g_input[629]), .B(e_input[0]), .Z(n2444) );
  AND U2450 ( .A(g_input[628]), .B(e_input[0]), .Z(n2445) );
  AND U2451 ( .A(g_input[627]), .B(e_input[0]), .Z(n2446) );
  AND U2452 ( .A(g_input[626]), .B(e_input[0]), .Z(n2447) );
  AND U2453 ( .A(g_input[625]), .B(e_input[0]), .Z(n2448) );
  AND U2454 ( .A(g_input[624]), .B(e_input[0]), .Z(n2449) );
  AND U2455 ( .A(g_input[623]), .B(e_input[0]), .Z(n2450) );
  AND U2456 ( .A(g_input[622]), .B(e_input[0]), .Z(n2451) );
  AND U2457 ( .A(g_input[621]), .B(e_input[0]), .Z(n2452) );
  AND U2458 ( .A(g_input[620]), .B(e_input[0]), .Z(n2453) );
  AND U2459 ( .A(g_input[619]), .B(e_input[0]), .Z(n2454) );
  AND U2460 ( .A(g_input[618]), .B(e_input[0]), .Z(n2455) );
  AND U2461 ( .A(g_input[617]), .B(e_input[0]), .Z(n2456) );
  AND U2462 ( .A(g_input[616]), .B(e_input[0]), .Z(n2457) );
  AND U2463 ( .A(g_input[615]), .B(e_input[0]), .Z(n2458) );
  AND U2464 ( .A(g_input[614]), .B(e_input[0]), .Z(n2459) );
  AND U2465 ( .A(g_input[613]), .B(e_input[0]), .Z(n2460) );
  AND U2466 ( .A(g_input[612]), .B(e_input[0]), .Z(n2461) );
  AND U2467 ( .A(g_input[611]), .B(e_input[0]), .Z(n2462) );
  AND U2468 ( .A(g_input[610]), .B(e_input[0]), .Z(n2463) );
  AND U2469 ( .A(g_input[609]), .B(e_input[0]), .Z(n2464) );
  AND U2470 ( .A(g_input[608]), .B(e_input[0]), .Z(n2465) );
  AND U2471 ( .A(g_input[607]), .B(e_input[0]), .Z(n2466) );
  AND U2472 ( .A(g_input[606]), .B(e_input[0]), .Z(n2467) );
  AND U2473 ( .A(g_input[605]), .B(e_input[0]), .Z(n2468) );
  AND U2474 ( .A(g_input[604]), .B(e_input[0]), .Z(n2469) );
  AND U2475 ( .A(g_input[603]), .B(e_input[0]), .Z(n2470) );
  AND U2476 ( .A(g_input[602]), .B(e_input[0]), .Z(n2471) );
  AND U2477 ( .A(g_input[601]), .B(e_input[0]), .Z(n2472) );
  AND U2478 ( .A(g_input[600]), .B(e_input[0]), .Z(n2473) );
  AND U2479 ( .A(g_input[599]), .B(e_input[0]), .Z(n2474) );
  AND U2480 ( .A(g_input[598]), .B(e_input[0]), .Z(n2475) );
  AND U2481 ( .A(g_input[597]), .B(e_input[0]), .Z(n2476) );
  AND U2482 ( .A(g_input[596]), .B(e_input[0]), .Z(n2477) );
  AND U2483 ( .A(g_input[595]), .B(e_input[0]), .Z(n2478) );
  AND U2484 ( .A(g_input[594]), .B(e_input[0]), .Z(n2479) );
  AND U2485 ( .A(g_input[593]), .B(e_input[0]), .Z(n2480) );
  AND U2486 ( .A(g_input[592]), .B(e_input[0]), .Z(n2481) );
  AND U2487 ( .A(g_input[591]), .B(e_input[0]), .Z(n2482) );
  AND U2488 ( .A(g_input[590]), .B(e_input[0]), .Z(n2483) );
  AND U2489 ( .A(g_input[589]), .B(e_input[0]), .Z(n2484) );
  AND U2490 ( .A(g_input[588]), .B(e_input[0]), .Z(n2485) );
  AND U2491 ( .A(g_input[587]), .B(e_input[0]), .Z(n2486) );
  AND U2492 ( .A(g_input[586]), .B(e_input[0]), .Z(n2487) );
  AND U2493 ( .A(g_input[585]), .B(e_input[0]), .Z(n2488) );
  AND U2494 ( .A(g_input[584]), .B(e_input[0]), .Z(n2489) );
  AND U2495 ( .A(g_input[583]), .B(e_input[0]), .Z(n2490) );
  AND U2496 ( .A(g_input[582]), .B(e_input[0]), .Z(n2491) );
  AND U2497 ( .A(g_input[581]), .B(e_input[0]), .Z(n2492) );
  AND U2498 ( .A(g_input[580]), .B(e_input[0]), .Z(n2493) );
  AND U2499 ( .A(g_input[579]), .B(e_input[0]), .Z(n2494) );
  AND U2500 ( .A(g_input[578]), .B(e_input[0]), .Z(n2495) );
  AND U2501 ( .A(g_input[577]), .B(e_input[0]), .Z(n2496) );
  AND U2502 ( .A(g_input[576]), .B(e_input[0]), .Z(n2497) );
  AND U2503 ( .A(g_input[575]), .B(e_input[0]), .Z(n2498) );
  AND U2504 ( .A(g_input[574]), .B(e_input[0]), .Z(n2499) );
  AND U2505 ( .A(g_input[573]), .B(e_input[0]), .Z(n2500) );
  AND U2506 ( .A(g_input[572]), .B(e_input[0]), .Z(n2501) );
  AND U2507 ( .A(g_input[571]), .B(e_input[0]), .Z(n2502) );
  AND U2508 ( .A(g_input[570]), .B(e_input[0]), .Z(n2503) );
  AND U2509 ( .A(g_input[569]), .B(e_input[0]), .Z(n2504) );
  AND U2510 ( .A(g_input[568]), .B(e_input[0]), .Z(n2505) );
  AND U2511 ( .A(g_input[567]), .B(e_input[0]), .Z(n2506) );
  AND U2512 ( .A(g_input[566]), .B(e_input[0]), .Z(n2507) );
  AND U2513 ( .A(g_input[565]), .B(e_input[0]), .Z(n2508) );
  AND U2514 ( .A(g_input[564]), .B(e_input[0]), .Z(n2509) );
  AND U2515 ( .A(g_input[563]), .B(e_input[0]), .Z(n2510) );
  AND U2516 ( .A(g_input[562]), .B(e_input[0]), .Z(n2511) );
  AND U2517 ( .A(g_input[561]), .B(e_input[0]), .Z(n2512) );
  AND U2518 ( .A(g_input[560]), .B(e_input[0]), .Z(n2513) );
  AND U2519 ( .A(g_input[559]), .B(e_input[0]), .Z(n2514) );
  AND U2520 ( .A(g_input[558]), .B(e_input[0]), .Z(n2515) );
  AND U2521 ( .A(g_input[557]), .B(e_input[0]), .Z(n2516) );
  AND U2522 ( .A(g_input[556]), .B(e_input[0]), .Z(n2517) );
  AND U2523 ( .A(g_input[555]), .B(e_input[0]), .Z(n2518) );
  AND U2524 ( .A(g_input[554]), .B(e_input[0]), .Z(n2519) );
  AND U2525 ( .A(g_input[553]), .B(e_input[0]), .Z(n2520) );
  AND U2526 ( .A(g_input[552]), .B(e_input[0]), .Z(n2521) );
  AND U2527 ( .A(g_input[551]), .B(e_input[0]), .Z(n2522) );
  AND U2528 ( .A(g_input[550]), .B(e_input[0]), .Z(n2523) );
  AND U2529 ( .A(g_input[549]), .B(e_input[0]), .Z(n2524) );
  AND U2530 ( .A(g_input[548]), .B(e_input[0]), .Z(n2525) );
  AND U2531 ( .A(g_input[547]), .B(e_input[0]), .Z(n2526) );
  AND U2532 ( .A(g_input[546]), .B(e_input[0]), .Z(n2527) );
  AND U2533 ( .A(g_input[545]), .B(e_input[0]), .Z(n2528) );
  AND U2534 ( .A(g_input[544]), .B(e_input[0]), .Z(n2529) );
  AND U2535 ( .A(g_input[543]), .B(e_input[0]), .Z(n2530) );
  AND U2536 ( .A(g_input[542]), .B(e_input[0]), .Z(n2531) );
  AND U2537 ( .A(g_input[541]), .B(e_input[0]), .Z(n2532) );
  AND U2538 ( .A(g_input[540]), .B(e_input[0]), .Z(n2533) );
  AND U2539 ( .A(g_input[539]), .B(e_input[0]), .Z(n2534) );
  AND U2540 ( .A(g_input[538]), .B(e_input[0]), .Z(n2535) );
  AND U2541 ( .A(g_input[537]), .B(e_input[0]), .Z(n2536) );
  AND U2542 ( .A(g_input[536]), .B(e_input[0]), .Z(n2537) );
  AND U2543 ( .A(g_input[535]), .B(e_input[0]), .Z(n2538) );
  AND U2544 ( .A(g_input[534]), .B(e_input[0]), .Z(n2539) );
  AND U2545 ( .A(g_input[533]), .B(e_input[0]), .Z(n2540) );
  AND U2546 ( .A(g_input[532]), .B(e_input[0]), .Z(n2541) );
  AND U2547 ( .A(g_input[531]), .B(e_input[0]), .Z(n2542) );
  AND U2548 ( .A(g_input[530]), .B(e_input[0]), .Z(n2543) );
  AND U2549 ( .A(g_input[529]), .B(e_input[0]), .Z(n2544) );
  AND U2550 ( .A(g_input[528]), .B(e_input[0]), .Z(n2545) );
  AND U2551 ( .A(g_input[527]), .B(e_input[0]), .Z(n2546) );
  AND U2552 ( .A(g_input[526]), .B(e_input[0]), .Z(n2547) );
  AND U2553 ( .A(g_input[525]), .B(e_input[0]), .Z(n2548) );
  AND U2554 ( .A(g_input[524]), .B(e_input[0]), .Z(n2549) );
  AND U2555 ( .A(g_input[523]), .B(e_input[0]), .Z(n2550) );
  AND U2556 ( .A(g_input[522]), .B(e_input[0]), .Z(n2551) );
  AND U2557 ( .A(g_input[521]), .B(e_input[0]), .Z(n2552) );
  AND U2558 ( .A(g_input[520]), .B(e_input[0]), .Z(n2553) );
  AND U2559 ( .A(g_input[519]), .B(e_input[0]), .Z(n2554) );
  AND U2560 ( .A(g_input[518]), .B(e_input[0]), .Z(n2555) );
  AND U2561 ( .A(g_input[517]), .B(e_input[0]), .Z(n2556) );
  AND U2562 ( .A(g_input[516]), .B(e_input[0]), .Z(n2557) );
  AND U2563 ( .A(g_input[515]), .B(e_input[0]), .Z(n2558) );
  AND U2564 ( .A(g_input[514]), .B(e_input[0]), .Z(n2559) );
  AND U2565 ( .A(g_input[513]), .B(e_input[0]), .Z(n2560) );
  AND U2566 ( .A(g_input[512]), .B(e_input[0]), .Z(n2561) );
  AND U2567 ( .A(g_input[511]), .B(e_input[0]), .Z(n2562) );
  AND U2568 ( .A(g_input[510]), .B(e_input[0]), .Z(n2563) );
  AND U2569 ( .A(g_input[509]), .B(e_input[0]), .Z(n2564) );
  AND U2570 ( .A(g_input[508]), .B(e_input[0]), .Z(n2565) );
  AND U2571 ( .A(g_input[507]), .B(e_input[0]), .Z(n2566) );
  AND U2572 ( .A(g_input[506]), .B(e_input[0]), .Z(n2567) );
  AND U2573 ( .A(g_input[505]), .B(e_input[0]), .Z(n2568) );
  AND U2574 ( .A(g_input[504]), .B(e_input[0]), .Z(n2569) );
  AND U2575 ( .A(g_input[503]), .B(e_input[0]), .Z(n2570) );
  AND U2576 ( .A(g_input[502]), .B(e_input[0]), .Z(n2571) );
  AND U2577 ( .A(g_input[501]), .B(e_input[0]), .Z(n2572) );
  AND U2578 ( .A(g_input[500]), .B(e_input[0]), .Z(n2573) );
  AND U2579 ( .A(g_input[499]), .B(e_input[0]), .Z(n2574) );
  AND U2580 ( .A(g_input[498]), .B(e_input[0]), .Z(n2575) );
  AND U2581 ( .A(g_input[497]), .B(e_input[0]), .Z(n2576) );
  AND U2582 ( .A(g_input[496]), .B(e_input[0]), .Z(n2577) );
  AND U2583 ( .A(g_input[495]), .B(e_input[0]), .Z(n2578) );
  AND U2584 ( .A(g_input[494]), .B(e_input[0]), .Z(n2579) );
  AND U2585 ( .A(g_input[493]), .B(e_input[0]), .Z(n2580) );
  AND U2586 ( .A(g_input[492]), .B(e_input[0]), .Z(n2581) );
  AND U2587 ( .A(g_input[491]), .B(e_input[0]), .Z(n2582) );
  AND U2588 ( .A(g_input[490]), .B(e_input[0]), .Z(n2583) );
  AND U2589 ( .A(g_input[489]), .B(e_input[0]), .Z(n2584) );
  AND U2590 ( .A(g_input[488]), .B(e_input[0]), .Z(n2585) );
  AND U2591 ( .A(g_input[487]), .B(e_input[0]), .Z(n2586) );
  AND U2592 ( .A(g_input[486]), .B(e_input[0]), .Z(n2587) );
  AND U2593 ( .A(g_input[485]), .B(e_input[0]), .Z(n2588) );
  AND U2594 ( .A(g_input[484]), .B(e_input[0]), .Z(n2589) );
  AND U2595 ( .A(g_input[483]), .B(e_input[0]), .Z(n2590) );
  AND U2596 ( .A(g_input[482]), .B(e_input[0]), .Z(n2591) );
  AND U2597 ( .A(g_input[481]), .B(e_input[0]), .Z(n2592) );
  AND U2598 ( .A(g_input[480]), .B(e_input[0]), .Z(n2593) );
  AND U2599 ( .A(g_input[479]), .B(e_input[0]), .Z(n2594) );
  AND U2600 ( .A(g_input[478]), .B(e_input[0]), .Z(n2595) );
  AND U2601 ( .A(g_input[477]), .B(e_input[0]), .Z(n2596) );
  AND U2602 ( .A(g_input[476]), .B(e_input[0]), .Z(n2597) );
  AND U2603 ( .A(g_input[475]), .B(e_input[0]), .Z(n2598) );
  AND U2604 ( .A(g_input[474]), .B(e_input[0]), .Z(n2599) );
  AND U2605 ( .A(g_input[473]), .B(e_input[0]), .Z(n2600) );
  AND U2606 ( .A(g_input[472]), .B(e_input[0]), .Z(n2601) );
  AND U2607 ( .A(g_input[471]), .B(e_input[0]), .Z(n2602) );
  AND U2608 ( .A(g_input[470]), .B(e_input[0]), .Z(n2603) );
  AND U2609 ( .A(g_input[469]), .B(e_input[0]), .Z(n2604) );
  AND U2610 ( .A(g_input[468]), .B(e_input[0]), .Z(n2605) );
  AND U2611 ( .A(g_input[467]), .B(e_input[0]), .Z(n2606) );
  AND U2612 ( .A(g_input[466]), .B(e_input[0]), .Z(n2607) );
  AND U2613 ( .A(g_input[465]), .B(e_input[0]), .Z(n2608) );
  AND U2614 ( .A(g_input[464]), .B(e_input[0]), .Z(n2609) );
  AND U2615 ( .A(g_input[463]), .B(e_input[0]), .Z(n2610) );
  AND U2616 ( .A(g_input[462]), .B(e_input[0]), .Z(n2611) );
  AND U2617 ( .A(g_input[461]), .B(e_input[0]), .Z(n2612) );
  AND U2618 ( .A(g_input[460]), .B(e_input[0]), .Z(n2613) );
  AND U2619 ( .A(g_input[459]), .B(e_input[0]), .Z(n2614) );
  AND U2620 ( .A(g_input[458]), .B(e_input[0]), .Z(n2615) );
  AND U2621 ( .A(g_input[457]), .B(e_input[0]), .Z(n2616) );
  AND U2622 ( .A(g_input[456]), .B(e_input[0]), .Z(n2617) );
  AND U2623 ( .A(g_input[455]), .B(e_input[0]), .Z(n2618) );
  AND U2624 ( .A(g_input[454]), .B(e_input[0]), .Z(n2619) );
  AND U2625 ( .A(g_input[453]), .B(e_input[0]), .Z(n2620) );
  AND U2626 ( .A(g_input[452]), .B(e_input[0]), .Z(n2621) );
  AND U2627 ( .A(g_input[451]), .B(e_input[0]), .Z(n2622) );
  AND U2628 ( .A(g_input[450]), .B(e_input[0]), .Z(n2623) );
  AND U2629 ( .A(g_input[449]), .B(e_input[0]), .Z(n2624) );
  AND U2630 ( .A(g_input[448]), .B(e_input[0]), .Z(n2625) );
  AND U2631 ( .A(g_input[447]), .B(e_input[0]), .Z(n2626) );
  AND U2632 ( .A(g_input[446]), .B(e_input[0]), .Z(n2627) );
  AND U2633 ( .A(g_input[445]), .B(e_input[0]), .Z(n2628) );
  AND U2634 ( .A(g_input[444]), .B(e_input[0]), .Z(n2629) );
  AND U2635 ( .A(g_input[443]), .B(e_input[0]), .Z(n2630) );
  AND U2636 ( .A(g_input[442]), .B(e_input[0]), .Z(n2631) );
  AND U2637 ( .A(g_input[441]), .B(e_input[0]), .Z(n2632) );
  AND U2638 ( .A(g_input[440]), .B(e_input[0]), .Z(n2633) );
  AND U2639 ( .A(g_input[439]), .B(e_input[0]), .Z(n2634) );
  AND U2640 ( .A(g_input[438]), .B(e_input[0]), .Z(n2635) );
  AND U2641 ( .A(g_input[437]), .B(e_input[0]), .Z(n2636) );
  AND U2642 ( .A(g_input[436]), .B(e_input[0]), .Z(n2637) );
  AND U2643 ( .A(g_input[435]), .B(e_input[0]), .Z(n2638) );
  AND U2644 ( .A(g_input[434]), .B(e_input[0]), .Z(n2639) );
  AND U2645 ( .A(g_input[433]), .B(e_input[0]), .Z(n2640) );
  AND U2646 ( .A(g_input[432]), .B(e_input[0]), .Z(n2641) );
  AND U2647 ( .A(g_input[431]), .B(e_input[0]), .Z(n2642) );
  AND U2648 ( .A(g_input[430]), .B(e_input[0]), .Z(n2643) );
  AND U2649 ( .A(g_input[429]), .B(e_input[0]), .Z(n2644) );
  AND U2650 ( .A(g_input[428]), .B(e_input[0]), .Z(n2645) );
  AND U2651 ( .A(g_input[427]), .B(e_input[0]), .Z(n2646) );
  AND U2652 ( .A(g_input[426]), .B(e_input[0]), .Z(n2647) );
  AND U2653 ( .A(g_input[425]), .B(e_input[0]), .Z(n2648) );
  AND U2654 ( .A(g_input[424]), .B(e_input[0]), .Z(n2649) );
  AND U2655 ( .A(g_input[423]), .B(e_input[0]), .Z(n2650) );
  AND U2656 ( .A(g_input[422]), .B(e_input[0]), .Z(n2651) );
  AND U2657 ( .A(g_input[421]), .B(e_input[0]), .Z(n2652) );
  AND U2658 ( .A(g_input[420]), .B(e_input[0]), .Z(n2653) );
  AND U2659 ( .A(g_input[419]), .B(e_input[0]), .Z(n2654) );
  AND U2660 ( .A(g_input[418]), .B(e_input[0]), .Z(n2655) );
  AND U2661 ( .A(g_input[417]), .B(e_input[0]), .Z(n2656) );
  AND U2662 ( .A(g_input[416]), .B(e_input[0]), .Z(n2657) );
  AND U2663 ( .A(g_input[415]), .B(e_input[0]), .Z(n2658) );
  AND U2664 ( .A(g_input[414]), .B(e_input[0]), .Z(n2659) );
  AND U2665 ( .A(g_input[413]), .B(e_input[0]), .Z(n2660) );
  AND U2666 ( .A(g_input[412]), .B(e_input[0]), .Z(n2661) );
  AND U2667 ( .A(g_input[411]), .B(e_input[0]), .Z(n2662) );
  AND U2668 ( .A(g_input[410]), .B(e_input[0]), .Z(n2663) );
  AND U2669 ( .A(g_input[409]), .B(e_input[0]), .Z(n2664) );
  AND U2670 ( .A(g_input[408]), .B(e_input[0]), .Z(n2665) );
  AND U2671 ( .A(g_input[407]), .B(e_input[0]), .Z(n2666) );
  AND U2672 ( .A(g_input[406]), .B(e_input[0]), .Z(n2667) );
  AND U2673 ( .A(g_input[405]), .B(e_input[0]), .Z(n2668) );
  AND U2674 ( .A(g_input[404]), .B(e_input[0]), .Z(n2669) );
  AND U2675 ( .A(g_input[403]), .B(e_input[0]), .Z(n2670) );
  AND U2676 ( .A(g_input[402]), .B(e_input[0]), .Z(n2671) );
  AND U2677 ( .A(g_input[401]), .B(e_input[0]), .Z(n2672) );
  AND U2678 ( .A(g_input[400]), .B(e_input[0]), .Z(n2673) );
  AND U2679 ( .A(g_input[399]), .B(e_input[0]), .Z(n2674) );
  AND U2680 ( .A(g_input[398]), .B(e_input[0]), .Z(n2675) );
  AND U2681 ( .A(g_input[397]), .B(e_input[0]), .Z(n2676) );
  AND U2682 ( .A(g_input[396]), .B(e_input[0]), .Z(n2677) );
  AND U2683 ( .A(g_input[395]), .B(e_input[0]), .Z(n2678) );
  AND U2684 ( .A(g_input[394]), .B(e_input[0]), .Z(n2679) );
  AND U2685 ( .A(g_input[393]), .B(e_input[0]), .Z(n2680) );
  AND U2686 ( .A(g_input[392]), .B(e_input[0]), .Z(n2681) );
  AND U2687 ( .A(g_input[391]), .B(e_input[0]), .Z(n2682) );
  AND U2688 ( .A(g_input[390]), .B(e_input[0]), .Z(n2683) );
  AND U2689 ( .A(g_input[389]), .B(e_input[0]), .Z(n2684) );
  AND U2690 ( .A(g_input[388]), .B(e_input[0]), .Z(n2685) );
  AND U2691 ( .A(g_input[387]), .B(e_input[0]), .Z(n2686) );
  AND U2692 ( .A(g_input[386]), .B(e_input[0]), .Z(n2687) );
  AND U2693 ( .A(g_input[385]), .B(e_input[0]), .Z(n2688) );
  AND U2694 ( .A(g_input[384]), .B(e_input[0]), .Z(n2689) );
  AND U2695 ( .A(g_input[383]), .B(e_input[0]), .Z(n2690) );
  AND U2696 ( .A(g_input[382]), .B(e_input[0]), .Z(n2691) );
  AND U2697 ( .A(g_input[381]), .B(e_input[0]), .Z(n2692) );
  AND U2698 ( .A(g_input[380]), .B(e_input[0]), .Z(n2693) );
  AND U2699 ( .A(g_input[379]), .B(e_input[0]), .Z(n2694) );
  AND U2700 ( .A(g_input[378]), .B(e_input[0]), .Z(n2695) );
  AND U2701 ( .A(g_input[377]), .B(e_input[0]), .Z(n2696) );
  AND U2702 ( .A(g_input[376]), .B(e_input[0]), .Z(n2697) );
  AND U2703 ( .A(g_input[375]), .B(e_input[0]), .Z(n2698) );
  AND U2704 ( .A(g_input[374]), .B(e_input[0]), .Z(n2699) );
  AND U2705 ( .A(g_input[373]), .B(e_input[0]), .Z(n2700) );
  AND U2706 ( .A(g_input[372]), .B(e_input[0]), .Z(n2701) );
  AND U2707 ( .A(g_input[371]), .B(e_input[0]), .Z(n2702) );
  AND U2708 ( .A(g_input[370]), .B(e_input[0]), .Z(n2703) );
  AND U2709 ( .A(g_input[369]), .B(e_input[0]), .Z(n2704) );
  AND U2710 ( .A(g_input[368]), .B(e_input[0]), .Z(n2705) );
  AND U2711 ( .A(g_input[367]), .B(e_input[0]), .Z(n2706) );
  AND U2712 ( .A(g_input[366]), .B(e_input[0]), .Z(n2707) );
  AND U2713 ( .A(g_input[365]), .B(e_input[0]), .Z(n2708) );
  AND U2714 ( .A(g_input[364]), .B(e_input[0]), .Z(n2709) );
  AND U2715 ( .A(g_input[363]), .B(e_input[0]), .Z(n2710) );
  AND U2716 ( .A(g_input[362]), .B(e_input[0]), .Z(n2711) );
  AND U2717 ( .A(g_input[361]), .B(e_input[0]), .Z(n2712) );
  AND U2718 ( .A(g_input[360]), .B(e_input[0]), .Z(n2713) );
  AND U2719 ( .A(g_input[359]), .B(e_input[0]), .Z(n2714) );
  AND U2720 ( .A(g_input[358]), .B(e_input[0]), .Z(n2715) );
  AND U2721 ( .A(g_input[357]), .B(e_input[0]), .Z(n2716) );
  AND U2722 ( .A(g_input[356]), .B(e_input[0]), .Z(n2717) );
  AND U2723 ( .A(g_input[355]), .B(e_input[0]), .Z(n2718) );
  AND U2724 ( .A(g_input[354]), .B(e_input[0]), .Z(n2719) );
  AND U2725 ( .A(g_input[353]), .B(e_input[0]), .Z(n2720) );
  AND U2726 ( .A(g_input[352]), .B(e_input[0]), .Z(n2721) );
  AND U2727 ( .A(g_input[351]), .B(e_input[0]), .Z(n2722) );
  AND U2728 ( .A(g_input[350]), .B(e_input[0]), .Z(n2723) );
  AND U2729 ( .A(g_input[349]), .B(e_input[0]), .Z(n2724) );
  AND U2730 ( .A(g_input[348]), .B(e_input[0]), .Z(n2725) );
  AND U2731 ( .A(g_input[347]), .B(e_input[0]), .Z(n2726) );
  AND U2732 ( .A(g_input[346]), .B(e_input[0]), .Z(n2727) );
  AND U2733 ( .A(g_input[345]), .B(e_input[0]), .Z(n2728) );
  AND U2734 ( .A(g_input[344]), .B(e_input[0]), .Z(n2729) );
  AND U2735 ( .A(g_input[343]), .B(e_input[0]), .Z(n2730) );
  AND U2736 ( .A(g_input[342]), .B(e_input[0]), .Z(n2731) );
  AND U2737 ( .A(g_input[341]), .B(e_input[0]), .Z(n2732) );
  AND U2738 ( .A(g_input[340]), .B(e_input[0]), .Z(n2733) );
  AND U2739 ( .A(g_input[339]), .B(e_input[0]), .Z(n2734) );
  AND U2740 ( .A(g_input[338]), .B(e_input[0]), .Z(n2735) );
  AND U2741 ( .A(g_input[337]), .B(e_input[0]), .Z(n2736) );
  AND U2742 ( .A(g_input[336]), .B(e_input[0]), .Z(n2737) );
  AND U2743 ( .A(g_input[335]), .B(e_input[0]), .Z(n2738) );
  AND U2744 ( .A(g_input[334]), .B(e_input[0]), .Z(n2739) );
  AND U2745 ( .A(g_input[333]), .B(e_input[0]), .Z(n2740) );
  AND U2746 ( .A(g_input[332]), .B(e_input[0]), .Z(n2741) );
  AND U2747 ( .A(g_input[331]), .B(e_input[0]), .Z(n2742) );
  AND U2748 ( .A(g_input[330]), .B(e_input[0]), .Z(n2743) );
  AND U2749 ( .A(g_input[329]), .B(e_input[0]), .Z(n2744) );
  AND U2750 ( .A(g_input[328]), .B(e_input[0]), .Z(n2745) );
  AND U2751 ( .A(g_input[327]), .B(e_input[0]), .Z(n2746) );
  AND U2752 ( .A(g_input[326]), .B(e_input[0]), .Z(n2747) );
  AND U2753 ( .A(g_input[325]), .B(e_input[0]), .Z(n2748) );
  AND U2754 ( .A(g_input[324]), .B(e_input[0]), .Z(n2749) );
  AND U2755 ( .A(g_input[323]), .B(e_input[0]), .Z(n2750) );
  AND U2756 ( .A(g_input[322]), .B(e_input[0]), .Z(n2751) );
  AND U2757 ( .A(g_input[321]), .B(e_input[0]), .Z(n2752) );
  AND U2758 ( .A(g_input[320]), .B(e_input[0]), .Z(n2753) );
  AND U2759 ( .A(g_input[319]), .B(e_input[0]), .Z(n2754) );
  AND U2760 ( .A(g_input[318]), .B(e_input[0]), .Z(n2755) );
  AND U2761 ( .A(g_input[317]), .B(e_input[0]), .Z(n2756) );
  AND U2762 ( .A(g_input[316]), .B(e_input[0]), .Z(n2757) );
  AND U2763 ( .A(g_input[315]), .B(e_input[0]), .Z(n2758) );
  AND U2764 ( .A(g_input[314]), .B(e_input[0]), .Z(n2759) );
  AND U2765 ( .A(g_input[313]), .B(e_input[0]), .Z(n2760) );
  AND U2766 ( .A(g_input[312]), .B(e_input[0]), .Z(n2761) );
  AND U2767 ( .A(g_input[311]), .B(e_input[0]), .Z(n2762) );
  AND U2768 ( .A(g_input[310]), .B(e_input[0]), .Z(n2763) );
  AND U2769 ( .A(g_input[309]), .B(e_input[0]), .Z(n2764) );
  AND U2770 ( .A(g_input[308]), .B(e_input[0]), .Z(n2765) );
  AND U2771 ( .A(g_input[307]), .B(e_input[0]), .Z(n2766) );
  AND U2772 ( .A(g_input[306]), .B(e_input[0]), .Z(n2767) );
  AND U2773 ( .A(g_input[305]), .B(e_input[0]), .Z(n2768) );
  AND U2774 ( .A(g_input[304]), .B(e_input[0]), .Z(n2769) );
  AND U2775 ( .A(g_input[303]), .B(e_input[0]), .Z(n2770) );
  AND U2776 ( .A(g_input[302]), .B(e_input[0]), .Z(n2771) );
  AND U2777 ( .A(g_input[301]), .B(e_input[0]), .Z(n2772) );
  AND U2778 ( .A(g_input[300]), .B(e_input[0]), .Z(n2773) );
  AND U2779 ( .A(g_input[299]), .B(e_input[0]), .Z(n2774) );
  AND U2780 ( .A(g_input[298]), .B(e_input[0]), .Z(n2775) );
  AND U2781 ( .A(g_input[297]), .B(e_input[0]), .Z(n2776) );
  AND U2782 ( .A(g_input[296]), .B(e_input[0]), .Z(n2777) );
  AND U2783 ( .A(g_input[295]), .B(e_input[0]), .Z(n2778) );
  AND U2784 ( .A(g_input[294]), .B(e_input[0]), .Z(n2779) );
  AND U2785 ( .A(g_input[293]), .B(e_input[0]), .Z(n2780) );
  AND U2786 ( .A(g_input[292]), .B(e_input[0]), .Z(n2781) );
  AND U2787 ( .A(g_input[291]), .B(e_input[0]), .Z(n2782) );
  AND U2788 ( .A(g_input[290]), .B(e_input[0]), .Z(n2783) );
  AND U2789 ( .A(g_input[289]), .B(e_input[0]), .Z(n2784) );
  AND U2790 ( .A(g_input[288]), .B(e_input[0]), .Z(n2785) );
  AND U2791 ( .A(g_input[287]), .B(e_input[0]), .Z(n2786) );
  AND U2792 ( .A(g_input[286]), .B(e_input[0]), .Z(n2787) );
  AND U2793 ( .A(g_input[285]), .B(e_input[0]), .Z(n2788) );
  AND U2794 ( .A(g_input[284]), .B(e_input[0]), .Z(n2789) );
  AND U2795 ( .A(g_input[283]), .B(e_input[0]), .Z(n2790) );
  AND U2796 ( .A(g_input[282]), .B(e_input[0]), .Z(n2791) );
  AND U2797 ( .A(g_input[281]), .B(e_input[0]), .Z(n2792) );
  AND U2798 ( .A(g_input[280]), .B(e_input[0]), .Z(n2793) );
  AND U2799 ( .A(g_input[279]), .B(e_input[0]), .Z(n2794) );
  AND U2800 ( .A(g_input[278]), .B(e_input[0]), .Z(n2795) );
  AND U2801 ( .A(g_input[277]), .B(e_input[0]), .Z(n2796) );
  AND U2802 ( .A(g_input[276]), .B(e_input[0]), .Z(n2797) );
  AND U2803 ( .A(g_input[275]), .B(e_input[0]), .Z(n2798) );
  AND U2804 ( .A(g_input[274]), .B(e_input[0]), .Z(n2799) );
  AND U2805 ( .A(g_input[273]), .B(e_input[0]), .Z(n2800) );
  AND U2806 ( .A(g_input[272]), .B(e_input[0]), .Z(n2801) );
  AND U2807 ( .A(g_input[271]), .B(e_input[0]), .Z(n2802) );
  AND U2808 ( .A(g_input[270]), .B(e_input[0]), .Z(n2803) );
  AND U2809 ( .A(g_input[269]), .B(e_input[0]), .Z(n2804) );
  AND U2810 ( .A(g_input[268]), .B(e_input[0]), .Z(n2805) );
  AND U2811 ( .A(g_input[267]), .B(e_input[0]), .Z(n2806) );
  AND U2812 ( .A(g_input[266]), .B(e_input[0]), .Z(n2807) );
  AND U2813 ( .A(g_input[265]), .B(e_input[0]), .Z(n2808) );
  AND U2814 ( .A(g_input[264]), .B(e_input[0]), .Z(n2809) );
  AND U2815 ( .A(g_input[263]), .B(e_input[0]), .Z(n2810) );
  AND U2816 ( .A(g_input[262]), .B(e_input[0]), .Z(n2811) );
  AND U2817 ( .A(g_input[261]), .B(e_input[0]), .Z(n2812) );
  AND U2818 ( .A(g_input[260]), .B(e_input[0]), .Z(n2813) );
  AND U2819 ( .A(g_input[259]), .B(e_input[0]), .Z(n2814) );
  AND U2820 ( .A(g_input[258]), .B(e_input[0]), .Z(n2815) );
  AND U2821 ( .A(g_input[257]), .B(e_input[0]), .Z(n2816) );
  AND U2822 ( .A(g_input[256]), .B(e_input[0]), .Z(n2817) );
  AND U2823 ( .A(g_input[255]), .B(e_input[0]), .Z(n2818) );
  AND U2824 ( .A(g_input[254]), .B(e_input[0]), .Z(n2819) );
  AND U2825 ( .A(g_input[253]), .B(e_input[0]), .Z(n2820) );
  AND U2826 ( .A(g_input[252]), .B(e_input[0]), .Z(n2821) );
  AND U2827 ( .A(g_input[251]), .B(e_input[0]), .Z(n2822) );
  AND U2828 ( .A(g_input[250]), .B(e_input[0]), .Z(n2823) );
  AND U2829 ( .A(g_input[249]), .B(e_input[0]), .Z(n2824) );
  AND U2830 ( .A(g_input[248]), .B(e_input[0]), .Z(n2825) );
  AND U2831 ( .A(g_input[247]), .B(e_input[0]), .Z(n2826) );
  AND U2832 ( .A(g_input[246]), .B(e_input[0]), .Z(n2827) );
  AND U2833 ( .A(g_input[245]), .B(e_input[0]), .Z(n2828) );
  AND U2834 ( .A(g_input[244]), .B(e_input[0]), .Z(n2829) );
  AND U2835 ( .A(g_input[243]), .B(e_input[0]), .Z(n2830) );
  AND U2836 ( .A(g_input[242]), .B(e_input[0]), .Z(n2831) );
  AND U2837 ( .A(g_input[241]), .B(e_input[0]), .Z(n2832) );
  AND U2838 ( .A(g_input[240]), .B(e_input[0]), .Z(n2833) );
  AND U2839 ( .A(g_input[239]), .B(e_input[0]), .Z(n2834) );
  AND U2840 ( .A(g_input[238]), .B(e_input[0]), .Z(n2835) );
  AND U2841 ( .A(g_input[237]), .B(e_input[0]), .Z(n2836) );
  AND U2842 ( .A(g_input[236]), .B(e_input[0]), .Z(n2837) );
  AND U2843 ( .A(g_input[235]), .B(e_input[0]), .Z(n2838) );
  AND U2844 ( .A(g_input[234]), .B(e_input[0]), .Z(n2839) );
  AND U2845 ( .A(g_input[233]), .B(e_input[0]), .Z(n2840) );
  AND U2846 ( .A(g_input[232]), .B(e_input[0]), .Z(n2841) );
  AND U2847 ( .A(g_input[231]), .B(e_input[0]), .Z(n2842) );
  AND U2848 ( .A(g_input[230]), .B(e_input[0]), .Z(n2843) );
  AND U2849 ( .A(g_input[229]), .B(e_input[0]), .Z(n2844) );
  AND U2850 ( .A(g_input[228]), .B(e_input[0]), .Z(n2845) );
  AND U2851 ( .A(g_input[227]), .B(e_input[0]), .Z(n2846) );
  AND U2852 ( .A(g_input[226]), .B(e_input[0]), .Z(n2847) );
  AND U2853 ( .A(g_input[225]), .B(e_input[0]), .Z(n2848) );
  AND U2854 ( .A(g_input[224]), .B(e_input[0]), .Z(n2849) );
  AND U2855 ( .A(g_input[223]), .B(e_input[0]), .Z(n2850) );
  AND U2856 ( .A(g_input[222]), .B(e_input[0]), .Z(n2851) );
  AND U2857 ( .A(g_input[221]), .B(e_input[0]), .Z(n2852) );
  AND U2858 ( .A(g_input[220]), .B(e_input[0]), .Z(n2853) );
  AND U2859 ( .A(g_input[219]), .B(e_input[0]), .Z(n2854) );
  AND U2860 ( .A(g_input[218]), .B(e_input[0]), .Z(n2855) );
  AND U2861 ( .A(g_input[217]), .B(e_input[0]), .Z(n2856) );
  AND U2862 ( .A(g_input[216]), .B(e_input[0]), .Z(n2857) );
  AND U2863 ( .A(g_input[215]), .B(e_input[0]), .Z(n2858) );
  AND U2864 ( .A(g_input[214]), .B(e_input[0]), .Z(n2859) );
  AND U2865 ( .A(g_input[213]), .B(e_input[0]), .Z(n2860) );
  AND U2866 ( .A(g_input[212]), .B(e_input[0]), .Z(n2861) );
  AND U2867 ( .A(g_input[211]), .B(e_input[0]), .Z(n2862) );
  AND U2868 ( .A(g_input[210]), .B(e_input[0]), .Z(n2863) );
  AND U2869 ( .A(g_input[209]), .B(e_input[0]), .Z(n2864) );
  AND U2870 ( .A(g_input[208]), .B(e_input[0]), .Z(n2865) );
  AND U2871 ( .A(g_input[207]), .B(e_input[0]), .Z(n2866) );
  AND U2872 ( .A(g_input[206]), .B(e_input[0]), .Z(n2867) );
  AND U2873 ( .A(g_input[205]), .B(e_input[0]), .Z(n2868) );
  AND U2874 ( .A(g_input[204]), .B(e_input[0]), .Z(n2869) );
  AND U2875 ( .A(g_input[203]), .B(e_input[0]), .Z(n2870) );
  AND U2876 ( .A(g_input[202]), .B(e_input[0]), .Z(n2871) );
  AND U2877 ( .A(g_input[201]), .B(e_input[0]), .Z(n2872) );
  AND U2878 ( .A(g_input[200]), .B(e_input[0]), .Z(n2873) );
  AND U2879 ( .A(g_input[199]), .B(e_input[0]), .Z(n2874) );
  AND U2880 ( .A(g_input[198]), .B(e_input[0]), .Z(n2875) );
  AND U2881 ( .A(g_input[197]), .B(e_input[0]), .Z(n2876) );
  AND U2882 ( .A(g_input[196]), .B(e_input[0]), .Z(n2877) );
  AND U2883 ( .A(g_input[195]), .B(e_input[0]), .Z(n2878) );
  AND U2884 ( .A(g_input[194]), .B(e_input[0]), .Z(n2879) );
  AND U2885 ( .A(g_input[193]), .B(e_input[0]), .Z(n2880) );
  AND U2886 ( .A(g_input[192]), .B(e_input[0]), .Z(n2881) );
  AND U2887 ( .A(g_input[191]), .B(e_input[0]), .Z(n2882) );
  AND U2888 ( .A(g_input[190]), .B(e_input[0]), .Z(n2883) );
  AND U2889 ( .A(g_input[189]), .B(e_input[0]), .Z(n2884) );
  AND U2890 ( .A(g_input[188]), .B(e_input[0]), .Z(n2885) );
  AND U2891 ( .A(g_input[187]), .B(e_input[0]), .Z(n2886) );
  AND U2892 ( .A(g_input[186]), .B(e_input[0]), .Z(n2887) );
  AND U2893 ( .A(g_input[185]), .B(e_input[0]), .Z(n2888) );
  AND U2894 ( .A(g_input[184]), .B(e_input[0]), .Z(n2889) );
  AND U2895 ( .A(g_input[183]), .B(e_input[0]), .Z(n2890) );
  AND U2896 ( .A(g_input[182]), .B(e_input[0]), .Z(n2891) );
  AND U2897 ( .A(g_input[181]), .B(e_input[0]), .Z(n2892) );
  AND U2898 ( .A(g_input[180]), .B(e_input[0]), .Z(n2893) );
  AND U2899 ( .A(g_input[179]), .B(e_input[0]), .Z(n2894) );
  AND U2900 ( .A(g_input[178]), .B(e_input[0]), .Z(n2895) );
  AND U2901 ( .A(g_input[177]), .B(e_input[0]), .Z(n2896) );
  AND U2902 ( .A(g_input[176]), .B(e_input[0]), .Z(n2897) );
  AND U2903 ( .A(g_input[175]), .B(e_input[0]), .Z(n2898) );
  AND U2904 ( .A(g_input[174]), .B(e_input[0]), .Z(n2899) );
  AND U2905 ( .A(g_input[173]), .B(e_input[0]), .Z(n2900) );
  AND U2906 ( .A(g_input[172]), .B(e_input[0]), .Z(n2901) );
  AND U2907 ( .A(g_input[171]), .B(e_input[0]), .Z(n2902) );
  AND U2908 ( .A(g_input[170]), .B(e_input[0]), .Z(n2903) );
  AND U2909 ( .A(g_input[169]), .B(e_input[0]), .Z(n2904) );
  AND U2910 ( .A(g_input[168]), .B(e_input[0]), .Z(n2905) );
  AND U2911 ( .A(g_input[167]), .B(e_input[0]), .Z(n2906) );
  AND U2912 ( .A(g_input[166]), .B(e_input[0]), .Z(n2907) );
  AND U2913 ( .A(g_input[165]), .B(e_input[0]), .Z(n2908) );
  AND U2914 ( .A(g_input[164]), .B(e_input[0]), .Z(n2909) );
  AND U2915 ( .A(g_input[163]), .B(e_input[0]), .Z(n2910) );
  AND U2916 ( .A(g_input[162]), .B(e_input[0]), .Z(n2911) );
  AND U2917 ( .A(g_input[161]), .B(e_input[0]), .Z(n2912) );
  AND U2918 ( .A(g_input[160]), .B(e_input[0]), .Z(n2913) );
  AND U2919 ( .A(g_input[159]), .B(e_input[0]), .Z(n2914) );
  AND U2920 ( .A(g_input[158]), .B(e_input[0]), .Z(n2915) );
  AND U2921 ( .A(g_input[157]), .B(e_input[0]), .Z(n2916) );
  AND U2922 ( .A(g_input[156]), .B(e_input[0]), .Z(n2917) );
  AND U2923 ( .A(g_input[155]), .B(e_input[0]), .Z(n2918) );
  AND U2924 ( .A(g_input[154]), .B(e_input[0]), .Z(n2919) );
  AND U2925 ( .A(g_input[153]), .B(e_input[0]), .Z(n2920) );
  AND U2926 ( .A(g_input[152]), .B(e_input[0]), .Z(n2921) );
  AND U2927 ( .A(g_input[151]), .B(e_input[0]), .Z(n2922) );
  AND U2928 ( .A(g_input[150]), .B(e_input[0]), .Z(n2923) );
  AND U2929 ( .A(g_input[149]), .B(e_input[0]), .Z(n2924) );
  AND U2930 ( .A(g_input[148]), .B(e_input[0]), .Z(n2925) );
  AND U2931 ( .A(g_input[147]), .B(e_input[0]), .Z(n2926) );
  AND U2932 ( .A(g_input[146]), .B(e_input[0]), .Z(n2927) );
  AND U2933 ( .A(g_input[145]), .B(e_input[0]), .Z(n2928) );
  AND U2934 ( .A(g_input[144]), .B(e_input[0]), .Z(n2929) );
  AND U2935 ( .A(g_input[143]), .B(e_input[0]), .Z(n2930) );
  AND U2936 ( .A(g_input[142]), .B(e_input[0]), .Z(n2931) );
  AND U2937 ( .A(g_input[141]), .B(e_input[0]), .Z(n2932) );
  AND U2938 ( .A(g_input[140]), .B(e_input[0]), .Z(n2933) );
  AND U2939 ( .A(g_input[139]), .B(e_input[0]), .Z(n2934) );
  AND U2940 ( .A(g_input[138]), .B(e_input[0]), .Z(n2935) );
  AND U2941 ( .A(g_input[137]), .B(e_input[0]), .Z(n2936) );
  AND U2942 ( .A(g_input[136]), .B(e_input[0]), .Z(n2937) );
  AND U2943 ( .A(g_input[135]), .B(e_input[0]), .Z(n2938) );
  AND U2944 ( .A(g_input[134]), .B(e_input[0]), .Z(n2939) );
  AND U2945 ( .A(g_input[133]), .B(e_input[0]), .Z(n2940) );
  AND U2946 ( .A(g_input[132]), .B(e_input[0]), .Z(n2941) );
  AND U2947 ( .A(g_input[131]), .B(e_input[0]), .Z(n2942) );
  AND U2948 ( .A(g_input[130]), .B(e_input[0]), .Z(n2943) );
  AND U2949 ( .A(g_input[129]), .B(e_input[0]), .Z(n2944) );
  AND U2950 ( .A(g_input[128]), .B(e_input[0]), .Z(n2945) );
  AND U2951 ( .A(g_input[127]), .B(e_input[0]), .Z(n2946) );
  AND U2952 ( .A(g_input[126]), .B(e_input[0]), .Z(n2947) );
  AND U2953 ( .A(g_input[125]), .B(e_input[0]), .Z(n2948) );
  AND U2954 ( .A(g_input[124]), .B(e_input[0]), .Z(n2949) );
  AND U2955 ( .A(g_input[123]), .B(e_input[0]), .Z(n2950) );
  AND U2956 ( .A(g_input[122]), .B(e_input[0]), .Z(n2951) );
  AND U2957 ( .A(g_input[121]), .B(e_input[0]), .Z(n2952) );
  AND U2958 ( .A(g_input[120]), .B(e_input[0]), .Z(n2953) );
  AND U2959 ( .A(g_input[119]), .B(e_input[0]), .Z(n2954) );
  AND U2960 ( .A(g_input[118]), .B(e_input[0]), .Z(n2955) );
  AND U2961 ( .A(g_input[117]), .B(e_input[0]), .Z(n2956) );
  AND U2962 ( .A(g_input[116]), .B(e_input[0]), .Z(n2957) );
  AND U2963 ( .A(g_input[115]), .B(e_input[0]), .Z(n2958) );
  AND U2964 ( .A(g_input[114]), .B(e_input[0]), .Z(n2959) );
  AND U2965 ( .A(g_input[113]), .B(e_input[0]), .Z(n2960) );
  AND U2966 ( .A(g_input[112]), .B(e_input[0]), .Z(n2961) );
  AND U2967 ( .A(g_input[111]), .B(e_input[0]), .Z(n2962) );
  AND U2968 ( .A(g_input[110]), .B(e_input[0]), .Z(n2963) );
  AND U2969 ( .A(g_input[109]), .B(e_input[0]), .Z(n2964) );
  AND U2970 ( .A(g_input[108]), .B(e_input[0]), .Z(n2965) );
  AND U2971 ( .A(g_input[107]), .B(e_input[0]), .Z(n2966) );
  AND U2972 ( .A(g_input[106]), .B(e_input[0]), .Z(n2967) );
  AND U2973 ( .A(g_input[105]), .B(e_input[0]), .Z(n2968) );
  AND U2974 ( .A(g_input[104]), .B(e_input[0]), .Z(n2969) );
  AND U2975 ( .A(g_input[103]), .B(e_input[0]), .Z(n2970) );
  AND U2976 ( .A(g_input[102]), .B(e_input[0]), .Z(n2971) );
  AND U2977 ( .A(g_input[101]), .B(e_input[0]), .Z(n2972) );
  AND U2978 ( .A(g_input[100]), .B(e_input[0]), .Z(n2973) );
  AND U2979 ( .A(g_input[99]), .B(e_input[0]), .Z(n2974) );
  AND U2980 ( .A(g_input[98]), .B(e_input[0]), .Z(n2975) );
  AND U2981 ( .A(g_input[97]), .B(e_input[0]), .Z(n2976) );
  AND U2982 ( .A(g_input[96]), .B(e_input[0]), .Z(n2977) );
  AND U2983 ( .A(g_input[95]), .B(e_input[0]), .Z(n2978) );
  AND U2984 ( .A(g_input[94]), .B(e_input[0]), .Z(n2979) );
  AND U2985 ( .A(g_input[93]), .B(e_input[0]), .Z(n2980) );
  AND U2986 ( .A(g_input[92]), .B(e_input[0]), .Z(n2981) );
  AND U2987 ( .A(g_input[91]), .B(e_input[0]), .Z(n2982) );
  AND U2988 ( .A(g_input[90]), .B(e_input[0]), .Z(n2983) );
  AND U2989 ( .A(g_input[89]), .B(e_input[0]), .Z(n2984) );
  AND U2990 ( .A(g_input[88]), .B(e_input[0]), .Z(n2985) );
  AND U2991 ( .A(g_input[87]), .B(e_input[0]), .Z(n2986) );
  AND U2992 ( .A(g_input[86]), .B(e_input[0]), .Z(n2987) );
  AND U2993 ( .A(g_input[85]), .B(e_input[0]), .Z(n2988) );
  AND U2994 ( .A(g_input[84]), .B(e_input[0]), .Z(n2989) );
  AND U2995 ( .A(g_input[83]), .B(e_input[0]), .Z(n2990) );
  AND U2996 ( .A(g_input[82]), .B(e_input[0]), .Z(n2991) );
  AND U2997 ( .A(g_input[81]), .B(e_input[0]), .Z(n2992) );
  AND U2998 ( .A(g_input[80]), .B(e_input[0]), .Z(n2993) );
  AND U2999 ( .A(g_input[79]), .B(e_input[0]), .Z(n2994) );
  AND U3000 ( .A(g_input[78]), .B(e_input[0]), .Z(n2995) );
  AND U3001 ( .A(g_input[77]), .B(e_input[0]), .Z(n2996) );
  AND U3002 ( .A(g_input[76]), .B(e_input[0]), .Z(n2997) );
  AND U3003 ( .A(g_input[75]), .B(e_input[0]), .Z(n2998) );
  AND U3004 ( .A(g_input[74]), .B(e_input[0]), .Z(n2999) );
  AND U3005 ( .A(g_input[73]), .B(e_input[0]), .Z(n3000) );
  AND U3006 ( .A(g_input[72]), .B(e_input[0]), .Z(n3001) );
  AND U3007 ( .A(g_input[71]), .B(e_input[0]), .Z(n3002) );
  AND U3008 ( .A(g_input[70]), .B(e_input[0]), .Z(n3003) );
  AND U3009 ( .A(g_input[69]), .B(e_input[0]), .Z(n3004) );
  AND U3010 ( .A(g_input[68]), .B(e_input[0]), .Z(n3005) );
  AND U3011 ( .A(g_input[67]), .B(e_input[0]), .Z(n3006) );
  AND U3012 ( .A(g_input[66]), .B(e_input[0]), .Z(n3007) );
  AND U3013 ( .A(g_input[65]), .B(e_input[0]), .Z(n3008) );
  AND U3014 ( .A(g_input[64]), .B(e_input[0]), .Z(n3009) );
  AND U3015 ( .A(g_input[63]), .B(e_input[0]), .Z(n3010) );
  AND U3016 ( .A(g_input[62]), .B(e_input[0]), .Z(n3011) );
  AND U3017 ( .A(g_input[61]), .B(e_input[0]), .Z(n3012) );
  AND U3018 ( .A(g_input[60]), .B(e_input[0]), .Z(n3013) );
  AND U3019 ( .A(g_input[59]), .B(e_input[0]), .Z(n3014) );
  AND U3020 ( .A(g_input[58]), .B(e_input[0]), .Z(n3015) );
  AND U3021 ( .A(g_input[57]), .B(e_input[0]), .Z(n3016) );
  AND U3022 ( .A(g_input[56]), .B(e_input[0]), .Z(n3017) );
  AND U3023 ( .A(g_input[55]), .B(e_input[0]), .Z(n3018) );
  AND U3024 ( .A(g_input[54]), .B(e_input[0]), .Z(n3019) );
  AND U3025 ( .A(g_input[53]), .B(e_input[0]), .Z(n3020) );
  AND U3026 ( .A(g_input[52]), .B(e_input[0]), .Z(n3021) );
  AND U3027 ( .A(g_input[51]), .B(e_input[0]), .Z(n3022) );
  AND U3028 ( .A(g_input[50]), .B(e_input[0]), .Z(n3023) );
  AND U3029 ( .A(g_input[49]), .B(e_input[0]), .Z(n3024) );
  AND U3030 ( .A(g_input[48]), .B(e_input[0]), .Z(n3025) );
  AND U3031 ( .A(g_input[47]), .B(e_input[0]), .Z(n3026) );
  AND U3032 ( .A(g_input[46]), .B(e_input[0]), .Z(n3027) );
  AND U3033 ( .A(g_input[45]), .B(e_input[0]), .Z(n3028) );
  AND U3034 ( .A(g_input[44]), .B(e_input[0]), .Z(n3029) );
  AND U3035 ( .A(g_input[43]), .B(e_input[0]), .Z(n3030) );
  AND U3036 ( .A(g_input[42]), .B(e_input[0]), .Z(n3031) );
  AND U3037 ( .A(g_input[41]), .B(e_input[0]), .Z(n3032) );
  AND U3038 ( .A(g_input[40]), .B(e_input[0]), .Z(n3033) );
  AND U3039 ( .A(g_input[39]), .B(e_input[0]), .Z(n3034) );
  AND U3040 ( .A(g_input[38]), .B(e_input[0]), .Z(n3035) );
  AND U3041 ( .A(g_input[37]), .B(e_input[0]), .Z(n3036) );
  AND U3042 ( .A(g_input[36]), .B(e_input[0]), .Z(n3037) );
  AND U3043 ( .A(g_input[35]), .B(e_input[0]), .Z(n3038) );
  AND U3044 ( .A(g_input[34]), .B(e_input[0]), .Z(n3039) );
  AND U3045 ( .A(g_input[33]), .B(e_input[0]), .Z(n3040) );
  AND U3046 ( .A(g_input[32]), .B(e_input[0]), .Z(n3041) );
  AND U3047 ( .A(g_input[31]), .B(e_input[0]), .Z(n3042) );
  AND U3048 ( .A(g_input[30]), .B(e_input[0]), .Z(n3043) );
  AND U3049 ( .A(g_input[29]), .B(e_input[0]), .Z(n3044) );
  AND U3050 ( .A(g_input[28]), .B(e_input[0]), .Z(n3045) );
  AND U3051 ( .A(g_input[27]), .B(e_input[0]), .Z(n3046) );
  AND U3052 ( .A(g_input[26]), .B(e_input[0]), .Z(n3047) );
  AND U3053 ( .A(g_input[25]), .B(e_input[0]), .Z(n3048) );
  AND U3054 ( .A(g_input[24]), .B(e_input[0]), .Z(n3049) );
  AND U3055 ( .A(g_input[23]), .B(e_input[0]), .Z(n3050) );
  AND U3056 ( .A(g_input[22]), .B(e_input[0]), .Z(n3051) );
  AND U3057 ( .A(g_input[21]), .B(e_input[0]), .Z(n3052) );
  AND U3058 ( .A(g_input[20]), .B(e_input[0]), .Z(n3053) );
  AND U3059 ( .A(g_input[19]), .B(e_input[0]), .Z(n3054) );
  AND U3060 ( .A(g_input[18]), .B(e_input[0]), .Z(n3055) );
  AND U3061 ( .A(g_input[17]), .B(e_input[0]), .Z(n3056) );
  AND U3062 ( .A(g_input[16]), .B(e_input[0]), .Z(n3057) );
  AND U3063 ( .A(g_input[15]), .B(e_input[0]), .Z(n3058) );
  AND U3064 ( .A(g_input[14]), .B(e_input[0]), .Z(n3059) );
  AND U3065 ( .A(g_input[13]), .B(e_input[0]), .Z(n3060) );
  AND U3066 ( .A(g_input[12]), .B(e_input[0]), .Z(n3061) );
  AND U3067 ( .A(g_input[11]), .B(e_input[0]), .Z(n3062) );
  AND U3068 ( .A(g_input[10]), .B(e_input[0]), .Z(n3063) );
  AND U3069 ( .A(g_input[9]), .B(e_input[0]), .Z(n3064) );
  AND U3070 ( .A(g_input[8]), .B(e_input[0]), .Z(n3065) );
  AND U3071 ( .A(g_input[7]), .B(e_input[0]), .Z(n3066) );
  AND U3072 ( .A(g_input[6]), .B(e_input[0]), .Z(n3067) );
  AND U3073 ( .A(g_input[5]), .B(e_input[0]), .Z(n3068) );
  AND U3074 ( .A(g_input[4]), .B(e_input[0]), .Z(n3069) );
  AND U3075 ( .A(g_input[3]), .B(e_input[0]), .Z(n3070) );
  AND U3076 ( .A(g_input[2]), .B(e_input[0]), .Z(n3071) );
  AND U3077 ( .A(g_input[1]), .B(e_input[0]), .Z(n3072) );
  AND U3078 ( .A(g_input[0]), .B(e_input[0]), .Z(n3073) );
endmodule

