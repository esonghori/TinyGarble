
module matrix_mult_N_M_3_N8_M32 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507;
  wire   [31:0] oi;

  DFF \o_reg[0]  ( .D(oi[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[0]) );
  DFF \o_reg[1]  ( .D(oi[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[1]) );
  DFF \o_reg[2]  ( .D(oi[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[2]) );
  DFF \o_reg[3]  ( .D(oi[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[3]) );
  DFF \o_reg[4]  ( .D(oi[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[4]) );
  DFF \o_reg[5]  ( .D(oi[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[5]) );
  DFF \o_reg[6]  ( .D(oi[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[6]) );
  DFF \o_reg[7]  ( .D(oi[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[7]) );
  DFF \o_reg[8]  ( .D(oi[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[8]) );
  DFF \o_reg[9]  ( .D(oi[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[9]) );
  DFF \o_reg[10]  ( .D(oi[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[10]) );
  DFF \o_reg[11]  ( .D(oi[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[11]) );
  DFF \o_reg[12]  ( .D(oi[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[12]) );
  DFF \o_reg[13]  ( .D(oi[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[13]) );
  DFF \o_reg[14]  ( .D(oi[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[14]) );
  DFF \o_reg[15]  ( .D(oi[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[15]) );
  DFF \o_reg[16]  ( .D(oi[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[16]) );
  DFF \o_reg[17]  ( .D(oi[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[17]) );
  DFF \o_reg[18]  ( .D(oi[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[18]) );
  DFF \o_reg[19]  ( .D(oi[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[19]) );
  DFF \o_reg[20]  ( .D(oi[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[20]) );
  DFF \o_reg[21]  ( .D(oi[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[21]) );
  DFF \o_reg[22]  ( .D(oi[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[22]) );
  DFF \o_reg[23]  ( .D(oi[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[23]) );
  DFF \o_reg[24]  ( .D(oi[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[24]) );
  DFF \o_reg[25]  ( .D(oi[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[25]) );
  DFF \o_reg[26]  ( .D(oi[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[26]) );
  DFF \o_reg[27]  ( .D(oi[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[27]) );
  DFF \o_reg[28]  ( .D(oi[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[28]) );
  DFF \o_reg[29]  ( .D(oi[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[29]) );
  DFF \o_reg[30]  ( .D(oi[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[30]) );
  DFF \o_reg[31]  ( .D(oi[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[31]) );
  MUX U35 ( .IN0(n33), .IN1(n1526), .SEL(n1527), .F(n1434) );
  IV U36 ( .A(n1528), .Z(n33) );
  MUX U37 ( .IN0(n1512), .IN1(n34), .SEL(n1513), .F(n1422) );
  IV U38 ( .A(n1514), .Z(n34) );
  MUX U39 ( .IN0(n1504), .IN1(n35), .SEL(n1505), .F(n1410) );
  IV U40 ( .A(n1506), .Z(n35) );
  XNOR U41 ( .A(n892), .B(n891), .Z(n888) );
  MUX U42 ( .IN0(n1298), .IN1(n36), .SEL(n1299), .F(n1196) );
  IV U43 ( .A(n1300), .Z(n36) );
  MUX U44 ( .IN0(n995), .IN1(n37), .SEL(n996), .F(n882) );
  IV U45 ( .A(n997), .Z(n37) );
  XNOR U46 ( .A(n876), .B(n875), .Z(n872) );
  MUX U47 ( .IN0(n979), .IN1(n38), .SEL(n980), .F(n866) );
  IV U48 ( .A(n981), .Z(n38) );
  MUX U49 ( .IN0(n1380), .IN1(n39), .SEL(n1381), .F(n1284) );
  IV U50 ( .A(n1382), .Z(n39) );
  XNOR U51 ( .A(n860), .B(n859), .Z(n856) );
  MUX U52 ( .IN0(n963), .IN1(n40), .SEL(n964), .F(n850) );
  IV U53 ( .A(n965), .Z(n40) );
  XNOR U54 ( .A(n844), .B(n843), .Z(n840) );
  MUX U55 ( .IN0(n1162), .IN1(n41), .SEL(n1163), .F(n1052) );
  IV U56 ( .A(n1164), .Z(n41) );
  MUX U57 ( .IN0(n947), .IN1(n42), .SEL(n948), .F(n834) );
  IV U58 ( .A(n949), .Z(n42) );
  MUX U59 ( .IN0(n1044), .IN1(n43), .SEL(n1045), .F(n934) );
  IV U60 ( .A(n1046), .Z(n43) );
  MUX U61 ( .IN0(n44), .IN1(n2431), .SEL(n2406), .F(n2288) );
  IV U62 ( .A(n2405), .Z(n44) );
  XNOR U63 ( .A(n820), .B(n819), .Z(n816) );
  MUX U64 ( .IN0(n922), .IN1(n45), .SEL(n923), .F(n810) );
  IV U65 ( .A(n924), .Z(n45) );
  MUX U66 ( .IN0(n2360), .IN1(n2362), .SEL(n2361), .F(n2276) );
  MUX U67 ( .IN0(n2413), .IN1(n2415), .SEL(n2414), .F(n2407) );
  MUX U68 ( .IN0(n46), .IN1(n2447), .SEL(n2426), .F(n2443) );
  IV U69 ( .A(n2425), .Z(n46) );
  MUX U70 ( .IN0(n803), .IN1(n379), .SEL(n802), .F(n47) );
  IV U71 ( .A(n47), .Z(n685) );
  MUX U72 ( .IN0(n2345), .IN1(n2353), .SEL(n2346), .F(n48) );
  IV U73 ( .A(n48), .Z(n2348) );
  MUX U74 ( .IN0(n2375), .IN1(n2395), .SEL(n2376), .F(n49) );
  IV U75 ( .A(n49), .Z(n2389) );
  MUX U76 ( .IN0(n50), .IN1(n2304), .SEL(n382), .F(n2300) );
  IV U77 ( .A(o[8]), .Z(n50) );
  MUX U78 ( .IN0(n51), .IN1(n2320), .SEL(n386), .F(n2316) );
  IV U79 ( .A(o[4]), .Z(n51) );
  MUX U80 ( .IN0(n1522), .IN1(n1524), .SEL(n1523), .F(n1430) );
  MUX U81 ( .IN0(n1422), .IN1(n52), .SEL(n1423), .F(n1322) );
  IV U82 ( .A(n1424), .Z(n52) );
  MUX U83 ( .IN0(n1596), .IN1(n53), .SEL(n1597), .F(n1508) );
  IV U84 ( .A(n1598), .Z(n53) );
  MUX U85 ( .IN0(n1406), .IN1(n54), .SEL(n1407), .F(n1310) );
  IV U86 ( .A(n1408), .Z(n54) );
  MUX U87 ( .IN0(n1979), .IN1(n1981), .SEL(n1980), .F(n1913) );
  MUX U88 ( .IN0(n1302), .IN1(n55), .SEL(n1303), .F(n1200) );
  IV U89 ( .A(n1304), .Z(n55) );
  MUX U90 ( .IN0(n1003), .IN1(n56), .SEL(n1004), .F(n890) );
  IV U91 ( .A(n1005), .Z(n56) );
  MUX U92 ( .IN0(n991), .IN1(n57), .SEL(n992), .F(n878) );
  IV U93 ( .A(n993), .Z(n57) );
  MUX U94 ( .IN0(n1488), .IN1(n58), .SEL(n1489), .F(n1392) );
  IV U95 ( .A(n1490), .Z(n58) );
  MUX U96 ( .IN0(n1666), .IN1(n59), .SEL(n1667), .F(n1584) );
  IV U97 ( .A(n1668), .Z(n59) );
  XNOR U98 ( .A(n771), .B(n770), .Z(n767) );
  MUX U99 ( .IN0(n1184), .IN1(n60), .SEL(n1185), .F(n1076) );
  IV U100 ( .A(n1186), .Z(n60) );
  MUX U101 ( .IN0(n975), .IN1(n61), .SEL(n976), .F(n862) );
  IV U102 ( .A(n977), .Z(n61) );
  MUX U103 ( .IN0(n1963), .IN1(n62), .SEL(n1964), .F(n1897) );
  IV U104 ( .A(n1965), .Z(n62) );
  MUX U105 ( .IN0(n2149), .IN1(n63), .SEL(n2150), .F(n2095) );
  IV U106 ( .A(n2151), .Z(n63) );
  XNOR U107 ( .A(n755), .B(n754), .Z(n751) );
  MUX U108 ( .IN0(n959), .IN1(n64), .SEL(n960), .F(n846) );
  IV U109 ( .A(n961), .Z(n64) );
  MUX U110 ( .IN0(n1270), .IN1(n65), .SEL(n1271), .F(n1172) );
  IV U111 ( .A(n1272), .Z(n65) );
  MUX U112 ( .IN0(n1472), .IN1(n66), .SEL(n1473), .F(n1376) );
  IV U113 ( .A(n1474), .Z(n66) );
  MUX U114 ( .IN0(n1650), .IN1(n67), .SEL(n1651), .F(n1568) );
  IV U115 ( .A(n1652), .Z(n67) );
  MUX U116 ( .IN0(n1811), .IN1(n68), .SEL(n1812), .F(n1736) );
  IV U117 ( .A(n1813), .Z(n68) );
  MUX U118 ( .IN0(n1955), .IN1(n69), .SEL(n1956), .F(n1889) );
  IV U119 ( .A(n1957), .Z(n69) );
  MUX U120 ( .IN0(n2141), .IN1(n70), .SEL(n2142), .F(n2087) );
  IV U121 ( .A(n2143), .Z(n70) );
  XNOR U122 ( .A(n739), .B(n738), .Z(n735) );
  MUX U123 ( .IN0(n2242), .IN1(n71), .SEL(n2243), .F(n2195) );
  IV U124 ( .A(n2244), .Z(n71) );
  MUX U125 ( .IN0(n943), .IN1(n72), .SEL(n944), .F(n830) );
  IV U126 ( .A(n945), .Z(n72) );
  MUX U127 ( .IN0(n2133), .IN1(n73), .SEL(n2134), .F(n2079) );
  IV U128 ( .A(n2135), .Z(n73) );
  MUX U129 ( .IN0(n74), .IN1(n2462), .SEL(n2438), .F(n2458) );
  IV U130 ( .A(n2437), .Z(n74) );
  XNOR U131 ( .A(n723), .B(n722), .Z(n719) );
  MUX U132 ( .IN0(n1150), .IN1(n75), .SEL(n1151), .F(n1038) );
  IV U133 ( .A(n1152), .Z(n75) );
  MUX U134 ( .IN0(n1356), .IN1(n76), .SEL(n1357), .F(n1258) );
  IV U135 ( .A(n1358), .Z(n76) );
  MUX U136 ( .IN0(n1548), .IN1(n77), .SEL(n1549), .F(n1460) );
  IV U137 ( .A(n1550), .Z(n77) );
  MUX U138 ( .IN0(n1716), .IN1(n78), .SEL(n1717), .F(n1638) );
  IV U139 ( .A(n1718), .Z(n78) );
  MUX U140 ( .IN0(n1869), .IN1(n79), .SEL(n1870), .F(n1799) );
  IV U141 ( .A(n1871), .Z(n79) );
  MUX U142 ( .IN0(n2005), .IN1(n80), .SEL(n2006), .F(n1943) );
  IV U143 ( .A(n2007), .Z(n80) );
  MUX U144 ( .IN0(n2125), .IN1(n81), .SEL(n2126), .F(n2071) );
  IV U145 ( .A(n2127), .Z(n81) );
  XNOR U146 ( .A(n707), .B(n706), .Z(n703) );
  XNOR U147 ( .A(n816), .B(n815), .Z(n812) );
  MUX U148 ( .IN0(n2384), .IN1(n2386), .SEL(n2385), .F(n2378) );
  MUX U149 ( .IN0(n2348), .IN1(n2350), .SEL(n2349), .F(n2272) );
  MUX U150 ( .IN0(n82), .IN1(n2480), .SEL(n2453), .F(n2476) );
  IV U151 ( .A(n2452), .Z(n82) );
  MUX U152 ( .IN0(n796), .IN1(n907), .SEL(n797), .F(n680) );
  XNOR U153 ( .A(n691), .B(n690), .Z(n687) );
  MUX U154 ( .IN0(n2357), .IN1(n2371), .SEL(n2358), .F(n83) );
  IV U155 ( .A(n83), .Z(n2365) );
  MUX U156 ( .IN0(n2399), .IN1(n2424), .SEL(n2400), .F(n84) );
  IV U157 ( .A(n84), .Z(n2418) );
  MUX U158 ( .IN0(n85), .IN1(n2308), .SEL(n383), .F(n2304) );
  IV U159 ( .A(o[7]), .Z(n85) );
  MUX U160 ( .IN0(n86), .IN1(n2324), .SEL(n387), .F(n2320) );
  IV U161 ( .A(o[3]), .Z(n86) );
  MUX U162 ( .IN0(n1430), .IN1(n1432), .SEL(n1431), .F(n1330) );
  MUX U163 ( .IN0(n87), .IN1(n1772), .SEL(n1773), .F(n1694) );
  IV U164 ( .A(n1774), .Z(n87) );
  MUX U165 ( .IN0(n1322), .IN1(n88), .SEL(n1323), .F(n1220) );
  IV U166 ( .A(n1324), .Z(n88) );
  MUX U167 ( .IN0(n1764), .IN1(n89), .SEL(n1765), .F(n1686) );
  IV U168 ( .A(n1766), .Z(n89) );
  MUX U169 ( .IN0(n1314), .IN1(n90), .SEL(n1315), .F(n1212) );
  IV U170 ( .A(n1316), .Z(n90) );
  MUX U171 ( .IN0(n1120), .IN1(n91), .SEL(n1121), .F(n1003) );
  IV U172 ( .A(n1122), .Z(n91) );
  MUX U173 ( .IN0(n1306), .IN1(n92), .SEL(n1307), .F(n1204) );
  IV U174 ( .A(n1308), .Z(n92) );
  MUX U175 ( .IN0(n1756), .IN1(n93), .SEL(n1757), .F(n1678) );
  IV U176 ( .A(n1758), .Z(n93) );
  MUX U177 ( .IN0(n94), .IN1(n2045), .SEL(n2046), .F(n1983) );
  IV U178 ( .A(n2047), .Z(n94) );
  MUX U179 ( .IN0(n95), .IN1(n894), .SEL(n895), .F(n777) );
  IV U180 ( .A(n896), .Z(n95) );
  XNOR U181 ( .A(n888), .B(n887), .Z(n884) );
  MUX U182 ( .IN0(n1388), .IN1(n96), .SEL(n1389), .F(n1294) );
  IV U183 ( .A(n1390), .Z(n96) );
  MUX U184 ( .IN0(n1580), .IN1(n97), .SEL(n1581), .F(n1492) );
  IV U185 ( .A(n1582), .Z(n97) );
  MUX U186 ( .IN0(n1748), .IN1(n98), .SEL(n1749), .F(n1670) );
  IV U187 ( .A(n1750), .Z(n98) );
  MUX U188 ( .IN0(n1971), .IN1(n99), .SEL(n1972), .F(n1905) );
  IV U189 ( .A(n1973), .Z(n99) );
  MUX U190 ( .IN0(n987), .IN1(n100), .SEL(n988), .F(n874) );
  IV U191 ( .A(n989), .Z(n100) );
  XNOR U192 ( .A(n872), .B(n871), .Z(n868) );
  XNOR U193 ( .A(n763), .B(n762), .Z(n759) );
  MUX U194 ( .IN0(n1180), .IN1(n101), .SEL(n1181), .F(n1072) );
  IV U195 ( .A(n1182), .Z(n101) );
  MUX U196 ( .IN0(n2203), .IN1(n2205), .SEL(n2204), .F(n2153) );
  MUX U197 ( .IN0(n971), .IN1(n102), .SEL(n972), .F(n858) );
  IV U198 ( .A(n973), .Z(n102) );
  XNOR U199 ( .A(n856), .B(n855), .Z(n852) );
  XNOR U200 ( .A(n747), .B(n746), .Z(n743) );
  MUX U201 ( .IN0(n1372), .IN1(n103), .SEL(n1373), .F(n1274) );
  IV U202 ( .A(n1374), .Z(n103) );
  MUX U203 ( .IN0(n1564), .IN1(n104), .SEL(n1565), .F(n1476) );
  IV U204 ( .A(n1566), .Z(n104) );
  MUX U205 ( .IN0(n1732), .IN1(n105), .SEL(n1733), .F(n1654) );
  IV U206 ( .A(n1734), .Z(n105) );
  MUX U207 ( .IN0(n1885), .IN1(n106), .SEL(n1886), .F(n1815) );
  IV U208 ( .A(n1887), .Z(n106) );
  MUX U209 ( .IN0(n2021), .IN1(n107), .SEL(n2022), .F(n1959) );
  IV U210 ( .A(n2023), .Z(n107) );
  MUX U211 ( .IN0(n108), .IN1(n2491), .SEL(n2460), .F(n2296) );
  IV U212 ( .A(n2461), .Z(n108) );
  MUX U213 ( .IN0(n1058), .IN1(n109), .SEL(n1059), .F(n947) );
  IV U214 ( .A(n1060), .Z(n109) );
  MUX U215 ( .IN0(n955), .IN1(n110), .SEL(n956), .F(n842) );
  IV U216 ( .A(n957), .Z(n110) );
  XNOR U217 ( .A(n840), .B(n839), .Z(n836) );
  XNOR U218 ( .A(n731), .B(n730), .Z(n727) );
  MUX U219 ( .IN0(n2187), .IN1(n111), .SEL(n2188), .F(n2137) );
  IV U220 ( .A(n2189), .Z(n111) );
  MUX U221 ( .IN0(n939), .IN1(n112), .SEL(n940), .F(n826) );
  IV U222 ( .A(n941), .Z(n112) );
  MUX U223 ( .IN0(n2402), .IN1(n2404), .SEL(n2403), .F(n2284) );
  XNOR U224 ( .A(n824), .B(n823), .Z(n820) );
  XNOR U225 ( .A(n715), .B(n714), .Z(n711) );
  MUX U226 ( .IN0(n1034), .IN1(n113), .SEL(n1035), .F(n926) );
  IV U227 ( .A(n1036), .Z(n113) );
  MUX U228 ( .IN0(n1254), .IN1(n114), .SEL(n1255), .F(n1154) );
  IV U229 ( .A(n1256), .Z(n114) );
  MUX U230 ( .IN0(n1456), .IN1(n115), .SEL(n1457), .F(n1360) );
  IV U231 ( .A(n1458), .Z(n115) );
  MUX U232 ( .IN0(n1634), .IN1(n116), .SEL(n1635), .F(n1552) );
  IV U233 ( .A(n1636), .Z(n116) );
  MUX U234 ( .IN0(n1795), .IN1(n117), .SEL(n1796), .F(n1720) );
  IV U235 ( .A(n1797), .Z(n117) );
  MUX U236 ( .IN0(n1939), .IN1(n118), .SEL(n1940), .F(n1873) );
  IV U237 ( .A(n1941), .Z(n118) );
  MUX U238 ( .IN0(n2067), .IN1(n119), .SEL(n2068), .F(n2009) );
  IV U239 ( .A(n2069), .Z(n119) );
  MUX U240 ( .IN0(n2225), .IN1(n2267), .SEL(n2227), .F(n2179) );
  MUX U241 ( .IN0(n120), .IN1(n2476), .SEL(n2450), .F(n2470) );
  IV U242 ( .A(n2449), .Z(n120) );
  XNOR U243 ( .A(n699), .B(n698), .Z(n695) );
  MUX U244 ( .IN0(n805), .IN1(n915), .SEL(n806), .F(n689) );
  MUX U245 ( .IN0(n2266), .IN1(n2264), .SEL(n2265), .F(n2221) );
  MUX U246 ( .IN0(n121), .IN1(n2451), .SEL(n2429), .F(n2447) );
  IV U247 ( .A(n2428), .Z(n121) );
  MUX U248 ( .IN0(n794), .IN1(n792), .SEL(n793), .F(n676) );
  MUX U249 ( .IN0(n680), .IN1(n795), .SEL(n681), .F(n437) );
  XNOR U250 ( .A(n2351), .B(n2352), .Z(n2342) );
  XNOR U251 ( .A(n2393), .B(n2394), .Z(n2372) );
  MUX U252 ( .IN0(n122), .IN1(n2312), .SEL(n384), .F(n2308) );
  IV U253 ( .A(o[6]), .Z(n122) );
  MUX U254 ( .IN0(n2328), .IN1(n123), .SEL(n784), .F(n2324) );
  IV U255 ( .A(o[2]), .Z(n123) );
  MUX U256 ( .IN0(n124), .IN1(n1694), .SEL(n1695), .F(n1612) );
  IV U257 ( .A(n1696), .Z(n124) );
  MUX U258 ( .IN0(n1604), .IN1(n125), .SEL(n1605), .F(n1516) );
  IV U259 ( .A(n1606), .Z(n125) );
  MUX U260 ( .IN0(n1330), .IN1(n1332), .SEL(n1331), .F(n1228) );
  MUX U261 ( .IN0(n1843), .IN1(n1845), .SEL(n1844), .F(n1768) );
  MUX U262 ( .IN0(n1318), .IN1(n126), .SEL(n1319), .F(n1216) );
  IV U263 ( .A(n1320), .Z(n126) );
  MUX U264 ( .IN0(n127), .IN1(n1128), .SEL(n1129), .F(n1011) );
  IV U265 ( .A(n1130), .Z(n127) );
  MUX U266 ( .IN0(n1116), .IN1(n128), .SEL(n1117), .F(n999) );
  IV U267 ( .A(n1118), .Z(n128) );
  MUX U268 ( .IN0(n1588), .IN1(n129), .SEL(n1589), .F(n1500) );
  IV U269 ( .A(n1590), .Z(n129) );
  MUX U270 ( .IN0(n1835), .IN1(n130), .SEL(n1836), .F(n1760) );
  IV U271 ( .A(n1837), .Z(n130) );
  MUX U272 ( .IN0(n1108), .IN1(n131), .SEL(n1109), .F(n991) );
  IV U273 ( .A(n1110), .Z(n131) );
  MUX U274 ( .IN0(n1492), .IN1(n132), .SEL(n1493), .F(n1396) );
  IV U275 ( .A(n1494), .Z(n132) );
  MUX U276 ( .IN0(n1294), .IN1(n133), .SEL(n1295), .F(n1192) );
  IV U277 ( .A(n1296), .Z(n133) );
  XNOR U278 ( .A(n775), .B(n774), .Z(n771) );
  XNOR U279 ( .A(n884), .B(n883), .Z(n880) );
  MUX U280 ( .IN0(n1098), .IN1(n134), .SEL(n1099), .F(n983) );
  IV U281 ( .A(n1100), .Z(n134) );
  MUX U282 ( .IN0(n1827), .IN1(n135), .SEL(n1828), .F(n1752) );
  IV U283 ( .A(n1829), .Z(n135) );
  MUX U284 ( .IN0(n2037), .IN1(n136), .SEL(n2038), .F(n1975) );
  IV U285 ( .A(n2039), .Z(n136) );
  MUX U286 ( .IN0(n137), .IN1(n2157), .SEL(n2158), .F(n2103) );
  IV U287 ( .A(n2159), .Z(n137) );
  MUX U288 ( .IN0(n1090), .IN1(n138), .SEL(n1091), .F(n975) );
  IV U289 ( .A(n1092), .Z(n138) );
  XNOR U290 ( .A(n759), .B(n758), .Z(n755) );
  XNOR U291 ( .A(n868), .B(n867), .Z(n864) );
  MUX U292 ( .IN0(n1080), .IN1(n139), .SEL(n1081), .F(n967) );
  IV U293 ( .A(n1082), .Z(n139) );
  MUX U294 ( .IN0(n1480), .IN1(n140), .SEL(n1481), .F(n1384) );
  IV U295 ( .A(n1482), .Z(n140) );
  MUX U296 ( .IN0(n1658), .IN1(n141), .SEL(n1659), .F(n1576) );
  IV U297 ( .A(n1660), .Z(n141) );
  MUX U298 ( .IN0(n1819), .IN1(n142), .SEL(n1820), .F(n1744) );
  IV U299 ( .A(n1821), .Z(n142) );
  MUX U300 ( .IN0(n2029), .IN1(n143), .SEL(n2030), .F(n1967) );
  IV U301 ( .A(n2031), .Z(n143) );
  MUX U302 ( .IN0(n1072), .IN1(n144), .SEL(n1073), .F(n959) );
  IV U303 ( .A(n1074), .Z(n144) );
  XNOR U304 ( .A(n743), .B(n742), .Z(n739) );
  XNOR U305 ( .A(n852), .B(n851), .Z(n848) );
  MUX U306 ( .IN0(n1062), .IN1(n145), .SEL(n1063), .F(n951) );
  IV U307 ( .A(n1064), .Z(n145) );
  MUX U308 ( .IN0(n2195), .IN1(n146), .SEL(n2196), .F(n2145) );
  IV U309 ( .A(n2197), .Z(n146) );
  MUX U310 ( .IN0(n2292), .IN1(n2294), .SEL(n2293), .F(n2250) );
  MUX U311 ( .IN0(n1048), .IN1(n147), .SEL(n1049), .F(n939) );
  IV U312 ( .A(n1050), .Z(n147) );
  XNOR U313 ( .A(n727), .B(n726), .Z(n723) );
  XNOR U314 ( .A(n836), .B(n835), .Z(n832) );
  MUX U315 ( .IN0(n1262), .IN1(n148), .SEL(n1263), .F(n1162) );
  IV U316 ( .A(n1264), .Z(n148) );
  MUX U317 ( .IN0(n1464), .IN1(n149), .SEL(n1465), .F(n1368) );
  IV U318 ( .A(n1466), .Z(n149) );
  MUX U319 ( .IN0(n1642), .IN1(n150), .SEL(n1643), .F(n1560) );
  IV U320 ( .A(n1644), .Z(n150) );
  MUX U321 ( .IN0(n1803), .IN1(n151), .SEL(n1804), .F(n1728) );
  IV U322 ( .A(n1805), .Z(n151) );
  MUX U323 ( .IN0(n1947), .IN1(n152), .SEL(n1948), .F(n1881) );
  IV U324 ( .A(n1949), .Z(n152) );
  MUX U325 ( .IN0(n2075), .IN1(n153), .SEL(n2076), .F(n2017) );
  IV U326 ( .A(n2077), .Z(n153) );
  MUX U327 ( .IN0(n154), .IN1(n2495), .SEL(n2468), .F(n2493) );
  IV U328 ( .A(n2469), .Z(n154) );
  MUX U329 ( .IN0(n2280), .IN1(n155), .SEL(n2281), .F(n2238) );
  IV U330 ( .A(n2282), .Z(n155) );
  MUX U331 ( .IN0(n156), .IN1(n2435), .SEL(n2412), .F(n2431) );
  IV U332 ( .A(n2411), .Z(n156) );
  MUX U333 ( .IN0(n930), .IN1(n157), .SEL(n931), .F(n818) );
  IV U334 ( .A(n932), .Z(n157) );
  XNOR U335 ( .A(n711), .B(n710), .Z(n707) );
  MUX U336 ( .IN0(n2230), .IN1(n158), .SEL(n2231), .F(n2183) );
  IV U337 ( .A(n2232), .Z(n158) );
  MUX U338 ( .IN0(n159), .IN1(n814), .SEL(n815), .F(n697) );
  IV U339 ( .A(n816), .Z(n159) );
  MUX U340 ( .IN0(n1029), .IN1(n1141), .SEL(n1031), .F(n922) );
  XNOR U341 ( .A(n695), .B(n694), .Z(n691) );
  MUX U342 ( .IN0(n1246), .IN1(n1248), .SEL(n1247), .F(n160) );
  IV U343 ( .A(n160), .Z(n1146) );
  MUX U344 ( .IN0(n1448), .IN1(n1450), .SEL(n1449), .F(n161) );
  IV U345 ( .A(n161), .Z(n1352) );
  MUX U346 ( .IN0(n1626), .IN1(n1628), .SEL(n1627), .F(n162) );
  IV U347 ( .A(n162), .Z(n1544) );
  MUX U348 ( .IN0(n1787), .IN1(n1789), .SEL(n1788), .F(n163) );
  IV U349 ( .A(n163), .Z(n1712) );
  MUX U350 ( .IN0(n1931), .IN1(n1933), .SEL(n1932), .F(n164) );
  IV U351 ( .A(n164), .Z(n1865) );
  MUX U352 ( .IN0(n2059), .IN1(n2061), .SEL(n2060), .F(n165) );
  IV U353 ( .A(n165), .Z(n2001) );
  MUX U354 ( .IN0(n2171), .IN1(n2173), .SEL(n2172), .F(n166) );
  IV U355 ( .A(n166), .Z(n2121) );
  MUX U356 ( .IN0(n2486), .IN1(n2503), .SEL(n2485), .F(n167) );
  IV U357 ( .A(n167), .Z(n2501) );
  XNOR U358 ( .A(n808), .B(n807), .Z(n803) );
  MUX U359 ( .IN0(n1023), .IN1(n1021), .SEL(n1022), .F(n912) );
  MUX U360 ( .IN0(n2338), .IN1(n2341), .SEL(n2339), .F(n2268) );
  XNOR U361 ( .A(n2369), .B(n2370), .Z(n2354) );
  XNOR U362 ( .A(n2422), .B(n2423), .Z(n2396) );
  MUX U363 ( .IN0(n676), .IN1(n678), .SEL(n677), .F(n168) );
  IV U364 ( .A(n168), .Z(n421) );
  MUX U365 ( .IN0(o[29]), .IN1(n666), .SEL(n667), .F(n424) );
  MUX U366 ( .IN0(o[25]), .IN1(n1132), .SEL(n1133), .F(n1015) );
  MUX U367 ( .IN0(o[21]), .IN1(n1530), .SEL(n1531), .F(n1438) );
  MUX U368 ( .IN0(o[17]), .IN1(n1851), .SEL(n1852), .F(n1777) );
  MUX U369 ( .IN0(o[13]), .IN1(n2107), .SEL(n2108), .F(n2049) );
  MUX U370 ( .IN0(o[9]), .IN1(n169), .SEL(n381), .F(n2258) );
  IV U371 ( .A(n2300), .Z(n169) );
  MUX U372 ( .IN0(n170), .IN1(n2316), .SEL(n385), .F(n2312) );
  IV U373 ( .A(o[5]), .Z(n170) );
  MUX U374 ( .IN0(n171), .IN1(n2332), .SEL(n1775), .F(n2328) );
  IV U375 ( .A(o[1]), .Z(n171) );
  MUX U376 ( .IN0(n172), .IN1(n1612), .SEL(n1613), .F(n1526) );
  IV U377 ( .A(n1614), .Z(n172) );
  MUX U378 ( .IN0(n1690), .IN1(n1692), .SEL(n1691), .F(n1608) );
  MUX U379 ( .IN0(n1508), .IN1(n173), .SEL(n1509), .F(n1416) );
  IV U380 ( .A(n1510), .Z(n173) );
  MUX U381 ( .IN0(n174), .IN1(n1232), .SEL(n1233), .F(n1128) );
  IV U382 ( .A(n1234), .Z(n174) );
  MUX U383 ( .IN0(n1682), .IN1(n175), .SEL(n1683), .F(n1600) );
  IV U384 ( .A(n1684), .Z(n175) );
  MUX U385 ( .IN0(n176), .IN1(n1917), .SEL(n1918), .F(n1847) );
  IV U386 ( .A(n1919), .Z(n176) );
  MUX U387 ( .IN0(n1224), .IN1(n177), .SEL(n1225), .F(n1120) );
  IV U388 ( .A(n1226), .Z(n177) );
  MUX U389 ( .IN0(n1310), .IN1(n178), .SEL(n1311), .F(n1208) );
  IV U390 ( .A(n1312), .Z(n178) );
  MUX U391 ( .IN0(n1007), .IN1(n1009), .SEL(n1008), .F(n894) );
  MUX U392 ( .IN0(n1496), .IN1(n179), .SEL(n1497), .F(n1402) );
  IV U393 ( .A(n1498), .Z(n179) );
  MUX U394 ( .IN0(n1674), .IN1(n180), .SEL(n1675), .F(n1592) );
  IV U395 ( .A(n1676), .Z(n180) );
  MUX U396 ( .IN0(n1909), .IN1(n181), .SEL(n1910), .F(n1839) );
  IV U397 ( .A(n1911), .Z(n181) );
  MUX U398 ( .IN0(n1112), .IN1(n182), .SEL(n1113), .F(n995) );
  IV U399 ( .A(n1114), .Z(n182) );
  MUX U400 ( .IN0(n999), .IN1(n183), .SEL(n1000), .F(n886) );
  IV U401 ( .A(n1001), .Z(n183) );
  MUX U402 ( .IN0(n1392), .IN1(n184), .SEL(n1393), .F(n1298) );
  IV U403 ( .A(n1394), .Z(n184) );
  MUX U404 ( .IN0(n783), .IN1(n185), .SEL(n782), .F(n514) );
  IV U405 ( .A(n781), .Z(n185) );
  MUX U406 ( .IN0(n1901), .IN1(n186), .SEL(n1902), .F(n1831) );
  IV U407 ( .A(n1903), .Z(n186) );
  MUX U408 ( .IN0(n2099), .IN1(n2101), .SEL(n2100), .F(n2041) );
  MUX U409 ( .IN0(n1094), .IN1(n187), .SEL(n1095), .F(n979) );
  IV U410 ( .A(n1096), .Z(n187) );
  XNOR U411 ( .A(n880), .B(n879), .Z(n876) );
  XNOR U412 ( .A(n767), .B(n766), .Z(n763) );
  MUX U413 ( .IN0(n983), .IN1(n188), .SEL(n984), .F(n870) );
  IV U414 ( .A(n985), .Z(n188) );
  MUX U415 ( .IN0(n1572), .IN1(n189), .SEL(n1573), .F(n1484) );
  IV U416 ( .A(n1574), .Z(n189) );
  MUX U417 ( .IN0(n1740), .IN1(n190), .SEL(n1741), .F(n1662) );
  IV U418 ( .A(n1742), .Z(n190) );
  MUX U419 ( .IN0(n1893), .IN1(n191), .SEL(n1894), .F(n1823) );
  IV U420 ( .A(n1895), .Z(n191) );
  MUX U421 ( .IN0(n2091), .IN1(n192), .SEL(n2092), .F(n2033) );
  IV U422 ( .A(n2093), .Z(n192) );
  MUX U423 ( .IN0(n193), .IN1(n2254), .SEL(n2255), .F(n2207) );
  IV U424 ( .A(n2256), .Z(n193) );
  MUX U425 ( .IN0(n1176), .IN1(n194), .SEL(n1177), .F(n1066) );
  IV U426 ( .A(n1178), .Z(n194) );
  MUX U427 ( .IN0(n1076), .IN1(n195), .SEL(n1077), .F(n963) );
  IV U428 ( .A(n1078), .Z(n195) );
  XNOR U429 ( .A(n864), .B(n863), .Z(n860) );
  XNOR U430 ( .A(n751), .B(n750), .Z(n747) );
  MUX U431 ( .IN0(n967), .IN1(n196), .SEL(n968), .F(n854) );
  IV U432 ( .A(n969), .Z(n196) );
  MUX U433 ( .IN0(n2083), .IN1(n197), .SEL(n2084), .F(n2025) );
  IV U434 ( .A(n2085), .Z(n197) );
  MUX U435 ( .IN0(n2246), .IN1(n198), .SEL(n2247), .F(n2199) );
  IV U436 ( .A(n2248), .Z(n198) );
  XNOR U437 ( .A(n848), .B(n847), .Z(n844) );
  XNOR U438 ( .A(n735), .B(n734), .Z(n731) );
  MUX U439 ( .IN0(n951), .IN1(n199), .SEL(n952), .F(n838) );
  IV U440 ( .A(n953), .Z(n199) );
  MUX U441 ( .IN0(n1158), .IN1(n200), .SEL(n1159), .F(n1048) );
  IV U442 ( .A(n1160), .Z(n200) );
  MUX U443 ( .IN0(n1364), .IN1(n201), .SEL(n1365), .F(n1266) );
  IV U444 ( .A(n1366), .Z(n201) );
  MUX U445 ( .IN0(n1556), .IN1(n202), .SEL(n1557), .F(n1468) );
  IV U446 ( .A(n1558), .Z(n202) );
  MUX U447 ( .IN0(n1724), .IN1(n203), .SEL(n1725), .F(n1646) );
  IV U448 ( .A(n1726), .Z(n203) );
  MUX U449 ( .IN0(n1877), .IN1(n204), .SEL(n1878), .F(n1807) );
  IV U450 ( .A(n1879), .Z(n204) );
  MUX U451 ( .IN0(n2013), .IN1(n205), .SEL(n2014), .F(n1951) );
  IV U452 ( .A(n2015), .Z(n205) );
  MUX U453 ( .IN0(n2238), .IN1(n206), .SEL(n2239), .F(n2191) );
  IV U454 ( .A(n2240), .Z(n206) );
  XNOR U455 ( .A(n832), .B(n831), .Z(n828) );
  XNOR U456 ( .A(n719), .B(n718), .Z(n715) );
  MUX U457 ( .IN0(n934), .IN1(n207), .SEL(n935), .F(n822) );
  IV U458 ( .A(n936), .Z(n207) );
  MUX U459 ( .IN0(n208), .IN1(n2497), .SEL(n2474), .F(n2495) );
  IV U460 ( .A(n2475), .Z(n208) );
  MUX U461 ( .IN0(n926), .IN1(n209), .SEL(n927), .F(n814) );
  IV U462 ( .A(n928), .Z(n209) );
  MUX U463 ( .IN0(n2179), .IN1(n210), .SEL(n2180), .F(n2129) );
  IV U464 ( .A(n2181), .Z(n210) );
  MUX U465 ( .IN0(n2276), .IN1(n211), .SEL(n2277), .F(n2234) );
  IV U466 ( .A(n2278), .Z(n211) );
  XNOR U467 ( .A(n703), .B(n702), .Z(n699) );
  XNOR U468 ( .A(n2405), .B(n2406), .Z(n2382) );
  XNOR U469 ( .A(n812), .B(n811), .Z(n808) );
  MUX U470 ( .IN0(n1142), .IN1(n1144), .SEL(n1143), .F(n212) );
  IV U471 ( .A(n212), .Z(n1029) );
  MUX U472 ( .IN0(n1348), .IN1(n1350), .SEL(n1349), .F(n213) );
  IV U473 ( .A(n213), .Z(n1250) );
  MUX U474 ( .IN0(n1540), .IN1(n1542), .SEL(n1541), .F(n214) );
  IV U475 ( .A(n214), .Z(n1452) );
  MUX U476 ( .IN0(n1708), .IN1(n1710), .SEL(n1709), .F(n215) );
  IV U477 ( .A(n215), .Z(n1630) );
  MUX U478 ( .IN0(n1861), .IN1(n1863), .SEL(n1862), .F(n216) );
  IV U479 ( .A(n216), .Z(n1791) );
  MUX U480 ( .IN0(n1997), .IN1(n1999), .SEL(n1998), .F(n217) );
  IV U481 ( .A(n217), .Z(n1935) );
  MUX U482 ( .IN0(n2117), .IN1(n2119), .SEL(n2118), .F(n218) );
  IV U483 ( .A(n218), .Z(n2063) );
  MUX U484 ( .IN0(n2221), .IN1(n2223), .SEL(n2222), .F(n219) );
  IV U485 ( .A(n219), .Z(n2175) );
  XNOR U486 ( .A(n2411), .B(n2412), .Z(n2387) );
  MUX U487 ( .IN0(n220), .IN1(n908), .SEL(n909), .F(n796) );
  IV U488 ( .A(n910), .Z(n220) );
  XNOR U489 ( .A(n2416), .B(n2417), .Z(n2393) );
  MUX U490 ( .IN0(n221), .IN1(n2484), .SEL(n2456), .F(n2480) );
  IV U491 ( .A(n2455), .Z(n221) );
  MUX U492 ( .IN0(n222), .IN1(n685), .SEL(n686), .F(n443) );
  IV U493 ( .A(n687), .Z(n222) );
  MUX U494 ( .IN0(n223), .IN1(n672), .SEL(n673), .F(n415) );
  IV U495 ( .A(n674), .Z(n223) );
  XNOR U496 ( .A(n2342), .B(n2343), .Z(n2338) );
  XNOR U497 ( .A(n2396), .B(n2397), .Z(n2375) );
  MUX U498 ( .IN0(o[26]), .IN1(n1015), .SEL(n1016), .F(n902) );
  MUX U499 ( .IN0(o[22]), .IN1(n1438), .SEL(n1439), .F(n1338) );
  MUX U500 ( .IN0(o[18]), .IN1(n1777), .SEL(n1778), .F(n1698) );
  MUX U501 ( .IN0(o[14]), .IN1(n2049), .SEL(n2050), .F(n1987) );
  MUX U502 ( .IN0(o[10]), .IN1(n2258), .SEL(n2259), .F(n2211) );
  XNOR U503 ( .A(n2345), .B(n2346), .Z(n2306) );
  XNOR U504 ( .A(n2399), .B(n2400), .Z(n2318) );
  XNOR U505 ( .A(n2308), .B(n2311), .Z(n2309) );
  XNOR U506 ( .A(n2320), .B(n2323), .Z(n2321) );
  MUX U507 ( .IN0(n1608), .IN1(n1610), .SEL(n1609), .F(n1522) );
  MUX U508 ( .IN0(n224), .IN1(n1334), .SEL(n1335), .F(n1232) );
  IV U509 ( .A(n1336), .Z(n224) );
  MUX U510 ( .IN0(n1686), .IN1(n225), .SEL(n1687), .F(n1604) );
  IV U511 ( .A(n1688), .Z(n225) );
  MUX U512 ( .IN0(n226), .IN1(n1847), .SEL(n1848), .F(n1772) );
  IV U513 ( .A(n1849), .Z(n226) );
  MUX U514 ( .IN0(n1326), .IN1(n227), .SEL(n1327), .F(n1224) );
  IV U515 ( .A(n1328), .Z(n227) );
  MUX U516 ( .IN0(n1124), .IN1(n1126), .SEL(n1125), .F(n1007) );
  MUX U517 ( .IN0(n1402), .IN1(n228), .SEL(n1403), .F(n1306) );
  IV U518 ( .A(n1404), .Z(n228) );
  MUX U519 ( .IN0(n1592), .IN1(n229), .SEL(n1593), .F(n1504) );
  IV U520 ( .A(n1594), .Z(n229) );
  MUX U521 ( .IN0(n1760), .IN1(n230), .SEL(n1761), .F(n1682) );
  IV U522 ( .A(n1762), .Z(n230) );
  MUX U523 ( .IN0(n1913), .IN1(n1915), .SEL(n1914), .F(n1843) );
  MUX U524 ( .IN0(n1216), .IN1(n231), .SEL(n1217), .F(n1112) );
  IV U525 ( .A(n1218), .Z(n231) );
  MUX U526 ( .IN0(n1208), .IN1(n232), .SEL(n1209), .F(n1102) );
  IV U527 ( .A(n1210), .Z(n232) );
  MUX U528 ( .IN0(n233), .IN1(n898), .SEL(n899), .F(n781) );
  IV U529 ( .A(n900), .Z(n233) );
  MUX U530 ( .IN0(n1670), .IN1(n234), .SEL(n1671), .F(n1588) );
  IV U531 ( .A(n1672), .Z(n234) );
  MUX U532 ( .IN0(n1831), .IN1(n235), .SEL(n1832), .F(n1756) );
  IV U533 ( .A(n1833), .Z(n235) );
  MUX U534 ( .IN0(n1975), .IN1(n236), .SEL(n1976), .F(n1909) );
  IV U535 ( .A(n1977), .Z(n236) );
  MUX U536 ( .IN0(n237), .IN1(n2103), .SEL(n2104), .F(n2045) );
  IV U537 ( .A(n2105), .Z(n237) );
  MUX U538 ( .IN0(n1200), .IN1(n238), .SEL(n1201), .F(n1094) );
  IV U539 ( .A(n1202), .Z(n238) );
  MUX U540 ( .IN0(n239), .IN1(n886), .SEL(n887), .F(n769) );
  IV U541 ( .A(n888), .Z(n239) );
  MUX U542 ( .IN0(n1192), .IN1(n240), .SEL(n1193), .F(n1084) );
  IV U543 ( .A(n1194), .Z(n240) );
  MUX U544 ( .IN0(n241), .IN1(n773), .SEL(n774), .F(n517) );
  IV U545 ( .A(n775), .Z(n241) );
  MUX U546 ( .IN0(n242), .IN1(n878), .SEL(n879), .F(n761) );
  IV U547 ( .A(n880), .Z(n242) );
  MUX U548 ( .IN0(n1384), .IN1(n243), .SEL(n1385), .F(n1288) );
  IV U549 ( .A(n1386), .Z(n243) );
  MUX U550 ( .IN0(n1576), .IN1(n244), .SEL(n1577), .F(n1488) );
  IV U551 ( .A(n1578), .Z(n244) );
  MUX U552 ( .IN0(n1744), .IN1(n245), .SEL(n1745), .F(n1666) );
  IV U553 ( .A(n1746), .Z(n245) );
  MUX U554 ( .IN0(n1897), .IN1(n246), .SEL(n1898), .F(n1827) );
  IV U555 ( .A(n1899), .Z(n246) );
  MUX U556 ( .IN0(n2033), .IN1(n247), .SEL(n2034), .F(n1971) );
  IV U557 ( .A(n2035), .Z(n247) );
  MUX U558 ( .IN0(n2153), .IN1(n2155), .SEL(n2154), .F(n2099) );
  MUX U559 ( .IN0(n248), .IN1(n765), .SEL(n766), .F(n509) );
  IV U560 ( .A(n767), .Z(n248) );
  MUX U561 ( .IN0(n249), .IN1(n870), .SEL(n871), .F(n753) );
  IV U562 ( .A(n872), .Z(n249) );
  MUX U563 ( .IN0(n250), .IN1(n757), .SEL(n758), .F(n503) );
  IV U564 ( .A(n759), .Z(n250) );
  MUX U565 ( .IN0(n251), .IN1(n862), .SEL(n863), .F(n745) );
  IV U566 ( .A(n864), .Z(n251) );
  MUX U567 ( .IN0(n1274), .IN1(n252), .SEL(n1275), .F(n1176) );
  IV U568 ( .A(n1276), .Z(n252) );
  MUX U569 ( .IN0(n1476), .IN1(n253), .SEL(n1477), .F(n1380) );
  IV U570 ( .A(n1478), .Z(n253) );
  MUX U571 ( .IN0(n1654), .IN1(n254), .SEL(n1655), .F(n1572) );
  IV U572 ( .A(n1656), .Z(n254) );
  MUX U573 ( .IN0(n1815), .IN1(n255), .SEL(n1816), .F(n1740) );
  IV U574 ( .A(n1817), .Z(n255) );
  MUX U575 ( .IN0(n1959), .IN1(n256), .SEL(n1960), .F(n1893) );
  IV U576 ( .A(n1961), .Z(n256) );
  MUX U577 ( .IN0(n2087), .IN1(n257), .SEL(n2088), .F(n2029) );
  IV U578 ( .A(n2089), .Z(n257) );
  MUX U579 ( .IN0(n2199), .IN1(n258), .SEL(n2200), .F(n2149) );
  IV U580 ( .A(n2201), .Z(n258) );
  MUX U581 ( .IN0(n259), .IN1(n2296), .SEL(n2297), .F(n2254) );
  IV U582 ( .A(n2298), .Z(n259) );
  MUX U583 ( .IN0(n260), .IN1(n749), .SEL(n750), .F(n497) );
  IV U584 ( .A(n751), .Z(n260) );
  MUX U585 ( .IN0(n261), .IN1(n854), .SEL(n855), .F(n737) );
  IV U586 ( .A(n856), .Z(n261) );
  MUX U587 ( .IN0(n262), .IN1(n741), .SEL(n742), .F(n491) );
  IV U588 ( .A(n743), .Z(n262) );
  MUX U589 ( .IN0(n263), .IN1(n846), .SEL(n847), .F(n729) );
  IV U590 ( .A(n848), .Z(n263) );
  MUX U591 ( .IN0(n1368), .IN1(n264), .SEL(n1369), .F(n1270) );
  IV U592 ( .A(n1370), .Z(n264) );
  MUX U593 ( .IN0(n1560), .IN1(n265), .SEL(n1561), .F(n1472) );
  IV U594 ( .A(n1562), .Z(n265) );
  MUX U595 ( .IN0(n1728), .IN1(n266), .SEL(n1729), .F(n1650) );
  IV U596 ( .A(n1730), .Z(n266) );
  MUX U597 ( .IN0(n1881), .IN1(n267), .SEL(n1882), .F(n1811) );
  IV U598 ( .A(n1883), .Z(n267) );
  MUX U599 ( .IN0(n2017), .IN1(n268), .SEL(n2018), .F(n1955) );
  IV U600 ( .A(n2019), .Z(n268) );
  MUX U601 ( .IN0(n2137), .IN1(n269), .SEL(n2138), .F(n2083) );
  IV U602 ( .A(n2139), .Z(n269) );
  MUX U603 ( .IN0(n270), .IN1(n2458), .SEL(n2434), .F(n2292) );
  IV U604 ( .A(n2433), .Z(n270) );
  MUX U605 ( .IN0(n271), .IN1(n733), .SEL(n734), .F(n485) );
  IV U606 ( .A(n735), .Z(n271) );
  MUX U607 ( .IN0(n272), .IN1(n838), .SEL(n839), .F(n721) );
  IV U608 ( .A(n840), .Z(n272) );
  MUX U609 ( .IN0(n2284), .IN1(n273), .SEL(n2285), .F(n2242) );
  IV U610 ( .A(n2286), .Z(n273) );
  MUX U611 ( .IN0(n274), .IN1(n725), .SEL(n726), .F(n479) );
  IV U612 ( .A(n727), .Z(n274) );
  MUX U613 ( .IN0(n275), .IN1(n830), .SEL(n831), .F(n713) );
  IV U614 ( .A(n832), .Z(n275) );
  MUX U615 ( .IN0(n1258), .IN1(n276), .SEL(n1259), .F(n1158) );
  IV U616 ( .A(n1260), .Z(n276) );
  MUX U617 ( .IN0(n1460), .IN1(n277), .SEL(n1461), .F(n1364) );
  IV U618 ( .A(n1462), .Z(n277) );
  MUX U619 ( .IN0(n1638), .IN1(n278), .SEL(n1639), .F(n1556) );
  IV U620 ( .A(n1640), .Z(n278) );
  MUX U621 ( .IN0(n1799), .IN1(n279), .SEL(n1800), .F(n1724) );
  IV U622 ( .A(n1801), .Z(n279) );
  MUX U623 ( .IN0(n1943), .IN1(n280), .SEL(n1944), .F(n1877) );
  IV U624 ( .A(n1945), .Z(n280) );
  MUX U625 ( .IN0(n2071), .IN1(n281), .SEL(n2072), .F(n2013) );
  IV U626 ( .A(n2073), .Z(n281) );
  MUX U627 ( .IN0(n2183), .IN1(n282), .SEL(n2184), .F(n2133) );
  IV U628 ( .A(n2185), .Z(n282) );
  MUX U629 ( .IN0(n283), .IN1(n717), .SEL(n718), .F(n473) );
  IV U630 ( .A(n719), .Z(n283) );
  MUX U631 ( .IN0(n284), .IN1(n822), .SEL(n823), .F(n705) );
  IV U632 ( .A(n824), .Z(n284) );
  MUX U633 ( .IN0(n285), .IN1(n2439), .SEL(n2417), .F(n2435) );
  IV U634 ( .A(n2416), .Z(n285) );
  MUX U635 ( .IN0(n286), .IN1(n2499), .SEL(n2478), .F(n2497) );
  IV U636 ( .A(n2479), .Z(n286) );
  MUX U637 ( .IN0(n287), .IN1(n709), .SEL(n710), .F(n467) );
  IV U638 ( .A(n711), .Z(n287) );
  MUX U639 ( .IN0(n1146), .IN1(n288), .SEL(n1147), .F(n1034) );
  IV U640 ( .A(n1148), .Z(n288) );
  MUX U641 ( .IN0(n1352), .IN1(n289), .SEL(n1353), .F(n1254) );
  IV U642 ( .A(n1354), .Z(n289) );
  MUX U643 ( .IN0(n1544), .IN1(n290), .SEL(n1545), .F(n1456) );
  IV U644 ( .A(n1546), .Z(n290) );
  MUX U645 ( .IN0(n1712), .IN1(n291), .SEL(n1713), .F(n1634) );
  IV U646 ( .A(n1714), .Z(n291) );
  MUX U647 ( .IN0(n1865), .IN1(n292), .SEL(n1866), .F(n1795) );
  IV U648 ( .A(n1867), .Z(n292) );
  MUX U649 ( .IN0(n2001), .IN1(n293), .SEL(n2002), .F(n1939) );
  IV U650 ( .A(n2003), .Z(n293) );
  MUX U651 ( .IN0(n2121), .IN1(n294), .SEL(n2122), .F(n2067) );
  IV U652 ( .A(n2123), .Z(n294) );
  MUX U653 ( .IN0(n295), .IN1(n701), .SEL(n702), .F(n461) );
  IV U654 ( .A(n703), .Z(n295) );
  MUX U655 ( .IN0(n1025), .IN1(n1027), .SEL(n1026), .F(n296) );
  IV U656 ( .A(n296), .Z(n916) );
  MUX U657 ( .IN0(n2268), .IN1(n2270), .SEL(n2269), .F(n297) );
  IV U658 ( .A(n297), .Z(n2225) );
  MUX U659 ( .IN0(n298), .IN1(n693), .SEL(n694), .F(n455) );
  IV U660 ( .A(n695), .Z(n298) );
  XNOR U661 ( .A(n687), .B(n686), .Z(n683) );
  MUX U662 ( .IN0(n1244), .IN1(n1242), .SEL(n1243), .F(n1142) );
  MUX U663 ( .IN0(n1446), .IN1(n1444), .SEL(n1445), .F(n1348) );
  MUX U664 ( .IN0(n1624), .IN1(n1622), .SEL(n1623), .F(n1540) );
  MUX U665 ( .IN0(n1785), .IN1(n1783), .SEL(n1784), .F(n1708) );
  MUX U666 ( .IN0(n1929), .IN1(n1927), .SEL(n1928), .F(n1861) );
  MUX U667 ( .IN0(n2057), .IN1(n2055), .SEL(n2056), .F(n1997) );
  MUX U668 ( .IN0(n2169), .IN1(n2167), .SEL(n2168), .F(n2117) );
  XNOR U669 ( .A(n2363), .B(n2364), .Z(n2351) );
  XNOR U670 ( .A(n803), .B(n802), .Z(n799) );
  XNOR U671 ( .A(n2354), .B(n2355), .Z(n2345) );
  XNOR U672 ( .A(n2425), .B(n2426), .Z(n2399) );
  AND U673 ( .A(g_input[1]), .B(n2506), .Z(n2507) );
  XNOR U674 ( .A(n414), .B(n413), .Z(n396) );
  MUX U675 ( .IN0(o[28]), .IN1(n786), .SEL(n787), .F(n666) );
  MUX U676 ( .IN0(o[24]), .IN1(n1236), .SEL(n1237), .F(n1132) );
  MUX U677 ( .IN0(o[20]), .IN1(n1616), .SEL(n1617), .F(n1530) );
  MUX U678 ( .IN0(o[16]), .IN1(n1921), .SEL(n1922), .F(n1851) );
  MUX U679 ( .IN0(o[12]), .IN1(n2161), .SEL(n2162), .F(n2107) );
  XNOR U680 ( .A(n2357), .B(n2358), .Z(n2310) );
  XNOR U681 ( .A(n2428), .B(n2429), .Z(n2322) );
  XNOR U682 ( .A(n2300), .B(n2303), .Z(n2301) );
  XNOR U683 ( .A(n2312), .B(n2315), .Z(n2313) );
  XNOR U684 ( .A(n2324), .B(n2327), .Z(n2325) );
  MUX U685 ( .IN0(n299), .IN1(n1434), .SEL(n1435), .F(n1334) );
  IV U686 ( .A(n1436), .Z(n299) );
  MUX U687 ( .IN0(n1426), .IN1(n300), .SEL(n1427), .F(n1326) );
  IV U688 ( .A(n1428), .Z(n300) );
  MUX U689 ( .IN0(n1600), .IN1(n301), .SEL(n1601), .F(n1512) );
  IV U690 ( .A(n1602), .Z(n301) );
  MUX U691 ( .IN0(n1768), .IN1(n1770), .SEL(n1769), .F(n1690) );
  MUX U692 ( .IN0(n1228), .IN1(n1230), .SEL(n1229), .F(n1124) );
  MUX U693 ( .IN0(n1220), .IN1(n302), .SEL(n1221), .F(n1116) );
  IV U694 ( .A(n1222), .Z(n302) );
  MUX U695 ( .IN0(n1500), .IN1(n303), .SEL(n1501), .F(n1406) );
  IV U696 ( .A(n1502), .Z(n303) );
  MUX U697 ( .IN0(n1678), .IN1(n304), .SEL(n1679), .F(n1596) );
  IV U698 ( .A(n1680), .Z(n304) );
  MUX U699 ( .IN0(n1839), .IN1(n305), .SEL(n1840), .F(n1764) );
  IV U700 ( .A(n1841), .Z(n305) );
  MUX U701 ( .IN0(n306), .IN1(n1983), .SEL(n1984), .F(n1917) );
  IV U702 ( .A(n1985), .Z(n306) );
  MUX U703 ( .IN0(n307), .IN1(n1011), .SEL(n1012), .F(n898) );
  IV U704 ( .A(n1013), .Z(n307) );
  MUX U705 ( .IN0(n1212), .IN1(n308), .SEL(n1213), .F(n1108) );
  IV U706 ( .A(n1214), .Z(n308) );
  MUX U707 ( .IN0(n1204), .IN1(n309), .SEL(n1205), .F(n1098) );
  IV U708 ( .A(n1206), .Z(n309) );
  MUX U709 ( .IN0(n1584), .IN1(n310), .SEL(n1585), .F(n1496) );
  IV U710 ( .A(n1586), .Z(n310) );
  MUX U711 ( .IN0(n1752), .IN1(n311), .SEL(n1753), .F(n1674) );
  IV U712 ( .A(n1754), .Z(n311) );
  MUX U713 ( .IN0(n1905), .IN1(n312), .SEL(n1906), .F(n1835) );
  IV U714 ( .A(n1907), .Z(n312) );
  MUX U715 ( .IN0(n2041), .IN1(n2043), .SEL(n2042), .F(n1979) );
  MUX U716 ( .IN0(n313), .IN1(n890), .SEL(n891), .F(n773) );
  IV U717 ( .A(n892), .Z(n313) );
  MUX U718 ( .IN0(n314), .IN1(n777), .SEL(n778), .F(n519) );
  IV U719 ( .A(n779), .Z(n314) );
  MUX U720 ( .IN0(n1196), .IN1(n315), .SEL(n1197), .F(n1090) );
  IV U721 ( .A(n1198), .Z(n315) );
  MUX U722 ( .IN0(n316), .IN1(n882), .SEL(n883), .F(n765) );
  IV U723 ( .A(n884), .Z(n316) );
  MUX U724 ( .IN0(n317), .IN1(n769), .SEL(n770), .F(n516) );
  IV U725 ( .A(n771), .Z(n317) );
  MUX U726 ( .IN0(n1188), .IN1(n318), .SEL(n1189), .F(n1080) );
  IV U727 ( .A(n1190), .Z(n318) );
  MUX U728 ( .IN0(n1284), .IN1(n319), .SEL(n1285), .F(n1184) );
  IV U729 ( .A(n1286), .Z(n319) );
  MUX U730 ( .IN0(n1484), .IN1(n320), .SEL(n1485), .F(n1388) );
  IV U731 ( .A(n1486), .Z(n320) );
  MUX U732 ( .IN0(n1662), .IN1(n321), .SEL(n1663), .F(n1580) );
  IV U733 ( .A(n1664), .Z(n321) );
  MUX U734 ( .IN0(n1823), .IN1(n322), .SEL(n1824), .F(n1748) );
  IV U735 ( .A(n1825), .Z(n322) );
  MUX U736 ( .IN0(n1967), .IN1(n323), .SEL(n1968), .F(n1901) );
  IV U737 ( .A(n1969), .Z(n323) );
  MUX U738 ( .IN0(n2095), .IN1(n324), .SEL(n2096), .F(n2037) );
  IV U739 ( .A(n2097), .Z(n324) );
  MUX U740 ( .IN0(n325), .IN1(n2207), .SEL(n2208), .F(n2157) );
  IV U741 ( .A(n2209), .Z(n325) );
  MUX U742 ( .IN0(n326), .IN1(n874), .SEL(n875), .F(n757) );
  IV U743 ( .A(n876), .Z(n326) );
  MUX U744 ( .IN0(n327), .IN1(n761), .SEL(n762), .F(n508) );
  IV U745 ( .A(n763), .Z(n327) );
  MUX U746 ( .IN0(n328), .IN1(n866), .SEL(n867), .F(n749) );
  IV U747 ( .A(n868), .Z(n328) );
  MUX U748 ( .IN0(n329), .IN1(n753), .SEL(n754), .F(n502) );
  IV U749 ( .A(n755), .Z(n329) );
  MUX U750 ( .IN0(n1172), .IN1(n330), .SEL(n1173), .F(n1062) );
  IV U751 ( .A(n1174), .Z(n330) );
  MUX U752 ( .IN0(n1376), .IN1(n331), .SEL(n1377), .F(n1278) );
  IV U753 ( .A(n1378), .Z(n331) );
  MUX U754 ( .IN0(n1568), .IN1(n332), .SEL(n1569), .F(n1480) );
  IV U755 ( .A(n1570), .Z(n332) );
  MUX U756 ( .IN0(n1736), .IN1(n333), .SEL(n1737), .F(n1658) );
  IV U757 ( .A(n1738), .Z(n333) );
  MUX U758 ( .IN0(n1889), .IN1(n334), .SEL(n1890), .F(n1819) );
  IV U759 ( .A(n1891), .Z(n334) );
  MUX U760 ( .IN0(n2025), .IN1(n335), .SEL(n2026), .F(n1963) );
  IV U761 ( .A(n2027), .Z(n335) );
  MUX U762 ( .IN0(n2145), .IN1(n336), .SEL(n2146), .F(n2091) );
  IV U763 ( .A(n2147), .Z(n336) );
  MUX U764 ( .IN0(n2250), .IN1(n2252), .SEL(n2251), .F(n2203) );
  MUX U765 ( .IN0(n337), .IN1(n858), .SEL(n859), .F(n741) );
  IV U766 ( .A(n860), .Z(n337) );
  MUX U767 ( .IN0(n338), .IN1(n745), .SEL(n746), .F(n496) );
  IV U768 ( .A(n747), .Z(n338) );
  MUX U769 ( .IN0(n339), .IN1(n850), .SEL(n851), .F(n733) );
  IV U770 ( .A(n852), .Z(n339) );
  MUX U771 ( .IN0(n340), .IN1(n737), .SEL(n738), .F(n490) );
  IV U772 ( .A(n739), .Z(n340) );
  MUX U773 ( .IN0(n1266), .IN1(n341), .SEL(n1267), .F(n1166) );
  IV U774 ( .A(n1268), .Z(n341) );
  MUX U775 ( .IN0(n1468), .IN1(n342), .SEL(n1469), .F(n1372) );
  IV U776 ( .A(n1470), .Z(n342) );
  MUX U777 ( .IN0(n1646), .IN1(n343), .SEL(n1647), .F(n1564) );
  IV U778 ( .A(n1648), .Z(n343) );
  MUX U779 ( .IN0(n1807), .IN1(n344), .SEL(n1808), .F(n1732) );
  IV U780 ( .A(n1809), .Z(n344) );
  MUX U781 ( .IN0(n1951), .IN1(n345), .SEL(n1952), .F(n1885) );
  IV U782 ( .A(n1953), .Z(n345) );
  MUX U783 ( .IN0(n2079), .IN1(n346), .SEL(n2080), .F(n2021) );
  IV U784 ( .A(n2081), .Z(n346) );
  MUX U785 ( .IN0(n2191), .IN1(n347), .SEL(n2192), .F(n2141) );
  IV U786 ( .A(n2193), .Z(n347) );
  MUX U787 ( .IN0(n2288), .IN1(n348), .SEL(n2289), .F(n2246) );
  IV U788 ( .A(n2290), .Z(n348) );
  MUX U789 ( .IN0(n349), .IN1(n2493), .SEL(n2464), .F(n2491) );
  IV U790 ( .A(n2465), .Z(n349) );
  MUX U791 ( .IN0(n350), .IN1(n842), .SEL(n843), .F(n725) );
  IV U792 ( .A(n844), .Z(n350) );
  MUX U793 ( .IN0(n351), .IN1(n729), .SEL(n730), .F(n484) );
  IV U794 ( .A(n731), .Z(n351) );
  MUX U795 ( .IN0(n352), .IN1(n834), .SEL(n835), .F(n717) );
  IV U796 ( .A(n836), .Z(n352) );
  MUX U797 ( .IN0(n353), .IN1(n721), .SEL(n722), .F(n478) );
  IV U798 ( .A(n723), .Z(n353) );
  MUX U799 ( .IN0(n1154), .IN1(n354), .SEL(n1155), .F(n1044) );
  IV U800 ( .A(n1156), .Z(n354) );
  MUX U801 ( .IN0(n1360), .IN1(n355), .SEL(n1361), .F(n1262) );
  IV U802 ( .A(n1362), .Z(n355) );
  MUX U803 ( .IN0(n1552), .IN1(n356), .SEL(n1553), .F(n1464) );
  IV U804 ( .A(n1554), .Z(n356) );
  MUX U805 ( .IN0(n1720), .IN1(n357), .SEL(n1721), .F(n1642) );
  IV U806 ( .A(n1722), .Z(n357) );
  MUX U807 ( .IN0(n1873), .IN1(n358), .SEL(n1874), .F(n1803) );
  IV U808 ( .A(n1875), .Z(n358) );
  MUX U809 ( .IN0(n2009), .IN1(n359), .SEL(n2010), .F(n1947) );
  IV U810 ( .A(n2011), .Z(n359) );
  MUX U811 ( .IN0(n2129), .IN1(n360), .SEL(n2130), .F(n2075) );
  IV U812 ( .A(n2131), .Z(n360) );
  MUX U813 ( .IN0(n2234), .IN1(n361), .SEL(n2235), .F(n2187) );
  IV U814 ( .A(n2236), .Z(n361) );
  MUX U815 ( .IN0(n362), .IN1(n2466), .SEL(n2442), .F(n2462) );
  IV U816 ( .A(n2441), .Z(n362) );
  MUX U817 ( .IN0(n363), .IN1(n826), .SEL(n827), .F(n709) );
  IV U818 ( .A(n828), .Z(n363) );
  MUX U819 ( .IN0(n364), .IN1(n713), .SEL(n714), .F(n472) );
  IV U820 ( .A(n715), .Z(n364) );
  MUX U821 ( .IN0(n365), .IN1(n818), .SEL(n819), .F(n701) );
  IV U822 ( .A(n820), .Z(n365) );
  MUX U823 ( .IN0(n366), .IN1(n705), .SEL(n706), .F(n466) );
  IV U824 ( .A(n707), .Z(n366) );
  MUX U825 ( .IN0(n1250), .IN1(n367), .SEL(n1251), .F(n1150) );
  IV U826 ( .A(n1252), .Z(n367) );
  MUX U827 ( .IN0(n1452), .IN1(n368), .SEL(n1453), .F(n1356) );
  IV U828 ( .A(n1454), .Z(n368) );
  MUX U829 ( .IN0(n1630), .IN1(n369), .SEL(n1631), .F(n1548) );
  IV U830 ( .A(n1632), .Z(n369) );
  MUX U831 ( .IN0(n1791), .IN1(n370), .SEL(n1792), .F(n1716) );
  IV U832 ( .A(n1793), .Z(n370) );
  MUX U833 ( .IN0(n1935), .IN1(n371), .SEL(n1936), .F(n1869) );
  IV U834 ( .A(n1937), .Z(n371) );
  MUX U835 ( .IN0(n2063), .IN1(n372), .SEL(n2064), .F(n2005) );
  IV U836 ( .A(n2065), .Z(n372) );
  MUX U837 ( .IN0(n2175), .IN1(n373), .SEL(n2176), .F(n2125) );
  IV U838 ( .A(n2177), .Z(n373) );
  MUX U839 ( .IN0(n2272), .IN1(n374), .SEL(n2273), .F(n2230) );
  IV U840 ( .A(n2274), .Z(n374) );
  MUX U841 ( .IN0(n375), .IN1(n2443), .SEL(n2423), .F(n2439) );
  IV U842 ( .A(n2422), .Z(n375) );
  MUX U843 ( .IN0(n376), .IN1(n2501), .SEL(n2482), .F(n2499) );
  IV U844 ( .A(n2483), .Z(n376) );
  MUX U845 ( .IN0(n377), .IN1(n810), .SEL(n811), .F(n693) );
  IV U846 ( .A(n812), .Z(n377) );
  MUX U847 ( .IN0(n378), .IN1(n697), .SEL(n698), .F(n460) );
  IV U848 ( .A(n699), .Z(n378) );
  MUX U849 ( .IN0(n912), .IN1(n914), .SEL(n913), .F(n379) );
  IV U850 ( .A(n379), .Z(n801) );
  XNOR U851 ( .A(n2382), .B(n2383), .Z(n2363) );
  MUX U852 ( .IN0(n380), .IN1(n689), .SEL(n690), .F(n454) );
  IV U853 ( .A(n691), .Z(n380) );
  MUX U854 ( .IN0(n1140), .IN1(n1138), .SEL(n1139), .F(n1025) );
  MUX U855 ( .IN0(n1346), .IN1(n1344), .SEL(n1345), .F(n1246) );
  MUX U856 ( .IN0(n1538), .IN1(n1536), .SEL(n1537), .F(n1448) );
  MUX U857 ( .IN0(n1706), .IN1(n1704), .SEL(n1705), .F(n1626) );
  MUX U858 ( .IN0(n1859), .IN1(n1857), .SEL(n1858), .F(n1787) );
  MUX U859 ( .IN0(n1995), .IN1(n1993), .SEL(n1994), .F(n1931) );
  MUX U860 ( .IN0(n2115), .IN1(n2113), .SEL(n2114), .F(n2059) );
  MUX U861 ( .IN0(n2219), .IN1(n2217), .SEL(n2218), .F(n2171) );
  XNOR U862 ( .A(n2387), .B(n2388), .Z(n2369) );
  XNOR U863 ( .A(n683), .B(n682), .Z(n678) );
  XNOR U864 ( .A(n799), .B(n798), .Z(n794) );
  XNOR U865 ( .A(n2372), .B(n2373), .Z(n2357) );
  XNOR U866 ( .A(n396), .B(n395), .Z(n403) );
  MUX U867 ( .IN0(o[27]), .IN1(n902), .SEL(n903), .F(n786) );
  MUX U868 ( .IN0(o[23]), .IN1(n1338), .SEL(n1339), .F(n1236) );
  MUX U869 ( .IN0(o[19]), .IN1(n1698), .SEL(n1699), .F(n1616) );
  MUX U870 ( .IN0(o[15]), .IN1(n1987), .SEL(n1988), .F(n1921) );
  MUX U871 ( .IN0(o[11]), .IN1(n2211), .SEL(n2212), .F(n2161) );
  XNOR U872 ( .A(n2338), .B(n2339), .Z(n2302) );
  XNOR U873 ( .A(n2375), .B(n2376), .Z(n2314) );
  XOR U874 ( .A(n2455), .B(n2456), .Z(n2326) );
  XNOR U875 ( .A(n2304), .B(n2307), .Z(n2305) );
  XNOR U876 ( .A(n2316), .B(n2319), .Z(n2317) );
  XOR U877 ( .A(n2329), .B(n2330), .Z(n784) );
  XNOR U878 ( .A(n381), .B(o[9]), .Z(oi[9]) );
  XNOR U879 ( .A(n382), .B(o[8]), .Z(oi[8]) );
  XNOR U880 ( .A(n383), .B(o[7]), .Z(oi[7]) );
  XNOR U881 ( .A(n384), .B(o[6]), .Z(oi[6]) );
  XNOR U882 ( .A(n385), .B(o[5]), .Z(oi[5]) );
  XNOR U883 ( .A(n386), .B(o[4]), .Z(oi[4]) );
  XNOR U884 ( .A(n387), .B(o[3]), .Z(oi[3]) );
  XOR U885 ( .A(n388), .B(n389), .Z(oi[31]) );
  XOR U886 ( .A(n390), .B(n391), .Z(n389) );
  XOR U887 ( .A(n392), .B(n393), .Z(n391) );
  AND U888 ( .A(e_input[2]), .B(g_input[29]), .Z(n393) );
  ANDN U889 ( .A(n394), .B(n395), .Z(n392) );
  XOR U890 ( .A(n396), .B(n397), .Z(n394) );
  XNOR U891 ( .A(o[31]), .B(n397), .Z(n390) );
  XOR U892 ( .A(n398), .B(n399), .Z(n388) );
  XOR U893 ( .A(n400), .B(n401), .Z(n399) );
  AND U894 ( .A(e_input[1]), .B(g_input[30]), .Z(n401) );
  NOR U895 ( .A(n402), .B(n403), .Z(n400) );
  XOR U896 ( .A(n404), .B(n405), .Z(n398) );
  AND U897 ( .A(g_input[31]), .B(e_input[0]), .Z(n405) );
  XOR U898 ( .A(n406), .B(n407), .Z(n404) );
  XOR U899 ( .A(n408), .B(n409), .Z(n407) );
  XOR U900 ( .A(n410), .B(n411), .Z(n409) );
  ANDN U901 ( .A(n412), .B(n413), .Z(n411) );
  XNOR U902 ( .A(n414), .B(n415), .Z(n412) );
  AND U903 ( .A(e_input[4]), .B(g_input[27]), .Z(n410) );
  XOR U904 ( .A(n416), .B(n417), .Z(n408) );
  ANDN U905 ( .A(n418), .B(n419), .Z(n417) );
  XNOR U906 ( .A(n420), .B(n421), .Z(n418) );
  AND U907 ( .A(n422), .B(n423), .Z(n416) );
  XOR U908 ( .A(o[30]), .B(n424), .Z(n423) );
  XOR U909 ( .A(n425), .B(n424), .Z(n406) );
  XOR U910 ( .A(n426), .B(n427), .Z(n425) );
  AND U911 ( .A(e_input[3]), .B(g_input[28]), .Z(n427) );
  XOR U912 ( .A(n428), .B(n429), .Z(n426) );
  XOR U913 ( .A(n430), .B(n431), .Z(n429) );
  XOR U914 ( .A(n432), .B(n433), .Z(n431) );
  AND U915 ( .A(e_input[5]), .B(g_input[26]), .Z(n433) );
  AND U916 ( .A(n434), .B(n435), .Z(n432) );
  XNOR U917 ( .A(n436), .B(n437), .Z(n435) );
  XOR U918 ( .A(n438), .B(n439), .Z(n430) );
  AND U919 ( .A(e_input[6]), .B(g_input[25]), .Z(n439) );
  AND U920 ( .A(n440), .B(n441), .Z(n438) );
  XNOR U921 ( .A(n442), .B(n443), .Z(n441) );
  XOR U922 ( .A(n444), .B(n445), .Z(n428) );
  XOR U923 ( .A(n446), .B(n447), .Z(n445) );
  XOR U924 ( .A(n448), .B(n449), .Z(n447) );
  XOR U925 ( .A(n437), .B(n443), .Z(n449) );
  XOR U926 ( .A(n450), .B(n451), .Z(n448) );
  XOR U927 ( .A(n452), .B(n453), .Z(n451) );
  XOR U928 ( .A(n454), .B(n455), .Z(n453) );
  XOR U929 ( .A(n456), .B(n457), .Z(n452) );
  XOR U930 ( .A(n458), .B(n459), .Z(n457) );
  XOR U931 ( .A(n460), .B(n461), .Z(n459) );
  XOR U932 ( .A(n462), .B(n463), .Z(n458) );
  XOR U933 ( .A(n464), .B(n465), .Z(n463) );
  XOR U934 ( .A(n466), .B(n467), .Z(n465) );
  XOR U935 ( .A(n468), .B(n469), .Z(n464) );
  XOR U936 ( .A(n470), .B(n471), .Z(n469) );
  XOR U937 ( .A(n472), .B(n473), .Z(n471) );
  XOR U938 ( .A(n474), .B(n475), .Z(n470) );
  XOR U939 ( .A(n476), .B(n477), .Z(n475) );
  XOR U940 ( .A(n478), .B(n479), .Z(n477) );
  XOR U941 ( .A(n480), .B(n481), .Z(n476) );
  XOR U942 ( .A(n482), .B(n483), .Z(n481) );
  XOR U943 ( .A(n484), .B(n485), .Z(n483) );
  XOR U944 ( .A(n486), .B(n487), .Z(n482) );
  XOR U945 ( .A(n488), .B(n489), .Z(n487) );
  XOR U946 ( .A(n490), .B(n491), .Z(n489) );
  XOR U947 ( .A(n492), .B(n493), .Z(n488) );
  XOR U948 ( .A(n494), .B(n495), .Z(n493) );
  XOR U949 ( .A(n496), .B(n497), .Z(n495) );
  XOR U950 ( .A(n498), .B(n499), .Z(n494) );
  XOR U951 ( .A(n500), .B(n501), .Z(n499) );
  XOR U952 ( .A(n502), .B(n503), .Z(n501) );
  XOR U953 ( .A(n504), .B(n505), .Z(n500) );
  XOR U954 ( .A(n506), .B(n507), .Z(n505) );
  XOR U955 ( .A(n508), .B(n509), .Z(n507) );
  XOR U956 ( .A(n510), .B(n511), .Z(n506) );
  XOR U957 ( .A(n512), .B(n513), .Z(n511) );
  XOR U958 ( .A(n514), .B(n515), .Z(n513) );
  XOR U959 ( .A(n516), .B(n517), .Z(n515) );
  XOR U960 ( .A(n518), .B(n519), .Z(n512) );
  AND U961 ( .A(g_input[2]), .B(e_input[29]), .Z(n518) );
  XOR U962 ( .A(n520), .B(n521), .Z(n510) );
  XOR U963 ( .A(n522), .B(n523), .Z(n521) );
  ANDN U964 ( .A(n524), .B(n525), .Z(n523) );
  XNOR U965 ( .A(n526), .B(n519), .Z(n524) );
  AND U966 ( .A(g_input[1]), .B(e_input[30]), .Z(n522) );
  XOR U967 ( .A(n527), .B(n528), .Z(n520) );
  ANDN U968 ( .A(n529), .B(n530), .Z(n528) );
  XOR U969 ( .A(n514), .B(n531), .Z(n529) );
  ANDN U970 ( .A(e_input[31]), .B(n532), .Z(n527) );
  XOR U971 ( .A(n533), .B(n534), .Z(n504) );
  XOR U972 ( .A(n535), .B(n536), .Z(n534) );
  AND U973 ( .A(g_input[4]), .B(e_input[27]), .Z(n536) );
  ANDN U974 ( .A(n537), .B(n538), .Z(n535) );
  XNOR U975 ( .A(n539), .B(n516), .Z(n537) );
  XOR U976 ( .A(n540), .B(n541), .Z(n533) );
  AND U977 ( .A(g_input[3]), .B(e_input[28]), .Z(n541) );
  ANDN U978 ( .A(n542), .B(n543), .Z(n540) );
  XNOR U979 ( .A(n544), .B(n517), .Z(n542) );
  XOR U980 ( .A(n545), .B(n546), .Z(n498) );
  XOR U981 ( .A(n547), .B(n548), .Z(n546) );
  AND U982 ( .A(g_input[6]), .B(e_input[25]), .Z(n548) );
  ANDN U983 ( .A(n549), .B(n550), .Z(n547) );
  XNOR U984 ( .A(n551), .B(n508), .Z(n549) );
  XOR U985 ( .A(n552), .B(n553), .Z(n545) );
  AND U986 ( .A(g_input[5]), .B(e_input[26]), .Z(n553) );
  ANDN U987 ( .A(n554), .B(n555), .Z(n552) );
  XNOR U988 ( .A(n556), .B(n509), .Z(n554) );
  XOR U989 ( .A(n557), .B(n558), .Z(n492) );
  XOR U990 ( .A(n559), .B(n560), .Z(n558) );
  AND U991 ( .A(g_input[8]), .B(e_input[23]), .Z(n560) );
  ANDN U992 ( .A(n561), .B(n562), .Z(n559) );
  XNOR U993 ( .A(n563), .B(n502), .Z(n561) );
  XOR U994 ( .A(n564), .B(n565), .Z(n557) );
  AND U995 ( .A(g_input[7]), .B(e_input[24]), .Z(n565) );
  ANDN U996 ( .A(n566), .B(n567), .Z(n564) );
  XNOR U997 ( .A(n568), .B(n503), .Z(n566) );
  XOR U998 ( .A(n569), .B(n570), .Z(n486) );
  XOR U999 ( .A(n571), .B(n572), .Z(n570) );
  AND U1000 ( .A(g_input[10]), .B(e_input[21]), .Z(n572) );
  ANDN U1001 ( .A(n573), .B(n574), .Z(n571) );
  XNOR U1002 ( .A(n575), .B(n496), .Z(n573) );
  XOR U1003 ( .A(n576), .B(n577), .Z(n569) );
  AND U1004 ( .A(g_input[9]), .B(e_input[22]), .Z(n577) );
  ANDN U1005 ( .A(n578), .B(n579), .Z(n576) );
  XNOR U1006 ( .A(n580), .B(n497), .Z(n578) );
  XOR U1007 ( .A(n581), .B(n582), .Z(n480) );
  XOR U1008 ( .A(n583), .B(n584), .Z(n582) );
  AND U1009 ( .A(g_input[12]), .B(e_input[19]), .Z(n584) );
  ANDN U1010 ( .A(n585), .B(n586), .Z(n583) );
  XNOR U1011 ( .A(n587), .B(n490), .Z(n585) );
  XOR U1012 ( .A(n588), .B(n589), .Z(n581) );
  AND U1013 ( .A(g_input[11]), .B(e_input[20]), .Z(n589) );
  ANDN U1014 ( .A(n590), .B(n591), .Z(n588) );
  XNOR U1015 ( .A(n592), .B(n491), .Z(n590) );
  XOR U1016 ( .A(n593), .B(n594), .Z(n474) );
  XOR U1017 ( .A(n595), .B(n596), .Z(n594) );
  AND U1018 ( .A(g_input[14]), .B(e_input[17]), .Z(n596) );
  ANDN U1019 ( .A(n597), .B(n598), .Z(n595) );
  XNOR U1020 ( .A(n599), .B(n484), .Z(n597) );
  XOR U1021 ( .A(n600), .B(n601), .Z(n593) );
  AND U1022 ( .A(g_input[13]), .B(e_input[18]), .Z(n601) );
  ANDN U1023 ( .A(n602), .B(n603), .Z(n600) );
  XNOR U1024 ( .A(n604), .B(n485), .Z(n602) );
  XOR U1025 ( .A(n605), .B(n606), .Z(n468) );
  XOR U1026 ( .A(n607), .B(n608), .Z(n606) );
  AND U1027 ( .A(g_input[16]), .B(e_input[15]), .Z(n608) );
  ANDN U1028 ( .A(n609), .B(n610), .Z(n607) );
  XNOR U1029 ( .A(n611), .B(n478), .Z(n609) );
  XOR U1030 ( .A(n612), .B(n613), .Z(n605) );
  AND U1031 ( .A(g_input[15]), .B(e_input[16]), .Z(n613) );
  ANDN U1032 ( .A(n614), .B(n615), .Z(n612) );
  XNOR U1033 ( .A(n616), .B(n479), .Z(n614) );
  XOR U1034 ( .A(n617), .B(n618), .Z(n462) );
  XOR U1035 ( .A(n619), .B(n620), .Z(n618) );
  AND U1036 ( .A(g_input[18]), .B(e_input[13]), .Z(n620) );
  ANDN U1037 ( .A(n621), .B(n622), .Z(n619) );
  XNOR U1038 ( .A(n623), .B(n472), .Z(n621) );
  XOR U1039 ( .A(n624), .B(n625), .Z(n617) );
  AND U1040 ( .A(g_input[17]), .B(e_input[14]), .Z(n625) );
  ANDN U1041 ( .A(n626), .B(n627), .Z(n624) );
  XNOR U1042 ( .A(n628), .B(n473), .Z(n626) );
  XOR U1043 ( .A(n629), .B(n630), .Z(n456) );
  XOR U1044 ( .A(n631), .B(n632), .Z(n630) );
  AND U1045 ( .A(g_input[20]), .B(e_input[11]), .Z(n632) );
  ANDN U1046 ( .A(n633), .B(n634), .Z(n631) );
  XNOR U1047 ( .A(n635), .B(n466), .Z(n633) );
  XOR U1048 ( .A(n636), .B(n637), .Z(n629) );
  AND U1049 ( .A(g_input[19]), .B(e_input[12]), .Z(n637) );
  ANDN U1050 ( .A(n638), .B(n639), .Z(n636) );
  XNOR U1051 ( .A(n640), .B(n467), .Z(n638) );
  XOR U1052 ( .A(n641), .B(n642), .Z(n450) );
  XOR U1053 ( .A(n643), .B(n644), .Z(n642) );
  AND U1054 ( .A(e_input[9]), .B(g_input[22]), .Z(n644) );
  ANDN U1055 ( .A(n645), .B(n646), .Z(n643) );
  XNOR U1056 ( .A(n647), .B(n460), .Z(n645) );
  XOR U1057 ( .A(n648), .B(n649), .Z(n641) );
  AND U1058 ( .A(g_input[21]), .B(e_input[10]), .Z(n649) );
  ANDN U1059 ( .A(n650), .B(n651), .Z(n648) );
  XNOR U1060 ( .A(n652), .B(n461), .Z(n650) );
  XOR U1061 ( .A(n653), .B(n654), .Z(n446) );
  XOR U1062 ( .A(n655), .B(n656), .Z(n654) );
  AND U1063 ( .A(e_input[7]), .B(g_input[24]), .Z(n656) );
  AND U1064 ( .A(n657), .B(n658), .Z(n655) );
  XNOR U1065 ( .A(n659), .B(n454), .Z(n658) );
  XOR U1066 ( .A(n660), .B(n661), .Z(n653) );
  AND U1067 ( .A(e_input[8]), .B(g_input[23]), .Z(n661) );
  AND U1068 ( .A(n662), .B(n663), .Z(n660) );
  XNOR U1069 ( .A(n664), .B(n455), .Z(n663) );
  XNOR U1070 ( .A(n421), .B(n415), .Z(n444) );
  XOR U1071 ( .A(n422), .B(o[30]), .Z(oi[30]) );
  XOR U1072 ( .A(n665), .B(n424), .Z(n422) );
  XOR U1073 ( .A(n403), .B(n402), .Z(n665) );
  NAND U1074 ( .A(g_input[30]), .B(e_input[0]), .Z(n402) );
  XNOR U1075 ( .A(n668), .B(n397), .Z(n395) );
  NANDN U1076 ( .B(n669), .A(n670), .Z(n397) );
  NAND U1077 ( .A(e_input[1]), .B(g_input[29]), .Z(n668) );
  XNOR U1078 ( .A(n415), .B(n671), .Z(n413) );
  AND U1079 ( .A(e_input[2]), .B(g_input[28]), .Z(n671) );
  XNOR U1080 ( .A(n420), .B(n419), .Z(n414) );
  XNOR U1081 ( .A(n421), .B(n675), .Z(n419) );
  AND U1082 ( .A(e_input[3]), .B(g_input[27]), .Z(n675) );
  XOR U1083 ( .A(n436), .B(n434), .Z(n420) );
  XOR U1084 ( .A(n437), .B(n679), .Z(n434) );
  AND U1085 ( .A(e_input[4]), .B(g_input[26]), .Z(n679) );
  XNOR U1086 ( .A(n683), .B(n680), .Z(n681) );
  XOR U1087 ( .A(n442), .B(n440), .Z(n436) );
  XOR U1088 ( .A(n443), .B(n684), .Z(n440) );
  AND U1089 ( .A(e_input[5]), .B(g_input[25]), .Z(n684) );
  XOR U1090 ( .A(n659), .B(n657), .Z(n442) );
  XOR U1091 ( .A(n454), .B(n688), .Z(n657) );
  AND U1092 ( .A(e_input[6]), .B(g_input[24]), .Z(n688) );
  XOR U1093 ( .A(n664), .B(n662), .Z(n659) );
  XOR U1094 ( .A(n455), .B(n692), .Z(n662) );
  AND U1095 ( .A(e_input[7]), .B(g_input[23]), .Z(n692) );
  XNOR U1096 ( .A(n647), .B(n646), .Z(n664) );
  XNOR U1097 ( .A(n460), .B(n696), .Z(n646) );
  AND U1098 ( .A(e_input[8]), .B(g_input[22]), .Z(n696) );
  XNOR U1099 ( .A(n652), .B(n651), .Z(n647) );
  XNOR U1100 ( .A(n461), .B(n700), .Z(n651) );
  AND U1101 ( .A(e_input[9]), .B(g_input[21]), .Z(n700) );
  XNOR U1102 ( .A(n635), .B(n634), .Z(n652) );
  XNOR U1103 ( .A(n466), .B(n704), .Z(n634) );
  AND U1104 ( .A(g_input[20]), .B(e_input[10]), .Z(n704) );
  XNOR U1105 ( .A(n640), .B(n639), .Z(n635) );
  XNOR U1106 ( .A(n467), .B(n708), .Z(n639) );
  AND U1107 ( .A(g_input[19]), .B(e_input[11]), .Z(n708) );
  XNOR U1108 ( .A(n623), .B(n622), .Z(n640) );
  XNOR U1109 ( .A(n472), .B(n712), .Z(n622) );
  AND U1110 ( .A(g_input[18]), .B(e_input[12]), .Z(n712) );
  XNOR U1111 ( .A(n628), .B(n627), .Z(n623) );
  XNOR U1112 ( .A(n473), .B(n716), .Z(n627) );
  AND U1113 ( .A(g_input[17]), .B(e_input[13]), .Z(n716) );
  XNOR U1114 ( .A(n611), .B(n610), .Z(n628) );
  XNOR U1115 ( .A(n478), .B(n720), .Z(n610) );
  AND U1116 ( .A(g_input[16]), .B(e_input[14]), .Z(n720) );
  XNOR U1117 ( .A(n616), .B(n615), .Z(n611) );
  XNOR U1118 ( .A(n479), .B(n724), .Z(n615) );
  AND U1119 ( .A(g_input[15]), .B(e_input[15]), .Z(n724) );
  XNOR U1120 ( .A(n599), .B(n598), .Z(n616) );
  XNOR U1121 ( .A(n484), .B(n728), .Z(n598) );
  AND U1122 ( .A(g_input[14]), .B(e_input[16]), .Z(n728) );
  XNOR U1123 ( .A(n604), .B(n603), .Z(n599) );
  XNOR U1124 ( .A(n485), .B(n732), .Z(n603) );
  AND U1125 ( .A(g_input[13]), .B(e_input[17]), .Z(n732) );
  XNOR U1126 ( .A(n587), .B(n586), .Z(n604) );
  XNOR U1127 ( .A(n490), .B(n736), .Z(n586) );
  AND U1128 ( .A(g_input[12]), .B(e_input[18]), .Z(n736) );
  XNOR U1129 ( .A(n592), .B(n591), .Z(n587) );
  XNOR U1130 ( .A(n491), .B(n740), .Z(n591) );
  AND U1131 ( .A(g_input[11]), .B(e_input[19]), .Z(n740) );
  XNOR U1132 ( .A(n575), .B(n574), .Z(n592) );
  XNOR U1133 ( .A(n496), .B(n744), .Z(n574) );
  AND U1134 ( .A(g_input[10]), .B(e_input[20]), .Z(n744) );
  XNOR U1135 ( .A(n580), .B(n579), .Z(n575) );
  XNOR U1136 ( .A(n497), .B(n748), .Z(n579) );
  AND U1137 ( .A(g_input[9]), .B(e_input[21]), .Z(n748) );
  XNOR U1138 ( .A(n563), .B(n562), .Z(n580) );
  XNOR U1139 ( .A(n502), .B(n752), .Z(n562) );
  AND U1140 ( .A(g_input[8]), .B(e_input[22]), .Z(n752) );
  XNOR U1141 ( .A(n568), .B(n567), .Z(n563) );
  XNOR U1142 ( .A(n503), .B(n756), .Z(n567) );
  AND U1143 ( .A(g_input[7]), .B(e_input[23]), .Z(n756) );
  XNOR U1144 ( .A(n551), .B(n550), .Z(n568) );
  XNOR U1145 ( .A(n508), .B(n760), .Z(n550) );
  AND U1146 ( .A(g_input[6]), .B(e_input[24]), .Z(n760) );
  XNOR U1147 ( .A(n556), .B(n555), .Z(n551) );
  XNOR U1148 ( .A(n509), .B(n764), .Z(n555) );
  AND U1149 ( .A(g_input[5]), .B(e_input[25]), .Z(n764) );
  XNOR U1150 ( .A(n539), .B(n538), .Z(n556) );
  XNOR U1151 ( .A(n516), .B(n768), .Z(n538) );
  AND U1152 ( .A(g_input[4]), .B(e_input[26]), .Z(n768) );
  XNOR U1153 ( .A(n544), .B(n543), .Z(n539) );
  XNOR U1154 ( .A(n517), .B(n772), .Z(n543) );
  AND U1155 ( .A(g_input[3]), .B(e_input[27]), .Z(n772) );
  XNOR U1156 ( .A(n526), .B(n525), .Z(n544) );
  XNOR U1157 ( .A(n519), .B(n776), .Z(n525) );
  AND U1158 ( .A(g_input[2]), .B(e_input[28]), .Z(n776) );
  XNOR U1159 ( .A(n530), .B(n531), .Z(n526) );
  NANDN U1160 ( .B(n532), .A(e_input[30]), .Z(n531) );
  XOR U1161 ( .A(n514), .B(n780), .Z(n530) );
  AND U1162 ( .A(g_input[1]), .B(e_input[29]), .Z(n780) );
  XOR U1163 ( .A(o[2]), .B(n784), .Z(oi[2]) );
  XNOR U1164 ( .A(n667), .B(o[29]), .Z(oi[29]) );
  XNOR U1165 ( .A(n785), .B(n666), .Z(n667) );
  XNOR U1166 ( .A(n670), .B(n669), .Z(n785) );
  NAND U1167 ( .A(g_input[29]), .B(e_input[0]), .Z(n669) );
  XOR U1168 ( .A(n674), .B(n673), .Z(n670) );
  XOR U1169 ( .A(n788), .B(n672), .Z(n673) );
  ANDN U1170 ( .A(n789), .B(n790), .Z(n672) );
  NAND U1171 ( .A(e_input[1]), .B(g_input[28]), .Z(n788) );
  XOR U1172 ( .A(n678), .B(n677), .Z(n674) );
  XNOR U1173 ( .A(n676), .B(n791), .Z(n677) );
  AND U1174 ( .A(e_input[2]), .B(g_input[27]), .Z(n791) );
  XNOR U1175 ( .A(n680), .B(n795), .Z(n682) );
  AND U1176 ( .A(e_input[3]), .B(g_input[26]), .Z(n795) );
  XNOR U1177 ( .A(n799), .B(n796), .Z(n797) );
  XNOR U1178 ( .A(n685), .B(n800), .Z(n686) );
  AND U1179 ( .A(e_input[4]), .B(g_input[25]), .Z(n800) );
  XNOR U1180 ( .A(n689), .B(n804), .Z(n690) );
  AND U1181 ( .A(e_input[5]), .B(g_input[24]), .Z(n804) );
  XNOR U1182 ( .A(n808), .B(n805), .Z(n806) );
  XNOR U1183 ( .A(n693), .B(n809), .Z(n694) );
  AND U1184 ( .A(e_input[6]), .B(g_input[23]), .Z(n809) );
  XNOR U1185 ( .A(n697), .B(n813), .Z(n698) );
  AND U1186 ( .A(e_input[7]), .B(g_input[22]), .Z(n813) );
  XNOR U1187 ( .A(n701), .B(n817), .Z(n702) );
  AND U1188 ( .A(e_input[8]), .B(g_input[21]), .Z(n817) );
  XNOR U1189 ( .A(n705), .B(n821), .Z(n706) );
  AND U1190 ( .A(e_input[9]), .B(g_input[20]), .Z(n821) );
  XNOR U1191 ( .A(n709), .B(n825), .Z(n710) );
  AND U1192 ( .A(g_input[19]), .B(e_input[10]), .Z(n825) );
  XNOR U1193 ( .A(n713), .B(n829), .Z(n714) );
  AND U1194 ( .A(g_input[18]), .B(e_input[11]), .Z(n829) );
  XNOR U1195 ( .A(n717), .B(n833), .Z(n718) );
  AND U1196 ( .A(g_input[17]), .B(e_input[12]), .Z(n833) );
  XNOR U1197 ( .A(n721), .B(n837), .Z(n722) );
  AND U1198 ( .A(g_input[16]), .B(e_input[13]), .Z(n837) );
  XNOR U1199 ( .A(n725), .B(n841), .Z(n726) );
  AND U1200 ( .A(g_input[15]), .B(e_input[14]), .Z(n841) );
  XNOR U1201 ( .A(n729), .B(n845), .Z(n730) );
  AND U1202 ( .A(g_input[14]), .B(e_input[15]), .Z(n845) );
  XNOR U1203 ( .A(n733), .B(n849), .Z(n734) );
  AND U1204 ( .A(g_input[13]), .B(e_input[16]), .Z(n849) );
  XNOR U1205 ( .A(n737), .B(n853), .Z(n738) );
  AND U1206 ( .A(g_input[12]), .B(e_input[17]), .Z(n853) );
  XNOR U1207 ( .A(n741), .B(n857), .Z(n742) );
  AND U1208 ( .A(g_input[11]), .B(e_input[18]), .Z(n857) );
  XNOR U1209 ( .A(n745), .B(n861), .Z(n746) );
  AND U1210 ( .A(g_input[10]), .B(e_input[19]), .Z(n861) );
  XNOR U1211 ( .A(n749), .B(n865), .Z(n750) );
  AND U1212 ( .A(g_input[9]), .B(e_input[20]), .Z(n865) );
  XNOR U1213 ( .A(n753), .B(n869), .Z(n754) );
  AND U1214 ( .A(g_input[8]), .B(e_input[21]), .Z(n869) );
  XNOR U1215 ( .A(n757), .B(n873), .Z(n758) );
  AND U1216 ( .A(g_input[7]), .B(e_input[22]), .Z(n873) );
  XNOR U1217 ( .A(n761), .B(n877), .Z(n762) );
  AND U1218 ( .A(g_input[6]), .B(e_input[23]), .Z(n877) );
  XNOR U1219 ( .A(n765), .B(n881), .Z(n766) );
  AND U1220 ( .A(g_input[5]), .B(e_input[24]), .Z(n881) );
  XNOR U1221 ( .A(n769), .B(n885), .Z(n770) );
  AND U1222 ( .A(g_input[4]), .B(e_input[25]), .Z(n885) );
  XNOR U1223 ( .A(n773), .B(n889), .Z(n774) );
  AND U1224 ( .A(g_input[3]), .B(e_input[26]), .Z(n889) );
  XNOR U1225 ( .A(n779), .B(n778), .Z(n775) );
  XNOR U1226 ( .A(n777), .B(n893), .Z(n778) );
  AND U1227 ( .A(g_input[2]), .B(e_input[27]), .Z(n893) );
  XNOR U1228 ( .A(n782), .B(n783), .Z(n779) );
  NANDN U1229 ( .B(n532), .A(e_input[29]), .Z(n783) );
  XNOR U1230 ( .A(n781), .B(n897), .Z(n782) );
  AND U1231 ( .A(g_input[1]), .B(e_input[28]), .Z(n897) );
  XNOR U1232 ( .A(n787), .B(o[28]), .Z(oi[28]) );
  XNOR U1233 ( .A(n901), .B(n786), .Z(n787) );
  XNOR U1234 ( .A(n789), .B(n790), .Z(n901) );
  NAND U1235 ( .A(g_input[28]), .B(e_input[0]), .Z(n790) );
  XOR U1236 ( .A(n794), .B(n793), .Z(n789) );
  XNOR U1237 ( .A(n904), .B(n792), .Z(n793) );
  NANDN U1238 ( .B(n905), .A(n906), .Z(n792) );
  NAND U1239 ( .A(e_input[1]), .B(g_input[27]), .Z(n904) );
  XNOR U1240 ( .A(n796), .B(n907), .Z(n798) );
  AND U1241 ( .A(e_input[2]), .B(g_input[26]), .Z(n907) );
  XNOR U1242 ( .A(n801), .B(n911), .Z(n802) );
  AND U1243 ( .A(e_input[3]), .B(g_input[25]), .Z(n911) );
  XNOR U1244 ( .A(n805), .B(n915), .Z(n807) );
  AND U1245 ( .A(e_input[4]), .B(g_input[24]), .Z(n915) );
  XOR U1246 ( .A(n916), .B(n917), .Z(n805) );
  AND U1247 ( .A(n918), .B(n919), .Z(n917) );
  XNOR U1248 ( .A(n920), .B(n916), .Z(n919) );
  XNOR U1249 ( .A(n810), .B(n921), .Z(n811) );
  AND U1250 ( .A(e_input[5]), .B(g_input[23]), .Z(n921) );
  XNOR U1251 ( .A(n814), .B(n925), .Z(n815) );
  AND U1252 ( .A(e_input[6]), .B(g_input[22]), .Z(n925) );
  XNOR U1253 ( .A(n818), .B(n929), .Z(n819) );
  AND U1254 ( .A(e_input[7]), .B(g_input[21]), .Z(n929) );
  XNOR U1255 ( .A(n822), .B(n933), .Z(n823) );
  AND U1256 ( .A(e_input[8]), .B(g_input[20]), .Z(n933) );
  XOR U1257 ( .A(n828), .B(n937), .Z(n824) );
  IV U1258 ( .A(n827), .Z(n937) );
  XNOR U1259 ( .A(n826), .B(n938), .Z(n827) );
  AND U1260 ( .A(e_input[9]), .B(g_input[19]), .Z(n938) );
  XNOR U1261 ( .A(n830), .B(n942), .Z(n831) );
  AND U1262 ( .A(g_input[18]), .B(e_input[10]), .Z(n942) );
  XNOR U1263 ( .A(n834), .B(n946), .Z(n835) );
  AND U1264 ( .A(g_input[17]), .B(e_input[11]), .Z(n946) );
  XNOR U1265 ( .A(n838), .B(n950), .Z(n839) );
  AND U1266 ( .A(g_input[16]), .B(e_input[12]), .Z(n950) );
  XNOR U1267 ( .A(n842), .B(n954), .Z(n843) );
  AND U1268 ( .A(g_input[15]), .B(e_input[13]), .Z(n954) );
  XNOR U1269 ( .A(n846), .B(n958), .Z(n847) );
  AND U1270 ( .A(g_input[14]), .B(e_input[14]), .Z(n958) );
  XNOR U1271 ( .A(n850), .B(n962), .Z(n851) );
  AND U1272 ( .A(g_input[13]), .B(e_input[15]), .Z(n962) );
  XNOR U1273 ( .A(n854), .B(n966), .Z(n855) );
  AND U1274 ( .A(g_input[12]), .B(e_input[16]), .Z(n966) );
  XNOR U1275 ( .A(n858), .B(n970), .Z(n859) );
  AND U1276 ( .A(g_input[11]), .B(e_input[17]), .Z(n970) );
  XNOR U1277 ( .A(n862), .B(n974), .Z(n863) );
  AND U1278 ( .A(g_input[10]), .B(e_input[18]), .Z(n974) );
  XNOR U1279 ( .A(n866), .B(n978), .Z(n867) );
  AND U1280 ( .A(g_input[9]), .B(e_input[19]), .Z(n978) );
  XNOR U1281 ( .A(n870), .B(n982), .Z(n871) );
  AND U1282 ( .A(g_input[8]), .B(e_input[20]), .Z(n982) );
  XNOR U1283 ( .A(n874), .B(n986), .Z(n875) );
  AND U1284 ( .A(g_input[7]), .B(e_input[21]), .Z(n986) );
  XNOR U1285 ( .A(n878), .B(n990), .Z(n879) );
  AND U1286 ( .A(g_input[6]), .B(e_input[22]), .Z(n990) );
  XNOR U1287 ( .A(n882), .B(n994), .Z(n883) );
  AND U1288 ( .A(g_input[5]), .B(e_input[23]), .Z(n994) );
  XNOR U1289 ( .A(n886), .B(n998), .Z(n887) );
  AND U1290 ( .A(g_input[4]), .B(e_input[24]), .Z(n998) );
  XNOR U1291 ( .A(n890), .B(n1002), .Z(n891) );
  AND U1292 ( .A(g_input[3]), .B(e_input[25]), .Z(n1002) );
  XNOR U1293 ( .A(n896), .B(n895), .Z(n892) );
  XNOR U1294 ( .A(n894), .B(n1006), .Z(n895) );
  AND U1295 ( .A(g_input[2]), .B(e_input[26]), .Z(n1006) );
  XNOR U1296 ( .A(n899), .B(n900), .Z(n896) );
  NANDN U1297 ( .B(n532), .A(e_input[28]), .Z(n900) );
  XNOR U1298 ( .A(n898), .B(n1010), .Z(n899) );
  AND U1299 ( .A(g_input[1]), .B(e_input[27]), .Z(n1010) );
  XNOR U1300 ( .A(n903), .B(o[27]), .Z(oi[27]) );
  XNOR U1301 ( .A(n1014), .B(n902), .Z(n903) );
  XNOR U1302 ( .A(n906), .B(n905), .Z(n1014) );
  NAND U1303 ( .A(g_input[27]), .B(e_input[0]), .Z(n905) );
  XOR U1304 ( .A(n910), .B(n909), .Z(n906) );
  XOR U1305 ( .A(n1017), .B(n908), .Z(n909) );
  ANDN U1306 ( .A(n1018), .B(n1019), .Z(n908) );
  NAND U1307 ( .A(e_input[1]), .B(g_input[26]), .Z(n1017) );
  XOR U1308 ( .A(n914), .B(n913), .Z(n910) );
  XNOR U1309 ( .A(n912), .B(n1020), .Z(n913) );
  AND U1310 ( .A(e_input[2]), .B(g_input[25]), .Z(n1020) );
  XOR U1311 ( .A(n920), .B(n918), .Z(n914) );
  XOR U1312 ( .A(n916), .B(n1024), .Z(n918) );
  AND U1313 ( .A(e_input[3]), .B(g_input[24]), .Z(n1024) );
  XOR U1314 ( .A(n924), .B(n923), .Z(n920) );
  XOR U1315 ( .A(n922), .B(n1028), .Z(n923) );
  AND U1316 ( .A(e_input[4]), .B(g_input[23]), .Z(n1028) );
  XNOR U1317 ( .A(n1032), .B(n1029), .Z(n1031) );
  XOR U1318 ( .A(n928), .B(n927), .Z(n924) );
  XOR U1319 ( .A(n926), .B(n1033), .Z(n927) );
  AND U1320 ( .A(e_input[5]), .B(g_input[22]), .Z(n1033) );
  XOR U1321 ( .A(n932), .B(n931), .Z(n928) );
  XOR U1322 ( .A(n930), .B(n1037), .Z(n931) );
  AND U1323 ( .A(e_input[6]), .B(g_input[21]), .Z(n1037) );
  XOR U1324 ( .A(n1038), .B(n1039), .Z(n930) );
  AND U1325 ( .A(n1040), .B(n1041), .Z(n1039) );
  XNOR U1326 ( .A(n1042), .B(n1038), .Z(n1041) );
  XOR U1327 ( .A(n936), .B(n935), .Z(n932) );
  XOR U1328 ( .A(n934), .B(n1043), .Z(n935) );
  AND U1329 ( .A(e_input[7]), .B(g_input[20]), .Z(n1043) );
  XOR U1330 ( .A(n941), .B(n940), .Z(n936) );
  XOR U1331 ( .A(n939), .B(n1047), .Z(n940) );
  AND U1332 ( .A(e_input[8]), .B(g_input[19]), .Z(n1047) );
  XOR U1333 ( .A(n945), .B(n944), .Z(n941) );
  XOR U1334 ( .A(n943), .B(n1051), .Z(n944) );
  AND U1335 ( .A(e_input[9]), .B(g_input[18]), .Z(n1051) );
  XOR U1336 ( .A(n1052), .B(n1053), .Z(n943) );
  AND U1337 ( .A(n1054), .B(n1055), .Z(n1053) );
  XNOR U1338 ( .A(n1056), .B(n1052), .Z(n1055) );
  XOR U1339 ( .A(n949), .B(n948), .Z(n945) );
  XOR U1340 ( .A(n947), .B(n1057), .Z(n948) );
  AND U1341 ( .A(g_input[17]), .B(e_input[10]), .Z(n1057) );
  XOR U1342 ( .A(n953), .B(n952), .Z(n949) );
  XOR U1343 ( .A(n951), .B(n1061), .Z(n952) );
  AND U1344 ( .A(g_input[16]), .B(e_input[11]), .Z(n1061) );
  XOR U1345 ( .A(n957), .B(n956), .Z(n953) );
  XOR U1346 ( .A(n955), .B(n1065), .Z(n956) );
  AND U1347 ( .A(g_input[15]), .B(e_input[12]), .Z(n1065) );
  XOR U1348 ( .A(n1066), .B(n1067), .Z(n955) );
  AND U1349 ( .A(n1068), .B(n1069), .Z(n1067) );
  XNOR U1350 ( .A(n1070), .B(n1066), .Z(n1069) );
  XOR U1351 ( .A(n961), .B(n960), .Z(n957) );
  XOR U1352 ( .A(n959), .B(n1071), .Z(n960) );
  AND U1353 ( .A(g_input[14]), .B(e_input[13]), .Z(n1071) );
  XOR U1354 ( .A(n965), .B(n964), .Z(n961) );
  XOR U1355 ( .A(n963), .B(n1075), .Z(n964) );
  AND U1356 ( .A(g_input[13]), .B(e_input[14]), .Z(n1075) );
  XOR U1357 ( .A(n969), .B(n968), .Z(n965) );
  XOR U1358 ( .A(n967), .B(n1079), .Z(n968) );
  AND U1359 ( .A(g_input[12]), .B(e_input[15]), .Z(n1079) );
  XOR U1360 ( .A(n973), .B(n972), .Z(n969) );
  XOR U1361 ( .A(n971), .B(n1083), .Z(n972) );
  AND U1362 ( .A(g_input[11]), .B(e_input[16]), .Z(n1083) );
  XOR U1363 ( .A(n1084), .B(n1085), .Z(n971) );
  AND U1364 ( .A(n1086), .B(n1087), .Z(n1085) );
  XNOR U1365 ( .A(n1088), .B(n1084), .Z(n1087) );
  XOR U1366 ( .A(n977), .B(n976), .Z(n973) );
  XOR U1367 ( .A(n975), .B(n1089), .Z(n976) );
  AND U1368 ( .A(g_input[10]), .B(e_input[17]), .Z(n1089) );
  XOR U1369 ( .A(n981), .B(n980), .Z(n977) );
  XOR U1370 ( .A(n979), .B(n1093), .Z(n980) );
  AND U1371 ( .A(g_input[9]), .B(e_input[18]), .Z(n1093) );
  XOR U1372 ( .A(n985), .B(n984), .Z(n981) );
  XOR U1373 ( .A(n983), .B(n1097), .Z(n984) );
  AND U1374 ( .A(g_input[8]), .B(e_input[19]), .Z(n1097) );
  XOR U1375 ( .A(n989), .B(n988), .Z(n985) );
  XOR U1376 ( .A(n987), .B(n1101), .Z(n988) );
  AND U1377 ( .A(g_input[7]), .B(e_input[20]), .Z(n1101) );
  XOR U1378 ( .A(n1102), .B(n1103), .Z(n987) );
  AND U1379 ( .A(n1104), .B(n1105), .Z(n1103) );
  XNOR U1380 ( .A(n1106), .B(n1102), .Z(n1105) );
  XOR U1381 ( .A(n993), .B(n992), .Z(n989) );
  XOR U1382 ( .A(n991), .B(n1107), .Z(n992) );
  AND U1383 ( .A(g_input[6]), .B(e_input[21]), .Z(n1107) );
  XOR U1384 ( .A(n997), .B(n996), .Z(n993) );
  XOR U1385 ( .A(n995), .B(n1111), .Z(n996) );
  AND U1386 ( .A(g_input[5]), .B(e_input[22]), .Z(n1111) );
  XOR U1387 ( .A(n1001), .B(n1000), .Z(n997) );
  XOR U1388 ( .A(n999), .B(n1115), .Z(n1000) );
  AND U1389 ( .A(g_input[4]), .B(e_input[23]), .Z(n1115) );
  XOR U1390 ( .A(n1005), .B(n1004), .Z(n1001) );
  XOR U1391 ( .A(n1003), .B(n1119), .Z(n1004) );
  AND U1392 ( .A(g_input[3]), .B(e_input[24]), .Z(n1119) );
  XNOR U1393 ( .A(n1009), .B(n1008), .Z(n1005) );
  XOR U1394 ( .A(n1007), .B(n1123), .Z(n1008) );
  AND U1395 ( .A(g_input[2]), .B(e_input[25]), .Z(n1123) );
  XOR U1396 ( .A(n1012), .B(n1013), .Z(n1009) );
  NANDN U1397 ( .B(n532), .A(e_input[27]), .Z(n1013) );
  XNOR U1398 ( .A(n1011), .B(n1127), .Z(n1012) );
  AND U1399 ( .A(g_input[1]), .B(e_input[26]), .Z(n1127) );
  XNOR U1400 ( .A(n1016), .B(o[26]), .Z(oi[26]) );
  XNOR U1401 ( .A(n1131), .B(n1015), .Z(n1016) );
  XNOR U1402 ( .A(n1018), .B(n1019), .Z(n1131) );
  NAND U1403 ( .A(g_input[26]), .B(e_input[0]), .Z(n1019) );
  XOR U1404 ( .A(n1023), .B(n1022), .Z(n1018) );
  XNOR U1405 ( .A(n1134), .B(n1021), .Z(n1022) );
  NANDN U1406 ( .B(n1135), .A(n1136), .Z(n1021) );
  NAND U1407 ( .A(e_input[1]), .B(g_input[25]), .Z(n1134) );
  XOR U1408 ( .A(n1027), .B(n1026), .Z(n1023) );
  XNOR U1409 ( .A(n1025), .B(n1137), .Z(n1026) );
  AND U1410 ( .A(e_input[2]), .B(g_input[24]), .Z(n1137) );
  XOR U1411 ( .A(n1032), .B(n1030), .Z(n1027) );
  XOR U1412 ( .A(n1029), .B(n1141), .Z(n1030) );
  AND U1413 ( .A(e_input[3]), .B(g_input[23]), .Z(n1141) );
  XOR U1414 ( .A(n1036), .B(n1035), .Z(n1032) );
  XOR U1415 ( .A(n1034), .B(n1145), .Z(n1035) );
  AND U1416 ( .A(e_input[4]), .B(g_input[22]), .Z(n1145) );
  XOR U1417 ( .A(n1042), .B(n1040), .Z(n1036) );
  XOR U1418 ( .A(n1038), .B(n1149), .Z(n1040) );
  AND U1419 ( .A(e_input[5]), .B(g_input[21]), .Z(n1149) );
  XOR U1420 ( .A(n1046), .B(n1045), .Z(n1042) );
  XOR U1421 ( .A(n1044), .B(n1153), .Z(n1045) );
  AND U1422 ( .A(e_input[6]), .B(g_input[20]), .Z(n1153) );
  XOR U1423 ( .A(n1050), .B(n1049), .Z(n1046) );
  XOR U1424 ( .A(n1048), .B(n1157), .Z(n1049) );
  AND U1425 ( .A(e_input[7]), .B(g_input[19]), .Z(n1157) );
  XOR U1426 ( .A(n1056), .B(n1054), .Z(n1050) );
  XOR U1427 ( .A(n1052), .B(n1161), .Z(n1054) );
  AND U1428 ( .A(e_input[8]), .B(g_input[18]), .Z(n1161) );
  XOR U1429 ( .A(n1060), .B(n1059), .Z(n1056) );
  XOR U1430 ( .A(n1058), .B(n1165), .Z(n1059) );
  AND U1431 ( .A(e_input[9]), .B(g_input[17]), .Z(n1165) );
  XOR U1432 ( .A(n1166), .B(n1167), .Z(n1058) );
  AND U1433 ( .A(n1168), .B(n1169), .Z(n1167) );
  XNOR U1434 ( .A(n1170), .B(n1166), .Z(n1169) );
  XOR U1435 ( .A(n1064), .B(n1063), .Z(n1060) );
  XOR U1436 ( .A(n1062), .B(n1171), .Z(n1063) );
  AND U1437 ( .A(g_input[16]), .B(e_input[10]), .Z(n1171) );
  XOR U1438 ( .A(n1070), .B(n1068), .Z(n1064) );
  XOR U1439 ( .A(n1066), .B(n1175), .Z(n1068) );
  AND U1440 ( .A(g_input[15]), .B(e_input[11]), .Z(n1175) );
  XOR U1441 ( .A(n1074), .B(n1073), .Z(n1070) );
  XOR U1442 ( .A(n1072), .B(n1179), .Z(n1073) );
  AND U1443 ( .A(g_input[14]), .B(e_input[12]), .Z(n1179) );
  XOR U1444 ( .A(n1078), .B(n1077), .Z(n1074) );
  XOR U1445 ( .A(n1076), .B(n1183), .Z(n1077) );
  AND U1446 ( .A(g_input[13]), .B(e_input[13]), .Z(n1183) );
  XOR U1447 ( .A(n1082), .B(n1081), .Z(n1078) );
  XOR U1448 ( .A(n1080), .B(n1187), .Z(n1081) );
  AND U1449 ( .A(g_input[12]), .B(e_input[14]), .Z(n1187) );
  XOR U1450 ( .A(n1088), .B(n1086), .Z(n1082) );
  XOR U1451 ( .A(n1084), .B(n1191), .Z(n1086) );
  AND U1452 ( .A(g_input[11]), .B(e_input[15]), .Z(n1191) );
  XOR U1453 ( .A(n1092), .B(n1091), .Z(n1088) );
  XOR U1454 ( .A(n1090), .B(n1195), .Z(n1091) );
  AND U1455 ( .A(g_input[10]), .B(e_input[16]), .Z(n1195) );
  XOR U1456 ( .A(n1096), .B(n1095), .Z(n1092) );
  XOR U1457 ( .A(n1094), .B(n1199), .Z(n1095) );
  AND U1458 ( .A(g_input[9]), .B(e_input[17]), .Z(n1199) );
  XOR U1459 ( .A(n1100), .B(n1099), .Z(n1096) );
  XOR U1460 ( .A(n1098), .B(n1203), .Z(n1099) );
  AND U1461 ( .A(g_input[8]), .B(e_input[18]), .Z(n1203) );
  XOR U1462 ( .A(n1106), .B(n1104), .Z(n1100) );
  XOR U1463 ( .A(n1102), .B(n1207), .Z(n1104) );
  AND U1464 ( .A(g_input[7]), .B(e_input[19]), .Z(n1207) );
  XOR U1465 ( .A(n1110), .B(n1109), .Z(n1106) );
  XOR U1466 ( .A(n1108), .B(n1211), .Z(n1109) );
  AND U1467 ( .A(g_input[6]), .B(e_input[20]), .Z(n1211) );
  XOR U1468 ( .A(n1114), .B(n1113), .Z(n1110) );
  XOR U1469 ( .A(n1112), .B(n1215), .Z(n1113) );
  AND U1470 ( .A(g_input[5]), .B(e_input[21]), .Z(n1215) );
  XOR U1471 ( .A(n1118), .B(n1117), .Z(n1114) );
  XOR U1472 ( .A(n1116), .B(n1219), .Z(n1117) );
  AND U1473 ( .A(g_input[4]), .B(e_input[22]), .Z(n1219) );
  XOR U1474 ( .A(n1122), .B(n1121), .Z(n1118) );
  XOR U1475 ( .A(n1120), .B(n1223), .Z(n1121) );
  AND U1476 ( .A(g_input[3]), .B(e_input[23]), .Z(n1223) );
  XNOR U1477 ( .A(n1126), .B(n1125), .Z(n1122) );
  XOR U1478 ( .A(n1124), .B(n1227), .Z(n1125) );
  AND U1479 ( .A(g_input[2]), .B(e_input[24]), .Z(n1227) );
  XOR U1480 ( .A(n1129), .B(n1130), .Z(n1126) );
  NANDN U1481 ( .B(n532), .A(e_input[26]), .Z(n1130) );
  XNOR U1482 ( .A(n1128), .B(n1231), .Z(n1129) );
  AND U1483 ( .A(g_input[1]), .B(e_input[25]), .Z(n1231) );
  XNOR U1484 ( .A(n1133), .B(o[25]), .Z(oi[25]) );
  XNOR U1485 ( .A(n1235), .B(n1132), .Z(n1133) );
  XNOR U1486 ( .A(n1136), .B(n1135), .Z(n1235) );
  NAND U1487 ( .A(g_input[25]), .B(e_input[0]), .Z(n1135) );
  XOR U1488 ( .A(n1140), .B(n1139), .Z(n1136) );
  XNOR U1489 ( .A(n1238), .B(n1138), .Z(n1139) );
  NANDN U1490 ( .B(n1239), .A(n1240), .Z(n1138) );
  NAND U1491 ( .A(e_input[1]), .B(g_input[24]), .Z(n1238) );
  XOR U1492 ( .A(n1144), .B(n1143), .Z(n1140) );
  XNOR U1493 ( .A(n1142), .B(n1241), .Z(n1143) );
  AND U1494 ( .A(e_input[2]), .B(g_input[23]), .Z(n1241) );
  XOR U1495 ( .A(n1148), .B(n1147), .Z(n1144) );
  XOR U1496 ( .A(n1146), .B(n1245), .Z(n1147) );
  AND U1497 ( .A(e_input[3]), .B(g_input[22]), .Z(n1245) );
  XOR U1498 ( .A(n1152), .B(n1151), .Z(n1148) );
  XOR U1499 ( .A(n1150), .B(n1249), .Z(n1151) );
  AND U1500 ( .A(e_input[4]), .B(g_input[21]), .Z(n1249) );
  XOR U1501 ( .A(n1156), .B(n1155), .Z(n1152) );
  XOR U1502 ( .A(n1154), .B(n1253), .Z(n1155) );
  AND U1503 ( .A(e_input[5]), .B(g_input[20]), .Z(n1253) );
  XOR U1504 ( .A(n1160), .B(n1159), .Z(n1156) );
  XOR U1505 ( .A(n1158), .B(n1257), .Z(n1159) );
  AND U1506 ( .A(e_input[6]), .B(g_input[19]), .Z(n1257) );
  XOR U1507 ( .A(n1164), .B(n1163), .Z(n1160) );
  XOR U1508 ( .A(n1162), .B(n1261), .Z(n1163) );
  AND U1509 ( .A(e_input[7]), .B(g_input[18]), .Z(n1261) );
  XOR U1510 ( .A(n1170), .B(n1168), .Z(n1164) );
  XOR U1511 ( .A(n1166), .B(n1265), .Z(n1168) );
  AND U1512 ( .A(e_input[8]), .B(g_input[17]), .Z(n1265) );
  XOR U1513 ( .A(n1174), .B(n1173), .Z(n1170) );
  XOR U1514 ( .A(n1172), .B(n1269), .Z(n1173) );
  AND U1515 ( .A(e_input[9]), .B(g_input[16]), .Z(n1269) );
  XOR U1516 ( .A(n1178), .B(n1177), .Z(n1174) );
  XOR U1517 ( .A(n1176), .B(n1273), .Z(n1177) );
  AND U1518 ( .A(g_input[15]), .B(e_input[10]), .Z(n1273) );
  XOR U1519 ( .A(n1182), .B(n1181), .Z(n1178) );
  XOR U1520 ( .A(n1180), .B(n1277), .Z(n1181) );
  AND U1521 ( .A(g_input[14]), .B(e_input[11]), .Z(n1277) );
  XOR U1522 ( .A(n1278), .B(n1279), .Z(n1180) );
  AND U1523 ( .A(n1280), .B(n1281), .Z(n1279) );
  XNOR U1524 ( .A(n1282), .B(n1278), .Z(n1281) );
  XOR U1525 ( .A(n1186), .B(n1185), .Z(n1182) );
  XOR U1526 ( .A(n1184), .B(n1283), .Z(n1185) );
  AND U1527 ( .A(g_input[13]), .B(e_input[12]), .Z(n1283) );
  XOR U1528 ( .A(n1190), .B(n1189), .Z(n1186) );
  XOR U1529 ( .A(n1188), .B(n1287), .Z(n1189) );
  AND U1530 ( .A(g_input[12]), .B(e_input[13]), .Z(n1287) );
  XOR U1531 ( .A(n1288), .B(n1289), .Z(n1188) );
  AND U1532 ( .A(n1290), .B(n1291), .Z(n1289) );
  XNOR U1533 ( .A(n1292), .B(n1288), .Z(n1291) );
  XOR U1534 ( .A(n1194), .B(n1193), .Z(n1190) );
  XOR U1535 ( .A(n1192), .B(n1293), .Z(n1193) );
  AND U1536 ( .A(g_input[11]), .B(e_input[14]), .Z(n1293) );
  XOR U1537 ( .A(n1198), .B(n1197), .Z(n1194) );
  XOR U1538 ( .A(n1196), .B(n1297), .Z(n1197) );
  AND U1539 ( .A(g_input[10]), .B(e_input[15]), .Z(n1297) );
  XOR U1540 ( .A(n1202), .B(n1201), .Z(n1198) );
  XOR U1541 ( .A(n1200), .B(n1301), .Z(n1201) );
  AND U1542 ( .A(g_input[9]), .B(e_input[16]), .Z(n1301) );
  XOR U1543 ( .A(n1206), .B(n1205), .Z(n1202) );
  XOR U1544 ( .A(n1204), .B(n1305), .Z(n1205) );
  AND U1545 ( .A(g_input[8]), .B(e_input[17]), .Z(n1305) );
  XOR U1546 ( .A(n1210), .B(n1209), .Z(n1206) );
  XOR U1547 ( .A(n1208), .B(n1309), .Z(n1209) );
  AND U1548 ( .A(g_input[7]), .B(e_input[18]), .Z(n1309) );
  XOR U1549 ( .A(n1214), .B(n1213), .Z(n1210) );
  XOR U1550 ( .A(n1212), .B(n1313), .Z(n1213) );
  AND U1551 ( .A(g_input[6]), .B(e_input[19]), .Z(n1313) );
  XOR U1552 ( .A(n1218), .B(n1217), .Z(n1214) );
  XOR U1553 ( .A(n1216), .B(n1317), .Z(n1217) );
  AND U1554 ( .A(g_input[5]), .B(e_input[20]), .Z(n1317) );
  XOR U1555 ( .A(n1222), .B(n1221), .Z(n1218) );
  XOR U1556 ( .A(n1220), .B(n1321), .Z(n1221) );
  AND U1557 ( .A(g_input[4]), .B(e_input[21]), .Z(n1321) );
  XOR U1558 ( .A(n1226), .B(n1225), .Z(n1222) );
  XOR U1559 ( .A(n1224), .B(n1325), .Z(n1225) );
  AND U1560 ( .A(g_input[3]), .B(e_input[22]), .Z(n1325) );
  XNOR U1561 ( .A(n1230), .B(n1229), .Z(n1226) );
  XOR U1562 ( .A(n1228), .B(n1329), .Z(n1229) );
  AND U1563 ( .A(g_input[2]), .B(e_input[23]), .Z(n1329) );
  XOR U1564 ( .A(n1233), .B(n1234), .Z(n1230) );
  NANDN U1565 ( .B(n532), .A(e_input[25]), .Z(n1234) );
  XNOR U1566 ( .A(n1232), .B(n1333), .Z(n1233) );
  AND U1567 ( .A(g_input[1]), .B(e_input[24]), .Z(n1333) );
  XNOR U1568 ( .A(n1237), .B(o[24]), .Z(oi[24]) );
  XNOR U1569 ( .A(n1337), .B(n1236), .Z(n1237) );
  XNOR U1570 ( .A(n1240), .B(n1239), .Z(n1337) );
  NAND U1571 ( .A(g_input[24]), .B(e_input[0]), .Z(n1239) );
  XOR U1572 ( .A(n1244), .B(n1243), .Z(n1240) );
  XNOR U1573 ( .A(n1340), .B(n1242), .Z(n1243) );
  NANDN U1574 ( .B(n1341), .A(n1342), .Z(n1242) );
  NAND U1575 ( .A(e_input[1]), .B(g_input[23]), .Z(n1340) );
  XOR U1576 ( .A(n1248), .B(n1247), .Z(n1244) );
  XNOR U1577 ( .A(n1246), .B(n1343), .Z(n1247) );
  AND U1578 ( .A(e_input[2]), .B(g_input[22]), .Z(n1343) );
  XOR U1579 ( .A(n1252), .B(n1251), .Z(n1248) );
  XOR U1580 ( .A(n1250), .B(n1347), .Z(n1251) );
  AND U1581 ( .A(e_input[3]), .B(g_input[21]), .Z(n1347) );
  XOR U1582 ( .A(n1256), .B(n1255), .Z(n1252) );
  XOR U1583 ( .A(n1254), .B(n1351), .Z(n1255) );
  AND U1584 ( .A(e_input[4]), .B(g_input[20]), .Z(n1351) );
  XOR U1585 ( .A(n1260), .B(n1259), .Z(n1256) );
  XOR U1586 ( .A(n1258), .B(n1355), .Z(n1259) );
  AND U1587 ( .A(e_input[5]), .B(g_input[19]), .Z(n1355) );
  XOR U1588 ( .A(n1264), .B(n1263), .Z(n1260) );
  XOR U1589 ( .A(n1262), .B(n1359), .Z(n1263) );
  AND U1590 ( .A(e_input[6]), .B(g_input[18]), .Z(n1359) );
  XOR U1591 ( .A(n1268), .B(n1267), .Z(n1264) );
  XOR U1592 ( .A(n1266), .B(n1363), .Z(n1267) );
  AND U1593 ( .A(e_input[7]), .B(g_input[17]), .Z(n1363) );
  XOR U1594 ( .A(n1272), .B(n1271), .Z(n1268) );
  XOR U1595 ( .A(n1270), .B(n1367), .Z(n1271) );
  AND U1596 ( .A(e_input[8]), .B(g_input[16]), .Z(n1367) );
  XOR U1597 ( .A(n1276), .B(n1275), .Z(n1272) );
  XOR U1598 ( .A(n1274), .B(n1371), .Z(n1275) );
  AND U1599 ( .A(e_input[9]), .B(g_input[15]), .Z(n1371) );
  XOR U1600 ( .A(n1282), .B(n1280), .Z(n1276) );
  XOR U1601 ( .A(n1278), .B(n1375), .Z(n1280) );
  AND U1602 ( .A(g_input[14]), .B(e_input[10]), .Z(n1375) );
  XOR U1603 ( .A(n1286), .B(n1285), .Z(n1282) );
  XOR U1604 ( .A(n1284), .B(n1379), .Z(n1285) );
  AND U1605 ( .A(g_input[13]), .B(e_input[11]), .Z(n1379) );
  XOR U1606 ( .A(n1292), .B(n1290), .Z(n1286) );
  XOR U1607 ( .A(n1288), .B(n1383), .Z(n1290) );
  AND U1608 ( .A(g_input[12]), .B(e_input[12]), .Z(n1383) );
  XOR U1609 ( .A(n1296), .B(n1295), .Z(n1292) );
  XOR U1610 ( .A(n1294), .B(n1387), .Z(n1295) );
  AND U1611 ( .A(g_input[11]), .B(e_input[13]), .Z(n1387) );
  XOR U1612 ( .A(n1300), .B(n1299), .Z(n1296) );
  XOR U1613 ( .A(n1298), .B(n1391), .Z(n1299) );
  AND U1614 ( .A(g_input[10]), .B(e_input[14]), .Z(n1391) );
  XOR U1615 ( .A(n1304), .B(n1303), .Z(n1300) );
  XOR U1616 ( .A(n1302), .B(n1395), .Z(n1303) );
  AND U1617 ( .A(g_input[9]), .B(e_input[15]), .Z(n1395) );
  XOR U1618 ( .A(n1396), .B(n1397), .Z(n1302) );
  AND U1619 ( .A(n1398), .B(n1399), .Z(n1397) );
  XNOR U1620 ( .A(n1400), .B(n1396), .Z(n1399) );
  XOR U1621 ( .A(n1308), .B(n1307), .Z(n1304) );
  XOR U1622 ( .A(n1306), .B(n1401), .Z(n1307) );
  AND U1623 ( .A(g_input[8]), .B(e_input[16]), .Z(n1401) );
  XOR U1624 ( .A(n1312), .B(n1311), .Z(n1308) );
  XOR U1625 ( .A(n1310), .B(n1405), .Z(n1311) );
  AND U1626 ( .A(g_input[7]), .B(e_input[17]), .Z(n1405) );
  XOR U1627 ( .A(n1316), .B(n1315), .Z(n1312) );
  XOR U1628 ( .A(n1314), .B(n1409), .Z(n1315) );
  AND U1629 ( .A(g_input[6]), .B(e_input[18]), .Z(n1409) );
  XOR U1630 ( .A(n1410), .B(n1411), .Z(n1314) );
  AND U1631 ( .A(n1412), .B(n1413), .Z(n1411) );
  XNOR U1632 ( .A(n1414), .B(n1410), .Z(n1413) );
  XOR U1633 ( .A(n1320), .B(n1319), .Z(n1316) );
  XOR U1634 ( .A(n1318), .B(n1415), .Z(n1319) );
  AND U1635 ( .A(g_input[5]), .B(e_input[19]), .Z(n1415) );
  XOR U1636 ( .A(n1416), .B(n1417), .Z(n1318) );
  AND U1637 ( .A(n1418), .B(n1419), .Z(n1417) );
  XNOR U1638 ( .A(n1420), .B(n1416), .Z(n1419) );
  XOR U1639 ( .A(n1324), .B(n1323), .Z(n1320) );
  XOR U1640 ( .A(n1322), .B(n1421), .Z(n1323) );
  AND U1641 ( .A(g_input[4]), .B(e_input[20]), .Z(n1421) );
  XOR U1642 ( .A(n1328), .B(n1327), .Z(n1324) );
  XOR U1643 ( .A(n1326), .B(n1425), .Z(n1327) );
  AND U1644 ( .A(g_input[3]), .B(e_input[21]), .Z(n1425) );
  XNOR U1645 ( .A(n1332), .B(n1331), .Z(n1328) );
  XOR U1646 ( .A(n1330), .B(n1429), .Z(n1331) );
  AND U1647 ( .A(g_input[2]), .B(e_input[22]), .Z(n1429) );
  XOR U1648 ( .A(n1335), .B(n1336), .Z(n1332) );
  NANDN U1649 ( .B(n532), .A(e_input[24]), .Z(n1336) );
  XNOR U1650 ( .A(n1334), .B(n1433), .Z(n1335) );
  AND U1651 ( .A(g_input[1]), .B(e_input[23]), .Z(n1433) );
  XNOR U1652 ( .A(n1339), .B(o[23]), .Z(oi[23]) );
  XNOR U1653 ( .A(n1437), .B(n1338), .Z(n1339) );
  XNOR U1654 ( .A(n1342), .B(n1341), .Z(n1437) );
  NAND U1655 ( .A(g_input[23]), .B(e_input[0]), .Z(n1341) );
  XOR U1656 ( .A(n1346), .B(n1345), .Z(n1342) );
  XNOR U1657 ( .A(n1440), .B(n1344), .Z(n1345) );
  NANDN U1658 ( .B(n1441), .A(n1442), .Z(n1344) );
  NAND U1659 ( .A(e_input[1]), .B(g_input[22]), .Z(n1440) );
  XOR U1660 ( .A(n1350), .B(n1349), .Z(n1346) );
  XNOR U1661 ( .A(n1348), .B(n1443), .Z(n1349) );
  AND U1662 ( .A(e_input[2]), .B(g_input[21]), .Z(n1443) );
  XOR U1663 ( .A(n1354), .B(n1353), .Z(n1350) );
  XOR U1664 ( .A(n1352), .B(n1447), .Z(n1353) );
  AND U1665 ( .A(e_input[3]), .B(g_input[20]), .Z(n1447) );
  XOR U1666 ( .A(n1358), .B(n1357), .Z(n1354) );
  XOR U1667 ( .A(n1356), .B(n1451), .Z(n1357) );
  AND U1668 ( .A(e_input[4]), .B(g_input[19]), .Z(n1451) );
  XOR U1669 ( .A(n1362), .B(n1361), .Z(n1358) );
  XOR U1670 ( .A(n1360), .B(n1455), .Z(n1361) );
  AND U1671 ( .A(e_input[5]), .B(g_input[18]), .Z(n1455) );
  XOR U1672 ( .A(n1366), .B(n1365), .Z(n1362) );
  XOR U1673 ( .A(n1364), .B(n1459), .Z(n1365) );
  AND U1674 ( .A(e_input[6]), .B(g_input[17]), .Z(n1459) );
  XOR U1675 ( .A(n1370), .B(n1369), .Z(n1366) );
  XOR U1676 ( .A(n1368), .B(n1463), .Z(n1369) );
  AND U1677 ( .A(e_input[7]), .B(g_input[16]), .Z(n1463) );
  XOR U1678 ( .A(n1374), .B(n1373), .Z(n1370) );
  XOR U1679 ( .A(n1372), .B(n1467), .Z(n1373) );
  AND U1680 ( .A(e_input[8]), .B(g_input[15]), .Z(n1467) );
  XOR U1681 ( .A(n1378), .B(n1377), .Z(n1374) );
  XOR U1682 ( .A(n1376), .B(n1471), .Z(n1377) );
  AND U1683 ( .A(e_input[9]), .B(g_input[14]), .Z(n1471) );
  XOR U1684 ( .A(n1382), .B(n1381), .Z(n1378) );
  XOR U1685 ( .A(n1380), .B(n1475), .Z(n1381) );
  AND U1686 ( .A(g_input[13]), .B(e_input[10]), .Z(n1475) );
  XOR U1687 ( .A(n1386), .B(n1385), .Z(n1382) );
  XOR U1688 ( .A(n1384), .B(n1479), .Z(n1385) );
  AND U1689 ( .A(g_input[12]), .B(e_input[11]), .Z(n1479) );
  XOR U1690 ( .A(n1390), .B(n1389), .Z(n1386) );
  XOR U1691 ( .A(n1388), .B(n1483), .Z(n1389) );
  AND U1692 ( .A(g_input[11]), .B(e_input[12]), .Z(n1483) );
  XOR U1693 ( .A(n1394), .B(n1393), .Z(n1390) );
  XOR U1694 ( .A(n1392), .B(n1487), .Z(n1393) );
  AND U1695 ( .A(g_input[10]), .B(e_input[13]), .Z(n1487) );
  XOR U1696 ( .A(n1400), .B(n1398), .Z(n1394) );
  XOR U1697 ( .A(n1396), .B(n1491), .Z(n1398) );
  AND U1698 ( .A(g_input[9]), .B(e_input[14]), .Z(n1491) );
  XOR U1699 ( .A(n1404), .B(n1403), .Z(n1400) );
  XOR U1700 ( .A(n1402), .B(n1495), .Z(n1403) );
  AND U1701 ( .A(g_input[8]), .B(e_input[15]), .Z(n1495) );
  XOR U1702 ( .A(n1408), .B(n1407), .Z(n1404) );
  XOR U1703 ( .A(n1406), .B(n1499), .Z(n1407) );
  AND U1704 ( .A(g_input[7]), .B(e_input[16]), .Z(n1499) );
  XOR U1705 ( .A(n1414), .B(n1412), .Z(n1408) );
  XOR U1706 ( .A(n1410), .B(n1503), .Z(n1412) );
  AND U1707 ( .A(g_input[6]), .B(e_input[17]), .Z(n1503) );
  XOR U1708 ( .A(n1420), .B(n1418), .Z(n1414) );
  XOR U1709 ( .A(n1416), .B(n1507), .Z(n1418) );
  AND U1710 ( .A(g_input[5]), .B(e_input[18]), .Z(n1507) );
  XOR U1711 ( .A(n1424), .B(n1423), .Z(n1420) );
  XOR U1712 ( .A(n1422), .B(n1511), .Z(n1423) );
  AND U1713 ( .A(g_input[4]), .B(e_input[19]), .Z(n1511) );
  XOR U1714 ( .A(n1428), .B(n1427), .Z(n1424) );
  XOR U1715 ( .A(n1426), .B(n1515), .Z(n1427) );
  AND U1716 ( .A(g_input[3]), .B(e_input[20]), .Z(n1515) );
  XOR U1717 ( .A(n1516), .B(n1517), .Z(n1426) );
  AND U1718 ( .A(n1518), .B(n1519), .Z(n1517) );
  XNOR U1719 ( .A(n1520), .B(n1516), .Z(n1519) );
  XNOR U1720 ( .A(n1432), .B(n1431), .Z(n1428) );
  XOR U1721 ( .A(n1430), .B(n1521), .Z(n1431) );
  AND U1722 ( .A(g_input[2]), .B(e_input[21]), .Z(n1521) );
  XOR U1723 ( .A(n1435), .B(n1436), .Z(n1432) );
  NANDN U1724 ( .B(n532), .A(e_input[23]), .Z(n1436) );
  XNOR U1725 ( .A(n1434), .B(n1525), .Z(n1435) );
  AND U1726 ( .A(g_input[1]), .B(e_input[22]), .Z(n1525) );
  XNOR U1727 ( .A(n1439), .B(o[22]), .Z(oi[22]) );
  XNOR U1728 ( .A(n1529), .B(n1438), .Z(n1439) );
  XNOR U1729 ( .A(n1442), .B(n1441), .Z(n1529) );
  NAND U1730 ( .A(g_input[22]), .B(e_input[0]), .Z(n1441) );
  XOR U1731 ( .A(n1446), .B(n1445), .Z(n1442) );
  XNOR U1732 ( .A(n1532), .B(n1444), .Z(n1445) );
  NANDN U1733 ( .B(n1533), .A(n1534), .Z(n1444) );
  NAND U1734 ( .A(e_input[1]), .B(g_input[21]), .Z(n1532) );
  XOR U1735 ( .A(n1450), .B(n1449), .Z(n1446) );
  XNOR U1736 ( .A(n1448), .B(n1535), .Z(n1449) );
  AND U1737 ( .A(e_input[2]), .B(g_input[20]), .Z(n1535) );
  XOR U1738 ( .A(n1454), .B(n1453), .Z(n1450) );
  XOR U1739 ( .A(n1452), .B(n1539), .Z(n1453) );
  AND U1740 ( .A(e_input[3]), .B(g_input[19]), .Z(n1539) );
  XOR U1741 ( .A(n1458), .B(n1457), .Z(n1454) );
  XOR U1742 ( .A(n1456), .B(n1543), .Z(n1457) );
  AND U1743 ( .A(e_input[4]), .B(g_input[18]), .Z(n1543) );
  XOR U1744 ( .A(n1462), .B(n1461), .Z(n1458) );
  XOR U1745 ( .A(n1460), .B(n1547), .Z(n1461) );
  AND U1746 ( .A(e_input[5]), .B(g_input[17]), .Z(n1547) );
  XOR U1747 ( .A(n1466), .B(n1465), .Z(n1462) );
  XOR U1748 ( .A(n1464), .B(n1551), .Z(n1465) );
  AND U1749 ( .A(e_input[6]), .B(g_input[16]), .Z(n1551) );
  XOR U1750 ( .A(n1470), .B(n1469), .Z(n1466) );
  XOR U1751 ( .A(n1468), .B(n1555), .Z(n1469) );
  AND U1752 ( .A(e_input[7]), .B(g_input[15]), .Z(n1555) );
  XOR U1753 ( .A(n1474), .B(n1473), .Z(n1470) );
  XOR U1754 ( .A(n1472), .B(n1559), .Z(n1473) );
  AND U1755 ( .A(e_input[8]), .B(g_input[14]), .Z(n1559) );
  XOR U1756 ( .A(n1478), .B(n1477), .Z(n1474) );
  XOR U1757 ( .A(n1476), .B(n1563), .Z(n1477) );
  AND U1758 ( .A(e_input[9]), .B(g_input[13]), .Z(n1563) );
  XOR U1759 ( .A(n1482), .B(n1481), .Z(n1478) );
  XOR U1760 ( .A(n1480), .B(n1567), .Z(n1481) );
  AND U1761 ( .A(g_input[12]), .B(e_input[10]), .Z(n1567) );
  XOR U1762 ( .A(n1486), .B(n1485), .Z(n1482) );
  XOR U1763 ( .A(n1484), .B(n1571), .Z(n1485) );
  AND U1764 ( .A(g_input[11]), .B(e_input[11]), .Z(n1571) );
  XOR U1765 ( .A(n1490), .B(n1489), .Z(n1486) );
  XOR U1766 ( .A(n1488), .B(n1575), .Z(n1489) );
  AND U1767 ( .A(g_input[10]), .B(e_input[12]), .Z(n1575) );
  XOR U1768 ( .A(n1494), .B(n1493), .Z(n1490) );
  XOR U1769 ( .A(n1492), .B(n1579), .Z(n1493) );
  AND U1770 ( .A(g_input[9]), .B(e_input[13]), .Z(n1579) );
  XOR U1771 ( .A(n1498), .B(n1497), .Z(n1494) );
  XOR U1772 ( .A(n1496), .B(n1583), .Z(n1497) );
  AND U1773 ( .A(g_input[8]), .B(e_input[14]), .Z(n1583) );
  XOR U1774 ( .A(n1502), .B(n1501), .Z(n1498) );
  XOR U1775 ( .A(n1500), .B(n1587), .Z(n1501) );
  AND U1776 ( .A(g_input[7]), .B(e_input[15]), .Z(n1587) );
  XOR U1777 ( .A(n1506), .B(n1505), .Z(n1502) );
  XOR U1778 ( .A(n1504), .B(n1591), .Z(n1505) );
  AND U1779 ( .A(g_input[6]), .B(e_input[16]), .Z(n1591) );
  XOR U1780 ( .A(n1510), .B(n1509), .Z(n1506) );
  XOR U1781 ( .A(n1508), .B(n1595), .Z(n1509) );
  AND U1782 ( .A(g_input[5]), .B(e_input[17]), .Z(n1595) );
  XOR U1783 ( .A(n1514), .B(n1513), .Z(n1510) );
  XOR U1784 ( .A(n1512), .B(n1599), .Z(n1513) );
  AND U1785 ( .A(g_input[4]), .B(e_input[18]), .Z(n1599) );
  XOR U1786 ( .A(n1520), .B(n1518), .Z(n1514) );
  XOR U1787 ( .A(n1516), .B(n1603), .Z(n1518) );
  AND U1788 ( .A(g_input[3]), .B(e_input[19]), .Z(n1603) );
  XNOR U1789 ( .A(n1524), .B(n1523), .Z(n1520) );
  XOR U1790 ( .A(n1522), .B(n1607), .Z(n1523) );
  AND U1791 ( .A(g_input[2]), .B(e_input[20]), .Z(n1607) );
  XOR U1792 ( .A(n1527), .B(n1528), .Z(n1524) );
  NANDN U1793 ( .B(n532), .A(e_input[22]), .Z(n1528) );
  XNOR U1794 ( .A(n1526), .B(n1611), .Z(n1527) );
  AND U1795 ( .A(g_input[1]), .B(e_input[21]), .Z(n1611) );
  XNOR U1796 ( .A(n1531), .B(o[21]), .Z(oi[21]) );
  XNOR U1797 ( .A(n1615), .B(n1530), .Z(n1531) );
  XNOR U1798 ( .A(n1534), .B(n1533), .Z(n1615) );
  NAND U1799 ( .A(g_input[21]), .B(e_input[0]), .Z(n1533) );
  XOR U1800 ( .A(n1538), .B(n1537), .Z(n1534) );
  XNOR U1801 ( .A(n1618), .B(n1536), .Z(n1537) );
  NANDN U1802 ( .B(n1619), .A(n1620), .Z(n1536) );
  NAND U1803 ( .A(e_input[1]), .B(g_input[20]), .Z(n1618) );
  XOR U1804 ( .A(n1542), .B(n1541), .Z(n1538) );
  XNOR U1805 ( .A(n1540), .B(n1621), .Z(n1541) );
  AND U1806 ( .A(e_input[2]), .B(g_input[19]), .Z(n1621) );
  XOR U1807 ( .A(n1546), .B(n1545), .Z(n1542) );
  XOR U1808 ( .A(n1544), .B(n1625), .Z(n1545) );
  AND U1809 ( .A(e_input[3]), .B(g_input[18]), .Z(n1625) );
  XOR U1810 ( .A(n1550), .B(n1549), .Z(n1546) );
  XOR U1811 ( .A(n1548), .B(n1629), .Z(n1549) );
  AND U1812 ( .A(e_input[4]), .B(g_input[17]), .Z(n1629) );
  XOR U1813 ( .A(n1554), .B(n1553), .Z(n1550) );
  XOR U1814 ( .A(n1552), .B(n1633), .Z(n1553) );
  AND U1815 ( .A(e_input[5]), .B(g_input[16]), .Z(n1633) );
  XOR U1816 ( .A(n1558), .B(n1557), .Z(n1554) );
  XOR U1817 ( .A(n1556), .B(n1637), .Z(n1557) );
  AND U1818 ( .A(e_input[6]), .B(g_input[15]), .Z(n1637) );
  XOR U1819 ( .A(n1562), .B(n1561), .Z(n1558) );
  XOR U1820 ( .A(n1560), .B(n1641), .Z(n1561) );
  AND U1821 ( .A(e_input[7]), .B(g_input[14]), .Z(n1641) );
  XOR U1822 ( .A(n1566), .B(n1565), .Z(n1562) );
  XOR U1823 ( .A(n1564), .B(n1645), .Z(n1565) );
  AND U1824 ( .A(e_input[8]), .B(g_input[13]), .Z(n1645) );
  XOR U1825 ( .A(n1570), .B(n1569), .Z(n1566) );
  XOR U1826 ( .A(n1568), .B(n1649), .Z(n1569) );
  AND U1827 ( .A(e_input[9]), .B(g_input[12]), .Z(n1649) );
  XOR U1828 ( .A(n1574), .B(n1573), .Z(n1570) );
  XOR U1829 ( .A(n1572), .B(n1653), .Z(n1573) );
  AND U1830 ( .A(g_input[11]), .B(e_input[10]), .Z(n1653) );
  XOR U1831 ( .A(n1578), .B(n1577), .Z(n1574) );
  XOR U1832 ( .A(n1576), .B(n1657), .Z(n1577) );
  AND U1833 ( .A(g_input[10]), .B(e_input[11]), .Z(n1657) );
  XOR U1834 ( .A(n1582), .B(n1581), .Z(n1578) );
  XOR U1835 ( .A(n1580), .B(n1661), .Z(n1581) );
  AND U1836 ( .A(g_input[9]), .B(e_input[12]), .Z(n1661) );
  XOR U1837 ( .A(n1586), .B(n1585), .Z(n1582) );
  XOR U1838 ( .A(n1584), .B(n1665), .Z(n1585) );
  AND U1839 ( .A(g_input[8]), .B(e_input[13]), .Z(n1665) );
  XOR U1840 ( .A(n1590), .B(n1589), .Z(n1586) );
  XOR U1841 ( .A(n1588), .B(n1669), .Z(n1589) );
  AND U1842 ( .A(g_input[7]), .B(e_input[14]), .Z(n1669) );
  XOR U1843 ( .A(n1594), .B(n1593), .Z(n1590) );
  XOR U1844 ( .A(n1592), .B(n1673), .Z(n1593) );
  AND U1845 ( .A(g_input[6]), .B(e_input[15]), .Z(n1673) );
  XOR U1846 ( .A(n1598), .B(n1597), .Z(n1594) );
  XOR U1847 ( .A(n1596), .B(n1677), .Z(n1597) );
  AND U1848 ( .A(g_input[5]), .B(e_input[16]), .Z(n1677) );
  XOR U1849 ( .A(n1602), .B(n1601), .Z(n1598) );
  XOR U1850 ( .A(n1600), .B(n1681), .Z(n1601) );
  AND U1851 ( .A(g_input[4]), .B(e_input[17]), .Z(n1681) );
  XOR U1852 ( .A(n1606), .B(n1605), .Z(n1602) );
  XOR U1853 ( .A(n1604), .B(n1685), .Z(n1605) );
  AND U1854 ( .A(g_input[3]), .B(e_input[18]), .Z(n1685) );
  XNOR U1855 ( .A(n1610), .B(n1609), .Z(n1606) );
  XOR U1856 ( .A(n1608), .B(n1689), .Z(n1609) );
  AND U1857 ( .A(g_input[2]), .B(e_input[19]), .Z(n1689) );
  XOR U1858 ( .A(n1613), .B(n1614), .Z(n1610) );
  NANDN U1859 ( .B(n532), .A(e_input[21]), .Z(n1614) );
  XNOR U1860 ( .A(n1612), .B(n1693), .Z(n1613) );
  AND U1861 ( .A(g_input[1]), .B(e_input[20]), .Z(n1693) );
  XNOR U1862 ( .A(n1617), .B(o[20]), .Z(oi[20]) );
  XNOR U1863 ( .A(n1697), .B(n1616), .Z(n1617) );
  XNOR U1864 ( .A(n1620), .B(n1619), .Z(n1697) );
  NAND U1865 ( .A(g_input[20]), .B(e_input[0]), .Z(n1619) );
  XOR U1866 ( .A(n1624), .B(n1623), .Z(n1620) );
  XNOR U1867 ( .A(n1700), .B(n1622), .Z(n1623) );
  NANDN U1868 ( .B(n1701), .A(n1702), .Z(n1622) );
  NAND U1869 ( .A(e_input[1]), .B(g_input[19]), .Z(n1700) );
  XOR U1870 ( .A(n1628), .B(n1627), .Z(n1624) );
  XNOR U1871 ( .A(n1626), .B(n1703), .Z(n1627) );
  AND U1872 ( .A(e_input[2]), .B(g_input[18]), .Z(n1703) );
  XOR U1873 ( .A(n1632), .B(n1631), .Z(n1628) );
  XOR U1874 ( .A(n1630), .B(n1707), .Z(n1631) );
  AND U1875 ( .A(e_input[3]), .B(g_input[17]), .Z(n1707) );
  XOR U1876 ( .A(n1636), .B(n1635), .Z(n1632) );
  XOR U1877 ( .A(n1634), .B(n1711), .Z(n1635) );
  AND U1878 ( .A(e_input[4]), .B(g_input[16]), .Z(n1711) );
  XOR U1879 ( .A(n1640), .B(n1639), .Z(n1636) );
  XOR U1880 ( .A(n1638), .B(n1715), .Z(n1639) );
  AND U1881 ( .A(e_input[5]), .B(g_input[15]), .Z(n1715) );
  XOR U1882 ( .A(n1644), .B(n1643), .Z(n1640) );
  XOR U1883 ( .A(n1642), .B(n1719), .Z(n1643) );
  AND U1884 ( .A(e_input[6]), .B(g_input[14]), .Z(n1719) );
  XOR U1885 ( .A(n1648), .B(n1647), .Z(n1644) );
  XOR U1886 ( .A(n1646), .B(n1723), .Z(n1647) );
  AND U1887 ( .A(e_input[7]), .B(g_input[13]), .Z(n1723) );
  XOR U1888 ( .A(n1652), .B(n1651), .Z(n1648) );
  XOR U1889 ( .A(n1650), .B(n1727), .Z(n1651) );
  AND U1890 ( .A(e_input[8]), .B(g_input[12]), .Z(n1727) );
  XOR U1891 ( .A(n1656), .B(n1655), .Z(n1652) );
  XOR U1892 ( .A(n1654), .B(n1731), .Z(n1655) );
  AND U1893 ( .A(e_input[9]), .B(g_input[11]), .Z(n1731) );
  XOR U1894 ( .A(n1660), .B(n1659), .Z(n1656) );
  XOR U1895 ( .A(n1658), .B(n1735), .Z(n1659) );
  AND U1896 ( .A(g_input[10]), .B(e_input[10]), .Z(n1735) );
  XOR U1897 ( .A(n1664), .B(n1663), .Z(n1660) );
  XOR U1898 ( .A(n1662), .B(n1739), .Z(n1663) );
  AND U1899 ( .A(g_input[9]), .B(e_input[11]), .Z(n1739) );
  XOR U1900 ( .A(n1668), .B(n1667), .Z(n1664) );
  XOR U1901 ( .A(n1666), .B(n1743), .Z(n1667) );
  AND U1902 ( .A(g_input[8]), .B(e_input[12]), .Z(n1743) );
  XOR U1903 ( .A(n1672), .B(n1671), .Z(n1668) );
  XOR U1904 ( .A(n1670), .B(n1747), .Z(n1671) );
  AND U1905 ( .A(g_input[7]), .B(e_input[13]), .Z(n1747) );
  XOR U1906 ( .A(n1676), .B(n1675), .Z(n1672) );
  XOR U1907 ( .A(n1674), .B(n1751), .Z(n1675) );
  AND U1908 ( .A(g_input[6]), .B(e_input[14]), .Z(n1751) );
  XOR U1909 ( .A(n1680), .B(n1679), .Z(n1676) );
  XOR U1910 ( .A(n1678), .B(n1755), .Z(n1679) );
  AND U1911 ( .A(g_input[5]), .B(e_input[15]), .Z(n1755) );
  XOR U1912 ( .A(n1684), .B(n1683), .Z(n1680) );
  XOR U1913 ( .A(n1682), .B(n1759), .Z(n1683) );
  AND U1914 ( .A(g_input[4]), .B(e_input[16]), .Z(n1759) );
  XOR U1915 ( .A(n1688), .B(n1687), .Z(n1684) );
  XOR U1916 ( .A(n1686), .B(n1763), .Z(n1687) );
  AND U1917 ( .A(g_input[3]), .B(e_input[17]), .Z(n1763) );
  XNOR U1918 ( .A(n1692), .B(n1691), .Z(n1688) );
  XOR U1919 ( .A(n1690), .B(n1767), .Z(n1691) );
  AND U1920 ( .A(g_input[2]), .B(e_input[18]), .Z(n1767) );
  XOR U1921 ( .A(n1695), .B(n1696), .Z(n1692) );
  NANDN U1922 ( .B(n532), .A(e_input[20]), .Z(n1696) );
  XNOR U1923 ( .A(n1694), .B(n1771), .Z(n1695) );
  AND U1924 ( .A(g_input[1]), .B(e_input[19]), .Z(n1771) );
  XNOR U1925 ( .A(o[1]), .B(n1775), .Z(oi[1]) );
  XNOR U1926 ( .A(n1699), .B(o[19]), .Z(oi[19]) );
  XNOR U1927 ( .A(n1776), .B(n1698), .Z(n1699) );
  XNOR U1928 ( .A(n1702), .B(n1701), .Z(n1776) );
  NAND U1929 ( .A(g_input[19]), .B(e_input[0]), .Z(n1701) );
  XOR U1930 ( .A(n1706), .B(n1705), .Z(n1702) );
  XNOR U1931 ( .A(n1779), .B(n1704), .Z(n1705) );
  NANDN U1932 ( .B(n1780), .A(n1781), .Z(n1704) );
  NAND U1933 ( .A(e_input[1]), .B(g_input[18]), .Z(n1779) );
  XOR U1934 ( .A(n1710), .B(n1709), .Z(n1706) );
  XNOR U1935 ( .A(n1708), .B(n1782), .Z(n1709) );
  AND U1936 ( .A(e_input[2]), .B(g_input[17]), .Z(n1782) );
  XOR U1937 ( .A(n1714), .B(n1713), .Z(n1710) );
  XOR U1938 ( .A(n1712), .B(n1786), .Z(n1713) );
  AND U1939 ( .A(e_input[3]), .B(g_input[16]), .Z(n1786) );
  XOR U1940 ( .A(n1718), .B(n1717), .Z(n1714) );
  XOR U1941 ( .A(n1716), .B(n1790), .Z(n1717) );
  AND U1942 ( .A(e_input[4]), .B(g_input[15]), .Z(n1790) );
  XOR U1943 ( .A(n1722), .B(n1721), .Z(n1718) );
  XOR U1944 ( .A(n1720), .B(n1794), .Z(n1721) );
  AND U1945 ( .A(e_input[5]), .B(g_input[14]), .Z(n1794) );
  XOR U1946 ( .A(n1726), .B(n1725), .Z(n1722) );
  XOR U1947 ( .A(n1724), .B(n1798), .Z(n1725) );
  AND U1948 ( .A(e_input[6]), .B(g_input[13]), .Z(n1798) );
  XOR U1949 ( .A(n1730), .B(n1729), .Z(n1726) );
  XOR U1950 ( .A(n1728), .B(n1802), .Z(n1729) );
  AND U1951 ( .A(e_input[7]), .B(g_input[12]), .Z(n1802) );
  XOR U1952 ( .A(n1734), .B(n1733), .Z(n1730) );
  XOR U1953 ( .A(n1732), .B(n1806), .Z(n1733) );
  AND U1954 ( .A(e_input[8]), .B(g_input[11]), .Z(n1806) );
  XOR U1955 ( .A(n1738), .B(n1737), .Z(n1734) );
  XOR U1956 ( .A(n1736), .B(n1810), .Z(n1737) );
  AND U1957 ( .A(e_input[9]), .B(g_input[10]), .Z(n1810) );
  XOR U1958 ( .A(n1742), .B(n1741), .Z(n1738) );
  XOR U1959 ( .A(n1740), .B(n1814), .Z(n1741) );
  AND U1960 ( .A(g_input[9]), .B(e_input[10]), .Z(n1814) );
  XOR U1961 ( .A(n1746), .B(n1745), .Z(n1742) );
  XOR U1962 ( .A(n1744), .B(n1818), .Z(n1745) );
  AND U1963 ( .A(g_input[8]), .B(e_input[11]), .Z(n1818) );
  XOR U1964 ( .A(n1750), .B(n1749), .Z(n1746) );
  XOR U1965 ( .A(n1748), .B(n1822), .Z(n1749) );
  AND U1966 ( .A(g_input[7]), .B(e_input[12]), .Z(n1822) );
  XOR U1967 ( .A(n1754), .B(n1753), .Z(n1750) );
  XOR U1968 ( .A(n1752), .B(n1826), .Z(n1753) );
  AND U1969 ( .A(g_input[6]), .B(e_input[13]), .Z(n1826) );
  XOR U1970 ( .A(n1758), .B(n1757), .Z(n1754) );
  XOR U1971 ( .A(n1756), .B(n1830), .Z(n1757) );
  AND U1972 ( .A(g_input[5]), .B(e_input[14]), .Z(n1830) );
  XOR U1973 ( .A(n1762), .B(n1761), .Z(n1758) );
  XOR U1974 ( .A(n1760), .B(n1834), .Z(n1761) );
  AND U1975 ( .A(g_input[4]), .B(e_input[15]), .Z(n1834) );
  XOR U1976 ( .A(n1766), .B(n1765), .Z(n1762) );
  XOR U1977 ( .A(n1764), .B(n1838), .Z(n1765) );
  AND U1978 ( .A(g_input[3]), .B(e_input[16]), .Z(n1838) );
  XNOR U1979 ( .A(n1770), .B(n1769), .Z(n1766) );
  XOR U1980 ( .A(n1768), .B(n1842), .Z(n1769) );
  AND U1981 ( .A(g_input[2]), .B(e_input[17]), .Z(n1842) );
  XOR U1982 ( .A(n1773), .B(n1774), .Z(n1770) );
  NANDN U1983 ( .B(n532), .A(e_input[19]), .Z(n1774) );
  XNOR U1984 ( .A(n1772), .B(n1846), .Z(n1773) );
  AND U1985 ( .A(g_input[1]), .B(e_input[18]), .Z(n1846) );
  XNOR U1986 ( .A(n1778), .B(o[18]), .Z(oi[18]) );
  XNOR U1987 ( .A(n1850), .B(n1777), .Z(n1778) );
  XNOR U1988 ( .A(n1781), .B(n1780), .Z(n1850) );
  NAND U1989 ( .A(g_input[18]), .B(e_input[0]), .Z(n1780) );
  XOR U1990 ( .A(n1785), .B(n1784), .Z(n1781) );
  XNOR U1991 ( .A(n1853), .B(n1783), .Z(n1784) );
  NANDN U1992 ( .B(n1854), .A(n1855), .Z(n1783) );
  NAND U1993 ( .A(e_input[1]), .B(g_input[17]), .Z(n1853) );
  XOR U1994 ( .A(n1789), .B(n1788), .Z(n1785) );
  XNOR U1995 ( .A(n1787), .B(n1856), .Z(n1788) );
  AND U1996 ( .A(e_input[2]), .B(g_input[16]), .Z(n1856) );
  XOR U1997 ( .A(n1793), .B(n1792), .Z(n1789) );
  XOR U1998 ( .A(n1791), .B(n1860), .Z(n1792) );
  AND U1999 ( .A(e_input[3]), .B(g_input[15]), .Z(n1860) );
  XOR U2000 ( .A(n1797), .B(n1796), .Z(n1793) );
  XOR U2001 ( .A(n1795), .B(n1864), .Z(n1796) );
  AND U2002 ( .A(e_input[4]), .B(g_input[14]), .Z(n1864) );
  XOR U2003 ( .A(n1801), .B(n1800), .Z(n1797) );
  XOR U2004 ( .A(n1799), .B(n1868), .Z(n1800) );
  AND U2005 ( .A(e_input[5]), .B(g_input[13]), .Z(n1868) );
  XOR U2006 ( .A(n1805), .B(n1804), .Z(n1801) );
  XOR U2007 ( .A(n1803), .B(n1872), .Z(n1804) );
  AND U2008 ( .A(e_input[6]), .B(g_input[12]), .Z(n1872) );
  XOR U2009 ( .A(n1809), .B(n1808), .Z(n1805) );
  XOR U2010 ( .A(n1807), .B(n1876), .Z(n1808) );
  AND U2011 ( .A(e_input[7]), .B(g_input[11]), .Z(n1876) );
  XOR U2012 ( .A(n1813), .B(n1812), .Z(n1809) );
  XOR U2013 ( .A(n1811), .B(n1880), .Z(n1812) );
  AND U2014 ( .A(e_input[8]), .B(g_input[10]), .Z(n1880) );
  XOR U2015 ( .A(n1817), .B(n1816), .Z(n1813) );
  XOR U2016 ( .A(n1815), .B(n1884), .Z(n1816) );
  AND U2017 ( .A(g_input[9]), .B(e_input[9]), .Z(n1884) );
  XOR U2018 ( .A(n1821), .B(n1820), .Z(n1817) );
  XOR U2019 ( .A(n1819), .B(n1888), .Z(n1820) );
  AND U2020 ( .A(g_input[8]), .B(e_input[10]), .Z(n1888) );
  XOR U2021 ( .A(n1825), .B(n1824), .Z(n1821) );
  XOR U2022 ( .A(n1823), .B(n1892), .Z(n1824) );
  AND U2023 ( .A(g_input[7]), .B(e_input[11]), .Z(n1892) );
  XOR U2024 ( .A(n1829), .B(n1828), .Z(n1825) );
  XOR U2025 ( .A(n1827), .B(n1896), .Z(n1828) );
  AND U2026 ( .A(g_input[6]), .B(e_input[12]), .Z(n1896) );
  XOR U2027 ( .A(n1833), .B(n1832), .Z(n1829) );
  XOR U2028 ( .A(n1831), .B(n1900), .Z(n1832) );
  AND U2029 ( .A(g_input[5]), .B(e_input[13]), .Z(n1900) );
  XOR U2030 ( .A(n1837), .B(n1836), .Z(n1833) );
  XOR U2031 ( .A(n1835), .B(n1904), .Z(n1836) );
  AND U2032 ( .A(g_input[4]), .B(e_input[14]), .Z(n1904) );
  XOR U2033 ( .A(n1841), .B(n1840), .Z(n1837) );
  XOR U2034 ( .A(n1839), .B(n1908), .Z(n1840) );
  AND U2035 ( .A(g_input[3]), .B(e_input[15]), .Z(n1908) );
  XNOR U2036 ( .A(n1845), .B(n1844), .Z(n1841) );
  XOR U2037 ( .A(n1843), .B(n1912), .Z(n1844) );
  AND U2038 ( .A(g_input[2]), .B(e_input[16]), .Z(n1912) );
  XOR U2039 ( .A(n1848), .B(n1849), .Z(n1845) );
  NANDN U2040 ( .B(n532), .A(e_input[18]), .Z(n1849) );
  XNOR U2041 ( .A(n1847), .B(n1916), .Z(n1848) );
  AND U2042 ( .A(g_input[1]), .B(e_input[17]), .Z(n1916) );
  XNOR U2043 ( .A(n1852), .B(o[17]), .Z(oi[17]) );
  XNOR U2044 ( .A(n1920), .B(n1851), .Z(n1852) );
  XNOR U2045 ( .A(n1855), .B(n1854), .Z(n1920) );
  NAND U2046 ( .A(g_input[17]), .B(e_input[0]), .Z(n1854) );
  XOR U2047 ( .A(n1859), .B(n1858), .Z(n1855) );
  XNOR U2048 ( .A(n1923), .B(n1857), .Z(n1858) );
  NANDN U2049 ( .B(n1924), .A(n1925), .Z(n1857) );
  NAND U2050 ( .A(e_input[1]), .B(g_input[16]), .Z(n1923) );
  XOR U2051 ( .A(n1863), .B(n1862), .Z(n1859) );
  XNOR U2052 ( .A(n1861), .B(n1926), .Z(n1862) );
  AND U2053 ( .A(e_input[2]), .B(g_input[15]), .Z(n1926) );
  XOR U2054 ( .A(n1867), .B(n1866), .Z(n1863) );
  XOR U2055 ( .A(n1865), .B(n1930), .Z(n1866) );
  AND U2056 ( .A(e_input[3]), .B(g_input[14]), .Z(n1930) );
  XOR U2057 ( .A(n1871), .B(n1870), .Z(n1867) );
  XOR U2058 ( .A(n1869), .B(n1934), .Z(n1870) );
  AND U2059 ( .A(e_input[4]), .B(g_input[13]), .Z(n1934) );
  XOR U2060 ( .A(n1875), .B(n1874), .Z(n1871) );
  XOR U2061 ( .A(n1873), .B(n1938), .Z(n1874) );
  AND U2062 ( .A(e_input[5]), .B(g_input[12]), .Z(n1938) );
  XOR U2063 ( .A(n1879), .B(n1878), .Z(n1875) );
  XOR U2064 ( .A(n1877), .B(n1942), .Z(n1878) );
  AND U2065 ( .A(e_input[6]), .B(g_input[11]), .Z(n1942) );
  XOR U2066 ( .A(n1883), .B(n1882), .Z(n1879) );
  XOR U2067 ( .A(n1881), .B(n1946), .Z(n1882) );
  AND U2068 ( .A(e_input[7]), .B(g_input[10]), .Z(n1946) );
  XOR U2069 ( .A(n1887), .B(n1886), .Z(n1883) );
  XOR U2070 ( .A(n1885), .B(n1950), .Z(n1886) );
  AND U2071 ( .A(e_input[8]), .B(g_input[9]), .Z(n1950) );
  XOR U2072 ( .A(n1891), .B(n1890), .Z(n1887) );
  XOR U2073 ( .A(n1889), .B(n1954), .Z(n1890) );
  AND U2074 ( .A(g_input[8]), .B(e_input[9]), .Z(n1954) );
  XOR U2075 ( .A(n1895), .B(n1894), .Z(n1891) );
  XOR U2076 ( .A(n1893), .B(n1958), .Z(n1894) );
  AND U2077 ( .A(g_input[7]), .B(e_input[10]), .Z(n1958) );
  XOR U2078 ( .A(n1899), .B(n1898), .Z(n1895) );
  XOR U2079 ( .A(n1897), .B(n1962), .Z(n1898) );
  AND U2080 ( .A(g_input[6]), .B(e_input[11]), .Z(n1962) );
  XOR U2081 ( .A(n1903), .B(n1902), .Z(n1899) );
  XOR U2082 ( .A(n1901), .B(n1966), .Z(n1902) );
  AND U2083 ( .A(g_input[5]), .B(e_input[12]), .Z(n1966) );
  XOR U2084 ( .A(n1907), .B(n1906), .Z(n1903) );
  XOR U2085 ( .A(n1905), .B(n1970), .Z(n1906) );
  AND U2086 ( .A(g_input[4]), .B(e_input[13]), .Z(n1970) );
  XOR U2087 ( .A(n1911), .B(n1910), .Z(n1907) );
  XOR U2088 ( .A(n1909), .B(n1974), .Z(n1910) );
  AND U2089 ( .A(g_input[3]), .B(e_input[14]), .Z(n1974) );
  XNOR U2090 ( .A(n1915), .B(n1914), .Z(n1911) );
  XOR U2091 ( .A(n1913), .B(n1978), .Z(n1914) );
  AND U2092 ( .A(g_input[2]), .B(e_input[15]), .Z(n1978) );
  XOR U2093 ( .A(n1918), .B(n1919), .Z(n1915) );
  NANDN U2094 ( .B(n532), .A(e_input[17]), .Z(n1919) );
  XNOR U2095 ( .A(n1917), .B(n1982), .Z(n1918) );
  AND U2096 ( .A(g_input[1]), .B(e_input[16]), .Z(n1982) );
  XNOR U2097 ( .A(n1922), .B(o[16]), .Z(oi[16]) );
  XNOR U2098 ( .A(n1986), .B(n1921), .Z(n1922) );
  XNOR U2099 ( .A(n1925), .B(n1924), .Z(n1986) );
  NAND U2100 ( .A(g_input[16]), .B(e_input[0]), .Z(n1924) );
  XOR U2101 ( .A(n1929), .B(n1928), .Z(n1925) );
  XNOR U2102 ( .A(n1989), .B(n1927), .Z(n1928) );
  NANDN U2103 ( .B(n1990), .A(n1991), .Z(n1927) );
  NAND U2104 ( .A(e_input[1]), .B(g_input[15]), .Z(n1989) );
  XOR U2105 ( .A(n1933), .B(n1932), .Z(n1929) );
  XNOR U2106 ( .A(n1931), .B(n1992), .Z(n1932) );
  AND U2107 ( .A(e_input[2]), .B(g_input[14]), .Z(n1992) );
  XOR U2108 ( .A(n1937), .B(n1936), .Z(n1933) );
  XOR U2109 ( .A(n1935), .B(n1996), .Z(n1936) );
  AND U2110 ( .A(e_input[3]), .B(g_input[13]), .Z(n1996) );
  XOR U2111 ( .A(n1941), .B(n1940), .Z(n1937) );
  XOR U2112 ( .A(n1939), .B(n2000), .Z(n1940) );
  AND U2113 ( .A(e_input[4]), .B(g_input[12]), .Z(n2000) );
  XOR U2114 ( .A(n1945), .B(n1944), .Z(n1941) );
  XOR U2115 ( .A(n1943), .B(n2004), .Z(n1944) );
  AND U2116 ( .A(e_input[5]), .B(g_input[11]), .Z(n2004) );
  XOR U2117 ( .A(n1949), .B(n1948), .Z(n1945) );
  XOR U2118 ( .A(n1947), .B(n2008), .Z(n1948) );
  AND U2119 ( .A(e_input[6]), .B(g_input[10]), .Z(n2008) );
  XOR U2120 ( .A(n1953), .B(n1952), .Z(n1949) );
  XOR U2121 ( .A(n1951), .B(n2012), .Z(n1952) );
  AND U2122 ( .A(e_input[7]), .B(g_input[9]), .Z(n2012) );
  XOR U2123 ( .A(n1957), .B(n1956), .Z(n1953) );
  XOR U2124 ( .A(n1955), .B(n2016), .Z(n1956) );
  AND U2125 ( .A(g_input[8]), .B(e_input[8]), .Z(n2016) );
  XOR U2126 ( .A(n1961), .B(n1960), .Z(n1957) );
  XOR U2127 ( .A(n1959), .B(n2020), .Z(n1960) );
  AND U2128 ( .A(g_input[7]), .B(e_input[9]), .Z(n2020) );
  XOR U2129 ( .A(n1965), .B(n1964), .Z(n1961) );
  XOR U2130 ( .A(n1963), .B(n2024), .Z(n1964) );
  AND U2131 ( .A(g_input[6]), .B(e_input[10]), .Z(n2024) );
  XOR U2132 ( .A(n1969), .B(n1968), .Z(n1965) );
  XOR U2133 ( .A(n1967), .B(n2028), .Z(n1968) );
  AND U2134 ( .A(g_input[5]), .B(e_input[11]), .Z(n2028) );
  XOR U2135 ( .A(n1973), .B(n1972), .Z(n1969) );
  XOR U2136 ( .A(n1971), .B(n2032), .Z(n1972) );
  AND U2137 ( .A(g_input[4]), .B(e_input[12]), .Z(n2032) );
  XOR U2138 ( .A(n1977), .B(n1976), .Z(n1973) );
  XOR U2139 ( .A(n1975), .B(n2036), .Z(n1976) );
  AND U2140 ( .A(g_input[3]), .B(e_input[13]), .Z(n2036) );
  XNOR U2141 ( .A(n1981), .B(n1980), .Z(n1977) );
  XOR U2142 ( .A(n1979), .B(n2040), .Z(n1980) );
  AND U2143 ( .A(g_input[2]), .B(e_input[14]), .Z(n2040) );
  XOR U2144 ( .A(n1984), .B(n1985), .Z(n1981) );
  NANDN U2145 ( .B(n532), .A(e_input[16]), .Z(n1985) );
  XNOR U2146 ( .A(n1983), .B(n2044), .Z(n1984) );
  AND U2147 ( .A(g_input[1]), .B(e_input[15]), .Z(n2044) );
  XNOR U2148 ( .A(n1988), .B(o[15]), .Z(oi[15]) );
  XNOR U2149 ( .A(n2048), .B(n1987), .Z(n1988) );
  XNOR U2150 ( .A(n1991), .B(n1990), .Z(n2048) );
  NAND U2151 ( .A(g_input[15]), .B(e_input[0]), .Z(n1990) );
  XOR U2152 ( .A(n1995), .B(n1994), .Z(n1991) );
  XNOR U2153 ( .A(n2051), .B(n1993), .Z(n1994) );
  NANDN U2154 ( .B(n2052), .A(n2053), .Z(n1993) );
  NAND U2155 ( .A(e_input[1]), .B(g_input[14]), .Z(n2051) );
  XOR U2156 ( .A(n1999), .B(n1998), .Z(n1995) );
  XNOR U2157 ( .A(n1997), .B(n2054), .Z(n1998) );
  AND U2158 ( .A(e_input[2]), .B(g_input[13]), .Z(n2054) );
  XOR U2159 ( .A(n2003), .B(n2002), .Z(n1999) );
  XOR U2160 ( .A(n2001), .B(n2058), .Z(n2002) );
  AND U2161 ( .A(e_input[3]), .B(g_input[12]), .Z(n2058) );
  XOR U2162 ( .A(n2007), .B(n2006), .Z(n2003) );
  XOR U2163 ( .A(n2005), .B(n2062), .Z(n2006) );
  AND U2164 ( .A(e_input[4]), .B(g_input[11]), .Z(n2062) );
  XOR U2165 ( .A(n2011), .B(n2010), .Z(n2007) );
  XOR U2166 ( .A(n2009), .B(n2066), .Z(n2010) );
  AND U2167 ( .A(e_input[5]), .B(g_input[10]), .Z(n2066) );
  XOR U2168 ( .A(n2015), .B(n2014), .Z(n2011) );
  XOR U2169 ( .A(n2013), .B(n2070), .Z(n2014) );
  AND U2170 ( .A(e_input[6]), .B(g_input[9]), .Z(n2070) );
  XOR U2171 ( .A(n2019), .B(n2018), .Z(n2015) );
  XOR U2172 ( .A(n2017), .B(n2074), .Z(n2018) );
  AND U2173 ( .A(e_input[7]), .B(g_input[8]), .Z(n2074) );
  XOR U2174 ( .A(n2023), .B(n2022), .Z(n2019) );
  XOR U2175 ( .A(n2021), .B(n2078), .Z(n2022) );
  AND U2176 ( .A(g_input[7]), .B(e_input[8]), .Z(n2078) );
  XOR U2177 ( .A(n2027), .B(n2026), .Z(n2023) );
  XOR U2178 ( .A(n2025), .B(n2082), .Z(n2026) );
  AND U2179 ( .A(g_input[6]), .B(e_input[9]), .Z(n2082) );
  XOR U2180 ( .A(n2031), .B(n2030), .Z(n2027) );
  XOR U2181 ( .A(n2029), .B(n2086), .Z(n2030) );
  AND U2182 ( .A(g_input[5]), .B(e_input[10]), .Z(n2086) );
  XOR U2183 ( .A(n2035), .B(n2034), .Z(n2031) );
  XOR U2184 ( .A(n2033), .B(n2090), .Z(n2034) );
  AND U2185 ( .A(g_input[4]), .B(e_input[11]), .Z(n2090) );
  XOR U2186 ( .A(n2039), .B(n2038), .Z(n2035) );
  XOR U2187 ( .A(n2037), .B(n2094), .Z(n2038) );
  AND U2188 ( .A(g_input[3]), .B(e_input[12]), .Z(n2094) );
  XNOR U2189 ( .A(n2043), .B(n2042), .Z(n2039) );
  XOR U2190 ( .A(n2041), .B(n2098), .Z(n2042) );
  AND U2191 ( .A(g_input[2]), .B(e_input[13]), .Z(n2098) );
  XOR U2192 ( .A(n2046), .B(n2047), .Z(n2043) );
  NANDN U2193 ( .B(n532), .A(e_input[15]), .Z(n2047) );
  XNOR U2194 ( .A(n2045), .B(n2102), .Z(n2046) );
  AND U2195 ( .A(g_input[1]), .B(e_input[14]), .Z(n2102) );
  XNOR U2196 ( .A(n2050), .B(o[14]), .Z(oi[14]) );
  XNOR U2197 ( .A(n2106), .B(n2049), .Z(n2050) );
  XNOR U2198 ( .A(n2053), .B(n2052), .Z(n2106) );
  NAND U2199 ( .A(g_input[14]), .B(e_input[0]), .Z(n2052) );
  XOR U2200 ( .A(n2057), .B(n2056), .Z(n2053) );
  XNOR U2201 ( .A(n2109), .B(n2055), .Z(n2056) );
  NANDN U2202 ( .B(n2110), .A(n2111), .Z(n2055) );
  NAND U2203 ( .A(e_input[1]), .B(g_input[13]), .Z(n2109) );
  XOR U2204 ( .A(n2061), .B(n2060), .Z(n2057) );
  XNOR U2205 ( .A(n2059), .B(n2112), .Z(n2060) );
  AND U2206 ( .A(e_input[2]), .B(g_input[12]), .Z(n2112) );
  XOR U2207 ( .A(n2065), .B(n2064), .Z(n2061) );
  XOR U2208 ( .A(n2063), .B(n2116), .Z(n2064) );
  AND U2209 ( .A(e_input[3]), .B(g_input[11]), .Z(n2116) );
  XOR U2210 ( .A(n2069), .B(n2068), .Z(n2065) );
  XOR U2211 ( .A(n2067), .B(n2120), .Z(n2068) );
  AND U2212 ( .A(e_input[4]), .B(g_input[10]), .Z(n2120) );
  XOR U2213 ( .A(n2073), .B(n2072), .Z(n2069) );
  XOR U2214 ( .A(n2071), .B(n2124), .Z(n2072) );
  AND U2215 ( .A(e_input[5]), .B(g_input[9]), .Z(n2124) );
  XOR U2216 ( .A(n2077), .B(n2076), .Z(n2073) );
  XOR U2217 ( .A(n2075), .B(n2128), .Z(n2076) );
  AND U2218 ( .A(e_input[6]), .B(g_input[8]), .Z(n2128) );
  XOR U2219 ( .A(n2081), .B(n2080), .Z(n2077) );
  XOR U2220 ( .A(n2079), .B(n2132), .Z(n2080) );
  AND U2221 ( .A(g_input[7]), .B(e_input[7]), .Z(n2132) );
  XOR U2222 ( .A(n2085), .B(n2084), .Z(n2081) );
  XOR U2223 ( .A(n2083), .B(n2136), .Z(n2084) );
  AND U2224 ( .A(g_input[6]), .B(e_input[8]), .Z(n2136) );
  XOR U2225 ( .A(n2089), .B(n2088), .Z(n2085) );
  XOR U2226 ( .A(n2087), .B(n2140), .Z(n2088) );
  AND U2227 ( .A(g_input[5]), .B(e_input[9]), .Z(n2140) );
  XOR U2228 ( .A(n2093), .B(n2092), .Z(n2089) );
  XOR U2229 ( .A(n2091), .B(n2144), .Z(n2092) );
  AND U2230 ( .A(g_input[4]), .B(e_input[10]), .Z(n2144) );
  XOR U2231 ( .A(n2097), .B(n2096), .Z(n2093) );
  XOR U2232 ( .A(n2095), .B(n2148), .Z(n2096) );
  AND U2233 ( .A(g_input[3]), .B(e_input[11]), .Z(n2148) );
  XNOR U2234 ( .A(n2101), .B(n2100), .Z(n2097) );
  XOR U2235 ( .A(n2099), .B(n2152), .Z(n2100) );
  AND U2236 ( .A(g_input[2]), .B(e_input[12]), .Z(n2152) );
  XOR U2237 ( .A(n2104), .B(n2105), .Z(n2101) );
  NANDN U2238 ( .B(n532), .A(e_input[14]), .Z(n2105) );
  XNOR U2239 ( .A(n2103), .B(n2156), .Z(n2104) );
  AND U2240 ( .A(g_input[1]), .B(e_input[13]), .Z(n2156) );
  XNOR U2241 ( .A(n2108), .B(o[13]), .Z(oi[13]) );
  XNOR U2242 ( .A(n2160), .B(n2107), .Z(n2108) );
  XNOR U2243 ( .A(n2111), .B(n2110), .Z(n2160) );
  NAND U2244 ( .A(g_input[13]), .B(e_input[0]), .Z(n2110) );
  XOR U2245 ( .A(n2115), .B(n2114), .Z(n2111) );
  XNOR U2246 ( .A(n2163), .B(n2113), .Z(n2114) );
  NANDN U2247 ( .B(n2164), .A(n2165), .Z(n2113) );
  NAND U2248 ( .A(e_input[1]), .B(g_input[12]), .Z(n2163) );
  XOR U2249 ( .A(n2119), .B(n2118), .Z(n2115) );
  XNOR U2250 ( .A(n2117), .B(n2166), .Z(n2118) );
  AND U2251 ( .A(e_input[2]), .B(g_input[11]), .Z(n2166) );
  XOR U2252 ( .A(n2123), .B(n2122), .Z(n2119) );
  XOR U2253 ( .A(n2121), .B(n2170), .Z(n2122) );
  AND U2254 ( .A(e_input[3]), .B(g_input[10]), .Z(n2170) );
  XOR U2255 ( .A(n2127), .B(n2126), .Z(n2123) );
  XOR U2256 ( .A(n2125), .B(n2174), .Z(n2126) );
  AND U2257 ( .A(e_input[4]), .B(g_input[9]), .Z(n2174) );
  XOR U2258 ( .A(n2131), .B(n2130), .Z(n2127) );
  XOR U2259 ( .A(n2129), .B(n2178), .Z(n2130) );
  AND U2260 ( .A(e_input[5]), .B(g_input[8]), .Z(n2178) );
  XOR U2261 ( .A(n2135), .B(n2134), .Z(n2131) );
  XOR U2262 ( .A(n2133), .B(n2182), .Z(n2134) );
  AND U2263 ( .A(e_input[6]), .B(g_input[7]), .Z(n2182) );
  XOR U2264 ( .A(n2139), .B(n2138), .Z(n2135) );
  XOR U2265 ( .A(n2137), .B(n2186), .Z(n2138) );
  AND U2266 ( .A(g_input[6]), .B(e_input[7]), .Z(n2186) );
  XOR U2267 ( .A(n2143), .B(n2142), .Z(n2139) );
  XOR U2268 ( .A(n2141), .B(n2190), .Z(n2142) );
  AND U2269 ( .A(g_input[5]), .B(e_input[8]), .Z(n2190) );
  XOR U2270 ( .A(n2147), .B(n2146), .Z(n2143) );
  XOR U2271 ( .A(n2145), .B(n2194), .Z(n2146) );
  AND U2272 ( .A(g_input[4]), .B(e_input[9]), .Z(n2194) );
  XOR U2273 ( .A(n2151), .B(n2150), .Z(n2147) );
  XOR U2274 ( .A(n2149), .B(n2198), .Z(n2150) );
  AND U2275 ( .A(g_input[3]), .B(e_input[10]), .Z(n2198) );
  XNOR U2276 ( .A(n2155), .B(n2154), .Z(n2151) );
  XOR U2277 ( .A(n2153), .B(n2202), .Z(n2154) );
  AND U2278 ( .A(g_input[2]), .B(e_input[11]), .Z(n2202) );
  XOR U2279 ( .A(n2158), .B(n2159), .Z(n2155) );
  NANDN U2280 ( .B(n532), .A(e_input[13]), .Z(n2159) );
  XNOR U2281 ( .A(n2157), .B(n2206), .Z(n2158) );
  AND U2282 ( .A(g_input[1]), .B(e_input[12]), .Z(n2206) );
  XNOR U2283 ( .A(n2162), .B(o[12]), .Z(oi[12]) );
  XNOR U2284 ( .A(n2210), .B(n2161), .Z(n2162) );
  XNOR U2285 ( .A(n2165), .B(n2164), .Z(n2210) );
  NAND U2286 ( .A(g_input[12]), .B(e_input[0]), .Z(n2164) );
  XOR U2287 ( .A(n2169), .B(n2168), .Z(n2165) );
  XNOR U2288 ( .A(n2213), .B(n2167), .Z(n2168) );
  NANDN U2289 ( .B(n2214), .A(n2215), .Z(n2167) );
  NAND U2290 ( .A(e_input[1]), .B(g_input[11]), .Z(n2213) );
  XOR U2291 ( .A(n2173), .B(n2172), .Z(n2169) );
  XNOR U2292 ( .A(n2171), .B(n2216), .Z(n2172) );
  AND U2293 ( .A(e_input[2]), .B(g_input[10]), .Z(n2216) );
  XOR U2294 ( .A(n2177), .B(n2176), .Z(n2173) );
  XOR U2295 ( .A(n2175), .B(n2220), .Z(n2176) );
  AND U2296 ( .A(e_input[3]), .B(g_input[9]), .Z(n2220) );
  XOR U2297 ( .A(n2181), .B(n2180), .Z(n2177) );
  XOR U2298 ( .A(n2179), .B(n2224), .Z(n2180) );
  AND U2299 ( .A(e_input[4]), .B(g_input[8]), .Z(n2224) );
  XNOR U2300 ( .A(n2228), .B(n2225), .Z(n2227) );
  XOR U2301 ( .A(n2185), .B(n2184), .Z(n2181) );
  XOR U2302 ( .A(n2183), .B(n2229), .Z(n2184) );
  AND U2303 ( .A(e_input[5]), .B(g_input[7]), .Z(n2229) );
  XOR U2304 ( .A(n2189), .B(n2188), .Z(n2185) );
  XOR U2305 ( .A(n2187), .B(n2233), .Z(n2188) );
  AND U2306 ( .A(g_input[6]), .B(e_input[6]), .Z(n2233) );
  XOR U2307 ( .A(n2193), .B(n2192), .Z(n2189) );
  XOR U2308 ( .A(n2191), .B(n2237), .Z(n2192) );
  AND U2309 ( .A(g_input[5]), .B(e_input[7]), .Z(n2237) );
  XOR U2310 ( .A(n2197), .B(n2196), .Z(n2193) );
  XOR U2311 ( .A(n2195), .B(n2241), .Z(n2196) );
  AND U2312 ( .A(g_input[4]), .B(e_input[8]), .Z(n2241) );
  XOR U2313 ( .A(n2201), .B(n2200), .Z(n2197) );
  XOR U2314 ( .A(n2199), .B(n2245), .Z(n2200) );
  AND U2315 ( .A(g_input[3]), .B(e_input[9]), .Z(n2245) );
  XNOR U2316 ( .A(n2205), .B(n2204), .Z(n2201) );
  XOR U2317 ( .A(n2203), .B(n2249), .Z(n2204) );
  AND U2318 ( .A(g_input[2]), .B(e_input[10]), .Z(n2249) );
  XOR U2319 ( .A(n2208), .B(n2209), .Z(n2205) );
  NANDN U2320 ( .B(n532), .A(e_input[12]), .Z(n2209) );
  XNOR U2321 ( .A(n2207), .B(n2253), .Z(n2208) );
  AND U2322 ( .A(g_input[1]), .B(e_input[11]), .Z(n2253) );
  XNOR U2323 ( .A(n2212), .B(o[11]), .Z(oi[11]) );
  XNOR U2324 ( .A(n2257), .B(n2211), .Z(n2212) );
  XNOR U2325 ( .A(n2215), .B(n2214), .Z(n2257) );
  NAND U2326 ( .A(g_input[11]), .B(e_input[0]), .Z(n2214) );
  XOR U2327 ( .A(n2219), .B(n2218), .Z(n2215) );
  XNOR U2328 ( .A(n2260), .B(n2217), .Z(n2218) );
  NANDN U2329 ( .B(n2261), .A(n2262), .Z(n2217) );
  NAND U2330 ( .A(e_input[1]), .B(g_input[10]), .Z(n2260) );
  XOR U2331 ( .A(n2223), .B(n2222), .Z(n2219) );
  XNOR U2332 ( .A(n2221), .B(n2263), .Z(n2222) );
  AND U2333 ( .A(e_input[2]), .B(g_input[9]), .Z(n2263) );
  XOR U2334 ( .A(n2228), .B(n2226), .Z(n2223) );
  XOR U2335 ( .A(n2225), .B(n2267), .Z(n2226) );
  AND U2336 ( .A(e_input[3]), .B(g_input[8]), .Z(n2267) );
  XOR U2337 ( .A(n2232), .B(n2231), .Z(n2228) );
  XOR U2338 ( .A(n2230), .B(n2271), .Z(n2231) );
  AND U2339 ( .A(e_input[4]), .B(g_input[7]), .Z(n2271) );
  XOR U2340 ( .A(n2236), .B(n2235), .Z(n2232) );
  XOR U2341 ( .A(n2234), .B(n2275), .Z(n2235) );
  AND U2342 ( .A(e_input[5]), .B(g_input[6]), .Z(n2275) );
  XOR U2343 ( .A(n2240), .B(n2239), .Z(n2236) );
  XOR U2344 ( .A(n2238), .B(n2279), .Z(n2239) );
  AND U2345 ( .A(g_input[5]), .B(e_input[6]), .Z(n2279) );
  XOR U2346 ( .A(n2244), .B(n2243), .Z(n2240) );
  XOR U2347 ( .A(n2242), .B(n2283), .Z(n2243) );
  AND U2348 ( .A(g_input[4]), .B(e_input[7]), .Z(n2283) );
  XOR U2349 ( .A(n2248), .B(n2247), .Z(n2244) );
  XOR U2350 ( .A(n2246), .B(n2287), .Z(n2247) );
  AND U2351 ( .A(g_input[3]), .B(e_input[8]), .Z(n2287) );
  XNOR U2352 ( .A(n2252), .B(n2251), .Z(n2248) );
  XOR U2353 ( .A(n2250), .B(n2291), .Z(n2251) );
  AND U2354 ( .A(g_input[2]), .B(e_input[9]), .Z(n2291) );
  XOR U2355 ( .A(n2255), .B(n2256), .Z(n2252) );
  NANDN U2356 ( .B(n532), .A(e_input[11]), .Z(n2256) );
  XNOR U2357 ( .A(n2254), .B(n2295), .Z(n2255) );
  AND U2358 ( .A(g_input[1]), .B(e_input[10]), .Z(n2295) );
  XNOR U2359 ( .A(n2259), .B(o[10]), .Z(oi[10]) );
  XNOR U2360 ( .A(n2299), .B(n2258), .Z(n2259) );
  XNOR U2361 ( .A(n2301), .B(n2302), .Z(n381) );
  XNOR U2362 ( .A(n2305), .B(n2306), .Z(n382) );
  XNOR U2363 ( .A(n2309), .B(n2310), .Z(n383) );
  XNOR U2364 ( .A(n2313), .B(n2314), .Z(n384) );
  XNOR U2365 ( .A(n2317), .B(n2318), .Z(n385) );
  XNOR U2366 ( .A(n2321), .B(n2322), .Z(n386) );
  XOR U2367 ( .A(n2325), .B(n2326), .Z(n387) );
  XNOR U2368 ( .A(n2328), .B(n2331), .Z(n2329) );
  XNOR U2369 ( .A(n2333), .B(n2334), .Z(n1775) );
  XOR U2370 ( .A(n2335), .B(n2332), .Z(n2333) );
  NANDN U2371 ( .B(n2336), .A(o[0]), .Z(n2332) );
  XNOR U2372 ( .A(n2262), .B(n2261), .Z(n2299) );
  NAND U2373 ( .A(g_input[10]), .B(e_input[0]), .Z(n2261) );
  XOR U2374 ( .A(n2266), .B(n2265), .Z(n2262) );
  XNOR U2375 ( .A(n2337), .B(n2264), .Z(n2265) );
  OR U2376 ( .A(n2302), .B(n2303), .Z(n2264) );
  NAND U2377 ( .A(g_input[9]), .B(e_input[0]), .Z(n2303) );
  NAND U2378 ( .A(e_input[1]), .B(g_input[9]), .Z(n2337) );
  XOR U2379 ( .A(n2270), .B(n2269), .Z(n2266) );
  XNOR U2380 ( .A(n2268), .B(n2340), .Z(n2269) );
  AND U2381 ( .A(e_input[2]), .B(g_input[8]), .Z(n2340) );
  XNOR U2382 ( .A(n2344), .B(n2341), .Z(n2339) );
  OR U2383 ( .A(n2306), .B(n2307), .Z(n2341) );
  NAND U2384 ( .A(g_input[8]), .B(e_input[0]), .Z(n2307) );
  NAND U2385 ( .A(e_input[1]), .B(g_input[8]), .Z(n2344) );
  XOR U2386 ( .A(n2274), .B(n2273), .Z(n2270) );
  XOR U2387 ( .A(n2272), .B(n2347), .Z(n2273) );
  AND U2388 ( .A(e_input[3]), .B(g_input[7]), .Z(n2347) );
  XNOR U2389 ( .A(n2348), .B(n2350), .Z(n2343) );
  AND U2390 ( .A(e_input[2]), .B(g_input[7]), .Z(n2350) );
  XNOR U2391 ( .A(n2342), .B(n2348), .Z(n2349) );
  XNOR U2392 ( .A(n2356), .B(n2353), .Z(n2346) );
  OR U2393 ( .A(n2310), .B(n2311), .Z(n2353) );
  NAND U2394 ( .A(g_input[7]), .B(e_input[0]), .Z(n2311) );
  NAND U2395 ( .A(e_input[1]), .B(g_input[7]), .Z(n2356) );
  XOR U2396 ( .A(n2278), .B(n2277), .Z(n2274) );
  XOR U2397 ( .A(n2276), .B(n2359), .Z(n2277) );
  AND U2398 ( .A(e_input[4]), .B(g_input[6]), .Z(n2359) );
  XNOR U2399 ( .A(n2360), .B(n2362), .Z(n2352) );
  AND U2400 ( .A(e_input[3]), .B(g_input[6]), .Z(n2362) );
  XNOR U2401 ( .A(n2351), .B(n2360), .Z(n2361) );
  XOR U2402 ( .A(n2365), .B(n2366), .Z(n2360) );
  ANDN U2403 ( .A(n2367), .B(n2355), .Z(n2366) );
  XNOR U2404 ( .A(n2365), .B(n2368), .Z(n2355) );
  AND U2405 ( .A(e_input[2]), .B(g_input[6]), .Z(n2368) );
  XNOR U2406 ( .A(n2354), .B(n2365), .Z(n2367) );
  XNOR U2407 ( .A(n2374), .B(n2371), .Z(n2358) );
  OR U2408 ( .A(n2314), .B(n2315), .Z(n2371) );
  NAND U2409 ( .A(g_input[6]), .B(e_input[0]), .Z(n2315) );
  NAND U2410 ( .A(e_input[1]), .B(g_input[6]), .Z(n2374) );
  XOR U2411 ( .A(n2282), .B(n2281), .Z(n2278) );
  XOR U2412 ( .A(n2280), .B(n2377), .Z(n2281) );
  AND U2413 ( .A(g_input[5]), .B(e_input[5]), .Z(n2377) );
  XOR U2414 ( .A(n2378), .B(n2379), .Z(n2280) );
  ANDN U2415 ( .A(n2380), .B(n2364), .Z(n2379) );
  XNOR U2416 ( .A(n2378), .B(n2381), .Z(n2364) );
  AND U2417 ( .A(e_input[4]), .B(g_input[5]), .Z(n2381) );
  XNOR U2418 ( .A(n2363), .B(n2378), .Z(n2380) );
  XNOR U2419 ( .A(n2384), .B(n2386), .Z(n2370) );
  AND U2420 ( .A(e_input[3]), .B(g_input[5]), .Z(n2386) );
  XNOR U2421 ( .A(n2369), .B(n2384), .Z(n2385) );
  XOR U2422 ( .A(n2389), .B(n2390), .Z(n2384) );
  ANDN U2423 ( .A(n2391), .B(n2373), .Z(n2390) );
  XNOR U2424 ( .A(n2389), .B(n2392), .Z(n2373) );
  AND U2425 ( .A(e_input[2]), .B(g_input[5]), .Z(n2392) );
  XNOR U2426 ( .A(n2372), .B(n2389), .Z(n2391) );
  XNOR U2427 ( .A(n2398), .B(n2395), .Z(n2376) );
  OR U2428 ( .A(n2318), .B(n2319), .Z(n2395) );
  NAND U2429 ( .A(g_input[5]), .B(e_input[0]), .Z(n2319) );
  NAND U2430 ( .A(e_input[1]), .B(g_input[5]), .Z(n2398) );
  XOR U2431 ( .A(n2286), .B(n2285), .Z(n2282) );
  XOR U2432 ( .A(n2284), .B(n2401), .Z(n2285) );
  AND U2433 ( .A(g_input[4]), .B(e_input[6]), .Z(n2401) );
  XNOR U2434 ( .A(n2402), .B(n2404), .Z(n2383) );
  AND U2435 ( .A(g_input[4]), .B(e_input[5]), .Z(n2404) );
  XNOR U2436 ( .A(n2382), .B(n2402), .Z(n2403) );
  XOR U2437 ( .A(n2407), .B(n2408), .Z(n2402) );
  ANDN U2438 ( .A(n2409), .B(n2388), .Z(n2408) );
  XNOR U2439 ( .A(n2407), .B(n2410), .Z(n2388) );
  AND U2440 ( .A(g_input[4]), .B(e_input[4]), .Z(n2410) );
  XNOR U2441 ( .A(n2387), .B(n2407), .Z(n2409) );
  XNOR U2442 ( .A(n2413), .B(n2415), .Z(n2394) );
  AND U2443 ( .A(e_input[3]), .B(g_input[4]), .Z(n2415) );
  XNOR U2444 ( .A(n2393), .B(n2413), .Z(n2414) );
  XOR U2445 ( .A(n2418), .B(n2419), .Z(n2413) );
  ANDN U2446 ( .A(n2420), .B(n2397), .Z(n2419) );
  XNOR U2447 ( .A(n2418), .B(n2421), .Z(n2397) );
  AND U2448 ( .A(e_input[2]), .B(g_input[4]), .Z(n2421) );
  XNOR U2449 ( .A(n2396), .B(n2418), .Z(n2420) );
  XNOR U2450 ( .A(n2427), .B(n2424), .Z(n2400) );
  OR U2451 ( .A(n2322), .B(n2323), .Z(n2424) );
  NAND U2452 ( .A(g_input[4]), .B(e_input[0]), .Z(n2323) );
  NAND U2453 ( .A(e_input[1]), .B(g_input[4]), .Z(n2427) );
  XOR U2454 ( .A(n2290), .B(n2289), .Z(n2286) );
  XOR U2455 ( .A(n2288), .B(n2430), .Z(n2289) );
  AND U2456 ( .A(g_input[3]), .B(e_input[7]), .Z(n2430) );
  XNOR U2457 ( .A(n2431), .B(n2432), .Z(n2406) );
  AND U2458 ( .A(g_input[3]), .B(e_input[6]), .Z(n2432) );
  XNOR U2459 ( .A(n2433), .B(n2434), .Z(n2405) );
  XNOR U2460 ( .A(n2435), .B(n2436), .Z(n2412) );
  AND U2461 ( .A(g_input[3]), .B(e_input[5]), .Z(n2436) );
  XNOR U2462 ( .A(n2437), .B(n2438), .Z(n2411) );
  XNOR U2463 ( .A(n2439), .B(n2440), .Z(n2417) );
  AND U2464 ( .A(g_input[3]), .B(e_input[4]), .Z(n2440) );
  XNOR U2465 ( .A(n2441), .B(n2442), .Z(n2416) );
  XNOR U2466 ( .A(n2443), .B(n2444), .Z(n2423) );
  AND U2467 ( .A(g_input[3]), .B(e_input[3]), .Z(n2444) );
  XNOR U2468 ( .A(n2445), .B(n2446), .Z(n2422) );
  XNOR U2469 ( .A(n2447), .B(n2448), .Z(n2426) );
  AND U2470 ( .A(e_input[2]), .B(g_input[3]), .Z(n2448) );
  XNOR U2471 ( .A(n2449), .B(n2450), .Z(n2425) );
  XNOR U2472 ( .A(n2452), .B(n2453), .Z(n2428) );
  XOR U2473 ( .A(n2454), .B(n2451), .Z(n2429) );
  ANDN U2474 ( .A(n2326), .B(n2327), .Z(n2451) );
  NAND U2475 ( .A(g_input[3]), .B(e_input[0]), .Z(n2327) );
  NAND U2476 ( .A(e_input[1]), .B(g_input[3]), .Z(n2454) );
  XNOR U2477 ( .A(n2294), .B(n2293), .Z(n2290) );
  XOR U2478 ( .A(n2292), .B(n2457), .Z(n2293) );
  AND U2479 ( .A(g_input[2]), .B(e_input[8]), .Z(n2457) );
  XNOR U2480 ( .A(n2458), .B(n2459), .Z(n2434) );
  AND U2481 ( .A(g_input[2]), .B(e_input[7]), .Z(n2459) );
  XNOR U2482 ( .A(n2460), .B(n2461), .Z(n2433) );
  XNOR U2483 ( .A(n2462), .B(n2463), .Z(n2438) );
  AND U2484 ( .A(g_input[2]), .B(e_input[6]), .Z(n2463) );
  XNOR U2485 ( .A(n2464), .B(n2465), .Z(n2437) );
  XNOR U2486 ( .A(n2466), .B(n2467), .Z(n2442) );
  AND U2487 ( .A(g_input[2]), .B(e_input[5]), .Z(n2467) );
  XNOR U2488 ( .A(n2468), .B(n2469), .Z(n2441) );
  XOR U2489 ( .A(n2470), .B(n2471), .Z(n2466) );
  ANDN U2490 ( .A(n2472), .B(n2446), .Z(n2471) );
  XNOR U2491 ( .A(n2470), .B(n2473), .Z(n2446) );
  AND U2492 ( .A(g_input[2]), .B(e_input[4]), .Z(n2473) );
  XNOR U2493 ( .A(n2445), .B(n2470), .Z(n2472) );
  XNOR U2494 ( .A(n2474), .B(n2475), .Z(n2445) );
  XNOR U2495 ( .A(n2476), .B(n2477), .Z(n2450) );
  AND U2496 ( .A(g_input[2]), .B(e_input[3]), .Z(n2477) );
  XNOR U2497 ( .A(n2478), .B(n2479), .Z(n2449) );
  XNOR U2498 ( .A(n2480), .B(n2481), .Z(n2453) );
  AND U2499 ( .A(g_input[2]), .B(e_input[2]), .Z(n2481) );
  XNOR U2500 ( .A(n2482), .B(n2483), .Z(n2452) );
  XNOR U2501 ( .A(n2485), .B(n2486), .Z(n2455) );
  XOR U2502 ( .A(n2487), .B(n2484), .Z(n2456) );
  NOR U2503 ( .A(n2330), .B(n2331), .Z(n2484) );
  NAND U2504 ( .A(g_input[2]), .B(e_input[0]), .Z(n2331) );
  XOR U2505 ( .A(n2488), .B(n2489), .Z(n2330) );
  NAND U2506 ( .A(e_input[1]), .B(g_input[2]), .Z(n2487) );
  XOR U2507 ( .A(n2297), .B(n2298), .Z(n2294) );
  NANDN U2508 ( .B(n532), .A(e_input[10]), .Z(n2298) );
  XNOR U2509 ( .A(n2296), .B(n2490), .Z(n2297) );
  AND U2510 ( .A(g_input[1]), .B(e_input[9]), .Z(n2490) );
  XNOR U2511 ( .A(n2491), .B(n2492), .Z(n2460) );
  AND U2512 ( .A(g_input[1]), .B(e_input[8]), .Z(n2492) );
  NANDN U2513 ( .B(n532), .A(e_input[9]), .Z(n2461) );
  XNOR U2514 ( .A(n2493), .B(n2494), .Z(n2464) );
  AND U2515 ( .A(g_input[1]), .B(e_input[7]), .Z(n2494) );
  NANDN U2516 ( .B(n532), .A(e_input[8]), .Z(n2465) );
  XNOR U2517 ( .A(n2495), .B(n2496), .Z(n2468) );
  AND U2518 ( .A(g_input[1]), .B(e_input[6]), .Z(n2496) );
  NANDN U2519 ( .B(n532), .A(e_input[7]), .Z(n2469) );
  XNOR U2520 ( .A(n2497), .B(n2498), .Z(n2474) );
  AND U2521 ( .A(g_input[1]), .B(e_input[5]), .Z(n2498) );
  NANDN U2522 ( .B(n532), .A(e_input[6]), .Z(n2475) );
  XNOR U2523 ( .A(n2499), .B(n2500), .Z(n2478) );
  AND U2524 ( .A(g_input[1]), .B(e_input[4]), .Z(n2500) );
  NANDN U2525 ( .B(n532), .A(e_input[5]), .Z(n2479) );
  XNOR U2526 ( .A(n2501), .B(n2502), .Z(n2482) );
  AND U2527 ( .A(g_input[1]), .B(e_input[3]), .Z(n2502) );
  NANDN U2528 ( .B(n532), .A(e_input[4]), .Z(n2483) );
  XOR U2529 ( .A(n2503), .B(n2504), .Z(n2485) );
  AND U2530 ( .A(g_input[1]), .B(e_input[2]), .Z(n2504) );
  NANDN U2531 ( .B(n532), .A(e_input[3]), .Z(n2486) );
  AND U2532 ( .A(n2505), .B(n2506), .Z(n2503) );
  NANDN U2533 ( .B(n2489), .A(n2488), .Z(n2505) );
  AND U2534 ( .A(n2507), .B(e_input[1]), .Z(n2488) );
  NANDN U2535 ( .B(n2334), .A(n2335), .Z(n2506) );
  AND U2536 ( .A(e_input[1]), .B(g_input[0]), .Z(n2335) );
  NAND U2537 ( .A(g_input[1]), .B(e_input[0]), .Z(n2334) );
  NANDN U2538 ( .B(n532), .A(e_input[2]), .Z(n2489) );
  XNOR U2539 ( .A(o[0]), .B(n2336), .Z(oi[0]) );
  NANDN U2540 ( .B(n532), .A(e_input[0]), .Z(n2336) );
  IV U2541 ( .A(g_input[0]), .Z(n532) );
endmodule

