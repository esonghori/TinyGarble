
module sum_N256_CC2 ( clk, rst, a, b, c );
  input [127:0] a;
  input [127:0] b;
  output [127:0] c;
  input clk, rst;
  wire   N258, N259, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912;
  wire   [1:0] carry_on;

  DFF \carry_on_reg[1]  ( .D(N259), .CLK(clk), .RST(rst), .Q(carry_on[1]) );
  DFF \carry_on_reg[0]  ( .D(N258), .CLK(clk), .RST(rst), .Q(carry_on[0]) );
  DFF \rc_reg[127]  ( .D(n512), .CLK(clk), .RST(1'b0), .Q(c[127]) );
  DFF \rc_reg[126]  ( .D(n511), .CLK(clk), .RST(1'b0), .Q(c[126]) );
  DFF \rc_reg[125]  ( .D(n510), .CLK(clk), .RST(1'b0), .Q(c[125]) );
  DFF \rc_reg[124]  ( .D(n509), .CLK(clk), .RST(1'b0), .Q(c[124]) );
  DFF \rc_reg[123]  ( .D(n508), .CLK(clk), .RST(1'b0), .Q(c[123]) );
  DFF \rc_reg[122]  ( .D(n507), .CLK(clk), .RST(1'b0), .Q(c[122]) );
  DFF \rc_reg[121]  ( .D(n506), .CLK(clk), .RST(1'b0), .Q(c[121]) );
  DFF \rc_reg[120]  ( .D(n505), .CLK(clk), .RST(1'b0), .Q(c[120]) );
  DFF \rc_reg[119]  ( .D(n504), .CLK(clk), .RST(1'b0), .Q(c[119]) );
  DFF \rc_reg[118]  ( .D(n503), .CLK(clk), .RST(1'b0), .Q(c[118]) );
  DFF \rc_reg[117]  ( .D(n502), .CLK(clk), .RST(1'b0), .Q(c[117]) );
  DFF \rc_reg[116]  ( .D(n501), .CLK(clk), .RST(1'b0), .Q(c[116]) );
  DFF \rc_reg[115]  ( .D(n500), .CLK(clk), .RST(1'b0), .Q(c[115]) );
  DFF \rc_reg[114]  ( .D(n499), .CLK(clk), .RST(1'b0), .Q(c[114]) );
  DFF \rc_reg[113]  ( .D(n498), .CLK(clk), .RST(1'b0), .Q(c[113]) );
  DFF \rc_reg[112]  ( .D(n497), .CLK(clk), .RST(1'b0), .Q(c[112]) );
  DFF \rc_reg[111]  ( .D(n496), .CLK(clk), .RST(1'b0), .Q(c[111]) );
  DFF \rc_reg[110]  ( .D(n495), .CLK(clk), .RST(1'b0), .Q(c[110]) );
  DFF \rc_reg[109]  ( .D(n494), .CLK(clk), .RST(1'b0), .Q(c[109]) );
  DFF \rc_reg[108]  ( .D(n493), .CLK(clk), .RST(1'b0), .Q(c[108]) );
  DFF \rc_reg[107]  ( .D(n492), .CLK(clk), .RST(1'b0), .Q(c[107]) );
  DFF \rc_reg[106]  ( .D(n491), .CLK(clk), .RST(1'b0), .Q(c[106]) );
  DFF \rc_reg[105]  ( .D(n490), .CLK(clk), .RST(1'b0), .Q(c[105]) );
  DFF \rc_reg[104]  ( .D(n489), .CLK(clk), .RST(1'b0), .Q(c[104]) );
  DFF \rc_reg[103]  ( .D(n488), .CLK(clk), .RST(1'b0), .Q(c[103]) );
  DFF \rc_reg[102]  ( .D(n487), .CLK(clk), .RST(1'b0), .Q(c[102]) );
  DFF \rc_reg[101]  ( .D(n486), .CLK(clk), .RST(1'b0), .Q(c[101]) );
  DFF \rc_reg[100]  ( .D(n485), .CLK(clk), .RST(1'b0), .Q(c[100]) );
  DFF \rc_reg[99]  ( .D(n484), .CLK(clk), .RST(1'b0), .Q(c[99]) );
  DFF \rc_reg[98]  ( .D(n483), .CLK(clk), .RST(1'b0), .Q(c[98]) );
  DFF \rc_reg[97]  ( .D(n482), .CLK(clk), .RST(1'b0), .Q(c[97]) );
  DFF \rc_reg[96]  ( .D(n481), .CLK(clk), .RST(1'b0), .Q(c[96]) );
  DFF \rc_reg[95]  ( .D(n480), .CLK(clk), .RST(1'b0), .Q(c[95]) );
  DFF \rc_reg[94]  ( .D(n479), .CLK(clk), .RST(1'b0), .Q(c[94]) );
  DFF \rc_reg[93]  ( .D(n478), .CLK(clk), .RST(1'b0), .Q(c[93]) );
  DFF \rc_reg[92]  ( .D(n477), .CLK(clk), .RST(1'b0), .Q(c[92]) );
  DFF \rc_reg[91]  ( .D(n476), .CLK(clk), .RST(1'b0), .Q(c[91]) );
  DFF \rc_reg[90]  ( .D(n475), .CLK(clk), .RST(1'b0), .Q(c[90]) );
  DFF \rc_reg[89]  ( .D(n474), .CLK(clk), .RST(1'b0), .Q(c[89]) );
  DFF \rc_reg[88]  ( .D(n473), .CLK(clk), .RST(1'b0), .Q(c[88]) );
  DFF \rc_reg[87]  ( .D(n472), .CLK(clk), .RST(1'b0), .Q(c[87]) );
  DFF \rc_reg[86]  ( .D(n471), .CLK(clk), .RST(1'b0), .Q(c[86]) );
  DFF \rc_reg[85]  ( .D(n470), .CLK(clk), .RST(1'b0), .Q(c[85]) );
  DFF \rc_reg[84]  ( .D(n469), .CLK(clk), .RST(1'b0), .Q(c[84]) );
  DFF \rc_reg[83]  ( .D(n468), .CLK(clk), .RST(1'b0), .Q(c[83]) );
  DFF \rc_reg[82]  ( .D(n467), .CLK(clk), .RST(1'b0), .Q(c[82]) );
  DFF \rc_reg[81]  ( .D(n466), .CLK(clk), .RST(1'b0), .Q(c[81]) );
  DFF \rc_reg[80]  ( .D(n465), .CLK(clk), .RST(1'b0), .Q(c[80]) );
  DFF \rc_reg[79]  ( .D(n464), .CLK(clk), .RST(1'b0), .Q(c[79]) );
  DFF \rc_reg[78]  ( .D(n463), .CLK(clk), .RST(1'b0), .Q(c[78]) );
  DFF \rc_reg[77]  ( .D(n462), .CLK(clk), .RST(1'b0), .Q(c[77]) );
  DFF \rc_reg[76]  ( .D(n461), .CLK(clk), .RST(1'b0), .Q(c[76]) );
  DFF \rc_reg[75]  ( .D(n460), .CLK(clk), .RST(1'b0), .Q(c[75]) );
  DFF \rc_reg[74]  ( .D(n459), .CLK(clk), .RST(1'b0), .Q(c[74]) );
  DFF \rc_reg[73]  ( .D(n458), .CLK(clk), .RST(1'b0), .Q(c[73]) );
  DFF \rc_reg[72]  ( .D(n457), .CLK(clk), .RST(1'b0), .Q(c[72]) );
  DFF \rc_reg[71]  ( .D(n456), .CLK(clk), .RST(1'b0), .Q(c[71]) );
  DFF \rc_reg[70]  ( .D(n455), .CLK(clk), .RST(1'b0), .Q(c[70]) );
  DFF \rc_reg[69]  ( .D(n454), .CLK(clk), .RST(1'b0), .Q(c[69]) );
  DFF \rc_reg[68]  ( .D(n453), .CLK(clk), .RST(1'b0), .Q(c[68]) );
  DFF \rc_reg[67]  ( .D(n452), .CLK(clk), .RST(1'b0), .Q(c[67]) );
  DFF \rc_reg[66]  ( .D(n451), .CLK(clk), .RST(1'b0), .Q(c[66]) );
  DFF \rc_reg[65]  ( .D(n450), .CLK(clk), .RST(1'b0), .Q(c[65]) );
  DFF \rc_reg[64]  ( .D(n449), .CLK(clk), .RST(1'b0), .Q(c[64]) );
  DFF \rc_reg[63]  ( .D(n448), .CLK(clk), .RST(1'b0), .Q(c[63]) );
  DFF \rc_reg[62]  ( .D(n447), .CLK(clk), .RST(1'b0), .Q(c[62]) );
  DFF \rc_reg[61]  ( .D(n446), .CLK(clk), .RST(1'b0), .Q(c[61]) );
  DFF \rc_reg[60]  ( .D(n445), .CLK(clk), .RST(1'b0), .Q(c[60]) );
  DFF \rc_reg[59]  ( .D(n444), .CLK(clk), .RST(1'b0), .Q(c[59]) );
  DFF \rc_reg[58]  ( .D(n443), .CLK(clk), .RST(1'b0), .Q(c[58]) );
  DFF \rc_reg[57]  ( .D(n442), .CLK(clk), .RST(1'b0), .Q(c[57]) );
  DFF \rc_reg[56]  ( .D(n441), .CLK(clk), .RST(1'b0), .Q(c[56]) );
  DFF \rc_reg[55]  ( .D(n440), .CLK(clk), .RST(1'b0), .Q(c[55]) );
  DFF \rc_reg[54]  ( .D(n439), .CLK(clk), .RST(1'b0), .Q(c[54]) );
  DFF \rc_reg[53]  ( .D(n438), .CLK(clk), .RST(1'b0), .Q(c[53]) );
  DFF \rc_reg[52]  ( .D(n437), .CLK(clk), .RST(1'b0), .Q(c[52]) );
  DFF \rc_reg[51]  ( .D(n436), .CLK(clk), .RST(1'b0), .Q(c[51]) );
  DFF \rc_reg[50]  ( .D(n435), .CLK(clk), .RST(1'b0), .Q(c[50]) );
  DFF \rc_reg[49]  ( .D(n434), .CLK(clk), .RST(1'b0), .Q(c[49]) );
  DFF \rc_reg[48]  ( .D(n433), .CLK(clk), .RST(1'b0), .Q(c[48]) );
  DFF \rc_reg[47]  ( .D(n432), .CLK(clk), .RST(1'b0), .Q(c[47]) );
  DFF \rc_reg[46]  ( .D(n431), .CLK(clk), .RST(1'b0), .Q(c[46]) );
  DFF \rc_reg[45]  ( .D(n430), .CLK(clk), .RST(1'b0), .Q(c[45]) );
  DFF \rc_reg[44]  ( .D(n429), .CLK(clk), .RST(1'b0), .Q(c[44]) );
  DFF \rc_reg[43]  ( .D(n428), .CLK(clk), .RST(1'b0), .Q(c[43]) );
  DFF \rc_reg[42]  ( .D(n427), .CLK(clk), .RST(1'b0), .Q(c[42]) );
  DFF \rc_reg[41]  ( .D(n426), .CLK(clk), .RST(1'b0), .Q(c[41]) );
  DFF \rc_reg[40]  ( .D(n425), .CLK(clk), .RST(1'b0), .Q(c[40]) );
  DFF \rc_reg[39]  ( .D(n424), .CLK(clk), .RST(1'b0), .Q(c[39]) );
  DFF \rc_reg[38]  ( .D(n423), .CLK(clk), .RST(1'b0), .Q(c[38]) );
  DFF \rc_reg[37]  ( .D(n422), .CLK(clk), .RST(1'b0), .Q(c[37]) );
  DFF \rc_reg[36]  ( .D(n421), .CLK(clk), .RST(1'b0), .Q(c[36]) );
  DFF \rc_reg[35]  ( .D(n420), .CLK(clk), .RST(1'b0), .Q(c[35]) );
  DFF \rc_reg[34]  ( .D(n419), .CLK(clk), .RST(1'b0), .Q(c[34]) );
  DFF \rc_reg[33]  ( .D(n418), .CLK(clk), .RST(1'b0), .Q(c[33]) );
  DFF \rc_reg[32]  ( .D(n417), .CLK(clk), .RST(1'b0), .Q(c[32]) );
  DFF \rc_reg[31]  ( .D(n416), .CLK(clk), .RST(1'b0), .Q(c[31]) );
  DFF \rc_reg[30]  ( .D(n415), .CLK(clk), .RST(1'b0), .Q(c[30]) );
  DFF \rc_reg[29]  ( .D(n414), .CLK(clk), .RST(1'b0), .Q(c[29]) );
  DFF \rc_reg[28]  ( .D(n413), .CLK(clk), .RST(1'b0), .Q(c[28]) );
  DFF \rc_reg[27]  ( .D(n412), .CLK(clk), .RST(1'b0), .Q(c[27]) );
  DFF \rc_reg[26]  ( .D(n411), .CLK(clk), .RST(1'b0), .Q(c[26]) );
  DFF \rc_reg[25]  ( .D(n410), .CLK(clk), .RST(1'b0), .Q(c[25]) );
  DFF \rc_reg[24]  ( .D(n409), .CLK(clk), .RST(1'b0), .Q(c[24]) );
  DFF \rc_reg[23]  ( .D(n408), .CLK(clk), .RST(1'b0), .Q(c[23]) );
  DFF \rc_reg[22]  ( .D(n407), .CLK(clk), .RST(1'b0), .Q(c[22]) );
  DFF \rc_reg[21]  ( .D(n406), .CLK(clk), .RST(1'b0), .Q(c[21]) );
  DFF \rc_reg[20]  ( .D(n405), .CLK(clk), .RST(1'b0), .Q(c[20]) );
  DFF \rc_reg[19]  ( .D(n404), .CLK(clk), .RST(1'b0), .Q(c[19]) );
  DFF \rc_reg[18]  ( .D(n403), .CLK(clk), .RST(1'b0), .Q(c[18]) );
  DFF \rc_reg[17]  ( .D(n402), .CLK(clk), .RST(1'b0), .Q(c[17]) );
  DFF \rc_reg[16]  ( .D(n401), .CLK(clk), .RST(1'b0), .Q(c[16]) );
  DFF \rc_reg[15]  ( .D(n400), .CLK(clk), .RST(1'b0), .Q(c[15]) );
  DFF \rc_reg[14]  ( .D(n399), .CLK(clk), .RST(1'b0), .Q(c[14]) );
  DFF \rc_reg[13]  ( .D(n398), .CLK(clk), .RST(1'b0), .Q(c[13]) );
  DFF \rc_reg[12]  ( .D(n397), .CLK(clk), .RST(1'b0), .Q(c[12]) );
  DFF \rc_reg[11]  ( .D(n396), .CLK(clk), .RST(1'b0), .Q(c[11]) );
  DFF \rc_reg[10]  ( .D(n395), .CLK(clk), .RST(1'b0), .Q(c[10]) );
  DFF \rc_reg[9]  ( .D(n394), .CLK(clk), .RST(1'b0), .Q(c[9]) );
  DFF \rc_reg[8]  ( .D(n393), .CLK(clk), .RST(1'b0), .Q(c[8]) );
  DFF \rc_reg[7]  ( .D(n392), .CLK(clk), .RST(1'b0), .Q(c[7]) );
  DFF \rc_reg[6]  ( .D(n391), .CLK(clk), .RST(1'b0), .Q(c[6]) );
  DFF \rc_reg[5]  ( .D(n390), .CLK(clk), .RST(1'b0), .Q(c[5]) );
  DFF \rc_reg[4]  ( .D(n389), .CLK(clk), .RST(1'b0), .Q(c[4]) );
  DFF \rc_reg[3]  ( .D(n388), .CLK(clk), .RST(1'b0), .Q(c[3]) );
  DFF \rc_reg[2]  ( .D(n387), .CLK(clk), .RST(1'b0), .Q(c[2]) );
  DFF \rc_reg[1]  ( .D(n386), .CLK(clk), .RST(1'b0), .Q(c[1]) );
  DFF \rc_reg[0]  ( .D(n385), .CLK(clk), .RST(1'b0), .Q(c[0]) );
  NANDN U515 ( .A(n1265), .B(n1266), .Z(n513) );
  NANDN U516 ( .A(n1899), .B(n1898), .Z(n514) );
  AND U517 ( .A(n513), .B(n514), .Z(n515) );
  NAND U518 ( .A(n1904), .B(n1903), .Z(n516) );
  NANDN U519 ( .A(n515), .B(n1267), .Z(n517) );
  AND U520 ( .A(n516), .B(n517), .Z(n1268) );
  XOR U521 ( .A(n572), .B(n571), .Z(n1318) );
  XOR U522 ( .A(n596), .B(n595), .Z(n1338) );
  XOR U523 ( .A(n620), .B(n619), .Z(n1358) );
  XOR U524 ( .A(n644), .B(n643), .Z(n1378) );
  XOR U525 ( .A(n668), .B(n667), .Z(n1398) );
  XOR U526 ( .A(n692), .B(n691), .Z(n1418) );
  XOR U527 ( .A(n716), .B(n715), .Z(n1438) );
  XOR U528 ( .A(n740), .B(n739), .Z(n1458) );
  XOR U529 ( .A(n764), .B(n763), .Z(n1478) );
  XOR U530 ( .A(n788), .B(n787), .Z(n1498) );
  XOR U531 ( .A(n812), .B(n811), .Z(n1518) );
  XOR U532 ( .A(n836), .B(n835), .Z(n1538) );
  XOR U533 ( .A(n860), .B(n859), .Z(n1558) );
  XOR U534 ( .A(n884), .B(n883), .Z(n1578) );
  XOR U535 ( .A(n908), .B(n907), .Z(n1598) );
  XOR U536 ( .A(n932), .B(n931), .Z(n1618) );
  XOR U537 ( .A(n956), .B(n955), .Z(n1638) );
  XOR U538 ( .A(n980), .B(n979), .Z(n1658) );
  XOR U539 ( .A(n1004), .B(n1003), .Z(n1678) );
  XOR U540 ( .A(n1028), .B(n1027), .Z(n1698) );
  XOR U541 ( .A(n1052), .B(n1051), .Z(n1718) );
  XOR U542 ( .A(n1076), .B(n1075), .Z(n1738) );
  XOR U543 ( .A(n1100), .B(n1099), .Z(n1758) );
  XOR U544 ( .A(n1124), .B(n1123), .Z(n1778) );
  XOR U545 ( .A(n1148), .B(n1147), .Z(n1798) );
  XOR U546 ( .A(n1172), .B(n1171), .Z(n1818) );
  XOR U547 ( .A(n1196), .B(n1195), .Z(n1838) );
  XOR U548 ( .A(n1220), .B(n1219), .Z(n1858) );
  XOR U549 ( .A(n1244), .B(n1243), .Z(n1878) );
  XOR U550 ( .A(n535), .B(n534), .Z(n1288) );
  XOR U551 ( .A(n560), .B(n559), .Z(n1308) );
  XOR U552 ( .A(n584), .B(n583), .Z(n1328) );
  XOR U553 ( .A(n608), .B(n607), .Z(n1348) );
  XOR U554 ( .A(n632), .B(n631), .Z(n1368) );
  XOR U555 ( .A(n656), .B(n655), .Z(n1388) );
  XOR U556 ( .A(n680), .B(n679), .Z(n1408) );
  XOR U557 ( .A(n704), .B(n703), .Z(n1428) );
  XOR U558 ( .A(n728), .B(n727), .Z(n1448) );
  XOR U559 ( .A(n752), .B(n751), .Z(n1468) );
  XOR U560 ( .A(n776), .B(n775), .Z(n1488) );
  XOR U561 ( .A(n800), .B(n799), .Z(n1508) );
  XOR U562 ( .A(n824), .B(n823), .Z(n1528) );
  XOR U563 ( .A(n848), .B(n847), .Z(n1548) );
  XOR U564 ( .A(n872), .B(n871), .Z(n1568) );
  XOR U565 ( .A(n896), .B(n895), .Z(n1588) );
  XOR U566 ( .A(n920), .B(n919), .Z(n1608) );
  XOR U567 ( .A(n944), .B(n943), .Z(n1628) );
  XOR U568 ( .A(n968), .B(n967), .Z(n1648) );
  XOR U569 ( .A(n992), .B(n991), .Z(n1668) );
  XOR U570 ( .A(n1016), .B(n1015), .Z(n1688) );
  XOR U571 ( .A(n1040), .B(n1039), .Z(n1708) );
  XOR U572 ( .A(n1064), .B(n1063), .Z(n1728) );
  XOR U573 ( .A(n1088), .B(n1087), .Z(n1748) );
  XOR U574 ( .A(n1112), .B(n1111), .Z(n1768) );
  XOR U575 ( .A(n1136), .B(n1135), .Z(n1788) );
  XOR U576 ( .A(n1160), .B(n1159), .Z(n1808) );
  XOR U577 ( .A(n1184), .B(n1183), .Z(n1828) );
  XOR U578 ( .A(n1208), .B(n1207), .Z(n1848) );
  XOR U579 ( .A(n1232), .B(n1231), .Z(n1868) );
  XOR U580 ( .A(n1256), .B(n1255), .Z(n1888) );
  AND U581 ( .A(b[127]), .B(a[127]), .Z(n1273) );
  NAND U582 ( .A(a[125]), .B(b[125]), .Z(n1267) );
  AND U583 ( .A(a[124]), .B(b[124]), .Z(n1265) );
  XNOR U584 ( .A(a[1]), .B(b[1]), .Z(n520) );
  XNOR U585 ( .A(carry_on[1]), .B(n520), .Z(n1279) );
  NAND U586 ( .A(a[0]), .B(b[0]), .Z(n519) );
  XOR U587 ( .A(a[0]), .B(b[0]), .Z(n1274) );
  NAND U588 ( .A(n1274), .B(carry_on[0]), .Z(n518) );
  NAND U589 ( .A(n519), .B(n518), .Z(n1278) );
  NAND U590 ( .A(n1279), .B(n1278), .Z(n522) );
  ANDN U591 ( .B(carry_on[1]), .A(n520), .Z(n523) );
  ANDN U592 ( .B(n522), .A(n523), .Z(n521) );
  NAND U593 ( .A(a[1]), .B(b[1]), .Z(n524) );
  NAND U594 ( .A(n521), .B(n524), .Z(n528) );
  XNOR U595 ( .A(n524), .B(n522), .Z(n526) );
  NAND U596 ( .A(n524), .B(n523), .Z(n525) );
  NAND U597 ( .A(n526), .B(n525), .Z(n1284) );
  XNOR U598 ( .A(a[2]), .B(b[2]), .Z(n1283) );
  NAND U599 ( .A(n1284), .B(n1283), .Z(n527) );
  NAND U600 ( .A(n528), .B(n527), .Z(n534) );
  NAND U601 ( .A(a[2]), .B(b[2]), .Z(n535) );
  AND U602 ( .A(n534), .B(n535), .Z(n530) );
  XOR U603 ( .A(a[3]), .B(b[3]), .Z(n1289) );
  ANDN U604 ( .B(n1288), .A(n1289), .Z(n529) );
  OR U605 ( .A(n530), .B(n529), .Z(n531) );
  AND U606 ( .A(a[3]), .B(b[3]), .Z(n533) );
  ANDN U607 ( .B(n531), .A(n533), .Z(n540) );
  NOR U608 ( .A(n535), .B(n534), .Z(n532) );
  XNOR U609 ( .A(n533), .B(n532), .Z(n538) );
  XOR U610 ( .A(n535), .B(n534), .Z(n536) );
  NAND U611 ( .A(n536), .B(n1289), .Z(n537) );
  NAND U612 ( .A(n538), .B(n537), .Z(n1294) );
  XNOR U613 ( .A(a[4]), .B(b[4]), .Z(n1293) );
  NAND U614 ( .A(n1294), .B(n1293), .Z(n539) );
  NANDN U615 ( .A(n540), .B(n539), .Z(n547) );
  AND U616 ( .A(a[4]), .B(b[4]), .Z(n541) );
  IV U617 ( .A(n541), .Z(n548) );
  AND U618 ( .A(n547), .B(n548), .Z(n543) );
  XOR U619 ( .A(a[5]), .B(b[5]), .Z(n1299) );
  XNOR U620 ( .A(n541), .B(n547), .Z(n1298) );
  NANDN U621 ( .A(n1299), .B(n1298), .Z(n542) );
  NANDN U622 ( .A(n543), .B(n542), .Z(n544) );
  AND U623 ( .A(a[5]), .B(b[5]), .Z(n546) );
  ANDN U624 ( .B(n544), .A(n546), .Z(n553) );
  NOR U625 ( .A(n548), .B(n547), .Z(n545) );
  XNOR U626 ( .A(n546), .B(n545), .Z(n551) );
  XOR U627 ( .A(n548), .B(n547), .Z(n549) );
  NAND U628 ( .A(n549), .B(n1299), .Z(n550) );
  NAND U629 ( .A(n551), .B(n550), .Z(n1304) );
  XNOR U630 ( .A(a[6]), .B(b[6]), .Z(n1303) );
  NAND U631 ( .A(n1304), .B(n1303), .Z(n552) );
  NANDN U632 ( .A(n553), .B(n552), .Z(n559) );
  NAND U633 ( .A(a[6]), .B(b[6]), .Z(n560) );
  AND U634 ( .A(n559), .B(n560), .Z(n555) );
  XOR U635 ( .A(a[7]), .B(b[7]), .Z(n1309) );
  ANDN U636 ( .B(n1308), .A(n1309), .Z(n554) );
  OR U637 ( .A(n555), .B(n554), .Z(n556) );
  AND U638 ( .A(a[7]), .B(b[7]), .Z(n558) );
  ANDN U639 ( .B(n556), .A(n558), .Z(n565) );
  NOR U640 ( .A(n560), .B(n559), .Z(n557) );
  XNOR U641 ( .A(n558), .B(n557), .Z(n563) );
  XOR U642 ( .A(n560), .B(n559), .Z(n561) );
  NAND U643 ( .A(n561), .B(n1309), .Z(n562) );
  NAND U644 ( .A(n563), .B(n562), .Z(n1314) );
  XNOR U645 ( .A(a[8]), .B(b[8]), .Z(n1313) );
  NAND U646 ( .A(n1314), .B(n1313), .Z(n564) );
  NANDN U647 ( .A(n565), .B(n564), .Z(n571) );
  NAND U648 ( .A(a[8]), .B(b[8]), .Z(n572) );
  AND U649 ( .A(n571), .B(n572), .Z(n567) );
  XOR U650 ( .A(a[9]), .B(b[9]), .Z(n1319) );
  ANDN U651 ( .B(n1318), .A(n1319), .Z(n566) );
  OR U652 ( .A(n567), .B(n566), .Z(n568) );
  AND U653 ( .A(a[9]), .B(b[9]), .Z(n570) );
  ANDN U654 ( .B(n568), .A(n570), .Z(n577) );
  NOR U655 ( .A(n572), .B(n571), .Z(n569) );
  XNOR U656 ( .A(n570), .B(n569), .Z(n575) );
  XOR U657 ( .A(n572), .B(n571), .Z(n573) );
  NAND U658 ( .A(n573), .B(n1319), .Z(n574) );
  NAND U659 ( .A(n575), .B(n574), .Z(n1324) );
  XNOR U660 ( .A(a[10]), .B(b[10]), .Z(n1323) );
  NAND U661 ( .A(n1324), .B(n1323), .Z(n576) );
  NANDN U662 ( .A(n577), .B(n576), .Z(n583) );
  NAND U663 ( .A(a[10]), .B(b[10]), .Z(n584) );
  AND U664 ( .A(n583), .B(n584), .Z(n579) );
  XOR U665 ( .A(a[11]), .B(b[11]), .Z(n1329) );
  ANDN U666 ( .B(n1328), .A(n1329), .Z(n578) );
  OR U667 ( .A(n579), .B(n578), .Z(n580) );
  AND U668 ( .A(a[11]), .B(b[11]), .Z(n582) );
  ANDN U669 ( .B(n580), .A(n582), .Z(n589) );
  NOR U670 ( .A(n584), .B(n583), .Z(n581) );
  XNOR U671 ( .A(n582), .B(n581), .Z(n587) );
  XOR U672 ( .A(n584), .B(n583), .Z(n585) );
  NAND U673 ( .A(n585), .B(n1329), .Z(n586) );
  NAND U674 ( .A(n587), .B(n586), .Z(n1334) );
  XNOR U675 ( .A(a[12]), .B(b[12]), .Z(n1333) );
  NAND U676 ( .A(n1334), .B(n1333), .Z(n588) );
  NANDN U677 ( .A(n589), .B(n588), .Z(n595) );
  NAND U678 ( .A(a[12]), .B(b[12]), .Z(n596) );
  AND U679 ( .A(n595), .B(n596), .Z(n591) );
  XOR U680 ( .A(a[13]), .B(b[13]), .Z(n1339) );
  ANDN U681 ( .B(n1338), .A(n1339), .Z(n590) );
  OR U682 ( .A(n591), .B(n590), .Z(n592) );
  AND U683 ( .A(a[13]), .B(b[13]), .Z(n594) );
  ANDN U684 ( .B(n592), .A(n594), .Z(n601) );
  NOR U685 ( .A(n596), .B(n595), .Z(n593) );
  XNOR U686 ( .A(n594), .B(n593), .Z(n599) );
  XOR U687 ( .A(n596), .B(n595), .Z(n597) );
  NAND U688 ( .A(n597), .B(n1339), .Z(n598) );
  NAND U689 ( .A(n599), .B(n598), .Z(n1344) );
  XNOR U690 ( .A(a[14]), .B(b[14]), .Z(n1343) );
  NAND U691 ( .A(n1344), .B(n1343), .Z(n600) );
  NANDN U692 ( .A(n601), .B(n600), .Z(n607) );
  NAND U693 ( .A(a[14]), .B(b[14]), .Z(n608) );
  AND U694 ( .A(n607), .B(n608), .Z(n603) );
  XOR U695 ( .A(a[15]), .B(b[15]), .Z(n1349) );
  ANDN U696 ( .B(n1348), .A(n1349), .Z(n602) );
  OR U697 ( .A(n603), .B(n602), .Z(n604) );
  AND U698 ( .A(a[15]), .B(b[15]), .Z(n606) );
  ANDN U699 ( .B(n604), .A(n606), .Z(n613) );
  NOR U700 ( .A(n608), .B(n607), .Z(n605) );
  XNOR U701 ( .A(n606), .B(n605), .Z(n611) );
  XOR U702 ( .A(n608), .B(n607), .Z(n609) );
  NAND U703 ( .A(n609), .B(n1349), .Z(n610) );
  NAND U704 ( .A(n611), .B(n610), .Z(n1354) );
  XNOR U705 ( .A(a[16]), .B(b[16]), .Z(n1353) );
  NAND U706 ( .A(n1354), .B(n1353), .Z(n612) );
  NANDN U707 ( .A(n613), .B(n612), .Z(n619) );
  NAND U708 ( .A(a[16]), .B(b[16]), .Z(n620) );
  AND U709 ( .A(n619), .B(n620), .Z(n615) );
  XOR U710 ( .A(a[17]), .B(b[17]), .Z(n1359) );
  ANDN U711 ( .B(n1358), .A(n1359), .Z(n614) );
  OR U712 ( .A(n615), .B(n614), .Z(n616) );
  AND U713 ( .A(a[17]), .B(b[17]), .Z(n618) );
  ANDN U714 ( .B(n616), .A(n618), .Z(n625) );
  NOR U715 ( .A(n620), .B(n619), .Z(n617) );
  XNOR U716 ( .A(n618), .B(n617), .Z(n623) );
  XOR U717 ( .A(n620), .B(n619), .Z(n621) );
  NAND U718 ( .A(n621), .B(n1359), .Z(n622) );
  NAND U719 ( .A(n623), .B(n622), .Z(n1364) );
  XNOR U720 ( .A(a[18]), .B(b[18]), .Z(n1363) );
  NAND U721 ( .A(n1364), .B(n1363), .Z(n624) );
  NANDN U722 ( .A(n625), .B(n624), .Z(n631) );
  NAND U723 ( .A(a[18]), .B(b[18]), .Z(n632) );
  AND U724 ( .A(n631), .B(n632), .Z(n627) );
  XOR U725 ( .A(a[19]), .B(b[19]), .Z(n1369) );
  ANDN U726 ( .B(n1368), .A(n1369), .Z(n626) );
  OR U727 ( .A(n627), .B(n626), .Z(n628) );
  AND U728 ( .A(a[19]), .B(b[19]), .Z(n630) );
  ANDN U729 ( .B(n628), .A(n630), .Z(n637) );
  NOR U730 ( .A(n632), .B(n631), .Z(n629) );
  XNOR U731 ( .A(n630), .B(n629), .Z(n635) );
  XOR U732 ( .A(n632), .B(n631), .Z(n633) );
  NAND U733 ( .A(n633), .B(n1369), .Z(n634) );
  NAND U734 ( .A(n635), .B(n634), .Z(n1374) );
  XNOR U735 ( .A(a[20]), .B(b[20]), .Z(n1373) );
  NAND U736 ( .A(n1374), .B(n1373), .Z(n636) );
  NANDN U737 ( .A(n637), .B(n636), .Z(n643) );
  NAND U738 ( .A(a[20]), .B(b[20]), .Z(n644) );
  AND U739 ( .A(n643), .B(n644), .Z(n639) );
  XOR U740 ( .A(a[21]), .B(b[21]), .Z(n1379) );
  ANDN U741 ( .B(n1378), .A(n1379), .Z(n638) );
  OR U742 ( .A(n639), .B(n638), .Z(n640) );
  AND U743 ( .A(a[21]), .B(b[21]), .Z(n642) );
  ANDN U744 ( .B(n640), .A(n642), .Z(n649) );
  NOR U745 ( .A(n644), .B(n643), .Z(n641) );
  XNOR U746 ( .A(n642), .B(n641), .Z(n647) );
  XOR U747 ( .A(n644), .B(n643), .Z(n645) );
  NAND U748 ( .A(n645), .B(n1379), .Z(n646) );
  NAND U749 ( .A(n647), .B(n646), .Z(n1384) );
  XNOR U750 ( .A(a[22]), .B(b[22]), .Z(n1383) );
  NAND U751 ( .A(n1384), .B(n1383), .Z(n648) );
  NANDN U752 ( .A(n649), .B(n648), .Z(n655) );
  NAND U753 ( .A(a[22]), .B(b[22]), .Z(n656) );
  AND U754 ( .A(n655), .B(n656), .Z(n651) );
  XOR U755 ( .A(a[23]), .B(b[23]), .Z(n1389) );
  ANDN U756 ( .B(n1388), .A(n1389), .Z(n650) );
  OR U757 ( .A(n651), .B(n650), .Z(n652) );
  AND U758 ( .A(a[23]), .B(b[23]), .Z(n654) );
  ANDN U759 ( .B(n652), .A(n654), .Z(n661) );
  NOR U760 ( .A(n656), .B(n655), .Z(n653) );
  XNOR U761 ( .A(n654), .B(n653), .Z(n659) );
  XOR U762 ( .A(n656), .B(n655), .Z(n657) );
  NAND U763 ( .A(n657), .B(n1389), .Z(n658) );
  NAND U764 ( .A(n659), .B(n658), .Z(n1394) );
  XNOR U765 ( .A(a[24]), .B(b[24]), .Z(n1393) );
  NAND U766 ( .A(n1394), .B(n1393), .Z(n660) );
  NANDN U767 ( .A(n661), .B(n660), .Z(n667) );
  NAND U768 ( .A(a[24]), .B(b[24]), .Z(n668) );
  AND U769 ( .A(n667), .B(n668), .Z(n663) );
  XOR U770 ( .A(a[25]), .B(b[25]), .Z(n1399) );
  ANDN U771 ( .B(n1398), .A(n1399), .Z(n662) );
  OR U772 ( .A(n663), .B(n662), .Z(n664) );
  AND U773 ( .A(a[25]), .B(b[25]), .Z(n666) );
  ANDN U774 ( .B(n664), .A(n666), .Z(n673) );
  NOR U775 ( .A(n668), .B(n667), .Z(n665) );
  XNOR U776 ( .A(n666), .B(n665), .Z(n671) );
  XOR U777 ( .A(n668), .B(n667), .Z(n669) );
  NAND U778 ( .A(n669), .B(n1399), .Z(n670) );
  NAND U779 ( .A(n671), .B(n670), .Z(n1404) );
  XNOR U780 ( .A(a[26]), .B(b[26]), .Z(n1403) );
  NAND U781 ( .A(n1404), .B(n1403), .Z(n672) );
  NANDN U782 ( .A(n673), .B(n672), .Z(n679) );
  NAND U783 ( .A(a[26]), .B(b[26]), .Z(n680) );
  AND U784 ( .A(n679), .B(n680), .Z(n675) );
  XOR U785 ( .A(a[27]), .B(b[27]), .Z(n1409) );
  ANDN U786 ( .B(n1408), .A(n1409), .Z(n674) );
  OR U787 ( .A(n675), .B(n674), .Z(n676) );
  AND U788 ( .A(a[27]), .B(b[27]), .Z(n678) );
  ANDN U789 ( .B(n676), .A(n678), .Z(n685) );
  NOR U790 ( .A(n680), .B(n679), .Z(n677) );
  XNOR U791 ( .A(n678), .B(n677), .Z(n683) );
  XOR U792 ( .A(n680), .B(n679), .Z(n681) );
  NAND U793 ( .A(n681), .B(n1409), .Z(n682) );
  NAND U794 ( .A(n683), .B(n682), .Z(n1414) );
  XNOR U795 ( .A(a[28]), .B(b[28]), .Z(n1413) );
  NAND U796 ( .A(n1414), .B(n1413), .Z(n684) );
  NANDN U797 ( .A(n685), .B(n684), .Z(n691) );
  NAND U798 ( .A(a[28]), .B(b[28]), .Z(n692) );
  AND U799 ( .A(n691), .B(n692), .Z(n687) );
  XOR U800 ( .A(a[29]), .B(b[29]), .Z(n1419) );
  ANDN U801 ( .B(n1418), .A(n1419), .Z(n686) );
  OR U802 ( .A(n687), .B(n686), .Z(n688) );
  AND U803 ( .A(a[29]), .B(b[29]), .Z(n690) );
  ANDN U804 ( .B(n688), .A(n690), .Z(n697) );
  NOR U805 ( .A(n692), .B(n691), .Z(n689) );
  XNOR U806 ( .A(n690), .B(n689), .Z(n695) );
  XOR U807 ( .A(n692), .B(n691), .Z(n693) );
  NAND U808 ( .A(n693), .B(n1419), .Z(n694) );
  NAND U809 ( .A(n695), .B(n694), .Z(n1424) );
  XNOR U810 ( .A(a[30]), .B(b[30]), .Z(n1423) );
  NAND U811 ( .A(n1424), .B(n1423), .Z(n696) );
  NANDN U812 ( .A(n697), .B(n696), .Z(n703) );
  NAND U813 ( .A(a[30]), .B(b[30]), .Z(n704) );
  AND U814 ( .A(n703), .B(n704), .Z(n699) );
  XOR U815 ( .A(a[31]), .B(b[31]), .Z(n1429) );
  ANDN U816 ( .B(n1428), .A(n1429), .Z(n698) );
  OR U817 ( .A(n699), .B(n698), .Z(n700) );
  AND U818 ( .A(a[31]), .B(b[31]), .Z(n702) );
  ANDN U819 ( .B(n700), .A(n702), .Z(n709) );
  NOR U820 ( .A(n704), .B(n703), .Z(n701) );
  XNOR U821 ( .A(n702), .B(n701), .Z(n707) );
  XOR U822 ( .A(n704), .B(n703), .Z(n705) );
  NAND U823 ( .A(n705), .B(n1429), .Z(n706) );
  NAND U824 ( .A(n707), .B(n706), .Z(n1434) );
  XNOR U825 ( .A(a[32]), .B(b[32]), .Z(n1433) );
  NAND U826 ( .A(n1434), .B(n1433), .Z(n708) );
  NANDN U827 ( .A(n709), .B(n708), .Z(n715) );
  NAND U828 ( .A(a[32]), .B(b[32]), .Z(n716) );
  AND U829 ( .A(n715), .B(n716), .Z(n711) );
  XOR U830 ( .A(a[33]), .B(b[33]), .Z(n1439) );
  ANDN U831 ( .B(n1438), .A(n1439), .Z(n710) );
  OR U832 ( .A(n711), .B(n710), .Z(n712) );
  AND U833 ( .A(a[33]), .B(b[33]), .Z(n714) );
  ANDN U834 ( .B(n712), .A(n714), .Z(n721) );
  NOR U835 ( .A(n716), .B(n715), .Z(n713) );
  XNOR U836 ( .A(n714), .B(n713), .Z(n719) );
  XOR U837 ( .A(n716), .B(n715), .Z(n717) );
  NAND U838 ( .A(n717), .B(n1439), .Z(n718) );
  NAND U839 ( .A(n719), .B(n718), .Z(n1444) );
  XNOR U840 ( .A(a[34]), .B(b[34]), .Z(n1443) );
  NAND U841 ( .A(n1444), .B(n1443), .Z(n720) );
  NANDN U842 ( .A(n721), .B(n720), .Z(n727) );
  NAND U843 ( .A(a[34]), .B(b[34]), .Z(n728) );
  AND U844 ( .A(n727), .B(n728), .Z(n723) );
  XOR U845 ( .A(a[35]), .B(b[35]), .Z(n1449) );
  ANDN U846 ( .B(n1448), .A(n1449), .Z(n722) );
  OR U847 ( .A(n723), .B(n722), .Z(n724) );
  AND U848 ( .A(a[35]), .B(b[35]), .Z(n726) );
  ANDN U849 ( .B(n724), .A(n726), .Z(n733) );
  NOR U850 ( .A(n728), .B(n727), .Z(n725) );
  XNOR U851 ( .A(n726), .B(n725), .Z(n731) );
  XOR U852 ( .A(n728), .B(n727), .Z(n729) );
  NAND U853 ( .A(n729), .B(n1449), .Z(n730) );
  NAND U854 ( .A(n731), .B(n730), .Z(n1454) );
  XNOR U855 ( .A(a[36]), .B(b[36]), .Z(n1453) );
  NAND U856 ( .A(n1454), .B(n1453), .Z(n732) );
  NANDN U857 ( .A(n733), .B(n732), .Z(n739) );
  NAND U858 ( .A(a[36]), .B(b[36]), .Z(n740) );
  AND U859 ( .A(n739), .B(n740), .Z(n735) );
  XOR U860 ( .A(a[37]), .B(b[37]), .Z(n1459) );
  ANDN U861 ( .B(n1458), .A(n1459), .Z(n734) );
  OR U862 ( .A(n735), .B(n734), .Z(n736) );
  AND U863 ( .A(a[37]), .B(b[37]), .Z(n738) );
  ANDN U864 ( .B(n736), .A(n738), .Z(n745) );
  NOR U865 ( .A(n740), .B(n739), .Z(n737) );
  XNOR U866 ( .A(n738), .B(n737), .Z(n743) );
  XOR U867 ( .A(n740), .B(n739), .Z(n741) );
  NAND U868 ( .A(n741), .B(n1459), .Z(n742) );
  NAND U869 ( .A(n743), .B(n742), .Z(n1464) );
  XNOR U870 ( .A(a[38]), .B(b[38]), .Z(n1463) );
  NAND U871 ( .A(n1464), .B(n1463), .Z(n744) );
  NANDN U872 ( .A(n745), .B(n744), .Z(n751) );
  NAND U873 ( .A(a[38]), .B(b[38]), .Z(n752) );
  AND U874 ( .A(n751), .B(n752), .Z(n747) );
  XOR U875 ( .A(a[39]), .B(b[39]), .Z(n1469) );
  ANDN U876 ( .B(n1468), .A(n1469), .Z(n746) );
  OR U877 ( .A(n747), .B(n746), .Z(n748) );
  AND U878 ( .A(a[39]), .B(b[39]), .Z(n750) );
  ANDN U879 ( .B(n748), .A(n750), .Z(n757) );
  NOR U880 ( .A(n752), .B(n751), .Z(n749) );
  XNOR U881 ( .A(n750), .B(n749), .Z(n755) );
  XOR U882 ( .A(n752), .B(n751), .Z(n753) );
  NAND U883 ( .A(n753), .B(n1469), .Z(n754) );
  NAND U884 ( .A(n755), .B(n754), .Z(n1474) );
  XNOR U885 ( .A(a[40]), .B(b[40]), .Z(n1473) );
  NAND U886 ( .A(n1474), .B(n1473), .Z(n756) );
  NANDN U887 ( .A(n757), .B(n756), .Z(n763) );
  NAND U888 ( .A(a[40]), .B(b[40]), .Z(n764) );
  AND U889 ( .A(n763), .B(n764), .Z(n759) );
  XOR U890 ( .A(a[41]), .B(b[41]), .Z(n1479) );
  ANDN U891 ( .B(n1478), .A(n1479), .Z(n758) );
  OR U892 ( .A(n759), .B(n758), .Z(n760) );
  AND U893 ( .A(a[41]), .B(b[41]), .Z(n762) );
  ANDN U894 ( .B(n760), .A(n762), .Z(n769) );
  NOR U895 ( .A(n764), .B(n763), .Z(n761) );
  XNOR U896 ( .A(n762), .B(n761), .Z(n767) );
  XOR U897 ( .A(n764), .B(n763), .Z(n765) );
  NAND U898 ( .A(n765), .B(n1479), .Z(n766) );
  NAND U899 ( .A(n767), .B(n766), .Z(n1484) );
  XNOR U900 ( .A(a[42]), .B(b[42]), .Z(n1483) );
  NAND U901 ( .A(n1484), .B(n1483), .Z(n768) );
  NANDN U902 ( .A(n769), .B(n768), .Z(n775) );
  NAND U903 ( .A(a[42]), .B(b[42]), .Z(n776) );
  AND U904 ( .A(n775), .B(n776), .Z(n771) );
  XOR U905 ( .A(a[43]), .B(b[43]), .Z(n1489) );
  ANDN U906 ( .B(n1488), .A(n1489), .Z(n770) );
  OR U907 ( .A(n771), .B(n770), .Z(n772) );
  AND U908 ( .A(a[43]), .B(b[43]), .Z(n774) );
  ANDN U909 ( .B(n772), .A(n774), .Z(n781) );
  NOR U910 ( .A(n776), .B(n775), .Z(n773) );
  XNOR U911 ( .A(n774), .B(n773), .Z(n779) );
  XOR U912 ( .A(n776), .B(n775), .Z(n777) );
  NAND U913 ( .A(n777), .B(n1489), .Z(n778) );
  NAND U914 ( .A(n779), .B(n778), .Z(n1494) );
  XNOR U915 ( .A(a[44]), .B(b[44]), .Z(n1493) );
  NAND U916 ( .A(n1494), .B(n1493), .Z(n780) );
  NANDN U917 ( .A(n781), .B(n780), .Z(n787) );
  NAND U918 ( .A(a[44]), .B(b[44]), .Z(n788) );
  AND U919 ( .A(n787), .B(n788), .Z(n783) );
  XOR U920 ( .A(a[45]), .B(b[45]), .Z(n1499) );
  ANDN U921 ( .B(n1498), .A(n1499), .Z(n782) );
  OR U922 ( .A(n783), .B(n782), .Z(n784) );
  AND U923 ( .A(a[45]), .B(b[45]), .Z(n786) );
  ANDN U924 ( .B(n784), .A(n786), .Z(n793) );
  NOR U925 ( .A(n788), .B(n787), .Z(n785) );
  XNOR U926 ( .A(n786), .B(n785), .Z(n791) );
  XOR U927 ( .A(n788), .B(n787), .Z(n789) );
  NAND U928 ( .A(n789), .B(n1499), .Z(n790) );
  NAND U929 ( .A(n791), .B(n790), .Z(n1504) );
  XNOR U930 ( .A(a[46]), .B(b[46]), .Z(n1503) );
  NAND U931 ( .A(n1504), .B(n1503), .Z(n792) );
  NANDN U932 ( .A(n793), .B(n792), .Z(n799) );
  NAND U933 ( .A(a[46]), .B(b[46]), .Z(n800) );
  AND U934 ( .A(n799), .B(n800), .Z(n795) );
  XOR U935 ( .A(a[47]), .B(b[47]), .Z(n1509) );
  ANDN U936 ( .B(n1508), .A(n1509), .Z(n794) );
  OR U937 ( .A(n795), .B(n794), .Z(n796) );
  AND U938 ( .A(a[47]), .B(b[47]), .Z(n798) );
  ANDN U939 ( .B(n796), .A(n798), .Z(n805) );
  NOR U940 ( .A(n800), .B(n799), .Z(n797) );
  XNOR U941 ( .A(n798), .B(n797), .Z(n803) );
  XOR U942 ( .A(n800), .B(n799), .Z(n801) );
  NAND U943 ( .A(n801), .B(n1509), .Z(n802) );
  NAND U944 ( .A(n803), .B(n802), .Z(n1514) );
  XNOR U945 ( .A(a[48]), .B(b[48]), .Z(n1513) );
  NAND U946 ( .A(n1514), .B(n1513), .Z(n804) );
  NANDN U947 ( .A(n805), .B(n804), .Z(n811) );
  NAND U948 ( .A(a[48]), .B(b[48]), .Z(n812) );
  AND U949 ( .A(n811), .B(n812), .Z(n807) );
  XOR U950 ( .A(a[49]), .B(b[49]), .Z(n1519) );
  ANDN U951 ( .B(n1518), .A(n1519), .Z(n806) );
  OR U952 ( .A(n807), .B(n806), .Z(n808) );
  AND U953 ( .A(a[49]), .B(b[49]), .Z(n810) );
  ANDN U954 ( .B(n808), .A(n810), .Z(n817) );
  NOR U955 ( .A(n812), .B(n811), .Z(n809) );
  XNOR U956 ( .A(n810), .B(n809), .Z(n815) );
  XOR U957 ( .A(n812), .B(n811), .Z(n813) );
  NAND U958 ( .A(n813), .B(n1519), .Z(n814) );
  NAND U959 ( .A(n815), .B(n814), .Z(n1524) );
  XNOR U960 ( .A(a[50]), .B(b[50]), .Z(n1523) );
  NAND U961 ( .A(n1524), .B(n1523), .Z(n816) );
  NANDN U962 ( .A(n817), .B(n816), .Z(n823) );
  NAND U963 ( .A(a[50]), .B(b[50]), .Z(n824) );
  AND U964 ( .A(n823), .B(n824), .Z(n819) );
  XOR U965 ( .A(a[51]), .B(b[51]), .Z(n1529) );
  ANDN U966 ( .B(n1528), .A(n1529), .Z(n818) );
  OR U967 ( .A(n819), .B(n818), .Z(n820) );
  AND U968 ( .A(a[51]), .B(b[51]), .Z(n822) );
  ANDN U969 ( .B(n820), .A(n822), .Z(n829) );
  NOR U970 ( .A(n824), .B(n823), .Z(n821) );
  XNOR U971 ( .A(n822), .B(n821), .Z(n827) );
  XOR U972 ( .A(n824), .B(n823), .Z(n825) );
  NAND U973 ( .A(n825), .B(n1529), .Z(n826) );
  NAND U974 ( .A(n827), .B(n826), .Z(n1534) );
  XNOR U975 ( .A(a[52]), .B(b[52]), .Z(n1533) );
  NAND U976 ( .A(n1534), .B(n1533), .Z(n828) );
  NANDN U977 ( .A(n829), .B(n828), .Z(n835) );
  NAND U978 ( .A(a[52]), .B(b[52]), .Z(n836) );
  AND U979 ( .A(n835), .B(n836), .Z(n831) );
  XOR U980 ( .A(a[53]), .B(b[53]), .Z(n1539) );
  ANDN U981 ( .B(n1538), .A(n1539), .Z(n830) );
  OR U982 ( .A(n831), .B(n830), .Z(n832) );
  AND U983 ( .A(a[53]), .B(b[53]), .Z(n834) );
  ANDN U984 ( .B(n832), .A(n834), .Z(n841) );
  NOR U985 ( .A(n836), .B(n835), .Z(n833) );
  XNOR U986 ( .A(n834), .B(n833), .Z(n839) );
  XOR U987 ( .A(n836), .B(n835), .Z(n837) );
  NAND U988 ( .A(n837), .B(n1539), .Z(n838) );
  NAND U989 ( .A(n839), .B(n838), .Z(n1544) );
  XNOR U990 ( .A(a[54]), .B(b[54]), .Z(n1543) );
  NAND U991 ( .A(n1544), .B(n1543), .Z(n840) );
  NANDN U992 ( .A(n841), .B(n840), .Z(n847) );
  NAND U993 ( .A(a[54]), .B(b[54]), .Z(n848) );
  AND U994 ( .A(n847), .B(n848), .Z(n843) );
  XOR U995 ( .A(a[55]), .B(b[55]), .Z(n1549) );
  ANDN U996 ( .B(n1548), .A(n1549), .Z(n842) );
  OR U997 ( .A(n843), .B(n842), .Z(n844) );
  AND U998 ( .A(a[55]), .B(b[55]), .Z(n846) );
  ANDN U999 ( .B(n844), .A(n846), .Z(n853) );
  NOR U1000 ( .A(n848), .B(n847), .Z(n845) );
  XNOR U1001 ( .A(n846), .B(n845), .Z(n851) );
  XOR U1002 ( .A(n848), .B(n847), .Z(n849) );
  NAND U1003 ( .A(n849), .B(n1549), .Z(n850) );
  NAND U1004 ( .A(n851), .B(n850), .Z(n1554) );
  XNOR U1005 ( .A(a[56]), .B(b[56]), .Z(n1553) );
  NAND U1006 ( .A(n1554), .B(n1553), .Z(n852) );
  NANDN U1007 ( .A(n853), .B(n852), .Z(n859) );
  NAND U1008 ( .A(a[56]), .B(b[56]), .Z(n860) );
  AND U1009 ( .A(n859), .B(n860), .Z(n855) );
  XOR U1010 ( .A(a[57]), .B(b[57]), .Z(n1559) );
  ANDN U1011 ( .B(n1558), .A(n1559), .Z(n854) );
  OR U1012 ( .A(n855), .B(n854), .Z(n856) );
  AND U1013 ( .A(a[57]), .B(b[57]), .Z(n858) );
  ANDN U1014 ( .B(n856), .A(n858), .Z(n865) );
  NOR U1015 ( .A(n860), .B(n859), .Z(n857) );
  XNOR U1016 ( .A(n858), .B(n857), .Z(n863) );
  XOR U1017 ( .A(n860), .B(n859), .Z(n861) );
  NAND U1018 ( .A(n861), .B(n1559), .Z(n862) );
  NAND U1019 ( .A(n863), .B(n862), .Z(n1564) );
  XNOR U1020 ( .A(a[58]), .B(b[58]), .Z(n1563) );
  NAND U1021 ( .A(n1564), .B(n1563), .Z(n864) );
  NANDN U1022 ( .A(n865), .B(n864), .Z(n871) );
  NAND U1023 ( .A(a[58]), .B(b[58]), .Z(n872) );
  AND U1024 ( .A(n871), .B(n872), .Z(n867) );
  XOR U1025 ( .A(a[59]), .B(b[59]), .Z(n1569) );
  ANDN U1026 ( .B(n1568), .A(n1569), .Z(n866) );
  OR U1027 ( .A(n867), .B(n866), .Z(n868) );
  AND U1028 ( .A(a[59]), .B(b[59]), .Z(n870) );
  ANDN U1029 ( .B(n868), .A(n870), .Z(n877) );
  NOR U1030 ( .A(n872), .B(n871), .Z(n869) );
  XNOR U1031 ( .A(n870), .B(n869), .Z(n875) );
  XOR U1032 ( .A(n872), .B(n871), .Z(n873) );
  NAND U1033 ( .A(n873), .B(n1569), .Z(n874) );
  NAND U1034 ( .A(n875), .B(n874), .Z(n1574) );
  XNOR U1035 ( .A(a[60]), .B(b[60]), .Z(n1573) );
  NAND U1036 ( .A(n1574), .B(n1573), .Z(n876) );
  NANDN U1037 ( .A(n877), .B(n876), .Z(n883) );
  NAND U1038 ( .A(a[60]), .B(b[60]), .Z(n884) );
  AND U1039 ( .A(n883), .B(n884), .Z(n879) );
  XOR U1040 ( .A(a[61]), .B(b[61]), .Z(n1579) );
  ANDN U1041 ( .B(n1578), .A(n1579), .Z(n878) );
  OR U1042 ( .A(n879), .B(n878), .Z(n880) );
  AND U1043 ( .A(a[61]), .B(b[61]), .Z(n882) );
  ANDN U1044 ( .B(n880), .A(n882), .Z(n889) );
  NOR U1045 ( .A(n884), .B(n883), .Z(n881) );
  XNOR U1046 ( .A(n882), .B(n881), .Z(n887) );
  XOR U1047 ( .A(n884), .B(n883), .Z(n885) );
  NAND U1048 ( .A(n885), .B(n1579), .Z(n886) );
  NAND U1049 ( .A(n887), .B(n886), .Z(n1584) );
  XNOR U1050 ( .A(a[62]), .B(b[62]), .Z(n1583) );
  NAND U1051 ( .A(n1584), .B(n1583), .Z(n888) );
  NANDN U1052 ( .A(n889), .B(n888), .Z(n895) );
  NAND U1053 ( .A(a[62]), .B(b[62]), .Z(n896) );
  AND U1054 ( .A(n895), .B(n896), .Z(n891) );
  XOR U1055 ( .A(a[63]), .B(b[63]), .Z(n1589) );
  ANDN U1056 ( .B(n1588), .A(n1589), .Z(n890) );
  OR U1057 ( .A(n891), .B(n890), .Z(n892) );
  AND U1058 ( .A(a[63]), .B(b[63]), .Z(n894) );
  ANDN U1059 ( .B(n892), .A(n894), .Z(n901) );
  NOR U1060 ( .A(n896), .B(n895), .Z(n893) );
  XNOR U1061 ( .A(n894), .B(n893), .Z(n899) );
  XOR U1062 ( .A(n896), .B(n895), .Z(n897) );
  NAND U1063 ( .A(n897), .B(n1589), .Z(n898) );
  NAND U1064 ( .A(n899), .B(n898), .Z(n1594) );
  XNOR U1065 ( .A(a[64]), .B(b[64]), .Z(n1593) );
  NAND U1066 ( .A(n1594), .B(n1593), .Z(n900) );
  NANDN U1067 ( .A(n901), .B(n900), .Z(n907) );
  NAND U1068 ( .A(a[64]), .B(b[64]), .Z(n908) );
  AND U1069 ( .A(n907), .B(n908), .Z(n903) );
  XOR U1070 ( .A(a[65]), .B(b[65]), .Z(n1599) );
  ANDN U1071 ( .B(n1598), .A(n1599), .Z(n902) );
  OR U1072 ( .A(n903), .B(n902), .Z(n904) );
  AND U1073 ( .A(a[65]), .B(b[65]), .Z(n906) );
  ANDN U1074 ( .B(n904), .A(n906), .Z(n913) );
  NOR U1075 ( .A(n908), .B(n907), .Z(n905) );
  XNOR U1076 ( .A(n906), .B(n905), .Z(n911) );
  XOR U1077 ( .A(n908), .B(n907), .Z(n909) );
  NAND U1078 ( .A(n909), .B(n1599), .Z(n910) );
  NAND U1079 ( .A(n911), .B(n910), .Z(n1604) );
  XNOR U1080 ( .A(a[66]), .B(b[66]), .Z(n1603) );
  NAND U1081 ( .A(n1604), .B(n1603), .Z(n912) );
  NANDN U1082 ( .A(n913), .B(n912), .Z(n919) );
  NAND U1083 ( .A(a[66]), .B(b[66]), .Z(n920) );
  AND U1084 ( .A(n919), .B(n920), .Z(n915) );
  XOR U1085 ( .A(a[67]), .B(b[67]), .Z(n1609) );
  ANDN U1086 ( .B(n1608), .A(n1609), .Z(n914) );
  OR U1087 ( .A(n915), .B(n914), .Z(n916) );
  AND U1088 ( .A(a[67]), .B(b[67]), .Z(n918) );
  ANDN U1089 ( .B(n916), .A(n918), .Z(n925) );
  NOR U1090 ( .A(n920), .B(n919), .Z(n917) );
  XNOR U1091 ( .A(n918), .B(n917), .Z(n923) );
  XOR U1092 ( .A(n920), .B(n919), .Z(n921) );
  NAND U1093 ( .A(n921), .B(n1609), .Z(n922) );
  NAND U1094 ( .A(n923), .B(n922), .Z(n1614) );
  XNOR U1095 ( .A(a[68]), .B(b[68]), .Z(n1613) );
  NAND U1096 ( .A(n1614), .B(n1613), .Z(n924) );
  NANDN U1097 ( .A(n925), .B(n924), .Z(n931) );
  NAND U1098 ( .A(a[68]), .B(b[68]), .Z(n932) );
  AND U1099 ( .A(n931), .B(n932), .Z(n927) );
  XOR U1100 ( .A(a[69]), .B(b[69]), .Z(n1619) );
  ANDN U1101 ( .B(n1618), .A(n1619), .Z(n926) );
  OR U1102 ( .A(n927), .B(n926), .Z(n928) );
  AND U1103 ( .A(a[69]), .B(b[69]), .Z(n930) );
  ANDN U1104 ( .B(n928), .A(n930), .Z(n937) );
  NOR U1105 ( .A(n932), .B(n931), .Z(n929) );
  XNOR U1106 ( .A(n930), .B(n929), .Z(n935) );
  XOR U1107 ( .A(n932), .B(n931), .Z(n933) );
  NAND U1108 ( .A(n933), .B(n1619), .Z(n934) );
  NAND U1109 ( .A(n935), .B(n934), .Z(n1624) );
  XNOR U1110 ( .A(a[70]), .B(b[70]), .Z(n1623) );
  NAND U1111 ( .A(n1624), .B(n1623), .Z(n936) );
  NANDN U1112 ( .A(n937), .B(n936), .Z(n943) );
  NAND U1113 ( .A(a[70]), .B(b[70]), .Z(n944) );
  AND U1114 ( .A(n943), .B(n944), .Z(n939) );
  XOR U1115 ( .A(a[71]), .B(b[71]), .Z(n1629) );
  ANDN U1116 ( .B(n1628), .A(n1629), .Z(n938) );
  OR U1117 ( .A(n939), .B(n938), .Z(n940) );
  AND U1118 ( .A(a[71]), .B(b[71]), .Z(n942) );
  ANDN U1119 ( .B(n940), .A(n942), .Z(n949) );
  NOR U1120 ( .A(n944), .B(n943), .Z(n941) );
  XNOR U1121 ( .A(n942), .B(n941), .Z(n947) );
  XOR U1122 ( .A(n944), .B(n943), .Z(n945) );
  NAND U1123 ( .A(n945), .B(n1629), .Z(n946) );
  NAND U1124 ( .A(n947), .B(n946), .Z(n1634) );
  XNOR U1125 ( .A(a[72]), .B(b[72]), .Z(n1633) );
  NAND U1126 ( .A(n1634), .B(n1633), .Z(n948) );
  NANDN U1127 ( .A(n949), .B(n948), .Z(n955) );
  NAND U1128 ( .A(a[72]), .B(b[72]), .Z(n956) );
  AND U1129 ( .A(n955), .B(n956), .Z(n951) );
  XOR U1130 ( .A(a[73]), .B(b[73]), .Z(n1639) );
  ANDN U1131 ( .B(n1638), .A(n1639), .Z(n950) );
  OR U1132 ( .A(n951), .B(n950), .Z(n952) );
  AND U1133 ( .A(a[73]), .B(b[73]), .Z(n954) );
  ANDN U1134 ( .B(n952), .A(n954), .Z(n961) );
  NOR U1135 ( .A(n956), .B(n955), .Z(n953) );
  XNOR U1136 ( .A(n954), .B(n953), .Z(n959) );
  XOR U1137 ( .A(n956), .B(n955), .Z(n957) );
  NAND U1138 ( .A(n957), .B(n1639), .Z(n958) );
  NAND U1139 ( .A(n959), .B(n958), .Z(n1644) );
  XNOR U1140 ( .A(a[74]), .B(b[74]), .Z(n1643) );
  NAND U1141 ( .A(n1644), .B(n1643), .Z(n960) );
  NANDN U1142 ( .A(n961), .B(n960), .Z(n967) );
  NAND U1143 ( .A(a[74]), .B(b[74]), .Z(n968) );
  AND U1144 ( .A(n967), .B(n968), .Z(n963) );
  XOR U1145 ( .A(a[75]), .B(b[75]), .Z(n1649) );
  ANDN U1146 ( .B(n1648), .A(n1649), .Z(n962) );
  OR U1147 ( .A(n963), .B(n962), .Z(n964) );
  AND U1148 ( .A(a[75]), .B(b[75]), .Z(n966) );
  ANDN U1149 ( .B(n964), .A(n966), .Z(n973) );
  NOR U1150 ( .A(n968), .B(n967), .Z(n965) );
  XNOR U1151 ( .A(n966), .B(n965), .Z(n971) );
  XOR U1152 ( .A(n968), .B(n967), .Z(n969) );
  NAND U1153 ( .A(n969), .B(n1649), .Z(n970) );
  NAND U1154 ( .A(n971), .B(n970), .Z(n1654) );
  XNOR U1155 ( .A(a[76]), .B(b[76]), .Z(n1653) );
  NAND U1156 ( .A(n1654), .B(n1653), .Z(n972) );
  NANDN U1157 ( .A(n973), .B(n972), .Z(n979) );
  NAND U1158 ( .A(a[76]), .B(b[76]), .Z(n980) );
  AND U1159 ( .A(n979), .B(n980), .Z(n975) );
  XOR U1160 ( .A(a[77]), .B(b[77]), .Z(n1659) );
  ANDN U1161 ( .B(n1658), .A(n1659), .Z(n974) );
  OR U1162 ( .A(n975), .B(n974), .Z(n976) );
  AND U1163 ( .A(a[77]), .B(b[77]), .Z(n978) );
  ANDN U1164 ( .B(n976), .A(n978), .Z(n985) );
  NOR U1165 ( .A(n980), .B(n979), .Z(n977) );
  XNOR U1166 ( .A(n978), .B(n977), .Z(n983) );
  XOR U1167 ( .A(n980), .B(n979), .Z(n981) );
  NAND U1168 ( .A(n981), .B(n1659), .Z(n982) );
  NAND U1169 ( .A(n983), .B(n982), .Z(n1664) );
  XNOR U1170 ( .A(a[78]), .B(b[78]), .Z(n1663) );
  NAND U1171 ( .A(n1664), .B(n1663), .Z(n984) );
  NANDN U1172 ( .A(n985), .B(n984), .Z(n991) );
  NAND U1173 ( .A(a[78]), .B(b[78]), .Z(n992) );
  AND U1174 ( .A(n991), .B(n992), .Z(n987) );
  XOR U1175 ( .A(a[79]), .B(b[79]), .Z(n1669) );
  ANDN U1176 ( .B(n1668), .A(n1669), .Z(n986) );
  OR U1177 ( .A(n987), .B(n986), .Z(n988) );
  AND U1178 ( .A(a[79]), .B(b[79]), .Z(n990) );
  ANDN U1179 ( .B(n988), .A(n990), .Z(n997) );
  NOR U1180 ( .A(n992), .B(n991), .Z(n989) );
  XNOR U1181 ( .A(n990), .B(n989), .Z(n995) );
  XOR U1182 ( .A(n992), .B(n991), .Z(n993) );
  NAND U1183 ( .A(n993), .B(n1669), .Z(n994) );
  NAND U1184 ( .A(n995), .B(n994), .Z(n1674) );
  XNOR U1185 ( .A(a[80]), .B(b[80]), .Z(n1673) );
  NAND U1186 ( .A(n1674), .B(n1673), .Z(n996) );
  NANDN U1187 ( .A(n997), .B(n996), .Z(n1003) );
  NAND U1188 ( .A(a[80]), .B(b[80]), .Z(n1004) );
  AND U1189 ( .A(n1003), .B(n1004), .Z(n999) );
  XOR U1190 ( .A(a[81]), .B(b[81]), .Z(n1679) );
  ANDN U1191 ( .B(n1678), .A(n1679), .Z(n998) );
  OR U1192 ( .A(n999), .B(n998), .Z(n1000) );
  AND U1193 ( .A(a[81]), .B(b[81]), .Z(n1002) );
  ANDN U1194 ( .B(n1000), .A(n1002), .Z(n1009) );
  NOR U1195 ( .A(n1004), .B(n1003), .Z(n1001) );
  XNOR U1196 ( .A(n1002), .B(n1001), .Z(n1007) );
  XOR U1197 ( .A(n1004), .B(n1003), .Z(n1005) );
  NAND U1198 ( .A(n1005), .B(n1679), .Z(n1006) );
  NAND U1199 ( .A(n1007), .B(n1006), .Z(n1684) );
  XNOR U1200 ( .A(a[82]), .B(b[82]), .Z(n1683) );
  NAND U1201 ( .A(n1684), .B(n1683), .Z(n1008) );
  NANDN U1202 ( .A(n1009), .B(n1008), .Z(n1015) );
  NAND U1203 ( .A(a[82]), .B(b[82]), .Z(n1016) );
  AND U1204 ( .A(n1015), .B(n1016), .Z(n1011) );
  XOR U1205 ( .A(a[83]), .B(b[83]), .Z(n1689) );
  ANDN U1206 ( .B(n1688), .A(n1689), .Z(n1010) );
  OR U1207 ( .A(n1011), .B(n1010), .Z(n1012) );
  AND U1208 ( .A(a[83]), .B(b[83]), .Z(n1014) );
  ANDN U1209 ( .B(n1012), .A(n1014), .Z(n1021) );
  NOR U1210 ( .A(n1016), .B(n1015), .Z(n1013) );
  XNOR U1211 ( .A(n1014), .B(n1013), .Z(n1019) );
  XOR U1212 ( .A(n1016), .B(n1015), .Z(n1017) );
  NAND U1213 ( .A(n1017), .B(n1689), .Z(n1018) );
  NAND U1214 ( .A(n1019), .B(n1018), .Z(n1694) );
  XNOR U1215 ( .A(a[84]), .B(b[84]), .Z(n1693) );
  NAND U1216 ( .A(n1694), .B(n1693), .Z(n1020) );
  NANDN U1217 ( .A(n1021), .B(n1020), .Z(n1027) );
  NAND U1218 ( .A(a[84]), .B(b[84]), .Z(n1028) );
  AND U1219 ( .A(n1027), .B(n1028), .Z(n1023) );
  XOR U1220 ( .A(a[85]), .B(b[85]), .Z(n1699) );
  ANDN U1221 ( .B(n1698), .A(n1699), .Z(n1022) );
  OR U1222 ( .A(n1023), .B(n1022), .Z(n1024) );
  AND U1223 ( .A(a[85]), .B(b[85]), .Z(n1026) );
  ANDN U1224 ( .B(n1024), .A(n1026), .Z(n1033) );
  NOR U1225 ( .A(n1028), .B(n1027), .Z(n1025) );
  XNOR U1226 ( .A(n1026), .B(n1025), .Z(n1031) );
  XOR U1227 ( .A(n1028), .B(n1027), .Z(n1029) );
  NAND U1228 ( .A(n1029), .B(n1699), .Z(n1030) );
  NAND U1229 ( .A(n1031), .B(n1030), .Z(n1704) );
  XNOR U1230 ( .A(a[86]), .B(b[86]), .Z(n1703) );
  NAND U1231 ( .A(n1704), .B(n1703), .Z(n1032) );
  NANDN U1232 ( .A(n1033), .B(n1032), .Z(n1039) );
  NAND U1233 ( .A(a[86]), .B(b[86]), .Z(n1040) );
  AND U1234 ( .A(n1039), .B(n1040), .Z(n1035) );
  XOR U1235 ( .A(a[87]), .B(b[87]), .Z(n1709) );
  ANDN U1236 ( .B(n1708), .A(n1709), .Z(n1034) );
  OR U1237 ( .A(n1035), .B(n1034), .Z(n1036) );
  AND U1238 ( .A(a[87]), .B(b[87]), .Z(n1038) );
  ANDN U1239 ( .B(n1036), .A(n1038), .Z(n1045) );
  NOR U1240 ( .A(n1040), .B(n1039), .Z(n1037) );
  XNOR U1241 ( .A(n1038), .B(n1037), .Z(n1043) );
  XOR U1242 ( .A(n1040), .B(n1039), .Z(n1041) );
  NAND U1243 ( .A(n1041), .B(n1709), .Z(n1042) );
  NAND U1244 ( .A(n1043), .B(n1042), .Z(n1714) );
  XNOR U1245 ( .A(a[88]), .B(b[88]), .Z(n1713) );
  NAND U1246 ( .A(n1714), .B(n1713), .Z(n1044) );
  NANDN U1247 ( .A(n1045), .B(n1044), .Z(n1051) );
  NAND U1248 ( .A(a[88]), .B(b[88]), .Z(n1052) );
  AND U1249 ( .A(n1051), .B(n1052), .Z(n1047) );
  XOR U1250 ( .A(a[89]), .B(b[89]), .Z(n1719) );
  ANDN U1251 ( .B(n1718), .A(n1719), .Z(n1046) );
  OR U1252 ( .A(n1047), .B(n1046), .Z(n1048) );
  AND U1253 ( .A(a[89]), .B(b[89]), .Z(n1050) );
  ANDN U1254 ( .B(n1048), .A(n1050), .Z(n1057) );
  NOR U1255 ( .A(n1052), .B(n1051), .Z(n1049) );
  XNOR U1256 ( .A(n1050), .B(n1049), .Z(n1055) );
  XOR U1257 ( .A(n1052), .B(n1051), .Z(n1053) );
  NAND U1258 ( .A(n1053), .B(n1719), .Z(n1054) );
  NAND U1259 ( .A(n1055), .B(n1054), .Z(n1724) );
  XNOR U1260 ( .A(a[90]), .B(b[90]), .Z(n1723) );
  NAND U1261 ( .A(n1724), .B(n1723), .Z(n1056) );
  NANDN U1262 ( .A(n1057), .B(n1056), .Z(n1063) );
  NAND U1263 ( .A(a[90]), .B(b[90]), .Z(n1064) );
  AND U1264 ( .A(n1063), .B(n1064), .Z(n1059) );
  XOR U1265 ( .A(a[91]), .B(b[91]), .Z(n1729) );
  ANDN U1266 ( .B(n1728), .A(n1729), .Z(n1058) );
  OR U1267 ( .A(n1059), .B(n1058), .Z(n1060) );
  AND U1268 ( .A(a[91]), .B(b[91]), .Z(n1062) );
  ANDN U1269 ( .B(n1060), .A(n1062), .Z(n1069) );
  NOR U1270 ( .A(n1064), .B(n1063), .Z(n1061) );
  XNOR U1271 ( .A(n1062), .B(n1061), .Z(n1067) );
  XOR U1272 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1273 ( .A(n1065), .B(n1729), .Z(n1066) );
  NAND U1274 ( .A(n1067), .B(n1066), .Z(n1734) );
  XNOR U1275 ( .A(a[92]), .B(b[92]), .Z(n1733) );
  NAND U1276 ( .A(n1734), .B(n1733), .Z(n1068) );
  NANDN U1277 ( .A(n1069), .B(n1068), .Z(n1075) );
  NAND U1278 ( .A(a[92]), .B(b[92]), .Z(n1076) );
  AND U1279 ( .A(n1075), .B(n1076), .Z(n1071) );
  XOR U1280 ( .A(a[93]), .B(b[93]), .Z(n1739) );
  ANDN U1281 ( .B(n1738), .A(n1739), .Z(n1070) );
  OR U1282 ( .A(n1071), .B(n1070), .Z(n1072) );
  AND U1283 ( .A(a[93]), .B(b[93]), .Z(n1074) );
  ANDN U1284 ( .B(n1072), .A(n1074), .Z(n1081) );
  NOR U1285 ( .A(n1076), .B(n1075), .Z(n1073) );
  XNOR U1286 ( .A(n1074), .B(n1073), .Z(n1079) );
  XOR U1287 ( .A(n1076), .B(n1075), .Z(n1077) );
  NAND U1288 ( .A(n1077), .B(n1739), .Z(n1078) );
  NAND U1289 ( .A(n1079), .B(n1078), .Z(n1744) );
  XNOR U1290 ( .A(a[94]), .B(b[94]), .Z(n1743) );
  NAND U1291 ( .A(n1744), .B(n1743), .Z(n1080) );
  NANDN U1292 ( .A(n1081), .B(n1080), .Z(n1087) );
  NAND U1293 ( .A(a[94]), .B(b[94]), .Z(n1088) );
  AND U1294 ( .A(n1087), .B(n1088), .Z(n1083) );
  XOR U1295 ( .A(a[95]), .B(b[95]), .Z(n1749) );
  ANDN U1296 ( .B(n1748), .A(n1749), .Z(n1082) );
  OR U1297 ( .A(n1083), .B(n1082), .Z(n1084) );
  AND U1298 ( .A(a[95]), .B(b[95]), .Z(n1086) );
  ANDN U1299 ( .B(n1084), .A(n1086), .Z(n1093) );
  NOR U1300 ( .A(n1088), .B(n1087), .Z(n1085) );
  XNOR U1301 ( .A(n1086), .B(n1085), .Z(n1091) );
  XOR U1302 ( .A(n1088), .B(n1087), .Z(n1089) );
  NAND U1303 ( .A(n1089), .B(n1749), .Z(n1090) );
  NAND U1304 ( .A(n1091), .B(n1090), .Z(n1754) );
  XNOR U1305 ( .A(a[96]), .B(b[96]), .Z(n1753) );
  NAND U1306 ( .A(n1754), .B(n1753), .Z(n1092) );
  NANDN U1307 ( .A(n1093), .B(n1092), .Z(n1099) );
  NAND U1308 ( .A(a[96]), .B(b[96]), .Z(n1100) );
  AND U1309 ( .A(n1099), .B(n1100), .Z(n1095) );
  XOR U1310 ( .A(a[97]), .B(b[97]), .Z(n1759) );
  ANDN U1311 ( .B(n1758), .A(n1759), .Z(n1094) );
  OR U1312 ( .A(n1095), .B(n1094), .Z(n1096) );
  AND U1313 ( .A(a[97]), .B(b[97]), .Z(n1098) );
  ANDN U1314 ( .B(n1096), .A(n1098), .Z(n1105) );
  NOR U1315 ( .A(n1100), .B(n1099), .Z(n1097) );
  XNOR U1316 ( .A(n1098), .B(n1097), .Z(n1103) );
  XOR U1317 ( .A(n1100), .B(n1099), .Z(n1101) );
  NAND U1318 ( .A(n1101), .B(n1759), .Z(n1102) );
  NAND U1319 ( .A(n1103), .B(n1102), .Z(n1764) );
  XNOR U1320 ( .A(a[98]), .B(b[98]), .Z(n1763) );
  NAND U1321 ( .A(n1764), .B(n1763), .Z(n1104) );
  NANDN U1322 ( .A(n1105), .B(n1104), .Z(n1111) );
  NAND U1323 ( .A(a[98]), .B(b[98]), .Z(n1112) );
  AND U1324 ( .A(n1111), .B(n1112), .Z(n1107) );
  XOR U1325 ( .A(a[99]), .B(b[99]), .Z(n1769) );
  ANDN U1326 ( .B(n1768), .A(n1769), .Z(n1106) );
  OR U1327 ( .A(n1107), .B(n1106), .Z(n1108) );
  AND U1328 ( .A(a[99]), .B(b[99]), .Z(n1110) );
  ANDN U1329 ( .B(n1108), .A(n1110), .Z(n1117) );
  NOR U1330 ( .A(n1112), .B(n1111), .Z(n1109) );
  XNOR U1331 ( .A(n1110), .B(n1109), .Z(n1115) );
  XOR U1332 ( .A(n1112), .B(n1111), .Z(n1113) );
  NAND U1333 ( .A(n1113), .B(n1769), .Z(n1114) );
  NAND U1334 ( .A(n1115), .B(n1114), .Z(n1774) );
  XNOR U1335 ( .A(a[100]), .B(b[100]), .Z(n1773) );
  NAND U1336 ( .A(n1774), .B(n1773), .Z(n1116) );
  NANDN U1337 ( .A(n1117), .B(n1116), .Z(n1123) );
  NAND U1338 ( .A(a[100]), .B(b[100]), .Z(n1124) );
  AND U1339 ( .A(n1123), .B(n1124), .Z(n1119) );
  XOR U1340 ( .A(a[101]), .B(b[101]), .Z(n1779) );
  ANDN U1341 ( .B(n1778), .A(n1779), .Z(n1118) );
  OR U1342 ( .A(n1119), .B(n1118), .Z(n1120) );
  AND U1343 ( .A(a[101]), .B(b[101]), .Z(n1122) );
  ANDN U1344 ( .B(n1120), .A(n1122), .Z(n1129) );
  NOR U1345 ( .A(n1124), .B(n1123), .Z(n1121) );
  XNOR U1346 ( .A(n1122), .B(n1121), .Z(n1127) );
  XOR U1347 ( .A(n1124), .B(n1123), .Z(n1125) );
  NAND U1348 ( .A(n1125), .B(n1779), .Z(n1126) );
  NAND U1349 ( .A(n1127), .B(n1126), .Z(n1784) );
  XNOR U1350 ( .A(a[102]), .B(b[102]), .Z(n1783) );
  NAND U1351 ( .A(n1784), .B(n1783), .Z(n1128) );
  NANDN U1352 ( .A(n1129), .B(n1128), .Z(n1135) );
  NAND U1353 ( .A(a[102]), .B(b[102]), .Z(n1136) );
  AND U1354 ( .A(n1135), .B(n1136), .Z(n1131) );
  XOR U1355 ( .A(a[103]), .B(b[103]), .Z(n1789) );
  ANDN U1356 ( .B(n1788), .A(n1789), .Z(n1130) );
  OR U1357 ( .A(n1131), .B(n1130), .Z(n1132) );
  AND U1358 ( .A(a[103]), .B(b[103]), .Z(n1134) );
  ANDN U1359 ( .B(n1132), .A(n1134), .Z(n1141) );
  NOR U1360 ( .A(n1136), .B(n1135), .Z(n1133) );
  XNOR U1361 ( .A(n1134), .B(n1133), .Z(n1139) );
  XOR U1362 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U1363 ( .A(n1137), .B(n1789), .Z(n1138) );
  NAND U1364 ( .A(n1139), .B(n1138), .Z(n1794) );
  XNOR U1365 ( .A(a[104]), .B(b[104]), .Z(n1793) );
  NAND U1366 ( .A(n1794), .B(n1793), .Z(n1140) );
  NANDN U1367 ( .A(n1141), .B(n1140), .Z(n1147) );
  NAND U1368 ( .A(a[104]), .B(b[104]), .Z(n1148) );
  AND U1369 ( .A(n1147), .B(n1148), .Z(n1143) );
  XOR U1370 ( .A(a[105]), .B(b[105]), .Z(n1799) );
  ANDN U1371 ( .B(n1798), .A(n1799), .Z(n1142) );
  OR U1372 ( .A(n1143), .B(n1142), .Z(n1144) );
  AND U1373 ( .A(a[105]), .B(b[105]), .Z(n1146) );
  ANDN U1374 ( .B(n1144), .A(n1146), .Z(n1153) );
  NOR U1375 ( .A(n1148), .B(n1147), .Z(n1145) );
  XNOR U1376 ( .A(n1146), .B(n1145), .Z(n1151) );
  XOR U1377 ( .A(n1148), .B(n1147), .Z(n1149) );
  NAND U1378 ( .A(n1149), .B(n1799), .Z(n1150) );
  NAND U1379 ( .A(n1151), .B(n1150), .Z(n1804) );
  XNOR U1380 ( .A(a[106]), .B(b[106]), .Z(n1803) );
  NAND U1381 ( .A(n1804), .B(n1803), .Z(n1152) );
  NANDN U1382 ( .A(n1153), .B(n1152), .Z(n1159) );
  NAND U1383 ( .A(a[106]), .B(b[106]), .Z(n1160) );
  AND U1384 ( .A(n1159), .B(n1160), .Z(n1155) );
  XOR U1385 ( .A(a[107]), .B(b[107]), .Z(n1809) );
  ANDN U1386 ( .B(n1808), .A(n1809), .Z(n1154) );
  OR U1387 ( .A(n1155), .B(n1154), .Z(n1156) );
  AND U1388 ( .A(a[107]), .B(b[107]), .Z(n1158) );
  ANDN U1389 ( .B(n1156), .A(n1158), .Z(n1165) );
  NOR U1390 ( .A(n1160), .B(n1159), .Z(n1157) );
  XNOR U1391 ( .A(n1158), .B(n1157), .Z(n1163) );
  XOR U1392 ( .A(n1160), .B(n1159), .Z(n1161) );
  NAND U1393 ( .A(n1161), .B(n1809), .Z(n1162) );
  NAND U1394 ( .A(n1163), .B(n1162), .Z(n1814) );
  XNOR U1395 ( .A(a[108]), .B(b[108]), .Z(n1813) );
  NAND U1396 ( .A(n1814), .B(n1813), .Z(n1164) );
  NANDN U1397 ( .A(n1165), .B(n1164), .Z(n1171) );
  NAND U1398 ( .A(a[108]), .B(b[108]), .Z(n1172) );
  AND U1399 ( .A(n1171), .B(n1172), .Z(n1167) );
  XOR U1400 ( .A(a[109]), .B(b[109]), .Z(n1819) );
  ANDN U1401 ( .B(n1818), .A(n1819), .Z(n1166) );
  OR U1402 ( .A(n1167), .B(n1166), .Z(n1168) );
  AND U1403 ( .A(a[109]), .B(b[109]), .Z(n1170) );
  ANDN U1404 ( .B(n1168), .A(n1170), .Z(n1177) );
  NOR U1405 ( .A(n1172), .B(n1171), .Z(n1169) );
  XNOR U1406 ( .A(n1170), .B(n1169), .Z(n1175) );
  XOR U1407 ( .A(n1172), .B(n1171), .Z(n1173) );
  NAND U1408 ( .A(n1173), .B(n1819), .Z(n1174) );
  NAND U1409 ( .A(n1175), .B(n1174), .Z(n1824) );
  XNOR U1410 ( .A(a[110]), .B(b[110]), .Z(n1823) );
  NAND U1411 ( .A(n1824), .B(n1823), .Z(n1176) );
  NANDN U1412 ( .A(n1177), .B(n1176), .Z(n1183) );
  NAND U1413 ( .A(a[110]), .B(b[110]), .Z(n1184) );
  AND U1414 ( .A(n1183), .B(n1184), .Z(n1179) );
  XOR U1415 ( .A(a[111]), .B(b[111]), .Z(n1829) );
  ANDN U1416 ( .B(n1828), .A(n1829), .Z(n1178) );
  OR U1417 ( .A(n1179), .B(n1178), .Z(n1180) );
  AND U1418 ( .A(a[111]), .B(b[111]), .Z(n1182) );
  ANDN U1419 ( .B(n1180), .A(n1182), .Z(n1189) );
  NOR U1420 ( .A(n1184), .B(n1183), .Z(n1181) );
  XNOR U1421 ( .A(n1182), .B(n1181), .Z(n1187) );
  XOR U1422 ( .A(n1184), .B(n1183), .Z(n1185) );
  NAND U1423 ( .A(n1185), .B(n1829), .Z(n1186) );
  NAND U1424 ( .A(n1187), .B(n1186), .Z(n1834) );
  XNOR U1425 ( .A(a[112]), .B(b[112]), .Z(n1833) );
  NAND U1426 ( .A(n1834), .B(n1833), .Z(n1188) );
  NANDN U1427 ( .A(n1189), .B(n1188), .Z(n1195) );
  NAND U1428 ( .A(a[112]), .B(b[112]), .Z(n1196) );
  AND U1429 ( .A(n1195), .B(n1196), .Z(n1191) );
  XOR U1430 ( .A(a[113]), .B(b[113]), .Z(n1839) );
  ANDN U1431 ( .B(n1838), .A(n1839), .Z(n1190) );
  OR U1432 ( .A(n1191), .B(n1190), .Z(n1192) );
  AND U1433 ( .A(a[113]), .B(b[113]), .Z(n1194) );
  ANDN U1434 ( .B(n1192), .A(n1194), .Z(n1201) );
  NOR U1435 ( .A(n1196), .B(n1195), .Z(n1193) );
  XNOR U1436 ( .A(n1194), .B(n1193), .Z(n1199) );
  XOR U1437 ( .A(n1196), .B(n1195), .Z(n1197) );
  NAND U1438 ( .A(n1197), .B(n1839), .Z(n1198) );
  NAND U1439 ( .A(n1199), .B(n1198), .Z(n1844) );
  XNOR U1440 ( .A(a[114]), .B(b[114]), .Z(n1843) );
  NAND U1441 ( .A(n1844), .B(n1843), .Z(n1200) );
  NANDN U1442 ( .A(n1201), .B(n1200), .Z(n1207) );
  NAND U1443 ( .A(a[114]), .B(b[114]), .Z(n1208) );
  AND U1444 ( .A(n1207), .B(n1208), .Z(n1203) );
  XOR U1445 ( .A(a[115]), .B(b[115]), .Z(n1849) );
  ANDN U1446 ( .B(n1848), .A(n1849), .Z(n1202) );
  OR U1447 ( .A(n1203), .B(n1202), .Z(n1204) );
  AND U1448 ( .A(a[115]), .B(b[115]), .Z(n1206) );
  ANDN U1449 ( .B(n1204), .A(n1206), .Z(n1213) );
  NOR U1450 ( .A(n1208), .B(n1207), .Z(n1205) );
  XNOR U1451 ( .A(n1206), .B(n1205), .Z(n1211) );
  XOR U1452 ( .A(n1208), .B(n1207), .Z(n1209) );
  NAND U1453 ( .A(n1209), .B(n1849), .Z(n1210) );
  NAND U1454 ( .A(n1211), .B(n1210), .Z(n1854) );
  XNOR U1455 ( .A(a[116]), .B(b[116]), .Z(n1853) );
  NAND U1456 ( .A(n1854), .B(n1853), .Z(n1212) );
  NANDN U1457 ( .A(n1213), .B(n1212), .Z(n1219) );
  NAND U1458 ( .A(a[116]), .B(b[116]), .Z(n1220) );
  AND U1459 ( .A(n1219), .B(n1220), .Z(n1215) );
  XOR U1460 ( .A(a[117]), .B(b[117]), .Z(n1859) );
  ANDN U1461 ( .B(n1858), .A(n1859), .Z(n1214) );
  OR U1462 ( .A(n1215), .B(n1214), .Z(n1216) );
  AND U1463 ( .A(a[117]), .B(b[117]), .Z(n1218) );
  ANDN U1464 ( .B(n1216), .A(n1218), .Z(n1225) );
  NOR U1465 ( .A(n1220), .B(n1219), .Z(n1217) );
  XNOR U1466 ( .A(n1218), .B(n1217), .Z(n1223) );
  XOR U1467 ( .A(n1220), .B(n1219), .Z(n1221) );
  NAND U1468 ( .A(n1221), .B(n1859), .Z(n1222) );
  NAND U1469 ( .A(n1223), .B(n1222), .Z(n1864) );
  XNOR U1470 ( .A(a[118]), .B(b[118]), .Z(n1863) );
  NAND U1471 ( .A(n1864), .B(n1863), .Z(n1224) );
  NANDN U1472 ( .A(n1225), .B(n1224), .Z(n1231) );
  NAND U1473 ( .A(a[118]), .B(b[118]), .Z(n1232) );
  AND U1474 ( .A(n1231), .B(n1232), .Z(n1227) );
  XOR U1475 ( .A(a[119]), .B(b[119]), .Z(n1869) );
  ANDN U1476 ( .B(n1868), .A(n1869), .Z(n1226) );
  OR U1477 ( .A(n1227), .B(n1226), .Z(n1228) );
  AND U1478 ( .A(a[119]), .B(b[119]), .Z(n1230) );
  ANDN U1479 ( .B(n1228), .A(n1230), .Z(n1237) );
  NOR U1480 ( .A(n1232), .B(n1231), .Z(n1229) );
  XNOR U1481 ( .A(n1230), .B(n1229), .Z(n1235) );
  XOR U1482 ( .A(n1232), .B(n1231), .Z(n1233) );
  NAND U1483 ( .A(n1233), .B(n1869), .Z(n1234) );
  NAND U1484 ( .A(n1235), .B(n1234), .Z(n1874) );
  XNOR U1485 ( .A(a[120]), .B(b[120]), .Z(n1873) );
  NAND U1486 ( .A(n1874), .B(n1873), .Z(n1236) );
  NANDN U1487 ( .A(n1237), .B(n1236), .Z(n1243) );
  NAND U1488 ( .A(a[120]), .B(b[120]), .Z(n1244) );
  AND U1489 ( .A(n1243), .B(n1244), .Z(n1239) );
  XOR U1490 ( .A(a[121]), .B(b[121]), .Z(n1879) );
  ANDN U1491 ( .B(n1878), .A(n1879), .Z(n1238) );
  OR U1492 ( .A(n1239), .B(n1238), .Z(n1240) );
  AND U1493 ( .A(a[121]), .B(b[121]), .Z(n1242) );
  ANDN U1494 ( .B(n1240), .A(n1242), .Z(n1249) );
  NOR U1495 ( .A(n1244), .B(n1243), .Z(n1241) );
  XNOR U1496 ( .A(n1242), .B(n1241), .Z(n1247) );
  XOR U1497 ( .A(n1244), .B(n1243), .Z(n1245) );
  NAND U1498 ( .A(n1245), .B(n1879), .Z(n1246) );
  NAND U1499 ( .A(n1247), .B(n1246), .Z(n1884) );
  XNOR U1500 ( .A(a[122]), .B(b[122]), .Z(n1883) );
  NAND U1501 ( .A(n1884), .B(n1883), .Z(n1248) );
  NANDN U1502 ( .A(n1249), .B(n1248), .Z(n1255) );
  NAND U1503 ( .A(a[122]), .B(b[122]), .Z(n1256) );
  AND U1504 ( .A(n1255), .B(n1256), .Z(n1251) );
  XOR U1505 ( .A(a[123]), .B(b[123]), .Z(n1889) );
  ANDN U1506 ( .B(n1888), .A(n1889), .Z(n1250) );
  OR U1507 ( .A(n1251), .B(n1250), .Z(n1252) );
  AND U1508 ( .A(a[123]), .B(b[123]), .Z(n1254) );
  ANDN U1509 ( .B(n1252), .A(n1254), .Z(n1261) );
  NOR U1510 ( .A(n1256), .B(n1255), .Z(n1253) );
  XNOR U1511 ( .A(n1254), .B(n1253), .Z(n1259) );
  XOR U1512 ( .A(n1256), .B(n1255), .Z(n1257) );
  NAND U1513 ( .A(n1257), .B(n1889), .Z(n1258) );
  NAND U1514 ( .A(n1259), .B(n1258), .Z(n1894) );
  XNOR U1515 ( .A(a[124]), .B(b[124]), .Z(n1893) );
  NAND U1516 ( .A(n1894), .B(n1893), .Z(n1260) );
  NANDN U1517 ( .A(n1261), .B(n1260), .Z(n1266) );
  ANDN U1518 ( .B(n1265), .A(n1266), .Z(n1262) );
  XOR U1519 ( .A(n1267), .B(n1262), .Z(n1264) );
  XOR U1520 ( .A(a[125]), .B(b[125]), .Z(n1899) );
  XNOR U1521 ( .A(n1265), .B(n1266), .Z(n1898) );
  NAND U1522 ( .A(n1899), .B(n1898), .Z(n1263) );
  NAND U1523 ( .A(n1264), .B(n1263), .Z(n1904) );
  XNOR U1524 ( .A(a[126]), .B(b[126]), .Z(n1903) );
  NAND U1525 ( .A(a[126]), .B(b[126]), .Z(n1269) );
  ANDN U1526 ( .B(n1268), .A(n1269), .Z(n1272) );
  XNOR U1527 ( .A(n1273), .B(n1272), .Z(n1271) );
  XNOR U1528 ( .A(n1269), .B(n1268), .Z(n1908) );
  XOR U1529 ( .A(b[127]), .B(a[127]), .Z(n1909) );
  NAND U1530 ( .A(n1908), .B(n1909), .Z(n1270) );
  NAND U1531 ( .A(n1271), .B(n1270), .Z(N258) );
  AND U1532 ( .A(n1273), .B(n1272), .Z(N259) );
  NAND U1534 ( .A(c[0]), .B(rst), .Z(n1277) );
  XOR U1535 ( .A(n1274), .B(carry_on[0]), .Z(n1275) );
  NANDN U1536 ( .A(rst), .B(n1275), .Z(n1276) );
  NAND U1537 ( .A(n1277), .B(n1276), .Z(n385) );
  NAND U1538 ( .A(c[1]), .B(rst), .Z(n1282) );
  XOR U1539 ( .A(n1279), .B(n1278), .Z(n1280) );
  NANDN U1540 ( .A(rst), .B(n1280), .Z(n1281) );
  NAND U1541 ( .A(n1282), .B(n1281), .Z(n386) );
  NAND U1542 ( .A(c[2]), .B(rst), .Z(n1287) );
  XNOR U1543 ( .A(n1284), .B(n1283), .Z(n1285) );
  NANDN U1544 ( .A(rst), .B(n1285), .Z(n1286) );
  NAND U1545 ( .A(n1287), .B(n1286), .Z(n387) );
  NAND U1546 ( .A(c[3]), .B(rst), .Z(n1292) );
  XOR U1547 ( .A(n1289), .B(n1288), .Z(n1290) );
  NANDN U1548 ( .A(rst), .B(n1290), .Z(n1291) );
  NAND U1549 ( .A(n1292), .B(n1291), .Z(n388) );
  NAND U1550 ( .A(c[4]), .B(rst), .Z(n1297) );
  XNOR U1551 ( .A(n1294), .B(n1293), .Z(n1295) );
  NANDN U1552 ( .A(rst), .B(n1295), .Z(n1296) );
  NAND U1553 ( .A(n1297), .B(n1296), .Z(n389) );
  NAND U1554 ( .A(c[5]), .B(rst), .Z(n1302) );
  XOR U1555 ( .A(n1299), .B(n1298), .Z(n1300) );
  NANDN U1556 ( .A(rst), .B(n1300), .Z(n1301) );
  NAND U1557 ( .A(n1302), .B(n1301), .Z(n390) );
  NAND U1558 ( .A(c[6]), .B(rst), .Z(n1307) );
  XNOR U1559 ( .A(n1304), .B(n1303), .Z(n1305) );
  NANDN U1560 ( .A(rst), .B(n1305), .Z(n1306) );
  NAND U1561 ( .A(n1307), .B(n1306), .Z(n391) );
  NAND U1562 ( .A(c[7]), .B(rst), .Z(n1312) );
  XOR U1563 ( .A(n1309), .B(n1308), .Z(n1310) );
  NANDN U1564 ( .A(rst), .B(n1310), .Z(n1311) );
  NAND U1565 ( .A(n1312), .B(n1311), .Z(n392) );
  NAND U1566 ( .A(c[8]), .B(rst), .Z(n1317) );
  XNOR U1567 ( .A(n1314), .B(n1313), .Z(n1315) );
  NANDN U1568 ( .A(rst), .B(n1315), .Z(n1316) );
  NAND U1569 ( .A(n1317), .B(n1316), .Z(n393) );
  NAND U1570 ( .A(c[9]), .B(rst), .Z(n1322) );
  XOR U1571 ( .A(n1319), .B(n1318), .Z(n1320) );
  NANDN U1572 ( .A(rst), .B(n1320), .Z(n1321) );
  NAND U1573 ( .A(n1322), .B(n1321), .Z(n394) );
  NAND U1574 ( .A(c[10]), .B(rst), .Z(n1327) );
  XNOR U1575 ( .A(n1324), .B(n1323), .Z(n1325) );
  NANDN U1576 ( .A(rst), .B(n1325), .Z(n1326) );
  NAND U1577 ( .A(n1327), .B(n1326), .Z(n395) );
  NAND U1578 ( .A(c[11]), .B(rst), .Z(n1332) );
  XOR U1579 ( .A(n1329), .B(n1328), .Z(n1330) );
  NANDN U1580 ( .A(rst), .B(n1330), .Z(n1331) );
  NAND U1581 ( .A(n1332), .B(n1331), .Z(n396) );
  NAND U1582 ( .A(c[12]), .B(rst), .Z(n1337) );
  XNOR U1583 ( .A(n1334), .B(n1333), .Z(n1335) );
  NANDN U1584 ( .A(rst), .B(n1335), .Z(n1336) );
  NAND U1585 ( .A(n1337), .B(n1336), .Z(n397) );
  NAND U1586 ( .A(c[13]), .B(rst), .Z(n1342) );
  XOR U1587 ( .A(n1339), .B(n1338), .Z(n1340) );
  NANDN U1588 ( .A(rst), .B(n1340), .Z(n1341) );
  NAND U1589 ( .A(n1342), .B(n1341), .Z(n398) );
  NAND U1590 ( .A(c[14]), .B(rst), .Z(n1347) );
  XNOR U1591 ( .A(n1344), .B(n1343), .Z(n1345) );
  NANDN U1592 ( .A(rst), .B(n1345), .Z(n1346) );
  NAND U1593 ( .A(n1347), .B(n1346), .Z(n399) );
  NAND U1594 ( .A(c[15]), .B(rst), .Z(n1352) );
  XOR U1595 ( .A(n1349), .B(n1348), .Z(n1350) );
  NANDN U1596 ( .A(rst), .B(n1350), .Z(n1351) );
  NAND U1597 ( .A(n1352), .B(n1351), .Z(n400) );
  NAND U1598 ( .A(c[16]), .B(rst), .Z(n1357) );
  XNOR U1599 ( .A(n1354), .B(n1353), .Z(n1355) );
  NANDN U1600 ( .A(rst), .B(n1355), .Z(n1356) );
  NAND U1601 ( .A(n1357), .B(n1356), .Z(n401) );
  NAND U1602 ( .A(c[17]), .B(rst), .Z(n1362) );
  XOR U1603 ( .A(n1359), .B(n1358), .Z(n1360) );
  NANDN U1604 ( .A(rst), .B(n1360), .Z(n1361) );
  NAND U1605 ( .A(n1362), .B(n1361), .Z(n402) );
  NAND U1606 ( .A(c[18]), .B(rst), .Z(n1367) );
  XNOR U1607 ( .A(n1364), .B(n1363), .Z(n1365) );
  NANDN U1608 ( .A(rst), .B(n1365), .Z(n1366) );
  NAND U1609 ( .A(n1367), .B(n1366), .Z(n403) );
  NAND U1610 ( .A(c[19]), .B(rst), .Z(n1372) );
  XOR U1611 ( .A(n1369), .B(n1368), .Z(n1370) );
  NANDN U1612 ( .A(rst), .B(n1370), .Z(n1371) );
  NAND U1613 ( .A(n1372), .B(n1371), .Z(n404) );
  NAND U1614 ( .A(c[20]), .B(rst), .Z(n1377) );
  XNOR U1615 ( .A(n1374), .B(n1373), .Z(n1375) );
  NANDN U1616 ( .A(rst), .B(n1375), .Z(n1376) );
  NAND U1617 ( .A(n1377), .B(n1376), .Z(n405) );
  NAND U1618 ( .A(c[21]), .B(rst), .Z(n1382) );
  XOR U1619 ( .A(n1379), .B(n1378), .Z(n1380) );
  NANDN U1620 ( .A(rst), .B(n1380), .Z(n1381) );
  NAND U1621 ( .A(n1382), .B(n1381), .Z(n406) );
  NAND U1622 ( .A(c[22]), .B(rst), .Z(n1387) );
  XNOR U1623 ( .A(n1384), .B(n1383), .Z(n1385) );
  NANDN U1624 ( .A(rst), .B(n1385), .Z(n1386) );
  NAND U1625 ( .A(n1387), .B(n1386), .Z(n407) );
  NAND U1626 ( .A(c[23]), .B(rst), .Z(n1392) );
  XOR U1627 ( .A(n1389), .B(n1388), .Z(n1390) );
  NANDN U1628 ( .A(rst), .B(n1390), .Z(n1391) );
  NAND U1629 ( .A(n1392), .B(n1391), .Z(n408) );
  NAND U1630 ( .A(c[24]), .B(rst), .Z(n1397) );
  XNOR U1631 ( .A(n1394), .B(n1393), .Z(n1395) );
  NANDN U1632 ( .A(rst), .B(n1395), .Z(n1396) );
  NAND U1633 ( .A(n1397), .B(n1396), .Z(n409) );
  NAND U1634 ( .A(c[25]), .B(rst), .Z(n1402) );
  XOR U1635 ( .A(n1399), .B(n1398), .Z(n1400) );
  NANDN U1636 ( .A(rst), .B(n1400), .Z(n1401) );
  NAND U1637 ( .A(n1402), .B(n1401), .Z(n410) );
  NAND U1638 ( .A(c[26]), .B(rst), .Z(n1407) );
  XNOR U1639 ( .A(n1404), .B(n1403), .Z(n1405) );
  NANDN U1640 ( .A(rst), .B(n1405), .Z(n1406) );
  NAND U1641 ( .A(n1407), .B(n1406), .Z(n411) );
  NAND U1642 ( .A(c[27]), .B(rst), .Z(n1412) );
  XOR U1643 ( .A(n1409), .B(n1408), .Z(n1410) );
  NANDN U1644 ( .A(rst), .B(n1410), .Z(n1411) );
  NAND U1645 ( .A(n1412), .B(n1411), .Z(n412) );
  NAND U1646 ( .A(c[28]), .B(rst), .Z(n1417) );
  XNOR U1647 ( .A(n1414), .B(n1413), .Z(n1415) );
  NANDN U1648 ( .A(rst), .B(n1415), .Z(n1416) );
  NAND U1649 ( .A(n1417), .B(n1416), .Z(n413) );
  NAND U1650 ( .A(c[29]), .B(rst), .Z(n1422) );
  XOR U1651 ( .A(n1419), .B(n1418), .Z(n1420) );
  NANDN U1652 ( .A(rst), .B(n1420), .Z(n1421) );
  NAND U1653 ( .A(n1422), .B(n1421), .Z(n414) );
  NAND U1654 ( .A(c[30]), .B(rst), .Z(n1427) );
  XNOR U1655 ( .A(n1424), .B(n1423), .Z(n1425) );
  NANDN U1656 ( .A(rst), .B(n1425), .Z(n1426) );
  NAND U1657 ( .A(n1427), .B(n1426), .Z(n415) );
  NAND U1658 ( .A(c[31]), .B(rst), .Z(n1432) );
  XOR U1659 ( .A(n1429), .B(n1428), .Z(n1430) );
  NANDN U1660 ( .A(rst), .B(n1430), .Z(n1431) );
  NAND U1661 ( .A(n1432), .B(n1431), .Z(n416) );
  NAND U1662 ( .A(c[32]), .B(rst), .Z(n1437) );
  XNOR U1663 ( .A(n1434), .B(n1433), .Z(n1435) );
  NANDN U1664 ( .A(rst), .B(n1435), .Z(n1436) );
  NAND U1665 ( .A(n1437), .B(n1436), .Z(n417) );
  NAND U1666 ( .A(c[33]), .B(rst), .Z(n1442) );
  XOR U1667 ( .A(n1439), .B(n1438), .Z(n1440) );
  NANDN U1668 ( .A(rst), .B(n1440), .Z(n1441) );
  NAND U1669 ( .A(n1442), .B(n1441), .Z(n418) );
  NAND U1670 ( .A(c[34]), .B(rst), .Z(n1447) );
  XNOR U1671 ( .A(n1444), .B(n1443), .Z(n1445) );
  NANDN U1672 ( .A(rst), .B(n1445), .Z(n1446) );
  NAND U1673 ( .A(n1447), .B(n1446), .Z(n419) );
  NAND U1674 ( .A(c[35]), .B(rst), .Z(n1452) );
  XOR U1675 ( .A(n1449), .B(n1448), .Z(n1450) );
  NANDN U1676 ( .A(rst), .B(n1450), .Z(n1451) );
  NAND U1677 ( .A(n1452), .B(n1451), .Z(n420) );
  NAND U1678 ( .A(c[36]), .B(rst), .Z(n1457) );
  XNOR U1679 ( .A(n1454), .B(n1453), .Z(n1455) );
  NANDN U1680 ( .A(rst), .B(n1455), .Z(n1456) );
  NAND U1681 ( .A(n1457), .B(n1456), .Z(n421) );
  NAND U1682 ( .A(c[37]), .B(rst), .Z(n1462) );
  XOR U1683 ( .A(n1459), .B(n1458), .Z(n1460) );
  NANDN U1684 ( .A(rst), .B(n1460), .Z(n1461) );
  NAND U1685 ( .A(n1462), .B(n1461), .Z(n422) );
  NAND U1686 ( .A(c[38]), .B(rst), .Z(n1467) );
  XNOR U1687 ( .A(n1464), .B(n1463), .Z(n1465) );
  NANDN U1688 ( .A(rst), .B(n1465), .Z(n1466) );
  NAND U1689 ( .A(n1467), .B(n1466), .Z(n423) );
  NAND U1690 ( .A(c[39]), .B(rst), .Z(n1472) );
  XOR U1691 ( .A(n1469), .B(n1468), .Z(n1470) );
  NANDN U1692 ( .A(rst), .B(n1470), .Z(n1471) );
  NAND U1693 ( .A(n1472), .B(n1471), .Z(n424) );
  NAND U1694 ( .A(c[40]), .B(rst), .Z(n1477) );
  XNOR U1695 ( .A(n1474), .B(n1473), .Z(n1475) );
  NANDN U1696 ( .A(rst), .B(n1475), .Z(n1476) );
  NAND U1697 ( .A(n1477), .B(n1476), .Z(n425) );
  NAND U1698 ( .A(c[41]), .B(rst), .Z(n1482) );
  XOR U1699 ( .A(n1479), .B(n1478), .Z(n1480) );
  NANDN U1700 ( .A(rst), .B(n1480), .Z(n1481) );
  NAND U1701 ( .A(n1482), .B(n1481), .Z(n426) );
  NAND U1702 ( .A(c[42]), .B(rst), .Z(n1487) );
  XNOR U1703 ( .A(n1484), .B(n1483), .Z(n1485) );
  NANDN U1704 ( .A(rst), .B(n1485), .Z(n1486) );
  NAND U1705 ( .A(n1487), .B(n1486), .Z(n427) );
  NAND U1706 ( .A(c[43]), .B(rst), .Z(n1492) );
  XOR U1707 ( .A(n1489), .B(n1488), .Z(n1490) );
  NANDN U1708 ( .A(rst), .B(n1490), .Z(n1491) );
  NAND U1709 ( .A(n1492), .B(n1491), .Z(n428) );
  NAND U1710 ( .A(c[44]), .B(rst), .Z(n1497) );
  XNOR U1711 ( .A(n1494), .B(n1493), .Z(n1495) );
  NANDN U1712 ( .A(rst), .B(n1495), .Z(n1496) );
  NAND U1713 ( .A(n1497), .B(n1496), .Z(n429) );
  NAND U1714 ( .A(c[45]), .B(rst), .Z(n1502) );
  XOR U1715 ( .A(n1499), .B(n1498), .Z(n1500) );
  NANDN U1716 ( .A(rst), .B(n1500), .Z(n1501) );
  NAND U1717 ( .A(n1502), .B(n1501), .Z(n430) );
  NAND U1718 ( .A(c[46]), .B(rst), .Z(n1507) );
  XNOR U1719 ( .A(n1504), .B(n1503), .Z(n1505) );
  NANDN U1720 ( .A(rst), .B(n1505), .Z(n1506) );
  NAND U1721 ( .A(n1507), .B(n1506), .Z(n431) );
  NAND U1722 ( .A(c[47]), .B(rst), .Z(n1512) );
  XOR U1723 ( .A(n1509), .B(n1508), .Z(n1510) );
  NANDN U1724 ( .A(rst), .B(n1510), .Z(n1511) );
  NAND U1725 ( .A(n1512), .B(n1511), .Z(n432) );
  NAND U1726 ( .A(c[48]), .B(rst), .Z(n1517) );
  XNOR U1727 ( .A(n1514), .B(n1513), .Z(n1515) );
  NANDN U1728 ( .A(rst), .B(n1515), .Z(n1516) );
  NAND U1729 ( .A(n1517), .B(n1516), .Z(n433) );
  NAND U1730 ( .A(c[49]), .B(rst), .Z(n1522) );
  XOR U1731 ( .A(n1519), .B(n1518), .Z(n1520) );
  NANDN U1732 ( .A(rst), .B(n1520), .Z(n1521) );
  NAND U1733 ( .A(n1522), .B(n1521), .Z(n434) );
  NAND U1734 ( .A(c[50]), .B(rst), .Z(n1527) );
  XNOR U1735 ( .A(n1524), .B(n1523), .Z(n1525) );
  NANDN U1736 ( .A(rst), .B(n1525), .Z(n1526) );
  NAND U1737 ( .A(n1527), .B(n1526), .Z(n435) );
  NAND U1738 ( .A(c[51]), .B(rst), .Z(n1532) );
  XOR U1739 ( .A(n1529), .B(n1528), .Z(n1530) );
  NANDN U1740 ( .A(rst), .B(n1530), .Z(n1531) );
  NAND U1741 ( .A(n1532), .B(n1531), .Z(n436) );
  NAND U1742 ( .A(c[52]), .B(rst), .Z(n1537) );
  XNOR U1743 ( .A(n1534), .B(n1533), .Z(n1535) );
  NANDN U1744 ( .A(rst), .B(n1535), .Z(n1536) );
  NAND U1745 ( .A(n1537), .B(n1536), .Z(n437) );
  NAND U1746 ( .A(c[53]), .B(rst), .Z(n1542) );
  XOR U1747 ( .A(n1539), .B(n1538), .Z(n1540) );
  NANDN U1748 ( .A(rst), .B(n1540), .Z(n1541) );
  NAND U1749 ( .A(n1542), .B(n1541), .Z(n438) );
  NAND U1750 ( .A(c[54]), .B(rst), .Z(n1547) );
  XNOR U1751 ( .A(n1544), .B(n1543), .Z(n1545) );
  NANDN U1752 ( .A(rst), .B(n1545), .Z(n1546) );
  NAND U1753 ( .A(n1547), .B(n1546), .Z(n439) );
  NAND U1754 ( .A(c[55]), .B(rst), .Z(n1552) );
  XOR U1755 ( .A(n1549), .B(n1548), .Z(n1550) );
  NANDN U1756 ( .A(rst), .B(n1550), .Z(n1551) );
  NAND U1757 ( .A(n1552), .B(n1551), .Z(n440) );
  NAND U1758 ( .A(c[56]), .B(rst), .Z(n1557) );
  XNOR U1759 ( .A(n1554), .B(n1553), .Z(n1555) );
  NANDN U1760 ( .A(rst), .B(n1555), .Z(n1556) );
  NAND U1761 ( .A(n1557), .B(n1556), .Z(n441) );
  NAND U1762 ( .A(c[57]), .B(rst), .Z(n1562) );
  XOR U1763 ( .A(n1559), .B(n1558), .Z(n1560) );
  NANDN U1764 ( .A(rst), .B(n1560), .Z(n1561) );
  NAND U1765 ( .A(n1562), .B(n1561), .Z(n442) );
  NAND U1766 ( .A(c[58]), .B(rst), .Z(n1567) );
  XNOR U1767 ( .A(n1564), .B(n1563), .Z(n1565) );
  NANDN U1768 ( .A(rst), .B(n1565), .Z(n1566) );
  NAND U1769 ( .A(n1567), .B(n1566), .Z(n443) );
  NAND U1770 ( .A(c[59]), .B(rst), .Z(n1572) );
  XOR U1771 ( .A(n1569), .B(n1568), .Z(n1570) );
  NANDN U1772 ( .A(rst), .B(n1570), .Z(n1571) );
  NAND U1773 ( .A(n1572), .B(n1571), .Z(n444) );
  NAND U1774 ( .A(c[60]), .B(rst), .Z(n1577) );
  XNOR U1775 ( .A(n1574), .B(n1573), .Z(n1575) );
  NANDN U1776 ( .A(rst), .B(n1575), .Z(n1576) );
  NAND U1777 ( .A(n1577), .B(n1576), .Z(n445) );
  NAND U1778 ( .A(c[61]), .B(rst), .Z(n1582) );
  XOR U1779 ( .A(n1579), .B(n1578), .Z(n1580) );
  NANDN U1780 ( .A(rst), .B(n1580), .Z(n1581) );
  NAND U1781 ( .A(n1582), .B(n1581), .Z(n446) );
  NAND U1782 ( .A(c[62]), .B(rst), .Z(n1587) );
  XNOR U1783 ( .A(n1584), .B(n1583), .Z(n1585) );
  NANDN U1784 ( .A(rst), .B(n1585), .Z(n1586) );
  NAND U1785 ( .A(n1587), .B(n1586), .Z(n447) );
  NAND U1786 ( .A(c[63]), .B(rst), .Z(n1592) );
  XOR U1787 ( .A(n1589), .B(n1588), .Z(n1590) );
  NANDN U1788 ( .A(rst), .B(n1590), .Z(n1591) );
  NAND U1789 ( .A(n1592), .B(n1591), .Z(n448) );
  NAND U1790 ( .A(c[64]), .B(rst), .Z(n1597) );
  XNOR U1791 ( .A(n1594), .B(n1593), .Z(n1595) );
  NANDN U1792 ( .A(rst), .B(n1595), .Z(n1596) );
  NAND U1793 ( .A(n1597), .B(n1596), .Z(n449) );
  NAND U1794 ( .A(c[65]), .B(rst), .Z(n1602) );
  XOR U1795 ( .A(n1599), .B(n1598), .Z(n1600) );
  NANDN U1796 ( .A(rst), .B(n1600), .Z(n1601) );
  NAND U1797 ( .A(n1602), .B(n1601), .Z(n450) );
  NAND U1798 ( .A(c[66]), .B(rst), .Z(n1607) );
  XNOR U1799 ( .A(n1604), .B(n1603), .Z(n1605) );
  NANDN U1800 ( .A(rst), .B(n1605), .Z(n1606) );
  NAND U1801 ( .A(n1607), .B(n1606), .Z(n451) );
  NAND U1802 ( .A(c[67]), .B(rst), .Z(n1612) );
  XOR U1803 ( .A(n1609), .B(n1608), .Z(n1610) );
  NANDN U1804 ( .A(rst), .B(n1610), .Z(n1611) );
  NAND U1805 ( .A(n1612), .B(n1611), .Z(n452) );
  NAND U1806 ( .A(c[68]), .B(rst), .Z(n1617) );
  XNOR U1807 ( .A(n1614), .B(n1613), .Z(n1615) );
  NANDN U1808 ( .A(rst), .B(n1615), .Z(n1616) );
  NAND U1809 ( .A(n1617), .B(n1616), .Z(n453) );
  NAND U1810 ( .A(c[69]), .B(rst), .Z(n1622) );
  XOR U1811 ( .A(n1619), .B(n1618), .Z(n1620) );
  NANDN U1812 ( .A(rst), .B(n1620), .Z(n1621) );
  NAND U1813 ( .A(n1622), .B(n1621), .Z(n454) );
  NAND U1814 ( .A(c[70]), .B(rst), .Z(n1627) );
  XNOR U1815 ( .A(n1624), .B(n1623), .Z(n1625) );
  NANDN U1816 ( .A(rst), .B(n1625), .Z(n1626) );
  NAND U1817 ( .A(n1627), .B(n1626), .Z(n455) );
  NAND U1818 ( .A(c[71]), .B(rst), .Z(n1632) );
  XOR U1819 ( .A(n1629), .B(n1628), .Z(n1630) );
  NANDN U1820 ( .A(rst), .B(n1630), .Z(n1631) );
  NAND U1821 ( .A(n1632), .B(n1631), .Z(n456) );
  NAND U1822 ( .A(c[72]), .B(rst), .Z(n1637) );
  XNOR U1823 ( .A(n1634), .B(n1633), .Z(n1635) );
  NANDN U1824 ( .A(rst), .B(n1635), .Z(n1636) );
  NAND U1825 ( .A(n1637), .B(n1636), .Z(n457) );
  NAND U1826 ( .A(c[73]), .B(rst), .Z(n1642) );
  XOR U1827 ( .A(n1639), .B(n1638), .Z(n1640) );
  NANDN U1828 ( .A(rst), .B(n1640), .Z(n1641) );
  NAND U1829 ( .A(n1642), .B(n1641), .Z(n458) );
  NAND U1830 ( .A(c[74]), .B(rst), .Z(n1647) );
  XNOR U1831 ( .A(n1644), .B(n1643), .Z(n1645) );
  NANDN U1832 ( .A(rst), .B(n1645), .Z(n1646) );
  NAND U1833 ( .A(n1647), .B(n1646), .Z(n459) );
  NAND U1834 ( .A(c[75]), .B(rst), .Z(n1652) );
  XOR U1835 ( .A(n1649), .B(n1648), .Z(n1650) );
  NANDN U1836 ( .A(rst), .B(n1650), .Z(n1651) );
  NAND U1837 ( .A(n1652), .B(n1651), .Z(n460) );
  NAND U1838 ( .A(c[76]), .B(rst), .Z(n1657) );
  XNOR U1839 ( .A(n1654), .B(n1653), .Z(n1655) );
  NANDN U1840 ( .A(rst), .B(n1655), .Z(n1656) );
  NAND U1841 ( .A(n1657), .B(n1656), .Z(n461) );
  NAND U1842 ( .A(c[77]), .B(rst), .Z(n1662) );
  XOR U1843 ( .A(n1659), .B(n1658), .Z(n1660) );
  NANDN U1844 ( .A(rst), .B(n1660), .Z(n1661) );
  NAND U1845 ( .A(n1662), .B(n1661), .Z(n462) );
  NAND U1846 ( .A(c[78]), .B(rst), .Z(n1667) );
  XNOR U1847 ( .A(n1664), .B(n1663), .Z(n1665) );
  NANDN U1848 ( .A(rst), .B(n1665), .Z(n1666) );
  NAND U1849 ( .A(n1667), .B(n1666), .Z(n463) );
  NAND U1850 ( .A(c[79]), .B(rst), .Z(n1672) );
  XOR U1851 ( .A(n1669), .B(n1668), .Z(n1670) );
  NANDN U1852 ( .A(rst), .B(n1670), .Z(n1671) );
  NAND U1853 ( .A(n1672), .B(n1671), .Z(n464) );
  NAND U1854 ( .A(c[80]), .B(rst), .Z(n1677) );
  XNOR U1855 ( .A(n1674), .B(n1673), .Z(n1675) );
  NANDN U1856 ( .A(rst), .B(n1675), .Z(n1676) );
  NAND U1857 ( .A(n1677), .B(n1676), .Z(n465) );
  NAND U1858 ( .A(c[81]), .B(rst), .Z(n1682) );
  XOR U1859 ( .A(n1679), .B(n1678), .Z(n1680) );
  NANDN U1860 ( .A(rst), .B(n1680), .Z(n1681) );
  NAND U1861 ( .A(n1682), .B(n1681), .Z(n466) );
  NAND U1862 ( .A(c[82]), .B(rst), .Z(n1687) );
  XNOR U1863 ( .A(n1684), .B(n1683), .Z(n1685) );
  NANDN U1864 ( .A(rst), .B(n1685), .Z(n1686) );
  NAND U1865 ( .A(n1687), .B(n1686), .Z(n467) );
  NAND U1866 ( .A(c[83]), .B(rst), .Z(n1692) );
  XOR U1867 ( .A(n1689), .B(n1688), .Z(n1690) );
  NANDN U1868 ( .A(rst), .B(n1690), .Z(n1691) );
  NAND U1869 ( .A(n1692), .B(n1691), .Z(n468) );
  NAND U1870 ( .A(c[84]), .B(rst), .Z(n1697) );
  XNOR U1871 ( .A(n1694), .B(n1693), .Z(n1695) );
  NANDN U1872 ( .A(rst), .B(n1695), .Z(n1696) );
  NAND U1873 ( .A(n1697), .B(n1696), .Z(n469) );
  NAND U1874 ( .A(c[85]), .B(rst), .Z(n1702) );
  XOR U1875 ( .A(n1699), .B(n1698), .Z(n1700) );
  NANDN U1876 ( .A(rst), .B(n1700), .Z(n1701) );
  NAND U1877 ( .A(n1702), .B(n1701), .Z(n470) );
  NAND U1878 ( .A(c[86]), .B(rst), .Z(n1707) );
  XNOR U1879 ( .A(n1704), .B(n1703), .Z(n1705) );
  NANDN U1880 ( .A(rst), .B(n1705), .Z(n1706) );
  NAND U1881 ( .A(n1707), .B(n1706), .Z(n471) );
  NAND U1882 ( .A(c[87]), .B(rst), .Z(n1712) );
  XOR U1883 ( .A(n1709), .B(n1708), .Z(n1710) );
  NANDN U1884 ( .A(rst), .B(n1710), .Z(n1711) );
  NAND U1885 ( .A(n1712), .B(n1711), .Z(n472) );
  NAND U1886 ( .A(c[88]), .B(rst), .Z(n1717) );
  XNOR U1887 ( .A(n1714), .B(n1713), .Z(n1715) );
  NANDN U1888 ( .A(rst), .B(n1715), .Z(n1716) );
  NAND U1889 ( .A(n1717), .B(n1716), .Z(n473) );
  NAND U1890 ( .A(c[89]), .B(rst), .Z(n1722) );
  XOR U1891 ( .A(n1719), .B(n1718), .Z(n1720) );
  NANDN U1892 ( .A(rst), .B(n1720), .Z(n1721) );
  NAND U1893 ( .A(n1722), .B(n1721), .Z(n474) );
  NAND U1894 ( .A(c[90]), .B(rst), .Z(n1727) );
  XNOR U1895 ( .A(n1724), .B(n1723), .Z(n1725) );
  NANDN U1896 ( .A(rst), .B(n1725), .Z(n1726) );
  NAND U1897 ( .A(n1727), .B(n1726), .Z(n475) );
  NAND U1898 ( .A(c[91]), .B(rst), .Z(n1732) );
  XOR U1899 ( .A(n1729), .B(n1728), .Z(n1730) );
  NANDN U1900 ( .A(rst), .B(n1730), .Z(n1731) );
  NAND U1901 ( .A(n1732), .B(n1731), .Z(n476) );
  NAND U1902 ( .A(c[92]), .B(rst), .Z(n1737) );
  XNOR U1903 ( .A(n1734), .B(n1733), .Z(n1735) );
  NANDN U1904 ( .A(rst), .B(n1735), .Z(n1736) );
  NAND U1905 ( .A(n1737), .B(n1736), .Z(n477) );
  NAND U1906 ( .A(c[93]), .B(rst), .Z(n1742) );
  XOR U1907 ( .A(n1739), .B(n1738), .Z(n1740) );
  NANDN U1908 ( .A(rst), .B(n1740), .Z(n1741) );
  NAND U1909 ( .A(n1742), .B(n1741), .Z(n478) );
  NAND U1910 ( .A(c[94]), .B(rst), .Z(n1747) );
  XNOR U1911 ( .A(n1744), .B(n1743), .Z(n1745) );
  NANDN U1912 ( .A(rst), .B(n1745), .Z(n1746) );
  NAND U1913 ( .A(n1747), .B(n1746), .Z(n479) );
  NAND U1914 ( .A(c[95]), .B(rst), .Z(n1752) );
  XOR U1915 ( .A(n1749), .B(n1748), .Z(n1750) );
  NANDN U1916 ( .A(rst), .B(n1750), .Z(n1751) );
  NAND U1917 ( .A(n1752), .B(n1751), .Z(n480) );
  NAND U1918 ( .A(c[96]), .B(rst), .Z(n1757) );
  XNOR U1919 ( .A(n1754), .B(n1753), .Z(n1755) );
  NANDN U1920 ( .A(rst), .B(n1755), .Z(n1756) );
  NAND U1921 ( .A(n1757), .B(n1756), .Z(n481) );
  NAND U1922 ( .A(c[97]), .B(rst), .Z(n1762) );
  XOR U1923 ( .A(n1759), .B(n1758), .Z(n1760) );
  NANDN U1924 ( .A(rst), .B(n1760), .Z(n1761) );
  NAND U1925 ( .A(n1762), .B(n1761), .Z(n482) );
  NAND U1926 ( .A(c[98]), .B(rst), .Z(n1767) );
  XNOR U1927 ( .A(n1764), .B(n1763), .Z(n1765) );
  NANDN U1928 ( .A(rst), .B(n1765), .Z(n1766) );
  NAND U1929 ( .A(n1767), .B(n1766), .Z(n483) );
  NAND U1930 ( .A(c[99]), .B(rst), .Z(n1772) );
  XOR U1931 ( .A(n1769), .B(n1768), .Z(n1770) );
  NANDN U1932 ( .A(rst), .B(n1770), .Z(n1771) );
  NAND U1933 ( .A(n1772), .B(n1771), .Z(n484) );
  NAND U1934 ( .A(c[100]), .B(rst), .Z(n1777) );
  XNOR U1935 ( .A(n1774), .B(n1773), .Z(n1775) );
  NANDN U1936 ( .A(rst), .B(n1775), .Z(n1776) );
  NAND U1937 ( .A(n1777), .B(n1776), .Z(n485) );
  NAND U1938 ( .A(c[101]), .B(rst), .Z(n1782) );
  XOR U1939 ( .A(n1779), .B(n1778), .Z(n1780) );
  NANDN U1940 ( .A(rst), .B(n1780), .Z(n1781) );
  NAND U1941 ( .A(n1782), .B(n1781), .Z(n486) );
  NAND U1942 ( .A(c[102]), .B(rst), .Z(n1787) );
  XNOR U1943 ( .A(n1784), .B(n1783), .Z(n1785) );
  NANDN U1944 ( .A(rst), .B(n1785), .Z(n1786) );
  NAND U1945 ( .A(n1787), .B(n1786), .Z(n487) );
  NAND U1946 ( .A(c[103]), .B(rst), .Z(n1792) );
  XOR U1947 ( .A(n1789), .B(n1788), .Z(n1790) );
  NANDN U1948 ( .A(rst), .B(n1790), .Z(n1791) );
  NAND U1949 ( .A(n1792), .B(n1791), .Z(n488) );
  NAND U1950 ( .A(c[104]), .B(rst), .Z(n1797) );
  XNOR U1951 ( .A(n1794), .B(n1793), .Z(n1795) );
  NANDN U1952 ( .A(rst), .B(n1795), .Z(n1796) );
  NAND U1953 ( .A(n1797), .B(n1796), .Z(n489) );
  NAND U1954 ( .A(c[105]), .B(rst), .Z(n1802) );
  XOR U1955 ( .A(n1799), .B(n1798), .Z(n1800) );
  NANDN U1956 ( .A(rst), .B(n1800), .Z(n1801) );
  NAND U1957 ( .A(n1802), .B(n1801), .Z(n490) );
  NAND U1958 ( .A(c[106]), .B(rst), .Z(n1807) );
  XNOR U1959 ( .A(n1804), .B(n1803), .Z(n1805) );
  NANDN U1960 ( .A(rst), .B(n1805), .Z(n1806) );
  NAND U1961 ( .A(n1807), .B(n1806), .Z(n491) );
  NAND U1962 ( .A(c[107]), .B(rst), .Z(n1812) );
  XOR U1963 ( .A(n1809), .B(n1808), .Z(n1810) );
  NANDN U1964 ( .A(rst), .B(n1810), .Z(n1811) );
  NAND U1965 ( .A(n1812), .B(n1811), .Z(n492) );
  NAND U1966 ( .A(c[108]), .B(rst), .Z(n1817) );
  XNOR U1967 ( .A(n1814), .B(n1813), .Z(n1815) );
  NANDN U1968 ( .A(rst), .B(n1815), .Z(n1816) );
  NAND U1969 ( .A(n1817), .B(n1816), .Z(n493) );
  NAND U1970 ( .A(c[109]), .B(rst), .Z(n1822) );
  XOR U1971 ( .A(n1819), .B(n1818), .Z(n1820) );
  NANDN U1972 ( .A(rst), .B(n1820), .Z(n1821) );
  NAND U1973 ( .A(n1822), .B(n1821), .Z(n494) );
  NAND U1974 ( .A(c[110]), .B(rst), .Z(n1827) );
  XNOR U1975 ( .A(n1824), .B(n1823), .Z(n1825) );
  NANDN U1976 ( .A(rst), .B(n1825), .Z(n1826) );
  NAND U1977 ( .A(n1827), .B(n1826), .Z(n495) );
  NAND U1978 ( .A(c[111]), .B(rst), .Z(n1832) );
  XOR U1979 ( .A(n1829), .B(n1828), .Z(n1830) );
  NANDN U1980 ( .A(rst), .B(n1830), .Z(n1831) );
  NAND U1981 ( .A(n1832), .B(n1831), .Z(n496) );
  NAND U1982 ( .A(c[112]), .B(rst), .Z(n1837) );
  XNOR U1983 ( .A(n1834), .B(n1833), .Z(n1835) );
  NANDN U1984 ( .A(rst), .B(n1835), .Z(n1836) );
  NAND U1985 ( .A(n1837), .B(n1836), .Z(n497) );
  NAND U1986 ( .A(c[113]), .B(rst), .Z(n1842) );
  XOR U1987 ( .A(n1839), .B(n1838), .Z(n1840) );
  NANDN U1988 ( .A(rst), .B(n1840), .Z(n1841) );
  NAND U1989 ( .A(n1842), .B(n1841), .Z(n498) );
  NAND U1990 ( .A(c[114]), .B(rst), .Z(n1847) );
  XNOR U1991 ( .A(n1844), .B(n1843), .Z(n1845) );
  NANDN U1992 ( .A(rst), .B(n1845), .Z(n1846) );
  NAND U1993 ( .A(n1847), .B(n1846), .Z(n499) );
  NAND U1994 ( .A(c[115]), .B(rst), .Z(n1852) );
  XOR U1995 ( .A(n1849), .B(n1848), .Z(n1850) );
  NANDN U1996 ( .A(rst), .B(n1850), .Z(n1851) );
  NAND U1997 ( .A(n1852), .B(n1851), .Z(n500) );
  NAND U1998 ( .A(c[116]), .B(rst), .Z(n1857) );
  XNOR U1999 ( .A(n1854), .B(n1853), .Z(n1855) );
  NANDN U2000 ( .A(rst), .B(n1855), .Z(n1856) );
  NAND U2001 ( .A(n1857), .B(n1856), .Z(n501) );
  NAND U2002 ( .A(c[117]), .B(rst), .Z(n1862) );
  XOR U2003 ( .A(n1859), .B(n1858), .Z(n1860) );
  NANDN U2004 ( .A(rst), .B(n1860), .Z(n1861) );
  NAND U2005 ( .A(n1862), .B(n1861), .Z(n502) );
  NAND U2006 ( .A(c[118]), .B(rst), .Z(n1867) );
  XNOR U2007 ( .A(n1864), .B(n1863), .Z(n1865) );
  NANDN U2008 ( .A(rst), .B(n1865), .Z(n1866) );
  NAND U2009 ( .A(n1867), .B(n1866), .Z(n503) );
  NAND U2010 ( .A(c[119]), .B(rst), .Z(n1872) );
  XOR U2011 ( .A(n1869), .B(n1868), .Z(n1870) );
  NANDN U2012 ( .A(rst), .B(n1870), .Z(n1871) );
  NAND U2013 ( .A(n1872), .B(n1871), .Z(n504) );
  NAND U2014 ( .A(c[120]), .B(rst), .Z(n1877) );
  XNOR U2015 ( .A(n1874), .B(n1873), .Z(n1875) );
  NANDN U2016 ( .A(rst), .B(n1875), .Z(n1876) );
  NAND U2017 ( .A(n1877), .B(n1876), .Z(n505) );
  NAND U2018 ( .A(c[121]), .B(rst), .Z(n1882) );
  XOR U2019 ( .A(n1879), .B(n1878), .Z(n1880) );
  NANDN U2020 ( .A(rst), .B(n1880), .Z(n1881) );
  NAND U2021 ( .A(n1882), .B(n1881), .Z(n506) );
  NAND U2022 ( .A(c[122]), .B(rst), .Z(n1887) );
  XNOR U2023 ( .A(n1884), .B(n1883), .Z(n1885) );
  NANDN U2024 ( .A(rst), .B(n1885), .Z(n1886) );
  NAND U2025 ( .A(n1887), .B(n1886), .Z(n507) );
  NAND U2026 ( .A(c[123]), .B(rst), .Z(n1892) );
  XOR U2027 ( .A(n1889), .B(n1888), .Z(n1890) );
  NANDN U2028 ( .A(rst), .B(n1890), .Z(n1891) );
  NAND U2029 ( .A(n1892), .B(n1891), .Z(n508) );
  NAND U2030 ( .A(c[124]), .B(rst), .Z(n1897) );
  XNOR U2031 ( .A(n1894), .B(n1893), .Z(n1895) );
  NANDN U2032 ( .A(rst), .B(n1895), .Z(n1896) );
  NAND U2033 ( .A(n1897), .B(n1896), .Z(n509) );
  NAND U2034 ( .A(c[125]), .B(rst), .Z(n1902) );
  XOR U2035 ( .A(n1899), .B(n1898), .Z(n1900) );
  NANDN U2036 ( .A(rst), .B(n1900), .Z(n1901) );
  NAND U2037 ( .A(n1902), .B(n1901), .Z(n510) );
  NAND U2038 ( .A(c[126]), .B(rst), .Z(n1907) );
  XNOR U2039 ( .A(n1904), .B(n1903), .Z(n1905) );
  NANDN U2040 ( .A(rst), .B(n1905), .Z(n1906) );
  NAND U2041 ( .A(n1907), .B(n1906), .Z(n511) );
  NAND U2042 ( .A(c[127]), .B(rst), .Z(n1912) );
  XOR U2043 ( .A(n1909), .B(n1908), .Z(n1910) );
  NANDN U2044 ( .A(rst), .B(n1910), .Z(n1911) );
  NAND U2045 ( .A(n1912), .B(n1911), .Z(n512) );
endmodule

